module basic_1500_15000_2000_5_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_631,In_1383);
nor U1 (N_1,In_1335,In_627);
and U2 (N_2,In_1426,In_678);
or U3 (N_3,In_185,In_816);
or U4 (N_4,In_665,In_593);
nor U5 (N_5,In_827,In_1217);
nor U6 (N_6,In_1241,In_757);
or U7 (N_7,In_1023,In_856);
and U8 (N_8,In_194,In_895);
or U9 (N_9,In_51,In_1171);
nor U10 (N_10,In_57,In_971);
nand U11 (N_11,In_523,In_1083);
nand U12 (N_12,In_739,In_1100);
or U13 (N_13,In_78,In_573);
nand U14 (N_14,In_464,In_606);
or U15 (N_15,In_1040,In_369);
nand U16 (N_16,In_1461,In_1416);
and U17 (N_17,In_802,In_90);
nand U18 (N_18,In_134,In_1033);
nand U19 (N_19,In_1482,In_1251);
and U20 (N_20,In_1265,In_970);
nand U21 (N_21,In_370,In_1065);
or U22 (N_22,In_311,In_434);
or U23 (N_23,In_43,In_1285);
nand U24 (N_24,In_611,In_1225);
or U25 (N_25,In_1364,In_1196);
and U26 (N_26,In_1096,In_422);
and U27 (N_27,In_406,In_985);
nand U28 (N_28,In_968,In_1245);
and U29 (N_29,In_1288,In_474);
and U30 (N_30,In_495,In_753);
nand U31 (N_31,In_1291,In_694);
nand U32 (N_32,In_663,In_1256);
and U33 (N_33,In_522,In_377);
or U34 (N_34,In_1290,In_513);
nor U35 (N_35,In_1376,In_1191);
nor U36 (N_36,In_438,In_295);
and U37 (N_37,In_969,In_1438);
nand U38 (N_38,In_661,In_813);
and U39 (N_39,In_1200,In_17);
nor U40 (N_40,In_845,In_430);
nor U41 (N_41,In_1456,In_419);
nor U42 (N_42,In_65,In_1323);
and U43 (N_43,In_1113,In_404);
nand U44 (N_44,In_756,In_817);
nand U45 (N_45,In_1237,In_1);
nor U46 (N_46,In_1247,In_1347);
or U47 (N_47,In_1390,In_1109);
xor U48 (N_48,In_149,In_892);
nor U49 (N_49,In_153,In_922);
nor U50 (N_50,In_75,In_1341);
nor U51 (N_51,In_893,In_614);
or U52 (N_52,In_159,In_583);
nor U53 (N_53,In_30,In_318);
and U54 (N_54,In_374,In_931);
and U55 (N_55,In_32,In_420);
nor U56 (N_56,In_619,In_274);
nor U57 (N_57,In_1136,In_446);
nand U58 (N_58,In_1402,In_300);
nor U59 (N_59,In_1302,In_632);
or U60 (N_60,In_339,In_166);
nor U61 (N_61,In_834,In_996);
and U62 (N_62,In_643,In_1398);
nand U63 (N_63,In_267,In_579);
and U64 (N_64,In_1469,In_447);
nand U65 (N_65,In_516,In_1355);
or U66 (N_66,In_784,In_1278);
nor U67 (N_67,In_467,In_239);
nor U68 (N_68,In_995,In_225);
or U69 (N_69,In_1253,In_29);
nor U70 (N_70,In_454,In_1007);
nor U71 (N_71,In_1373,In_992);
or U72 (N_72,In_1326,In_854);
nor U73 (N_73,In_72,In_515);
or U74 (N_74,In_183,In_1233);
or U75 (N_75,In_825,In_1216);
or U76 (N_76,In_1316,In_695);
nand U77 (N_77,In_914,In_1235);
and U78 (N_78,In_23,In_308);
nand U79 (N_79,In_1126,In_538);
nand U80 (N_80,In_729,In_1258);
or U81 (N_81,In_286,In_1473);
xnor U82 (N_82,In_62,In_820);
xor U83 (N_83,In_868,In_1173);
nand U84 (N_84,In_533,In_258);
and U85 (N_85,In_1440,In_655);
nor U86 (N_86,In_63,In_246);
nor U87 (N_87,In_1344,In_340);
nand U88 (N_88,In_1465,In_459);
nand U89 (N_89,In_1429,In_261);
and U90 (N_90,In_918,In_1379);
nand U91 (N_91,In_1084,In_243);
nor U92 (N_92,In_659,In_11);
or U93 (N_93,In_810,In_206);
nand U94 (N_94,In_1161,In_81);
nand U95 (N_95,In_38,In_1218);
nand U96 (N_96,In_507,In_751);
nor U97 (N_97,In_129,In_1139);
nor U98 (N_98,In_385,In_731);
and U99 (N_99,In_1018,In_469);
or U100 (N_100,In_1066,In_955);
or U101 (N_101,In_1399,In_691);
nand U102 (N_102,In_1181,In_26);
nand U103 (N_103,In_237,In_1377);
nand U104 (N_104,In_965,In_1006);
and U105 (N_105,In_587,In_875);
xor U106 (N_106,In_889,In_765);
or U107 (N_107,In_463,In_1491);
nand U108 (N_108,In_759,In_602);
nand U109 (N_109,In_122,In_1021);
and U110 (N_110,In_491,In_241);
nand U111 (N_111,In_64,In_843);
nand U112 (N_112,In_131,In_577);
and U113 (N_113,In_568,In_209);
nand U114 (N_114,In_508,In_371);
and U115 (N_115,In_74,In_618);
or U116 (N_116,In_52,In_972);
and U117 (N_117,In_1219,In_716);
nand U118 (N_118,In_857,In_1299);
nor U119 (N_119,In_1063,In_444);
and U120 (N_120,In_1035,In_326);
and U121 (N_121,In_1486,In_228);
nor U122 (N_122,In_73,In_737);
nor U123 (N_123,In_544,In_141);
nor U124 (N_124,In_1481,In_1274);
nor U125 (N_125,In_1411,In_233);
and U126 (N_126,In_806,In_599);
and U127 (N_127,In_40,In_624);
nor U128 (N_128,In_104,In_1490);
and U129 (N_129,In_1356,In_324);
nor U130 (N_130,In_1188,In_499);
and U131 (N_131,In_1273,In_645);
and U132 (N_132,In_160,In_672);
nor U133 (N_133,In_204,In_863);
and U134 (N_134,In_407,In_1127);
nor U135 (N_135,In_9,In_270);
or U136 (N_136,In_890,In_539);
and U137 (N_137,In_94,In_750);
nand U138 (N_138,In_709,In_60);
nor U139 (N_139,In_708,In_1480);
nand U140 (N_140,In_200,In_1050);
nor U141 (N_141,In_1076,In_1346);
nor U142 (N_142,In_1037,In_788);
or U143 (N_143,In_1002,In_487);
nor U144 (N_144,In_993,In_470);
xor U145 (N_145,In_651,In_835);
nor U146 (N_146,In_54,In_1110);
nand U147 (N_147,In_83,In_220);
nor U148 (N_148,In_964,In_829);
nor U149 (N_149,In_99,In_1078);
and U150 (N_150,In_217,In_101);
nand U151 (N_151,In_908,In_502);
or U152 (N_152,In_435,In_903);
or U153 (N_153,In_238,In_126);
or U154 (N_154,In_1085,In_667);
nand U155 (N_155,In_1387,In_178);
and U156 (N_156,In_1466,In_634);
nand U157 (N_157,In_1406,In_550);
nor U158 (N_158,In_15,In_654);
nand U159 (N_159,In_685,In_1361);
nor U160 (N_160,In_1107,In_836);
nand U161 (N_161,In_831,In_608);
nand U162 (N_162,In_506,In_296);
or U163 (N_163,In_1255,In_367);
xor U164 (N_164,In_18,In_984);
nand U165 (N_165,In_668,In_1052);
or U166 (N_166,In_58,In_1182);
nand U167 (N_167,In_749,In_1305);
nor U168 (N_168,In_31,In_97);
or U169 (N_169,In_773,In_1234);
nand U170 (N_170,In_1282,In_986);
or U171 (N_171,In_403,In_1322);
or U172 (N_172,In_457,In_325);
and U173 (N_173,In_222,In_763);
and U174 (N_174,In_1008,In_1250);
or U175 (N_175,In_1163,In_548);
and U176 (N_176,In_1178,In_881);
nand U177 (N_177,In_1280,In_113);
or U178 (N_178,In_1319,In_235);
or U179 (N_179,In_743,In_924);
nor U180 (N_180,In_425,In_537);
and U181 (N_181,In_1381,In_1343);
nand U182 (N_182,In_219,In_299);
and U183 (N_183,In_1444,In_120);
nor U184 (N_184,In_1362,In_1211);
nor U185 (N_185,In_738,In_1039);
and U186 (N_186,In_6,In_285);
nor U187 (N_187,In_357,In_617);
nor U188 (N_188,In_226,In_1333);
and U189 (N_189,In_382,In_264);
nor U190 (N_190,In_1276,In_1164);
xor U191 (N_191,In_1293,In_1449);
or U192 (N_192,In_27,In_501);
nand U193 (N_193,In_1442,In_1430);
or U194 (N_194,In_56,In_1358);
xor U195 (N_195,In_952,In_331);
and U196 (N_196,In_215,In_398);
and U197 (N_197,In_1423,In_509);
nand U198 (N_198,In_555,In_1170);
nor U199 (N_199,In_1014,In_347);
and U200 (N_200,In_201,In_683);
and U201 (N_201,In_884,In_41);
nor U202 (N_202,In_115,In_973);
nand U203 (N_203,In_327,In_861);
and U204 (N_204,In_163,In_888);
and U205 (N_205,In_1378,In_704);
nor U206 (N_206,In_188,In_473);
or U207 (N_207,In_77,In_894);
nand U208 (N_208,In_553,In_630);
nor U209 (N_209,In_1297,In_42);
nor U210 (N_210,In_88,In_1311);
nor U211 (N_211,In_623,In_298);
xnor U212 (N_212,In_1104,In_152);
or U213 (N_213,In_864,In_1206);
nor U214 (N_214,In_556,In_811);
and U215 (N_215,In_291,In_859);
or U216 (N_216,In_679,In_1254);
or U217 (N_217,In_316,In_850);
or U218 (N_218,In_1156,In_823);
or U219 (N_219,In_1227,In_1261);
or U220 (N_220,In_517,In_728);
nand U221 (N_221,In_1309,In_1318);
nand U222 (N_222,In_313,In_1000);
nor U223 (N_223,In_794,In_361);
and U224 (N_224,In_91,In_28);
nor U225 (N_225,In_334,In_1408);
or U226 (N_226,In_584,In_1207);
nand U227 (N_227,In_703,In_658);
and U228 (N_228,In_229,In_448);
or U229 (N_229,In_1352,In_1422);
nand U230 (N_230,In_1393,In_1244);
or U231 (N_231,In_391,In_36);
and U232 (N_232,In_724,In_748);
nor U233 (N_233,In_629,In_1374);
nand U234 (N_234,In_1224,In_1435);
nor U235 (N_235,In_1419,In_976);
and U236 (N_236,In_1150,In_140);
or U237 (N_237,In_828,In_1412);
and U238 (N_238,In_1354,In_789);
and U239 (N_239,In_1238,In_365);
or U240 (N_240,In_1324,In_575);
nor U241 (N_241,In_1329,In_1044);
and U242 (N_242,In_1199,In_1303);
nor U243 (N_243,In_730,In_108);
nor U244 (N_244,In_991,In_1151);
or U245 (N_245,In_1146,In_839);
nor U246 (N_246,In_671,In_89);
nand U247 (N_247,In_518,In_176);
and U248 (N_248,In_844,In_946);
and U249 (N_249,In_769,In_1108);
or U250 (N_250,In_701,In_597);
and U251 (N_251,In_589,In_1048);
xor U252 (N_252,In_528,In_307);
xor U253 (N_253,In_150,In_718);
or U254 (N_254,In_1272,In_1407);
nand U255 (N_255,In_1013,In_997);
nor U256 (N_256,In_352,In_151);
or U257 (N_257,In_1116,In_277);
nand U258 (N_258,In_330,In_1057);
nor U259 (N_259,In_1089,In_375);
xnor U260 (N_260,In_781,In_251);
and U261 (N_261,In_111,In_208);
and U262 (N_262,In_851,In_755);
xnor U263 (N_263,In_356,In_1101);
nor U264 (N_264,In_1472,In_275);
or U265 (N_265,In_14,In_37);
nor U266 (N_266,In_390,In_1198);
nand U267 (N_267,In_840,In_1121);
or U268 (N_268,In_1162,In_1431);
xnor U269 (N_269,In_492,In_412);
and U270 (N_270,In_343,In_527);
nor U271 (N_271,In_943,In_1103);
and U272 (N_272,In_493,In_653);
xnor U273 (N_273,In_462,In_768);
and U274 (N_274,In_1301,In_429);
or U275 (N_275,In_164,In_196);
nand U276 (N_276,In_342,In_1079);
nand U277 (N_277,In_269,In_842);
nor U278 (N_278,In_929,In_388);
or U279 (N_279,In_1143,In_1372);
nand U280 (N_280,In_39,In_1118);
or U281 (N_281,In_1165,In_1215);
and U282 (N_282,In_80,In_1029);
nor U283 (N_283,In_1401,In_292);
or U284 (N_284,In_96,In_1231);
or U285 (N_285,In_721,In_248);
or U286 (N_286,In_1180,In_564);
nor U287 (N_287,In_284,In_921);
nor U288 (N_288,In_1155,In_916);
and U289 (N_289,In_345,In_882);
xor U290 (N_290,In_871,In_1495);
or U291 (N_291,In_268,In_912);
or U292 (N_292,In_783,In_1175);
nand U293 (N_293,In_1203,In_1294);
nand U294 (N_294,In_127,In_621);
or U295 (N_295,In_562,In_471);
nand U296 (N_296,In_1153,In_287);
nor U297 (N_297,In_428,In_353);
nand U298 (N_298,In_1289,In_67);
nor U299 (N_299,In_93,In_932);
nor U300 (N_300,In_1296,In_4);
or U301 (N_301,In_1051,In_319);
or U302 (N_302,In_1034,In_1192);
nand U303 (N_303,In_620,In_951);
nor U304 (N_304,In_959,In_503);
or U305 (N_305,In_1026,In_417);
or U306 (N_306,In_869,In_725);
and U307 (N_307,In_578,In_116);
or U308 (N_308,In_936,In_937);
or U309 (N_309,In_732,In_221);
or U310 (N_310,In_880,In_572);
and U311 (N_311,In_705,In_966);
or U312 (N_312,In_994,In_1221);
nor U313 (N_313,In_637,In_213);
nand U314 (N_314,In_1005,In_472);
nand U315 (N_315,In_689,In_690);
nand U316 (N_316,In_1371,In_478);
nand U317 (N_317,In_1471,In_1365);
nand U318 (N_318,In_273,In_254);
xnor U319 (N_319,In_379,In_1312);
nand U320 (N_320,In_558,In_1105);
and U321 (N_321,In_1142,In_436);
and U322 (N_322,In_1112,In_1072);
nor U323 (N_323,In_230,In_867);
or U324 (N_324,In_787,In_1117);
or U325 (N_325,In_443,In_144);
and U326 (N_326,In_139,In_551);
or U327 (N_327,In_698,In_1396);
and U328 (N_328,In_913,In_1269);
or U329 (N_329,In_402,In_1194);
or U330 (N_330,In_494,In_1457);
nand U331 (N_331,In_734,In_950);
or U332 (N_332,In_198,In_1030);
nor U333 (N_333,In_543,In_639);
or U334 (N_334,In_920,In_1487);
or U335 (N_335,In_649,In_1093);
and U336 (N_336,In_1332,In_423);
nor U337 (N_337,In_1214,In_1141);
or U338 (N_338,In_190,In_1060);
or U339 (N_339,In_796,In_758);
and U340 (N_340,In_511,In_68);
nor U341 (N_341,In_1493,In_455);
nand U342 (N_342,In_271,In_1123);
and U343 (N_343,In_944,In_949);
nand U344 (N_344,In_184,In_1268);
nand U345 (N_345,In_574,In_1330);
nand U346 (N_346,In_186,In_272);
and U347 (N_347,In_1425,In_779);
xnor U348 (N_348,In_1054,In_540);
nand U349 (N_349,In_745,In_767);
nor U350 (N_350,In_673,In_1357);
and U351 (N_351,In_1334,In_899);
nor U352 (N_352,In_1190,In_1031);
and U353 (N_353,In_309,In_1152);
and U354 (N_354,In_580,In_211);
nand U355 (N_355,In_1331,In_329);
nor U356 (N_356,In_468,In_592);
nor U357 (N_357,In_322,In_317);
and U358 (N_358,In_987,In_498);
or U359 (N_359,In_337,In_328);
nor U360 (N_360,In_1080,In_1479);
and U361 (N_361,In_1366,In_107);
xnor U362 (N_362,In_740,In_216);
and U363 (N_363,In_625,In_245);
and U364 (N_364,In_1284,In_87);
and U365 (N_365,In_85,In_1147);
nand U366 (N_366,In_1277,In_69);
or U367 (N_367,In_1160,In_250);
nand U368 (N_368,In_911,In_302);
or U369 (N_369,In_1228,In_263);
nand U370 (N_370,In_699,In_961);
or U371 (N_371,In_376,In_764);
or U372 (N_372,In_978,In_189);
nor U373 (N_373,In_642,In_1345);
or U374 (N_374,In_1025,In_900);
nand U375 (N_375,In_392,In_977);
and U376 (N_376,In_8,In_1375);
nand U377 (N_377,In_1022,In_855);
or U378 (N_378,In_803,In_1315);
or U379 (N_379,In_321,In_124);
and U380 (N_380,In_338,In_335);
nand U381 (N_381,In_804,In_290);
or U382 (N_382,In_866,In_1092);
nand U383 (N_383,In_191,In_1226);
or U384 (N_384,In_680,In_383);
nand U385 (N_385,In_1483,In_179);
and U386 (N_386,In_110,In_956);
nand U387 (N_387,In_635,In_297);
xnor U388 (N_388,In_82,In_336);
nor U389 (N_389,In_1154,In_891);
or U390 (N_390,In_1458,In_1240);
or U391 (N_391,In_860,In_1003);
nand U392 (N_392,In_1132,In_761);
nand U393 (N_393,In_1016,In_465);
nor U394 (N_394,In_760,In_5);
or U395 (N_395,In_1414,In_306);
and U396 (N_396,In_848,In_524);
nand U397 (N_397,In_1140,In_1115);
nor U398 (N_398,In_933,In_195);
and U399 (N_399,In_368,In_1403);
nor U400 (N_400,In_982,In_16);
and U401 (N_401,In_925,In_1270);
and U402 (N_402,In_847,In_1494);
and U403 (N_403,In_1232,In_741);
nand U404 (N_404,In_1447,In_628);
and U405 (N_405,In_214,In_904);
nor U406 (N_406,In_10,In_289);
xnor U407 (N_407,In_320,In_853);
or U408 (N_408,In_117,In_766);
nand U409 (N_409,In_1236,In_693);
nand U410 (N_410,In_1338,In_826);
or U411 (N_411,In_874,In_181);
or U412 (N_412,In_410,In_514);
nor U413 (N_413,In_646,In_1070);
nor U414 (N_414,In_421,In_838);
nand U415 (N_415,In_280,In_1073);
or U416 (N_416,In_175,In_870);
and U417 (N_417,In_143,In_1114);
nand U418 (N_418,In_118,In_983);
and U419 (N_419,In_939,In_1300);
nand U420 (N_420,In_165,In_736);
and U421 (N_421,In_1004,In_2);
nor U422 (N_422,In_1367,In_1159);
nor U423 (N_423,In_610,In_1202);
nand U424 (N_424,In_591,In_598);
nor U425 (N_425,In_84,In_301);
nand U426 (N_426,In_169,In_1340);
nand U427 (N_427,In_1012,In_341);
and U428 (N_428,In_452,In_1463);
or U429 (N_429,In_824,In_1488);
or U430 (N_430,In_293,In_1475);
nand U431 (N_431,In_706,In_461);
nor U432 (N_432,In_657,In_947);
or U433 (N_433,In_581,In_1197);
or U434 (N_434,In_1454,In_24);
or U435 (N_435,In_535,In_1125);
nor U436 (N_436,In_354,In_1271);
and U437 (N_437,In_771,In_1418);
or U438 (N_438,In_541,In_413);
or U439 (N_439,In_333,In_1468);
or U440 (N_440,In_224,In_415);
nand U441 (N_441,In_519,In_1389);
nor U442 (N_442,In_106,In_401);
nor U443 (N_443,In_25,In_565);
or U444 (N_444,In_1336,In_1496);
and U445 (N_445,In_1097,In_265);
and U446 (N_446,In_227,In_1353);
nor U447 (N_447,In_1424,In_381);
xor U448 (N_448,In_1395,In_1460);
nand U449 (N_449,In_1497,In_61);
and U450 (N_450,In_1212,In_1055);
nand U451 (N_451,In_1138,In_133);
or U452 (N_452,In_373,In_879);
nor U453 (N_453,In_386,In_79);
xnor U454 (N_454,In_752,In_7);
and U455 (N_455,In_1452,In_358);
and U456 (N_456,In_887,In_442);
or U457 (N_457,In_930,In_362);
nand U458 (N_458,In_50,In_147);
nor U459 (N_459,In_1492,In_719);
or U460 (N_460,In_427,In_1038);
and U461 (N_461,In_1009,In_247);
nand U462 (N_462,In_666,In_98);
or U463 (N_463,In_798,In_782);
and U464 (N_464,In_33,In_726);
nand U465 (N_465,In_1091,In_1045);
xor U466 (N_466,In_1246,In_86);
nor U467 (N_467,In_545,In_232);
or U468 (N_468,In_1020,In_1382);
nor U469 (N_469,In_1130,In_431);
or U470 (N_470,In_44,In_1281);
or U471 (N_471,In_1075,In_1019);
nor U472 (N_472,In_554,In_510);
nor U473 (N_473,In_1094,In_1032);
and U474 (N_474,In_1386,In_1448);
or U475 (N_475,In_1043,In_563);
or U476 (N_476,In_138,In_1350);
and U477 (N_477,In_1432,In_1413);
nor U478 (N_478,In_418,In_234);
nand U479 (N_479,In_1176,In_648);
or U480 (N_480,In_1230,In_1433);
and U481 (N_481,In_915,In_445);
nand U482 (N_482,In_426,In_1133);
and U483 (N_483,In_662,In_529);
and U484 (N_484,In_1428,In_146);
nor U485 (N_485,In_549,In_348);
nand U486 (N_486,In_1462,In_1208);
nand U487 (N_487,In_720,In_256);
or U488 (N_488,In_962,In_490);
xnor U489 (N_489,In_136,In_1348);
or U490 (N_490,In_450,In_1455);
nor U491 (N_491,In_830,In_772);
nand U492 (N_492,In_832,In_1028);
or U493 (N_493,In_479,In_1252);
or U494 (N_494,In_512,In_1360);
and U495 (N_495,In_1242,In_92);
nand U496 (N_496,In_387,In_1388);
nand U497 (N_497,In_197,In_652);
nor U498 (N_498,In_1243,In_873);
nand U499 (N_499,In_70,In_546);
nand U500 (N_500,In_775,In_260);
and U501 (N_501,In_1087,In_733);
and U502 (N_502,In_1131,In_66);
nor U503 (N_503,In_762,In_609);
and U504 (N_504,In_1437,In_1148);
and U505 (N_505,In_744,In_1024);
and U506 (N_506,In_1351,In_980);
or U507 (N_507,In_346,In_1047);
xor U508 (N_508,In_440,In_650);
nor U509 (N_509,In_1223,In_561);
nor U510 (N_510,In_876,In_409);
nand U511 (N_511,In_1405,In_926);
nor U512 (N_512,In_47,In_483);
nand U513 (N_513,In_885,In_1174);
and U514 (N_514,In_821,In_156);
nand U515 (N_515,In_1400,In_1128);
or U516 (N_516,In_102,In_1077);
nand U517 (N_517,In_252,In_253);
or U518 (N_518,In_158,In_696);
or U519 (N_519,In_1177,In_180);
or U520 (N_520,In_281,In_534);
xor U521 (N_521,In_571,In_531);
nand U522 (N_522,In_49,In_485);
or U523 (N_523,In_596,In_1446);
nor U524 (N_524,In_162,In_525);
xnor U525 (N_525,In_1213,In_670);
nor U526 (N_526,In_998,In_109);
and U527 (N_527,In_323,In_960);
and U528 (N_528,In_1106,In_1384);
and U529 (N_529,In_1068,In_1453);
nand U530 (N_530,In_865,In_1187);
and U531 (N_531,In_594,In_458);
nor U532 (N_532,In_132,In_394);
nand U533 (N_533,In_95,In_148);
or U534 (N_534,In_590,In_818);
nand U535 (N_535,In_858,In_948);
nor U536 (N_536,In_456,In_199);
or U537 (N_537,In_1036,In_717);
and U538 (N_538,In_355,In_310);
and U539 (N_539,In_1179,In_841);
or U540 (N_540,In_205,In_928);
and U541 (N_541,In_774,In_1267);
nand U542 (N_542,In_727,In_1441);
nor U543 (N_543,In_276,In_242);
and U544 (N_544,In_849,In_938);
or U545 (N_545,In_877,In_942);
nor U546 (N_546,In_974,In_359);
nor U547 (N_547,In_1307,In_1168);
or U548 (N_548,In_552,In_786);
xnor U549 (N_549,In_1314,In_907);
xnor U550 (N_550,In_0,In_1010);
nor U551 (N_551,In_21,In_570);
and U552 (N_552,In_350,In_795);
nand U553 (N_553,In_807,In_906);
nand U554 (N_554,In_257,In_1157);
and U555 (N_555,In_697,In_793);
nand U556 (N_556,In_1337,In_747);
and U557 (N_557,In_1011,In_1485);
nor U558 (N_558,In_735,In_675);
nand U559 (N_559,In_1443,In_1474);
nor U560 (N_560,In_656,In_441);
and U561 (N_561,In_792,In_1263);
nand U562 (N_562,In_723,In_278);
or U563 (N_563,In_799,In_453);
nand U564 (N_564,In_1484,In_480);
nand U565 (N_565,In_360,In_687);
nor U566 (N_566,In_1415,In_1086);
or U567 (N_567,In_192,In_1209);
nor U568 (N_568,In_1279,In_1464);
nand U569 (N_569,In_1229,In_380);
nor U570 (N_570,In_1184,In_640);
and U571 (N_571,In_1102,In_615);
and U572 (N_572,In_114,In_218);
nand U573 (N_573,In_710,In_1321);
and U574 (N_574,In_3,In_677);
nor U575 (N_575,In_1193,In_770);
nor U576 (N_576,In_332,In_161);
nor U577 (N_577,In_1467,In_477);
nor U578 (N_578,In_400,In_722);
or U579 (N_579,In_259,In_520);
or U580 (N_580,In_603,In_975);
nand U581 (N_581,In_1262,In_536);
nor U582 (N_582,In_1222,In_569);
and U583 (N_583,In_702,In_935);
or U584 (N_584,In_351,In_344);
or U585 (N_585,In_288,In_203);
and U586 (N_586,In_1477,In_626);
nor U587 (N_587,In_1264,In_588);
or U588 (N_588,In_76,In_963);
nor U589 (N_589,In_71,In_1489);
and U590 (N_590,In_1186,In_1498);
and U591 (N_591,In_530,In_812);
nor U592 (N_592,In_940,In_1298);
nand U593 (N_593,In_1205,In_210);
nor U594 (N_594,In_638,In_754);
nand U595 (N_595,In_1328,In_954);
nor U596 (N_596,In_372,In_231);
and U597 (N_597,In_567,In_837);
and U598 (N_598,In_155,In_1292);
nor U599 (N_599,In_130,In_560);
and U600 (N_600,In_945,In_557);
or U601 (N_601,In_283,In_294);
nand U602 (N_602,In_898,In_1137);
nand U603 (N_603,In_22,In_776);
or U604 (N_604,In_305,In_1067);
nand U605 (N_605,In_1049,In_1074);
nor U606 (N_606,In_941,In_778);
nand U607 (N_607,In_100,In_59);
nand U608 (N_608,In_1410,In_187);
nand U609 (N_609,In_112,In_304);
xor U610 (N_610,In_366,In_700);
or U611 (N_611,In_173,In_157);
nand U612 (N_612,In_1027,In_633);
and U613 (N_613,In_714,In_1082);
nand U614 (N_614,In_746,In_1476);
and U615 (N_615,In_1041,In_636);
or U616 (N_616,In_1172,In_1239);
nand U617 (N_617,In_674,In_170);
nand U618 (N_618,In_1062,In_585);
and U619 (N_619,In_896,In_497);
and U620 (N_620,In_1380,In_886);
or U621 (N_621,In_128,In_505);
and U622 (N_622,In_466,In_1166);
and U623 (N_623,In_902,In_1042);
and U624 (N_624,In_1451,In_432);
nor U625 (N_625,In_1445,In_154);
and U626 (N_626,In_125,In_262);
xor U627 (N_627,In_999,In_1342);
nand U628 (N_628,In_910,In_616);
nand U629 (N_629,In_780,In_193);
nor U630 (N_630,In_1427,In_282);
nor U631 (N_631,In_814,In_612);
xnor U632 (N_632,In_1450,In_364);
nand U633 (N_633,In_664,In_1306);
nor U634 (N_634,In_207,In_411);
nand U635 (N_635,In_715,In_1120);
xnor U636 (N_636,In_488,In_1088);
nand U637 (N_637,In_19,In_55);
or U638 (N_638,In_1210,In_681);
nand U639 (N_639,In_486,In_405);
and U640 (N_640,In_979,In_53);
nor U641 (N_641,In_526,In_500);
nand U642 (N_642,In_1095,In_121);
and U643 (N_643,In_1061,In_439);
nor U644 (N_644,In_713,In_1417);
or U645 (N_645,In_1325,In_660);
and U646 (N_646,In_927,In_46);
and U647 (N_647,In_312,In_1169);
and U648 (N_648,In_396,In_669);
or U649 (N_649,In_363,In_1368);
nand U650 (N_650,In_800,In_1220);
and U651 (N_651,In_601,In_1283);
and U652 (N_652,In_711,In_1059);
or U653 (N_653,In_1359,In_958);
nand U654 (N_654,In_1201,In_142);
or U655 (N_655,In_647,In_989);
nor U656 (N_656,In_437,In_909);
nand U657 (N_657,In_967,In_1391);
and U658 (N_658,In_1295,In_13);
nor U659 (N_659,In_20,In_1478);
or U660 (N_660,In_862,In_123);
nand U661 (N_661,In_236,In_35);
and U662 (N_662,In_676,In_1017);
nand U663 (N_663,In_1111,In_988);
nand U664 (N_664,In_1056,In_604);
and U665 (N_665,In_1144,In_1470);
or U666 (N_666,In_145,In_1145);
nand U667 (N_667,In_1327,In_482);
and U668 (N_668,In_1260,In_34);
nand U669 (N_669,In_1320,In_1363);
xnor U670 (N_670,In_408,In_1124);
nor U671 (N_671,In_688,In_883);
nor U672 (N_672,In_1249,In_809);
or U673 (N_673,In_103,In_1158);
nor U674 (N_674,In_622,In_1204);
and U675 (N_675,In_923,In_1134);
and U676 (N_676,In_475,In_416);
nand U677 (N_677,In_167,In_742);
nand U678 (N_678,In_1317,In_600);
nand U679 (N_679,In_897,In_315);
or U680 (N_680,In_1001,In_1287);
and U681 (N_681,In_785,In_819);
nor U682 (N_682,In_878,In_605);
nand U683 (N_683,In_981,In_801);
nand U684 (N_684,In_12,In_953);
nor U685 (N_685,In_1266,In_934);
nor U686 (N_686,In_1420,In_547);
xnor U687 (N_687,In_174,In_349);
xnor U688 (N_688,In_255,In_1099);
nand U689 (N_689,In_901,In_1122);
or U690 (N_690,In_1167,In_1394);
nor U691 (N_691,In_1081,In_460);
nand U692 (N_692,In_389,In_613);
nor U693 (N_693,In_135,In_1436);
and U694 (N_694,In_815,In_212);
nand U695 (N_695,In_1069,In_1119);
nor U696 (N_696,In_1149,In_1183);
xnor U697 (N_697,In_266,In_644);
nor U698 (N_698,In_576,In_1349);
nand U699 (N_699,In_45,In_990);
nor U700 (N_700,In_303,In_1409);
nand U701 (N_701,In_595,In_1286);
or U702 (N_702,In_607,In_1129);
or U703 (N_703,In_805,In_692);
nor U704 (N_704,In_244,In_504);
nand U705 (N_705,In_393,In_1310);
or U706 (N_706,In_395,In_542);
xnor U707 (N_707,In_808,In_476);
and U708 (N_708,In_684,In_1339);
nor U709 (N_709,In_449,In_1185);
or U710 (N_710,In_1369,In_314);
and U711 (N_711,In_1308,In_397);
nor U712 (N_712,In_240,In_712);
nor U713 (N_713,In_424,In_686);
or U714 (N_714,In_171,In_1135);
nand U715 (N_715,In_48,In_790);
and U716 (N_716,In_586,In_1071);
nand U717 (N_717,In_797,In_378);
or U718 (N_718,In_822,In_919);
and U719 (N_719,In_917,In_1098);
nand U720 (N_720,In_777,In_1439);
or U721 (N_721,In_399,In_707);
or U722 (N_722,In_872,In_1275);
and U723 (N_723,In_484,In_682);
or U724 (N_724,In_1259,In_521);
nand U725 (N_725,In_957,In_1434);
nand U726 (N_726,In_1189,In_119);
nor U727 (N_727,In_249,In_532);
nor U728 (N_728,In_1257,In_1046);
and U729 (N_729,In_566,In_489);
nand U730 (N_730,In_1058,In_223);
xor U731 (N_731,In_177,In_1404);
and U732 (N_732,In_1499,In_279);
nor U733 (N_733,In_202,In_1370);
nand U734 (N_734,In_137,In_1385);
and U735 (N_735,In_172,In_1195);
or U736 (N_736,In_1397,In_433);
or U737 (N_737,In_182,In_414);
nor U738 (N_738,In_1304,In_582);
or U739 (N_739,In_496,In_1053);
or U740 (N_740,In_384,In_641);
nand U741 (N_741,In_168,In_559);
nand U742 (N_742,In_905,In_1313);
nor U743 (N_743,In_1015,In_1421);
nor U744 (N_744,In_1459,In_1248);
nand U745 (N_745,In_1392,In_451);
and U746 (N_746,In_846,In_1064);
nand U747 (N_747,In_105,In_481);
nand U748 (N_748,In_791,In_1090);
nand U749 (N_749,In_833,In_852);
or U750 (N_750,In_761,In_336);
or U751 (N_751,In_1083,In_1191);
or U752 (N_752,In_43,In_1234);
xor U753 (N_753,In_1415,In_1031);
or U754 (N_754,In_977,In_1457);
or U755 (N_755,In_447,In_200);
nor U756 (N_756,In_1060,In_1303);
or U757 (N_757,In_1417,In_884);
nor U758 (N_758,In_749,In_73);
nand U759 (N_759,In_879,In_773);
and U760 (N_760,In_123,In_1429);
xor U761 (N_761,In_4,In_532);
nor U762 (N_762,In_757,In_970);
nand U763 (N_763,In_861,In_1361);
or U764 (N_764,In_398,In_1147);
or U765 (N_765,In_709,In_829);
nor U766 (N_766,In_1327,In_1102);
or U767 (N_767,In_1036,In_101);
or U768 (N_768,In_114,In_1116);
and U769 (N_769,In_1021,In_453);
nor U770 (N_770,In_1006,In_349);
nor U771 (N_771,In_865,In_1258);
nand U772 (N_772,In_1328,In_868);
nand U773 (N_773,In_412,In_1287);
or U774 (N_774,In_1461,In_1045);
or U775 (N_775,In_959,In_1485);
or U776 (N_776,In_817,In_272);
and U777 (N_777,In_1436,In_1076);
nand U778 (N_778,In_897,In_216);
or U779 (N_779,In_293,In_15);
and U780 (N_780,In_1333,In_730);
nor U781 (N_781,In_397,In_791);
or U782 (N_782,In_444,In_587);
nor U783 (N_783,In_618,In_443);
nand U784 (N_784,In_427,In_310);
nand U785 (N_785,In_145,In_112);
and U786 (N_786,In_1107,In_628);
and U787 (N_787,In_590,In_787);
or U788 (N_788,In_194,In_1079);
nand U789 (N_789,In_1081,In_1450);
and U790 (N_790,In_421,In_725);
and U791 (N_791,In_675,In_193);
xnor U792 (N_792,In_25,In_553);
nand U793 (N_793,In_1398,In_1272);
and U794 (N_794,In_178,In_482);
or U795 (N_795,In_1284,In_1013);
and U796 (N_796,In_1280,In_1168);
nor U797 (N_797,In_1254,In_1203);
nand U798 (N_798,In_1049,In_804);
or U799 (N_799,In_214,In_1143);
and U800 (N_800,In_1434,In_158);
nand U801 (N_801,In_192,In_894);
nor U802 (N_802,In_1115,In_263);
and U803 (N_803,In_988,In_274);
nor U804 (N_804,In_213,In_1373);
xor U805 (N_805,In_1409,In_1049);
or U806 (N_806,In_1033,In_990);
and U807 (N_807,In_172,In_102);
or U808 (N_808,In_1210,In_1226);
or U809 (N_809,In_524,In_1196);
nand U810 (N_810,In_49,In_613);
or U811 (N_811,In_761,In_462);
or U812 (N_812,In_609,In_982);
nand U813 (N_813,In_1325,In_1409);
or U814 (N_814,In_1265,In_378);
nor U815 (N_815,In_1156,In_1351);
and U816 (N_816,In_393,In_38);
or U817 (N_817,In_261,In_510);
nand U818 (N_818,In_196,In_1135);
or U819 (N_819,In_679,In_908);
nor U820 (N_820,In_929,In_499);
xnor U821 (N_821,In_911,In_1117);
nand U822 (N_822,In_840,In_1194);
nand U823 (N_823,In_1422,In_580);
nand U824 (N_824,In_1169,In_1151);
nand U825 (N_825,In_145,In_262);
xor U826 (N_826,In_486,In_1439);
or U827 (N_827,In_544,In_1062);
nor U828 (N_828,In_1038,In_402);
or U829 (N_829,In_645,In_1199);
and U830 (N_830,In_504,In_393);
and U831 (N_831,In_376,In_403);
nand U832 (N_832,In_802,In_747);
nand U833 (N_833,In_666,In_1442);
and U834 (N_834,In_12,In_749);
nand U835 (N_835,In_152,In_1437);
nand U836 (N_836,In_854,In_1274);
or U837 (N_837,In_229,In_1482);
and U838 (N_838,In_771,In_1471);
nor U839 (N_839,In_1245,In_1164);
nor U840 (N_840,In_1180,In_833);
nand U841 (N_841,In_520,In_410);
nand U842 (N_842,In_371,In_818);
or U843 (N_843,In_883,In_761);
nor U844 (N_844,In_943,In_85);
nand U845 (N_845,In_186,In_55);
and U846 (N_846,In_1412,In_1190);
or U847 (N_847,In_955,In_909);
nor U848 (N_848,In_1379,In_102);
nor U849 (N_849,In_674,In_287);
nor U850 (N_850,In_1336,In_55);
and U851 (N_851,In_542,In_42);
nor U852 (N_852,In_1436,In_177);
and U853 (N_853,In_900,In_321);
nor U854 (N_854,In_1157,In_425);
nand U855 (N_855,In_307,In_1022);
nor U856 (N_856,In_550,In_1262);
nor U857 (N_857,In_1127,In_555);
xor U858 (N_858,In_1147,In_114);
and U859 (N_859,In_1302,In_633);
and U860 (N_860,In_1480,In_1152);
and U861 (N_861,In_270,In_750);
nand U862 (N_862,In_682,In_133);
nand U863 (N_863,In_209,In_807);
nor U864 (N_864,In_254,In_1390);
and U865 (N_865,In_1482,In_715);
nor U866 (N_866,In_1454,In_759);
xor U867 (N_867,In_1039,In_773);
nor U868 (N_868,In_682,In_353);
nor U869 (N_869,In_1387,In_952);
nand U870 (N_870,In_1131,In_473);
or U871 (N_871,In_781,In_1365);
and U872 (N_872,In_74,In_1345);
and U873 (N_873,In_1212,In_321);
or U874 (N_874,In_676,In_602);
and U875 (N_875,In_71,In_1472);
nand U876 (N_876,In_475,In_51);
and U877 (N_877,In_354,In_1474);
nand U878 (N_878,In_205,In_373);
or U879 (N_879,In_779,In_1326);
nand U880 (N_880,In_90,In_475);
and U881 (N_881,In_1169,In_920);
nor U882 (N_882,In_891,In_1339);
or U883 (N_883,In_1458,In_463);
nand U884 (N_884,In_943,In_1021);
or U885 (N_885,In_10,In_1407);
nor U886 (N_886,In_1000,In_498);
or U887 (N_887,In_471,In_969);
and U888 (N_888,In_1438,In_267);
nand U889 (N_889,In_1248,In_698);
and U890 (N_890,In_778,In_1395);
nand U891 (N_891,In_446,In_924);
nor U892 (N_892,In_1319,In_892);
nand U893 (N_893,In_971,In_699);
nor U894 (N_894,In_51,In_1044);
nand U895 (N_895,In_175,In_1407);
and U896 (N_896,In_58,In_161);
nor U897 (N_897,In_594,In_726);
or U898 (N_898,In_434,In_669);
nand U899 (N_899,In_466,In_249);
nor U900 (N_900,In_1332,In_1485);
and U901 (N_901,In_73,In_530);
and U902 (N_902,In_1416,In_610);
nand U903 (N_903,In_658,In_99);
or U904 (N_904,In_874,In_1194);
or U905 (N_905,In_1277,In_856);
nand U906 (N_906,In_1137,In_88);
or U907 (N_907,In_1094,In_17);
nand U908 (N_908,In_263,In_557);
nor U909 (N_909,In_658,In_405);
nor U910 (N_910,In_120,In_925);
or U911 (N_911,In_589,In_277);
nand U912 (N_912,In_455,In_1050);
or U913 (N_913,In_203,In_339);
nand U914 (N_914,In_911,In_605);
or U915 (N_915,In_893,In_165);
or U916 (N_916,In_542,In_52);
and U917 (N_917,In_1392,In_73);
nor U918 (N_918,In_129,In_978);
xor U919 (N_919,In_1424,In_524);
or U920 (N_920,In_654,In_670);
nor U921 (N_921,In_1425,In_278);
nor U922 (N_922,In_180,In_1070);
and U923 (N_923,In_1172,In_1189);
nand U924 (N_924,In_591,In_909);
xor U925 (N_925,In_1302,In_42);
and U926 (N_926,In_72,In_1402);
nand U927 (N_927,In_690,In_865);
nor U928 (N_928,In_1287,In_568);
nor U929 (N_929,In_540,In_79);
nor U930 (N_930,In_839,In_1391);
or U931 (N_931,In_1031,In_294);
nand U932 (N_932,In_1275,In_502);
and U933 (N_933,In_185,In_644);
nor U934 (N_934,In_1041,In_413);
or U935 (N_935,In_377,In_1025);
nor U936 (N_936,In_167,In_1184);
or U937 (N_937,In_164,In_348);
and U938 (N_938,In_623,In_681);
nor U939 (N_939,In_813,In_754);
nor U940 (N_940,In_649,In_278);
nand U941 (N_941,In_1464,In_1010);
or U942 (N_942,In_953,In_1);
or U943 (N_943,In_263,In_665);
or U944 (N_944,In_467,In_725);
and U945 (N_945,In_739,In_1172);
and U946 (N_946,In_1189,In_543);
nor U947 (N_947,In_605,In_942);
and U948 (N_948,In_68,In_299);
nand U949 (N_949,In_1183,In_94);
and U950 (N_950,In_1233,In_1479);
nor U951 (N_951,In_1439,In_427);
or U952 (N_952,In_485,In_220);
nand U953 (N_953,In_1181,In_285);
xor U954 (N_954,In_1350,In_898);
or U955 (N_955,In_460,In_909);
or U956 (N_956,In_286,In_732);
or U957 (N_957,In_904,In_345);
and U958 (N_958,In_1117,In_1076);
and U959 (N_959,In_1407,In_968);
or U960 (N_960,In_592,In_1418);
and U961 (N_961,In_1075,In_893);
or U962 (N_962,In_784,In_284);
and U963 (N_963,In_331,In_1282);
nand U964 (N_964,In_1391,In_78);
xor U965 (N_965,In_1253,In_536);
or U966 (N_966,In_339,In_1362);
nor U967 (N_967,In_998,In_213);
nand U968 (N_968,In_216,In_491);
or U969 (N_969,In_1349,In_1468);
nor U970 (N_970,In_111,In_1218);
nand U971 (N_971,In_1430,In_961);
nand U972 (N_972,In_530,In_334);
xnor U973 (N_973,In_30,In_759);
nor U974 (N_974,In_448,In_1268);
xnor U975 (N_975,In_210,In_1090);
nand U976 (N_976,In_1275,In_104);
nand U977 (N_977,In_537,In_1454);
nand U978 (N_978,In_1346,In_651);
nor U979 (N_979,In_750,In_1474);
nand U980 (N_980,In_1021,In_567);
nand U981 (N_981,In_934,In_233);
and U982 (N_982,In_862,In_1330);
or U983 (N_983,In_1314,In_120);
nand U984 (N_984,In_510,In_48);
and U985 (N_985,In_226,In_1413);
nand U986 (N_986,In_285,In_126);
nand U987 (N_987,In_1171,In_983);
nor U988 (N_988,In_114,In_1349);
nor U989 (N_989,In_467,In_373);
nand U990 (N_990,In_811,In_1376);
nor U991 (N_991,In_375,In_740);
or U992 (N_992,In_404,In_1082);
and U993 (N_993,In_1026,In_673);
and U994 (N_994,In_560,In_638);
and U995 (N_995,In_700,In_1122);
nor U996 (N_996,In_933,In_657);
and U997 (N_997,In_317,In_928);
nor U998 (N_998,In_818,In_1034);
and U999 (N_999,In_242,In_2);
or U1000 (N_1000,In_985,In_105);
or U1001 (N_1001,In_322,In_910);
or U1002 (N_1002,In_214,In_27);
or U1003 (N_1003,In_1198,In_330);
and U1004 (N_1004,In_700,In_1277);
nand U1005 (N_1005,In_1240,In_500);
nor U1006 (N_1006,In_520,In_1438);
or U1007 (N_1007,In_1386,In_1200);
nor U1008 (N_1008,In_155,In_525);
nand U1009 (N_1009,In_1459,In_951);
and U1010 (N_1010,In_954,In_1493);
nor U1011 (N_1011,In_1354,In_479);
xnor U1012 (N_1012,In_245,In_700);
xor U1013 (N_1013,In_772,In_1015);
and U1014 (N_1014,In_51,In_1267);
nand U1015 (N_1015,In_1256,In_482);
xnor U1016 (N_1016,In_993,In_1057);
nand U1017 (N_1017,In_59,In_434);
or U1018 (N_1018,In_469,In_682);
or U1019 (N_1019,In_1069,In_542);
or U1020 (N_1020,In_179,In_386);
and U1021 (N_1021,In_1016,In_344);
and U1022 (N_1022,In_268,In_1201);
nor U1023 (N_1023,In_539,In_87);
nand U1024 (N_1024,In_307,In_611);
nand U1025 (N_1025,In_1041,In_219);
nor U1026 (N_1026,In_223,In_819);
nand U1027 (N_1027,In_410,In_56);
nand U1028 (N_1028,In_87,In_1106);
nor U1029 (N_1029,In_831,In_898);
xor U1030 (N_1030,In_1307,In_1131);
nor U1031 (N_1031,In_522,In_929);
or U1032 (N_1032,In_105,In_1287);
nor U1033 (N_1033,In_636,In_1123);
nor U1034 (N_1034,In_1385,In_855);
nor U1035 (N_1035,In_1127,In_204);
nor U1036 (N_1036,In_1184,In_595);
nand U1037 (N_1037,In_89,In_731);
nor U1038 (N_1038,In_166,In_24);
or U1039 (N_1039,In_1094,In_1492);
or U1040 (N_1040,In_1425,In_1282);
nand U1041 (N_1041,In_215,In_981);
nor U1042 (N_1042,In_236,In_1039);
nor U1043 (N_1043,In_189,In_512);
nand U1044 (N_1044,In_40,In_1171);
and U1045 (N_1045,In_1183,In_421);
or U1046 (N_1046,In_580,In_1458);
or U1047 (N_1047,In_1205,In_65);
nor U1048 (N_1048,In_158,In_1179);
nand U1049 (N_1049,In_244,In_765);
nor U1050 (N_1050,In_959,In_255);
and U1051 (N_1051,In_318,In_1237);
nand U1052 (N_1052,In_1063,In_123);
nor U1053 (N_1053,In_951,In_834);
and U1054 (N_1054,In_445,In_554);
nor U1055 (N_1055,In_1366,In_363);
nor U1056 (N_1056,In_1221,In_1314);
and U1057 (N_1057,In_305,In_582);
nor U1058 (N_1058,In_1151,In_1414);
xnor U1059 (N_1059,In_297,In_22);
nor U1060 (N_1060,In_173,In_925);
or U1061 (N_1061,In_1389,In_996);
or U1062 (N_1062,In_681,In_1135);
and U1063 (N_1063,In_1023,In_651);
nor U1064 (N_1064,In_1421,In_615);
and U1065 (N_1065,In_1368,In_1376);
nand U1066 (N_1066,In_68,In_1153);
nor U1067 (N_1067,In_685,In_709);
and U1068 (N_1068,In_1377,In_1270);
nand U1069 (N_1069,In_1107,In_1445);
nand U1070 (N_1070,In_825,In_974);
nor U1071 (N_1071,In_1385,In_560);
or U1072 (N_1072,In_1260,In_1358);
nand U1073 (N_1073,In_791,In_148);
or U1074 (N_1074,In_354,In_1435);
nor U1075 (N_1075,In_723,In_286);
or U1076 (N_1076,In_308,In_684);
nor U1077 (N_1077,In_166,In_633);
or U1078 (N_1078,In_250,In_1217);
nand U1079 (N_1079,In_209,In_293);
nor U1080 (N_1080,In_876,In_1277);
and U1081 (N_1081,In_146,In_1402);
nor U1082 (N_1082,In_1016,In_1204);
or U1083 (N_1083,In_1447,In_1415);
nor U1084 (N_1084,In_869,In_750);
nor U1085 (N_1085,In_1104,In_293);
nand U1086 (N_1086,In_263,In_993);
xor U1087 (N_1087,In_247,In_841);
nand U1088 (N_1088,In_1111,In_744);
nand U1089 (N_1089,In_1483,In_329);
nor U1090 (N_1090,In_1279,In_283);
or U1091 (N_1091,In_578,In_286);
and U1092 (N_1092,In_676,In_354);
nor U1093 (N_1093,In_767,In_1394);
nor U1094 (N_1094,In_446,In_258);
and U1095 (N_1095,In_574,In_900);
nand U1096 (N_1096,In_1162,In_638);
and U1097 (N_1097,In_963,In_247);
or U1098 (N_1098,In_1458,In_843);
and U1099 (N_1099,In_1279,In_1189);
or U1100 (N_1100,In_89,In_782);
nand U1101 (N_1101,In_348,In_321);
and U1102 (N_1102,In_220,In_1142);
nor U1103 (N_1103,In_505,In_347);
nand U1104 (N_1104,In_603,In_1488);
nor U1105 (N_1105,In_1074,In_315);
nand U1106 (N_1106,In_933,In_518);
xnor U1107 (N_1107,In_731,In_746);
nor U1108 (N_1108,In_983,In_1390);
nor U1109 (N_1109,In_977,In_201);
nand U1110 (N_1110,In_423,In_821);
or U1111 (N_1111,In_1016,In_1220);
nand U1112 (N_1112,In_456,In_274);
nand U1113 (N_1113,In_245,In_999);
and U1114 (N_1114,In_915,In_265);
or U1115 (N_1115,In_36,In_207);
and U1116 (N_1116,In_856,In_589);
or U1117 (N_1117,In_777,In_1068);
nor U1118 (N_1118,In_82,In_297);
or U1119 (N_1119,In_667,In_85);
or U1120 (N_1120,In_1453,In_443);
or U1121 (N_1121,In_685,In_762);
and U1122 (N_1122,In_968,In_816);
nand U1123 (N_1123,In_815,In_1471);
and U1124 (N_1124,In_1165,In_1048);
nand U1125 (N_1125,In_936,In_906);
nand U1126 (N_1126,In_53,In_1233);
nand U1127 (N_1127,In_1474,In_1024);
nand U1128 (N_1128,In_1375,In_520);
nand U1129 (N_1129,In_887,In_937);
xor U1130 (N_1130,In_974,In_1292);
and U1131 (N_1131,In_570,In_444);
and U1132 (N_1132,In_468,In_1347);
and U1133 (N_1133,In_84,In_1360);
and U1134 (N_1134,In_686,In_1282);
and U1135 (N_1135,In_1461,In_238);
or U1136 (N_1136,In_826,In_1237);
or U1137 (N_1137,In_13,In_136);
or U1138 (N_1138,In_138,In_1010);
nand U1139 (N_1139,In_42,In_1480);
nand U1140 (N_1140,In_1169,In_638);
nor U1141 (N_1141,In_154,In_1163);
nor U1142 (N_1142,In_261,In_1423);
and U1143 (N_1143,In_428,In_1013);
and U1144 (N_1144,In_435,In_1022);
and U1145 (N_1145,In_1245,In_16);
and U1146 (N_1146,In_1035,In_537);
nor U1147 (N_1147,In_443,In_623);
nand U1148 (N_1148,In_976,In_943);
or U1149 (N_1149,In_897,In_562);
and U1150 (N_1150,In_1305,In_551);
or U1151 (N_1151,In_222,In_613);
or U1152 (N_1152,In_728,In_774);
nand U1153 (N_1153,In_687,In_323);
or U1154 (N_1154,In_35,In_1441);
or U1155 (N_1155,In_557,In_748);
nor U1156 (N_1156,In_831,In_1175);
nand U1157 (N_1157,In_1193,In_227);
and U1158 (N_1158,In_852,In_92);
and U1159 (N_1159,In_875,In_65);
and U1160 (N_1160,In_808,In_1264);
nand U1161 (N_1161,In_1006,In_1117);
nor U1162 (N_1162,In_791,In_1178);
or U1163 (N_1163,In_749,In_1138);
nand U1164 (N_1164,In_1128,In_1081);
and U1165 (N_1165,In_415,In_342);
nor U1166 (N_1166,In_155,In_378);
nor U1167 (N_1167,In_1262,In_1354);
and U1168 (N_1168,In_801,In_587);
nor U1169 (N_1169,In_884,In_1472);
or U1170 (N_1170,In_1398,In_1261);
nor U1171 (N_1171,In_758,In_827);
and U1172 (N_1172,In_57,In_1495);
nand U1173 (N_1173,In_152,In_519);
and U1174 (N_1174,In_1404,In_230);
and U1175 (N_1175,In_497,In_1339);
nor U1176 (N_1176,In_1233,In_1);
xnor U1177 (N_1177,In_273,In_1066);
and U1178 (N_1178,In_785,In_106);
nand U1179 (N_1179,In_1188,In_600);
and U1180 (N_1180,In_939,In_456);
and U1181 (N_1181,In_360,In_885);
or U1182 (N_1182,In_1065,In_966);
nor U1183 (N_1183,In_1389,In_289);
or U1184 (N_1184,In_1156,In_960);
nand U1185 (N_1185,In_870,In_884);
nor U1186 (N_1186,In_326,In_1221);
nor U1187 (N_1187,In_588,In_433);
xor U1188 (N_1188,In_35,In_1434);
nor U1189 (N_1189,In_634,In_594);
nor U1190 (N_1190,In_1334,In_1406);
and U1191 (N_1191,In_1149,In_1169);
nand U1192 (N_1192,In_515,In_1454);
nor U1193 (N_1193,In_1218,In_1194);
and U1194 (N_1194,In_1012,In_1382);
nand U1195 (N_1195,In_1407,In_127);
nor U1196 (N_1196,In_1301,In_1235);
and U1197 (N_1197,In_873,In_72);
nand U1198 (N_1198,In_967,In_224);
or U1199 (N_1199,In_1088,In_811);
or U1200 (N_1200,In_1161,In_1255);
or U1201 (N_1201,In_828,In_1437);
or U1202 (N_1202,In_1420,In_1493);
nand U1203 (N_1203,In_1187,In_338);
and U1204 (N_1204,In_1029,In_1344);
nand U1205 (N_1205,In_797,In_788);
nor U1206 (N_1206,In_174,In_477);
nand U1207 (N_1207,In_1257,In_339);
or U1208 (N_1208,In_720,In_1346);
nand U1209 (N_1209,In_711,In_1219);
or U1210 (N_1210,In_286,In_859);
nand U1211 (N_1211,In_875,In_1020);
and U1212 (N_1212,In_713,In_732);
nor U1213 (N_1213,In_745,In_1104);
or U1214 (N_1214,In_228,In_1309);
nor U1215 (N_1215,In_335,In_480);
nand U1216 (N_1216,In_757,In_877);
or U1217 (N_1217,In_509,In_1210);
nand U1218 (N_1218,In_762,In_314);
nand U1219 (N_1219,In_1150,In_578);
nor U1220 (N_1220,In_495,In_531);
and U1221 (N_1221,In_726,In_1448);
nand U1222 (N_1222,In_249,In_1098);
nand U1223 (N_1223,In_1127,In_224);
nor U1224 (N_1224,In_503,In_1244);
nand U1225 (N_1225,In_274,In_804);
or U1226 (N_1226,In_1329,In_1135);
or U1227 (N_1227,In_1448,In_122);
xor U1228 (N_1228,In_713,In_503);
nand U1229 (N_1229,In_16,In_580);
nor U1230 (N_1230,In_976,In_1321);
and U1231 (N_1231,In_599,In_304);
nor U1232 (N_1232,In_788,In_700);
and U1233 (N_1233,In_956,In_1400);
nor U1234 (N_1234,In_693,In_160);
and U1235 (N_1235,In_961,In_554);
nand U1236 (N_1236,In_512,In_637);
and U1237 (N_1237,In_54,In_446);
or U1238 (N_1238,In_52,In_511);
nor U1239 (N_1239,In_904,In_210);
nor U1240 (N_1240,In_126,In_907);
nor U1241 (N_1241,In_216,In_723);
nor U1242 (N_1242,In_7,In_156);
nor U1243 (N_1243,In_237,In_1093);
or U1244 (N_1244,In_223,In_532);
and U1245 (N_1245,In_1266,In_651);
and U1246 (N_1246,In_725,In_523);
and U1247 (N_1247,In_7,In_223);
nand U1248 (N_1248,In_18,In_1198);
xor U1249 (N_1249,In_966,In_803);
and U1250 (N_1250,In_48,In_1178);
and U1251 (N_1251,In_1498,In_56);
nand U1252 (N_1252,In_1241,In_907);
nand U1253 (N_1253,In_519,In_888);
nor U1254 (N_1254,In_115,In_393);
nor U1255 (N_1255,In_706,In_51);
nand U1256 (N_1256,In_1448,In_1054);
nor U1257 (N_1257,In_961,In_331);
and U1258 (N_1258,In_790,In_1017);
nor U1259 (N_1259,In_1438,In_1426);
and U1260 (N_1260,In_1343,In_1101);
nand U1261 (N_1261,In_1374,In_1483);
or U1262 (N_1262,In_647,In_1290);
or U1263 (N_1263,In_1400,In_1224);
nand U1264 (N_1264,In_127,In_101);
or U1265 (N_1265,In_322,In_959);
nor U1266 (N_1266,In_1176,In_229);
and U1267 (N_1267,In_780,In_1161);
nor U1268 (N_1268,In_702,In_824);
nor U1269 (N_1269,In_1412,In_900);
or U1270 (N_1270,In_1288,In_1154);
and U1271 (N_1271,In_480,In_298);
nand U1272 (N_1272,In_1266,In_379);
nand U1273 (N_1273,In_958,In_568);
nand U1274 (N_1274,In_847,In_434);
xor U1275 (N_1275,In_1021,In_613);
nand U1276 (N_1276,In_518,In_471);
and U1277 (N_1277,In_853,In_375);
nand U1278 (N_1278,In_473,In_523);
and U1279 (N_1279,In_476,In_917);
and U1280 (N_1280,In_782,In_181);
or U1281 (N_1281,In_1212,In_1124);
nand U1282 (N_1282,In_49,In_566);
or U1283 (N_1283,In_556,In_903);
nand U1284 (N_1284,In_1106,In_317);
nand U1285 (N_1285,In_1406,In_1057);
nor U1286 (N_1286,In_942,In_299);
or U1287 (N_1287,In_682,In_667);
nand U1288 (N_1288,In_131,In_1040);
nand U1289 (N_1289,In_82,In_760);
xor U1290 (N_1290,In_98,In_1104);
and U1291 (N_1291,In_1426,In_88);
or U1292 (N_1292,In_604,In_821);
and U1293 (N_1293,In_541,In_890);
nand U1294 (N_1294,In_751,In_927);
nand U1295 (N_1295,In_1446,In_213);
or U1296 (N_1296,In_1131,In_328);
or U1297 (N_1297,In_1364,In_263);
nor U1298 (N_1298,In_1162,In_52);
nand U1299 (N_1299,In_770,In_1053);
xor U1300 (N_1300,In_448,In_852);
nor U1301 (N_1301,In_432,In_1299);
nor U1302 (N_1302,In_1474,In_147);
nor U1303 (N_1303,In_1445,In_836);
and U1304 (N_1304,In_1064,In_837);
or U1305 (N_1305,In_157,In_1493);
and U1306 (N_1306,In_887,In_766);
nand U1307 (N_1307,In_489,In_280);
nor U1308 (N_1308,In_871,In_997);
and U1309 (N_1309,In_1429,In_713);
or U1310 (N_1310,In_978,In_756);
nand U1311 (N_1311,In_156,In_59);
nand U1312 (N_1312,In_817,In_1335);
or U1313 (N_1313,In_869,In_566);
nor U1314 (N_1314,In_901,In_829);
nor U1315 (N_1315,In_42,In_742);
nand U1316 (N_1316,In_1460,In_357);
or U1317 (N_1317,In_850,In_846);
nor U1318 (N_1318,In_622,In_189);
nor U1319 (N_1319,In_1469,In_1491);
and U1320 (N_1320,In_588,In_231);
and U1321 (N_1321,In_519,In_1238);
or U1322 (N_1322,In_859,In_221);
nor U1323 (N_1323,In_151,In_48);
and U1324 (N_1324,In_366,In_441);
and U1325 (N_1325,In_1046,In_364);
nor U1326 (N_1326,In_425,In_1254);
nor U1327 (N_1327,In_454,In_804);
and U1328 (N_1328,In_306,In_158);
nand U1329 (N_1329,In_1276,In_221);
nor U1330 (N_1330,In_1185,In_677);
nor U1331 (N_1331,In_1371,In_272);
nand U1332 (N_1332,In_517,In_1085);
and U1333 (N_1333,In_1118,In_486);
nand U1334 (N_1334,In_1325,In_888);
nor U1335 (N_1335,In_1450,In_1172);
nor U1336 (N_1336,In_1001,In_732);
or U1337 (N_1337,In_867,In_848);
nand U1338 (N_1338,In_556,In_724);
nor U1339 (N_1339,In_874,In_612);
nor U1340 (N_1340,In_1009,In_1058);
nand U1341 (N_1341,In_1369,In_720);
nor U1342 (N_1342,In_1239,In_713);
nor U1343 (N_1343,In_515,In_511);
nand U1344 (N_1344,In_1128,In_805);
and U1345 (N_1345,In_249,In_642);
nor U1346 (N_1346,In_1430,In_610);
and U1347 (N_1347,In_127,In_1204);
or U1348 (N_1348,In_1068,In_595);
nor U1349 (N_1349,In_460,In_591);
and U1350 (N_1350,In_1082,In_34);
or U1351 (N_1351,In_1448,In_1164);
nand U1352 (N_1352,In_1068,In_370);
nor U1353 (N_1353,In_990,In_1263);
and U1354 (N_1354,In_34,In_1320);
or U1355 (N_1355,In_429,In_820);
nand U1356 (N_1356,In_958,In_1224);
nor U1357 (N_1357,In_290,In_1188);
and U1358 (N_1358,In_702,In_169);
nand U1359 (N_1359,In_669,In_29);
nand U1360 (N_1360,In_512,In_257);
or U1361 (N_1361,In_1439,In_334);
and U1362 (N_1362,In_1328,In_5);
nand U1363 (N_1363,In_677,In_1402);
nand U1364 (N_1364,In_1478,In_200);
and U1365 (N_1365,In_641,In_214);
nor U1366 (N_1366,In_1095,In_17);
nand U1367 (N_1367,In_1167,In_1303);
nand U1368 (N_1368,In_470,In_915);
and U1369 (N_1369,In_712,In_637);
nand U1370 (N_1370,In_985,In_761);
and U1371 (N_1371,In_595,In_1498);
or U1372 (N_1372,In_1361,In_1224);
nand U1373 (N_1373,In_733,In_189);
nor U1374 (N_1374,In_132,In_1091);
or U1375 (N_1375,In_916,In_258);
and U1376 (N_1376,In_846,In_1171);
nor U1377 (N_1377,In_4,In_864);
or U1378 (N_1378,In_1236,In_235);
nor U1379 (N_1379,In_478,In_1473);
nand U1380 (N_1380,In_704,In_1135);
or U1381 (N_1381,In_461,In_903);
or U1382 (N_1382,In_789,In_129);
and U1383 (N_1383,In_9,In_1046);
xor U1384 (N_1384,In_916,In_391);
or U1385 (N_1385,In_1384,In_1072);
xnor U1386 (N_1386,In_1407,In_582);
or U1387 (N_1387,In_1400,In_900);
and U1388 (N_1388,In_207,In_891);
nand U1389 (N_1389,In_1464,In_58);
and U1390 (N_1390,In_151,In_303);
nor U1391 (N_1391,In_933,In_1280);
nor U1392 (N_1392,In_168,In_30);
nor U1393 (N_1393,In_558,In_752);
nand U1394 (N_1394,In_249,In_100);
or U1395 (N_1395,In_157,In_211);
nor U1396 (N_1396,In_953,In_1026);
and U1397 (N_1397,In_1044,In_103);
nand U1398 (N_1398,In_1212,In_66);
and U1399 (N_1399,In_57,In_112);
and U1400 (N_1400,In_612,In_889);
or U1401 (N_1401,In_442,In_979);
or U1402 (N_1402,In_1499,In_466);
and U1403 (N_1403,In_73,In_76);
and U1404 (N_1404,In_1376,In_1306);
and U1405 (N_1405,In_91,In_1119);
or U1406 (N_1406,In_29,In_292);
nand U1407 (N_1407,In_499,In_19);
or U1408 (N_1408,In_523,In_1228);
nor U1409 (N_1409,In_22,In_622);
nand U1410 (N_1410,In_488,In_444);
and U1411 (N_1411,In_1219,In_1473);
nor U1412 (N_1412,In_67,In_510);
and U1413 (N_1413,In_380,In_1021);
nor U1414 (N_1414,In_900,In_855);
nor U1415 (N_1415,In_1205,In_732);
nand U1416 (N_1416,In_326,In_463);
xnor U1417 (N_1417,In_951,In_715);
nor U1418 (N_1418,In_52,In_1247);
or U1419 (N_1419,In_472,In_960);
xnor U1420 (N_1420,In_805,In_663);
nor U1421 (N_1421,In_1140,In_131);
nor U1422 (N_1422,In_226,In_959);
and U1423 (N_1423,In_1267,In_944);
and U1424 (N_1424,In_322,In_886);
and U1425 (N_1425,In_363,In_685);
and U1426 (N_1426,In_947,In_370);
nand U1427 (N_1427,In_1474,In_662);
nand U1428 (N_1428,In_1363,In_969);
nor U1429 (N_1429,In_1457,In_206);
and U1430 (N_1430,In_136,In_993);
or U1431 (N_1431,In_9,In_292);
or U1432 (N_1432,In_682,In_1153);
and U1433 (N_1433,In_1483,In_1059);
or U1434 (N_1434,In_810,In_1226);
nor U1435 (N_1435,In_222,In_1111);
and U1436 (N_1436,In_1236,In_1422);
nor U1437 (N_1437,In_636,In_1457);
and U1438 (N_1438,In_940,In_782);
xor U1439 (N_1439,In_965,In_383);
nor U1440 (N_1440,In_259,In_500);
nand U1441 (N_1441,In_1140,In_389);
nand U1442 (N_1442,In_163,In_1066);
nand U1443 (N_1443,In_772,In_413);
nand U1444 (N_1444,In_1455,In_6);
nand U1445 (N_1445,In_565,In_1410);
xor U1446 (N_1446,In_584,In_933);
or U1447 (N_1447,In_868,In_883);
nand U1448 (N_1448,In_954,In_1010);
and U1449 (N_1449,In_1128,In_91);
or U1450 (N_1450,In_422,In_523);
nand U1451 (N_1451,In_1469,In_1018);
or U1452 (N_1452,In_547,In_298);
or U1453 (N_1453,In_739,In_1182);
and U1454 (N_1454,In_1132,In_367);
nand U1455 (N_1455,In_1150,In_702);
nor U1456 (N_1456,In_54,In_741);
or U1457 (N_1457,In_662,In_899);
or U1458 (N_1458,In_118,In_962);
nand U1459 (N_1459,In_1300,In_2);
nand U1460 (N_1460,In_927,In_511);
and U1461 (N_1461,In_48,In_431);
or U1462 (N_1462,In_1319,In_279);
nand U1463 (N_1463,In_613,In_713);
nor U1464 (N_1464,In_285,In_1046);
or U1465 (N_1465,In_889,In_309);
nand U1466 (N_1466,In_1338,In_1046);
or U1467 (N_1467,In_588,In_816);
nand U1468 (N_1468,In_1321,In_1073);
nand U1469 (N_1469,In_1095,In_506);
nor U1470 (N_1470,In_472,In_1066);
nor U1471 (N_1471,In_1065,In_182);
and U1472 (N_1472,In_298,In_571);
nor U1473 (N_1473,In_291,In_1019);
nor U1474 (N_1474,In_802,In_969);
nand U1475 (N_1475,In_353,In_396);
nor U1476 (N_1476,In_575,In_1138);
nor U1477 (N_1477,In_779,In_1031);
and U1478 (N_1478,In_653,In_553);
nor U1479 (N_1479,In_168,In_270);
nand U1480 (N_1480,In_686,In_601);
nor U1481 (N_1481,In_776,In_665);
and U1482 (N_1482,In_117,In_508);
nor U1483 (N_1483,In_829,In_955);
nor U1484 (N_1484,In_161,In_809);
nor U1485 (N_1485,In_465,In_871);
nor U1486 (N_1486,In_1185,In_1082);
nor U1487 (N_1487,In_819,In_1407);
nand U1488 (N_1488,In_782,In_198);
and U1489 (N_1489,In_1165,In_1294);
nand U1490 (N_1490,In_259,In_1115);
nor U1491 (N_1491,In_1211,In_9);
nor U1492 (N_1492,In_231,In_841);
and U1493 (N_1493,In_995,In_1038);
or U1494 (N_1494,In_641,In_397);
xor U1495 (N_1495,In_494,In_398);
nand U1496 (N_1496,In_610,In_782);
xor U1497 (N_1497,In_958,In_309);
nor U1498 (N_1498,In_291,In_888);
or U1499 (N_1499,In_325,In_536);
nor U1500 (N_1500,In_230,In_801);
and U1501 (N_1501,In_1402,In_912);
nand U1502 (N_1502,In_273,In_62);
nand U1503 (N_1503,In_377,In_1244);
nor U1504 (N_1504,In_201,In_175);
and U1505 (N_1505,In_699,In_1067);
nand U1506 (N_1506,In_759,In_1033);
xor U1507 (N_1507,In_1303,In_300);
or U1508 (N_1508,In_1187,In_391);
nor U1509 (N_1509,In_1055,In_765);
or U1510 (N_1510,In_690,In_396);
nor U1511 (N_1511,In_428,In_384);
nand U1512 (N_1512,In_874,In_480);
and U1513 (N_1513,In_946,In_35);
and U1514 (N_1514,In_337,In_12);
nand U1515 (N_1515,In_197,In_1338);
or U1516 (N_1516,In_1305,In_279);
or U1517 (N_1517,In_835,In_309);
and U1518 (N_1518,In_683,In_948);
nor U1519 (N_1519,In_233,In_575);
nand U1520 (N_1520,In_0,In_786);
and U1521 (N_1521,In_1278,In_987);
and U1522 (N_1522,In_453,In_602);
and U1523 (N_1523,In_1494,In_838);
or U1524 (N_1524,In_795,In_345);
and U1525 (N_1525,In_1150,In_1452);
or U1526 (N_1526,In_447,In_1444);
nor U1527 (N_1527,In_572,In_1424);
nand U1528 (N_1528,In_1459,In_165);
or U1529 (N_1529,In_1000,In_921);
nand U1530 (N_1530,In_810,In_446);
and U1531 (N_1531,In_173,In_993);
nor U1532 (N_1532,In_1247,In_1495);
or U1533 (N_1533,In_502,In_124);
or U1534 (N_1534,In_425,In_1457);
or U1535 (N_1535,In_760,In_1080);
or U1536 (N_1536,In_98,In_211);
and U1537 (N_1537,In_1437,In_199);
nor U1538 (N_1538,In_614,In_48);
nor U1539 (N_1539,In_1325,In_417);
nor U1540 (N_1540,In_1286,In_631);
or U1541 (N_1541,In_141,In_1314);
and U1542 (N_1542,In_407,In_898);
and U1543 (N_1543,In_62,In_1206);
nor U1544 (N_1544,In_1145,In_9);
or U1545 (N_1545,In_830,In_626);
or U1546 (N_1546,In_1174,In_82);
xor U1547 (N_1547,In_1027,In_752);
nand U1548 (N_1548,In_504,In_781);
nand U1549 (N_1549,In_1469,In_1430);
nor U1550 (N_1550,In_1098,In_549);
and U1551 (N_1551,In_1179,In_1215);
or U1552 (N_1552,In_399,In_85);
nand U1553 (N_1553,In_189,In_637);
nor U1554 (N_1554,In_245,In_614);
nand U1555 (N_1555,In_1318,In_1249);
or U1556 (N_1556,In_1354,In_1269);
nand U1557 (N_1557,In_521,In_654);
nand U1558 (N_1558,In_413,In_1259);
nand U1559 (N_1559,In_731,In_1178);
nor U1560 (N_1560,In_605,In_198);
and U1561 (N_1561,In_587,In_54);
and U1562 (N_1562,In_581,In_77);
and U1563 (N_1563,In_1257,In_1474);
or U1564 (N_1564,In_548,In_1437);
nor U1565 (N_1565,In_904,In_635);
or U1566 (N_1566,In_1429,In_420);
and U1567 (N_1567,In_62,In_676);
or U1568 (N_1568,In_1253,In_1393);
nand U1569 (N_1569,In_1036,In_435);
nand U1570 (N_1570,In_1439,In_739);
nand U1571 (N_1571,In_180,In_1354);
or U1572 (N_1572,In_178,In_1425);
nand U1573 (N_1573,In_1283,In_590);
and U1574 (N_1574,In_1337,In_619);
nand U1575 (N_1575,In_597,In_298);
or U1576 (N_1576,In_1337,In_960);
nor U1577 (N_1577,In_787,In_918);
or U1578 (N_1578,In_1312,In_987);
nor U1579 (N_1579,In_817,In_1205);
xnor U1580 (N_1580,In_924,In_149);
nor U1581 (N_1581,In_1115,In_351);
or U1582 (N_1582,In_180,In_234);
nand U1583 (N_1583,In_461,In_273);
nand U1584 (N_1584,In_86,In_1426);
nor U1585 (N_1585,In_821,In_621);
or U1586 (N_1586,In_396,In_1481);
nor U1587 (N_1587,In_1493,In_124);
nor U1588 (N_1588,In_174,In_577);
nor U1589 (N_1589,In_1484,In_508);
nor U1590 (N_1590,In_1473,In_765);
and U1591 (N_1591,In_16,In_566);
nor U1592 (N_1592,In_1261,In_905);
and U1593 (N_1593,In_847,In_803);
or U1594 (N_1594,In_428,In_1261);
or U1595 (N_1595,In_879,In_438);
nor U1596 (N_1596,In_734,In_9);
nand U1597 (N_1597,In_849,In_179);
nor U1598 (N_1598,In_1404,In_546);
or U1599 (N_1599,In_1265,In_679);
nand U1600 (N_1600,In_328,In_348);
and U1601 (N_1601,In_435,In_19);
nor U1602 (N_1602,In_1049,In_176);
and U1603 (N_1603,In_885,In_222);
or U1604 (N_1604,In_682,In_519);
and U1605 (N_1605,In_298,In_963);
nor U1606 (N_1606,In_222,In_787);
or U1607 (N_1607,In_500,In_191);
or U1608 (N_1608,In_1232,In_370);
nor U1609 (N_1609,In_1279,In_1466);
nand U1610 (N_1610,In_1434,In_688);
nor U1611 (N_1611,In_607,In_1309);
nand U1612 (N_1612,In_1249,In_1319);
nand U1613 (N_1613,In_1284,In_985);
or U1614 (N_1614,In_1294,In_911);
nand U1615 (N_1615,In_1256,In_1456);
nor U1616 (N_1616,In_1275,In_291);
and U1617 (N_1617,In_1303,In_36);
nor U1618 (N_1618,In_687,In_480);
nand U1619 (N_1619,In_253,In_564);
and U1620 (N_1620,In_608,In_837);
nor U1621 (N_1621,In_1355,In_722);
and U1622 (N_1622,In_1265,In_359);
nor U1623 (N_1623,In_950,In_187);
or U1624 (N_1624,In_434,In_561);
and U1625 (N_1625,In_72,In_85);
nor U1626 (N_1626,In_1096,In_1316);
or U1627 (N_1627,In_1015,In_929);
or U1628 (N_1628,In_1120,In_1057);
and U1629 (N_1629,In_952,In_60);
or U1630 (N_1630,In_51,In_1067);
or U1631 (N_1631,In_1323,In_936);
and U1632 (N_1632,In_1174,In_50);
and U1633 (N_1633,In_1218,In_339);
nor U1634 (N_1634,In_507,In_641);
nand U1635 (N_1635,In_695,In_1347);
nand U1636 (N_1636,In_326,In_1245);
or U1637 (N_1637,In_203,In_631);
nand U1638 (N_1638,In_1218,In_608);
and U1639 (N_1639,In_665,In_299);
and U1640 (N_1640,In_409,In_1033);
xor U1641 (N_1641,In_675,In_1310);
and U1642 (N_1642,In_221,In_621);
and U1643 (N_1643,In_15,In_1432);
and U1644 (N_1644,In_1110,In_1184);
or U1645 (N_1645,In_1411,In_1158);
nand U1646 (N_1646,In_671,In_643);
nor U1647 (N_1647,In_977,In_289);
nand U1648 (N_1648,In_1341,In_238);
nor U1649 (N_1649,In_1415,In_518);
nor U1650 (N_1650,In_1384,In_967);
or U1651 (N_1651,In_920,In_475);
nor U1652 (N_1652,In_144,In_799);
nand U1653 (N_1653,In_1218,In_1462);
nor U1654 (N_1654,In_862,In_1419);
nor U1655 (N_1655,In_278,In_1212);
nor U1656 (N_1656,In_462,In_380);
or U1657 (N_1657,In_1173,In_667);
nand U1658 (N_1658,In_35,In_1466);
nand U1659 (N_1659,In_667,In_128);
nand U1660 (N_1660,In_1321,In_1399);
or U1661 (N_1661,In_712,In_1402);
nand U1662 (N_1662,In_1202,In_369);
and U1663 (N_1663,In_1434,In_849);
and U1664 (N_1664,In_1138,In_459);
nand U1665 (N_1665,In_1147,In_1479);
and U1666 (N_1666,In_1245,In_918);
or U1667 (N_1667,In_1459,In_431);
nand U1668 (N_1668,In_869,In_30);
nand U1669 (N_1669,In_985,In_1416);
or U1670 (N_1670,In_273,In_1236);
or U1671 (N_1671,In_1193,In_304);
nand U1672 (N_1672,In_837,In_412);
or U1673 (N_1673,In_1172,In_650);
and U1674 (N_1674,In_650,In_279);
or U1675 (N_1675,In_258,In_1292);
nand U1676 (N_1676,In_350,In_524);
nand U1677 (N_1677,In_641,In_538);
or U1678 (N_1678,In_1292,In_372);
or U1679 (N_1679,In_1263,In_63);
or U1680 (N_1680,In_1335,In_1291);
or U1681 (N_1681,In_1360,In_773);
nor U1682 (N_1682,In_484,In_824);
or U1683 (N_1683,In_1486,In_57);
nand U1684 (N_1684,In_304,In_1063);
and U1685 (N_1685,In_317,In_876);
and U1686 (N_1686,In_398,In_1336);
and U1687 (N_1687,In_555,In_323);
nand U1688 (N_1688,In_1415,In_555);
and U1689 (N_1689,In_1435,In_862);
and U1690 (N_1690,In_1060,In_601);
nor U1691 (N_1691,In_29,In_228);
or U1692 (N_1692,In_1012,In_1480);
or U1693 (N_1693,In_3,In_2);
and U1694 (N_1694,In_1089,In_1084);
and U1695 (N_1695,In_732,In_291);
nand U1696 (N_1696,In_725,In_811);
and U1697 (N_1697,In_1400,In_1488);
xor U1698 (N_1698,In_1451,In_848);
or U1699 (N_1699,In_1426,In_1262);
nor U1700 (N_1700,In_979,In_961);
and U1701 (N_1701,In_485,In_571);
nor U1702 (N_1702,In_594,In_530);
and U1703 (N_1703,In_695,In_1261);
nor U1704 (N_1704,In_847,In_858);
nand U1705 (N_1705,In_291,In_967);
nand U1706 (N_1706,In_214,In_452);
nor U1707 (N_1707,In_152,In_385);
nand U1708 (N_1708,In_586,In_790);
nor U1709 (N_1709,In_1156,In_1185);
or U1710 (N_1710,In_1128,In_307);
and U1711 (N_1711,In_724,In_1435);
or U1712 (N_1712,In_699,In_151);
or U1713 (N_1713,In_751,In_1407);
and U1714 (N_1714,In_1049,In_1232);
or U1715 (N_1715,In_1189,In_1392);
xor U1716 (N_1716,In_160,In_176);
nand U1717 (N_1717,In_392,In_68);
and U1718 (N_1718,In_1122,In_34);
or U1719 (N_1719,In_46,In_618);
nor U1720 (N_1720,In_159,In_821);
nand U1721 (N_1721,In_57,In_897);
nor U1722 (N_1722,In_1024,In_526);
nor U1723 (N_1723,In_779,In_520);
or U1724 (N_1724,In_86,In_1455);
or U1725 (N_1725,In_1154,In_123);
or U1726 (N_1726,In_1113,In_511);
nand U1727 (N_1727,In_872,In_1387);
nand U1728 (N_1728,In_481,In_1285);
nor U1729 (N_1729,In_739,In_962);
and U1730 (N_1730,In_1194,In_777);
or U1731 (N_1731,In_560,In_1313);
and U1732 (N_1732,In_1450,In_1226);
nor U1733 (N_1733,In_269,In_1416);
or U1734 (N_1734,In_539,In_1094);
or U1735 (N_1735,In_742,In_377);
and U1736 (N_1736,In_743,In_261);
nand U1737 (N_1737,In_367,In_806);
or U1738 (N_1738,In_625,In_1081);
xor U1739 (N_1739,In_1211,In_794);
nor U1740 (N_1740,In_187,In_1218);
nand U1741 (N_1741,In_315,In_1083);
nand U1742 (N_1742,In_925,In_162);
and U1743 (N_1743,In_963,In_1112);
and U1744 (N_1744,In_968,In_554);
and U1745 (N_1745,In_164,In_222);
or U1746 (N_1746,In_559,In_630);
or U1747 (N_1747,In_1348,In_398);
and U1748 (N_1748,In_923,In_1125);
nor U1749 (N_1749,In_753,In_929);
xor U1750 (N_1750,In_848,In_1351);
and U1751 (N_1751,In_1454,In_9);
nor U1752 (N_1752,In_485,In_94);
nor U1753 (N_1753,In_1058,In_274);
nand U1754 (N_1754,In_134,In_537);
nor U1755 (N_1755,In_23,In_731);
and U1756 (N_1756,In_376,In_861);
nand U1757 (N_1757,In_670,In_515);
nand U1758 (N_1758,In_1188,In_1249);
nor U1759 (N_1759,In_484,In_1278);
or U1760 (N_1760,In_880,In_1426);
nand U1761 (N_1761,In_595,In_446);
or U1762 (N_1762,In_1146,In_1358);
or U1763 (N_1763,In_977,In_1431);
nor U1764 (N_1764,In_445,In_503);
and U1765 (N_1765,In_92,In_86);
and U1766 (N_1766,In_563,In_1247);
nand U1767 (N_1767,In_102,In_1247);
nor U1768 (N_1768,In_1422,In_103);
or U1769 (N_1769,In_61,In_626);
nor U1770 (N_1770,In_1275,In_518);
or U1771 (N_1771,In_581,In_145);
nand U1772 (N_1772,In_875,In_100);
nand U1773 (N_1773,In_685,In_1454);
and U1774 (N_1774,In_763,In_946);
and U1775 (N_1775,In_673,In_1221);
and U1776 (N_1776,In_1132,In_705);
and U1777 (N_1777,In_1450,In_767);
nand U1778 (N_1778,In_632,In_284);
or U1779 (N_1779,In_799,In_310);
nor U1780 (N_1780,In_306,In_1473);
nand U1781 (N_1781,In_980,In_1421);
and U1782 (N_1782,In_1001,In_180);
and U1783 (N_1783,In_849,In_1157);
and U1784 (N_1784,In_382,In_1190);
and U1785 (N_1785,In_740,In_1018);
or U1786 (N_1786,In_497,In_371);
nand U1787 (N_1787,In_515,In_414);
nor U1788 (N_1788,In_558,In_1072);
nor U1789 (N_1789,In_1359,In_256);
or U1790 (N_1790,In_972,In_1018);
and U1791 (N_1791,In_651,In_690);
nand U1792 (N_1792,In_306,In_117);
or U1793 (N_1793,In_504,In_1195);
or U1794 (N_1794,In_1264,In_710);
nand U1795 (N_1795,In_654,In_967);
and U1796 (N_1796,In_1241,In_48);
nand U1797 (N_1797,In_1480,In_1426);
nor U1798 (N_1798,In_310,In_1234);
nor U1799 (N_1799,In_1158,In_163);
nand U1800 (N_1800,In_1163,In_587);
and U1801 (N_1801,In_725,In_108);
and U1802 (N_1802,In_463,In_1464);
or U1803 (N_1803,In_1023,In_238);
nor U1804 (N_1804,In_1467,In_99);
nand U1805 (N_1805,In_216,In_1231);
and U1806 (N_1806,In_48,In_192);
nor U1807 (N_1807,In_451,In_532);
and U1808 (N_1808,In_501,In_773);
nand U1809 (N_1809,In_519,In_1493);
or U1810 (N_1810,In_844,In_851);
nor U1811 (N_1811,In_1039,In_1231);
nand U1812 (N_1812,In_1177,In_612);
nand U1813 (N_1813,In_310,In_400);
nor U1814 (N_1814,In_1241,In_1222);
or U1815 (N_1815,In_1269,In_383);
xor U1816 (N_1816,In_1327,In_264);
and U1817 (N_1817,In_544,In_531);
nand U1818 (N_1818,In_414,In_220);
xor U1819 (N_1819,In_1452,In_186);
nand U1820 (N_1820,In_157,In_963);
and U1821 (N_1821,In_310,In_990);
or U1822 (N_1822,In_354,In_289);
nand U1823 (N_1823,In_969,In_547);
nor U1824 (N_1824,In_1370,In_1368);
nor U1825 (N_1825,In_107,In_1251);
and U1826 (N_1826,In_503,In_1057);
nand U1827 (N_1827,In_259,In_1246);
nor U1828 (N_1828,In_428,In_1058);
and U1829 (N_1829,In_139,In_1471);
nand U1830 (N_1830,In_1105,In_1343);
nand U1831 (N_1831,In_1020,In_823);
and U1832 (N_1832,In_447,In_99);
nand U1833 (N_1833,In_1255,In_179);
xnor U1834 (N_1834,In_1440,In_43);
or U1835 (N_1835,In_911,In_189);
nand U1836 (N_1836,In_42,In_1086);
nor U1837 (N_1837,In_62,In_1400);
and U1838 (N_1838,In_361,In_292);
and U1839 (N_1839,In_659,In_1444);
or U1840 (N_1840,In_1284,In_1115);
nor U1841 (N_1841,In_1113,In_903);
nand U1842 (N_1842,In_619,In_1476);
nand U1843 (N_1843,In_1011,In_273);
nand U1844 (N_1844,In_672,In_1126);
nand U1845 (N_1845,In_1196,In_1414);
and U1846 (N_1846,In_537,In_255);
nor U1847 (N_1847,In_1170,In_1351);
and U1848 (N_1848,In_838,In_1247);
nand U1849 (N_1849,In_1111,In_1194);
nor U1850 (N_1850,In_248,In_831);
and U1851 (N_1851,In_634,In_1122);
nor U1852 (N_1852,In_1139,In_1312);
or U1853 (N_1853,In_821,In_445);
or U1854 (N_1854,In_979,In_660);
or U1855 (N_1855,In_1233,In_89);
nor U1856 (N_1856,In_1030,In_1132);
nor U1857 (N_1857,In_323,In_542);
nor U1858 (N_1858,In_531,In_796);
or U1859 (N_1859,In_575,In_1283);
and U1860 (N_1860,In_1125,In_756);
or U1861 (N_1861,In_802,In_1446);
and U1862 (N_1862,In_1265,In_1313);
nor U1863 (N_1863,In_654,In_1091);
nand U1864 (N_1864,In_1438,In_405);
nor U1865 (N_1865,In_967,In_812);
nor U1866 (N_1866,In_127,In_204);
or U1867 (N_1867,In_129,In_1487);
nor U1868 (N_1868,In_388,In_31);
and U1869 (N_1869,In_648,In_160);
and U1870 (N_1870,In_275,In_1087);
nor U1871 (N_1871,In_130,In_1463);
or U1872 (N_1872,In_983,In_758);
nor U1873 (N_1873,In_391,In_954);
or U1874 (N_1874,In_338,In_890);
nor U1875 (N_1875,In_761,In_1057);
and U1876 (N_1876,In_640,In_383);
and U1877 (N_1877,In_1361,In_1086);
or U1878 (N_1878,In_618,In_316);
and U1879 (N_1879,In_912,In_299);
nand U1880 (N_1880,In_657,In_227);
and U1881 (N_1881,In_255,In_1147);
nand U1882 (N_1882,In_600,In_519);
or U1883 (N_1883,In_866,In_824);
or U1884 (N_1884,In_1487,In_1101);
or U1885 (N_1885,In_923,In_190);
nor U1886 (N_1886,In_926,In_665);
and U1887 (N_1887,In_981,In_746);
and U1888 (N_1888,In_1204,In_1258);
nor U1889 (N_1889,In_348,In_1099);
or U1890 (N_1890,In_15,In_128);
and U1891 (N_1891,In_964,In_1268);
nand U1892 (N_1892,In_1338,In_1139);
nor U1893 (N_1893,In_1412,In_271);
and U1894 (N_1894,In_481,In_779);
nand U1895 (N_1895,In_1111,In_310);
nor U1896 (N_1896,In_687,In_767);
or U1897 (N_1897,In_1280,In_763);
nor U1898 (N_1898,In_792,In_1399);
and U1899 (N_1899,In_331,In_461);
nor U1900 (N_1900,In_323,In_783);
nor U1901 (N_1901,In_481,In_1143);
nor U1902 (N_1902,In_195,In_722);
and U1903 (N_1903,In_408,In_926);
nor U1904 (N_1904,In_1142,In_122);
xor U1905 (N_1905,In_462,In_38);
nor U1906 (N_1906,In_249,In_1151);
nand U1907 (N_1907,In_327,In_1070);
nand U1908 (N_1908,In_579,In_1062);
or U1909 (N_1909,In_659,In_1356);
nor U1910 (N_1910,In_701,In_535);
xor U1911 (N_1911,In_4,In_599);
or U1912 (N_1912,In_84,In_965);
or U1913 (N_1913,In_291,In_1408);
or U1914 (N_1914,In_11,In_548);
nor U1915 (N_1915,In_1499,In_910);
nand U1916 (N_1916,In_339,In_852);
and U1917 (N_1917,In_562,In_1416);
nor U1918 (N_1918,In_308,In_960);
nor U1919 (N_1919,In_852,In_102);
nand U1920 (N_1920,In_313,In_66);
nand U1921 (N_1921,In_349,In_692);
nor U1922 (N_1922,In_743,In_813);
xnor U1923 (N_1923,In_938,In_399);
or U1924 (N_1924,In_482,In_721);
nor U1925 (N_1925,In_752,In_323);
nand U1926 (N_1926,In_728,In_313);
and U1927 (N_1927,In_997,In_141);
nor U1928 (N_1928,In_393,In_1346);
nand U1929 (N_1929,In_985,In_1178);
nor U1930 (N_1930,In_1254,In_225);
and U1931 (N_1931,In_1325,In_743);
nor U1932 (N_1932,In_903,In_190);
nand U1933 (N_1933,In_954,In_911);
and U1934 (N_1934,In_290,In_894);
and U1935 (N_1935,In_919,In_409);
nand U1936 (N_1936,In_1370,In_888);
and U1937 (N_1937,In_1463,In_1352);
nor U1938 (N_1938,In_1010,In_1095);
and U1939 (N_1939,In_908,In_1311);
or U1940 (N_1940,In_347,In_237);
and U1941 (N_1941,In_980,In_253);
nor U1942 (N_1942,In_116,In_1307);
or U1943 (N_1943,In_1061,In_1407);
nor U1944 (N_1944,In_1166,In_843);
and U1945 (N_1945,In_343,In_1367);
nand U1946 (N_1946,In_1025,In_1014);
and U1947 (N_1947,In_416,In_337);
nand U1948 (N_1948,In_1299,In_327);
nand U1949 (N_1949,In_1318,In_600);
and U1950 (N_1950,In_125,In_1368);
or U1951 (N_1951,In_845,In_905);
and U1952 (N_1952,In_725,In_485);
nor U1953 (N_1953,In_943,In_683);
and U1954 (N_1954,In_210,In_605);
nand U1955 (N_1955,In_1053,In_1490);
nand U1956 (N_1956,In_1022,In_1492);
nand U1957 (N_1957,In_561,In_1079);
nor U1958 (N_1958,In_1471,In_9);
nand U1959 (N_1959,In_996,In_872);
nand U1960 (N_1960,In_1006,In_1063);
and U1961 (N_1961,In_1267,In_218);
or U1962 (N_1962,In_98,In_1049);
nand U1963 (N_1963,In_123,In_997);
nor U1964 (N_1964,In_100,In_47);
and U1965 (N_1965,In_996,In_271);
or U1966 (N_1966,In_470,In_205);
and U1967 (N_1967,In_228,In_155);
or U1968 (N_1968,In_783,In_835);
nor U1969 (N_1969,In_19,In_932);
nand U1970 (N_1970,In_1290,In_1030);
nor U1971 (N_1971,In_16,In_1127);
nor U1972 (N_1972,In_716,In_727);
and U1973 (N_1973,In_648,In_1006);
nor U1974 (N_1974,In_105,In_900);
nand U1975 (N_1975,In_720,In_1012);
nor U1976 (N_1976,In_1087,In_1067);
or U1977 (N_1977,In_474,In_723);
and U1978 (N_1978,In_1059,In_1164);
or U1979 (N_1979,In_1198,In_34);
nand U1980 (N_1980,In_107,In_1347);
nor U1981 (N_1981,In_1260,In_333);
or U1982 (N_1982,In_899,In_640);
nor U1983 (N_1983,In_41,In_301);
or U1984 (N_1984,In_91,In_707);
xnor U1985 (N_1985,In_1271,In_258);
nor U1986 (N_1986,In_904,In_1156);
nand U1987 (N_1987,In_1480,In_1489);
or U1988 (N_1988,In_870,In_1155);
nand U1989 (N_1989,In_282,In_1292);
and U1990 (N_1990,In_659,In_1408);
or U1991 (N_1991,In_784,In_1181);
nor U1992 (N_1992,In_1007,In_440);
or U1993 (N_1993,In_1346,In_646);
or U1994 (N_1994,In_722,In_1340);
nor U1995 (N_1995,In_674,In_1012);
nor U1996 (N_1996,In_1237,In_1010);
and U1997 (N_1997,In_1486,In_116);
nor U1998 (N_1998,In_520,In_513);
nand U1999 (N_1999,In_278,In_694);
nand U2000 (N_2000,In_815,In_1315);
or U2001 (N_2001,In_1099,In_83);
nor U2002 (N_2002,In_627,In_783);
and U2003 (N_2003,In_260,In_1122);
or U2004 (N_2004,In_501,In_343);
or U2005 (N_2005,In_996,In_405);
nand U2006 (N_2006,In_1277,In_1363);
nand U2007 (N_2007,In_951,In_1015);
nand U2008 (N_2008,In_835,In_1488);
nand U2009 (N_2009,In_1187,In_960);
and U2010 (N_2010,In_887,In_129);
and U2011 (N_2011,In_304,In_783);
or U2012 (N_2012,In_962,In_1418);
or U2013 (N_2013,In_721,In_303);
or U2014 (N_2014,In_658,In_746);
or U2015 (N_2015,In_60,In_1146);
or U2016 (N_2016,In_1241,In_899);
and U2017 (N_2017,In_663,In_972);
and U2018 (N_2018,In_678,In_835);
nand U2019 (N_2019,In_40,In_284);
nor U2020 (N_2020,In_670,In_37);
nand U2021 (N_2021,In_1142,In_1419);
nand U2022 (N_2022,In_752,In_1238);
nand U2023 (N_2023,In_1141,In_959);
or U2024 (N_2024,In_1246,In_279);
and U2025 (N_2025,In_1377,In_758);
and U2026 (N_2026,In_342,In_1399);
nor U2027 (N_2027,In_904,In_45);
and U2028 (N_2028,In_16,In_657);
nand U2029 (N_2029,In_1310,In_413);
nand U2030 (N_2030,In_947,In_1245);
or U2031 (N_2031,In_1053,In_1465);
nand U2032 (N_2032,In_173,In_1499);
and U2033 (N_2033,In_1472,In_626);
nand U2034 (N_2034,In_936,In_102);
nor U2035 (N_2035,In_685,In_1469);
nand U2036 (N_2036,In_763,In_1198);
nor U2037 (N_2037,In_765,In_994);
nor U2038 (N_2038,In_1310,In_929);
or U2039 (N_2039,In_168,In_767);
or U2040 (N_2040,In_131,In_614);
nand U2041 (N_2041,In_111,In_465);
nor U2042 (N_2042,In_1155,In_694);
nor U2043 (N_2043,In_953,In_1214);
nor U2044 (N_2044,In_136,In_486);
and U2045 (N_2045,In_868,In_1196);
or U2046 (N_2046,In_1202,In_487);
and U2047 (N_2047,In_476,In_599);
nand U2048 (N_2048,In_314,In_1306);
xnor U2049 (N_2049,In_877,In_608);
or U2050 (N_2050,In_1310,In_1454);
and U2051 (N_2051,In_932,In_1197);
or U2052 (N_2052,In_221,In_930);
or U2053 (N_2053,In_720,In_1414);
nand U2054 (N_2054,In_101,In_362);
and U2055 (N_2055,In_812,In_487);
nor U2056 (N_2056,In_846,In_587);
or U2057 (N_2057,In_863,In_831);
and U2058 (N_2058,In_1028,In_308);
or U2059 (N_2059,In_51,In_828);
and U2060 (N_2060,In_766,In_328);
nand U2061 (N_2061,In_330,In_1112);
or U2062 (N_2062,In_876,In_371);
nor U2063 (N_2063,In_283,In_1001);
nand U2064 (N_2064,In_46,In_797);
nand U2065 (N_2065,In_157,In_133);
or U2066 (N_2066,In_541,In_593);
or U2067 (N_2067,In_1420,In_1031);
and U2068 (N_2068,In_266,In_1464);
nand U2069 (N_2069,In_316,In_227);
and U2070 (N_2070,In_396,In_701);
or U2071 (N_2071,In_91,In_247);
nor U2072 (N_2072,In_1245,In_1221);
nor U2073 (N_2073,In_1337,In_560);
nand U2074 (N_2074,In_83,In_209);
nand U2075 (N_2075,In_309,In_178);
and U2076 (N_2076,In_1176,In_1081);
nor U2077 (N_2077,In_4,In_706);
nand U2078 (N_2078,In_363,In_954);
and U2079 (N_2079,In_1462,In_871);
and U2080 (N_2080,In_586,In_1296);
nand U2081 (N_2081,In_1100,In_810);
nand U2082 (N_2082,In_982,In_176);
and U2083 (N_2083,In_1302,In_445);
nand U2084 (N_2084,In_154,In_1217);
nand U2085 (N_2085,In_1185,In_80);
or U2086 (N_2086,In_350,In_687);
xor U2087 (N_2087,In_755,In_564);
and U2088 (N_2088,In_498,In_1411);
nor U2089 (N_2089,In_350,In_1028);
nor U2090 (N_2090,In_11,In_724);
or U2091 (N_2091,In_195,In_408);
nor U2092 (N_2092,In_713,In_90);
nor U2093 (N_2093,In_997,In_578);
nor U2094 (N_2094,In_892,In_1138);
nor U2095 (N_2095,In_1282,In_656);
or U2096 (N_2096,In_1225,In_1063);
nor U2097 (N_2097,In_1273,In_1223);
or U2098 (N_2098,In_14,In_1280);
or U2099 (N_2099,In_1033,In_1198);
and U2100 (N_2100,In_846,In_1048);
nor U2101 (N_2101,In_1377,In_286);
nand U2102 (N_2102,In_1157,In_1111);
and U2103 (N_2103,In_641,In_763);
and U2104 (N_2104,In_620,In_538);
nand U2105 (N_2105,In_7,In_334);
or U2106 (N_2106,In_1357,In_1011);
and U2107 (N_2107,In_1445,In_1212);
nand U2108 (N_2108,In_1494,In_358);
nand U2109 (N_2109,In_629,In_444);
or U2110 (N_2110,In_587,In_632);
or U2111 (N_2111,In_442,In_1221);
nand U2112 (N_2112,In_275,In_146);
nor U2113 (N_2113,In_308,In_682);
or U2114 (N_2114,In_287,In_1139);
nand U2115 (N_2115,In_472,In_110);
nor U2116 (N_2116,In_407,In_808);
or U2117 (N_2117,In_1279,In_524);
nand U2118 (N_2118,In_407,In_1253);
and U2119 (N_2119,In_1083,In_247);
nand U2120 (N_2120,In_203,In_68);
nand U2121 (N_2121,In_1003,In_1415);
and U2122 (N_2122,In_859,In_483);
and U2123 (N_2123,In_579,In_188);
xor U2124 (N_2124,In_580,In_704);
nand U2125 (N_2125,In_924,In_1352);
nor U2126 (N_2126,In_1461,In_1310);
nand U2127 (N_2127,In_1071,In_649);
or U2128 (N_2128,In_1046,In_1105);
or U2129 (N_2129,In_1032,In_883);
nand U2130 (N_2130,In_756,In_781);
xor U2131 (N_2131,In_242,In_597);
or U2132 (N_2132,In_35,In_1355);
nand U2133 (N_2133,In_860,In_588);
nor U2134 (N_2134,In_1307,In_442);
xnor U2135 (N_2135,In_117,In_435);
or U2136 (N_2136,In_1056,In_1376);
nand U2137 (N_2137,In_311,In_686);
or U2138 (N_2138,In_173,In_408);
nand U2139 (N_2139,In_1186,In_1120);
nand U2140 (N_2140,In_541,In_834);
or U2141 (N_2141,In_289,In_1309);
xor U2142 (N_2142,In_1177,In_780);
nor U2143 (N_2143,In_1347,In_782);
or U2144 (N_2144,In_1206,In_277);
or U2145 (N_2145,In_532,In_142);
nand U2146 (N_2146,In_379,In_700);
or U2147 (N_2147,In_1061,In_942);
and U2148 (N_2148,In_1371,In_1498);
nor U2149 (N_2149,In_763,In_1091);
and U2150 (N_2150,In_453,In_32);
and U2151 (N_2151,In_1445,In_1357);
nor U2152 (N_2152,In_303,In_266);
nand U2153 (N_2153,In_745,In_1095);
nand U2154 (N_2154,In_72,In_512);
nand U2155 (N_2155,In_1499,In_169);
nand U2156 (N_2156,In_721,In_898);
nand U2157 (N_2157,In_1072,In_486);
nor U2158 (N_2158,In_5,In_63);
or U2159 (N_2159,In_39,In_444);
and U2160 (N_2160,In_562,In_1307);
nand U2161 (N_2161,In_1399,In_111);
nor U2162 (N_2162,In_455,In_649);
nand U2163 (N_2163,In_1048,In_576);
and U2164 (N_2164,In_1282,In_1023);
nand U2165 (N_2165,In_791,In_192);
or U2166 (N_2166,In_235,In_1065);
or U2167 (N_2167,In_1110,In_1284);
nand U2168 (N_2168,In_14,In_1242);
xnor U2169 (N_2169,In_917,In_174);
nand U2170 (N_2170,In_19,In_341);
nor U2171 (N_2171,In_648,In_830);
nor U2172 (N_2172,In_287,In_764);
or U2173 (N_2173,In_820,In_27);
nor U2174 (N_2174,In_765,In_18);
and U2175 (N_2175,In_1032,In_699);
nor U2176 (N_2176,In_1423,In_1006);
nand U2177 (N_2177,In_363,In_1483);
nand U2178 (N_2178,In_13,In_1145);
xnor U2179 (N_2179,In_1016,In_638);
nand U2180 (N_2180,In_1295,In_480);
or U2181 (N_2181,In_924,In_13);
nor U2182 (N_2182,In_1125,In_467);
and U2183 (N_2183,In_629,In_1158);
nor U2184 (N_2184,In_1406,In_1207);
nor U2185 (N_2185,In_460,In_1257);
nand U2186 (N_2186,In_1330,In_1006);
nor U2187 (N_2187,In_1118,In_1029);
and U2188 (N_2188,In_422,In_1313);
and U2189 (N_2189,In_522,In_1129);
nand U2190 (N_2190,In_1300,In_757);
nand U2191 (N_2191,In_383,In_356);
and U2192 (N_2192,In_1389,In_1300);
and U2193 (N_2193,In_733,In_615);
nor U2194 (N_2194,In_257,In_1358);
and U2195 (N_2195,In_13,In_622);
or U2196 (N_2196,In_326,In_690);
nor U2197 (N_2197,In_399,In_670);
and U2198 (N_2198,In_916,In_1203);
and U2199 (N_2199,In_982,In_650);
and U2200 (N_2200,In_976,In_449);
nand U2201 (N_2201,In_877,In_1236);
or U2202 (N_2202,In_476,In_1047);
and U2203 (N_2203,In_783,In_206);
nand U2204 (N_2204,In_1219,In_591);
nand U2205 (N_2205,In_921,In_673);
nor U2206 (N_2206,In_686,In_1386);
nor U2207 (N_2207,In_138,In_1219);
xor U2208 (N_2208,In_1048,In_331);
nor U2209 (N_2209,In_646,In_727);
nor U2210 (N_2210,In_182,In_1328);
xnor U2211 (N_2211,In_1293,In_369);
nor U2212 (N_2212,In_431,In_220);
nand U2213 (N_2213,In_50,In_957);
xor U2214 (N_2214,In_1362,In_133);
and U2215 (N_2215,In_1295,In_749);
and U2216 (N_2216,In_1093,In_1424);
nand U2217 (N_2217,In_1292,In_432);
nor U2218 (N_2218,In_1287,In_1201);
nand U2219 (N_2219,In_370,In_1371);
and U2220 (N_2220,In_223,In_1362);
nand U2221 (N_2221,In_435,In_1312);
and U2222 (N_2222,In_724,In_344);
and U2223 (N_2223,In_160,In_1229);
nor U2224 (N_2224,In_1140,In_151);
and U2225 (N_2225,In_1344,In_527);
or U2226 (N_2226,In_1098,In_1216);
nand U2227 (N_2227,In_716,In_381);
nand U2228 (N_2228,In_1031,In_1116);
and U2229 (N_2229,In_1454,In_1128);
or U2230 (N_2230,In_1307,In_1498);
or U2231 (N_2231,In_938,In_1337);
and U2232 (N_2232,In_1200,In_1169);
and U2233 (N_2233,In_402,In_1383);
nand U2234 (N_2234,In_955,In_632);
xnor U2235 (N_2235,In_510,In_419);
or U2236 (N_2236,In_1118,In_1081);
or U2237 (N_2237,In_45,In_1317);
or U2238 (N_2238,In_1231,In_271);
nand U2239 (N_2239,In_937,In_156);
or U2240 (N_2240,In_1306,In_39);
nor U2241 (N_2241,In_1024,In_105);
or U2242 (N_2242,In_1200,In_71);
nand U2243 (N_2243,In_23,In_966);
or U2244 (N_2244,In_824,In_1410);
nor U2245 (N_2245,In_1266,In_334);
nor U2246 (N_2246,In_105,In_294);
nor U2247 (N_2247,In_482,In_668);
nor U2248 (N_2248,In_930,In_43);
or U2249 (N_2249,In_7,In_460);
nor U2250 (N_2250,In_1313,In_763);
nand U2251 (N_2251,In_1383,In_288);
nand U2252 (N_2252,In_1432,In_1062);
nor U2253 (N_2253,In_818,In_127);
nand U2254 (N_2254,In_873,In_544);
xnor U2255 (N_2255,In_1450,In_179);
and U2256 (N_2256,In_1493,In_1148);
and U2257 (N_2257,In_1380,In_338);
nand U2258 (N_2258,In_1283,In_1327);
nor U2259 (N_2259,In_1194,In_196);
nand U2260 (N_2260,In_1261,In_1119);
nor U2261 (N_2261,In_935,In_1299);
nor U2262 (N_2262,In_187,In_229);
nand U2263 (N_2263,In_307,In_564);
nand U2264 (N_2264,In_667,In_1125);
nor U2265 (N_2265,In_1403,In_324);
or U2266 (N_2266,In_1120,In_1448);
and U2267 (N_2267,In_149,In_1341);
or U2268 (N_2268,In_450,In_1329);
and U2269 (N_2269,In_441,In_1436);
nor U2270 (N_2270,In_534,In_1076);
and U2271 (N_2271,In_639,In_617);
nor U2272 (N_2272,In_668,In_1265);
nor U2273 (N_2273,In_435,In_358);
nor U2274 (N_2274,In_483,In_986);
and U2275 (N_2275,In_813,In_1013);
and U2276 (N_2276,In_258,In_1199);
or U2277 (N_2277,In_300,In_206);
and U2278 (N_2278,In_1090,In_604);
and U2279 (N_2279,In_400,In_1099);
nor U2280 (N_2280,In_755,In_872);
and U2281 (N_2281,In_677,In_645);
nor U2282 (N_2282,In_1001,In_782);
and U2283 (N_2283,In_181,In_1249);
and U2284 (N_2284,In_14,In_466);
or U2285 (N_2285,In_1277,In_422);
or U2286 (N_2286,In_1267,In_1383);
or U2287 (N_2287,In_501,In_226);
or U2288 (N_2288,In_995,In_417);
or U2289 (N_2289,In_1171,In_300);
xor U2290 (N_2290,In_70,In_399);
nor U2291 (N_2291,In_243,In_1054);
or U2292 (N_2292,In_346,In_871);
nor U2293 (N_2293,In_1123,In_121);
nand U2294 (N_2294,In_1476,In_1359);
nand U2295 (N_2295,In_1306,In_414);
and U2296 (N_2296,In_43,In_554);
and U2297 (N_2297,In_669,In_1494);
nand U2298 (N_2298,In_1279,In_948);
and U2299 (N_2299,In_1443,In_300);
nand U2300 (N_2300,In_1134,In_246);
nand U2301 (N_2301,In_267,In_1064);
or U2302 (N_2302,In_760,In_412);
nand U2303 (N_2303,In_637,In_819);
and U2304 (N_2304,In_1207,In_6);
nor U2305 (N_2305,In_744,In_530);
nand U2306 (N_2306,In_823,In_349);
nand U2307 (N_2307,In_972,In_169);
nor U2308 (N_2308,In_1013,In_1490);
nor U2309 (N_2309,In_384,In_271);
nor U2310 (N_2310,In_1350,In_640);
nor U2311 (N_2311,In_253,In_1111);
xnor U2312 (N_2312,In_874,In_1230);
nor U2313 (N_2313,In_1366,In_180);
xnor U2314 (N_2314,In_1051,In_1196);
nand U2315 (N_2315,In_1052,In_595);
and U2316 (N_2316,In_575,In_374);
nor U2317 (N_2317,In_659,In_510);
or U2318 (N_2318,In_241,In_1279);
nor U2319 (N_2319,In_1106,In_458);
and U2320 (N_2320,In_596,In_1092);
and U2321 (N_2321,In_1162,In_797);
xnor U2322 (N_2322,In_1476,In_11);
nand U2323 (N_2323,In_686,In_1362);
or U2324 (N_2324,In_178,In_67);
or U2325 (N_2325,In_873,In_445);
nand U2326 (N_2326,In_572,In_1191);
nand U2327 (N_2327,In_971,In_564);
and U2328 (N_2328,In_1329,In_147);
or U2329 (N_2329,In_1373,In_856);
or U2330 (N_2330,In_1049,In_213);
and U2331 (N_2331,In_598,In_1034);
nor U2332 (N_2332,In_1314,In_473);
and U2333 (N_2333,In_1,In_1360);
or U2334 (N_2334,In_1319,In_511);
and U2335 (N_2335,In_779,In_922);
nand U2336 (N_2336,In_490,In_583);
nor U2337 (N_2337,In_624,In_1145);
xnor U2338 (N_2338,In_1163,In_436);
xnor U2339 (N_2339,In_348,In_763);
xnor U2340 (N_2340,In_964,In_788);
nor U2341 (N_2341,In_423,In_397);
or U2342 (N_2342,In_1236,In_768);
or U2343 (N_2343,In_467,In_835);
and U2344 (N_2344,In_1453,In_1084);
and U2345 (N_2345,In_1491,In_1330);
nor U2346 (N_2346,In_645,In_1385);
nor U2347 (N_2347,In_886,In_527);
or U2348 (N_2348,In_131,In_597);
or U2349 (N_2349,In_852,In_317);
and U2350 (N_2350,In_0,In_364);
or U2351 (N_2351,In_982,In_69);
and U2352 (N_2352,In_1355,In_1294);
nor U2353 (N_2353,In_1193,In_248);
nor U2354 (N_2354,In_973,In_453);
and U2355 (N_2355,In_1048,In_355);
nand U2356 (N_2356,In_962,In_745);
nand U2357 (N_2357,In_286,In_972);
or U2358 (N_2358,In_335,In_754);
or U2359 (N_2359,In_797,In_1030);
nor U2360 (N_2360,In_332,In_796);
nor U2361 (N_2361,In_1031,In_664);
and U2362 (N_2362,In_1294,In_219);
or U2363 (N_2363,In_2,In_996);
and U2364 (N_2364,In_1039,In_1410);
or U2365 (N_2365,In_1443,In_1358);
or U2366 (N_2366,In_1221,In_422);
and U2367 (N_2367,In_289,In_1173);
nor U2368 (N_2368,In_207,In_561);
or U2369 (N_2369,In_356,In_876);
or U2370 (N_2370,In_1476,In_1448);
nand U2371 (N_2371,In_1326,In_929);
or U2372 (N_2372,In_70,In_765);
nand U2373 (N_2373,In_178,In_1223);
nand U2374 (N_2374,In_918,In_1412);
xnor U2375 (N_2375,In_1019,In_1227);
and U2376 (N_2376,In_156,In_820);
or U2377 (N_2377,In_863,In_1382);
and U2378 (N_2378,In_37,In_575);
and U2379 (N_2379,In_1403,In_128);
or U2380 (N_2380,In_134,In_674);
nand U2381 (N_2381,In_1064,In_725);
and U2382 (N_2382,In_119,In_1344);
or U2383 (N_2383,In_526,In_684);
nor U2384 (N_2384,In_1478,In_766);
nor U2385 (N_2385,In_52,In_353);
or U2386 (N_2386,In_300,In_260);
nor U2387 (N_2387,In_571,In_157);
nand U2388 (N_2388,In_445,In_254);
and U2389 (N_2389,In_808,In_241);
nor U2390 (N_2390,In_97,In_1205);
and U2391 (N_2391,In_970,In_938);
xor U2392 (N_2392,In_906,In_1447);
nor U2393 (N_2393,In_541,In_84);
nor U2394 (N_2394,In_653,In_1151);
nand U2395 (N_2395,In_296,In_1227);
or U2396 (N_2396,In_1364,In_1207);
or U2397 (N_2397,In_1362,In_1364);
nand U2398 (N_2398,In_1371,In_114);
nor U2399 (N_2399,In_923,In_850);
nand U2400 (N_2400,In_63,In_698);
or U2401 (N_2401,In_1248,In_935);
nor U2402 (N_2402,In_313,In_528);
and U2403 (N_2403,In_1028,In_132);
nand U2404 (N_2404,In_183,In_294);
and U2405 (N_2405,In_734,In_259);
nand U2406 (N_2406,In_727,In_384);
or U2407 (N_2407,In_314,In_1442);
and U2408 (N_2408,In_875,In_135);
or U2409 (N_2409,In_459,In_375);
or U2410 (N_2410,In_1015,In_335);
or U2411 (N_2411,In_229,In_1155);
or U2412 (N_2412,In_33,In_1457);
and U2413 (N_2413,In_1059,In_854);
and U2414 (N_2414,In_423,In_343);
nand U2415 (N_2415,In_894,In_1071);
or U2416 (N_2416,In_865,In_482);
nand U2417 (N_2417,In_894,In_1331);
xnor U2418 (N_2418,In_819,In_574);
nor U2419 (N_2419,In_887,In_1443);
nand U2420 (N_2420,In_537,In_773);
and U2421 (N_2421,In_549,In_1431);
nand U2422 (N_2422,In_620,In_537);
nand U2423 (N_2423,In_442,In_391);
nor U2424 (N_2424,In_914,In_1499);
or U2425 (N_2425,In_2,In_268);
or U2426 (N_2426,In_1365,In_830);
or U2427 (N_2427,In_59,In_413);
or U2428 (N_2428,In_885,In_1254);
nor U2429 (N_2429,In_1128,In_643);
nor U2430 (N_2430,In_1177,In_222);
or U2431 (N_2431,In_827,In_1088);
or U2432 (N_2432,In_1113,In_346);
or U2433 (N_2433,In_279,In_385);
nand U2434 (N_2434,In_748,In_164);
nand U2435 (N_2435,In_1294,In_533);
nor U2436 (N_2436,In_766,In_960);
nor U2437 (N_2437,In_335,In_1380);
or U2438 (N_2438,In_1005,In_1432);
nand U2439 (N_2439,In_10,In_68);
or U2440 (N_2440,In_299,In_1070);
nor U2441 (N_2441,In_1212,In_1401);
nor U2442 (N_2442,In_758,In_384);
and U2443 (N_2443,In_1090,In_726);
nor U2444 (N_2444,In_1179,In_57);
nor U2445 (N_2445,In_435,In_28);
nand U2446 (N_2446,In_601,In_310);
nand U2447 (N_2447,In_64,In_826);
or U2448 (N_2448,In_868,In_950);
and U2449 (N_2449,In_1135,In_472);
nand U2450 (N_2450,In_1416,In_379);
and U2451 (N_2451,In_1303,In_1454);
nor U2452 (N_2452,In_70,In_230);
and U2453 (N_2453,In_1197,In_1014);
nand U2454 (N_2454,In_54,In_407);
or U2455 (N_2455,In_1300,In_919);
nor U2456 (N_2456,In_1312,In_333);
nand U2457 (N_2457,In_49,In_96);
or U2458 (N_2458,In_914,In_212);
nand U2459 (N_2459,In_500,In_1348);
nor U2460 (N_2460,In_189,In_1353);
or U2461 (N_2461,In_971,In_1360);
nor U2462 (N_2462,In_712,In_1479);
nor U2463 (N_2463,In_473,In_320);
nand U2464 (N_2464,In_118,In_604);
and U2465 (N_2465,In_1402,In_470);
nor U2466 (N_2466,In_1177,In_1041);
nand U2467 (N_2467,In_951,In_635);
and U2468 (N_2468,In_1065,In_1372);
nand U2469 (N_2469,In_1000,In_303);
nor U2470 (N_2470,In_1310,In_230);
nor U2471 (N_2471,In_893,In_49);
nor U2472 (N_2472,In_1353,In_506);
nor U2473 (N_2473,In_96,In_475);
nand U2474 (N_2474,In_634,In_860);
nand U2475 (N_2475,In_439,In_934);
nor U2476 (N_2476,In_183,In_0);
and U2477 (N_2477,In_1261,In_1181);
and U2478 (N_2478,In_1115,In_964);
nand U2479 (N_2479,In_1030,In_903);
or U2480 (N_2480,In_876,In_301);
nor U2481 (N_2481,In_885,In_1460);
xor U2482 (N_2482,In_106,In_1400);
and U2483 (N_2483,In_168,In_157);
or U2484 (N_2484,In_1333,In_1480);
nand U2485 (N_2485,In_868,In_704);
nand U2486 (N_2486,In_504,In_517);
nand U2487 (N_2487,In_176,In_676);
or U2488 (N_2488,In_58,In_1189);
and U2489 (N_2489,In_1328,In_971);
or U2490 (N_2490,In_362,In_282);
nand U2491 (N_2491,In_829,In_291);
nor U2492 (N_2492,In_173,In_814);
nand U2493 (N_2493,In_386,In_131);
xnor U2494 (N_2494,In_1370,In_194);
and U2495 (N_2495,In_1003,In_1379);
and U2496 (N_2496,In_597,In_776);
nand U2497 (N_2497,In_414,In_1386);
and U2498 (N_2498,In_1021,In_468);
nor U2499 (N_2499,In_1446,In_782);
and U2500 (N_2500,In_1261,In_576);
xor U2501 (N_2501,In_1237,In_652);
nor U2502 (N_2502,In_634,In_445);
nor U2503 (N_2503,In_86,In_1381);
or U2504 (N_2504,In_461,In_1117);
or U2505 (N_2505,In_1356,In_385);
or U2506 (N_2506,In_1257,In_1123);
or U2507 (N_2507,In_210,In_979);
or U2508 (N_2508,In_1019,In_126);
or U2509 (N_2509,In_1136,In_1111);
nand U2510 (N_2510,In_933,In_1160);
nand U2511 (N_2511,In_531,In_342);
or U2512 (N_2512,In_584,In_70);
nand U2513 (N_2513,In_349,In_398);
nor U2514 (N_2514,In_348,In_563);
nand U2515 (N_2515,In_1044,In_467);
and U2516 (N_2516,In_1130,In_409);
and U2517 (N_2517,In_136,In_1423);
nand U2518 (N_2518,In_1163,In_1210);
nor U2519 (N_2519,In_435,In_137);
nor U2520 (N_2520,In_381,In_500);
and U2521 (N_2521,In_388,In_653);
nor U2522 (N_2522,In_527,In_1377);
and U2523 (N_2523,In_996,In_1141);
nand U2524 (N_2524,In_572,In_327);
or U2525 (N_2525,In_228,In_334);
or U2526 (N_2526,In_769,In_366);
nor U2527 (N_2527,In_17,In_877);
nor U2528 (N_2528,In_1338,In_1245);
nand U2529 (N_2529,In_426,In_79);
or U2530 (N_2530,In_1245,In_767);
and U2531 (N_2531,In_879,In_1358);
or U2532 (N_2532,In_336,In_279);
nor U2533 (N_2533,In_1459,In_1083);
nand U2534 (N_2534,In_1068,In_1218);
nand U2535 (N_2535,In_884,In_1475);
and U2536 (N_2536,In_313,In_854);
and U2537 (N_2537,In_1453,In_192);
and U2538 (N_2538,In_122,In_967);
nor U2539 (N_2539,In_1270,In_657);
or U2540 (N_2540,In_333,In_330);
nand U2541 (N_2541,In_1453,In_542);
or U2542 (N_2542,In_937,In_1361);
or U2543 (N_2543,In_1407,In_875);
nor U2544 (N_2544,In_652,In_778);
and U2545 (N_2545,In_841,In_311);
or U2546 (N_2546,In_1205,In_95);
nor U2547 (N_2547,In_992,In_1168);
nand U2548 (N_2548,In_1378,In_1073);
or U2549 (N_2549,In_837,In_1251);
and U2550 (N_2550,In_91,In_328);
or U2551 (N_2551,In_944,In_1007);
and U2552 (N_2552,In_605,In_230);
nand U2553 (N_2553,In_1246,In_1348);
nand U2554 (N_2554,In_1296,In_1187);
nor U2555 (N_2555,In_188,In_759);
nand U2556 (N_2556,In_1284,In_329);
nor U2557 (N_2557,In_897,In_1152);
nor U2558 (N_2558,In_578,In_900);
nand U2559 (N_2559,In_1317,In_968);
nand U2560 (N_2560,In_706,In_520);
nor U2561 (N_2561,In_1246,In_729);
and U2562 (N_2562,In_655,In_680);
xor U2563 (N_2563,In_962,In_1182);
or U2564 (N_2564,In_82,In_1091);
or U2565 (N_2565,In_8,In_1126);
or U2566 (N_2566,In_505,In_179);
or U2567 (N_2567,In_830,In_1487);
or U2568 (N_2568,In_530,In_746);
or U2569 (N_2569,In_1290,In_476);
or U2570 (N_2570,In_207,In_1022);
and U2571 (N_2571,In_679,In_209);
or U2572 (N_2572,In_6,In_950);
nand U2573 (N_2573,In_1392,In_1443);
and U2574 (N_2574,In_128,In_1270);
nor U2575 (N_2575,In_615,In_1375);
nor U2576 (N_2576,In_769,In_669);
and U2577 (N_2577,In_785,In_270);
and U2578 (N_2578,In_1170,In_834);
nand U2579 (N_2579,In_451,In_842);
nand U2580 (N_2580,In_515,In_1333);
or U2581 (N_2581,In_1302,In_35);
nand U2582 (N_2582,In_1412,In_344);
or U2583 (N_2583,In_106,In_51);
and U2584 (N_2584,In_1053,In_466);
and U2585 (N_2585,In_84,In_812);
and U2586 (N_2586,In_907,In_526);
and U2587 (N_2587,In_1144,In_821);
and U2588 (N_2588,In_425,In_498);
nand U2589 (N_2589,In_520,In_187);
or U2590 (N_2590,In_408,In_1434);
xnor U2591 (N_2591,In_1293,In_1226);
or U2592 (N_2592,In_41,In_317);
or U2593 (N_2593,In_967,In_90);
and U2594 (N_2594,In_152,In_420);
nor U2595 (N_2595,In_70,In_1026);
nand U2596 (N_2596,In_1360,In_328);
and U2597 (N_2597,In_493,In_999);
or U2598 (N_2598,In_178,In_1069);
nand U2599 (N_2599,In_473,In_993);
or U2600 (N_2600,In_840,In_666);
nand U2601 (N_2601,In_114,In_855);
nand U2602 (N_2602,In_1106,In_837);
or U2603 (N_2603,In_980,In_1384);
and U2604 (N_2604,In_561,In_1266);
or U2605 (N_2605,In_1431,In_422);
or U2606 (N_2606,In_15,In_1327);
and U2607 (N_2607,In_89,In_663);
and U2608 (N_2608,In_1390,In_336);
nor U2609 (N_2609,In_1032,In_271);
and U2610 (N_2610,In_531,In_221);
or U2611 (N_2611,In_1224,In_471);
nor U2612 (N_2612,In_877,In_867);
nand U2613 (N_2613,In_391,In_82);
nor U2614 (N_2614,In_691,In_406);
or U2615 (N_2615,In_428,In_1220);
or U2616 (N_2616,In_3,In_491);
or U2617 (N_2617,In_735,In_1407);
xor U2618 (N_2618,In_1252,In_1345);
and U2619 (N_2619,In_294,In_1320);
and U2620 (N_2620,In_692,In_1464);
nand U2621 (N_2621,In_1468,In_1309);
nand U2622 (N_2622,In_1243,In_1104);
nor U2623 (N_2623,In_1044,In_436);
nor U2624 (N_2624,In_831,In_417);
nand U2625 (N_2625,In_238,In_1319);
nor U2626 (N_2626,In_1310,In_1420);
xor U2627 (N_2627,In_851,In_980);
xor U2628 (N_2628,In_874,In_1413);
and U2629 (N_2629,In_6,In_1459);
nand U2630 (N_2630,In_396,In_774);
or U2631 (N_2631,In_655,In_1013);
nor U2632 (N_2632,In_202,In_791);
nand U2633 (N_2633,In_437,In_701);
nor U2634 (N_2634,In_1331,In_486);
and U2635 (N_2635,In_1290,In_427);
nor U2636 (N_2636,In_327,In_214);
and U2637 (N_2637,In_237,In_1221);
or U2638 (N_2638,In_210,In_926);
nor U2639 (N_2639,In_1375,In_1402);
or U2640 (N_2640,In_706,In_1342);
nand U2641 (N_2641,In_1496,In_608);
nand U2642 (N_2642,In_1167,In_632);
nor U2643 (N_2643,In_575,In_255);
or U2644 (N_2644,In_1184,In_599);
nand U2645 (N_2645,In_26,In_430);
and U2646 (N_2646,In_132,In_48);
and U2647 (N_2647,In_47,In_1043);
nor U2648 (N_2648,In_977,In_1004);
and U2649 (N_2649,In_69,In_1056);
and U2650 (N_2650,In_864,In_1139);
nor U2651 (N_2651,In_1379,In_906);
nand U2652 (N_2652,In_245,In_368);
nor U2653 (N_2653,In_1229,In_83);
nor U2654 (N_2654,In_168,In_59);
and U2655 (N_2655,In_867,In_931);
nand U2656 (N_2656,In_312,In_234);
nor U2657 (N_2657,In_863,In_287);
or U2658 (N_2658,In_1205,In_975);
nand U2659 (N_2659,In_698,In_605);
nand U2660 (N_2660,In_4,In_358);
and U2661 (N_2661,In_267,In_1462);
or U2662 (N_2662,In_359,In_377);
nor U2663 (N_2663,In_578,In_1025);
or U2664 (N_2664,In_322,In_343);
and U2665 (N_2665,In_455,In_890);
xor U2666 (N_2666,In_146,In_283);
or U2667 (N_2667,In_1019,In_35);
nor U2668 (N_2668,In_703,In_1257);
or U2669 (N_2669,In_424,In_323);
nand U2670 (N_2670,In_924,In_906);
or U2671 (N_2671,In_1,In_702);
and U2672 (N_2672,In_1375,In_394);
nand U2673 (N_2673,In_1423,In_1317);
nand U2674 (N_2674,In_423,In_837);
nor U2675 (N_2675,In_1377,In_222);
nand U2676 (N_2676,In_618,In_660);
or U2677 (N_2677,In_1091,In_1475);
and U2678 (N_2678,In_752,In_872);
nor U2679 (N_2679,In_950,In_546);
or U2680 (N_2680,In_71,In_453);
and U2681 (N_2681,In_744,In_706);
nand U2682 (N_2682,In_663,In_1441);
nand U2683 (N_2683,In_143,In_853);
nor U2684 (N_2684,In_52,In_1437);
nor U2685 (N_2685,In_1408,In_611);
or U2686 (N_2686,In_978,In_1499);
nand U2687 (N_2687,In_1233,In_1032);
or U2688 (N_2688,In_1022,In_224);
nand U2689 (N_2689,In_1306,In_1484);
or U2690 (N_2690,In_349,In_1369);
nor U2691 (N_2691,In_997,In_52);
nor U2692 (N_2692,In_68,In_530);
nor U2693 (N_2693,In_1283,In_620);
nand U2694 (N_2694,In_1292,In_30);
or U2695 (N_2695,In_1182,In_19);
or U2696 (N_2696,In_961,In_342);
and U2697 (N_2697,In_1046,In_50);
or U2698 (N_2698,In_1290,In_919);
nor U2699 (N_2699,In_1130,In_310);
nand U2700 (N_2700,In_1387,In_811);
and U2701 (N_2701,In_1253,In_433);
nor U2702 (N_2702,In_234,In_605);
nand U2703 (N_2703,In_1297,In_261);
nand U2704 (N_2704,In_570,In_835);
nor U2705 (N_2705,In_1339,In_307);
and U2706 (N_2706,In_1314,In_332);
nand U2707 (N_2707,In_880,In_1131);
or U2708 (N_2708,In_758,In_139);
nand U2709 (N_2709,In_476,In_1235);
nor U2710 (N_2710,In_203,In_118);
and U2711 (N_2711,In_131,In_541);
and U2712 (N_2712,In_1165,In_632);
or U2713 (N_2713,In_1065,In_1196);
nor U2714 (N_2714,In_584,In_1377);
nor U2715 (N_2715,In_1237,In_834);
or U2716 (N_2716,In_1050,In_1003);
nor U2717 (N_2717,In_742,In_110);
and U2718 (N_2718,In_1364,In_436);
nor U2719 (N_2719,In_1424,In_1246);
and U2720 (N_2720,In_1456,In_325);
nor U2721 (N_2721,In_451,In_700);
nor U2722 (N_2722,In_576,In_557);
and U2723 (N_2723,In_718,In_403);
nand U2724 (N_2724,In_647,In_703);
nand U2725 (N_2725,In_503,In_1221);
and U2726 (N_2726,In_514,In_1281);
nor U2727 (N_2727,In_284,In_199);
nand U2728 (N_2728,In_750,In_1023);
nand U2729 (N_2729,In_995,In_36);
or U2730 (N_2730,In_321,In_235);
or U2731 (N_2731,In_876,In_1275);
nor U2732 (N_2732,In_15,In_367);
nor U2733 (N_2733,In_821,In_83);
nor U2734 (N_2734,In_215,In_32);
and U2735 (N_2735,In_92,In_38);
or U2736 (N_2736,In_938,In_299);
nand U2737 (N_2737,In_801,In_1013);
or U2738 (N_2738,In_1003,In_1388);
nor U2739 (N_2739,In_527,In_648);
and U2740 (N_2740,In_164,In_1043);
or U2741 (N_2741,In_1154,In_1072);
or U2742 (N_2742,In_1481,In_557);
and U2743 (N_2743,In_1136,In_83);
or U2744 (N_2744,In_281,In_639);
or U2745 (N_2745,In_1177,In_912);
and U2746 (N_2746,In_566,In_1318);
nand U2747 (N_2747,In_1148,In_1378);
and U2748 (N_2748,In_1266,In_846);
xor U2749 (N_2749,In_800,In_1013);
and U2750 (N_2750,In_675,In_812);
nand U2751 (N_2751,In_138,In_1179);
and U2752 (N_2752,In_240,In_342);
nand U2753 (N_2753,In_550,In_617);
nand U2754 (N_2754,In_11,In_1216);
nand U2755 (N_2755,In_76,In_1196);
and U2756 (N_2756,In_1402,In_448);
xor U2757 (N_2757,In_472,In_665);
and U2758 (N_2758,In_388,In_602);
nand U2759 (N_2759,In_1289,In_1356);
or U2760 (N_2760,In_91,In_906);
nor U2761 (N_2761,In_1139,In_749);
xor U2762 (N_2762,In_193,In_85);
and U2763 (N_2763,In_160,In_280);
or U2764 (N_2764,In_1129,In_632);
nand U2765 (N_2765,In_404,In_282);
nand U2766 (N_2766,In_505,In_1491);
nor U2767 (N_2767,In_629,In_1395);
or U2768 (N_2768,In_1277,In_428);
nand U2769 (N_2769,In_844,In_1043);
and U2770 (N_2770,In_274,In_528);
nor U2771 (N_2771,In_1143,In_1426);
nor U2772 (N_2772,In_1472,In_1252);
and U2773 (N_2773,In_1232,In_51);
nor U2774 (N_2774,In_827,In_992);
xnor U2775 (N_2775,In_1298,In_1196);
or U2776 (N_2776,In_46,In_793);
nor U2777 (N_2777,In_794,In_933);
nand U2778 (N_2778,In_553,In_1479);
nor U2779 (N_2779,In_489,In_740);
and U2780 (N_2780,In_1341,In_1183);
nor U2781 (N_2781,In_591,In_220);
nand U2782 (N_2782,In_342,In_645);
nand U2783 (N_2783,In_960,In_695);
and U2784 (N_2784,In_454,In_1280);
or U2785 (N_2785,In_1200,In_1326);
nor U2786 (N_2786,In_552,In_154);
or U2787 (N_2787,In_1169,In_1189);
or U2788 (N_2788,In_441,In_1369);
nand U2789 (N_2789,In_161,In_894);
or U2790 (N_2790,In_694,In_706);
nor U2791 (N_2791,In_1109,In_1021);
nand U2792 (N_2792,In_1278,In_1061);
and U2793 (N_2793,In_204,In_284);
and U2794 (N_2794,In_1299,In_246);
nand U2795 (N_2795,In_304,In_620);
xnor U2796 (N_2796,In_1165,In_646);
nand U2797 (N_2797,In_628,In_338);
nor U2798 (N_2798,In_591,In_238);
nand U2799 (N_2799,In_1288,In_81);
and U2800 (N_2800,In_783,In_1071);
xnor U2801 (N_2801,In_50,In_799);
and U2802 (N_2802,In_607,In_1095);
nor U2803 (N_2803,In_873,In_448);
or U2804 (N_2804,In_1405,In_497);
and U2805 (N_2805,In_607,In_493);
nand U2806 (N_2806,In_69,In_1201);
nor U2807 (N_2807,In_286,In_939);
and U2808 (N_2808,In_565,In_880);
or U2809 (N_2809,In_831,In_1401);
or U2810 (N_2810,In_1099,In_1115);
and U2811 (N_2811,In_1179,In_575);
and U2812 (N_2812,In_1330,In_1130);
nor U2813 (N_2813,In_570,In_1402);
or U2814 (N_2814,In_1069,In_1271);
nand U2815 (N_2815,In_109,In_1070);
and U2816 (N_2816,In_841,In_1176);
xnor U2817 (N_2817,In_1259,In_1489);
or U2818 (N_2818,In_833,In_30);
and U2819 (N_2819,In_1114,In_248);
xor U2820 (N_2820,In_1042,In_500);
and U2821 (N_2821,In_921,In_134);
or U2822 (N_2822,In_1320,In_1402);
and U2823 (N_2823,In_1123,In_1177);
nand U2824 (N_2824,In_698,In_1201);
and U2825 (N_2825,In_439,In_19);
or U2826 (N_2826,In_211,In_266);
or U2827 (N_2827,In_817,In_1029);
nor U2828 (N_2828,In_883,In_1086);
and U2829 (N_2829,In_283,In_123);
or U2830 (N_2830,In_977,In_99);
and U2831 (N_2831,In_1250,In_1184);
and U2832 (N_2832,In_1154,In_657);
and U2833 (N_2833,In_644,In_666);
nand U2834 (N_2834,In_761,In_928);
or U2835 (N_2835,In_942,In_1416);
nand U2836 (N_2836,In_248,In_313);
or U2837 (N_2837,In_402,In_628);
and U2838 (N_2838,In_1077,In_401);
nand U2839 (N_2839,In_1083,In_489);
nand U2840 (N_2840,In_110,In_105);
or U2841 (N_2841,In_228,In_1412);
nor U2842 (N_2842,In_572,In_1352);
nand U2843 (N_2843,In_670,In_560);
nor U2844 (N_2844,In_866,In_1030);
and U2845 (N_2845,In_464,In_481);
nor U2846 (N_2846,In_1453,In_444);
nand U2847 (N_2847,In_1082,In_308);
and U2848 (N_2848,In_1101,In_186);
nor U2849 (N_2849,In_1125,In_107);
or U2850 (N_2850,In_1143,In_805);
and U2851 (N_2851,In_1360,In_1266);
or U2852 (N_2852,In_1104,In_1202);
or U2853 (N_2853,In_875,In_877);
or U2854 (N_2854,In_448,In_564);
or U2855 (N_2855,In_359,In_588);
or U2856 (N_2856,In_1050,In_1452);
or U2857 (N_2857,In_754,In_961);
or U2858 (N_2858,In_1003,In_903);
nor U2859 (N_2859,In_1149,In_327);
or U2860 (N_2860,In_1313,In_396);
and U2861 (N_2861,In_252,In_1233);
and U2862 (N_2862,In_1476,In_969);
and U2863 (N_2863,In_82,In_380);
or U2864 (N_2864,In_93,In_1076);
and U2865 (N_2865,In_939,In_828);
nand U2866 (N_2866,In_894,In_1413);
nand U2867 (N_2867,In_849,In_1005);
and U2868 (N_2868,In_384,In_1133);
nor U2869 (N_2869,In_1247,In_1033);
or U2870 (N_2870,In_917,In_1056);
nor U2871 (N_2871,In_360,In_1487);
or U2872 (N_2872,In_153,In_559);
nand U2873 (N_2873,In_39,In_472);
and U2874 (N_2874,In_1211,In_571);
nand U2875 (N_2875,In_377,In_240);
nor U2876 (N_2876,In_216,In_1087);
nor U2877 (N_2877,In_1258,In_943);
nor U2878 (N_2878,In_130,In_688);
xnor U2879 (N_2879,In_787,In_1348);
nor U2880 (N_2880,In_1019,In_1191);
nand U2881 (N_2881,In_719,In_146);
and U2882 (N_2882,In_1080,In_940);
nand U2883 (N_2883,In_232,In_237);
nor U2884 (N_2884,In_444,In_121);
nor U2885 (N_2885,In_390,In_4);
nor U2886 (N_2886,In_637,In_210);
nand U2887 (N_2887,In_712,In_772);
nor U2888 (N_2888,In_36,In_502);
and U2889 (N_2889,In_1455,In_114);
and U2890 (N_2890,In_1029,In_206);
and U2891 (N_2891,In_587,In_1071);
and U2892 (N_2892,In_518,In_1369);
nand U2893 (N_2893,In_1253,In_1228);
nor U2894 (N_2894,In_1420,In_1171);
or U2895 (N_2895,In_571,In_94);
or U2896 (N_2896,In_1444,In_673);
nand U2897 (N_2897,In_1034,In_558);
or U2898 (N_2898,In_732,In_1223);
and U2899 (N_2899,In_373,In_713);
and U2900 (N_2900,In_3,In_830);
xnor U2901 (N_2901,In_434,In_1492);
and U2902 (N_2902,In_527,In_96);
nor U2903 (N_2903,In_1352,In_130);
nand U2904 (N_2904,In_1438,In_353);
and U2905 (N_2905,In_334,In_1032);
nand U2906 (N_2906,In_369,In_367);
nand U2907 (N_2907,In_296,In_1101);
nand U2908 (N_2908,In_1302,In_1443);
nor U2909 (N_2909,In_175,In_415);
or U2910 (N_2910,In_789,In_1144);
nand U2911 (N_2911,In_432,In_745);
and U2912 (N_2912,In_358,In_279);
nor U2913 (N_2913,In_998,In_1140);
and U2914 (N_2914,In_125,In_616);
nand U2915 (N_2915,In_735,In_531);
nor U2916 (N_2916,In_616,In_1056);
nand U2917 (N_2917,In_342,In_398);
xnor U2918 (N_2918,In_1281,In_524);
or U2919 (N_2919,In_1213,In_609);
xnor U2920 (N_2920,In_361,In_1441);
nand U2921 (N_2921,In_1084,In_892);
nor U2922 (N_2922,In_153,In_1373);
and U2923 (N_2923,In_207,In_1065);
nor U2924 (N_2924,In_1123,In_969);
xnor U2925 (N_2925,In_817,In_1142);
nand U2926 (N_2926,In_786,In_887);
and U2927 (N_2927,In_122,In_958);
or U2928 (N_2928,In_1033,In_915);
or U2929 (N_2929,In_859,In_1464);
and U2930 (N_2930,In_212,In_19);
or U2931 (N_2931,In_264,In_81);
nand U2932 (N_2932,In_391,In_1253);
nor U2933 (N_2933,In_1087,In_919);
nand U2934 (N_2934,In_1487,In_974);
nor U2935 (N_2935,In_650,In_1194);
nor U2936 (N_2936,In_99,In_97);
nor U2937 (N_2937,In_1367,In_377);
nor U2938 (N_2938,In_1079,In_1405);
xor U2939 (N_2939,In_1214,In_322);
or U2940 (N_2940,In_1299,In_1306);
nand U2941 (N_2941,In_74,In_526);
or U2942 (N_2942,In_982,In_170);
nor U2943 (N_2943,In_359,In_146);
or U2944 (N_2944,In_937,In_1124);
and U2945 (N_2945,In_327,In_1315);
nand U2946 (N_2946,In_763,In_1376);
or U2947 (N_2947,In_326,In_667);
nand U2948 (N_2948,In_1296,In_1365);
or U2949 (N_2949,In_270,In_1444);
or U2950 (N_2950,In_936,In_241);
nor U2951 (N_2951,In_854,In_861);
and U2952 (N_2952,In_511,In_1187);
nand U2953 (N_2953,In_172,In_939);
nor U2954 (N_2954,In_187,In_637);
nand U2955 (N_2955,In_1262,In_92);
and U2956 (N_2956,In_1256,In_430);
nor U2957 (N_2957,In_271,In_226);
and U2958 (N_2958,In_988,In_72);
nand U2959 (N_2959,In_632,In_1330);
nand U2960 (N_2960,In_262,In_965);
nand U2961 (N_2961,In_1469,In_1255);
nor U2962 (N_2962,In_1480,In_649);
nor U2963 (N_2963,In_163,In_641);
nor U2964 (N_2964,In_4,In_1350);
nor U2965 (N_2965,In_183,In_1249);
nand U2966 (N_2966,In_971,In_454);
nor U2967 (N_2967,In_1357,In_596);
nor U2968 (N_2968,In_463,In_1381);
or U2969 (N_2969,In_42,In_433);
nor U2970 (N_2970,In_440,In_1408);
nand U2971 (N_2971,In_399,In_47);
and U2972 (N_2972,In_1114,In_1354);
nand U2973 (N_2973,In_512,In_1389);
or U2974 (N_2974,In_356,In_1256);
or U2975 (N_2975,In_191,In_1481);
nand U2976 (N_2976,In_259,In_152);
and U2977 (N_2977,In_1266,In_248);
or U2978 (N_2978,In_986,In_3);
or U2979 (N_2979,In_638,In_1481);
or U2980 (N_2980,In_899,In_65);
nand U2981 (N_2981,In_1319,In_1181);
nand U2982 (N_2982,In_1287,In_402);
nand U2983 (N_2983,In_980,In_1474);
nor U2984 (N_2984,In_1225,In_233);
or U2985 (N_2985,In_73,In_449);
nor U2986 (N_2986,In_1033,In_646);
and U2987 (N_2987,In_796,In_42);
and U2988 (N_2988,In_1182,In_1389);
and U2989 (N_2989,In_1229,In_1334);
or U2990 (N_2990,In_1371,In_219);
nor U2991 (N_2991,In_593,In_1239);
or U2992 (N_2992,In_1331,In_927);
nor U2993 (N_2993,In_255,In_911);
or U2994 (N_2994,In_752,In_643);
nor U2995 (N_2995,In_1390,In_307);
and U2996 (N_2996,In_875,In_1028);
nand U2997 (N_2997,In_911,In_318);
nand U2998 (N_2998,In_1008,In_666);
nor U2999 (N_2999,In_586,In_1054);
or U3000 (N_3000,N_1858,N_293);
nand U3001 (N_3001,N_2013,N_1318);
or U3002 (N_3002,N_2335,N_629);
nor U3003 (N_3003,N_525,N_550);
and U3004 (N_3004,N_335,N_1669);
nand U3005 (N_3005,N_2077,N_1113);
or U3006 (N_3006,N_985,N_2041);
and U3007 (N_3007,N_1056,N_2214);
nand U3008 (N_3008,N_250,N_2368);
or U3009 (N_3009,N_2930,N_92);
and U3010 (N_3010,N_2536,N_1547);
nor U3011 (N_3011,N_387,N_414);
nand U3012 (N_3012,N_1041,N_401);
nand U3013 (N_3013,N_999,N_695);
or U3014 (N_3014,N_1257,N_2140);
nand U3015 (N_3015,N_1554,N_2120);
xor U3016 (N_3016,N_505,N_2730);
and U3017 (N_3017,N_1484,N_1921);
or U3018 (N_3018,N_273,N_2142);
nand U3019 (N_3019,N_616,N_1292);
nor U3020 (N_3020,N_1181,N_2322);
or U3021 (N_3021,N_2807,N_1987);
or U3022 (N_3022,N_2566,N_2055);
nand U3023 (N_3023,N_927,N_1444);
or U3024 (N_3024,N_1273,N_1710);
nand U3025 (N_3025,N_2644,N_2445);
nor U3026 (N_3026,N_2786,N_82);
nand U3027 (N_3027,N_1164,N_1007);
nand U3028 (N_3028,N_1751,N_2698);
nor U3029 (N_3029,N_2617,N_1127);
and U3030 (N_3030,N_957,N_1174);
nand U3031 (N_3031,N_309,N_1438);
nor U3032 (N_3032,N_2707,N_1765);
or U3033 (N_3033,N_344,N_2375);
or U3034 (N_3034,N_655,N_462);
nor U3035 (N_3035,N_1173,N_2020);
nor U3036 (N_3036,N_410,N_1551);
or U3037 (N_3037,N_2045,N_2560);
nand U3038 (N_3038,N_877,N_2752);
nand U3039 (N_3039,N_1842,N_1357);
or U3040 (N_3040,N_408,N_586);
nor U3041 (N_3041,N_1664,N_1381);
or U3042 (N_3042,N_640,N_2802);
and U3043 (N_3043,N_1199,N_1902);
or U3044 (N_3044,N_910,N_39);
nand U3045 (N_3045,N_1410,N_1186);
or U3046 (N_3046,N_2546,N_772);
nand U3047 (N_3047,N_576,N_1363);
and U3048 (N_3048,N_2917,N_2936);
nor U3049 (N_3049,N_1226,N_2921);
nor U3050 (N_3050,N_1562,N_1275);
or U3051 (N_3051,N_2902,N_1268);
or U3052 (N_3052,N_1740,N_2685);
nand U3053 (N_3053,N_2024,N_1465);
or U3054 (N_3054,N_946,N_1653);
nand U3055 (N_3055,N_1963,N_1420);
nor U3056 (N_3056,N_1689,N_2767);
and U3057 (N_3057,N_2282,N_2231);
nor U3058 (N_3058,N_1535,N_2486);
or U3059 (N_3059,N_533,N_933);
nor U3060 (N_3060,N_2117,N_1764);
nand U3061 (N_3061,N_1491,N_2172);
or U3062 (N_3062,N_2237,N_2671);
nor U3063 (N_3063,N_1757,N_995);
nor U3064 (N_3064,N_2725,N_376);
and U3065 (N_3065,N_1140,N_650);
and U3066 (N_3066,N_952,N_2704);
nand U3067 (N_3067,N_1838,N_1236);
nor U3068 (N_3068,N_1726,N_2190);
nor U3069 (N_3069,N_24,N_809);
nand U3070 (N_3070,N_276,N_1477);
and U3071 (N_3071,N_1213,N_291);
nand U3072 (N_3072,N_1623,N_1474);
nand U3073 (N_3073,N_1237,N_2145);
xor U3074 (N_3074,N_553,N_1175);
or U3075 (N_3075,N_2434,N_1069);
nand U3076 (N_3076,N_2580,N_1251);
or U3077 (N_3077,N_1681,N_2418);
and U3078 (N_3078,N_499,N_2880);
and U3079 (N_3079,N_581,N_1328);
or U3080 (N_3080,N_2683,N_1883);
and U3081 (N_3081,N_734,N_498);
and U3082 (N_3082,N_2895,N_2626);
nand U3083 (N_3083,N_1797,N_2052);
and U3084 (N_3084,N_2836,N_395);
nand U3085 (N_3085,N_1561,N_482);
and U3086 (N_3086,N_1261,N_2789);
or U3087 (N_3087,N_1933,N_256);
or U3088 (N_3088,N_1806,N_440);
nor U3089 (N_3089,N_1559,N_583);
nand U3090 (N_3090,N_1832,N_966);
nand U3091 (N_3091,N_2378,N_804);
nand U3092 (N_3092,N_449,N_2212);
nand U3093 (N_3093,N_2544,N_2497);
nor U3094 (N_3094,N_2977,N_980);
nand U3095 (N_3095,N_543,N_753);
nand U3096 (N_3096,N_2809,N_2998);
or U3097 (N_3097,N_1530,N_2135);
nor U3098 (N_3098,N_494,N_762);
and U3099 (N_3099,N_106,N_1055);
and U3100 (N_3100,N_1819,N_2596);
and U3101 (N_3101,N_422,N_302);
or U3102 (N_3102,N_2892,N_1560);
and U3103 (N_3103,N_2539,N_119);
and U3104 (N_3104,N_2840,N_987);
or U3105 (N_3105,N_1802,N_467);
nor U3106 (N_3106,N_638,N_204);
and U3107 (N_3107,N_920,N_2694);
or U3108 (N_3108,N_1163,N_763);
nor U3109 (N_3109,N_77,N_521);
and U3110 (N_3110,N_2496,N_1752);
and U3111 (N_3111,N_2124,N_856);
nand U3112 (N_3112,N_711,N_796);
or U3113 (N_3113,N_2687,N_2852);
nand U3114 (N_3114,N_2064,N_1239);
nor U3115 (N_3115,N_720,N_2974);
xnor U3116 (N_3116,N_2995,N_2473);
and U3117 (N_3117,N_1976,N_1855);
nand U3118 (N_3118,N_2218,N_1013);
nand U3119 (N_3119,N_802,N_1015);
or U3120 (N_3120,N_2967,N_163);
nand U3121 (N_3121,N_1729,N_2054);
nand U3122 (N_3122,N_2086,N_1049);
nand U3123 (N_3123,N_430,N_148);
and U3124 (N_3124,N_318,N_2563);
nor U3125 (N_3125,N_2913,N_2464);
nand U3126 (N_3126,N_798,N_2484);
nor U3127 (N_3127,N_384,N_1613);
nand U3128 (N_3128,N_1542,N_822);
or U3129 (N_3129,N_2303,N_1234);
nor U3130 (N_3130,N_2147,N_1338);
nand U3131 (N_3131,N_2529,N_1320);
and U3132 (N_3132,N_2527,N_2164);
nand U3133 (N_3133,N_974,N_2317);
nand U3134 (N_3134,N_951,N_277);
or U3135 (N_3135,N_2148,N_502);
nor U3136 (N_3136,N_1051,N_2273);
nor U3137 (N_3137,N_2586,N_1690);
nor U3138 (N_3138,N_765,N_1329);
nand U3139 (N_3139,N_630,N_2647);
or U3140 (N_3140,N_253,N_2106);
nor U3141 (N_3141,N_2310,N_2171);
and U3142 (N_3142,N_377,N_2449);
or U3143 (N_3143,N_1265,N_851);
or U3144 (N_3144,N_2990,N_1748);
or U3145 (N_3145,N_539,N_2396);
nand U3146 (N_3146,N_2177,N_1167);
nor U3147 (N_3147,N_1548,N_2069);
or U3148 (N_3148,N_345,N_2079);
or U3149 (N_3149,N_2391,N_2167);
nand U3150 (N_3150,N_1004,N_1367);
or U3151 (N_3151,N_2957,N_1467);
nand U3152 (N_3152,N_2621,N_2210);
nand U3153 (N_3153,N_90,N_797);
nor U3154 (N_3154,N_1433,N_216);
and U3155 (N_3155,N_1650,N_1938);
nor U3156 (N_3156,N_1878,N_1545);
and U3157 (N_3157,N_1035,N_903);
nand U3158 (N_3158,N_490,N_2379);
or U3159 (N_3159,N_777,N_371);
nand U3160 (N_3160,N_64,N_2111);
and U3161 (N_3161,N_1135,N_2451);
and U3162 (N_3162,N_1067,N_2143);
nor U3163 (N_3163,N_1179,N_676);
nor U3164 (N_3164,N_2792,N_2878);
xnor U3165 (N_3165,N_2255,N_1877);
nor U3166 (N_3166,N_2184,N_2315);
nand U3167 (N_3167,N_448,N_488);
or U3168 (N_3168,N_1362,N_34);
or U3169 (N_3169,N_2945,N_160);
nor U3170 (N_3170,N_2492,N_1820);
xor U3171 (N_3171,N_875,N_1032);
and U3172 (N_3172,N_2993,N_2651);
nand U3173 (N_3173,N_2485,N_2779);
nand U3174 (N_3174,N_1934,N_2562);
or U3175 (N_3175,N_2505,N_2059);
and U3176 (N_3176,N_1121,N_2600);
nand U3177 (N_3177,N_1852,N_218);
nor U3178 (N_3178,N_165,N_257);
and U3179 (N_3179,N_1045,N_694);
nand U3180 (N_3180,N_486,N_1612);
and U3181 (N_3181,N_2615,N_1808);
or U3182 (N_3182,N_2031,N_565);
and U3183 (N_3183,N_2851,N_2224);
or U3184 (N_3184,N_1380,N_1849);
or U3185 (N_3185,N_1603,N_1799);
nor U3186 (N_3186,N_69,N_2568);
or U3187 (N_3187,N_2264,N_1546);
nand U3188 (N_3188,N_1183,N_1622);
nor U3189 (N_3189,N_1458,N_1416);
nand U3190 (N_3190,N_2460,N_2886);
nor U3191 (N_3191,N_1598,N_2541);
nor U3192 (N_3192,N_2735,N_751);
nor U3193 (N_3193,N_579,N_2196);
nor U3194 (N_3194,N_1198,N_2215);
xnor U3195 (N_3195,N_2857,N_2405);
or U3196 (N_3196,N_2848,N_1582);
or U3197 (N_3197,N_1854,N_1024);
and U3198 (N_3198,N_2274,N_2818);
or U3199 (N_3199,N_1128,N_531);
and U3200 (N_3200,N_2718,N_2);
or U3201 (N_3201,N_632,N_342);
xor U3202 (N_3202,N_209,N_1117);
nor U3203 (N_3203,N_739,N_234);
or U3204 (N_3204,N_813,N_535);
nand U3205 (N_3205,N_2666,N_2979);
nand U3206 (N_3206,N_301,N_678);
nor U3207 (N_3207,N_2431,N_2994);
and U3208 (N_3208,N_364,N_465);
nor U3209 (N_3209,N_2858,N_284);
nand U3210 (N_3210,N_1993,N_577);
nor U3211 (N_3211,N_1897,N_807);
nor U3212 (N_3212,N_2668,N_1372);
nand U3213 (N_3213,N_1743,N_729);
nor U3214 (N_3214,N_1632,N_242);
and U3215 (N_3215,N_902,N_834);
nor U3216 (N_3216,N_2008,N_2442);
and U3217 (N_3217,N_2741,N_2720);
and U3218 (N_3218,N_955,N_808);
nor U3219 (N_3219,N_2844,N_1654);
nand U3220 (N_3220,N_456,N_123);
or U3221 (N_3221,N_76,N_2098);
nor U3222 (N_3222,N_2477,N_1633);
nand U3223 (N_3223,N_874,N_223);
or U3224 (N_3224,N_2897,N_2910);
nor U3225 (N_3225,N_2395,N_476);
and U3226 (N_3226,N_2161,N_2777);
nand U3227 (N_3227,N_1450,N_2991);
nor U3228 (N_3228,N_469,N_429);
and U3229 (N_3229,N_2480,N_2740);
and U3230 (N_3230,N_1626,N_596);
nor U3231 (N_3231,N_2987,N_1777);
and U3232 (N_3232,N_756,N_748);
nor U3233 (N_3233,N_2204,N_1886);
nand U3234 (N_3234,N_1973,N_95);
nor U3235 (N_3235,N_2307,N_1655);
nand U3236 (N_3236,N_1716,N_2016);
nor U3237 (N_3237,N_1759,N_1053);
or U3238 (N_3238,N_2642,N_2276);
and U3239 (N_3239,N_1801,N_1435);
and U3240 (N_3240,N_2467,N_71);
and U3241 (N_3241,N_1665,N_1766);
nand U3242 (N_3242,N_1659,N_259);
nand U3243 (N_3243,N_645,N_2891);
nor U3244 (N_3244,N_50,N_178);
and U3245 (N_3245,N_761,N_2810);
and U3246 (N_3246,N_668,N_198);
or U3247 (N_3247,N_471,N_764);
or U3248 (N_3248,N_194,N_725);
or U3249 (N_3249,N_2270,N_2854);
and U3250 (N_3250,N_479,N_1657);
nand U3251 (N_3251,N_2439,N_2823);
nor U3252 (N_3252,N_982,N_2554);
nor U3253 (N_3253,N_517,N_2244);
and U3254 (N_3254,N_2619,N_1577);
and U3255 (N_3255,N_1014,N_824);
nor U3256 (N_3256,N_262,N_799);
nor U3257 (N_3257,N_1621,N_846);
nand U3258 (N_3258,N_197,N_1103);
nand U3259 (N_3259,N_1374,N_1411);
and U3260 (N_3260,N_1925,N_681);
nor U3261 (N_3261,N_1619,N_2017);
nor U3262 (N_3262,N_2532,N_1953);
or U3263 (N_3263,N_2042,N_1489);
nand U3264 (N_3264,N_1722,N_2597);
or U3265 (N_3265,N_871,N_339);
or U3266 (N_3266,N_1494,N_1466);
nand U3267 (N_3267,N_2409,N_27);
and U3268 (N_3268,N_14,N_2387);
nor U3269 (N_3269,N_1475,N_286);
nand U3270 (N_3270,N_1090,N_2162);
or U3271 (N_3271,N_2417,N_2081);
and U3272 (N_3272,N_491,N_464);
or U3273 (N_3273,N_131,N_2334);
or U3274 (N_3274,N_2499,N_2129);
or U3275 (N_3275,N_2150,N_2869);
nor U3276 (N_3276,N_1735,N_1635);
nor U3277 (N_3277,N_1401,N_2940);
nor U3278 (N_3278,N_2345,N_1637);
or U3279 (N_3279,N_1991,N_2201);
and U3280 (N_3280,N_2461,N_812);
and U3281 (N_3281,N_1412,N_526);
nand U3282 (N_3282,N_1666,N_1238);
nand U3283 (N_3283,N_2385,N_1075);
or U3284 (N_3284,N_2281,N_2688);
nand U3285 (N_3285,N_512,N_1640);
nor U3286 (N_3286,N_727,N_1076);
xnor U3287 (N_3287,N_1217,N_65);
nor U3288 (N_3288,N_338,N_388);
and U3289 (N_3289,N_2843,N_778);
or U3290 (N_3290,N_2817,N_861);
xor U3291 (N_3291,N_914,N_436);
nand U3292 (N_3292,N_2080,N_573);
nor U3293 (N_3293,N_993,N_1916);
nor U3294 (N_3294,N_1483,N_1732);
and U3295 (N_3295,N_833,N_169);
nand U3296 (N_3296,N_2478,N_609);
nand U3297 (N_3297,N_1158,N_1442);
or U3298 (N_3298,N_1382,N_461);
or U3299 (N_3299,N_509,N_1296);
nand U3300 (N_3300,N_152,N_4);
nand U3301 (N_3301,N_439,N_2296);
nor U3302 (N_3302,N_2929,N_1606);
and U3303 (N_3303,N_1792,N_811);
nor U3304 (N_3304,N_2846,N_2234);
nor U3305 (N_3305,N_1638,N_1889);
nand U3306 (N_3306,N_1966,N_2382);
nor U3307 (N_3307,N_1011,N_225);
and U3308 (N_3308,N_879,N_287);
or U3309 (N_3309,N_357,N_2716);
nor U3310 (N_3310,N_2424,N_784);
nor U3311 (N_3311,N_696,N_1452);
nor U3312 (N_3312,N_417,N_2436);
nor U3313 (N_3313,N_2037,N_2877);
nand U3314 (N_3314,N_19,N_2804);
nor U3315 (N_3315,N_1769,N_1969);
nor U3316 (N_3316,N_1837,N_984);
and U3317 (N_3317,N_1846,N_1397);
or U3318 (N_3318,N_1333,N_2975);
nor U3319 (N_3319,N_1364,N_1611);
or U3320 (N_3320,N_1870,N_2305);
and U3321 (N_3321,N_891,N_2701);
xnor U3322 (N_3322,N_68,N_1624);
nor U3323 (N_3323,N_1376,N_2549);
or U3324 (N_3324,N_1768,N_1402);
and U3325 (N_3325,N_2404,N_2631);
or U3326 (N_3326,N_2186,N_682);
or U3327 (N_3327,N_1259,N_754);
nor U3328 (N_3328,N_1375,N_2118);
nor U3329 (N_3329,N_158,N_383);
or U3330 (N_3330,N_906,N_2113);
or U3331 (N_3331,N_94,N_487);
nor U3332 (N_3332,N_1157,N_2907);
nand U3333 (N_3333,N_1303,N_945);
nor U3334 (N_3334,N_1242,N_703);
and U3335 (N_3335,N_1573,N_298);
nor U3336 (N_3336,N_1074,N_102);
and U3337 (N_3337,N_2348,N_379);
or U3338 (N_3338,N_1980,N_2251);
and U3339 (N_3339,N_1636,N_1246);
and U3340 (N_3340,N_2376,N_567);
or U3341 (N_3341,N_1297,N_2446);
nor U3342 (N_3342,N_559,N_2125);
nand U3343 (N_3343,N_1124,N_380);
nor U3344 (N_3344,N_201,N_1027);
nand U3345 (N_3345,N_353,N_1605);
nor U3346 (N_3346,N_771,N_2828);
nand U3347 (N_3347,N_973,N_2452);
nor U3348 (N_3348,N_2301,N_1094);
nor U3349 (N_3349,N_1737,N_1901);
and U3350 (N_3350,N_1197,N_1988);
or U3351 (N_3351,N_1352,N_1531);
nand U3352 (N_3352,N_474,N_972);
nor U3353 (N_3353,N_1332,N_2483);
and U3354 (N_3354,N_2246,N_386);
nor U3355 (N_3355,N_2588,N_516);
and U3356 (N_3356,N_99,N_2547);
nor U3357 (N_3357,N_1724,N_2057);
xnor U3358 (N_3358,N_1025,N_2341);
nor U3359 (N_3359,N_2415,N_1460);
nand U3360 (N_3360,N_1077,N_2414);
and U3361 (N_3361,N_2225,N_31);
and U3362 (N_3362,N_975,N_1644);
and U3363 (N_3363,N_2742,N_2394);
and U3364 (N_3364,N_1267,N_2399);
or U3365 (N_3365,N_300,N_1063);
nor U3366 (N_3366,N_736,N_1778);
and U3367 (N_3367,N_661,N_504);
nand U3368 (N_3368,N_1698,N_2606);
nor U3369 (N_3369,N_2028,N_255);
or U3370 (N_3370,N_1335,N_263);
and U3371 (N_3371,N_1543,N_2298);
or U3372 (N_3372,N_1084,N_781);
or U3373 (N_3373,N_2984,N_237);
nor U3374 (N_3374,N_2796,N_2326);
nand U3375 (N_3375,N_1155,N_2715);
nand U3376 (N_3376,N_1862,N_919);
or U3377 (N_3377,N_229,N_2455);
and U3378 (N_3378,N_1346,N_2358);
nor U3379 (N_3379,N_1522,N_212);
or U3380 (N_3380,N_1307,N_1628);
and U3381 (N_3381,N_75,N_1447);
and U3382 (N_3382,N_2471,N_2472);
xnor U3383 (N_3383,N_1393,N_519);
nand U3384 (N_3384,N_2782,N_1874);
and U3385 (N_3385,N_1208,N_1699);
and U3386 (N_3386,N_2753,N_2738);
nor U3387 (N_3387,N_2812,N_1201);
nand U3388 (N_3388,N_375,N_1369);
or U3389 (N_3389,N_496,N_2952);
or U3390 (N_3390,N_2832,N_1001);
nor U3391 (N_3391,N_1756,N_817);
and U3392 (N_3392,N_2015,N_1436);
xor U3393 (N_3393,N_2912,N_1642);
nand U3394 (N_3394,N_1947,N_1895);
or U3395 (N_3395,N_2618,N_1274);
or U3396 (N_3396,N_1313,N_2170);
nand U3397 (N_3397,N_1232,N_2552);
nor U3398 (N_3398,N_2132,N_113);
and U3399 (N_3399,N_2528,N_43);
nand U3400 (N_3400,N_1919,N_1558);
nor U3401 (N_3401,N_825,N_2468);
nor U3402 (N_3402,N_2627,N_2493);
and U3403 (N_3403,N_1370,N_2515);
and U3404 (N_3404,N_742,N_1604);
nor U3405 (N_3405,N_717,N_1220);
nand U3406 (N_3406,N_1107,N_1342);
nand U3407 (N_3407,N_1351,N_271);
and U3408 (N_3408,N_1961,N_9);
and U3409 (N_3409,N_2924,N_647);
and U3410 (N_3410,N_2029,N_2357);
nand U3411 (N_3411,N_1763,N_447);
nand U3412 (N_3412,N_2141,N_2075);
nand U3413 (N_3413,N_1462,N_20);
or U3414 (N_3414,N_1137,N_2879);
nor U3415 (N_3415,N_1583,N_2463);
nor U3416 (N_3416,N_74,N_708);
or U3417 (N_3417,N_1569,N_832);
nand U3418 (N_3418,N_1060,N_1083);
or U3419 (N_3419,N_2337,N_254);
and U3420 (N_3420,N_2909,N_2352);
and U3421 (N_3421,N_981,N_1576);
and U3422 (N_3422,N_2798,N_1749);
nor U3423 (N_3423,N_407,N_1932);
nor U3424 (N_3424,N_592,N_1828);
nand U3425 (N_3425,N_200,N_1266);
nor U3426 (N_3426,N_455,N_1147);
or U3427 (N_3427,N_1200,N_783);
and U3428 (N_3428,N_107,N_325);
nand U3429 (N_3429,N_2302,N_2732);
nor U3430 (N_3430,N_768,N_2390);
nand U3431 (N_3431,N_2706,N_2850);
or U3432 (N_3432,N_1414,N_2628);
nand U3433 (N_3433,N_2689,N_2128);
nor U3434 (N_3434,N_1997,N_1168);
nand U3435 (N_3435,N_1229,N_1805);
nor U3436 (N_3436,N_1386,N_2585);
and U3437 (N_3437,N_176,N_847);
or U3438 (N_3438,N_2006,N_654);
nor U3439 (N_3439,N_954,N_2437);
nor U3440 (N_3440,N_177,N_1652);
or U3441 (N_3441,N_2938,N_2476);
and U3442 (N_3442,N_1610,N_775);
nand U3443 (N_3443,N_1817,N_454);
or U3444 (N_3444,N_359,N_855);
nor U3445 (N_3445,N_1728,N_740);
xnor U3446 (N_3446,N_484,N_129);
or U3447 (N_3447,N_1887,N_1368);
nand U3448 (N_3448,N_1575,N_208);
nor U3449 (N_3449,N_1913,N_998);
or U3450 (N_3450,N_988,N_556);
nand U3451 (N_3451,N_572,N_2510);
nand U3452 (N_3452,N_1290,N_406);
and U3453 (N_3453,N_1345,N_558);
or U3454 (N_3454,N_2905,N_2675);
nor U3455 (N_3455,N_721,N_1325);
nor U3456 (N_3456,N_862,N_2350);
and U3457 (N_3457,N_529,N_1946);
or U3458 (N_3458,N_697,N_295);
nor U3459 (N_3459,N_2520,N_2127);
nor U3460 (N_3460,N_1812,N_880);
xor U3461 (N_3461,N_1927,N_1711);
and U3462 (N_3462,N_2043,N_1072);
and U3463 (N_3463,N_425,N_1905);
nor U3464 (N_3464,N_930,N_1441);
xor U3465 (N_3465,N_265,N_44);
and U3466 (N_3466,N_1818,N_601);
nor U3467 (N_3467,N_953,N_402);
or U3468 (N_3468,N_1384,N_2887);
nand U3469 (N_3469,N_435,N_141);
nand U3470 (N_3470,N_1283,N_1373);
and U3471 (N_3471,N_1291,N_2205);
nand U3472 (N_3472,N_1086,N_1519);
nor U3473 (N_3473,N_1936,N_1831);
nand U3474 (N_3474,N_2316,N_2349);
or U3475 (N_3475,N_1774,N_1971);
nor U3476 (N_3476,N_1225,N_2433);
or U3477 (N_3477,N_2949,N_2920);
nor U3478 (N_3478,N_2790,N_2686);
nand U3479 (N_3479,N_2776,N_1151);
nand U3480 (N_3480,N_182,N_1761);
or U3481 (N_3481,N_937,N_2060);
nor U3482 (N_3482,N_52,N_1834);
nor U3483 (N_3483,N_1798,N_312);
nor U3484 (N_3484,N_787,N_566);
and U3485 (N_3485,N_792,N_2014);
nor U3486 (N_3486,N_2904,N_58);
nand U3487 (N_3487,N_1178,N_2049);
nor U3488 (N_3488,N_2440,N_665);
nor U3489 (N_3489,N_1288,N_372);
and U3490 (N_3490,N_602,N_1493);
nor U3491 (N_3491,N_2822,N_278);
or U3492 (N_3492,N_2491,N_2531);
nor U3493 (N_3493,N_1034,N_2503);
nor U3494 (N_3494,N_2507,N_622);
and U3495 (N_3495,N_2663,N_506);
nand U3496 (N_3496,N_1111,N_2643);
nand U3497 (N_3497,N_2392,N_1082);
or U3498 (N_3498,N_901,N_1129);
and U3499 (N_3499,N_260,N_213);
and U3500 (N_3500,N_2968,N_2681);
nand U3501 (N_3501,N_2226,N_1935);
or U3502 (N_3502,N_2837,N_2839);
and U3503 (N_3503,N_2784,N_2088);
nor U3504 (N_3504,N_1159,N_2038);
nor U3505 (N_3505,N_350,N_1144);
and U3506 (N_3506,N_472,N_1294);
and U3507 (N_3507,N_849,N_2992);
xnor U3508 (N_3508,N_1550,N_2650);
and U3509 (N_3509,N_36,N_2956);
or U3510 (N_3510,N_2153,N_673);
and U3511 (N_3511,N_1299,N_2228);
nand U3512 (N_3512,N_571,N_1341);
nand U3513 (N_3513,N_282,N_627);
nand U3514 (N_3514,N_1028,N_1281);
and U3515 (N_3515,N_230,N_2030);
or U3516 (N_3516,N_1675,N_2602);
or U3517 (N_3517,N_2785,N_1696);
nor U3518 (N_3518,N_1425,N_2122);
nor U3519 (N_3519,N_2459,N_2447);
nand U3520 (N_3520,N_2370,N_548);
nand U3521 (N_3521,N_2572,N_2457);
nand U3522 (N_3522,N_2428,N_1787);
or U3523 (N_3523,N_41,N_1920);
and U3524 (N_3524,N_1567,N_962);
and U3525 (N_3525,N_2939,N_1998);
nand U3526 (N_3526,N_2295,N_1745);
or U3527 (N_3527,N_1326,N_1205);
and U3528 (N_3528,N_1950,N_156);
nor U3529 (N_3529,N_299,N_267);
and U3530 (N_3530,N_468,N_2188);
nand U3531 (N_3531,N_2801,N_545);
nand U3532 (N_3532,N_233,N_1544);
nor U3533 (N_3533,N_2773,N_21);
nand U3534 (N_3534,N_716,N_2284);
nor U3535 (N_3535,N_1772,N_316);
and U3536 (N_3536,N_1776,N_170);
and U3537 (N_3537,N_2416,N_532);
nor U3538 (N_3538,N_2521,N_2328);
nand U3539 (N_3539,N_1956,N_2209);
or U3540 (N_3540,N_2517,N_800);
and U3541 (N_3541,N_1836,N_1058);
or U3542 (N_3542,N_1131,N_1276);
or U3543 (N_3543,N_1959,N_2285);
and U3544 (N_3544,N_823,N_1453);
nand U3545 (N_3545,N_83,N_1588);
and U3546 (N_3546,N_1746,N_378);
and U3547 (N_3547,N_1700,N_1826);
nor U3548 (N_3548,N_2748,N_2855);
or U3549 (N_3549,N_2591,N_28);
nand U3550 (N_3550,N_195,N_2356);
nand U3551 (N_3551,N_2479,N_1262);
and U3552 (N_3552,N_2641,N_292);
nand U3553 (N_3553,N_1955,N_791);
nand U3554 (N_3554,N_672,N_620);
nand U3555 (N_3555,N_244,N_2071);
or U3556 (N_3556,N_2422,N_719);
nand U3557 (N_3557,N_2981,N_442);
nor U3558 (N_3558,N_1909,N_597);
nor U3559 (N_3559,N_1521,N_173);
nand U3560 (N_3560,N_733,N_2737);
nor U3561 (N_3561,N_2781,N_1830);
or U3562 (N_3562,N_2100,N_838);
nand U3563 (N_3563,N_32,N_639);
nor U3564 (N_3564,N_473,N_614);
nor U3565 (N_3565,N_1784,N_2928);
nor U3566 (N_3566,N_2814,N_598);
nand U3567 (N_3567,N_1951,N_2793);
nor U3568 (N_3568,N_633,N_928);
nand U3569 (N_3569,N_2339,N_1230);
nor U3570 (N_3570,N_1507,N_2340);
or U3571 (N_3571,N_2096,N_1911);
and U3572 (N_3572,N_2900,N_104);
nand U3573 (N_3573,N_831,N_2859);
nand U3574 (N_3574,N_290,N_25);
nand U3575 (N_3575,N_652,N_2999);
nor U3576 (N_3576,N_2761,N_801);
nand U3577 (N_3577,N_1037,N_40);
or U3578 (N_3578,N_2714,N_365);
nand U3579 (N_3579,N_306,N_1468);
nand U3580 (N_3580,N_723,N_243);
xnor U3581 (N_3581,N_1813,N_1446);
nand U3582 (N_3582,N_382,N_2342);
nor U3583 (N_3583,N_687,N_636);
nor U3584 (N_3584,N_746,N_1093);
xor U3585 (N_3585,N_500,N_162);
nand U3586 (N_3586,N_1580,N_2512);
nand U3587 (N_3587,N_908,N_1356);
nor U3588 (N_3588,N_2267,N_2412);
nor U3589 (N_3589,N_432,N_1712);
and U3590 (N_3590,N_2667,N_251);
or U3591 (N_3591,N_362,N_575);
or U3592 (N_3592,N_730,N_2400);
xor U3593 (N_3593,N_1713,N_2526);
nand U3594 (N_3594,N_1378,N_2001);
nand U3595 (N_3595,N_1876,N_749);
or U3596 (N_3596,N_308,N_1884);
nand U3597 (N_3597,N_397,N_495);
nor U3598 (N_3598,N_1009,N_1840);
or U3599 (N_3599,N_1894,N_986);
or U3600 (N_3600,N_1678,N_893);
nor U3601 (N_3601,N_646,N_1859);
or U3602 (N_3602,N_2138,N_108);
or U3603 (N_3603,N_2766,N_1646);
and U3604 (N_3604,N_2709,N_112);
nor U3605 (N_3605,N_224,N_1195);
or U3606 (N_3606,N_1810,N_726);
and U3607 (N_3607,N_1277,N_853);
nor U3608 (N_3608,N_2941,N_2094);
nor U3609 (N_3609,N_1042,N_2548);
nand U3610 (N_3610,N_2578,N_1172);
nor U3611 (N_3611,N_2947,N_1114);
nand U3612 (N_3612,N_839,N_2297);
nand U3613 (N_3613,N_662,N_100);
nand U3614 (N_3614,N_207,N_2506);
nor U3615 (N_3615,N_667,N_1355);
nor U3616 (N_3616,N_1064,N_1353);
or U3617 (N_3617,N_1404,N_2131);
or U3618 (N_3618,N_2565,N_111);
nor U3619 (N_3619,N_2915,N_2009);
nor U3620 (N_3620,N_147,N_2241);
nor U3621 (N_3621,N_404,N_2420);
and U3622 (N_3622,N_315,N_2332);
or U3623 (N_3623,N_423,N_1882);
xor U3624 (N_3624,N_319,N_1112);
nor U3625 (N_3625,N_1252,N_1469);
and U3626 (N_3626,N_16,N_2469);
nand U3627 (N_3627,N_1890,N_1518);
nor U3628 (N_3628,N_1990,N_485);
nand U3629 (N_3629,N_2398,N_2545);
nor U3630 (N_3630,N_1499,N_564);
nor U3631 (N_3631,N_1501,N_1319);
nand U3632 (N_3632,N_1502,N_2533);
nor U3633 (N_3633,N_2432,N_2372);
xnor U3634 (N_3634,N_1327,N_1249);
or U3635 (N_3635,N_2306,N_1078);
nand U3636 (N_3636,N_2193,N_1944);
nand U3637 (N_3637,N_735,N_950);
or U3638 (N_3638,N_606,N_247);
nand U3639 (N_3639,N_1286,N_1349);
or U3640 (N_3640,N_2608,N_884);
or U3641 (N_3641,N_1440,N_618);
nor U3642 (N_3642,N_361,N_1218);
or U3643 (N_3643,N_453,N_1682);
nor U3644 (N_3644,N_1599,N_2583);
and U3645 (N_3645,N_235,N_1184);
nand U3646 (N_3646,N_2669,N_1254);
or U3647 (N_3647,N_1755,N_5);
and U3648 (N_3648,N_1485,N_2867);
and U3649 (N_3649,N_2965,N_1145);
and U3650 (N_3650,N_1136,N_2275);
nand U3651 (N_3651,N_2951,N_1779);
nor U3652 (N_3652,N_2652,N_1992);
nor U3653 (N_3653,N_297,N_887);
nor U3654 (N_3654,N_1010,N_2713);
or U3655 (N_3655,N_780,N_2727);
nor U3656 (N_3656,N_143,N_42);
nand U3657 (N_3657,N_1154,N_1981);
or U3658 (N_3658,N_2189,N_2438);
nor U3659 (N_3659,N_2937,N_390);
or U3660 (N_3660,N_6,N_2894);
nand U3661 (N_3661,N_2744,N_1594);
or U3662 (N_3662,N_1400,N_1348);
and U3663 (N_3663,N_2530,N_2622);
or U3664 (N_3664,N_1231,N_2197);
or U3665 (N_3665,N_89,N_1026);
nor U3666 (N_3666,N_960,N_1967);
or U3667 (N_3667,N_2645,N_1881);
or U3668 (N_3668,N_2351,N_2300);
nand U3669 (N_3669,N_2537,N_157);
or U3670 (N_3670,N_1043,N_621);
and U3671 (N_3671,N_2711,N_2072);
or U3672 (N_3672,N_2540,N_2318);
nor U3673 (N_3673,N_1046,N_759);
nand U3674 (N_3674,N_1203,N_2362);
or U3675 (N_3675,N_1202,N_611);
or U3676 (N_3676,N_416,N_2970);
nor U3677 (N_3677,N_1631,N_2635);
nor U3678 (N_3678,N_713,N_752);
or U3679 (N_3679,N_992,N_2654);
nand U3680 (N_3680,N_1566,N_1527);
nand U3681 (N_3681,N_1571,N_940);
or U3682 (N_3682,N_608,N_2755);
nor U3683 (N_3683,N_1461,N_1081);
nor U3684 (N_3684,N_1304,N_1708);
or U3685 (N_3685,N_956,N_261);
nor U3686 (N_3686,N_2988,N_557);
nand U3687 (N_3687,N_1487,N_2553);
and U3688 (N_3688,N_172,N_80);
nor U3689 (N_3689,N_1020,N_8);
and U3690 (N_3690,N_2063,N_1789);
nor U3691 (N_3691,N_2213,N_2805);
or U3692 (N_3692,N_2788,N_2119);
or U3693 (N_3693,N_96,N_84);
nor U3694 (N_3694,N_1321,N_2355);
and U3695 (N_3695,N_1736,N_1080);
nor U3696 (N_3696,N_2044,N_1017);
nor U3697 (N_3697,N_1428,N_2960);
and U3698 (N_3698,N_394,N_1358);
or U3699 (N_3699,N_1160,N_925);
and U3700 (N_3700,N_750,N_2638);
and U3701 (N_3701,N_2365,N_2908);
nor U3702 (N_3702,N_2616,N_1193);
nor U3703 (N_3703,N_549,N_527);
nand U3704 (N_3704,N_610,N_522);
and U3705 (N_3705,N_2249,N_334);
nand U3706 (N_3706,N_2065,N_1904);
nor U3707 (N_3707,N_2427,N_977);
nor U3708 (N_3708,N_1486,N_0);
nor U3709 (N_3709,N_79,N_470);
or U3710 (N_3710,N_2678,N_2056);
nor U3711 (N_3711,N_1116,N_897);
and U3712 (N_3712,N_1930,N_2319);
or U3713 (N_3713,N_743,N_2799);
nand U3714 (N_3714,N_1771,N_2211);
and U3715 (N_3715,N_2712,N_2233);
and U3716 (N_3716,N_2996,N_948);
nor U3717 (N_3717,N_2655,N_2893);
nand U3718 (N_3718,N_2890,N_607);
or U3719 (N_3719,N_821,N_1421);
nand U3720 (N_3720,N_314,N_2959);
or U3721 (N_3721,N_2759,N_1867);
or U3722 (N_3722,N_2444,N_568);
nand U3723 (N_3723,N_2159,N_1672);
xor U3724 (N_3724,N_1651,N_88);
and U3725 (N_3725,N_174,N_818);
and U3726 (N_3726,N_258,N_757);
or U3727 (N_3727,N_1783,N_2636);
and U3728 (N_3728,N_1134,N_2765);
or U3729 (N_3729,N_2856,N_2508);
nand U3730 (N_3730,N_1556,N_2625);
or U3731 (N_3731,N_248,N_2236);
xor U3732 (N_3732,N_2498,N_1343);
nor U3733 (N_3733,N_1744,N_674);
nor U3734 (N_3734,N_1541,N_904);
and U3735 (N_3735,N_497,N_547);
nor U3736 (N_3736,N_2961,N_1388);
nand U3737 (N_3737,N_1280,N_2983);
and U3738 (N_3738,N_1627,N_2815);
nand U3739 (N_3739,N_2884,N_59);
and U3740 (N_3740,N_231,N_623);
nor U3741 (N_3741,N_101,N_1945);
nor U3742 (N_3742,N_2603,N_2926);
and U3743 (N_3743,N_2286,N_2601);
and U3744 (N_3744,N_2487,N_2522);
nor U3745 (N_3745,N_2955,N_1601);
or U3746 (N_3746,N_2595,N_2156);
or U3747 (N_3747,N_1533,N_2263);
and U3748 (N_3748,N_252,N_1138);
xnor U3749 (N_3749,N_1845,N_1398);
and U3750 (N_3750,N_2613,N_2208);
or U3751 (N_3751,N_1399,N_227);
nor U3752 (N_3752,N_443,N_385);
nand U3753 (N_3753,N_1122,N_1788);
or U3754 (N_3754,N_922,N_1130);
xnor U3755 (N_3755,N_1000,N_2760);
or U3756 (N_3756,N_1317,N_916);
and U3757 (N_3757,N_2933,N_2734);
and U3758 (N_3758,N_1308,N_2191);
nand U3759 (N_3759,N_2216,N_1336);
xnor U3760 (N_3760,N_755,N_280);
or U3761 (N_3761,N_605,N_1141);
nor U3762 (N_3762,N_2495,N_2146);
or U3763 (N_3763,N_1182,N_183);
nor U3764 (N_3764,N_1092,N_758);
nand U3765 (N_3765,N_1108,N_2657);
and U3766 (N_3766,N_685,N_2731);
nor U3767 (N_3767,N_2018,N_2769);
and U3768 (N_3768,N_187,N_810);
nor U3769 (N_3769,N_426,N_1061);
nor U3770 (N_3770,N_1717,N_1169);
nand U3771 (N_3771,N_680,N_412);
and U3772 (N_3772,N_2323,N_1110);
and U3773 (N_3773,N_1431,N_2696);
nor U3774 (N_3774,N_2743,N_873);
nand U3775 (N_3775,N_441,N_2344);
and U3776 (N_3776,N_1389,N_1492);
nor U3777 (N_3777,N_2093,N_1120);
or U3778 (N_3778,N_2576,N_737);
and U3779 (N_3779,N_1525,N_1052);
nor U3780 (N_3780,N_2594,N_2719);
and U3781 (N_3781,N_570,N_2504);
nand U3782 (N_3782,N_859,N_684);
or U3783 (N_3783,N_1039,N_86);
nor U3784 (N_3784,N_2864,N_47);
or U3785 (N_3785,N_1608,N_2845);
nand U3786 (N_3786,N_515,N_2250);
nand U3787 (N_3787,N_63,N_202);
nor U3788 (N_3788,N_303,N_206);
or U3789 (N_3789,N_693,N_270);
or U3790 (N_3790,N_722,N_1455);
or U3791 (N_3791,N_1018,N_475);
and U3792 (N_3792,N_2927,N_1270);
and U3793 (N_3793,N_785,N_2333);
nand U3794 (N_3794,N_1038,N_1694);
or U3795 (N_3795,N_381,N_1228);
nand U3796 (N_3796,N_2314,N_2068);
or U3797 (N_3797,N_2881,N_1683);
and U3798 (N_3798,N_872,N_214);
nor U3799 (N_3799,N_1850,N_1718);
nor U3800 (N_3800,N_1423,N_30);
nor U3801 (N_3801,N_2430,N_1999);
nand U3802 (N_3802,N_1132,N_85);
nor U3803 (N_3803,N_1102,N_2559);
or U3804 (N_3804,N_1449,N_1824);
nor U3805 (N_3805,N_921,N_619);
nand U3806 (N_3806,N_2354,N_2012);
nand U3807 (N_3807,N_2311,N_1841);
or U3808 (N_3808,N_2862,N_689);
xor U3809 (N_3809,N_2841,N_2739);
nand U3810 (N_3810,N_1383,N_481);
nor U3811 (N_3811,N_283,N_782);
nand U3812 (N_3812,N_2353,N_420);
or U3813 (N_3813,N_648,N_1952);
or U3814 (N_3814,N_909,N_477);
or U3815 (N_3815,N_2587,N_2259);
nand U3816 (N_3816,N_351,N_411);
nand U3817 (N_3817,N_1719,N_1863);
and U3818 (N_3818,N_805,N_126);
or U3819 (N_3819,N_2062,N_1540);
nor U3820 (N_3820,N_815,N_1104);
nand U3821 (N_3821,N_907,N_1983);
nand U3822 (N_3822,N_328,N_2649);
nand U3823 (N_3823,N_2327,N_1923);
nand U3824 (N_3824,N_1534,N_1071);
nand U3825 (N_3825,N_2331,N_2728);
and U3826 (N_3826,N_268,N_2265);
xor U3827 (N_3827,N_1643,N_1773);
nor U3828 (N_3828,N_1324,N_155);
and U3829 (N_3829,N_2511,N_1807);
or U3830 (N_3830,N_541,N_2826);
and U3831 (N_3831,N_2040,N_2535);
or U3832 (N_3832,N_1725,N_2592);
nand U3833 (N_3833,N_615,N_1625);
or U3834 (N_3834,N_827,N_333);
nor U3835 (N_3835,N_540,N_2347);
or U3836 (N_3836,N_1618,N_2950);
and U3837 (N_3837,N_1793,N_709);
xor U3838 (N_3838,N_1365,N_1413);
nand U3839 (N_3839,N_2693,N_2574);
nand U3840 (N_3840,N_996,N_296);
and U3841 (N_3841,N_664,N_1480);
nor U3842 (N_3842,N_2198,N_327);
or U3843 (N_3843,N_538,N_2269);
nand U3844 (N_3844,N_210,N_446);
or U3845 (N_3845,N_1629,N_2972);
nand U3846 (N_3846,N_991,N_1677);
or U3847 (N_3847,N_2366,N_1315);
and U3848 (N_3848,N_2866,N_2726);
nand U3849 (N_3849,N_1508,N_2944);
and U3850 (N_3850,N_1942,N_2525);
nor U3851 (N_3851,N_53,N_1782);
nand U3852 (N_3852,N_978,N_203);
nor U3853 (N_3853,N_2555,N_1152);
or U3854 (N_3854,N_1579,N_1656);
nand U3855 (N_3855,N_374,N_1310);
and U3856 (N_3856,N_398,N_1591);
and U3857 (N_3857,N_1044,N_2813);
and U3858 (N_3858,N_272,N_2772);
nand U3859 (N_3859,N_2873,N_1962);
and U3860 (N_3860,N_2443,N_1350);
and U3861 (N_3861,N_2456,N_1451);
or U3862 (N_3862,N_1300,N_683);
and U3863 (N_3863,N_1800,N_331);
and U3864 (N_3864,N_1316,N_1896);
nor U3865 (N_3865,N_1371,N_1133);
nand U3866 (N_3866,N_105,N_2200);
nor U3867 (N_3867,N_166,N_604);
and U3868 (N_3868,N_1360,N_1247);
or U3869 (N_3869,N_2808,N_145);
and U3870 (N_3870,N_2453,N_1620);
nor U3871 (N_3871,N_1250,N_936);
nand U3872 (N_3872,N_1762,N_2919);
and U3873 (N_3873,N_2067,N_770);
and U3874 (N_3874,N_2109,N_2771);
nor U3875 (N_3875,N_2123,N_1091);
and U3876 (N_3876,N_1688,N_918);
nor U3877 (N_3877,N_38,N_1616);
nor U3878 (N_3878,N_2393,N_1427);
nand U3879 (N_3879,N_1240,N_2371);
or U3880 (N_3880,N_659,N_1301);
or U3881 (N_3881,N_1943,N_2922);
nand U3882 (N_3882,N_274,N_428);
and U3883 (N_3883,N_1741,N_1848);
nor U3884 (N_3884,N_690,N_1532);
and U3885 (N_3885,N_2407,N_2078);
nand U3886 (N_3886,N_2425,N_1853);
or U3887 (N_3887,N_580,N_2105);
and U3888 (N_3888,N_923,N_947);
or U3889 (N_3889,N_320,N_137);
nand U3890 (N_3890,N_2834,N_2219);
and U3891 (N_3891,N_33,N_317);
or U3892 (N_3892,N_699,N_1922);
nor U3893 (N_3893,N_2935,N_2973);
nand U3894 (N_3894,N_2160,N_2861);
nor U3895 (N_3895,N_2000,N_1279);
nor U3896 (N_3896,N_373,N_1795);
nand U3897 (N_3897,N_140,N_2003);
nor U3898 (N_3898,N_2542,N_1791);
nand U3899 (N_3899,N_1379,N_1517);
and U3900 (N_3900,N_2185,N_943);
or U3901 (N_3901,N_1330,N_1306);
or U3902 (N_3902,N_1293,N_1109);
nor U3903 (N_3903,N_241,N_2474);
and U3904 (N_3904,N_635,N_1478);
and U3905 (N_3905,N_840,N_2229);
nor U3906 (N_3906,N_889,N_321);
nand U3907 (N_3907,N_2780,N_2614);
and U3908 (N_3908,N_2325,N_2287);
or U3909 (N_3909,N_1503,N_1781);
nor U3910 (N_3910,N_837,N_890);
or U3911 (N_3911,N_326,N_1309);
nand U3912 (N_3912,N_841,N_900);
and U3913 (N_3913,N_91,N_1912);
or U3914 (N_3914,N_168,N_1065);
and U3915 (N_3915,N_2207,N_926);
and U3916 (N_3916,N_724,N_2611);
nor U3917 (N_3917,N_73,N_1538);
xnor U3918 (N_3918,N_1803,N_1258);
and U3919 (N_3919,N_1940,N_116);
nand U3920 (N_3920,N_2482,N_1245);
or U3921 (N_3921,N_118,N_562);
or U3922 (N_3922,N_2085,N_115);
nand U3923 (N_3923,N_1149,N_2833);
nand U3924 (N_3924,N_1068,N_2575);
and U3925 (N_3925,N_2646,N_2011);
and U3926 (N_3926,N_348,N_2346);
or U3927 (N_3927,N_2593,N_2304);
or U3928 (N_3928,N_1271,N_2166);
or U3929 (N_3929,N_67,N_1323);
nor U3930 (N_3930,N_970,N_1481);
or U3931 (N_3931,N_2598,N_2397);
or U3932 (N_3932,N_1269,N_1214);
and U3933 (N_3933,N_578,N_1190);
nand U3934 (N_3934,N_1012,N_1216);
or U3935 (N_3935,N_1523,N_2664);
or U3936 (N_3936,N_434,N_965);
or U3937 (N_3937,N_2756,N_1989);
nand U3938 (N_3938,N_1667,N_139);
and U3939 (N_3939,N_1641,N_1758);
nor U3940 (N_3940,N_1504,N_2083);
or U3941 (N_3941,N_2174,N_712);
nor U3942 (N_3942,N_2677,N_72);
and U3943 (N_3943,N_1865,N_2561);
nor U3944 (N_3944,N_1021,N_1191);
nor U3945 (N_3945,N_337,N_1472);
or U3946 (N_3946,N_288,N_2717);
nor U3947 (N_3947,N_1019,N_2381);
and U3948 (N_3948,N_103,N_845);
nand U3949 (N_3949,N_1898,N_2046);
nor U3950 (N_3950,N_285,N_1448);
nand U3951 (N_3951,N_843,N_2876);
or U3952 (N_3952,N_2110,N_190);
nor U3953 (N_3953,N_2985,N_707);
and U3954 (N_3954,N_1815,N_589);
nand U3955 (N_3955,N_1264,N_688);
nand U3956 (N_3956,N_1529,N_1505);
nand U3957 (N_3957,N_2426,N_924);
or U3958 (N_3958,N_2163,N_528);
nand U3959 (N_3959,N_1939,N_976);
nand U3960 (N_3960,N_1595,N_1322);
nor U3961 (N_3961,N_347,N_842);
nand U3962 (N_3962,N_2050,N_2888);
xor U3963 (N_3963,N_2702,N_626);
xor U3964 (N_3964,N_340,N_1106);
nand U3965 (N_3965,N_1443,N_2982);
nor U3966 (N_3966,N_1391,N_1958);
nand U3967 (N_3967,N_2639,N_1597);
or U3968 (N_3968,N_1490,N_1189);
nand U3969 (N_3969,N_2465,N_1003);
and U3970 (N_3970,N_2221,N_555);
and U3971 (N_3971,N_2564,N_2662);
or U3972 (N_3972,N_603,N_2454);
nand U3973 (N_3973,N_1066,N_125);
and U3974 (N_3974,N_1899,N_692);
or U3975 (N_3975,N_876,N_2612);
and U3976 (N_3976,N_127,N_2989);
or U3977 (N_3977,N_1422,N_294);
and U3978 (N_3978,N_2607,N_2757);
nand U3979 (N_3979,N_2624,N_2838);
nand U3980 (N_3980,N_1030,N_2178);
and U3981 (N_3981,N_2199,N_816);
nor U3982 (N_3982,N_1674,N_2010);
and U3983 (N_3983,N_2883,N_78);
nor U3984 (N_3984,N_2672,N_1298);
nand U3985 (N_3985,N_1437,N_489);
nor U3986 (N_3986,N_1387,N_2152);
and U3987 (N_3987,N_1903,N_392);
nand U3988 (N_3988,N_120,N_1287);
or U3989 (N_3989,N_1592,N_236);
nand U3990 (N_3990,N_1022,N_1185);
nand U3991 (N_3991,N_2175,N_1023);
or U3992 (N_3992,N_513,N_2590);
nor U3993 (N_3993,N_1790,N_2076);
and U3994 (N_3994,N_2934,N_1403);
or U3995 (N_3995,N_48,N_888);
or U3996 (N_3996,N_679,N_1347);
or U3997 (N_3997,N_651,N_2104);
xnor U3998 (N_3998,N_369,N_1098);
nand U3999 (N_3999,N_1426,N_701);
nor U4000 (N_4000,N_450,N_492);
or U4001 (N_4001,N_2514,N_1565);
nand U4002 (N_4002,N_2513,N_1814);
nand U4003 (N_4003,N_867,N_2746);
nor U4004 (N_4004,N_868,N_2558);
or U4005 (N_4005,N_915,N_1219);
nor U4006 (N_4006,N_852,N_1701);
and U4007 (N_4007,N_1419,N_2488);
nand U4008 (N_4008,N_281,N_144);
nor U4009 (N_4009,N_731,N_2870);
and U4010 (N_4010,N_2871,N_199);
or U4011 (N_4011,N_2865,N_523);
or U4012 (N_4012,N_959,N_2289);
nor U4013 (N_4013,N_971,N_2543);
and U4014 (N_4014,N_2126,N_2721);
nand U4015 (N_4015,N_794,N_2114);
and U4016 (N_4016,N_2579,N_2570);
nor U4017 (N_4017,N_2648,N_2291);
or U4018 (N_4018,N_1260,N_196);
and U4019 (N_4019,N_1339,N_2102);
and U4020 (N_4020,N_1706,N_17);
or U4021 (N_4021,N_2489,N_2256);
and U4022 (N_4022,N_221,N_98);
nand U4023 (N_4023,N_905,N_354);
xnor U4024 (N_4024,N_1822,N_2827);
nor U4025 (N_4025,N_2633,N_2066);
or U4026 (N_4026,N_1965,N_2980);
or U4027 (N_4027,N_1087,N_2500);
or U4028 (N_4028,N_2019,N_164);
nor U4029 (N_4029,N_2816,N_1454);
and U4030 (N_4030,N_1871,N_1471);
nor U4031 (N_4031,N_625,N_1639);
and U4032 (N_4032,N_2173,N_324);
xnor U4033 (N_4033,N_2516,N_738);
and U4034 (N_4034,N_1596,N_2026);
and U4035 (N_4035,N_2899,N_2299);
nand U4036 (N_4036,N_171,N_587);
and U4037 (N_4037,N_2946,N_2911);
and U4038 (N_4038,N_963,N_2524);
nor U4039 (N_4039,N_1101,N_1804);
nand U4040 (N_4040,N_304,N_1915);
nand U4041 (N_4041,N_114,N_1528);
and U4042 (N_4042,N_1875,N_1861);
nand U4043 (N_4043,N_2247,N_2048);
nand U4044 (N_4044,N_530,N_483);
and U4045 (N_4045,N_1097,N_2245);
or U4046 (N_4046,N_511,N_1385);
and U4047 (N_4047,N_355,N_2134);
or U4048 (N_4048,N_1497,N_1031);
or U4049 (N_4049,N_1704,N_2534);
nand U4050 (N_4050,N_2629,N_663);
or U4051 (N_4051,N_2690,N_2502);
nor U4052 (N_4052,N_2811,N_2569);
xor U4053 (N_4053,N_1816,N_1148);
or U4054 (N_4054,N_2494,N_1557);
or U4055 (N_4055,N_2421,N_2963);
nand U4056 (N_4056,N_1359,N_1974);
nor U4057 (N_4057,N_122,N_886);
nand U4058 (N_4058,N_1811,N_2058);
or U4059 (N_4059,N_289,N_2206);
nand U4060 (N_4060,N_1187,N_1407);
and U4061 (N_4061,N_1555,N_37);
or U4062 (N_4062,N_205,N_1119);
nor U4063 (N_4063,N_1907,N_830);
and U4064 (N_4064,N_13,N_1295);
and U4065 (N_4065,N_128,N_2386);
and U4066 (N_4066,N_2402,N_1906);
and U4067 (N_4067,N_2157,N_346);
nor U4068 (N_4068,N_2383,N_1931);
nand U4069 (N_4069,N_1964,N_593);
nor U4070 (N_4070,N_35,N_1515);
or U4071 (N_4071,N_704,N_863);
or U4072 (N_4072,N_341,N_1584);
or U4073 (N_4073,N_1839,N_870);
nor U4074 (N_4074,N_2971,N_1253);
xor U4075 (N_4075,N_1142,N_2158);
nand U4076 (N_4076,N_2004,N_698);
or U4077 (N_4077,N_1827,N_1607);
nor U4078 (N_4078,N_961,N_1668);
or U4079 (N_4079,N_892,N_617);
nand U4080 (N_4080,N_2700,N_12);
or U4081 (N_4081,N_2458,N_2149);
nor U4082 (N_4082,N_2023,N_702);
or U4083 (N_4083,N_2180,N_2948);
nor U4084 (N_4084,N_1680,N_2997);
and U4085 (N_4085,N_1753,N_514);
xor U4086 (N_4086,N_2824,N_23);
nor U4087 (N_4087,N_1459,N_658);
nand U4088 (N_4088,N_1702,N_424);
or U4089 (N_4089,N_2519,N_2906);
nor U4090 (N_4090,N_806,N_1630);
or U4091 (N_4091,N_1941,N_2501);
and U4092 (N_4092,N_2181,N_2768);
and U4093 (N_4093,N_2670,N_1509);
nand U4094 (N_4094,N_1524,N_911);
nand U4095 (N_4095,N_2179,N_2187);
xor U4096 (N_4096,N_669,N_70);
or U4097 (N_4097,N_2703,N_1312);
nand U4098 (N_4098,N_1570,N_2092);
nand U4099 (N_4099,N_2747,N_2573);
and U4100 (N_4100,N_1910,N_1123);
nand U4101 (N_4101,N_238,N_1986);
and U4102 (N_4102,N_1284,N_1223);
xnor U4103 (N_4103,N_2581,N_1334);
xor U4104 (N_4104,N_2775,N_2271);
xor U4105 (N_4105,N_1578,N_2419);
or U4106 (N_4106,N_2033,N_1118);
or U4107 (N_4107,N_1395,N_1243);
or U4108 (N_4108,N_894,N_1392);
or U4109 (N_4109,N_2121,N_1809);
nand U4110 (N_4110,N_433,N_1679);
nor U4111 (N_4111,N_2260,N_121);
nor U4112 (N_4112,N_186,N_913);
nand U4113 (N_4113,N_360,N_2235);
nand U4114 (N_4114,N_677,N_929);
or U4115 (N_4115,N_2691,N_2380);
nand U4116 (N_4116,N_932,N_1587);
or U4117 (N_4117,N_613,N_1676);
or U4118 (N_4118,N_29,N_2082);
or U4119 (N_4119,N_1775,N_1354);
nand U4120 (N_4120,N_2599,N_403);
or U4121 (N_4121,N_1222,N_643);
nand U4122 (N_4122,N_706,N_1340);
nand U4123 (N_4123,N_773,N_2223);
nor U4124 (N_4124,N_1552,N_188);
xor U4125 (N_4125,N_2373,N_524);
nand U4126 (N_4126,N_537,N_1196);
or U4127 (N_4127,N_191,N_2384);
nand U4128 (N_4128,N_958,N_2966);
or U4129 (N_4129,N_1553,N_15);
or U4130 (N_4130,N_2609,N_159);
or U4131 (N_4131,N_133,N_2288);
nand U4132 (N_4132,N_741,N_1662);
nor U4133 (N_4133,N_769,N_2875);
and U4134 (N_4134,N_1609,N_2330);
nand U4135 (N_4135,N_2803,N_1794);
or U4136 (N_4136,N_368,N_2435);
nor U4137 (N_4137,N_1040,N_2736);
or U4138 (N_4138,N_1,N_2665);
nor U4139 (N_4139,N_1536,N_463);
and U4140 (N_4140,N_2889,N_2336);
and U4141 (N_4141,N_1006,N_1464);
and U4142 (N_4142,N_2061,N_2674);
nand U4143 (N_4143,N_2032,N_2754);
and U4144 (N_4144,N_2238,N_1589);
nor U4145 (N_4145,N_1738,N_1005);
or U4146 (N_4146,N_1707,N_1212);
nand U4147 (N_4147,N_819,N_700);
nand U4148 (N_4148,N_356,N_1926);
and U4149 (N_4149,N_1600,N_2637);
or U4150 (N_4150,N_1661,N_1984);
or U4151 (N_4151,N_1995,N_62);
nand U4152 (N_4152,N_246,N_2272);
and U4153 (N_4153,N_2509,N_2022);
or U4154 (N_4154,N_2411,N_1498);
or U4155 (N_4155,N_22,N_2632);
nor U4156 (N_4156,N_363,N_1720);
or U4157 (N_4157,N_2266,N_1115);
nand U4158 (N_4158,N_1289,N_132);
nand U4159 (N_4159,N_767,N_793);
or U4160 (N_4160,N_1918,N_1496);
or U4161 (N_4161,N_2722,N_931);
or U4162 (N_4162,N_829,N_848);
nor U4163 (N_4163,N_117,N_1095);
nand U4164 (N_4164,N_1750,N_2222);
nand U4165 (N_4165,N_2361,N_1070);
or U4166 (N_4166,N_2133,N_1099);
or U4167 (N_4167,N_710,N_445);
nor U4168 (N_4168,N_1954,N_2490);
nand U4169 (N_4169,N_1073,N_1177);
nand U4170 (N_4170,N_419,N_2151);
or U4171 (N_4171,N_2280,N_1648);
or U4172 (N_4172,N_2182,N_149);
and U4173 (N_4173,N_399,N_2408);
nand U4174 (N_4174,N_1747,N_732);
nand U4175 (N_4175,N_949,N_1615);
nor U4176 (N_4176,N_2293,N_1206);
nor U4177 (N_4177,N_2462,N_2047);
xor U4178 (N_4178,N_1314,N_585);
nand U4179 (N_4179,N_1215,N_1439);
and U4180 (N_4180,N_2751,N_1739);
nor U4181 (N_4181,N_2551,N_2978);
and U4182 (N_4182,N_2708,N_1914);
nand U4183 (N_4183,N_670,N_2931);
nand U4184 (N_4184,N_2363,N_2227);
nor U4185 (N_4185,N_2115,N_790);
and U4186 (N_4186,N_1586,N_1526);
nand U4187 (N_4187,N_1645,N_574);
nand U4188 (N_4188,N_1166,N_466);
nor U4189 (N_4189,N_1456,N_2918);
nor U4190 (N_4190,N_409,N_2986);
and U4191 (N_4191,N_590,N_1139);
and U4192 (N_4192,N_2253,N_1302);
or U4193 (N_4193,N_744,N_997);
or U4194 (N_4194,N_1721,N_2087);
nand U4195 (N_4195,N_2661,N_2240);
or U4196 (N_4196,N_61,N_866);
nand U4197 (N_4197,N_899,N_49);
and U4198 (N_4198,N_935,N_2051);
or U4199 (N_4199,N_2923,N_774);
nand U4200 (N_4200,N_2002,N_1539);
nor U4201 (N_4201,N_1048,N_814);
nor U4202 (N_4202,N_2329,N_1059);
nor U4203 (N_4203,N_1715,N_452);
nor U4204 (N_4204,N_1564,N_1975);
nand U4205 (N_4205,N_2916,N_803);
nand U4206 (N_4206,N_934,N_2658);
nand U4207 (N_4207,N_134,N_2137);
and U4208 (N_4208,N_1255,N_1520);
nand U4209 (N_4209,N_2268,N_1344);
nand U4210 (N_4210,N_1866,N_715);
or U4211 (N_4211,N_1463,N_2729);
and U4212 (N_4212,N_1311,N_93);
nand U4213 (N_4213,N_332,N_1337);
or U4214 (N_4214,N_2448,N_2324);
or U4215 (N_4215,N_1062,N_1917);
or U4216 (N_4216,N_269,N_2243);
nor U4217 (N_4217,N_1476,N_2925);
nor U4218 (N_4218,N_666,N_391);
and U4219 (N_4219,N_896,N_1684);
nor U4220 (N_4220,N_1900,N_367);
or U4221 (N_4221,N_1979,N_2954);
nor U4222 (N_4222,N_192,N_1821);
nand U4223 (N_4223,N_967,N_520);
nand U4224 (N_4224,N_2860,N_10);
nor U4225 (N_4225,N_776,N_2309);
or U4226 (N_4226,N_653,N_599);
or U4227 (N_4227,N_1949,N_349);
nor U4228 (N_4228,N_882,N_1996);
nor U4229 (N_4229,N_1495,N_2254);
nand U4230 (N_4230,N_885,N_895);
or U4231 (N_4231,N_828,N_1057);
nor U4232 (N_4232,N_2682,N_3);
and U4233 (N_4233,N_2819,N_1864);
nand U4234 (N_4234,N_2550,N_228);
and U4235 (N_4235,N_142,N_503);
nor U4236 (N_4236,N_2112,N_1424);
and U4237 (N_4237,N_239,N_2853);
and U4238 (N_4238,N_508,N_2710);
nor U4239 (N_4239,N_226,N_1709);
nand U4240 (N_4240,N_421,N_1892);
and U4241 (N_4241,N_865,N_1734);
or U4242 (N_4242,N_2389,N_2169);
or U4243 (N_4243,N_1829,N_1396);
and U4244 (N_4244,N_542,N_642);
nand U4245 (N_4245,N_2733,N_1727);
nand U4246 (N_4246,N_938,N_2770);
nor U4247 (N_4247,N_1572,N_582);
and U4248 (N_4248,N_2095,N_964);
or U4249 (N_4249,N_2099,N_2097);
nand U4250 (N_4250,N_1929,N_844);
nor U4251 (N_4251,N_1432,N_1649);
nand U4252 (N_4252,N_864,N_2806);
nand U4253 (N_4253,N_1670,N_2144);
or U4254 (N_4254,N_2699,N_2279);
and U4255 (N_4255,N_1957,N_2829);
nor U4256 (N_4256,N_1248,N_1088);
and U4257 (N_4257,N_2953,N_1786);
xnor U4258 (N_4258,N_826,N_518);
nor U4259 (N_4259,N_2763,N_898);
and U4260 (N_4260,N_2958,N_2932);
nand U4261 (N_4261,N_2847,N_110);
nand U4262 (N_4262,N_1100,N_912);
or U4263 (N_4263,N_660,N_2901);
nand U4264 (N_4264,N_2567,N_1470);
nor U4265 (N_4265,N_1429,N_358);
xor U4266 (N_4266,N_2673,N_1394);
nor U4267 (N_4267,N_2290,N_2556);
or U4268 (N_4268,N_2518,N_1972);
nor U4269 (N_4269,N_1857,N_266);
nand U4270 (N_4270,N_275,N_2538);
nor U4271 (N_4271,N_552,N_2116);
nand U4272 (N_4272,N_836,N_2783);
and U4273 (N_4273,N_1125,N_167);
nor U4274 (N_4274,N_2338,N_1879);
nand U4275 (N_4275,N_2101,N_2242);
and U4276 (N_4276,N_2749,N_2090);
or U4277 (N_4277,N_1692,N_2914);
and U4278 (N_4278,N_857,N_1673);
or U4279 (N_4279,N_968,N_343);
nor U4280 (N_4280,N_766,N_2684);
or U4281 (N_4281,N_1658,N_264);
nand U4282 (N_4282,N_1192,N_2070);
nor U4283 (N_4283,N_2084,N_2778);
or U4284 (N_4284,N_1733,N_400);
nor U4285 (N_4285,N_138,N_2007);
nand U4286 (N_4286,N_1754,N_560);
and U4287 (N_4287,N_2429,N_2074);
or U4288 (N_4288,N_1978,N_2630);
nand U4289 (N_4289,N_1162,N_1851);
or U4290 (N_4290,N_1686,N_969);
and U4291 (N_4291,N_1016,N_675);
nand U4292 (N_4292,N_2025,N_1977);
nand U4293 (N_4293,N_2165,N_249);
and U4294 (N_4294,N_2195,N_788);
nor U4295 (N_4295,N_2604,N_1581);
nand U4296 (N_4296,N_2962,N_2258);
and U4297 (N_4297,N_860,N_97);
nor U4298 (N_4298,N_1510,N_2589);
nor U4299 (N_4299,N_1418,N_944);
xor U4300 (N_4300,N_1590,N_153);
and U4301 (N_4301,N_747,N_189);
nand U4302 (N_4302,N_180,N_1516);
nand U4303 (N_4303,N_51,N_1844);
or U4304 (N_4304,N_644,N_1143);
and U4305 (N_4305,N_2089,N_2292);
nand U4306 (N_4306,N_56,N_193);
and U4307 (N_4307,N_554,N_396);
nand U4308 (N_4308,N_1705,N_820);
or U4309 (N_4309,N_979,N_2800);
or U4310 (N_4310,N_2252,N_1513);
nand U4311 (N_4311,N_1697,N_2762);
xnor U4312 (N_4312,N_2969,N_2584);
nor U4313 (N_4313,N_1937,N_2239);
nor U4314 (N_4314,N_534,N_501);
xor U4315 (N_4315,N_2679,N_310);
nor U4316 (N_4316,N_1377,N_2825);
and U4317 (N_4317,N_2634,N_2369);
or U4318 (N_4318,N_1835,N_2872);
nand U4319 (N_4319,N_1549,N_219);
nand U4320 (N_4320,N_850,N_151);
xnor U4321 (N_4321,N_2107,N_2623);
or U4322 (N_4322,N_1366,N_2103);
or U4323 (N_4323,N_2320,N_1512);
and U4324 (N_4324,N_1417,N_1488);
and U4325 (N_4325,N_1244,N_1079);
nand U4326 (N_4326,N_1785,N_1153);
nor U4327 (N_4327,N_2403,N_1165);
nor U4328 (N_4328,N_858,N_1176);
nor U4329 (N_4329,N_136,N_561);
and U4330 (N_4330,N_2481,N_2475);
or U4331 (N_4331,N_444,N_1445);
or U4332 (N_4332,N_2640,N_2577);
and U4333 (N_4333,N_2964,N_779);
or U4334 (N_4334,N_2705,N_2278);
nand U4335 (N_4335,N_1430,N_1514);
or U4336 (N_4336,N_1968,N_1994);
nor U4337 (N_4337,N_135,N_1036);
nand U4338 (N_4338,N_2277,N_691);
nor U4339 (N_4339,N_2697,N_1085);
or U4340 (N_4340,N_881,N_1415);
nor U4341 (N_4341,N_427,N_2073);
and U4342 (N_4342,N_1703,N_2695);
and U4343 (N_4343,N_179,N_2863);
nor U4344 (N_4344,N_2723,N_2849);
and U4345 (N_4345,N_551,N_2898);
nor U4346 (N_4346,N_1767,N_150);
nor U4347 (N_4347,N_330,N_1207);
nand U4348 (N_4348,N_1563,N_588);
nand U4349 (N_4349,N_55,N_2155);
or U4350 (N_4350,N_389,N_18);
or U4351 (N_4351,N_185,N_2202);
nand U4352 (N_4352,N_989,N_493);
nor U4353 (N_4353,N_1885,N_459);
nor U4354 (N_4354,N_2359,N_2450);
or U4355 (N_4355,N_1482,N_2605);
or U4356 (N_4356,N_1235,N_1730);
and U4357 (N_4357,N_546,N_1888);
nor U4358 (N_4358,N_322,N_2835);
or U4359 (N_4359,N_1833,N_2896);
or U4360 (N_4360,N_2192,N_983);
nor U4361 (N_4361,N_311,N_942);
or U4362 (N_4362,N_624,N_1171);
or U4363 (N_4363,N_2724,N_2257);
nor U4364 (N_4364,N_1714,N_2820);
or U4365 (N_4365,N_2441,N_1924);
and U4366 (N_4366,N_1285,N_789);
nor U4367 (N_4367,N_1893,N_1002);
and U4368 (N_4368,N_45,N_795);
nand U4369 (N_4369,N_26,N_1908);
and U4370 (N_4370,N_2406,N_1457);
nor U4371 (N_4371,N_232,N_370);
nor U4372 (N_4372,N_2091,N_2874);
nand U4373 (N_4373,N_1241,N_1948);
nor U4374 (N_4374,N_1050,N_2168);
nor U4375 (N_4375,N_415,N_1390);
nor U4376 (N_4376,N_2610,N_60);
nor U4377 (N_4377,N_184,N_939);
nand U4378 (N_4378,N_2830,N_46);
xnor U4379 (N_4379,N_657,N_1872);
nand U4380 (N_4380,N_600,N_1150);
nor U4381 (N_4381,N_305,N_714);
or U4382 (N_4382,N_584,N_1970);
and U4383 (N_4383,N_1146,N_649);
nand U4384 (N_4384,N_1634,N_124);
nand U4385 (N_4385,N_1760,N_181);
xnor U4386 (N_4386,N_686,N_329);
and U4387 (N_4387,N_2294,N_451);
nand U4388 (N_4388,N_883,N_220);
nor U4389 (N_4389,N_307,N_510);
and U4390 (N_4390,N_2842,N_641);
nand U4391 (N_4391,N_54,N_1204);
nand U4392 (N_4392,N_366,N_2868);
and U4393 (N_4393,N_1731,N_1170);
nand U4394 (N_4394,N_1224,N_1770);
or U4395 (N_4395,N_2262,N_2401);
or U4396 (N_4396,N_1434,N_2039);
or U4397 (N_4397,N_2903,N_1574);
nor U4398 (N_4398,N_1691,N_1211);
nand U4399 (N_4399,N_146,N_1602);
and U4400 (N_4400,N_2139,N_1796);
nor U4401 (N_4401,N_2831,N_2217);
or U4402 (N_4402,N_2620,N_457);
xnor U4403 (N_4403,N_2660,N_1008);
and U4404 (N_4404,N_1780,N_536);
nor U4405 (N_4405,N_109,N_413);
and U4406 (N_4406,N_2027,N_2750);
nor U4407 (N_4407,N_2582,N_2758);
nand U4408 (N_4408,N_1585,N_1660);
nand U4409 (N_4409,N_1161,N_215);
nand U4410 (N_4410,N_2794,N_2364);
and U4411 (N_4411,N_1847,N_1096);
and U4412 (N_4412,N_175,N_2466);
nand U4413 (N_4413,N_1960,N_2183);
nor U4414 (N_4414,N_994,N_728);
or U4415 (N_4415,N_1617,N_1331);
nor U4416 (N_4416,N_563,N_2203);
and U4417 (N_4417,N_917,N_2821);
or U4418 (N_4418,N_431,N_2791);
nand U4419 (N_4419,N_7,N_2774);
nor U4420 (N_4420,N_569,N_2176);
nor U4421 (N_4421,N_1406,N_2377);
nand U4422 (N_4422,N_2308,N_2248);
or U4423 (N_4423,N_1671,N_2005);
nor U4424 (N_4424,N_1687,N_1221);
and U4425 (N_4425,N_1047,N_594);
nor U4426 (N_4426,N_1105,N_544);
nor U4427 (N_4427,N_1156,N_1500);
and U4428 (N_4428,N_460,N_869);
nor U4429 (N_4429,N_2942,N_1869);
nor U4430 (N_4430,N_507,N_1985);
and U4431 (N_4431,N_2676,N_2367);
nand U4432 (N_4432,N_1823,N_1825);
and U4433 (N_4433,N_2021,N_352);
and U4434 (N_4434,N_990,N_1663);
xnor U4435 (N_4435,N_2194,N_1723);
nand U4436 (N_4436,N_637,N_2313);
and U4437 (N_4437,N_1614,N_87);
nor U4438 (N_4438,N_222,N_1180);
nand U4439 (N_4439,N_1305,N_2882);
nand U4440 (N_4440,N_705,N_2232);
nand U4441 (N_4441,N_1537,N_634);
and U4442 (N_4442,N_2680,N_437);
nand U4443 (N_4443,N_1873,N_323);
or U4444 (N_4444,N_1194,N_2036);
or U4445 (N_4445,N_2745,N_1693);
and U4446 (N_4446,N_1272,N_2321);
nand U4447 (N_4447,N_2656,N_2261);
nor U4448 (N_4448,N_2154,N_161);
nor U4449 (N_4449,N_2943,N_313);
nand U4450 (N_4450,N_130,N_941);
nand U4451 (N_4451,N_1089,N_1860);
or U4452 (N_4452,N_1473,N_1868);
or U4453 (N_4453,N_1256,N_1685);
and U4454 (N_4454,N_1188,N_1054);
nand U4455 (N_4455,N_2653,N_2035);
and U4456 (N_4456,N_631,N_1856);
nor U4457 (N_4457,N_240,N_2108);
nor U4458 (N_4458,N_405,N_2976);
and U4459 (N_4459,N_1209,N_2571);
nand U4460 (N_4460,N_2388,N_656);
nor U4461 (N_4461,N_66,N_2423);
nand U4462 (N_4462,N_2034,N_211);
nor U4463 (N_4463,N_1408,N_1695);
nand U4464 (N_4464,N_1210,N_2523);
nand U4465 (N_4465,N_2557,N_2885);
nand U4466 (N_4466,N_1568,N_480);
nand U4467 (N_4467,N_760,N_2410);
and U4468 (N_4468,N_1029,N_878);
and U4469 (N_4469,N_745,N_2470);
nor U4470 (N_4470,N_835,N_2283);
nand U4471 (N_4471,N_2130,N_1928);
nand U4472 (N_4472,N_1647,N_57);
or U4473 (N_4473,N_2764,N_854);
or U4474 (N_4474,N_438,N_1033);
nor U4475 (N_4475,N_2374,N_1126);
or U4476 (N_4476,N_2659,N_217);
xnor U4477 (N_4477,N_1282,N_718);
nor U4478 (N_4478,N_2787,N_628);
nand U4479 (N_4479,N_2360,N_1233);
nor U4480 (N_4480,N_1361,N_2797);
nor U4481 (N_4481,N_2136,N_2343);
and U4482 (N_4482,N_393,N_1511);
nor U4483 (N_4483,N_786,N_2053);
or U4484 (N_4484,N_1843,N_11);
and U4485 (N_4485,N_1227,N_245);
nor U4486 (N_4486,N_1409,N_81);
or U4487 (N_4487,N_1278,N_2220);
nor U4488 (N_4488,N_612,N_1891);
or U4489 (N_4489,N_1880,N_2230);
nand U4490 (N_4490,N_2795,N_1593);
nand U4491 (N_4491,N_1982,N_671);
nand U4492 (N_4492,N_591,N_458);
and U4493 (N_4493,N_1263,N_279);
nor U4494 (N_4494,N_2692,N_1479);
or U4495 (N_4495,N_478,N_336);
nor U4496 (N_4496,N_2413,N_1506);
or U4497 (N_4497,N_1405,N_1742);
nor U4498 (N_4498,N_418,N_2312);
nor U4499 (N_4499,N_154,N_595);
or U4500 (N_4500,N_1,N_1533);
nor U4501 (N_4501,N_774,N_499);
nand U4502 (N_4502,N_542,N_2941);
nand U4503 (N_4503,N_1854,N_2265);
or U4504 (N_4504,N_262,N_1939);
nor U4505 (N_4505,N_184,N_1566);
nor U4506 (N_4506,N_1950,N_1877);
nor U4507 (N_4507,N_2858,N_606);
or U4508 (N_4508,N_2913,N_877);
nand U4509 (N_4509,N_1689,N_1064);
nand U4510 (N_4510,N_454,N_2438);
nor U4511 (N_4511,N_3,N_1634);
xnor U4512 (N_4512,N_1603,N_807);
nor U4513 (N_4513,N_580,N_1792);
nand U4514 (N_4514,N_2949,N_2596);
nor U4515 (N_4515,N_552,N_2135);
nand U4516 (N_4516,N_2500,N_2714);
nand U4517 (N_4517,N_1952,N_2166);
or U4518 (N_4518,N_1072,N_1447);
nand U4519 (N_4519,N_2963,N_2304);
and U4520 (N_4520,N_2999,N_2324);
nor U4521 (N_4521,N_2133,N_1428);
or U4522 (N_4522,N_646,N_1685);
xnor U4523 (N_4523,N_2136,N_831);
xnor U4524 (N_4524,N_955,N_2693);
nand U4525 (N_4525,N_2496,N_2305);
and U4526 (N_4526,N_2927,N_1468);
xor U4527 (N_4527,N_1188,N_2165);
nor U4528 (N_4528,N_1924,N_1838);
nand U4529 (N_4529,N_1641,N_513);
or U4530 (N_4530,N_2987,N_2216);
nor U4531 (N_4531,N_394,N_2754);
and U4532 (N_4532,N_1384,N_1756);
or U4533 (N_4533,N_2636,N_1124);
or U4534 (N_4534,N_1428,N_1265);
nand U4535 (N_4535,N_1091,N_1122);
nand U4536 (N_4536,N_2172,N_725);
or U4537 (N_4537,N_1577,N_2589);
nand U4538 (N_4538,N_536,N_2563);
or U4539 (N_4539,N_898,N_2140);
nor U4540 (N_4540,N_1448,N_2611);
nor U4541 (N_4541,N_726,N_1707);
nor U4542 (N_4542,N_1001,N_2907);
and U4543 (N_4543,N_2036,N_1590);
nand U4544 (N_4544,N_851,N_2561);
or U4545 (N_4545,N_1834,N_2359);
or U4546 (N_4546,N_2867,N_2883);
nand U4547 (N_4547,N_2611,N_1615);
nor U4548 (N_4548,N_1292,N_2270);
xor U4549 (N_4549,N_2232,N_2759);
or U4550 (N_4550,N_299,N_489);
and U4551 (N_4551,N_1563,N_246);
or U4552 (N_4552,N_1615,N_123);
nand U4553 (N_4553,N_722,N_25);
xnor U4554 (N_4554,N_2586,N_1425);
nor U4555 (N_4555,N_664,N_2237);
or U4556 (N_4556,N_1182,N_2407);
nor U4557 (N_4557,N_2000,N_2562);
and U4558 (N_4558,N_1980,N_1730);
or U4559 (N_4559,N_881,N_795);
nand U4560 (N_4560,N_43,N_399);
nor U4561 (N_4561,N_2801,N_1597);
nand U4562 (N_4562,N_428,N_1794);
and U4563 (N_4563,N_1590,N_2312);
nand U4564 (N_4564,N_804,N_407);
nor U4565 (N_4565,N_1884,N_1039);
nand U4566 (N_4566,N_141,N_1847);
and U4567 (N_4567,N_2943,N_1883);
and U4568 (N_4568,N_1291,N_121);
or U4569 (N_4569,N_1760,N_850);
or U4570 (N_4570,N_433,N_641);
nor U4571 (N_4571,N_1601,N_2608);
nor U4572 (N_4572,N_2335,N_564);
and U4573 (N_4573,N_711,N_733);
nor U4574 (N_4574,N_1554,N_893);
nand U4575 (N_4575,N_1307,N_2801);
or U4576 (N_4576,N_738,N_1089);
xnor U4577 (N_4577,N_898,N_2754);
and U4578 (N_4578,N_1041,N_1935);
and U4579 (N_4579,N_480,N_1718);
and U4580 (N_4580,N_39,N_2074);
nor U4581 (N_4581,N_988,N_960);
nand U4582 (N_4582,N_2769,N_388);
nand U4583 (N_4583,N_99,N_2014);
and U4584 (N_4584,N_1077,N_702);
or U4585 (N_4585,N_547,N_1973);
nor U4586 (N_4586,N_2171,N_1146);
xor U4587 (N_4587,N_476,N_1421);
and U4588 (N_4588,N_1484,N_2331);
and U4589 (N_4589,N_2592,N_43);
nand U4590 (N_4590,N_318,N_1601);
nand U4591 (N_4591,N_2893,N_314);
or U4592 (N_4592,N_167,N_629);
and U4593 (N_4593,N_1477,N_2498);
nor U4594 (N_4594,N_782,N_844);
or U4595 (N_4595,N_48,N_2235);
and U4596 (N_4596,N_2982,N_1293);
or U4597 (N_4597,N_246,N_2186);
or U4598 (N_4598,N_663,N_1665);
xor U4599 (N_4599,N_2640,N_273);
nor U4600 (N_4600,N_622,N_2442);
nand U4601 (N_4601,N_2396,N_367);
nand U4602 (N_4602,N_1498,N_2905);
nand U4603 (N_4603,N_1671,N_1841);
nand U4604 (N_4604,N_2072,N_2263);
and U4605 (N_4605,N_2151,N_224);
and U4606 (N_4606,N_2509,N_2444);
and U4607 (N_4607,N_2133,N_1244);
nor U4608 (N_4608,N_260,N_2513);
or U4609 (N_4609,N_554,N_2373);
nand U4610 (N_4610,N_1846,N_1896);
nand U4611 (N_4611,N_340,N_2834);
and U4612 (N_4612,N_208,N_1823);
or U4613 (N_4613,N_2820,N_666);
nand U4614 (N_4614,N_439,N_1493);
or U4615 (N_4615,N_1525,N_309);
or U4616 (N_4616,N_424,N_1749);
and U4617 (N_4617,N_1060,N_2090);
nor U4618 (N_4618,N_1728,N_799);
nor U4619 (N_4619,N_2822,N_872);
or U4620 (N_4620,N_2016,N_24);
or U4621 (N_4621,N_438,N_1611);
xnor U4622 (N_4622,N_102,N_929);
and U4623 (N_4623,N_783,N_1443);
nor U4624 (N_4624,N_1677,N_1416);
nand U4625 (N_4625,N_1183,N_48);
nand U4626 (N_4626,N_896,N_1932);
nand U4627 (N_4627,N_1280,N_602);
and U4628 (N_4628,N_2709,N_1473);
nand U4629 (N_4629,N_873,N_2711);
nand U4630 (N_4630,N_1798,N_2620);
nand U4631 (N_4631,N_2071,N_2903);
nand U4632 (N_4632,N_1483,N_650);
nor U4633 (N_4633,N_2895,N_1879);
nor U4634 (N_4634,N_1402,N_1401);
and U4635 (N_4635,N_1131,N_532);
nor U4636 (N_4636,N_841,N_1551);
nor U4637 (N_4637,N_2499,N_36);
nand U4638 (N_4638,N_2090,N_2614);
or U4639 (N_4639,N_766,N_2885);
nor U4640 (N_4640,N_91,N_1620);
or U4641 (N_4641,N_2284,N_1243);
and U4642 (N_4642,N_2132,N_1007);
nor U4643 (N_4643,N_1533,N_2495);
nand U4644 (N_4644,N_2824,N_708);
and U4645 (N_4645,N_971,N_2366);
or U4646 (N_4646,N_2994,N_2089);
nand U4647 (N_4647,N_296,N_1245);
and U4648 (N_4648,N_731,N_1618);
or U4649 (N_4649,N_916,N_294);
nor U4650 (N_4650,N_1296,N_780);
nand U4651 (N_4651,N_222,N_2956);
nor U4652 (N_4652,N_1163,N_117);
nor U4653 (N_4653,N_1976,N_2113);
nor U4654 (N_4654,N_1234,N_2376);
or U4655 (N_4655,N_683,N_1012);
nand U4656 (N_4656,N_1185,N_2249);
nor U4657 (N_4657,N_2554,N_1015);
or U4658 (N_4658,N_1181,N_2116);
or U4659 (N_4659,N_275,N_1285);
nor U4660 (N_4660,N_1143,N_852);
or U4661 (N_4661,N_2670,N_460);
nand U4662 (N_4662,N_97,N_2084);
nand U4663 (N_4663,N_543,N_951);
nand U4664 (N_4664,N_1684,N_2325);
nand U4665 (N_4665,N_561,N_2880);
nor U4666 (N_4666,N_1159,N_2082);
and U4667 (N_4667,N_1455,N_897);
or U4668 (N_4668,N_1868,N_1663);
nor U4669 (N_4669,N_1485,N_22);
nor U4670 (N_4670,N_2245,N_720);
or U4671 (N_4671,N_1734,N_2326);
nor U4672 (N_4672,N_1286,N_2394);
or U4673 (N_4673,N_551,N_220);
and U4674 (N_4674,N_999,N_2043);
nand U4675 (N_4675,N_57,N_2197);
nor U4676 (N_4676,N_2321,N_29);
or U4677 (N_4677,N_1831,N_2321);
nor U4678 (N_4678,N_1698,N_2628);
and U4679 (N_4679,N_382,N_1747);
and U4680 (N_4680,N_2095,N_277);
nor U4681 (N_4681,N_1696,N_302);
nand U4682 (N_4682,N_468,N_1455);
xnor U4683 (N_4683,N_9,N_1394);
and U4684 (N_4684,N_1447,N_2529);
nand U4685 (N_4685,N_2723,N_1285);
or U4686 (N_4686,N_182,N_940);
nor U4687 (N_4687,N_1495,N_1131);
nand U4688 (N_4688,N_2447,N_1291);
xnor U4689 (N_4689,N_803,N_1784);
nor U4690 (N_4690,N_1495,N_2835);
nor U4691 (N_4691,N_1982,N_1483);
nand U4692 (N_4692,N_2343,N_2728);
and U4693 (N_4693,N_1072,N_2915);
and U4694 (N_4694,N_777,N_2519);
nor U4695 (N_4695,N_2221,N_2637);
or U4696 (N_4696,N_1212,N_2292);
or U4697 (N_4697,N_592,N_141);
nand U4698 (N_4698,N_2460,N_591);
or U4699 (N_4699,N_1051,N_46);
and U4700 (N_4700,N_2353,N_2989);
nand U4701 (N_4701,N_1802,N_1656);
or U4702 (N_4702,N_1820,N_696);
nand U4703 (N_4703,N_709,N_1037);
nor U4704 (N_4704,N_1562,N_699);
and U4705 (N_4705,N_2415,N_1388);
or U4706 (N_4706,N_2898,N_1238);
and U4707 (N_4707,N_233,N_172);
or U4708 (N_4708,N_796,N_1174);
nor U4709 (N_4709,N_1079,N_2866);
and U4710 (N_4710,N_376,N_737);
nor U4711 (N_4711,N_160,N_2742);
nand U4712 (N_4712,N_2724,N_2427);
and U4713 (N_4713,N_679,N_978);
and U4714 (N_4714,N_581,N_1428);
nand U4715 (N_4715,N_1409,N_98);
or U4716 (N_4716,N_2959,N_2126);
and U4717 (N_4717,N_1461,N_1253);
nand U4718 (N_4718,N_1025,N_2917);
nor U4719 (N_4719,N_2290,N_2196);
and U4720 (N_4720,N_2844,N_1639);
or U4721 (N_4721,N_2925,N_2244);
nor U4722 (N_4722,N_614,N_2525);
nand U4723 (N_4723,N_2095,N_1760);
nor U4724 (N_4724,N_1227,N_1215);
nor U4725 (N_4725,N_2702,N_1935);
nor U4726 (N_4726,N_149,N_2465);
nor U4727 (N_4727,N_415,N_992);
nand U4728 (N_4728,N_1228,N_2378);
and U4729 (N_4729,N_2498,N_1570);
nor U4730 (N_4730,N_2386,N_1391);
and U4731 (N_4731,N_1071,N_2170);
xnor U4732 (N_4732,N_751,N_1132);
nor U4733 (N_4733,N_2974,N_2954);
or U4734 (N_4734,N_465,N_2987);
and U4735 (N_4735,N_2412,N_425);
and U4736 (N_4736,N_1800,N_1904);
nor U4737 (N_4737,N_183,N_2850);
nand U4738 (N_4738,N_1302,N_1732);
and U4739 (N_4739,N_757,N_2231);
and U4740 (N_4740,N_1255,N_2929);
nand U4741 (N_4741,N_2709,N_83);
or U4742 (N_4742,N_2209,N_1552);
nand U4743 (N_4743,N_1410,N_2283);
and U4744 (N_4744,N_1965,N_144);
nand U4745 (N_4745,N_2188,N_831);
and U4746 (N_4746,N_244,N_1165);
nor U4747 (N_4747,N_1559,N_2907);
nor U4748 (N_4748,N_1478,N_1766);
or U4749 (N_4749,N_2930,N_1457);
nor U4750 (N_4750,N_270,N_2980);
and U4751 (N_4751,N_1070,N_1226);
nor U4752 (N_4752,N_679,N_1558);
or U4753 (N_4753,N_67,N_282);
or U4754 (N_4754,N_2326,N_2355);
and U4755 (N_4755,N_2097,N_1458);
nor U4756 (N_4756,N_2389,N_2155);
nor U4757 (N_4757,N_2600,N_831);
nand U4758 (N_4758,N_255,N_561);
nand U4759 (N_4759,N_2898,N_762);
and U4760 (N_4760,N_1491,N_2998);
nand U4761 (N_4761,N_2586,N_1764);
xor U4762 (N_4762,N_610,N_1305);
nand U4763 (N_4763,N_1640,N_2865);
and U4764 (N_4764,N_420,N_2879);
nand U4765 (N_4765,N_1102,N_349);
and U4766 (N_4766,N_1812,N_1991);
or U4767 (N_4767,N_325,N_2142);
and U4768 (N_4768,N_291,N_2411);
nor U4769 (N_4769,N_2624,N_1396);
or U4770 (N_4770,N_1259,N_2013);
nor U4771 (N_4771,N_163,N_944);
nor U4772 (N_4772,N_389,N_2676);
or U4773 (N_4773,N_2959,N_102);
nand U4774 (N_4774,N_378,N_2657);
xnor U4775 (N_4775,N_2515,N_262);
nand U4776 (N_4776,N_1068,N_2411);
nand U4777 (N_4777,N_1093,N_1940);
nor U4778 (N_4778,N_129,N_1331);
nor U4779 (N_4779,N_2730,N_493);
or U4780 (N_4780,N_1845,N_1971);
nor U4781 (N_4781,N_183,N_1773);
nor U4782 (N_4782,N_1554,N_2124);
or U4783 (N_4783,N_441,N_1687);
nand U4784 (N_4784,N_2885,N_1282);
nand U4785 (N_4785,N_2564,N_1857);
nor U4786 (N_4786,N_1889,N_16);
nand U4787 (N_4787,N_774,N_1265);
and U4788 (N_4788,N_1933,N_2570);
xnor U4789 (N_4789,N_798,N_749);
nor U4790 (N_4790,N_1010,N_2646);
nand U4791 (N_4791,N_1246,N_2561);
or U4792 (N_4792,N_371,N_1438);
nand U4793 (N_4793,N_2341,N_1564);
nor U4794 (N_4794,N_1965,N_1122);
nor U4795 (N_4795,N_841,N_1942);
or U4796 (N_4796,N_248,N_2585);
or U4797 (N_4797,N_2261,N_273);
and U4798 (N_4798,N_2246,N_941);
and U4799 (N_4799,N_2939,N_2924);
or U4800 (N_4800,N_494,N_2364);
nand U4801 (N_4801,N_911,N_153);
nand U4802 (N_4802,N_1110,N_1559);
or U4803 (N_4803,N_1154,N_1936);
and U4804 (N_4804,N_945,N_406);
nand U4805 (N_4805,N_2431,N_2234);
or U4806 (N_4806,N_1970,N_2827);
and U4807 (N_4807,N_1122,N_2449);
nor U4808 (N_4808,N_1082,N_2044);
or U4809 (N_4809,N_2401,N_320);
nand U4810 (N_4810,N_959,N_1631);
and U4811 (N_4811,N_777,N_2982);
or U4812 (N_4812,N_212,N_2192);
nor U4813 (N_4813,N_2090,N_2248);
nand U4814 (N_4814,N_1067,N_730);
and U4815 (N_4815,N_2083,N_2923);
nand U4816 (N_4816,N_583,N_815);
nand U4817 (N_4817,N_1218,N_1217);
or U4818 (N_4818,N_1627,N_208);
xor U4819 (N_4819,N_2555,N_962);
or U4820 (N_4820,N_89,N_854);
nor U4821 (N_4821,N_2536,N_580);
or U4822 (N_4822,N_2033,N_353);
nor U4823 (N_4823,N_1506,N_2237);
or U4824 (N_4824,N_726,N_2148);
and U4825 (N_4825,N_173,N_621);
or U4826 (N_4826,N_2514,N_2303);
nand U4827 (N_4827,N_238,N_1170);
nor U4828 (N_4828,N_2782,N_1589);
and U4829 (N_4829,N_1007,N_530);
nand U4830 (N_4830,N_2380,N_2322);
xnor U4831 (N_4831,N_1681,N_2387);
or U4832 (N_4832,N_1473,N_2247);
and U4833 (N_4833,N_1467,N_453);
or U4834 (N_4834,N_2801,N_766);
nand U4835 (N_4835,N_347,N_1119);
nand U4836 (N_4836,N_1379,N_2481);
xor U4837 (N_4837,N_392,N_11);
nand U4838 (N_4838,N_287,N_176);
and U4839 (N_4839,N_459,N_1072);
nand U4840 (N_4840,N_651,N_862);
xor U4841 (N_4841,N_1971,N_226);
and U4842 (N_4842,N_2460,N_109);
or U4843 (N_4843,N_740,N_1474);
or U4844 (N_4844,N_1424,N_2363);
nor U4845 (N_4845,N_2773,N_1724);
and U4846 (N_4846,N_1440,N_164);
nand U4847 (N_4847,N_735,N_2749);
nor U4848 (N_4848,N_1328,N_723);
nor U4849 (N_4849,N_2507,N_1795);
nand U4850 (N_4850,N_1505,N_2426);
or U4851 (N_4851,N_975,N_2859);
nand U4852 (N_4852,N_2814,N_148);
and U4853 (N_4853,N_176,N_1280);
nor U4854 (N_4854,N_2216,N_2515);
and U4855 (N_4855,N_1415,N_968);
and U4856 (N_4856,N_563,N_67);
and U4857 (N_4857,N_31,N_946);
nand U4858 (N_4858,N_1123,N_638);
nand U4859 (N_4859,N_597,N_1334);
nand U4860 (N_4860,N_2347,N_2476);
or U4861 (N_4861,N_1887,N_1168);
and U4862 (N_4862,N_2390,N_2734);
nor U4863 (N_4863,N_1197,N_535);
and U4864 (N_4864,N_2329,N_624);
and U4865 (N_4865,N_1032,N_74);
or U4866 (N_4866,N_2998,N_647);
nand U4867 (N_4867,N_2644,N_2267);
and U4868 (N_4868,N_958,N_529);
or U4869 (N_4869,N_2382,N_2202);
nor U4870 (N_4870,N_1253,N_1457);
and U4871 (N_4871,N_2751,N_1696);
nand U4872 (N_4872,N_695,N_1677);
nand U4873 (N_4873,N_1674,N_2418);
nand U4874 (N_4874,N_745,N_2614);
nand U4875 (N_4875,N_2459,N_2369);
or U4876 (N_4876,N_33,N_2925);
xor U4877 (N_4877,N_1166,N_2726);
nand U4878 (N_4878,N_1215,N_917);
nand U4879 (N_4879,N_1804,N_909);
nor U4880 (N_4880,N_836,N_2750);
nand U4881 (N_4881,N_1470,N_1146);
and U4882 (N_4882,N_887,N_338);
nand U4883 (N_4883,N_1658,N_2826);
and U4884 (N_4884,N_2804,N_2107);
and U4885 (N_4885,N_2520,N_1398);
nand U4886 (N_4886,N_2176,N_464);
or U4887 (N_4887,N_989,N_1829);
or U4888 (N_4888,N_714,N_1468);
xor U4889 (N_4889,N_1813,N_111);
xnor U4890 (N_4890,N_1708,N_2209);
and U4891 (N_4891,N_1570,N_1593);
and U4892 (N_4892,N_1231,N_2089);
and U4893 (N_4893,N_514,N_1127);
nor U4894 (N_4894,N_2148,N_1647);
and U4895 (N_4895,N_1894,N_1619);
and U4896 (N_4896,N_1768,N_430);
nand U4897 (N_4897,N_219,N_181);
and U4898 (N_4898,N_1142,N_1995);
and U4899 (N_4899,N_569,N_2895);
and U4900 (N_4900,N_1183,N_1062);
nor U4901 (N_4901,N_1661,N_995);
and U4902 (N_4902,N_2794,N_1666);
and U4903 (N_4903,N_1647,N_1441);
and U4904 (N_4904,N_1433,N_860);
nand U4905 (N_4905,N_1488,N_2936);
and U4906 (N_4906,N_275,N_82);
nor U4907 (N_4907,N_2645,N_1417);
nand U4908 (N_4908,N_887,N_1734);
or U4909 (N_4909,N_2692,N_2970);
nand U4910 (N_4910,N_2674,N_758);
or U4911 (N_4911,N_690,N_2944);
nand U4912 (N_4912,N_2480,N_430);
or U4913 (N_4913,N_2345,N_360);
nand U4914 (N_4914,N_2440,N_2534);
nand U4915 (N_4915,N_2037,N_1015);
xor U4916 (N_4916,N_105,N_429);
nor U4917 (N_4917,N_2169,N_139);
or U4918 (N_4918,N_1633,N_1918);
and U4919 (N_4919,N_538,N_838);
nor U4920 (N_4920,N_2115,N_2791);
or U4921 (N_4921,N_1561,N_641);
nor U4922 (N_4922,N_2479,N_2321);
or U4923 (N_4923,N_1049,N_1587);
or U4924 (N_4924,N_295,N_2965);
nor U4925 (N_4925,N_1009,N_1788);
nand U4926 (N_4926,N_2226,N_1502);
and U4927 (N_4927,N_171,N_2287);
xnor U4928 (N_4928,N_232,N_591);
nand U4929 (N_4929,N_2148,N_1812);
and U4930 (N_4930,N_2634,N_2953);
and U4931 (N_4931,N_1159,N_1531);
nor U4932 (N_4932,N_1159,N_818);
or U4933 (N_4933,N_356,N_2213);
or U4934 (N_4934,N_1236,N_2577);
and U4935 (N_4935,N_1567,N_1054);
nor U4936 (N_4936,N_1068,N_688);
nand U4937 (N_4937,N_29,N_1751);
nand U4938 (N_4938,N_1091,N_40);
or U4939 (N_4939,N_1068,N_2975);
and U4940 (N_4940,N_1764,N_2725);
nand U4941 (N_4941,N_2412,N_1977);
or U4942 (N_4942,N_1808,N_2386);
nor U4943 (N_4943,N_600,N_513);
and U4944 (N_4944,N_2236,N_1697);
or U4945 (N_4945,N_1362,N_2265);
nor U4946 (N_4946,N_310,N_589);
nor U4947 (N_4947,N_2372,N_2573);
nor U4948 (N_4948,N_2900,N_832);
or U4949 (N_4949,N_733,N_849);
and U4950 (N_4950,N_2492,N_1055);
nor U4951 (N_4951,N_978,N_916);
nand U4952 (N_4952,N_185,N_968);
or U4953 (N_4953,N_2536,N_2753);
and U4954 (N_4954,N_259,N_2587);
and U4955 (N_4955,N_2091,N_1628);
and U4956 (N_4956,N_1450,N_1490);
and U4957 (N_4957,N_2431,N_1367);
or U4958 (N_4958,N_2996,N_689);
nor U4959 (N_4959,N_2276,N_2865);
nor U4960 (N_4960,N_2227,N_190);
or U4961 (N_4961,N_11,N_1911);
and U4962 (N_4962,N_43,N_1050);
or U4963 (N_4963,N_1372,N_1636);
and U4964 (N_4964,N_2759,N_416);
nand U4965 (N_4965,N_62,N_2647);
nor U4966 (N_4966,N_110,N_2699);
nor U4967 (N_4967,N_2508,N_1532);
nor U4968 (N_4968,N_1465,N_2172);
nor U4969 (N_4969,N_2386,N_1783);
nor U4970 (N_4970,N_520,N_2057);
nand U4971 (N_4971,N_1113,N_1538);
nand U4972 (N_4972,N_152,N_1135);
xnor U4973 (N_4973,N_1043,N_2508);
and U4974 (N_4974,N_946,N_125);
or U4975 (N_4975,N_2106,N_2447);
nand U4976 (N_4976,N_2293,N_1274);
nor U4977 (N_4977,N_276,N_2667);
or U4978 (N_4978,N_359,N_2190);
or U4979 (N_4979,N_1517,N_2739);
nand U4980 (N_4980,N_782,N_2087);
or U4981 (N_4981,N_1019,N_2550);
nor U4982 (N_4982,N_1909,N_2475);
nand U4983 (N_4983,N_2847,N_1397);
nor U4984 (N_4984,N_1713,N_839);
nand U4985 (N_4985,N_745,N_2910);
nor U4986 (N_4986,N_1760,N_1531);
or U4987 (N_4987,N_2957,N_390);
or U4988 (N_4988,N_2990,N_0);
nor U4989 (N_4989,N_69,N_268);
and U4990 (N_4990,N_2071,N_1003);
or U4991 (N_4991,N_2724,N_2366);
and U4992 (N_4992,N_2348,N_2625);
xnor U4993 (N_4993,N_1386,N_2408);
nand U4994 (N_4994,N_405,N_2314);
nor U4995 (N_4995,N_413,N_962);
nor U4996 (N_4996,N_2206,N_1579);
and U4997 (N_4997,N_2234,N_2133);
xor U4998 (N_4998,N_903,N_1103);
and U4999 (N_4999,N_2618,N_2038);
nor U5000 (N_5000,N_1537,N_452);
nand U5001 (N_5001,N_1009,N_2017);
and U5002 (N_5002,N_1561,N_584);
nor U5003 (N_5003,N_275,N_1289);
nand U5004 (N_5004,N_1870,N_732);
or U5005 (N_5005,N_2009,N_2176);
and U5006 (N_5006,N_1711,N_1845);
and U5007 (N_5007,N_2816,N_2304);
nand U5008 (N_5008,N_3,N_1100);
and U5009 (N_5009,N_2346,N_2954);
and U5010 (N_5010,N_1480,N_2895);
or U5011 (N_5011,N_38,N_1690);
nand U5012 (N_5012,N_749,N_865);
or U5013 (N_5013,N_2166,N_657);
nor U5014 (N_5014,N_688,N_1263);
or U5015 (N_5015,N_2427,N_178);
and U5016 (N_5016,N_612,N_1369);
or U5017 (N_5017,N_1415,N_1142);
nand U5018 (N_5018,N_2019,N_2488);
and U5019 (N_5019,N_225,N_2410);
nand U5020 (N_5020,N_2764,N_1542);
nand U5021 (N_5021,N_2606,N_1776);
nor U5022 (N_5022,N_2718,N_1087);
nand U5023 (N_5023,N_938,N_41);
nand U5024 (N_5024,N_86,N_2663);
nor U5025 (N_5025,N_2000,N_2604);
nor U5026 (N_5026,N_2712,N_660);
nor U5027 (N_5027,N_1623,N_2720);
nand U5028 (N_5028,N_928,N_987);
and U5029 (N_5029,N_2370,N_1171);
or U5030 (N_5030,N_492,N_2827);
and U5031 (N_5031,N_514,N_2956);
nor U5032 (N_5032,N_1034,N_1635);
and U5033 (N_5033,N_1270,N_1556);
nand U5034 (N_5034,N_2863,N_952);
nand U5035 (N_5035,N_2924,N_2121);
or U5036 (N_5036,N_374,N_1414);
nor U5037 (N_5037,N_1497,N_2685);
nor U5038 (N_5038,N_562,N_1661);
nor U5039 (N_5039,N_2689,N_1635);
nand U5040 (N_5040,N_304,N_923);
nand U5041 (N_5041,N_2905,N_2426);
nor U5042 (N_5042,N_281,N_893);
or U5043 (N_5043,N_325,N_427);
nor U5044 (N_5044,N_2409,N_458);
nor U5045 (N_5045,N_1491,N_1612);
and U5046 (N_5046,N_223,N_2705);
nand U5047 (N_5047,N_1458,N_85);
and U5048 (N_5048,N_127,N_1876);
nand U5049 (N_5049,N_491,N_1403);
or U5050 (N_5050,N_1275,N_832);
or U5051 (N_5051,N_1059,N_1169);
and U5052 (N_5052,N_871,N_1625);
or U5053 (N_5053,N_598,N_1916);
and U5054 (N_5054,N_2485,N_2027);
or U5055 (N_5055,N_1045,N_2438);
and U5056 (N_5056,N_444,N_240);
or U5057 (N_5057,N_888,N_1149);
nand U5058 (N_5058,N_2115,N_2605);
or U5059 (N_5059,N_2470,N_1506);
and U5060 (N_5060,N_2414,N_2798);
nor U5061 (N_5061,N_1694,N_2911);
nand U5062 (N_5062,N_1442,N_2653);
or U5063 (N_5063,N_2239,N_2870);
or U5064 (N_5064,N_2174,N_1199);
or U5065 (N_5065,N_2700,N_2878);
nand U5066 (N_5066,N_347,N_876);
and U5067 (N_5067,N_1883,N_723);
and U5068 (N_5068,N_1369,N_1483);
nand U5069 (N_5069,N_2812,N_2851);
or U5070 (N_5070,N_2582,N_511);
or U5071 (N_5071,N_2432,N_1646);
nand U5072 (N_5072,N_1847,N_1786);
nand U5073 (N_5073,N_2419,N_1904);
nor U5074 (N_5074,N_1317,N_913);
or U5075 (N_5075,N_2948,N_1917);
nor U5076 (N_5076,N_2077,N_1779);
nor U5077 (N_5077,N_1898,N_2033);
or U5078 (N_5078,N_445,N_1155);
nand U5079 (N_5079,N_2044,N_1562);
or U5080 (N_5080,N_2480,N_592);
and U5081 (N_5081,N_2383,N_674);
or U5082 (N_5082,N_710,N_365);
and U5083 (N_5083,N_2192,N_538);
nand U5084 (N_5084,N_1686,N_2370);
or U5085 (N_5085,N_1305,N_2556);
nand U5086 (N_5086,N_1213,N_2208);
or U5087 (N_5087,N_2031,N_2834);
or U5088 (N_5088,N_2482,N_2307);
nand U5089 (N_5089,N_1185,N_996);
and U5090 (N_5090,N_720,N_1160);
nand U5091 (N_5091,N_38,N_2887);
nand U5092 (N_5092,N_2410,N_1739);
and U5093 (N_5093,N_1164,N_1438);
and U5094 (N_5094,N_2626,N_1764);
xor U5095 (N_5095,N_1481,N_1310);
nand U5096 (N_5096,N_1959,N_2245);
nor U5097 (N_5097,N_367,N_1448);
and U5098 (N_5098,N_2251,N_2285);
and U5099 (N_5099,N_2159,N_1535);
and U5100 (N_5100,N_115,N_1592);
nor U5101 (N_5101,N_392,N_1397);
and U5102 (N_5102,N_2060,N_746);
nand U5103 (N_5103,N_2246,N_1759);
nand U5104 (N_5104,N_2958,N_2971);
nor U5105 (N_5105,N_1499,N_1637);
nand U5106 (N_5106,N_1647,N_1513);
nand U5107 (N_5107,N_729,N_871);
nand U5108 (N_5108,N_1570,N_1036);
or U5109 (N_5109,N_2071,N_1963);
and U5110 (N_5110,N_545,N_1262);
nand U5111 (N_5111,N_1829,N_2783);
nand U5112 (N_5112,N_1911,N_2309);
nor U5113 (N_5113,N_2471,N_1795);
nor U5114 (N_5114,N_2034,N_320);
nand U5115 (N_5115,N_2935,N_2706);
and U5116 (N_5116,N_2838,N_720);
xor U5117 (N_5117,N_1065,N_2046);
nor U5118 (N_5118,N_1304,N_778);
or U5119 (N_5119,N_2367,N_2388);
nand U5120 (N_5120,N_523,N_1489);
and U5121 (N_5121,N_2118,N_296);
nor U5122 (N_5122,N_1162,N_61);
xnor U5123 (N_5123,N_2013,N_2908);
nand U5124 (N_5124,N_261,N_1103);
nor U5125 (N_5125,N_2888,N_981);
nor U5126 (N_5126,N_2717,N_1122);
or U5127 (N_5127,N_458,N_1892);
and U5128 (N_5128,N_908,N_317);
nand U5129 (N_5129,N_2498,N_1080);
nor U5130 (N_5130,N_2411,N_1829);
nand U5131 (N_5131,N_2120,N_2481);
nand U5132 (N_5132,N_1030,N_1288);
and U5133 (N_5133,N_265,N_2721);
nor U5134 (N_5134,N_1293,N_1951);
or U5135 (N_5135,N_1520,N_2099);
or U5136 (N_5136,N_1196,N_2533);
and U5137 (N_5137,N_1250,N_2824);
or U5138 (N_5138,N_1153,N_414);
nand U5139 (N_5139,N_1432,N_2546);
or U5140 (N_5140,N_662,N_266);
or U5141 (N_5141,N_1502,N_1010);
and U5142 (N_5142,N_240,N_1987);
and U5143 (N_5143,N_1228,N_1387);
and U5144 (N_5144,N_1509,N_1333);
nand U5145 (N_5145,N_882,N_862);
and U5146 (N_5146,N_106,N_2604);
or U5147 (N_5147,N_1050,N_1834);
nand U5148 (N_5148,N_2867,N_2431);
and U5149 (N_5149,N_13,N_1576);
or U5150 (N_5150,N_1810,N_938);
or U5151 (N_5151,N_1936,N_1204);
nand U5152 (N_5152,N_1088,N_2697);
nor U5153 (N_5153,N_1377,N_1251);
or U5154 (N_5154,N_1774,N_1779);
nor U5155 (N_5155,N_1810,N_2525);
nor U5156 (N_5156,N_2879,N_2472);
xnor U5157 (N_5157,N_1251,N_2186);
nand U5158 (N_5158,N_960,N_1461);
nor U5159 (N_5159,N_691,N_1604);
nor U5160 (N_5160,N_2604,N_1414);
nor U5161 (N_5161,N_2440,N_1700);
and U5162 (N_5162,N_797,N_1169);
and U5163 (N_5163,N_2982,N_2909);
and U5164 (N_5164,N_2393,N_771);
nor U5165 (N_5165,N_2413,N_316);
nor U5166 (N_5166,N_2369,N_2141);
or U5167 (N_5167,N_1087,N_2201);
nor U5168 (N_5168,N_2700,N_1208);
nand U5169 (N_5169,N_2241,N_2773);
or U5170 (N_5170,N_992,N_2132);
and U5171 (N_5171,N_201,N_1796);
nand U5172 (N_5172,N_89,N_559);
or U5173 (N_5173,N_1530,N_1424);
nand U5174 (N_5174,N_922,N_115);
or U5175 (N_5175,N_1632,N_1848);
nor U5176 (N_5176,N_2412,N_271);
or U5177 (N_5177,N_227,N_1436);
or U5178 (N_5178,N_2955,N_305);
and U5179 (N_5179,N_1465,N_2599);
and U5180 (N_5180,N_528,N_1107);
nand U5181 (N_5181,N_789,N_153);
or U5182 (N_5182,N_1531,N_1873);
nand U5183 (N_5183,N_1824,N_2947);
nand U5184 (N_5184,N_2934,N_903);
or U5185 (N_5185,N_254,N_1163);
or U5186 (N_5186,N_1524,N_275);
nor U5187 (N_5187,N_1007,N_2221);
nand U5188 (N_5188,N_839,N_264);
nor U5189 (N_5189,N_45,N_2740);
nand U5190 (N_5190,N_1611,N_897);
nor U5191 (N_5191,N_644,N_1741);
and U5192 (N_5192,N_2525,N_2957);
or U5193 (N_5193,N_96,N_2732);
nor U5194 (N_5194,N_1683,N_2794);
nor U5195 (N_5195,N_1088,N_1235);
nor U5196 (N_5196,N_2763,N_152);
nor U5197 (N_5197,N_1698,N_2077);
or U5198 (N_5198,N_825,N_720);
or U5199 (N_5199,N_2966,N_965);
nand U5200 (N_5200,N_1658,N_2189);
xnor U5201 (N_5201,N_974,N_2827);
and U5202 (N_5202,N_844,N_390);
or U5203 (N_5203,N_772,N_2636);
nand U5204 (N_5204,N_641,N_2281);
or U5205 (N_5205,N_742,N_902);
nand U5206 (N_5206,N_2894,N_980);
xor U5207 (N_5207,N_1621,N_1878);
nor U5208 (N_5208,N_119,N_446);
and U5209 (N_5209,N_2518,N_2576);
nand U5210 (N_5210,N_2074,N_2932);
nor U5211 (N_5211,N_678,N_1721);
or U5212 (N_5212,N_705,N_1856);
nor U5213 (N_5213,N_1570,N_398);
and U5214 (N_5214,N_2819,N_396);
and U5215 (N_5215,N_2684,N_2439);
nor U5216 (N_5216,N_2251,N_847);
nor U5217 (N_5217,N_1341,N_1161);
and U5218 (N_5218,N_2139,N_1748);
or U5219 (N_5219,N_296,N_2074);
or U5220 (N_5220,N_1457,N_152);
nand U5221 (N_5221,N_993,N_1844);
and U5222 (N_5222,N_790,N_2073);
and U5223 (N_5223,N_1209,N_584);
and U5224 (N_5224,N_2989,N_1829);
and U5225 (N_5225,N_2620,N_2917);
and U5226 (N_5226,N_1129,N_3);
nand U5227 (N_5227,N_2997,N_476);
nor U5228 (N_5228,N_432,N_511);
nand U5229 (N_5229,N_2202,N_2330);
and U5230 (N_5230,N_1943,N_25);
or U5231 (N_5231,N_2322,N_1878);
nand U5232 (N_5232,N_1638,N_2453);
nand U5233 (N_5233,N_558,N_1139);
and U5234 (N_5234,N_1679,N_2325);
nor U5235 (N_5235,N_1505,N_154);
and U5236 (N_5236,N_79,N_2217);
nand U5237 (N_5237,N_1807,N_1482);
nand U5238 (N_5238,N_2037,N_2431);
or U5239 (N_5239,N_735,N_2430);
and U5240 (N_5240,N_2161,N_1008);
nor U5241 (N_5241,N_2293,N_619);
nand U5242 (N_5242,N_662,N_1334);
or U5243 (N_5243,N_2437,N_1773);
and U5244 (N_5244,N_713,N_2987);
nor U5245 (N_5245,N_372,N_175);
or U5246 (N_5246,N_88,N_2983);
nand U5247 (N_5247,N_971,N_2671);
or U5248 (N_5248,N_688,N_513);
or U5249 (N_5249,N_2999,N_625);
or U5250 (N_5250,N_484,N_2702);
and U5251 (N_5251,N_1390,N_1336);
nand U5252 (N_5252,N_1690,N_1050);
xor U5253 (N_5253,N_247,N_658);
and U5254 (N_5254,N_920,N_1567);
or U5255 (N_5255,N_2410,N_349);
or U5256 (N_5256,N_2061,N_389);
or U5257 (N_5257,N_2521,N_2357);
and U5258 (N_5258,N_2626,N_2226);
or U5259 (N_5259,N_22,N_1825);
nand U5260 (N_5260,N_2461,N_1524);
nor U5261 (N_5261,N_663,N_566);
nor U5262 (N_5262,N_1179,N_2060);
and U5263 (N_5263,N_1913,N_243);
or U5264 (N_5264,N_1902,N_713);
and U5265 (N_5265,N_556,N_2159);
xnor U5266 (N_5266,N_2493,N_2116);
nand U5267 (N_5267,N_900,N_521);
nor U5268 (N_5268,N_1284,N_2171);
nor U5269 (N_5269,N_2987,N_1092);
or U5270 (N_5270,N_2853,N_1364);
or U5271 (N_5271,N_1697,N_1621);
and U5272 (N_5272,N_1552,N_235);
or U5273 (N_5273,N_1557,N_1694);
nand U5274 (N_5274,N_2269,N_2647);
and U5275 (N_5275,N_2249,N_2843);
and U5276 (N_5276,N_762,N_1310);
and U5277 (N_5277,N_2317,N_1403);
or U5278 (N_5278,N_2698,N_2085);
nor U5279 (N_5279,N_1580,N_616);
and U5280 (N_5280,N_2873,N_1998);
and U5281 (N_5281,N_2048,N_1116);
nor U5282 (N_5282,N_217,N_480);
or U5283 (N_5283,N_610,N_296);
and U5284 (N_5284,N_1131,N_2519);
nor U5285 (N_5285,N_185,N_1971);
nand U5286 (N_5286,N_1157,N_257);
or U5287 (N_5287,N_547,N_1187);
nand U5288 (N_5288,N_425,N_2263);
nand U5289 (N_5289,N_1106,N_1647);
and U5290 (N_5290,N_2823,N_735);
or U5291 (N_5291,N_732,N_2029);
nor U5292 (N_5292,N_2357,N_605);
and U5293 (N_5293,N_2872,N_864);
or U5294 (N_5294,N_549,N_1995);
or U5295 (N_5295,N_857,N_533);
and U5296 (N_5296,N_366,N_354);
or U5297 (N_5297,N_1961,N_2602);
and U5298 (N_5298,N_726,N_2821);
and U5299 (N_5299,N_1578,N_224);
or U5300 (N_5300,N_189,N_645);
nor U5301 (N_5301,N_365,N_1842);
nand U5302 (N_5302,N_902,N_2228);
or U5303 (N_5303,N_119,N_1914);
nor U5304 (N_5304,N_1437,N_2947);
and U5305 (N_5305,N_2745,N_2811);
or U5306 (N_5306,N_2250,N_2191);
or U5307 (N_5307,N_1643,N_1182);
nor U5308 (N_5308,N_2850,N_237);
nand U5309 (N_5309,N_2229,N_1814);
nand U5310 (N_5310,N_2858,N_617);
nand U5311 (N_5311,N_59,N_2125);
and U5312 (N_5312,N_2593,N_924);
and U5313 (N_5313,N_2741,N_2521);
and U5314 (N_5314,N_2058,N_1929);
nand U5315 (N_5315,N_805,N_2505);
or U5316 (N_5316,N_504,N_1843);
and U5317 (N_5317,N_521,N_1221);
nand U5318 (N_5318,N_1863,N_522);
or U5319 (N_5319,N_540,N_1447);
or U5320 (N_5320,N_1807,N_278);
nand U5321 (N_5321,N_1214,N_2595);
nor U5322 (N_5322,N_2458,N_2477);
nand U5323 (N_5323,N_2656,N_2437);
nand U5324 (N_5324,N_142,N_1069);
nor U5325 (N_5325,N_955,N_52);
nor U5326 (N_5326,N_1809,N_170);
and U5327 (N_5327,N_1991,N_2204);
nor U5328 (N_5328,N_1448,N_1213);
nor U5329 (N_5329,N_1046,N_1149);
and U5330 (N_5330,N_1809,N_2204);
or U5331 (N_5331,N_417,N_1866);
or U5332 (N_5332,N_2941,N_2461);
or U5333 (N_5333,N_2614,N_1433);
or U5334 (N_5334,N_2934,N_2611);
nand U5335 (N_5335,N_601,N_1141);
nand U5336 (N_5336,N_2872,N_2881);
nor U5337 (N_5337,N_949,N_1677);
and U5338 (N_5338,N_294,N_55);
or U5339 (N_5339,N_1734,N_2788);
or U5340 (N_5340,N_2608,N_2153);
and U5341 (N_5341,N_893,N_697);
nor U5342 (N_5342,N_1534,N_242);
nor U5343 (N_5343,N_1297,N_497);
nand U5344 (N_5344,N_2870,N_2307);
nor U5345 (N_5345,N_1928,N_2509);
or U5346 (N_5346,N_2945,N_1255);
nand U5347 (N_5347,N_2167,N_1239);
nand U5348 (N_5348,N_1751,N_1349);
or U5349 (N_5349,N_419,N_1913);
and U5350 (N_5350,N_2199,N_1208);
nor U5351 (N_5351,N_1267,N_2454);
or U5352 (N_5352,N_2955,N_2177);
xnor U5353 (N_5353,N_1262,N_1290);
or U5354 (N_5354,N_2293,N_1355);
nand U5355 (N_5355,N_2728,N_201);
and U5356 (N_5356,N_635,N_167);
nor U5357 (N_5357,N_2765,N_383);
xnor U5358 (N_5358,N_1092,N_798);
and U5359 (N_5359,N_238,N_785);
nand U5360 (N_5360,N_1944,N_950);
or U5361 (N_5361,N_1855,N_148);
nor U5362 (N_5362,N_558,N_2506);
or U5363 (N_5363,N_707,N_2024);
and U5364 (N_5364,N_1769,N_2669);
and U5365 (N_5365,N_2981,N_2265);
nand U5366 (N_5366,N_1949,N_2514);
or U5367 (N_5367,N_217,N_2890);
nor U5368 (N_5368,N_373,N_711);
and U5369 (N_5369,N_830,N_1740);
xor U5370 (N_5370,N_2949,N_2448);
or U5371 (N_5371,N_1645,N_2499);
nand U5372 (N_5372,N_1067,N_1843);
nand U5373 (N_5373,N_1091,N_2302);
or U5374 (N_5374,N_14,N_2628);
nor U5375 (N_5375,N_2254,N_561);
or U5376 (N_5376,N_2601,N_210);
or U5377 (N_5377,N_279,N_2778);
or U5378 (N_5378,N_1805,N_1597);
or U5379 (N_5379,N_1727,N_1960);
nand U5380 (N_5380,N_763,N_1616);
or U5381 (N_5381,N_1264,N_596);
xor U5382 (N_5382,N_2441,N_98);
nand U5383 (N_5383,N_1328,N_1174);
xnor U5384 (N_5384,N_192,N_2766);
nor U5385 (N_5385,N_1531,N_1107);
nor U5386 (N_5386,N_313,N_275);
nor U5387 (N_5387,N_1348,N_1407);
or U5388 (N_5388,N_28,N_615);
and U5389 (N_5389,N_2011,N_19);
and U5390 (N_5390,N_2432,N_940);
and U5391 (N_5391,N_2573,N_2795);
nor U5392 (N_5392,N_2578,N_796);
and U5393 (N_5393,N_558,N_1570);
nand U5394 (N_5394,N_626,N_303);
and U5395 (N_5395,N_349,N_2121);
or U5396 (N_5396,N_573,N_2249);
nand U5397 (N_5397,N_764,N_1013);
and U5398 (N_5398,N_1972,N_2577);
nand U5399 (N_5399,N_2738,N_76);
or U5400 (N_5400,N_1381,N_1223);
nor U5401 (N_5401,N_562,N_2955);
and U5402 (N_5402,N_1416,N_2547);
or U5403 (N_5403,N_2901,N_1211);
and U5404 (N_5404,N_1149,N_2599);
and U5405 (N_5405,N_2146,N_808);
or U5406 (N_5406,N_1479,N_2997);
nor U5407 (N_5407,N_509,N_1682);
nor U5408 (N_5408,N_2134,N_941);
nand U5409 (N_5409,N_2024,N_2433);
nand U5410 (N_5410,N_1766,N_1721);
nor U5411 (N_5411,N_174,N_893);
and U5412 (N_5412,N_1495,N_1680);
nor U5413 (N_5413,N_2943,N_2665);
or U5414 (N_5414,N_1828,N_2304);
and U5415 (N_5415,N_2603,N_1702);
and U5416 (N_5416,N_294,N_2624);
nor U5417 (N_5417,N_2684,N_2073);
or U5418 (N_5418,N_2013,N_2063);
nand U5419 (N_5419,N_2671,N_1908);
nor U5420 (N_5420,N_2498,N_1526);
and U5421 (N_5421,N_1409,N_544);
or U5422 (N_5422,N_1497,N_231);
nand U5423 (N_5423,N_933,N_433);
nand U5424 (N_5424,N_911,N_2485);
or U5425 (N_5425,N_2393,N_105);
nor U5426 (N_5426,N_1212,N_2661);
nor U5427 (N_5427,N_2836,N_218);
or U5428 (N_5428,N_2017,N_273);
or U5429 (N_5429,N_2768,N_2907);
nor U5430 (N_5430,N_1671,N_2024);
nor U5431 (N_5431,N_1914,N_1977);
and U5432 (N_5432,N_567,N_494);
nand U5433 (N_5433,N_697,N_2457);
or U5434 (N_5434,N_2698,N_852);
and U5435 (N_5435,N_1234,N_1023);
or U5436 (N_5436,N_67,N_263);
nor U5437 (N_5437,N_1326,N_2762);
and U5438 (N_5438,N_2698,N_864);
nor U5439 (N_5439,N_1208,N_1692);
nand U5440 (N_5440,N_2128,N_1874);
and U5441 (N_5441,N_1576,N_2540);
or U5442 (N_5442,N_431,N_873);
and U5443 (N_5443,N_2033,N_2942);
nand U5444 (N_5444,N_1672,N_2094);
and U5445 (N_5445,N_78,N_978);
nand U5446 (N_5446,N_432,N_298);
nand U5447 (N_5447,N_132,N_1890);
or U5448 (N_5448,N_2050,N_2237);
or U5449 (N_5449,N_2273,N_403);
nor U5450 (N_5450,N_1251,N_2076);
or U5451 (N_5451,N_1366,N_153);
nor U5452 (N_5452,N_1824,N_1895);
nor U5453 (N_5453,N_1069,N_1801);
and U5454 (N_5454,N_2677,N_1853);
nor U5455 (N_5455,N_988,N_1227);
or U5456 (N_5456,N_1343,N_1743);
nand U5457 (N_5457,N_2151,N_1516);
and U5458 (N_5458,N_1159,N_1173);
and U5459 (N_5459,N_2721,N_1155);
nor U5460 (N_5460,N_2579,N_2242);
or U5461 (N_5461,N_2310,N_956);
xnor U5462 (N_5462,N_18,N_2874);
and U5463 (N_5463,N_1763,N_34);
nor U5464 (N_5464,N_1692,N_116);
nand U5465 (N_5465,N_139,N_1045);
or U5466 (N_5466,N_2437,N_769);
nand U5467 (N_5467,N_554,N_1718);
or U5468 (N_5468,N_377,N_613);
xor U5469 (N_5469,N_1471,N_1505);
or U5470 (N_5470,N_1834,N_2239);
nor U5471 (N_5471,N_2234,N_1496);
or U5472 (N_5472,N_134,N_2083);
nor U5473 (N_5473,N_599,N_2204);
nor U5474 (N_5474,N_206,N_1025);
nor U5475 (N_5475,N_1676,N_2591);
or U5476 (N_5476,N_1808,N_330);
nor U5477 (N_5477,N_1056,N_2079);
or U5478 (N_5478,N_1960,N_1094);
nand U5479 (N_5479,N_2603,N_2647);
and U5480 (N_5480,N_1728,N_2080);
nor U5481 (N_5481,N_2752,N_1210);
and U5482 (N_5482,N_1470,N_872);
and U5483 (N_5483,N_1601,N_1134);
nor U5484 (N_5484,N_716,N_1025);
nor U5485 (N_5485,N_900,N_64);
nor U5486 (N_5486,N_310,N_1207);
and U5487 (N_5487,N_2955,N_820);
or U5488 (N_5488,N_292,N_1702);
or U5489 (N_5489,N_2629,N_1051);
nor U5490 (N_5490,N_1223,N_859);
nor U5491 (N_5491,N_1814,N_1738);
nor U5492 (N_5492,N_457,N_372);
and U5493 (N_5493,N_395,N_2576);
nand U5494 (N_5494,N_2972,N_2024);
nand U5495 (N_5495,N_620,N_2737);
nand U5496 (N_5496,N_2531,N_342);
and U5497 (N_5497,N_2571,N_2982);
and U5498 (N_5498,N_2243,N_288);
or U5499 (N_5499,N_987,N_1987);
and U5500 (N_5500,N_1645,N_891);
nand U5501 (N_5501,N_1443,N_2239);
nand U5502 (N_5502,N_48,N_1737);
or U5503 (N_5503,N_1116,N_2925);
nor U5504 (N_5504,N_2317,N_928);
xor U5505 (N_5505,N_2895,N_417);
nor U5506 (N_5506,N_2789,N_1124);
nor U5507 (N_5507,N_2469,N_569);
nand U5508 (N_5508,N_1301,N_2416);
and U5509 (N_5509,N_2940,N_239);
nand U5510 (N_5510,N_1126,N_541);
and U5511 (N_5511,N_1530,N_670);
and U5512 (N_5512,N_1250,N_2947);
nand U5513 (N_5513,N_2447,N_1241);
and U5514 (N_5514,N_650,N_732);
or U5515 (N_5515,N_1095,N_763);
or U5516 (N_5516,N_2685,N_1655);
nor U5517 (N_5517,N_342,N_2392);
nor U5518 (N_5518,N_394,N_1385);
and U5519 (N_5519,N_408,N_1967);
nand U5520 (N_5520,N_634,N_520);
and U5521 (N_5521,N_1058,N_429);
xor U5522 (N_5522,N_26,N_1234);
and U5523 (N_5523,N_2089,N_493);
or U5524 (N_5524,N_48,N_1965);
or U5525 (N_5525,N_59,N_2608);
or U5526 (N_5526,N_1094,N_1765);
or U5527 (N_5527,N_5,N_2855);
nand U5528 (N_5528,N_517,N_1459);
nor U5529 (N_5529,N_1859,N_1130);
or U5530 (N_5530,N_2732,N_183);
nor U5531 (N_5531,N_1377,N_503);
and U5532 (N_5532,N_66,N_193);
and U5533 (N_5533,N_2354,N_523);
and U5534 (N_5534,N_2020,N_1148);
and U5535 (N_5535,N_51,N_940);
nand U5536 (N_5536,N_1777,N_1739);
nand U5537 (N_5537,N_209,N_1989);
or U5538 (N_5538,N_405,N_1500);
xor U5539 (N_5539,N_1510,N_1287);
and U5540 (N_5540,N_266,N_136);
or U5541 (N_5541,N_1850,N_1307);
and U5542 (N_5542,N_324,N_453);
and U5543 (N_5543,N_2536,N_1113);
nand U5544 (N_5544,N_906,N_1791);
and U5545 (N_5545,N_2719,N_572);
and U5546 (N_5546,N_2407,N_283);
and U5547 (N_5547,N_2045,N_2817);
nor U5548 (N_5548,N_1686,N_1108);
nor U5549 (N_5549,N_1694,N_2733);
nor U5550 (N_5550,N_2986,N_296);
nand U5551 (N_5551,N_2949,N_1633);
or U5552 (N_5552,N_1347,N_1861);
and U5553 (N_5553,N_1838,N_986);
nand U5554 (N_5554,N_1491,N_2145);
nor U5555 (N_5555,N_1413,N_2247);
nor U5556 (N_5556,N_1537,N_1977);
nand U5557 (N_5557,N_1084,N_3);
nor U5558 (N_5558,N_44,N_2637);
nand U5559 (N_5559,N_2434,N_348);
nand U5560 (N_5560,N_2141,N_1447);
nand U5561 (N_5561,N_33,N_2295);
and U5562 (N_5562,N_854,N_2413);
nor U5563 (N_5563,N_2181,N_1847);
and U5564 (N_5564,N_1549,N_2834);
nand U5565 (N_5565,N_2629,N_2758);
or U5566 (N_5566,N_1591,N_420);
nor U5567 (N_5567,N_1155,N_1902);
and U5568 (N_5568,N_515,N_615);
or U5569 (N_5569,N_823,N_660);
nor U5570 (N_5570,N_2037,N_1393);
or U5571 (N_5571,N_2821,N_1545);
or U5572 (N_5572,N_1054,N_151);
and U5573 (N_5573,N_1463,N_189);
nand U5574 (N_5574,N_136,N_2362);
or U5575 (N_5575,N_127,N_889);
nor U5576 (N_5576,N_2720,N_2129);
nand U5577 (N_5577,N_1233,N_2711);
or U5578 (N_5578,N_2994,N_2904);
nand U5579 (N_5579,N_985,N_897);
or U5580 (N_5580,N_362,N_1844);
nor U5581 (N_5581,N_838,N_863);
or U5582 (N_5582,N_2714,N_317);
or U5583 (N_5583,N_319,N_213);
nor U5584 (N_5584,N_1677,N_1259);
nand U5585 (N_5585,N_2588,N_2402);
and U5586 (N_5586,N_1730,N_2209);
or U5587 (N_5587,N_2705,N_622);
xor U5588 (N_5588,N_2342,N_1301);
and U5589 (N_5589,N_1533,N_77);
nand U5590 (N_5590,N_808,N_2503);
or U5591 (N_5591,N_916,N_1869);
nor U5592 (N_5592,N_342,N_1992);
and U5593 (N_5593,N_586,N_233);
or U5594 (N_5594,N_2033,N_1394);
nand U5595 (N_5595,N_2281,N_2679);
nor U5596 (N_5596,N_1489,N_1924);
nor U5597 (N_5597,N_2442,N_2973);
nand U5598 (N_5598,N_2213,N_837);
nand U5599 (N_5599,N_563,N_939);
and U5600 (N_5600,N_2253,N_1570);
nor U5601 (N_5601,N_2222,N_1044);
or U5602 (N_5602,N_2134,N_1848);
nor U5603 (N_5603,N_2799,N_81);
nor U5604 (N_5604,N_706,N_2389);
or U5605 (N_5605,N_1003,N_692);
or U5606 (N_5606,N_581,N_1831);
and U5607 (N_5607,N_300,N_671);
nor U5608 (N_5608,N_1591,N_967);
or U5609 (N_5609,N_2142,N_176);
and U5610 (N_5610,N_2056,N_2878);
nand U5611 (N_5611,N_925,N_1811);
nor U5612 (N_5612,N_157,N_1326);
nand U5613 (N_5613,N_1887,N_1175);
and U5614 (N_5614,N_495,N_2794);
or U5615 (N_5615,N_2735,N_2828);
or U5616 (N_5616,N_1755,N_2433);
nor U5617 (N_5617,N_1125,N_324);
and U5618 (N_5618,N_146,N_2248);
nor U5619 (N_5619,N_801,N_1096);
or U5620 (N_5620,N_1835,N_1213);
or U5621 (N_5621,N_863,N_1954);
or U5622 (N_5622,N_1747,N_467);
nor U5623 (N_5623,N_2973,N_2321);
nand U5624 (N_5624,N_2314,N_2278);
nand U5625 (N_5625,N_2663,N_2118);
and U5626 (N_5626,N_2467,N_1903);
nor U5627 (N_5627,N_286,N_27);
and U5628 (N_5628,N_1021,N_600);
nor U5629 (N_5629,N_141,N_455);
or U5630 (N_5630,N_2856,N_793);
xor U5631 (N_5631,N_1769,N_1614);
nand U5632 (N_5632,N_2531,N_56);
nand U5633 (N_5633,N_2383,N_909);
nand U5634 (N_5634,N_1563,N_756);
nand U5635 (N_5635,N_1423,N_1108);
nand U5636 (N_5636,N_2048,N_2877);
or U5637 (N_5637,N_1413,N_2740);
nand U5638 (N_5638,N_514,N_2199);
and U5639 (N_5639,N_1795,N_1003);
nor U5640 (N_5640,N_2194,N_216);
or U5641 (N_5641,N_1099,N_2575);
nand U5642 (N_5642,N_506,N_1208);
and U5643 (N_5643,N_2234,N_430);
and U5644 (N_5644,N_399,N_1273);
and U5645 (N_5645,N_946,N_776);
and U5646 (N_5646,N_1092,N_2967);
or U5647 (N_5647,N_2196,N_121);
nor U5648 (N_5648,N_886,N_1877);
nor U5649 (N_5649,N_1092,N_2850);
nand U5650 (N_5650,N_1601,N_698);
or U5651 (N_5651,N_1557,N_2216);
nor U5652 (N_5652,N_2058,N_1081);
nor U5653 (N_5653,N_9,N_282);
or U5654 (N_5654,N_1504,N_153);
or U5655 (N_5655,N_1940,N_902);
and U5656 (N_5656,N_633,N_340);
nor U5657 (N_5657,N_1287,N_17);
nand U5658 (N_5658,N_2464,N_308);
and U5659 (N_5659,N_1611,N_2641);
nor U5660 (N_5660,N_1169,N_55);
nor U5661 (N_5661,N_790,N_2685);
and U5662 (N_5662,N_2078,N_2677);
or U5663 (N_5663,N_338,N_370);
nand U5664 (N_5664,N_1606,N_1794);
nand U5665 (N_5665,N_2009,N_2624);
xor U5666 (N_5666,N_1482,N_1651);
nor U5667 (N_5667,N_1278,N_783);
nand U5668 (N_5668,N_1516,N_1187);
nand U5669 (N_5669,N_12,N_470);
and U5670 (N_5670,N_450,N_2373);
or U5671 (N_5671,N_25,N_2617);
or U5672 (N_5672,N_2398,N_818);
or U5673 (N_5673,N_2358,N_643);
or U5674 (N_5674,N_2927,N_346);
nor U5675 (N_5675,N_671,N_456);
and U5676 (N_5676,N_2175,N_1577);
or U5677 (N_5677,N_956,N_1922);
and U5678 (N_5678,N_2408,N_1523);
nor U5679 (N_5679,N_1586,N_1601);
nand U5680 (N_5680,N_1359,N_768);
nand U5681 (N_5681,N_2789,N_1335);
or U5682 (N_5682,N_2240,N_249);
nor U5683 (N_5683,N_555,N_2134);
nand U5684 (N_5684,N_1104,N_919);
nand U5685 (N_5685,N_1006,N_1899);
nand U5686 (N_5686,N_1274,N_2246);
nand U5687 (N_5687,N_673,N_1825);
nand U5688 (N_5688,N_24,N_735);
nor U5689 (N_5689,N_1788,N_2580);
nand U5690 (N_5690,N_864,N_2514);
and U5691 (N_5691,N_1759,N_2925);
nand U5692 (N_5692,N_101,N_147);
and U5693 (N_5693,N_2612,N_2135);
nand U5694 (N_5694,N_392,N_1727);
and U5695 (N_5695,N_2156,N_791);
nand U5696 (N_5696,N_2975,N_1226);
nor U5697 (N_5697,N_285,N_2792);
or U5698 (N_5698,N_254,N_375);
and U5699 (N_5699,N_196,N_942);
nor U5700 (N_5700,N_1211,N_2578);
nor U5701 (N_5701,N_474,N_2594);
nor U5702 (N_5702,N_1632,N_1322);
nand U5703 (N_5703,N_1363,N_379);
nand U5704 (N_5704,N_1332,N_382);
and U5705 (N_5705,N_487,N_514);
and U5706 (N_5706,N_2645,N_2512);
and U5707 (N_5707,N_2328,N_1407);
or U5708 (N_5708,N_986,N_2595);
and U5709 (N_5709,N_2212,N_2344);
xnor U5710 (N_5710,N_414,N_2594);
nand U5711 (N_5711,N_2555,N_1743);
and U5712 (N_5712,N_1740,N_2157);
or U5713 (N_5713,N_494,N_468);
and U5714 (N_5714,N_2357,N_2837);
xnor U5715 (N_5715,N_1382,N_532);
or U5716 (N_5716,N_2255,N_2432);
and U5717 (N_5717,N_418,N_2050);
or U5718 (N_5718,N_1664,N_2268);
or U5719 (N_5719,N_2496,N_775);
or U5720 (N_5720,N_327,N_2369);
and U5721 (N_5721,N_2361,N_858);
and U5722 (N_5722,N_467,N_1870);
nand U5723 (N_5723,N_807,N_2913);
nor U5724 (N_5724,N_2925,N_1826);
nor U5725 (N_5725,N_503,N_2310);
nor U5726 (N_5726,N_293,N_124);
nor U5727 (N_5727,N_2619,N_2922);
and U5728 (N_5728,N_2621,N_2135);
or U5729 (N_5729,N_352,N_2031);
or U5730 (N_5730,N_833,N_288);
and U5731 (N_5731,N_2456,N_1184);
or U5732 (N_5732,N_287,N_2934);
or U5733 (N_5733,N_2823,N_104);
or U5734 (N_5734,N_1827,N_418);
or U5735 (N_5735,N_815,N_1091);
nor U5736 (N_5736,N_125,N_1076);
nand U5737 (N_5737,N_1228,N_2694);
nand U5738 (N_5738,N_331,N_1938);
and U5739 (N_5739,N_315,N_426);
or U5740 (N_5740,N_1429,N_502);
and U5741 (N_5741,N_572,N_1138);
nand U5742 (N_5742,N_2864,N_1209);
nand U5743 (N_5743,N_1878,N_1719);
nor U5744 (N_5744,N_2490,N_2815);
nor U5745 (N_5745,N_574,N_1066);
nand U5746 (N_5746,N_552,N_1823);
nor U5747 (N_5747,N_772,N_2297);
nand U5748 (N_5748,N_626,N_1172);
xnor U5749 (N_5749,N_632,N_1154);
nor U5750 (N_5750,N_2177,N_1615);
and U5751 (N_5751,N_1392,N_2875);
or U5752 (N_5752,N_1727,N_1839);
nor U5753 (N_5753,N_2185,N_1353);
nor U5754 (N_5754,N_2039,N_578);
nor U5755 (N_5755,N_2703,N_2734);
and U5756 (N_5756,N_1360,N_1396);
or U5757 (N_5757,N_1872,N_1346);
and U5758 (N_5758,N_2334,N_2430);
and U5759 (N_5759,N_31,N_2756);
and U5760 (N_5760,N_152,N_2833);
nor U5761 (N_5761,N_1029,N_2014);
nand U5762 (N_5762,N_777,N_2546);
nand U5763 (N_5763,N_2803,N_1902);
and U5764 (N_5764,N_998,N_1064);
nor U5765 (N_5765,N_2264,N_2114);
and U5766 (N_5766,N_1469,N_297);
nor U5767 (N_5767,N_1630,N_1440);
or U5768 (N_5768,N_2514,N_1702);
and U5769 (N_5769,N_2330,N_2030);
and U5770 (N_5770,N_883,N_2130);
nand U5771 (N_5771,N_769,N_669);
and U5772 (N_5772,N_1556,N_743);
nor U5773 (N_5773,N_2339,N_45);
nor U5774 (N_5774,N_1557,N_536);
or U5775 (N_5775,N_2041,N_2186);
nor U5776 (N_5776,N_2503,N_938);
or U5777 (N_5777,N_2983,N_2923);
nor U5778 (N_5778,N_1941,N_348);
nor U5779 (N_5779,N_2715,N_344);
nor U5780 (N_5780,N_502,N_959);
nor U5781 (N_5781,N_1222,N_2028);
and U5782 (N_5782,N_1374,N_415);
or U5783 (N_5783,N_942,N_2713);
nand U5784 (N_5784,N_2150,N_1789);
nand U5785 (N_5785,N_2296,N_2558);
xor U5786 (N_5786,N_1802,N_1645);
nand U5787 (N_5787,N_1951,N_77);
nor U5788 (N_5788,N_1758,N_2074);
nand U5789 (N_5789,N_2154,N_2435);
nand U5790 (N_5790,N_2080,N_2399);
and U5791 (N_5791,N_1838,N_175);
or U5792 (N_5792,N_2216,N_445);
or U5793 (N_5793,N_1749,N_1745);
and U5794 (N_5794,N_929,N_2439);
or U5795 (N_5795,N_282,N_246);
nand U5796 (N_5796,N_2359,N_2646);
nor U5797 (N_5797,N_1230,N_1980);
or U5798 (N_5798,N_1005,N_770);
nand U5799 (N_5799,N_2074,N_1331);
and U5800 (N_5800,N_1402,N_2088);
nand U5801 (N_5801,N_2373,N_1234);
xor U5802 (N_5802,N_1242,N_2838);
nor U5803 (N_5803,N_125,N_780);
nor U5804 (N_5804,N_2212,N_349);
and U5805 (N_5805,N_888,N_96);
and U5806 (N_5806,N_2129,N_678);
nand U5807 (N_5807,N_2007,N_515);
nor U5808 (N_5808,N_918,N_2928);
nor U5809 (N_5809,N_848,N_2266);
nand U5810 (N_5810,N_86,N_1207);
nand U5811 (N_5811,N_2262,N_1921);
nand U5812 (N_5812,N_2113,N_1745);
nand U5813 (N_5813,N_1746,N_794);
or U5814 (N_5814,N_971,N_2461);
and U5815 (N_5815,N_2076,N_2558);
xnor U5816 (N_5816,N_917,N_1331);
and U5817 (N_5817,N_1459,N_2045);
nor U5818 (N_5818,N_2968,N_2693);
or U5819 (N_5819,N_1672,N_449);
or U5820 (N_5820,N_367,N_2227);
nand U5821 (N_5821,N_2945,N_2832);
or U5822 (N_5822,N_2520,N_1276);
or U5823 (N_5823,N_35,N_198);
nor U5824 (N_5824,N_2935,N_2400);
and U5825 (N_5825,N_1113,N_36);
or U5826 (N_5826,N_1270,N_1474);
nand U5827 (N_5827,N_2422,N_374);
and U5828 (N_5828,N_715,N_816);
nand U5829 (N_5829,N_579,N_1961);
or U5830 (N_5830,N_1834,N_1426);
or U5831 (N_5831,N_707,N_2613);
or U5832 (N_5832,N_2947,N_1866);
and U5833 (N_5833,N_1775,N_1479);
or U5834 (N_5834,N_2453,N_1390);
or U5835 (N_5835,N_1914,N_1311);
and U5836 (N_5836,N_140,N_2728);
and U5837 (N_5837,N_438,N_1978);
nand U5838 (N_5838,N_913,N_2355);
nand U5839 (N_5839,N_635,N_2781);
and U5840 (N_5840,N_495,N_1863);
or U5841 (N_5841,N_916,N_1915);
nor U5842 (N_5842,N_2165,N_418);
nor U5843 (N_5843,N_2494,N_218);
nand U5844 (N_5844,N_1900,N_97);
nor U5845 (N_5845,N_543,N_257);
nor U5846 (N_5846,N_1112,N_1971);
and U5847 (N_5847,N_626,N_1826);
and U5848 (N_5848,N_2709,N_2046);
and U5849 (N_5849,N_2366,N_2297);
nor U5850 (N_5850,N_2818,N_1991);
nand U5851 (N_5851,N_35,N_1740);
nor U5852 (N_5852,N_755,N_2257);
nor U5853 (N_5853,N_2335,N_2997);
nand U5854 (N_5854,N_2310,N_168);
and U5855 (N_5855,N_1397,N_151);
and U5856 (N_5856,N_1603,N_1074);
or U5857 (N_5857,N_70,N_224);
nand U5858 (N_5858,N_862,N_2407);
nand U5859 (N_5859,N_2971,N_377);
or U5860 (N_5860,N_2771,N_914);
nand U5861 (N_5861,N_2251,N_425);
nand U5862 (N_5862,N_2114,N_776);
nor U5863 (N_5863,N_1411,N_2077);
nor U5864 (N_5864,N_1994,N_1381);
or U5865 (N_5865,N_1667,N_827);
or U5866 (N_5866,N_1689,N_944);
and U5867 (N_5867,N_1577,N_1054);
nor U5868 (N_5868,N_455,N_113);
nor U5869 (N_5869,N_2044,N_465);
and U5870 (N_5870,N_1123,N_695);
or U5871 (N_5871,N_491,N_2286);
and U5872 (N_5872,N_1265,N_2596);
or U5873 (N_5873,N_1550,N_2473);
nor U5874 (N_5874,N_1545,N_1397);
nand U5875 (N_5875,N_2474,N_1025);
and U5876 (N_5876,N_866,N_2264);
nor U5877 (N_5877,N_2298,N_2820);
or U5878 (N_5878,N_983,N_100);
nand U5879 (N_5879,N_2294,N_1035);
or U5880 (N_5880,N_2181,N_1604);
and U5881 (N_5881,N_2187,N_2644);
nand U5882 (N_5882,N_1584,N_941);
and U5883 (N_5883,N_312,N_681);
and U5884 (N_5884,N_73,N_899);
nand U5885 (N_5885,N_1968,N_1146);
xnor U5886 (N_5886,N_2623,N_2698);
nand U5887 (N_5887,N_1467,N_2333);
nand U5888 (N_5888,N_2478,N_2355);
or U5889 (N_5889,N_2285,N_264);
nand U5890 (N_5890,N_1663,N_2842);
nand U5891 (N_5891,N_939,N_193);
nand U5892 (N_5892,N_2661,N_2546);
and U5893 (N_5893,N_2453,N_2759);
nand U5894 (N_5894,N_2647,N_1371);
nor U5895 (N_5895,N_2102,N_1944);
and U5896 (N_5896,N_1396,N_100);
nor U5897 (N_5897,N_1945,N_2404);
nand U5898 (N_5898,N_100,N_91);
nand U5899 (N_5899,N_695,N_2830);
nand U5900 (N_5900,N_2891,N_1661);
nor U5901 (N_5901,N_1843,N_1440);
nand U5902 (N_5902,N_2582,N_1551);
nor U5903 (N_5903,N_1840,N_1406);
and U5904 (N_5904,N_1187,N_2951);
nand U5905 (N_5905,N_850,N_2930);
xnor U5906 (N_5906,N_2677,N_633);
nor U5907 (N_5907,N_1197,N_2836);
and U5908 (N_5908,N_1191,N_462);
xnor U5909 (N_5909,N_1635,N_2669);
or U5910 (N_5910,N_2578,N_279);
and U5911 (N_5911,N_2011,N_480);
nor U5912 (N_5912,N_96,N_1614);
nor U5913 (N_5913,N_129,N_1414);
nand U5914 (N_5914,N_2674,N_1638);
or U5915 (N_5915,N_788,N_151);
nand U5916 (N_5916,N_838,N_1909);
and U5917 (N_5917,N_115,N_2514);
or U5918 (N_5918,N_1272,N_2417);
nand U5919 (N_5919,N_1995,N_2672);
nand U5920 (N_5920,N_2529,N_746);
and U5921 (N_5921,N_2642,N_1105);
or U5922 (N_5922,N_2488,N_373);
or U5923 (N_5923,N_1344,N_2399);
nand U5924 (N_5924,N_47,N_1237);
or U5925 (N_5925,N_1552,N_2395);
nor U5926 (N_5926,N_1316,N_1663);
and U5927 (N_5927,N_979,N_2152);
and U5928 (N_5928,N_872,N_1258);
or U5929 (N_5929,N_1271,N_284);
nor U5930 (N_5930,N_1663,N_489);
and U5931 (N_5931,N_18,N_1899);
or U5932 (N_5932,N_891,N_1208);
nor U5933 (N_5933,N_1241,N_2261);
nor U5934 (N_5934,N_560,N_2137);
nor U5935 (N_5935,N_2691,N_2892);
nand U5936 (N_5936,N_1699,N_2845);
nand U5937 (N_5937,N_1632,N_957);
or U5938 (N_5938,N_1026,N_2754);
nand U5939 (N_5939,N_581,N_1614);
nor U5940 (N_5940,N_168,N_2424);
and U5941 (N_5941,N_2368,N_2009);
nand U5942 (N_5942,N_1558,N_716);
nand U5943 (N_5943,N_1850,N_545);
nor U5944 (N_5944,N_2588,N_1736);
nor U5945 (N_5945,N_1140,N_2204);
nor U5946 (N_5946,N_2341,N_757);
and U5947 (N_5947,N_1399,N_1140);
nand U5948 (N_5948,N_2147,N_1161);
and U5949 (N_5949,N_1144,N_1789);
or U5950 (N_5950,N_1181,N_2209);
or U5951 (N_5951,N_29,N_2386);
nand U5952 (N_5952,N_1278,N_15);
and U5953 (N_5953,N_547,N_2972);
or U5954 (N_5954,N_721,N_2227);
or U5955 (N_5955,N_608,N_874);
or U5956 (N_5956,N_2602,N_905);
and U5957 (N_5957,N_1291,N_2538);
and U5958 (N_5958,N_707,N_254);
or U5959 (N_5959,N_2102,N_892);
or U5960 (N_5960,N_1463,N_589);
and U5961 (N_5961,N_816,N_2941);
or U5962 (N_5962,N_769,N_2517);
and U5963 (N_5963,N_2261,N_831);
or U5964 (N_5964,N_1409,N_2373);
nand U5965 (N_5965,N_2830,N_308);
and U5966 (N_5966,N_1873,N_2524);
or U5967 (N_5967,N_1797,N_1804);
or U5968 (N_5968,N_304,N_67);
and U5969 (N_5969,N_1863,N_2560);
nand U5970 (N_5970,N_2467,N_23);
and U5971 (N_5971,N_2669,N_2497);
and U5972 (N_5972,N_1505,N_436);
nand U5973 (N_5973,N_8,N_1021);
xor U5974 (N_5974,N_429,N_2412);
and U5975 (N_5975,N_2493,N_1802);
nor U5976 (N_5976,N_2682,N_1193);
nor U5977 (N_5977,N_2745,N_923);
or U5978 (N_5978,N_421,N_1506);
nand U5979 (N_5979,N_2980,N_724);
and U5980 (N_5980,N_1641,N_1412);
and U5981 (N_5981,N_2883,N_1611);
nand U5982 (N_5982,N_208,N_1771);
nor U5983 (N_5983,N_281,N_2402);
and U5984 (N_5984,N_52,N_732);
or U5985 (N_5985,N_1102,N_2354);
or U5986 (N_5986,N_2384,N_257);
or U5987 (N_5987,N_2089,N_889);
nand U5988 (N_5988,N_1781,N_2859);
nor U5989 (N_5989,N_1249,N_2326);
nand U5990 (N_5990,N_672,N_1761);
or U5991 (N_5991,N_1467,N_1297);
nor U5992 (N_5992,N_1845,N_706);
nor U5993 (N_5993,N_722,N_74);
nor U5994 (N_5994,N_757,N_1281);
and U5995 (N_5995,N_1712,N_595);
and U5996 (N_5996,N_2130,N_1383);
nor U5997 (N_5997,N_2510,N_2719);
and U5998 (N_5998,N_1504,N_1490);
nand U5999 (N_5999,N_1695,N_2131);
nand U6000 (N_6000,N_3431,N_3864);
nor U6001 (N_6001,N_4465,N_5650);
nand U6002 (N_6002,N_4976,N_5429);
and U6003 (N_6003,N_3418,N_3153);
and U6004 (N_6004,N_3128,N_5448);
and U6005 (N_6005,N_4677,N_5521);
and U6006 (N_6006,N_3387,N_3097);
or U6007 (N_6007,N_5337,N_3425);
and U6008 (N_6008,N_3770,N_4748);
or U6009 (N_6009,N_4602,N_5737);
nor U6010 (N_6010,N_3808,N_4512);
nor U6011 (N_6011,N_3565,N_4781);
and U6012 (N_6012,N_4992,N_3477);
and U6013 (N_6013,N_5717,N_5689);
or U6014 (N_6014,N_5946,N_3371);
nand U6015 (N_6015,N_5925,N_4296);
and U6016 (N_6016,N_4409,N_4298);
and U6017 (N_6017,N_3703,N_5499);
nand U6018 (N_6018,N_5502,N_3672);
nor U6019 (N_6019,N_3372,N_5687);
and U6020 (N_6020,N_4425,N_4339);
or U6021 (N_6021,N_5576,N_4620);
nand U6022 (N_6022,N_4305,N_5658);
nand U6023 (N_6023,N_5122,N_5057);
xnor U6024 (N_6024,N_5998,N_5046);
and U6025 (N_6025,N_4913,N_4098);
or U6026 (N_6026,N_5978,N_3675);
or U6027 (N_6027,N_5697,N_4700);
xnor U6028 (N_6028,N_5995,N_4529);
nor U6029 (N_6029,N_5535,N_5056);
and U6030 (N_6030,N_4875,N_3901);
and U6031 (N_6031,N_5515,N_5793);
and U6032 (N_6032,N_3424,N_3484);
and U6033 (N_6033,N_5136,N_4192);
and U6034 (N_6034,N_4009,N_3743);
or U6035 (N_6035,N_3405,N_4536);
nand U6036 (N_6036,N_5613,N_4396);
and U6037 (N_6037,N_3676,N_5917);
nor U6038 (N_6038,N_3699,N_5338);
xnor U6039 (N_6039,N_4208,N_4744);
nand U6040 (N_6040,N_4825,N_5764);
nor U6041 (N_6041,N_3615,N_5482);
and U6042 (N_6042,N_4914,N_4254);
nor U6043 (N_6043,N_4293,N_3444);
and U6044 (N_6044,N_3490,N_3148);
and U6045 (N_6045,N_5811,N_3359);
nand U6046 (N_6046,N_5966,N_3796);
or U6047 (N_6047,N_3756,N_3328);
and U6048 (N_6048,N_5761,N_4872);
and U6049 (N_6049,N_4854,N_4849);
and U6050 (N_6050,N_3280,N_4017);
or U6051 (N_6051,N_5087,N_5125);
nand U6052 (N_6052,N_5231,N_3798);
nor U6053 (N_6053,N_4874,N_4742);
nor U6054 (N_6054,N_5437,N_4406);
nor U6055 (N_6055,N_4091,N_3980);
or U6056 (N_6056,N_5100,N_4183);
nand U6057 (N_6057,N_5339,N_4460);
xor U6058 (N_6058,N_3242,N_5428);
nor U6059 (N_6059,N_5478,N_3227);
nand U6060 (N_6060,N_4845,N_4281);
and U6061 (N_6061,N_4149,N_5410);
nor U6062 (N_6062,N_4168,N_3177);
nand U6063 (N_6063,N_3077,N_4717);
or U6064 (N_6064,N_5935,N_5920);
nand U6065 (N_6065,N_4611,N_5038);
nand U6066 (N_6066,N_5710,N_4637);
nor U6067 (N_6067,N_5875,N_5147);
and U6068 (N_6068,N_5467,N_4654);
and U6069 (N_6069,N_3529,N_3584);
or U6070 (N_6070,N_3940,N_4736);
nand U6071 (N_6071,N_5417,N_3353);
nand U6072 (N_6072,N_5831,N_3246);
or U6073 (N_6073,N_5566,N_5116);
and U6074 (N_6074,N_3028,N_5076);
or U6075 (N_6075,N_3916,N_3524);
nand U6076 (N_6076,N_4881,N_3181);
nand U6077 (N_6077,N_3818,N_4222);
and U6078 (N_6078,N_5355,N_3067);
nand U6079 (N_6079,N_5074,N_3514);
nand U6080 (N_6080,N_4193,N_3084);
nor U6081 (N_6081,N_5716,N_4649);
nor U6082 (N_6082,N_3481,N_4360);
nand U6083 (N_6083,N_5483,N_4210);
nand U6084 (N_6084,N_4747,N_3283);
nand U6085 (N_6085,N_4295,N_4152);
nor U6086 (N_6086,N_5516,N_4123);
and U6087 (N_6087,N_3960,N_4978);
nand U6088 (N_6088,N_4911,N_3170);
nand U6089 (N_6089,N_5911,N_5440);
and U6090 (N_6090,N_4055,N_5111);
nor U6091 (N_6091,N_3972,N_4609);
nand U6092 (N_6092,N_4363,N_4566);
nor U6093 (N_6093,N_5738,N_4246);
nor U6094 (N_6094,N_5106,N_5735);
and U6095 (N_6095,N_5776,N_5285);
or U6096 (N_6096,N_3171,N_3889);
or U6097 (N_6097,N_3593,N_5987);
nor U6098 (N_6098,N_3741,N_3230);
nor U6099 (N_6099,N_4114,N_4738);
and U6100 (N_6100,N_4886,N_4767);
and U6101 (N_6101,N_4134,N_3637);
and U6102 (N_6102,N_3446,N_3517);
nand U6103 (N_6103,N_5117,N_4085);
and U6104 (N_6104,N_5442,N_5178);
nand U6105 (N_6105,N_5715,N_4993);
and U6106 (N_6106,N_5041,N_5379);
and U6107 (N_6107,N_4585,N_4335);
nor U6108 (N_6108,N_3755,N_4587);
nand U6109 (N_6109,N_3352,N_3852);
or U6110 (N_6110,N_5529,N_3695);
nor U6111 (N_6111,N_5809,N_5193);
nand U6112 (N_6112,N_3948,N_4682);
and U6113 (N_6113,N_4835,N_5629);
and U6114 (N_6114,N_5019,N_3961);
and U6115 (N_6115,N_4545,N_5077);
or U6116 (N_6116,N_5507,N_5278);
and U6117 (N_6117,N_3056,N_5272);
or U6118 (N_6118,N_5066,N_4066);
xor U6119 (N_6119,N_4142,N_4464);
nand U6120 (N_6120,N_4000,N_4773);
nor U6121 (N_6121,N_5684,N_5099);
and U6122 (N_6122,N_3156,N_4885);
xnor U6123 (N_6123,N_5534,N_5949);
nand U6124 (N_6124,N_4571,N_4975);
nor U6125 (N_6125,N_4211,N_3503);
nor U6126 (N_6126,N_5127,N_4701);
nor U6127 (N_6127,N_5146,N_4321);
nor U6128 (N_6128,N_3908,N_5196);
or U6129 (N_6129,N_5557,N_4236);
and U6130 (N_6130,N_3164,N_4184);
or U6131 (N_6131,N_5543,N_3971);
and U6132 (N_6132,N_4894,N_5739);
xor U6133 (N_6133,N_4974,N_4475);
and U6134 (N_6134,N_3689,N_5149);
nor U6135 (N_6135,N_5874,N_5208);
nor U6136 (N_6136,N_5003,N_5577);
nor U6137 (N_6137,N_4387,N_4564);
or U6138 (N_6138,N_5470,N_5651);
or U6139 (N_6139,N_4218,N_3992);
nor U6140 (N_6140,N_3112,N_3044);
nand U6141 (N_6141,N_3832,N_5936);
or U6142 (N_6142,N_3793,N_4954);
nand U6143 (N_6143,N_5441,N_3662);
nand U6144 (N_6144,N_4333,N_4697);
nor U6145 (N_6145,N_4725,N_4989);
nand U6146 (N_6146,N_4336,N_4837);
nor U6147 (N_6147,N_4382,N_5524);
and U6148 (N_6148,N_5645,N_5401);
or U6149 (N_6149,N_3654,N_5615);
or U6150 (N_6150,N_5519,N_3422);
nand U6151 (N_6151,N_4921,N_4521);
nand U6152 (N_6152,N_3567,N_4081);
and U6153 (N_6153,N_3188,N_4855);
nand U6154 (N_6154,N_4705,N_4803);
and U6155 (N_6155,N_3101,N_5675);
or U6156 (N_6156,N_5720,N_4526);
nor U6157 (N_6157,N_5606,N_5980);
and U6158 (N_6158,N_4122,N_4117);
and U6159 (N_6159,N_4719,N_4356);
or U6160 (N_6160,N_3554,N_3746);
and U6161 (N_6161,N_4371,N_3288);
nor U6162 (N_6162,N_5725,N_4005);
nand U6163 (N_6163,N_3473,N_4121);
nand U6164 (N_6164,N_3850,N_3111);
nand U6165 (N_6165,N_4935,N_3210);
nor U6166 (N_6166,N_5544,N_3863);
nor U6167 (N_6167,N_5086,N_3628);
nand U6168 (N_6168,N_3932,N_4088);
and U6169 (N_6169,N_5032,N_3344);
nand U6170 (N_6170,N_4632,N_3732);
nor U6171 (N_6171,N_4870,N_4801);
nor U6172 (N_6172,N_3393,N_4795);
and U6173 (N_6173,N_5113,N_5723);
nor U6174 (N_6174,N_4805,N_5702);
nor U6175 (N_6175,N_5150,N_5618);
or U6176 (N_6176,N_3331,N_5590);
nor U6177 (N_6177,N_3193,N_4096);
or U6178 (N_6178,N_4815,N_3778);
nor U6179 (N_6179,N_3933,N_5876);
and U6180 (N_6180,N_3979,N_4237);
nor U6181 (N_6181,N_3797,N_3358);
nor U6182 (N_6182,N_3356,N_4228);
nand U6183 (N_6183,N_3590,N_3069);
nor U6184 (N_6184,N_4033,N_4561);
and U6185 (N_6185,N_4482,N_5938);
nor U6186 (N_6186,N_3475,N_4752);
or U6187 (N_6187,N_3251,N_5414);
and U6188 (N_6188,N_4608,N_3526);
xor U6189 (N_6189,N_3127,N_3836);
or U6190 (N_6190,N_5387,N_4514);
or U6191 (N_6191,N_3286,N_3589);
nand U6192 (N_6192,N_5011,N_4770);
nor U6193 (N_6193,N_3854,N_3008);
and U6194 (N_6194,N_4645,N_5334);
or U6195 (N_6195,N_4588,N_5786);
nand U6196 (N_6196,N_3744,N_5202);
or U6197 (N_6197,N_5232,N_4289);
or U6198 (N_6198,N_4050,N_3792);
xnor U6199 (N_6199,N_5868,N_3160);
nand U6200 (N_6200,N_3644,N_5632);
and U6201 (N_6201,N_4554,N_4657);
and U6202 (N_6202,N_5413,N_4633);
and U6203 (N_6203,N_4397,N_3277);
nor U6204 (N_6204,N_3781,N_3244);
and U6205 (N_6205,N_4723,N_3178);
or U6206 (N_6206,N_5281,N_5489);
nor U6207 (N_6207,N_4515,N_3994);
or U6208 (N_6208,N_5732,N_3061);
nand U6209 (N_6209,N_4097,N_4120);
or U6210 (N_6210,N_3489,N_3624);
and U6211 (N_6211,N_4901,N_5678);
nor U6212 (N_6212,N_5291,N_4916);
nor U6213 (N_6213,N_5886,N_4337);
or U6214 (N_6214,N_5973,N_5797);
and U6215 (N_6215,N_3954,N_5711);
and U6216 (N_6216,N_4979,N_5770);
and U6217 (N_6217,N_4955,N_3935);
and U6218 (N_6218,N_3316,N_5135);
nor U6219 (N_6219,N_5906,N_5424);
and U6220 (N_6220,N_5423,N_3116);
nand U6221 (N_6221,N_5828,N_3395);
and U6222 (N_6222,N_3597,N_5888);
and U6223 (N_6223,N_3555,N_4500);
nor U6224 (N_6224,N_3301,N_5255);
nand U6225 (N_6225,N_4634,N_5696);
nand U6226 (N_6226,N_3812,N_4413);
or U6227 (N_6227,N_4613,N_4660);
or U6228 (N_6228,N_4900,N_3071);
or U6229 (N_6229,N_5840,N_5755);
xnor U6230 (N_6230,N_5071,N_5181);
nor U6231 (N_6231,N_5088,N_5343);
and U6232 (N_6232,N_5771,N_5913);
nor U6233 (N_6233,N_5060,N_3007);
nand U6234 (N_6234,N_5092,N_5815);
or U6235 (N_6235,N_4219,N_5598);
nor U6236 (N_6236,N_3791,N_3727);
nor U6237 (N_6237,N_4197,N_5533);
or U6238 (N_6238,N_5471,N_5638);
nor U6239 (N_6239,N_5054,N_4675);
xnor U6240 (N_6240,N_3373,N_5703);
and U6241 (N_6241,N_4313,N_4204);
and U6242 (N_6242,N_4386,N_3035);
nand U6243 (N_6243,N_5729,N_5950);
and U6244 (N_6244,N_3974,N_5139);
or U6245 (N_6245,N_4389,N_3085);
nor U6246 (N_6246,N_5295,N_3919);
nor U6247 (N_6247,N_5941,N_4572);
nor U6248 (N_6248,N_5070,N_5619);
or U6249 (N_6249,N_5760,N_5751);
and U6250 (N_6250,N_5922,N_3494);
or U6251 (N_6251,N_3773,N_3653);
xnor U6252 (N_6252,N_4285,N_5861);
nand U6253 (N_6253,N_4786,N_4902);
and U6254 (N_6254,N_4449,N_4473);
nand U6255 (N_6255,N_5848,N_4314);
or U6256 (N_6256,N_4531,N_4599);
nor U6257 (N_6257,N_3876,N_5241);
and U6258 (N_6258,N_4164,N_5806);
or U6259 (N_6259,N_3783,N_5276);
nor U6260 (N_6260,N_4113,N_4787);
nor U6261 (N_6261,N_5186,N_3264);
or U6262 (N_6262,N_4539,N_5227);
nor U6263 (N_6263,N_4368,N_5827);
nand U6264 (N_6264,N_3263,N_4398);
or U6265 (N_6265,N_5914,N_5513);
or U6266 (N_6266,N_5115,N_5787);
nand U6267 (N_6267,N_4630,N_5211);
and U6268 (N_6268,N_4733,N_3076);
nor U6269 (N_6269,N_5944,N_5934);
or U6270 (N_6270,N_3437,N_4560);
nor U6271 (N_6271,N_3849,N_5532);
nand U6272 (N_6272,N_5568,N_3369);
nand U6273 (N_6273,N_3175,N_3815);
nand U6274 (N_6274,N_5965,N_5096);
and U6275 (N_6275,N_4732,N_3273);
and U6276 (N_6276,N_3993,N_5319);
nor U6277 (N_6277,N_4361,N_4683);
or U6278 (N_6278,N_5592,N_4696);
nor U6279 (N_6279,N_3925,N_5915);
or U6280 (N_6280,N_4138,N_5091);
nand U6281 (N_6281,N_3274,N_5880);
and U6282 (N_6282,N_4619,N_5152);
nand U6283 (N_6283,N_4816,N_3313);
and U6284 (N_6284,N_3645,N_5020);
nor U6285 (N_6285,N_5604,N_4282);
and U6286 (N_6286,N_3066,N_3575);
and U6287 (N_6287,N_3327,N_3197);
nand U6288 (N_6288,N_5372,N_5652);
nor U6289 (N_6289,N_4109,N_4960);
and U6290 (N_6290,N_5169,N_4258);
or U6291 (N_6291,N_3296,N_4132);
xnor U6292 (N_6292,N_4022,N_5909);
nor U6293 (N_6293,N_3337,N_5389);
or U6294 (N_6294,N_4325,N_3633);
or U6295 (N_6295,N_5967,N_4294);
nor U6296 (N_6296,N_4411,N_5674);
nand U6297 (N_6297,N_3539,N_5258);
nand U6298 (N_6298,N_3894,N_3194);
nand U6299 (N_6299,N_5328,N_4330);
and U6300 (N_6300,N_5741,N_3949);
and U6301 (N_6301,N_5302,N_5539);
or U6302 (N_6302,N_3673,N_3687);
nand U6303 (N_6303,N_4140,N_3411);
nand U6304 (N_6304,N_4947,N_5745);
nand U6305 (N_6305,N_4372,N_3825);
or U6306 (N_6306,N_3043,N_3198);
and U6307 (N_6307,N_5602,N_3810);
and U6308 (N_6308,N_4474,N_4944);
or U6309 (N_6309,N_3135,N_5784);
nand U6310 (N_6310,N_5444,N_4766);
and U6311 (N_6311,N_4972,N_5154);
nand U6312 (N_6312,N_3239,N_5981);
nand U6313 (N_6313,N_3956,N_3113);
nand U6314 (N_6314,N_3325,N_4789);
and U6315 (N_6315,N_3310,N_5933);
and U6316 (N_6316,N_3142,N_4821);
or U6317 (N_6317,N_4812,N_3147);
or U6318 (N_6318,N_4135,N_5249);
nand U6319 (N_6319,N_5816,N_3159);
nand U6320 (N_6320,N_4999,N_5655);
and U6321 (N_6321,N_4235,N_4756);
nor U6322 (N_6322,N_4720,N_5537);
or U6323 (N_6323,N_4511,N_5826);
and U6324 (N_6324,N_3338,N_5744);
nand U6325 (N_6325,N_4390,N_4205);
nand U6326 (N_6326,N_4112,N_3723);
nor U6327 (N_6327,N_5841,N_4238);
or U6328 (N_6328,N_3784,N_3833);
nand U6329 (N_6329,N_5554,N_3132);
nand U6330 (N_6330,N_3218,N_5589);
nand U6331 (N_6331,N_4859,N_5182);
nor U6332 (N_6332,N_5986,N_5305);
and U6333 (N_6333,N_3285,N_4257);
and U6334 (N_6334,N_3923,N_5010);
and U6335 (N_6335,N_3718,N_4232);
xnor U6336 (N_6336,N_5224,N_5673);
xnor U6337 (N_6337,N_5048,N_5317);
and U6338 (N_6338,N_4353,N_4365);
nor U6339 (N_6339,N_3822,N_3724);
or U6340 (N_6340,N_3862,N_4148);
and U6341 (N_6341,N_5468,N_4563);
or U6342 (N_6342,N_5792,N_4250);
nand U6343 (N_6343,N_3143,N_5439);
nand U6344 (N_6344,N_5035,N_3501);
or U6345 (N_6345,N_3060,N_4702);
nor U6346 (N_6346,N_4968,N_5223);
nand U6347 (N_6347,N_3911,N_5392);
nor U6348 (N_6348,N_4497,N_5399);
nor U6349 (N_6349,N_3614,N_4084);
and U6350 (N_6350,N_3169,N_5068);
or U6351 (N_6351,N_4827,N_5871);
nor U6352 (N_6352,N_3802,N_4404);
nand U6353 (N_6353,N_4842,N_3449);
nor U6354 (N_6354,N_5594,N_3226);
nand U6355 (N_6355,N_4503,N_5203);
and U6356 (N_6356,N_5926,N_5120);
nor U6357 (N_6357,N_3383,N_3323);
nand U6358 (N_6358,N_3531,N_4590);
nand U6359 (N_6359,N_5904,N_5885);
and U6360 (N_6360,N_3070,N_5962);
or U6361 (N_6361,N_3161,N_5252);
and U6362 (N_6362,N_3895,N_4430);
or U6363 (N_6363,N_3311,N_3176);
nand U6364 (N_6364,N_4857,N_5310);
or U6365 (N_6365,N_4984,N_4492);
or U6366 (N_6366,N_5849,N_3528);
or U6367 (N_6367,N_5939,N_3467);
or U6368 (N_6368,N_5435,N_4057);
nor U6369 (N_6369,N_3938,N_4119);
and U6370 (N_6370,N_4950,N_4759);
and U6371 (N_6371,N_5833,N_5700);
or U6372 (N_6372,N_4791,N_3382);
or U6373 (N_6373,N_3749,N_3771);
nor U6374 (N_6374,N_4444,N_3155);
or U6375 (N_6375,N_4153,N_3618);
nand U6376 (N_6376,N_3655,N_4684);
nor U6377 (N_6377,N_4297,N_3537);
nor U6378 (N_6378,N_5599,N_5743);
nor U6379 (N_6379,N_4504,N_5426);
and U6380 (N_6380,N_5677,N_5336);
nand U6381 (N_6381,N_4056,N_4672);
or U6382 (N_6382,N_5930,N_3388);
nand U6383 (N_6383,N_4410,N_5190);
nand U6384 (N_6384,N_4259,N_4061);
nor U6385 (N_6385,N_3897,N_5553);
and U6386 (N_6386,N_3126,N_3611);
or U6387 (N_6387,N_5979,N_5897);
nor U6388 (N_6388,N_4871,N_4169);
and U6389 (N_6389,N_5958,N_4090);
nor U6390 (N_6390,N_5311,N_4170);
and U6391 (N_6391,N_5912,N_3282);
nor U6392 (N_6392,N_5402,N_4493);
and U6393 (N_6393,N_5664,N_5701);
or U6394 (N_6394,N_3920,N_5158);
and U6395 (N_6395,N_5342,N_5246);
or U6396 (N_6396,N_4039,N_5916);
nor U6397 (N_6397,N_3613,N_3879);
or U6398 (N_6398,N_3354,N_3728);
nand U6399 (N_6399,N_3694,N_3495);
and U6400 (N_6400,N_4663,N_5900);
nand U6401 (N_6401,N_5176,N_3601);
nor U6402 (N_6402,N_5090,N_5366);
nor U6403 (N_6403,N_4846,N_3981);
nor U6404 (N_6404,N_4762,N_4342);
nand U6405 (N_6405,N_5460,N_5405);
nor U6406 (N_6406,N_3406,N_4729);
nor U6407 (N_6407,N_4704,N_4334);
or U6408 (N_6408,N_5260,N_5692);
and U6409 (N_6409,N_3023,N_4015);
nor U6410 (N_6410,N_5518,N_3869);
or U6411 (N_6411,N_3572,N_4708);
nor U6412 (N_6412,N_5061,N_4195);
nand U6413 (N_6413,N_3267,N_3435);
nand U6414 (N_6414,N_5037,N_3020);
nor U6415 (N_6415,N_5514,N_3891);
or U6416 (N_6416,N_5321,N_3258);
nor U6417 (N_6417,N_4662,N_4376);
nor U6418 (N_6418,N_5271,N_4597);
and U6419 (N_6419,N_3394,N_5824);
nand U6420 (N_6420,N_3570,N_3224);
or U6421 (N_6421,N_4042,N_5982);
nor U6422 (N_6422,N_3685,N_5728);
or U6423 (N_6423,N_5330,N_3766);
or U6424 (N_6424,N_3396,N_5304);
nand U6425 (N_6425,N_4847,N_3721);
nor U6426 (N_6426,N_5298,N_3221);
and U6427 (N_6427,N_3105,N_4273);
and U6428 (N_6428,N_5286,N_5501);
and U6429 (N_6429,N_3408,N_4832);
or U6430 (N_6430,N_4127,N_4030);
and U6431 (N_6431,N_3650,N_3429);
nor U6432 (N_6432,N_3509,N_4668);
or U6433 (N_6433,N_4693,N_3217);
nand U6434 (N_6434,N_3299,N_4352);
nand U6435 (N_6435,N_5558,N_5836);
nor U6436 (N_6436,N_5381,N_4242);
or U6437 (N_6437,N_4740,N_3585);
nor U6438 (N_6438,N_3038,N_3760);
and U6439 (N_6439,N_5213,N_4679);
nor U6440 (N_6440,N_4291,N_4344);
and U6441 (N_6441,N_3631,N_5403);
and U6442 (N_6442,N_4179,N_4074);
xor U6443 (N_6443,N_3314,N_3366);
nor U6444 (N_6444,N_3269,N_3245);
nand U6445 (N_6445,N_3996,N_3541);
and U6446 (N_6446,N_3573,N_3208);
nand U6447 (N_6447,N_5660,N_3720);
or U6448 (N_6448,N_3426,N_5858);
and U6449 (N_6449,N_5376,N_3665);
and U6450 (N_6450,N_3779,N_3146);
and U6451 (N_6451,N_3834,N_5206);
nand U6452 (N_6452,N_3885,N_5477);
and U6453 (N_6453,N_4324,N_3152);
nand U6454 (N_6454,N_5026,N_4967);
nor U6455 (N_6455,N_4498,N_5726);
nand U6456 (N_6456,N_5431,N_4949);
or U6457 (N_6457,N_5487,N_4818);
xor U6458 (N_6458,N_4459,N_5550);
or U6459 (N_6459,N_3859,N_4472);
and U6460 (N_6460,N_3603,N_5970);
and U6461 (N_6461,N_4067,N_5000);
nor U6462 (N_6462,N_3478,N_3059);
or U6463 (N_6463,N_5004,N_4265);
or U6464 (N_6464,N_4369,N_3017);
or U6465 (N_6465,N_4438,N_3065);
xor U6466 (N_6466,N_4006,N_4480);
nor U6467 (N_6467,N_5765,N_4627);
or U6468 (N_6468,N_4661,N_3690);
nand U6469 (N_6469,N_4364,N_3738);
and U6470 (N_6470,N_3693,N_3364);
nor U6471 (N_6471,N_3691,N_3131);
or U6472 (N_6472,N_4605,N_4850);
and U6473 (N_6473,N_5782,N_3622);
or U6474 (N_6474,N_3204,N_4604);
nand U6475 (N_6475,N_3646,N_5842);
nand U6476 (N_6476,N_3875,N_3683);
nor U6477 (N_6477,N_4681,N_3647);
and U6478 (N_6478,N_5648,N_5546);
or U6479 (N_6479,N_4690,N_4167);
nor U6480 (N_6480,N_5924,N_3397);
or U6481 (N_6481,N_5772,N_5707);
and U6482 (N_6482,N_3936,N_3525);
or U6483 (N_6483,N_5869,N_3568);
and U6484 (N_6484,N_5974,N_4078);
or U6485 (N_6485,N_4552,N_5750);
nand U6486 (N_6486,N_4402,N_3360);
nor U6487 (N_6487,N_3707,N_5862);
or U6488 (N_6488,N_5264,N_3623);
or U6489 (N_6489,N_5894,N_5378);
nand U6490 (N_6490,N_3322,N_5945);
nor U6491 (N_6491,N_4505,N_4150);
and U6492 (N_6492,N_3817,N_3297);
nor U6493 (N_6493,N_5472,N_3203);
nor U6494 (N_6494,N_3835,N_3641);
nor U6495 (N_6495,N_4692,N_3051);
nand U6496 (N_6496,N_3074,N_3878);
or U6497 (N_6497,N_4519,N_3752);
nor U6498 (N_6498,N_4349,N_4118);
nor U6499 (N_6499,N_4549,N_5273);
nand U6500 (N_6500,N_3984,N_4403);
nor U6501 (N_6501,N_4087,N_5572);
nand U6502 (N_6502,N_4839,N_4893);
and U6503 (N_6503,N_4925,N_5957);
nor U6504 (N_6504,N_5891,N_5463);
nand U6505 (N_6505,N_4485,N_4929);
xnor U6506 (N_6506,N_5722,N_5433);
nand U6507 (N_6507,N_3368,N_4592);
and U6508 (N_6508,N_4730,N_3860);
and U6509 (N_6509,N_4421,N_3710);
nor U6510 (N_6510,N_3669,N_3047);
nor U6511 (N_6511,N_5261,N_4290);
nor U6512 (N_6512,N_4309,N_5996);
and U6513 (N_6513,N_5045,N_3305);
or U6514 (N_6514,N_4071,N_3440);
nor U6515 (N_6515,N_3384,N_4327);
nor U6516 (N_6516,N_3416,N_5051);
nand U6517 (N_6517,N_4046,N_4938);
and U6518 (N_6518,N_3341,N_5634);
nor U6519 (N_6519,N_4694,N_5835);
and U6520 (N_6520,N_3742,N_3846);
nor U6521 (N_6521,N_3332,N_4509);
nor U6522 (N_6522,N_4624,N_3540);
and U6523 (N_6523,N_5341,N_3172);
nor U6524 (N_6524,N_4674,N_4841);
and U6525 (N_6525,N_3913,N_5119);
nor U6526 (N_6526,N_4895,N_4125);
or U6527 (N_6527,N_5795,N_5657);
nand U6528 (N_6528,N_5306,N_4317);
nand U6529 (N_6529,N_3385,N_3390);
and U6530 (N_6530,N_5394,N_5465);
and U6531 (N_6531,N_5500,N_3480);
nor U6532 (N_6532,N_4367,N_3576);
nor U6533 (N_6533,N_3870,N_3026);
nand U6534 (N_6534,N_4276,N_4769);
and U6535 (N_6535,N_5665,N_3782);
xnor U6536 (N_6536,N_4920,N_5985);
or U6537 (N_6537,N_4016,N_4506);
or U6538 (N_6538,N_4058,N_5110);
and U6539 (N_6539,N_4185,N_3561);
and U6540 (N_6540,N_3963,N_4092);
nand U6541 (N_6541,N_4653,N_4049);
nand U6542 (N_6542,N_4277,N_5253);
and U6543 (N_6543,N_5571,N_3093);
nand U6544 (N_6544,N_5748,N_5156);
or U6545 (N_6545,N_4964,N_3536);
and U6546 (N_6546,N_3237,N_5617);
nand U6547 (N_6547,N_5714,N_5685);
or U6548 (N_6548,N_4200,N_5250);
and U6549 (N_6549,N_4023,N_4263);
nor U6550 (N_6550,N_4593,N_5391);
xnor U6551 (N_6551,N_5641,N_5427);
nor U6552 (N_6552,N_3518,N_3873);
and U6553 (N_6553,N_4959,N_4570);
nor U6554 (N_6554,N_3780,N_4130);
nand U6555 (N_6555,N_4555,N_3233);
nand U6556 (N_6556,N_3037,N_3110);
nor U6557 (N_6557,N_4378,N_5480);
or U6558 (N_6558,N_5730,N_3592);
xor U6559 (N_6559,N_4206,N_4230);
or U6560 (N_6560,N_3574,N_5560);
or U6561 (N_6561,N_3058,N_5455);
nor U6562 (N_6562,N_5575,N_5234);
or U6563 (N_6563,N_4685,N_4380);
nor U6564 (N_6564,N_3086,N_3365);
nor U6565 (N_6565,N_4477,N_3900);
and U6566 (N_6566,N_5733,N_3763);
nand U6567 (N_6567,N_4840,N_4798);
nand U6568 (N_6568,N_3019,N_3001);
nor U6569 (N_6569,N_4524,N_4707);
and U6570 (N_6570,N_4350,N_5370);
nor U6571 (N_6571,N_3123,N_5309);
nor U6572 (N_6572,N_4063,N_3904);
or U6573 (N_6573,N_3031,N_3166);
and U6574 (N_6574,N_3108,N_5012);
nand U6575 (N_6575,N_4343,N_5667);
nand U6576 (N_6576,N_3813,N_3626);
nand U6577 (N_6577,N_4621,N_3349);
nor U6578 (N_6578,N_5143,N_3287);
and U6579 (N_6579,N_4287,N_3636);
nand U6580 (N_6580,N_5721,N_5984);
nor U6581 (N_6581,N_3215,N_5199);
nor U6582 (N_6582,N_3458,N_5397);
and U6583 (N_6583,N_5121,N_5850);
or U6584 (N_6584,N_5138,N_5919);
nand U6585 (N_6585,N_4864,N_3519);
nor U6586 (N_6586,N_3289,N_3104);
nand U6587 (N_6587,N_4393,N_4182);
or U6588 (N_6588,N_3124,N_5595);
and U6589 (N_6589,N_3857,N_5420);
and U6590 (N_6590,N_5396,N_5819);
nor U6591 (N_6591,N_4256,N_4479);
nor U6592 (N_6592,N_4541,N_5623);
or U6593 (N_6593,N_5921,N_3887);
or U6594 (N_6594,N_3141,N_4836);
or U6595 (N_6595,N_3684,N_4507);
and U6596 (N_6596,N_4434,N_5857);
and U6597 (N_6597,N_3516,N_5541);
and U6598 (N_6598,N_4484,N_4248);
nor U6599 (N_6599,N_5503,N_5691);
and U6600 (N_6600,N_4688,N_3997);
nand U6601 (N_6601,N_5062,N_3604);
or U6602 (N_6602,N_3339,N_5931);
nor U6603 (N_6603,N_4312,N_3241);
nand U6604 (N_6604,N_4728,N_4936);
nand U6605 (N_6605,N_3621,N_4817);
and U6606 (N_6606,N_5422,N_4429);
nor U6607 (N_6607,N_5852,N_3415);
nor U6608 (N_6608,N_3229,N_4819);
or U6609 (N_6609,N_4851,N_4158);
and U6610 (N_6610,N_4251,N_5588);
nand U6611 (N_6611,N_5130,N_3520);
nor U6612 (N_6612,N_3988,N_5251);
nand U6613 (N_6613,N_5953,N_4809);
nor U6614 (N_6614,N_5614,N_5570);
nand U6615 (N_6615,N_4942,N_5326);
xnor U6616 (N_6616,N_4223,N_3046);
xnor U6617 (N_6617,N_5040,N_5450);
nor U6618 (N_6618,N_3423,N_4060);
nand U6619 (N_6619,N_5277,N_4869);
or U6620 (N_6620,N_3602,N_3795);
and U6621 (N_6621,N_5031,N_5959);
nor U6622 (N_6622,N_4043,N_5990);
and U6623 (N_6623,N_3004,N_5325);
or U6624 (N_6624,N_3206,N_4502);
nor U6625 (N_6625,N_3102,N_5740);
nor U6626 (N_6626,N_3542,N_3250);
nand U6627 (N_6627,N_3660,N_5168);
or U6628 (N_6628,N_4414,N_5228);
or U6629 (N_6629,N_3402,N_4601);
nand U6630 (N_6630,N_5591,N_3033);
or U6631 (N_6631,N_3133,N_4550);
nand U6632 (N_6632,N_4443,N_5633);
or U6633 (N_6633,N_3973,N_4777);
and U6634 (N_6634,N_3534,N_5690);
nor U6635 (N_6635,N_5663,N_5348);
nor U6636 (N_6636,N_3034,N_3048);
nor U6637 (N_6637,N_4930,N_4635);
and U6638 (N_6638,N_3522,N_5932);
nand U6639 (N_6639,N_3874,N_5453);
nand U6640 (N_6640,N_4014,N_3421);
and U6641 (N_6641,N_3309,N_3945);
and U6642 (N_6642,N_5177,N_3959);
nor U6643 (N_6643,N_3357,N_4626);
nand U6644 (N_6644,N_4909,N_5484);
nor U6645 (N_6645,N_5216,N_5447);
or U6646 (N_6646,N_5180,N_5351);
nand U6647 (N_6647,N_4147,N_4826);
nor U6648 (N_6648,N_3045,N_5574);
or U6649 (N_6649,N_5357,N_5905);
nand U6650 (N_6650,N_3042,N_5605);
nand U6651 (N_6651,N_5752,N_3000);
and U6652 (N_6652,N_5805,N_5044);
nor U6653 (N_6653,N_4904,N_5292);
and U6654 (N_6654,N_3191,N_5890);
nand U6655 (N_6655,N_4784,N_5621);
nand U6656 (N_6656,N_3591,N_3906);
or U6657 (N_6657,N_4143,N_3201);
and U6658 (N_6658,N_4532,N_4658);
and U6659 (N_6659,N_5364,N_3736);
or U6660 (N_6660,N_3543,N_5346);
or U6661 (N_6661,N_5775,N_5896);
or U6662 (N_6662,N_4165,N_4408);
and U6663 (N_6663,N_4220,N_5257);
or U6664 (N_6664,N_4062,N_5055);
or U6665 (N_6665,N_4155,N_4640);
nor U6666 (N_6666,N_5545,N_4173);
or U6667 (N_6667,N_5018,N_3951);
and U6668 (N_6668,N_4603,N_3082);
or U6669 (N_6669,N_4031,N_4244);
nor U6670 (N_6670,N_5065,N_3549);
or U6671 (N_6671,N_5625,N_5009);
nand U6672 (N_6672,N_5197,N_5324);
and U6673 (N_6673,N_4466,N_3329);
nor U6674 (N_6674,N_5390,N_4476);
or U6675 (N_6675,N_4086,N_5043);
and U6676 (N_6676,N_3612,N_5731);
and U6677 (N_6677,N_4568,N_4686);
and U6678 (N_6678,N_5354,N_4889);
nor U6679 (N_6679,N_3376,N_5385);
xor U6680 (N_6680,N_5800,N_3073);
nor U6681 (N_6681,N_5778,N_4734);
xor U6682 (N_6682,N_3789,N_5587);
or U6683 (N_6683,N_4037,N_4780);
nand U6684 (N_6684,N_3138,N_3452);
nor U6685 (N_6685,N_3137,N_5126);
nand U6686 (N_6686,N_4041,N_4065);
and U6687 (N_6687,N_4415,N_3991);
and U6688 (N_6688,N_4982,N_3697);
xnor U6689 (N_6689,N_3461,N_3014);
and U6690 (N_6690,N_3816,N_5411);
nand U6691 (N_6691,N_3187,N_4785);
or U6692 (N_6692,N_3335,N_4956);
nor U6693 (N_6693,N_5412,N_4024);
xor U6694 (N_6694,N_5129,N_4329);
and U6695 (N_6695,N_5893,N_5192);
nand U6696 (N_6696,N_3843,N_3312);
and U6697 (N_6697,N_5892,N_4530);
and U6698 (N_6698,N_5742,N_4618);
or U6699 (N_6699,N_3260,N_5215);
and U6700 (N_6700,N_4388,N_4743);
and U6701 (N_6701,N_3050,N_5308);
or U6702 (N_6702,N_4517,N_5832);
nor U6703 (N_6703,N_5872,N_4496);
or U6704 (N_6704,N_5331,N_3943);
and U6705 (N_6705,N_4928,N_3566);
nand U6706 (N_6706,N_5112,N_5218);
nand U6707 (N_6707,N_5993,N_5683);
or U6708 (N_6708,N_4012,N_3748);
or U6709 (N_6709,N_3404,N_3677);
nand U6710 (N_6710,N_5608,N_3100);
xor U6711 (N_6711,N_3212,N_4646);
and U6712 (N_6712,N_3702,N_4562);
nand U6713 (N_6713,N_5415,N_3451);
nand U6714 (N_6714,N_5548,N_4594);
nor U6715 (N_6715,N_5024,N_4581);
or U6716 (N_6716,N_4775,N_4412);
or U6717 (N_6717,N_3284,N_3807);
nand U6718 (N_6718,N_3346,N_4834);
nand U6719 (N_6719,N_3715,N_3454);
and U6720 (N_6720,N_3236,N_5407);
and U6721 (N_6721,N_4103,N_5166);
and U6722 (N_6722,N_3564,N_5290);
nor U6723 (N_6723,N_3302,N_3294);
nor U6724 (N_6724,N_4643,N_4101);
nor U6725 (N_6725,N_3207,N_4932);
or U6726 (N_6726,N_4283,N_3428);
and U6727 (N_6727,N_3381,N_4948);
nor U6728 (N_6728,N_3999,N_3083);
and U6729 (N_6729,N_3455,N_5404);
or U6730 (N_6730,N_3588,N_3064);
or U6731 (N_6731,N_3594,N_4946);
nand U6732 (N_6732,N_5746,N_4064);
and U6733 (N_6733,N_3546,N_5901);
or U6734 (N_6734,N_5466,N_4567);
or U6735 (N_6735,N_5694,N_5528);
nand U6736 (N_6736,N_4980,N_5363);
nor U6737 (N_6737,N_5994,N_4310);
or U6738 (N_6738,N_3121,N_5229);
xnor U6739 (N_6739,N_4796,N_3814);
or U6740 (N_6740,N_5016,N_4741);
or U6741 (N_6741,N_4939,N_3745);
or U6742 (N_6742,N_5918,N_3453);
or U6743 (N_6743,N_5159,N_5093);
nor U6744 (N_6744,N_4527,N_3513);
nand U6745 (N_6745,N_3103,N_3247);
and U6746 (N_6746,N_4797,N_4877);
and U6747 (N_6747,N_5860,N_4416);
or U6748 (N_6748,N_5194,N_5352);
nor U6749 (N_6749,N_5124,N_3717);
or U6750 (N_6750,N_4659,N_5774);
nand U6751 (N_6751,N_5567,N_4440);
or U6752 (N_6752,N_5353,N_4824);
or U6753 (N_6753,N_5347,N_3800);
nor U6754 (N_6754,N_4059,N_4912);
nand U6755 (N_6755,N_4216,N_4188);
nor U6756 (N_6756,N_5247,N_5386);
nand U6757 (N_6757,N_5844,N_5421);
and U6758 (N_6758,N_5165,N_5243);
and U6759 (N_6759,N_3506,N_4814);
or U6760 (N_6760,N_3538,N_3386);
nor U6761 (N_6761,N_3249,N_5406);
or U6762 (N_6762,N_5131,N_3839);
or U6763 (N_6763,N_4865,N_4320);
or U6764 (N_6764,N_5002,N_4452);
nor U6765 (N_6765,N_5790,N_4428);
and U6766 (N_6766,N_4028,N_5963);
nand U6767 (N_6767,N_3907,N_4266);
nand U6768 (N_6768,N_4478,N_4772);
nor U6769 (N_6769,N_5222,N_4115);
xnor U6770 (N_6770,N_3698,N_5219);
or U6771 (N_6771,N_5635,N_4670);
nor U6772 (N_6772,N_4420,N_3785);
or U6773 (N_6773,N_4625,N_4737);
nor U6774 (N_6774,N_5164,N_4927);
nand U6775 (N_6775,N_5854,N_5668);
nor U6776 (N_6776,N_3712,N_4831);
or U6777 (N_6777,N_3523,N_3605);
nor U6778 (N_6778,N_5525,N_5565);
nand U6779 (N_6779,N_4580,N_3184);
nand U6780 (N_6780,N_4198,N_5719);
and U6781 (N_6781,N_5903,N_5865);
nor U6782 (N_6782,N_4792,N_3186);
and U6783 (N_6783,N_5636,N_5174);
and U6784 (N_6784,N_4691,N_4802);
nand U6785 (N_6785,N_3747,N_3417);
xor U6786 (N_6786,N_4754,N_4953);
and U6787 (N_6787,N_3861,N_4746);
or U6788 (N_6788,N_5642,N_4957);
and U6789 (N_6789,N_3476,N_5624);
and U6790 (N_6790,N_3259,N_5148);
and U6791 (N_6791,N_3625,N_3295);
xnor U6792 (N_6792,N_4249,N_4366);
or U6793 (N_6793,N_4261,N_3595);
and U6794 (N_6794,N_3680,N_3947);
nand U6795 (N_6795,N_3255,N_4384);
nand U6796 (N_6796,N_3661,N_5462);
or U6797 (N_6797,N_3921,N_4243);
or U6798 (N_6798,N_5549,N_5493);
nand U6799 (N_6799,N_4271,N_4997);
nor U6800 (N_6800,N_4212,N_5230);
and U6801 (N_6801,N_4800,N_5887);
nor U6802 (N_6802,N_4718,N_3504);
or U6803 (N_6803,N_5670,N_3829);
nor U6804 (N_6804,N_4508,N_4713);
and U6805 (N_6805,N_4664,N_3753);
nand U6806 (N_6806,N_3521,N_5244);
and U6807 (N_6807,N_5369,N_5820);
and U6808 (N_6808,N_5847,N_3010);
nand U6809 (N_6809,N_5578,N_5382);
nor U6810 (N_6810,N_3180,N_5001);
and U6811 (N_6811,N_5713,N_3096);
nand U6812 (N_6812,N_4447,N_4906);
nand U6813 (N_6813,N_5559,N_5107);
nor U6814 (N_6814,N_3254,N_4848);
and U6815 (N_6815,N_5654,N_5322);
or U6816 (N_6816,N_4553,N_3788);
and U6817 (N_6817,N_3211,N_3235);
and U6818 (N_6818,N_5245,N_5889);
nand U6819 (N_6819,N_4075,N_5631);
and U6820 (N_6820,N_4272,N_4991);
and U6821 (N_6821,N_3893,N_3125);
nand U6822 (N_6822,N_5058,N_3596);
nor U6823 (N_6823,N_5416,N_5132);
and U6824 (N_6824,N_5028,N_3998);
nand U6825 (N_6825,N_4316,N_4615);
nand U6826 (N_6826,N_4610,N_3162);
nor U6827 (N_6827,N_3099,N_3505);
nor U6828 (N_6828,N_3149,N_4884);
nor U6829 (N_6829,N_4099,N_4896);
and U6830 (N_6830,N_3582,N_4094);
or U6831 (N_6831,N_4311,N_3776);
nor U6832 (N_6832,N_4917,N_5036);
nor U6833 (N_6833,N_4589,N_3205);
or U6834 (N_6834,N_3361,N_5821);
nand U6835 (N_6835,N_5289,N_5976);
nor U6836 (N_6836,N_4379,N_3847);
nor U6837 (N_6837,N_5895,N_3409);
and U6838 (N_6838,N_5204,N_5898);
and U6839 (N_6839,N_4996,N_5788);
nor U6840 (N_6840,N_5688,N_5103);
and U6841 (N_6841,N_3855,N_5195);
nand U6842 (N_6842,N_5084,N_4919);
nor U6843 (N_6843,N_3512,N_5022);
nor U6844 (N_6844,N_3826,N_5671);
nand U6845 (N_6845,N_3735,N_4757);
or U6846 (N_6846,N_5512,N_3087);
nor U6847 (N_6847,N_3374,N_4304);
nand U6848 (N_6848,N_5266,N_4002);
nand U6849 (N_6849,N_4551,N_4586);
nand U6850 (N_6850,N_4990,N_3620);
nor U6851 (N_6851,N_3530,N_3767);
and U6852 (N_6852,N_4547,N_5734);
nor U6853 (N_6853,N_4867,N_5556);
nor U6854 (N_6854,N_4162,N_5118);
nor U6855 (N_6855,N_3378,N_3130);
nor U6856 (N_6856,N_4491,N_4267);
or U6857 (N_6857,N_4345,N_5823);
nand U6858 (N_6858,N_3533,N_5207);
nand U6859 (N_6859,N_4348,N_4268);
or U6860 (N_6860,N_3214,N_4680);
and U6861 (N_6861,N_4776,N_5398);
nor U6862 (N_6862,N_4915,N_4790);
and U6863 (N_6863,N_5972,N_5552);
nor U6864 (N_6864,N_3682,N_3643);
or U6865 (N_6865,N_3560,N_5498);
nand U6866 (N_6866,N_5015,N_4401);
nor U6867 (N_6867,N_3163,N_5160);
and U6868 (N_6868,N_3970,N_3757);
nor U6869 (N_6869,N_4963,N_4518);
or U6870 (N_6870,N_5997,N_4001);
nand U6871 (N_6871,N_4623,N_4750);
and U6872 (N_6872,N_4987,N_4448);
nand U6873 (N_6873,N_3021,N_3270);
nor U6874 (N_6874,N_4076,N_3275);
nor U6875 (N_6875,N_4326,N_4004);
nor U6876 (N_6876,N_3158,N_3731);
nor U6877 (N_6877,N_3705,N_4883);
and U6878 (N_6878,N_5259,N_5454);
nand U6879 (N_6879,N_5479,N_4494);
and U6880 (N_6880,N_3571,N_5042);
or U6881 (N_6881,N_3734,N_4357);
and U6882 (N_6882,N_4131,N_4264);
and U6883 (N_6883,N_4910,N_5476);
nor U6884 (N_6884,N_5780,N_4537);
and U6885 (N_6885,N_4793,N_3090);
nand U6886 (N_6886,N_4375,N_3931);
or U6887 (N_6887,N_4862,N_5843);
nor U6888 (N_6888,N_5666,N_5017);
or U6889 (N_6889,N_4358,N_4522);
nor U6890 (N_6890,N_3929,N_3068);
or U6891 (N_6891,N_3168,N_4648);
nand U6892 (N_6892,N_4450,N_5075);
nor U6893 (N_6893,N_5240,N_4245);
nand U6894 (N_6894,N_4689,N_5530);
or U6895 (N_6895,N_3487,N_4897);
nor U6896 (N_6896,N_4923,N_4582);
nor U6897 (N_6897,N_4918,N_3003);
and U6898 (N_6898,N_4137,N_5133);
and U6899 (N_6899,N_3200,N_5474);
or U6900 (N_6900,N_3511,N_3029);
xnor U6901 (N_6901,N_3976,N_3304);
nand U6902 (N_6902,N_3196,N_4302);
nand U6903 (N_6903,N_5562,N_4985);
nand U6904 (N_6904,N_5777,N_4331);
nor U6905 (N_6905,N_3801,N_3510);
nor U6906 (N_6906,N_3252,N_5283);
nand U6907 (N_6907,N_3407,N_4647);
and U6908 (N_6908,N_5659,N_3674);
xor U6909 (N_6909,N_5083,N_4146);
nand U6910 (N_6910,N_5899,N_5262);
nand U6911 (N_6911,N_4600,N_3413);
and U6912 (N_6912,N_4124,N_4584);
nand U6913 (N_6913,N_4799,N_4217);
or U6914 (N_6914,N_5395,N_4712);
or U6915 (N_6915,N_4102,N_3351);
and U6916 (N_6916,N_4577,N_5686);
nand U6917 (N_6917,N_5486,N_3841);
nor U6918 (N_6918,N_3598,N_5345);
or U6919 (N_6919,N_4731,N_3696);
nor U6920 (N_6920,N_4810,N_5866);
and U6921 (N_6921,N_5983,N_5280);
or U6922 (N_6922,N_4988,N_3658);
nand U6923 (N_6923,N_4804,N_3828);
nand U6924 (N_6924,N_3412,N_5952);
or U6925 (N_6925,N_5072,N_3851);
or U6926 (N_6926,N_5881,N_3892);
and U6927 (N_6927,N_5145,N_5630);
and U6928 (N_6928,N_5628,N_5662);
and U6929 (N_6929,N_4616,N_3238);
nor U6930 (N_6930,N_3827,N_3671);
or U6931 (N_6931,N_5349,N_3983);
or U6932 (N_6932,N_3306,N_4163);
nor U6933 (N_6933,N_3787,N_4436);
and U6934 (N_6934,N_4860,N_5640);
or U6935 (N_6935,N_5940,N_4405);
nor U6936 (N_6936,N_5561,N_5316);
nand U6937 (N_6937,N_5242,N_4486);
and U6938 (N_6938,N_4698,N_5029);
or U6939 (N_6939,N_4467,N_5817);
nand U6940 (N_6940,N_5527,N_3318);
and U6941 (N_6941,N_3392,N_3942);
and U6942 (N_6942,N_5908,N_3737);
nand U6943 (N_6943,N_3502,N_3751);
nand U6944 (N_6944,N_4453,N_5078);
nor U6945 (N_6945,N_5430,N_5672);
or U6946 (N_6946,N_3279,N_5013);
and U6947 (N_6947,N_5644,N_3223);
nor U6948 (N_6948,N_4788,N_4079);
nor U6949 (N_6949,N_3032,N_3468);
nor U6950 (N_6950,N_5080,N_4047);
or U6951 (N_6951,N_5756,N_4481);
and U6952 (N_6952,N_4209,N_5142);
nand U6953 (N_6953,N_4642,N_3165);
or U6954 (N_6954,N_4341,N_5661);
or U6955 (N_6955,N_4073,N_4214);
or U6956 (N_6956,N_5753,N_5141);
and U6957 (N_6957,N_3678,N_4598);
and U6958 (N_6958,N_4710,N_3150);
or U6959 (N_6959,N_3587,N_4548);
nand U6960 (N_6960,N_4606,N_5569);
nand U6961 (N_6961,N_5864,N_4559);
and U6962 (N_6962,N_3089,N_4678);
nand U6963 (N_6963,N_4666,N_4829);
and U6964 (N_6964,N_3220,N_3556);
and U6965 (N_6965,N_5622,N_4247);
and U6966 (N_6966,N_5653,N_5157);
nand U6967 (N_6967,N_4445,N_3740);
or U6968 (N_6968,N_4558,N_5508);
nand U6969 (N_6969,N_4003,N_5977);
or U6970 (N_6970,N_5201,N_4171);
and U6971 (N_6971,N_4008,N_3081);
nor U6972 (N_6972,N_5799,N_4395);
or U6973 (N_6973,N_4026,N_4768);
and U6974 (N_6974,N_5269,N_4308);
nor U6975 (N_6975,N_5307,N_5923);
and U6976 (N_6976,N_3118,N_3079);
or U6977 (N_6977,N_4234,N_3450);
nor U6978 (N_6978,N_4089,N_4225);
or U6979 (N_6979,N_3507,N_5419);
xnor U6980 (N_6980,N_3462,N_4983);
and U6981 (N_6981,N_4040,N_5064);
nand U6982 (N_6982,N_5059,N_5344);
xor U6983 (N_6983,N_3552,N_3599);
nand U6984 (N_6984,N_4116,N_3469);
nand U6985 (N_6985,N_3145,N_3248);
and U6986 (N_6986,N_4262,N_5434);
or U6987 (N_6987,N_3750,N_5279);
and U6988 (N_6988,N_3199,N_3320);
and U6989 (N_6989,N_5669,N_5282);
nor U6990 (N_6990,N_4151,N_4866);
and U6991 (N_6991,N_3005,N_4546);
or U6992 (N_6992,N_3761,N_3053);
nor U6993 (N_6993,N_5303,N_3442);
and U6994 (N_6994,N_3030,N_4931);
and U6995 (N_6995,N_5600,N_5510);
or U6996 (N_6996,N_5927,N_4213);
nand U6997 (N_6997,N_4172,N_3094);
nor U6998 (N_6998,N_4178,N_5581);
and U6999 (N_6999,N_4890,N_5492);
nor U7000 (N_7000,N_3002,N_3765);
nand U7001 (N_7001,N_4461,N_4715);
nor U7002 (N_7002,N_4811,N_3419);
nor U7003 (N_7003,N_5473,N_3890);
or U7004 (N_7004,N_4676,N_3232);
and U7005 (N_7005,N_5189,N_3095);
or U7006 (N_7006,N_4673,N_5907);
nor U7007 (N_7007,N_4105,N_5371);
nor U7008 (N_7008,N_4435,N_3768);
or U7009 (N_7009,N_4355,N_3692);
or U7010 (N_7010,N_4032,N_3608);
and U7011 (N_7011,N_3225,N_3986);
nor U7012 (N_7012,N_5006,N_5265);
nand U7013 (N_7013,N_3837,N_5301);
xnor U7014 (N_7014,N_3298,N_5597);
and U7015 (N_7015,N_4301,N_5766);
or U7016 (N_7016,N_3363,N_5859);
and U7017 (N_7017,N_5708,N_4735);
or U7018 (N_7018,N_5239,N_3640);
nand U7019 (N_7019,N_5153,N_3884);
nand U7020 (N_7020,N_5948,N_3990);
and U7021 (N_7021,N_3326,N_3805);
and U7022 (N_7022,N_3950,N_3638);
nor U7023 (N_7023,N_5323,N_3324);
nor U7024 (N_7024,N_4332,N_4456);
and U7025 (N_7025,N_4761,N_3563);
xnor U7026 (N_7026,N_4418,N_5191);
and U7027 (N_7027,N_4011,N_5256);
nor U7028 (N_7028,N_5104,N_3185);
or U7029 (N_7029,N_5408,N_4583);
or U7030 (N_7030,N_3432,N_3527);
nand U7031 (N_7031,N_3485,N_4596);
and U7032 (N_7032,N_4727,N_4426);
nand U7033 (N_7033,N_3434,N_5807);
nor U7034 (N_7034,N_3977,N_3811);
and U7035 (N_7035,N_3321,N_5034);
and U7036 (N_7036,N_4892,N_4145);
nor U7037 (N_7037,N_5452,N_4431);
nor U7038 (N_7038,N_3651,N_4520);
nand U7039 (N_7039,N_5522,N_3291);
nor U7040 (N_7040,N_4201,N_4468);
or U7041 (N_7041,N_5027,N_5814);
or U7042 (N_7042,N_4903,N_4898);
nand U7043 (N_7043,N_5458,N_5804);
nor U7044 (N_7044,N_3939,N_4783);
or U7045 (N_7045,N_3315,N_5542);
nor U7046 (N_7046,N_4823,N_3819);
or U7047 (N_7047,N_5288,N_5951);
nand U7048 (N_7048,N_5079,N_4879);
nor U7049 (N_7049,N_5162,N_4053);
and U7050 (N_7050,N_5333,N_5151);
nand U7051 (N_7051,N_5547,N_5511);
or U7052 (N_7052,N_4578,N_5475);
nand U7053 (N_7053,N_4557,N_5073);
nand U7054 (N_7054,N_3649,N_5538);
or U7055 (N_7055,N_3441,N_4966);
and U7056 (N_7056,N_4513,N_5067);
and U7057 (N_7057,N_5679,N_3714);
nand U7058 (N_7058,N_3964,N_3183);
and U7059 (N_7059,N_3154,N_4489);
nand U7060 (N_7060,N_3982,N_3909);
or U7061 (N_7061,N_3726,N_4180);
or U7062 (N_7062,N_3062,N_4753);
or U7063 (N_7063,N_3821,N_3914);
xor U7064 (N_7064,N_5485,N_5436);
or U7065 (N_7065,N_3569,N_5656);
nand U7066 (N_7066,N_5724,N_3039);
or U7067 (N_7067,N_4340,N_5008);
nor U7068 (N_7068,N_5268,N_3856);
xnor U7069 (N_7069,N_5443,N_3619);
and U7070 (N_7070,N_4880,N_3234);
and U7071 (N_7071,N_4439,N_3927);
or U7072 (N_7072,N_3902,N_5205);
or U7073 (N_7073,N_3957,N_5198);
and U7074 (N_7074,N_5488,N_3054);
nor U7075 (N_7075,N_3844,N_4036);
xor U7076 (N_7076,N_3403,N_5627);
or U7077 (N_7077,N_4574,N_4538);
nand U7078 (N_7078,N_3281,N_3330);
nand U7079 (N_7079,N_5596,N_4020);
or U7080 (N_7080,N_3896,N_3930);
nor U7081 (N_7081,N_4882,N_5375);
xor U7082 (N_7082,N_3987,N_5300);
or U7083 (N_7083,N_5137,N_3157);
and U7084 (N_7084,N_5377,N_4051);
or U7085 (N_7085,N_4299,N_4044);
or U7086 (N_7086,N_3041,N_3762);
nor U7087 (N_7087,N_4160,N_5975);
nand U7088 (N_7088,N_5968,N_4644);
nand U7089 (N_7089,N_3729,N_3799);
nor U7090 (N_7090,N_4128,N_4328);
or U7091 (N_7091,N_3853,N_4374);
nor U7092 (N_7092,N_4962,N_4462);
nand U7093 (N_7093,N_3725,N_3049);
xor U7094 (N_7094,N_3858,N_3656);
or U7095 (N_7095,N_5114,N_3944);
nor U7096 (N_7096,N_3400,N_5536);
nor U7097 (N_7097,N_4241,N_3464);
nand U7098 (N_7098,N_5551,N_4451);
and U7099 (N_7099,N_4794,N_3686);
nor U7100 (N_7100,N_4760,N_5579);
and U7101 (N_7101,N_3804,N_3340);
and U7102 (N_7102,N_3659,N_4072);
nor U7103 (N_7103,N_3209,N_5128);
and U7104 (N_7104,N_5616,N_5646);
and U7105 (N_7105,N_3491,N_3648);
xor U7106 (N_7106,N_4021,N_3535);
and U7107 (N_7107,N_4175,N_5768);
nor U7108 (N_7108,N_4981,N_3969);
nor U7109 (N_7109,N_5226,N_5109);
and U7110 (N_7110,N_3577,N_4833);
nand U7111 (N_7111,N_4922,N_5884);
or U7112 (N_7112,N_3436,N_4226);
or U7113 (N_7113,N_5081,N_4080);
or U7114 (N_7114,N_4828,N_4838);
and U7115 (N_7115,N_5049,N_3639);
or U7116 (N_7116,N_3018,N_3483);
nor U7117 (N_7117,N_5313,N_3117);
nand U7118 (N_7118,N_5356,N_3119);
or U7119 (N_7119,N_3262,N_5698);
nand U7120 (N_7120,N_3966,N_5971);
nand U7121 (N_7121,N_5098,N_5910);
or U7122 (N_7122,N_4714,N_4652);
nor U7123 (N_7123,N_3809,N_4779);
nand U7124 (N_7124,N_5225,N_4933);
and U7125 (N_7125,N_3459,N_4362);
nand U7126 (N_7126,N_3934,N_3883);
or U7127 (N_7127,N_4965,N_5586);
or U7128 (N_7128,N_4417,N_5813);
or U7129 (N_7129,N_5681,N_3557);
and U7130 (N_7130,N_3012,N_4233);
and U7131 (N_7131,N_3410,N_4108);
and U7132 (N_7132,N_3257,N_4240);
nor U7133 (N_7133,N_5736,N_3006);
or U7134 (N_7134,N_3022,N_3271);
nor U7135 (N_7135,N_5161,N_5763);
and U7136 (N_7136,N_3343,N_5102);
nor U7137 (N_7137,N_5425,N_5637);
nor U7138 (N_7138,N_4278,N_5089);
or U7139 (N_7139,N_4844,N_3664);
nor U7140 (N_7140,N_3292,N_5163);
or U7141 (N_7141,N_4199,N_5520);
nand U7142 (N_7142,N_5643,N_3398);
or U7143 (N_7143,N_3544,N_4191);
nor U7144 (N_7144,N_3080,N_3965);
and U7145 (N_7145,N_4136,N_4994);
or U7146 (N_7146,N_5754,N_3498);
or U7147 (N_7147,N_5214,N_5144);
and U7148 (N_7148,N_4292,N_3439);
nor U7149 (N_7149,N_3448,N_4229);
or U7150 (N_7150,N_4534,N_3016);
and U7151 (N_7151,N_4628,N_5855);
nor U7152 (N_7152,N_3025,N_3380);
and U7153 (N_7153,N_4542,N_3414);
and U7154 (N_7154,N_5878,N_3009);
or U7155 (N_7155,N_4764,N_4029);
nand U7156 (N_7156,N_3377,N_5749);
and U7157 (N_7157,N_4973,N_4863);
and U7158 (N_7158,N_4083,N_4280);
or U7159 (N_7159,N_3910,N_5451);
or U7160 (N_7160,N_5233,N_4544);
nor U7161 (N_7161,N_4573,N_4027);
nor U7162 (N_7162,N_3917,N_5297);
or U7163 (N_7163,N_3739,N_5988);
nor U7164 (N_7164,N_3276,N_3775);
and U7165 (N_7165,N_5789,N_3293);
or U7166 (N_7166,N_4495,N_4951);
and U7167 (N_7167,N_4569,N_3820);
nor U7168 (N_7168,N_5796,N_5185);
nor U7169 (N_7169,N_3882,N_3975);
nand U7170 (N_7170,N_5610,N_4899);
or U7171 (N_7171,N_5825,N_5094);
or U7172 (N_7172,N_5582,N_5759);
or U7173 (N_7173,N_4176,N_4528);
nor U7174 (N_7174,N_3774,N_3865);
nand U7175 (N_7175,N_5747,N_4018);
nor U7176 (N_7176,N_4457,N_3794);
and U7177 (N_7177,N_3580,N_4174);
and U7178 (N_7178,N_4399,N_4667);
and U7179 (N_7179,N_5005,N_5446);
nand U7180 (N_7180,N_5496,N_4763);
nor U7181 (N_7181,N_4370,N_4575);
nor U7182 (N_7182,N_3222,N_3013);
nor U7183 (N_7183,N_4636,N_4007);
and U7184 (N_7184,N_3120,N_5781);
nand U7185 (N_7185,N_3553,N_3231);
and U7186 (N_7186,N_5505,N_5695);
and U7187 (N_7187,N_4252,N_3179);
or U7188 (N_7188,N_3362,N_4591);
or U7189 (N_7189,N_4100,N_5095);
nand U7190 (N_7190,N_3139,N_5937);
nor U7191 (N_7191,N_4303,N_5853);
and U7192 (N_7192,N_3508,N_3806);
nand U7193 (N_7193,N_3722,N_4157);
nor U7194 (N_7194,N_3642,N_5461);
or U7195 (N_7195,N_3905,N_4458);
and U7196 (N_7196,N_5757,N_5209);
nand U7197 (N_7197,N_5173,N_3667);
nor U7198 (N_7198,N_4069,N_3610);
nor U7199 (N_7199,N_5942,N_4106);
nor U7200 (N_7200,N_4808,N_3838);
nand U7201 (N_7201,N_4052,N_4454);
and U7202 (N_7202,N_5954,N_3627);
nor U7203 (N_7203,N_3136,N_3558);
or U7204 (N_7204,N_3515,N_5564);
nand U7205 (N_7205,N_5082,N_3350);
and U7206 (N_7206,N_5812,N_3300);
nor U7207 (N_7207,N_5235,N_4487);
xnor U7208 (N_7208,N_5350,N_4595);
nor U7209 (N_7209,N_4306,N_3027);
nor U7210 (N_7210,N_5517,N_5607);
or U7211 (N_7211,N_4813,N_5947);
nor U7212 (N_7212,N_5829,N_5263);
nand U7213 (N_7213,N_3190,N_4381);
nor U7214 (N_7214,N_3562,N_5047);
nand U7215 (N_7215,N_5495,N_4639);
nor U7216 (N_7216,N_3848,N_4490);
or U7217 (N_7217,N_4154,N_4156);
nor U7218 (N_7218,N_5801,N_4187);
or U7219 (N_7219,N_3915,N_5682);
or U7220 (N_7220,N_3548,N_3427);
nor U7221 (N_7221,N_5053,N_3098);
nand U7222 (N_7222,N_3872,N_5155);
nor U7223 (N_7223,N_4622,N_3606);
nor U7224 (N_7224,N_4190,N_4858);
and U7225 (N_7225,N_3052,N_3488);
or U7226 (N_7226,N_4139,N_5989);
nand U7227 (N_7227,N_3466,N_5237);
or U7228 (N_7228,N_3877,N_4822);
and U7229 (N_7229,N_4279,N_3926);
nor U7230 (N_7230,N_3342,N_5845);
nand U7231 (N_7231,N_4873,N_3823);
nor U7232 (N_7232,N_5293,N_3115);
nor U7233 (N_7233,N_5851,N_3040);
nand U7234 (N_7234,N_3579,N_4631);
or U7235 (N_7235,N_3272,N_4669);
nand U7236 (N_7236,N_5943,N_5284);
nand U7237 (N_7237,N_3334,N_3866);
or U7238 (N_7238,N_4275,N_4565);
nand U7239 (N_7239,N_5400,N_4806);
nor U7240 (N_7240,N_3629,N_3347);
nand U7241 (N_7241,N_3668,N_5867);
nand U7242 (N_7242,N_5818,N_4315);
or U7243 (N_7243,N_3995,N_4203);
and U7244 (N_7244,N_3550,N_4274);
nor U7245 (N_7245,N_3399,N_4765);
nand U7246 (N_7246,N_3946,N_4470);
and U7247 (N_7247,N_4054,N_3824);
xor U7248 (N_7248,N_4351,N_5928);
and U7249 (N_7249,N_5601,N_5808);
nor U7250 (N_7250,N_5418,N_5490);
nand U7251 (N_7251,N_5810,N_4424);
nor U7252 (N_7252,N_4077,N_4861);
nor U7253 (N_7253,N_4995,N_3240);
nor U7254 (N_7254,N_3109,N_4721);
and U7255 (N_7255,N_3547,N_4013);
nand U7256 (N_7256,N_5315,N_3881);
nand U7257 (N_7257,N_5175,N_4758);
and U7258 (N_7258,N_4782,N_4699);
nor U7259 (N_7259,N_4830,N_3303);
or U7260 (N_7260,N_5409,N_5540);
nand U7261 (N_7261,N_3868,N_3011);
nand U7262 (N_7262,N_4427,N_5108);
or U7263 (N_7263,N_4133,N_4469);
or U7264 (N_7264,N_3688,N_3308);
nand U7265 (N_7265,N_5839,N_3496);
or U7266 (N_7266,N_3075,N_3989);
nor U7267 (N_7267,N_3290,N_4391);
or U7268 (N_7268,N_3106,N_3666);
and U7269 (N_7269,N_3151,N_3888);
and U7270 (N_7270,N_5929,N_3898);
or U7271 (N_7271,N_5327,N_4166);
nand U7272 (N_7272,N_4523,N_5838);
and U7273 (N_7273,N_3268,N_5140);
and U7274 (N_7274,N_5870,N_4419);
and U7275 (N_7275,N_4144,N_3670);
nor U7276 (N_7276,N_5822,N_3319);
nor U7277 (N_7277,N_3024,N_5879);
nand U7278 (N_7278,N_5105,N_3055);
and U7279 (N_7279,N_3129,N_4876);
and U7280 (N_7280,N_4432,N_4186);
nand U7281 (N_7281,N_5609,N_5676);
nor U7282 (N_7282,N_3213,N_5791);
nand U7283 (N_7283,N_4945,N_5383);
nand U7284 (N_7284,N_5523,N_4253);
and U7285 (N_7285,N_3830,N_4941);
xor U7286 (N_7286,N_5709,N_4359);
and U7287 (N_7287,N_4300,N_3317);
nand U7288 (N_7288,N_4739,N_3706);
nand U7289 (N_7289,N_3078,N_5365);
nand U7290 (N_7290,N_4433,N_3144);
nor U7291 (N_7291,N_4471,N_3379);
and U7292 (N_7292,N_4161,N_5170);
nand U7293 (N_7293,N_4853,N_4231);
and U7294 (N_7294,N_3336,N_3134);
and U7295 (N_7295,N_4709,N_5846);
nor U7296 (N_7296,N_5248,N_3189);
nor U7297 (N_7297,N_4656,N_5007);
nor U7298 (N_7298,N_5050,N_3173);
and U7299 (N_7299,N_4891,N_3880);
and U7300 (N_7300,N_4971,N_3140);
nand U7301 (N_7301,N_4535,N_3978);
nor U7302 (N_7302,N_4711,N_5320);
and U7303 (N_7303,N_5294,N_5802);
or U7304 (N_7304,N_5069,N_3967);
and U7305 (N_7305,N_5393,N_4908);
and U7306 (N_7306,N_3438,N_4284);
and U7307 (N_7307,N_4888,N_4441);
and U7308 (N_7308,N_3433,N_5481);
nand U7309 (N_7309,N_5773,N_5384);
nand U7310 (N_7310,N_4576,N_5464);
or U7311 (N_7311,N_5785,N_3716);
or U7312 (N_7312,N_4207,N_4843);
and U7313 (N_7313,N_3375,N_4755);
or U7314 (N_7314,N_5960,N_3167);
or U7315 (N_7315,N_5432,N_3266);
xor U7316 (N_7316,N_3345,N_3367);
nand U7317 (N_7317,N_3551,N_4093);
nor U7318 (N_7318,N_5340,N_5873);
nand U7319 (N_7319,N_5039,N_5767);
and U7320 (N_7320,N_4961,N_3107);
or U7321 (N_7321,N_3772,N_3253);
and U7322 (N_7322,N_3842,N_4377);
nand U7323 (N_7323,N_5718,N_5254);
and U7324 (N_7324,N_5693,N_4820);
nor U7325 (N_7325,N_4392,N_4986);
nand U7326 (N_7326,N_5593,N_5583);
nor U7327 (N_7327,N_3924,N_3174);
and U7328 (N_7328,N_4651,N_3867);
nor U7329 (N_7329,N_3759,N_4129);
nand U7330 (N_7330,N_4614,N_5023);
nor U7331 (N_7331,N_5727,N_5172);
nor U7332 (N_7332,N_5834,N_5585);
nand U7333 (N_7333,N_3493,N_3456);
xor U7334 (N_7334,N_4952,N_4977);
nand U7335 (N_7335,N_3333,N_3733);
nor U7336 (N_7336,N_4194,N_5779);
and U7337 (N_7337,N_5362,N_4159);
nand U7338 (N_7338,N_4354,N_5318);
nor U7339 (N_7339,N_3202,N_3985);
nand U7340 (N_7340,N_3912,N_3036);
nor U7341 (N_7341,N_4338,N_3261);
nand U7342 (N_7342,N_3730,N_3216);
nand U7343 (N_7343,N_4286,N_5612);
and U7344 (N_7344,N_5956,N_5706);
or U7345 (N_7345,N_4407,N_3114);
nor U7346 (N_7346,N_4751,N_3474);
nor U7347 (N_7347,N_3711,N_4221);
or U7348 (N_7348,N_5332,N_4579);
nor U7349 (N_7349,N_5798,N_5187);
xor U7350 (N_7350,N_3630,N_3955);
or U7351 (N_7351,N_3719,N_5358);
nand U7352 (N_7352,N_3092,N_4488);
xor U7353 (N_7353,N_3445,N_5373);
nor U7354 (N_7354,N_4111,N_3777);
or U7355 (N_7355,N_5123,N_5509);
nor U7356 (N_7356,N_4307,N_3443);
or U7357 (N_7357,N_4035,N_4373);
nor U7358 (N_7358,N_5171,N_4437);
nand U7359 (N_7359,N_5361,N_3953);
nor U7360 (N_7360,N_3497,N_5267);
and U7361 (N_7361,N_4703,N_4095);
and U7362 (N_7362,N_3928,N_4687);
and U7363 (N_7363,N_5063,N_4878);
and U7364 (N_7364,N_5856,N_3057);
nand U7365 (N_7365,N_4322,N_3704);
xor U7366 (N_7366,N_4177,N_4215);
nand U7367 (N_7367,N_3401,N_5580);
nor U7368 (N_7368,N_3609,N_5210);
nor U7369 (N_7369,N_3600,N_5603);
and U7370 (N_7370,N_4189,N_5830);
nand U7371 (N_7371,N_4958,N_4695);
nor U7372 (N_7372,N_3182,N_5200);
or U7373 (N_7373,N_5085,N_5758);
and U7374 (N_7374,N_3256,N_4525);
and U7375 (N_7375,N_4346,N_5699);
xor U7376 (N_7376,N_5033,N_3545);
nor U7377 (N_7377,N_3941,N_3962);
nor U7378 (N_7378,N_5014,N_3918);
or U7379 (N_7379,N_4141,N_5179);
and U7380 (N_7380,N_5626,N_3709);
or U7381 (N_7381,N_5639,N_5584);
nand U7382 (N_7382,N_5329,N_4383);
nor U7383 (N_7383,N_3831,N_3472);
or U7384 (N_7384,N_3663,N_5712);
nor U7385 (N_7385,N_5573,N_3607);
and U7386 (N_7386,N_3758,N_4749);
and U7387 (N_7387,N_4724,N_4181);
nor U7388 (N_7388,N_4516,N_3532);
nor U7389 (N_7389,N_3457,N_4607);
and U7390 (N_7390,N_3420,N_3091);
and U7391 (N_7391,N_5221,N_4774);
nand U7392 (N_7392,N_4510,N_3465);
or U7393 (N_7393,N_3482,N_5236);
or U7394 (N_7394,N_3899,N_5531);
nand U7395 (N_7395,N_3348,N_4655);
and U7396 (N_7396,N_3632,N_4617);
nand U7397 (N_7397,N_4745,N_5367);
or U7398 (N_7398,N_3871,N_4543);
nor U7399 (N_7399,N_4887,N_5955);
and U7400 (N_7400,N_4905,N_5287);
xnor U7401 (N_7401,N_5837,N_5526);
or U7402 (N_7402,N_4010,N_3192);
and U7403 (N_7403,N_3952,N_5649);
xor U7404 (N_7404,N_3463,N_3486);
and U7405 (N_7405,N_3391,N_4288);
nor U7406 (N_7406,N_3500,N_4940);
nand U7407 (N_7407,N_5991,N_5902);
or U7408 (N_7408,N_4270,N_4255);
nor U7409 (N_7409,N_4934,N_4556);
nand U7410 (N_7410,N_4771,N_3430);
nor U7411 (N_7411,N_3122,N_5312);
and U7412 (N_7412,N_3389,N_5188);
nand U7413 (N_7413,N_5704,N_5863);
and U7414 (N_7414,N_5438,N_3786);
or U7415 (N_7415,N_5380,N_4629);
and U7416 (N_7416,N_3460,N_3063);
nand U7417 (N_7417,N_5769,N_4533);
or U7418 (N_7418,N_5275,N_5270);
nor U7419 (N_7419,N_5555,N_4726);
or U7420 (N_7420,N_5449,N_4196);
nand U7421 (N_7421,N_4716,N_3922);
or U7422 (N_7422,N_5497,N_3617);
nor U7423 (N_7423,N_4034,N_4943);
nand U7424 (N_7424,N_4260,N_3581);
and U7425 (N_7425,N_3652,N_5134);
or U7426 (N_7426,N_5314,N_4019);
nand U7427 (N_7427,N_3708,N_3701);
and U7428 (N_7428,N_4070,N_3370);
nor U7429 (N_7429,N_5877,N_4463);
xor U7430 (N_7430,N_3228,N_5335);
nor U7431 (N_7431,N_4924,N_5491);
xnor U7432 (N_7432,N_5882,N_5783);
xnor U7433 (N_7433,N_4868,N_4778);
and U7434 (N_7434,N_3195,N_4400);
nand U7435 (N_7435,N_5647,N_5359);
xnor U7436 (N_7436,N_3840,N_4665);
nand U7437 (N_7437,N_4722,N_3681);
nor U7438 (N_7438,N_3586,N_4038);
nor U7439 (N_7439,N_5680,N_4970);
nand U7440 (N_7440,N_5992,N_3754);
nor U7441 (N_7441,N_4501,N_4650);
and U7442 (N_7442,N_5999,N_3634);
nor U7443 (N_7443,N_4110,N_3499);
and U7444 (N_7444,N_5217,N_5445);
xnor U7445 (N_7445,N_5563,N_4082);
nor U7446 (N_7446,N_5611,N_5969);
and U7447 (N_7447,N_4706,N_4807);
xor U7448 (N_7448,N_3937,N_4852);
nand U7449 (N_7449,N_3072,N_3265);
nand U7450 (N_7450,N_5021,N_3886);
and U7451 (N_7451,N_5274,N_5762);
nand U7452 (N_7452,N_3764,N_3700);
nand U7453 (N_7453,N_5030,N_5494);
and U7454 (N_7454,N_3616,N_3088);
nand U7455 (N_7455,N_3803,N_4483);
and U7456 (N_7456,N_3479,N_5025);
and U7457 (N_7457,N_5705,N_4856);
and U7458 (N_7458,N_4540,N_3470);
and U7459 (N_7459,N_3578,N_5456);
nor U7460 (N_7460,N_3657,N_4202);
nand U7461 (N_7461,N_4455,N_5052);
and U7462 (N_7462,N_3635,N_3492);
and U7463 (N_7463,N_4394,N_3769);
nor U7464 (N_7464,N_4224,N_3471);
nand U7465 (N_7465,N_5167,N_5961);
nand U7466 (N_7466,N_5504,N_5457);
and U7467 (N_7467,N_4323,N_3015);
nand U7468 (N_7468,N_3583,N_5388);
nor U7469 (N_7469,N_4442,N_3968);
nor U7470 (N_7470,N_4025,N_4068);
nand U7471 (N_7471,N_5212,N_4638);
nand U7472 (N_7472,N_3559,N_5299);
xnor U7473 (N_7473,N_5883,N_4239);
and U7474 (N_7474,N_5620,N_5296);
and U7475 (N_7475,N_5097,N_4269);
nand U7476 (N_7476,N_4998,N_4045);
nand U7477 (N_7477,N_4318,N_4499);
and U7478 (N_7478,N_5459,N_5803);
and U7479 (N_7479,N_3679,N_5368);
xnor U7480 (N_7480,N_4926,N_4422);
nand U7481 (N_7481,N_3958,N_3278);
or U7482 (N_7482,N_5101,N_4423);
or U7483 (N_7483,N_3243,N_5794);
or U7484 (N_7484,N_5220,N_3790);
nor U7485 (N_7485,N_5506,N_4907);
and U7486 (N_7486,N_5469,N_4104);
nor U7487 (N_7487,N_5360,N_4937);
nor U7488 (N_7488,N_4446,N_5183);
and U7489 (N_7489,N_4612,N_3713);
and U7490 (N_7490,N_4969,N_3903);
nor U7491 (N_7491,N_5238,N_3845);
nand U7492 (N_7492,N_3355,N_5184);
nand U7493 (N_7493,N_4126,N_4048);
or U7494 (N_7494,N_5964,N_3307);
nor U7495 (N_7495,N_3447,N_4347);
and U7496 (N_7496,N_4319,N_4107);
nor U7497 (N_7497,N_4671,N_4385);
or U7498 (N_7498,N_3219,N_4227);
or U7499 (N_7499,N_4641,N_5374);
nor U7500 (N_7500,N_5118,N_5719);
xor U7501 (N_7501,N_5823,N_4254);
and U7502 (N_7502,N_4585,N_4574);
nand U7503 (N_7503,N_3365,N_4445);
and U7504 (N_7504,N_4041,N_4965);
or U7505 (N_7505,N_3173,N_4424);
and U7506 (N_7506,N_5259,N_4727);
and U7507 (N_7507,N_3582,N_5562);
nor U7508 (N_7508,N_3432,N_4374);
and U7509 (N_7509,N_3715,N_3909);
nand U7510 (N_7510,N_5169,N_5570);
nor U7511 (N_7511,N_3943,N_4223);
nand U7512 (N_7512,N_4954,N_3392);
or U7513 (N_7513,N_3791,N_4968);
and U7514 (N_7514,N_5007,N_4401);
and U7515 (N_7515,N_3482,N_4463);
or U7516 (N_7516,N_3832,N_4136);
nand U7517 (N_7517,N_5434,N_5593);
or U7518 (N_7518,N_4371,N_4953);
and U7519 (N_7519,N_3979,N_5565);
and U7520 (N_7520,N_3868,N_4563);
nand U7521 (N_7521,N_5726,N_5577);
or U7522 (N_7522,N_4144,N_3091);
nor U7523 (N_7523,N_3255,N_4453);
or U7524 (N_7524,N_5919,N_5612);
and U7525 (N_7525,N_5955,N_4641);
or U7526 (N_7526,N_3183,N_3062);
nor U7527 (N_7527,N_4440,N_4665);
nand U7528 (N_7528,N_3381,N_5664);
nand U7529 (N_7529,N_5208,N_3367);
and U7530 (N_7530,N_3812,N_5316);
nand U7531 (N_7531,N_3353,N_3352);
and U7532 (N_7532,N_3070,N_3390);
or U7533 (N_7533,N_3424,N_3644);
nand U7534 (N_7534,N_5461,N_3524);
or U7535 (N_7535,N_3302,N_4310);
nand U7536 (N_7536,N_5750,N_3289);
and U7537 (N_7537,N_5598,N_5195);
nor U7538 (N_7538,N_3793,N_4822);
and U7539 (N_7539,N_5688,N_5642);
or U7540 (N_7540,N_4618,N_3883);
and U7541 (N_7541,N_3173,N_3597);
and U7542 (N_7542,N_3706,N_5684);
nor U7543 (N_7543,N_4491,N_5118);
nor U7544 (N_7544,N_5950,N_3382);
nand U7545 (N_7545,N_4035,N_4536);
and U7546 (N_7546,N_4012,N_3760);
nand U7547 (N_7547,N_5761,N_5978);
nand U7548 (N_7548,N_4931,N_4426);
and U7549 (N_7549,N_3192,N_5570);
nor U7550 (N_7550,N_3726,N_3735);
nand U7551 (N_7551,N_4042,N_5746);
or U7552 (N_7552,N_4772,N_4647);
nor U7553 (N_7553,N_3012,N_3842);
or U7554 (N_7554,N_4108,N_5187);
and U7555 (N_7555,N_4791,N_5040);
nor U7556 (N_7556,N_4651,N_3403);
nand U7557 (N_7557,N_4485,N_4241);
xnor U7558 (N_7558,N_5661,N_5031);
nor U7559 (N_7559,N_4257,N_5241);
nor U7560 (N_7560,N_4786,N_5451);
nor U7561 (N_7561,N_3431,N_5814);
nand U7562 (N_7562,N_4659,N_4903);
nor U7563 (N_7563,N_4261,N_4116);
nor U7564 (N_7564,N_3084,N_4144);
nor U7565 (N_7565,N_3512,N_3661);
or U7566 (N_7566,N_5868,N_5071);
nand U7567 (N_7567,N_4852,N_5425);
nand U7568 (N_7568,N_4129,N_5025);
and U7569 (N_7569,N_3462,N_5450);
nor U7570 (N_7570,N_5572,N_5916);
nand U7571 (N_7571,N_3273,N_4867);
xor U7572 (N_7572,N_4699,N_5490);
nand U7573 (N_7573,N_5658,N_3668);
nand U7574 (N_7574,N_5975,N_3400);
nor U7575 (N_7575,N_5362,N_5443);
nor U7576 (N_7576,N_4078,N_5595);
or U7577 (N_7577,N_3189,N_3618);
nand U7578 (N_7578,N_4771,N_3721);
and U7579 (N_7579,N_3794,N_4153);
nand U7580 (N_7580,N_4127,N_4693);
or U7581 (N_7581,N_4505,N_5387);
nand U7582 (N_7582,N_3035,N_3289);
or U7583 (N_7583,N_3193,N_3346);
nand U7584 (N_7584,N_5065,N_4654);
xnor U7585 (N_7585,N_3088,N_4168);
and U7586 (N_7586,N_5075,N_4037);
or U7587 (N_7587,N_4644,N_4656);
or U7588 (N_7588,N_3081,N_5105);
and U7589 (N_7589,N_4882,N_3664);
nor U7590 (N_7590,N_3649,N_4139);
nand U7591 (N_7591,N_5275,N_4123);
nand U7592 (N_7592,N_4006,N_3845);
nand U7593 (N_7593,N_5620,N_5692);
xnor U7594 (N_7594,N_5857,N_4597);
and U7595 (N_7595,N_5167,N_5422);
nand U7596 (N_7596,N_5338,N_3186);
and U7597 (N_7597,N_3215,N_5660);
nor U7598 (N_7598,N_4100,N_3976);
nor U7599 (N_7599,N_3160,N_3652);
nor U7600 (N_7600,N_4314,N_4337);
and U7601 (N_7601,N_5647,N_5692);
nor U7602 (N_7602,N_5667,N_4512);
or U7603 (N_7603,N_3350,N_4295);
and U7604 (N_7604,N_3448,N_4953);
or U7605 (N_7605,N_4325,N_4742);
and U7606 (N_7606,N_5328,N_4900);
or U7607 (N_7607,N_4374,N_3070);
or U7608 (N_7608,N_5672,N_3117);
or U7609 (N_7609,N_3762,N_4184);
or U7610 (N_7610,N_4573,N_5296);
nand U7611 (N_7611,N_3129,N_3274);
and U7612 (N_7612,N_3740,N_5717);
nand U7613 (N_7613,N_5754,N_4037);
or U7614 (N_7614,N_5809,N_4862);
and U7615 (N_7615,N_4371,N_3161);
and U7616 (N_7616,N_4305,N_5932);
nand U7617 (N_7617,N_4208,N_4477);
nand U7618 (N_7618,N_3179,N_4421);
and U7619 (N_7619,N_4646,N_5951);
nor U7620 (N_7620,N_3301,N_3053);
or U7621 (N_7621,N_5759,N_4826);
or U7622 (N_7622,N_5124,N_4608);
nand U7623 (N_7623,N_4534,N_3342);
and U7624 (N_7624,N_5311,N_5459);
or U7625 (N_7625,N_4638,N_3632);
and U7626 (N_7626,N_3550,N_4746);
nand U7627 (N_7627,N_3374,N_3513);
nand U7628 (N_7628,N_4917,N_4050);
or U7629 (N_7629,N_4801,N_3669);
or U7630 (N_7630,N_3294,N_3910);
or U7631 (N_7631,N_3474,N_4306);
nor U7632 (N_7632,N_3784,N_5173);
or U7633 (N_7633,N_3399,N_5421);
nor U7634 (N_7634,N_5616,N_5601);
nand U7635 (N_7635,N_5418,N_5057);
or U7636 (N_7636,N_4567,N_4683);
nor U7637 (N_7637,N_5038,N_5365);
and U7638 (N_7638,N_3222,N_4976);
nor U7639 (N_7639,N_3408,N_5763);
and U7640 (N_7640,N_3529,N_4943);
nand U7641 (N_7641,N_3378,N_5871);
nor U7642 (N_7642,N_4849,N_5227);
nor U7643 (N_7643,N_5699,N_4271);
or U7644 (N_7644,N_3109,N_5136);
nor U7645 (N_7645,N_3879,N_5199);
nor U7646 (N_7646,N_5228,N_4143);
nand U7647 (N_7647,N_5594,N_4638);
and U7648 (N_7648,N_4119,N_3818);
and U7649 (N_7649,N_5070,N_5993);
nand U7650 (N_7650,N_3709,N_3297);
or U7651 (N_7651,N_3664,N_5004);
and U7652 (N_7652,N_3695,N_3544);
or U7653 (N_7653,N_3568,N_3561);
and U7654 (N_7654,N_4328,N_3411);
and U7655 (N_7655,N_5870,N_3957);
and U7656 (N_7656,N_5713,N_5914);
nor U7657 (N_7657,N_5032,N_5742);
or U7658 (N_7658,N_5731,N_4904);
or U7659 (N_7659,N_4834,N_4371);
nand U7660 (N_7660,N_3626,N_3400);
xnor U7661 (N_7661,N_4714,N_4247);
nor U7662 (N_7662,N_5828,N_5608);
nand U7663 (N_7663,N_4518,N_5657);
nand U7664 (N_7664,N_3222,N_3787);
xnor U7665 (N_7665,N_3531,N_3960);
nor U7666 (N_7666,N_5009,N_5858);
or U7667 (N_7667,N_3788,N_4301);
and U7668 (N_7668,N_4082,N_4937);
nor U7669 (N_7669,N_3002,N_3312);
or U7670 (N_7670,N_4386,N_4972);
or U7671 (N_7671,N_3875,N_5736);
and U7672 (N_7672,N_3043,N_5807);
nor U7673 (N_7673,N_4745,N_4982);
and U7674 (N_7674,N_3581,N_3639);
nand U7675 (N_7675,N_5546,N_4989);
nor U7676 (N_7676,N_4376,N_5491);
nor U7677 (N_7677,N_4450,N_5585);
nor U7678 (N_7678,N_5057,N_4681);
and U7679 (N_7679,N_3423,N_3202);
or U7680 (N_7680,N_5984,N_5383);
or U7681 (N_7681,N_5154,N_3537);
nor U7682 (N_7682,N_4559,N_3525);
nor U7683 (N_7683,N_3620,N_3197);
nor U7684 (N_7684,N_5806,N_5915);
nor U7685 (N_7685,N_4195,N_4532);
nor U7686 (N_7686,N_5366,N_5541);
nand U7687 (N_7687,N_3396,N_5043);
and U7688 (N_7688,N_4254,N_4436);
xnor U7689 (N_7689,N_5155,N_5817);
nor U7690 (N_7690,N_4474,N_3394);
nor U7691 (N_7691,N_5829,N_3198);
nand U7692 (N_7692,N_5088,N_5950);
nand U7693 (N_7693,N_4833,N_5062);
and U7694 (N_7694,N_4504,N_4722);
nor U7695 (N_7695,N_3518,N_3957);
and U7696 (N_7696,N_3902,N_4691);
nor U7697 (N_7697,N_3372,N_4462);
nand U7698 (N_7698,N_4833,N_4374);
and U7699 (N_7699,N_5622,N_5036);
and U7700 (N_7700,N_3095,N_4308);
nor U7701 (N_7701,N_5106,N_4133);
or U7702 (N_7702,N_3697,N_5662);
nand U7703 (N_7703,N_4335,N_4802);
and U7704 (N_7704,N_4722,N_4138);
and U7705 (N_7705,N_3329,N_3701);
and U7706 (N_7706,N_5075,N_3159);
and U7707 (N_7707,N_4611,N_4301);
nand U7708 (N_7708,N_5848,N_4724);
nand U7709 (N_7709,N_4918,N_4893);
nand U7710 (N_7710,N_4864,N_3701);
nor U7711 (N_7711,N_4908,N_5168);
nor U7712 (N_7712,N_4548,N_4974);
and U7713 (N_7713,N_3428,N_4436);
or U7714 (N_7714,N_4744,N_4218);
nor U7715 (N_7715,N_4177,N_3896);
and U7716 (N_7716,N_5816,N_5736);
nor U7717 (N_7717,N_3525,N_5946);
nand U7718 (N_7718,N_4579,N_5451);
or U7719 (N_7719,N_4315,N_3177);
nand U7720 (N_7720,N_3072,N_4415);
xnor U7721 (N_7721,N_4418,N_4147);
and U7722 (N_7722,N_4943,N_4091);
or U7723 (N_7723,N_3126,N_4776);
and U7724 (N_7724,N_3956,N_3344);
or U7725 (N_7725,N_3664,N_4684);
nor U7726 (N_7726,N_4074,N_4599);
and U7727 (N_7727,N_5507,N_3760);
nand U7728 (N_7728,N_3241,N_5106);
and U7729 (N_7729,N_5623,N_4998);
or U7730 (N_7730,N_4888,N_3381);
and U7731 (N_7731,N_3111,N_5900);
and U7732 (N_7732,N_5734,N_4419);
xor U7733 (N_7733,N_5513,N_5844);
and U7734 (N_7734,N_5580,N_3379);
nand U7735 (N_7735,N_4363,N_3269);
and U7736 (N_7736,N_5332,N_3191);
or U7737 (N_7737,N_3825,N_3411);
or U7738 (N_7738,N_4672,N_5284);
and U7739 (N_7739,N_5308,N_3922);
nand U7740 (N_7740,N_5397,N_4561);
nand U7741 (N_7741,N_4519,N_4140);
nand U7742 (N_7742,N_5964,N_5153);
or U7743 (N_7743,N_5213,N_4492);
nor U7744 (N_7744,N_4975,N_3911);
nand U7745 (N_7745,N_5743,N_3732);
or U7746 (N_7746,N_3526,N_4841);
nand U7747 (N_7747,N_4692,N_5748);
nor U7748 (N_7748,N_5913,N_5218);
nand U7749 (N_7749,N_4400,N_4215);
nor U7750 (N_7750,N_5748,N_4112);
nand U7751 (N_7751,N_3317,N_4536);
nor U7752 (N_7752,N_5385,N_5438);
nand U7753 (N_7753,N_5958,N_4062);
nand U7754 (N_7754,N_3317,N_4532);
and U7755 (N_7755,N_3485,N_4368);
nand U7756 (N_7756,N_4670,N_4492);
nand U7757 (N_7757,N_3875,N_3724);
nor U7758 (N_7758,N_5146,N_4747);
and U7759 (N_7759,N_3926,N_5201);
nand U7760 (N_7760,N_5987,N_4045);
nor U7761 (N_7761,N_3112,N_4821);
or U7762 (N_7762,N_5455,N_4365);
nand U7763 (N_7763,N_4546,N_3436);
nor U7764 (N_7764,N_3101,N_4329);
nor U7765 (N_7765,N_4625,N_5710);
nand U7766 (N_7766,N_4553,N_5263);
nand U7767 (N_7767,N_5899,N_5396);
and U7768 (N_7768,N_5755,N_3381);
or U7769 (N_7769,N_4335,N_4383);
and U7770 (N_7770,N_5625,N_4721);
or U7771 (N_7771,N_5757,N_5747);
nand U7772 (N_7772,N_4216,N_3962);
nand U7773 (N_7773,N_3016,N_4451);
xor U7774 (N_7774,N_5587,N_3081);
nand U7775 (N_7775,N_5039,N_4217);
nor U7776 (N_7776,N_5058,N_4096);
or U7777 (N_7777,N_4672,N_5463);
nand U7778 (N_7778,N_4401,N_5778);
nor U7779 (N_7779,N_4337,N_5756);
and U7780 (N_7780,N_4815,N_5564);
and U7781 (N_7781,N_3828,N_4374);
or U7782 (N_7782,N_3149,N_3439);
or U7783 (N_7783,N_5861,N_4714);
and U7784 (N_7784,N_3143,N_5038);
or U7785 (N_7785,N_4834,N_4766);
nor U7786 (N_7786,N_4286,N_5357);
nand U7787 (N_7787,N_3908,N_3413);
and U7788 (N_7788,N_4088,N_3305);
xor U7789 (N_7789,N_3658,N_4131);
and U7790 (N_7790,N_3876,N_3951);
nand U7791 (N_7791,N_3389,N_3015);
and U7792 (N_7792,N_3650,N_5153);
nor U7793 (N_7793,N_3479,N_4019);
and U7794 (N_7794,N_5140,N_3980);
or U7795 (N_7795,N_5607,N_4161);
nand U7796 (N_7796,N_3472,N_4723);
xnor U7797 (N_7797,N_5733,N_5143);
and U7798 (N_7798,N_5151,N_3120);
nor U7799 (N_7799,N_5956,N_4332);
or U7800 (N_7800,N_3951,N_5118);
nor U7801 (N_7801,N_4243,N_4671);
nand U7802 (N_7802,N_4154,N_3799);
nor U7803 (N_7803,N_4496,N_5514);
xor U7804 (N_7804,N_4068,N_3658);
and U7805 (N_7805,N_3443,N_4293);
and U7806 (N_7806,N_3148,N_5723);
or U7807 (N_7807,N_5642,N_5910);
nor U7808 (N_7808,N_4612,N_3617);
and U7809 (N_7809,N_5659,N_3382);
nor U7810 (N_7810,N_4836,N_3459);
nor U7811 (N_7811,N_3167,N_4517);
or U7812 (N_7812,N_4487,N_4892);
nor U7813 (N_7813,N_5071,N_4809);
and U7814 (N_7814,N_3197,N_3977);
or U7815 (N_7815,N_5858,N_3986);
nor U7816 (N_7816,N_4080,N_5318);
and U7817 (N_7817,N_4116,N_5860);
and U7818 (N_7818,N_3341,N_3954);
and U7819 (N_7819,N_3334,N_5417);
and U7820 (N_7820,N_3974,N_4630);
or U7821 (N_7821,N_4077,N_3413);
or U7822 (N_7822,N_3127,N_4482);
or U7823 (N_7823,N_4535,N_5372);
nor U7824 (N_7824,N_4996,N_4426);
or U7825 (N_7825,N_3050,N_3560);
and U7826 (N_7826,N_3788,N_3511);
nor U7827 (N_7827,N_5214,N_3124);
and U7828 (N_7828,N_4312,N_3070);
nor U7829 (N_7829,N_3456,N_4988);
and U7830 (N_7830,N_3851,N_4147);
xnor U7831 (N_7831,N_5464,N_5590);
nor U7832 (N_7832,N_3705,N_3232);
xor U7833 (N_7833,N_4959,N_4666);
or U7834 (N_7834,N_5705,N_3239);
nand U7835 (N_7835,N_3616,N_4997);
nand U7836 (N_7836,N_5407,N_5495);
nand U7837 (N_7837,N_4956,N_5246);
nor U7838 (N_7838,N_4760,N_3889);
and U7839 (N_7839,N_4753,N_4037);
or U7840 (N_7840,N_3068,N_3505);
nor U7841 (N_7841,N_4901,N_3038);
and U7842 (N_7842,N_4642,N_4358);
or U7843 (N_7843,N_4764,N_5409);
and U7844 (N_7844,N_5900,N_5528);
nand U7845 (N_7845,N_4808,N_4252);
nor U7846 (N_7846,N_3615,N_4598);
nor U7847 (N_7847,N_4394,N_4461);
or U7848 (N_7848,N_5833,N_5522);
or U7849 (N_7849,N_4568,N_3298);
nand U7850 (N_7850,N_5473,N_3132);
nor U7851 (N_7851,N_3669,N_5840);
or U7852 (N_7852,N_4749,N_4214);
and U7853 (N_7853,N_4301,N_3679);
and U7854 (N_7854,N_5881,N_5319);
xor U7855 (N_7855,N_3685,N_3264);
nand U7856 (N_7856,N_5313,N_4111);
nor U7857 (N_7857,N_4495,N_3980);
or U7858 (N_7858,N_5996,N_5355);
or U7859 (N_7859,N_4738,N_5141);
and U7860 (N_7860,N_4227,N_4686);
and U7861 (N_7861,N_4536,N_4237);
or U7862 (N_7862,N_3018,N_3866);
and U7863 (N_7863,N_5803,N_5097);
xor U7864 (N_7864,N_3526,N_5051);
nor U7865 (N_7865,N_3117,N_5401);
nand U7866 (N_7866,N_4190,N_3052);
nand U7867 (N_7867,N_4615,N_3531);
and U7868 (N_7868,N_5161,N_5130);
nor U7869 (N_7869,N_4087,N_4018);
or U7870 (N_7870,N_4876,N_4084);
and U7871 (N_7871,N_4963,N_5012);
nor U7872 (N_7872,N_3413,N_4617);
and U7873 (N_7873,N_4500,N_3344);
nand U7874 (N_7874,N_3162,N_5181);
nand U7875 (N_7875,N_3439,N_3590);
or U7876 (N_7876,N_4098,N_3397);
and U7877 (N_7877,N_4336,N_5136);
or U7878 (N_7878,N_4853,N_3019);
or U7879 (N_7879,N_3053,N_5997);
and U7880 (N_7880,N_4342,N_3366);
or U7881 (N_7881,N_4560,N_3369);
and U7882 (N_7882,N_5590,N_5088);
nand U7883 (N_7883,N_3144,N_5677);
nand U7884 (N_7884,N_3122,N_5913);
or U7885 (N_7885,N_5262,N_4645);
or U7886 (N_7886,N_5740,N_4384);
nand U7887 (N_7887,N_4002,N_3885);
nor U7888 (N_7888,N_3517,N_3439);
or U7889 (N_7889,N_3269,N_3635);
nand U7890 (N_7890,N_4612,N_3742);
or U7891 (N_7891,N_3650,N_3162);
nand U7892 (N_7892,N_5337,N_4884);
or U7893 (N_7893,N_5710,N_3655);
nand U7894 (N_7894,N_3174,N_5921);
or U7895 (N_7895,N_4527,N_3288);
nor U7896 (N_7896,N_3787,N_4521);
nor U7897 (N_7897,N_3142,N_3687);
xnor U7898 (N_7898,N_4129,N_5252);
nand U7899 (N_7899,N_4251,N_4670);
nor U7900 (N_7900,N_3545,N_3254);
nand U7901 (N_7901,N_3238,N_5070);
nor U7902 (N_7902,N_4650,N_4756);
nor U7903 (N_7903,N_5444,N_4391);
nor U7904 (N_7904,N_4220,N_4025);
nor U7905 (N_7905,N_5542,N_3520);
or U7906 (N_7906,N_3324,N_5055);
nor U7907 (N_7907,N_4996,N_3030);
and U7908 (N_7908,N_4803,N_3473);
and U7909 (N_7909,N_4157,N_3966);
and U7910 (N_7910,N_3894,N_4923);
nand U7911 (N_7911,N_3475,N_5393);
nand U7912 (N_7912,N_5157,N_4086);
or U7913 (N_7913,N_5320,N_3265);
nand U7914 (N_7914,N_5711,N_4726);
nor U7915 (N_7915,N_4730,N_4669);
nand U7916 (N_7916,N_4402,N_4821);
xnor U7917 (N_7917,N_5346,N_5621);
xnor U7918 (N_7918,N_4222,N_4612);
nand U7919 (N_7919,N_4244,N_4491);
and U7920 (N_7920,N_5820,N_3696);
nand U7921 (N_7921,N_3492,N_5724);
nand U7922 (N_7922,N_5376,N_4259);
and U7923 (N_7923,N_4564,N_4084);
and U7924 (N_7924,N_5010,N_4904);
nand U7925 (N_7925,N_4651,N_5118);
nor U7926 (N_7926,N_5377,N_5557);
nand U7927 (N_7927,N_4203,N_4109);
or U7928 (N_7928,N_5718,N_5800);
or U7929 (N_7929,N_5094,N_3166);
nor U7930 (N_7930,N_4998,N_4773);
or U7931 (N_7931,N_5495,N_4125);
or U7932 (N_7932,N_4184,N_5372);
nand U7933 (N_7933,N_5613,N_3025);
and U7934 (N_7934,N_4978,N_4028);
nor U7935 (N_7935,N_5509,N_5665);
and U7936 (N_7936,N_4373,N_3435);
nand U7937 (N_7937,N_4948,N_5635);
nor U7938 (N_7938,N_4790,N_3803);
nor U7939 (N_7939,N_5146,N_4022);
and U7940 (N_7940,N_4070,N_5400);
or U7941 (N_7941,N_5218,N_5944);
and U7942 (N_7942,N_5014,N_4512);
nand U7943 (N_7943,N_4460,N_5354);
and U7944 (N_7944,N_3227,N_5321);
nor U7945 (N_7945,N_5418,N_4748);
nor U7946 (N_7946,N_3783,N_4295);
or U7947 (N_7947,N_4593,N_3165);
nor U7948 (N_7948,N_3251,N_3907);
or U7949 (N_7949,N_3598,N_3734);
nor U7950 (N_7950,N_3566,N_4888);
nor U7951 (N_7951,N_3949,N_4123);
or U7952 (N_7952,N_3108,N_5805);
nor U7953 (N_7953,N_3366,N_4442);
xnor U7954 (N_7954,N_3455,N_5858);
or U7955 (N_7955,N_3666,N_4998);
or U7956 (N_7956,N_3456,N_4440);
nand U7957 (N_7957,N_4881,N_3488);
nand U7958 (N_7958,N_4457,N_3763);
and U7959 (N_7959,N_5444,N_5660);
nor U7960 (N_7960,N_4287,N_3634);
or U7961 (N_7961,N_4634,N_5429);
xor U7962 (N_7962,N_5565,N_3557);
and U7963 (N_7963,N_4923,N_3807);
and U7964 (N_7964,N_5178,N_5839);
or U7965 (N_7965,N_4130,N_4703);
or U7966 (N_7966,N_4664,N_3701);
nor U7967 (N_7967,N_5843,N_4755);
and U7968 (N_7968,N_4948,N_5601);
nor U7969 (N_7969,N_3514,N_3907);
nand U7970 (N_7970,N_5733,N_5173);
and U7971 (N_7971,N_5822,N_3146);
nor U7972 (N_7972,N_4655,N_5976);
nand U7973 (N_7973,N_4180,N_5481);
xor U7974 (N_7974,N_4896,N_3999);
and U7975 (N_7975,N_4508,N_4181);
and U7976 (N_7976,N_3285,N_5315);
xor U7977 (N_7977,N_5444,N_4103);
and U7978 (N_7978,N_5179,N_3540);
nand U7979 (N_7979,N_3975,N_5970);
nand U7980 (N_7980,N_3178,N_5237);
or U7981 (N_7981,N_3244,N_4582);
nand U7982 (N_7982,N_4485,N_5541);
nand U7983 (N_7983,N_4249,N_4691);
and U7984 (N_7984,N_3288,N_5452);
nand U7985 (N_7985,N_3579,N_4555);
xnor U7986 (N_7986,N_4357,N_4244);
or U7987 (N_7987,N_5418,N_4286);
nor U7988 (N_7988,N_5521,N_5701);
or U7989 (N_7989,N_5064,N_5036);
and U7990 (N_7990,N_4659,N_5558);
or U7991 (N_7991,N_5885,N_4737);
nor U7992 (N_7992,N_5527,N_4594);
or U7993 (N_7993,N_5520,N_4312);
nand U7994 (N_7994,N_5426,N_5031);
nand U7995 (N_7995,N_3434,N_3334);
nand U7996 (N_7996,N_5406,N_5666);
or U7997 (N_7997,N_3986,N_5348);
nor U7998 (N_7998,N_5999,N_4527);
xor U7999 (N_7999,N_5548,N_3043);
or U8000 (N_8000,N_3881,N_4560);
nand U8001 (N_8001,N_3630,N_5954);
or U8002 (N_8002,N_4046,N_4391);
and U8003 (N_8003,N_4831,N_5263);
nand U8004 (N_8004,N_4834,N_5124);
nand U8005 (N_8005,N_3163,N_4655);
or U8006 (N_8006,N_5221,N_5910);
and U8007 (N_8007,N_4940,N_3095);
xnor U8008 (N_8008,N_3524,N_5483);
and U8009 (N_8009,N_4833,N_3399);
and U8010 (N_8010,N_3131,N_5797);
and U8011 (N_8011,N_5058,N_5620);
nand U8012 (N_8012,N_5053,N_4080);
nand U8013 (N_8013,N_4708,N_5057);
and U8014 (N_8014,N_5613,N_4554);
and U8015 (N_8015,N_5596,N_3244);
or U8016 (N_8016,N_4578,N_5920);
nand U8017 (N_8017,N_3277,N_3113);
and U8018 (N_8018,N_4981,N_5475);
or U8019 (N_8019,N_3479,N_5580);
or U8020 (N_8020,N_4204,N_4560);
nor U8021 (N_8021,N_5058,N_5502);
and U8022 (N_8022,N_5117,N_5550);
and U8023 (N_8023,N_3270,N_5280);
or U8024 (N_8024,N_3241,N_4969);
nand U8025 (N_8025,N_3318,N_3882);
nand U8026 (N_8026,N_5853,N_5469);
nor U8027 (N_8027,N_5283,N_4304);
or U8028 (N_8028,N_3757,N_5506);
nor U8029 (N_8029,N_4747,N_4914);
nand U8030 (N_8030,N_3333,N_4544);
or U8031 (N_8031,N_4511,N_3410);
and U8032 (N_8032,N_4758,N_5425);
and U8033 (N_8033,N_3011,N_4128);
nand U8034 (N_8034,N_4560,N_4122);
and U8035 (N_8035,N_5452,N_5568);
nand U8036 (N_8036,N_4243,N_5428);
or U8037 (N_8037,N_3904,N_3958);
or U8038 (N_8038,N_3447,N_5269);
and U8039 (N_8039,N_3924,N_4322);
nand U8040 (N_8040,N_4740,N_4655);
nand U8041 (N_8041,N_4815,N_5591);
nand U8042 (N_8042,N_3353,N_3860);
or U8043 (N_8043,N_5613,N_5766);
nand U8044 (N_8044,N_5092,N_4784);
nor U8045 (N_8045,N_3941,N_5606);
nand U8046 (N_8046,N_5235,N_5787);
nor U8047 (N_8047,N_4367,N_5289);
and U8048 (N_8048,N_5178,N_3925);
nor U8049 (N_8049,N_4096,N_5621);
nand U8050 (N_8050,N_4065,N_3615);
nand U8051 (N_8051,N_4794,N_3010);
xor U8052 (N_8052,N_5880,N_3639);
or U8053 (N_8053,N_5336,N_4518);
nor U8054 (N_8054,N_4104,N_5985);
nand U8055 (N_8055,N_4068,N_5865);
and U8056 (N_8056,N_3935,N_3284);
or U8057 (N_8057,N_5087,N_3261);
and U8058 (N_8058,N_3578,N_3705);
and U8059 (N_8059,N_3102,N_5750);
nand U8060 (N_8060,N_5141,N_4801);
nor U8061 (N_8061,N_4904,N_4367);
nand U8062 (N_8062,N_5312,N_4051);
and U8063 (N_8063,N_4899,N_4477);
xor U8064 (N_8064,N_5506,N_4064);
nor U8065 (N_8065,N_4307,N_5479);
or U8066 (N_8066,N_3378,N_5232);
and U8067 (N_8067,N_5994,N_5891);
or U8068 (N_8068,N_5514,N_5524);
nand U8069 (N_8069,N_3517,N_5505);
nand U8070 (N_8070,N_3186,N_3288);
or U8071 (N_8071,N_5990,N_3113);
and U8072 (N_8072,N_3493,N_4326);
and U8073 (N_8073,N_5308,N_5555);
nor U8074 (N_8074,N_4141,N_5996);
nand U8075 (N_8075,N_5622,N_4773);
and U8076 (N_8076,N_4905,N_4186);
and U8077 (N_8077,N_3733,N_5465);
nand U8078 (N_8078,N_4782,N_5573);
and U8079 (N_8079,N_3982,N_4333);
or U8080 (N_8080,N_5497,N_5126);
nand U8081 (N_8081,N_3166,N_3088);
nand U8082 (N_8082,N_3570,N_4941);
or U8083 (N_8083,N_4091,N_3054);
or U8084 (N_8084,N_3593,N_4067);
nand U8085 (N_8085,N_5766,N_5983);
or U8086 (N_8086,N_5926,N_4852);
or U8087 (N_8087,N_4410,N_4746);
nor U8088 (N_8088,N_5408,N_4955);
nor U8089 (N_8089,N_5890,N_3213);
and U8090 (N_8090,N_4122,N_4709);
and U8091 (N_8091,N_5761,N_5942);
or U8092 (N_8092,N_4663,N_3119);
or U8093 (N_8093,N_3798,N_4938);
or U8094 (N_8094,N_4390,N_4578);
xnor U8095 (N_8095,N_3192,N_4649);
nor U8096 (N_8096,N_5332,N_4917);
nor U8097 (N_8097,N_3598,N_4145);
xnor U8098 (N_8098,N_5219,N_4893);
or U8099 (N_8099,N_5885,N_3237);
and U8100 (N_8100,N_5087,N_3526);
nor U8101 (N_8101,N_4056,N_3027);
nand U8102 (N_8102,N_3050,N_3940);
nand U8103 (N_8103,N_4777,N_4738);
or U8104 (N_8104,N_5896,N_3527);
or U8105 (N_8105,N_3147,N_3446);
nor U8106 (N_8106,N_3838,N_3604);
or U8107 (N_8107,N_4013,N_5406);
nor U8108 (N_8108,N_3616,N_3316);
or U8109 (N_8109,N_4611,N_3623);
and U8110 (N_8110,N_3112,N_4955);
or U8111 (N_8111,N_3358,N_5553);
nor U8112 (N_8112,N_4573,N_4271);
and U8113 (N_8113,N_4231,N_5710);
or U8114 (N_8114,N_4380,N_3388);
nor U8115 (N_8115,N_3416,N_5738);
nor U8116 (N_8116,N_3839,N_5262);
or U8117 (N_8117,N_5811,N_3518);
or U8118 (N_8118,N_3839,N_3873);
nand U8119 (N_8119,N_4945,N_5345);
and U8120 (N_8120,N_5174,N_5955);
or U8121 (N_8121,N_5245,N_3750);
and U8122 (N_8122,N_4893,N_5969);
or U8123 (N_8123,N_5513,N_5515);
or U8124 (N_8124,N_3998,N_4207);
nor U8125 (N_8125,N_5245,N_3373);
xnor U8126 (N_8126,N_5619,N_4532);
nor U8127 (N_8127,N_4272,N_3335);
nand U8128 (N_8128,N_4894,N_5761);
and U8129 (N_8129,N_5155,N_4592);
and U8130 (N_8130,N_3258,N_3304);
and U8131 (N_8131,N_4486,N_4516);
nand U8132 (N_8132,N_5648,N_4141);
nand U8133 (N_8133,N_4057,N_4698);
nor U8134 (N_8134,N_4283,N_5850);
nor U8135 (N_8135,N_3770,N_3450);
nand U8136 (N_8136,N_3936,N_3527);
nor U8137 (N_8137,N_4815,N_3850);
or U8138 (N_8138,N_5088,N_4810);
and U8139 (N_8139,N_4036,N_4263);
or U8140 (N_8140,N_4945,N_4879);
and U8141 (N_8141,N_3035,N_5958);
nand U8142 (N_8142,N_3350,N_3760);
nor U8143 (N_8143,N_3221,N_3910);
nand U8144 (N_8144,N_5327,N_4805);
nand U8145 (N_8145,N_3111,N_5943);
nand U8146 (N_8146,N_4536,N_4146);
nand U8147 (N_8147,N_4528,N_4841);
and U8148 (N_8148,N_4331,N_4813);
nor U8149 (N_8149,N_4877,N_4215);
nand U8150 (N_8150,N_5563,N_3730);
nor U8151 (N_8151,N_5775,N_5148);
nor U8152 (N_8152,N_5249,N_4454);
nor U8153 (N_8153,N_3401,N_3755);
nand U8154 (N_8154,N_4195,N_3186);
nor U8155 (N_8155,N_5707,N_3507);
and U8156 (N_8156,N_3646,N_3837);
and U8157 (N_8157,N_3906,N_5131);
nor U8158 (N_8158,N_4618,N_5721);
or U8159 (N_8159,N_3684,N_5762);
and U8160 (N_8160,N_3576,N_5736);
or U8161 (N_8161,N_3082,N_5062);
nand U8162 (N_8162,N_4340,N_5037);
nand U8163 (N_8163,N_4753,N_4537);
nand U8164 (N_8164,N_5741,N_5921);
xnor U8165 (N_8165,N_4228,N_5895);
nor U8166 (N_8166,N_4722,N_4271);
nor U8167 (N_8167,N_5962,N_3384);
and U8168 (N_8168,N_5283,N_5802);
nor U8169 (N_8169,N_4665,N_4226);
or U8170 (N_8170,N_5553,N_3233);
and U8171 (N_8171,N_4649,N_5384);
nand U8172 (N_8172,N_5286,N_5670);
or U8173 (N_8173,N_3820,N_3543);
nand U8174 (N_8174,N_4572,N_3522);
or U8175 (N_8175,N_3777,N_5374);
or U8176 (N_8176,N_5397,N_4079);
and U8177 (N_8177,N_4108,N_5198);
nor U8178 (N_8178,N_3149,N_5509);
or U8179 (N_8179,N_4811,N_4603);
xor U8180 (N_8180,N_4280,N_5633);
or U8181 (N_8181,N_4571,N_5348);
nand U8182 (N_8182,N_3285,N_3889);
or U8183 (N_8183,N_3559,N_4588);
nand U8184 (N_8184,N_3496,N_4681);
or U8185 (N_8185,N_4805,N_5144);
and U8186 (N_8186,N_5809,N_5840);
nor U8187 (N_8187,N_3871,N_3563);
or U8188 (N_8188,N_3437,N_4872);
and U8189 (N_8189,N_3994,N_3647);
nand U8190 (N_8190,N_4651,N_5537);
and U8191 (N_8191,N_3264,N_4341);
nand U8192 (N_8192,N_5298,N_4403);
nand U8193 (N_8193,N_4338,N_4278);
or U8194 (N_8194,N_3246,N_3846);
or U8195 (N_8195,N_4203,N_3226);
and U8196 (N_8196,N_3478,N_5409);
nor U8197 (N_8197,N_5627,N_5832);
or U8198 (N_8198,N_5305,N_4842);
nor U8199 (N_8199,N_4982,N_5366);
or U8200 (N_8200,N_5255,N_3224);
or U8201 (N_8201,N_4164,N_5410);
nor U8202 (N_8202,N_3928,N_3726);
or U8203 (N_8203,N_4105,N_5987);
nor U8204 (N_8204,N_5242,N_5595);
or U8205 (N_8205,N_3126,N_3968);
and U8206 (N_8206,N_5126,N_4348);
nand U8207 (N_8207,N_4870,N_3377);
and U8208 (N_8208,N_4101,N_3248);
nand U8209 (N_8209,N_4975,N_4521);
nor U8210 (N_8210,N_4395,N_5899);
xor U8211 (N_8211,N_4638,N_3818);
nor U8212 (N_8212,N_5111,N_4796);
and U8213 (N_8213,N_4703,N_4283);
nand U8214 (N_8214,N_4231,N_3761);
nand U8215 (N_8215,N_4862,N_3266);
nand U8216 (N_8216,N_4105,N_4632);
nor U8217 (N_8217,N_3070,N_4020);
nand U8218 (N_8218,N_4848,N_4516);
and U8219 (N_8219,N_4487,N_4668);
xor U8220 (N_8220,N_4450,N_4880);
nand U8221 (N_8221,N_4672,N_4417);
nor U8222 (N_8222,N_3303,N_3398);
or U8223 (N_8223,N_5432,N_5821);
nor U8224 (N_8224,N_5489,N_3969);
or U8225 (N_8225,N_4152,N_4323);
and U8226 (N_8226,N_3323,N_5554);
nor U8227 (N_8227,N_5384,N_5485);
nand U8228 (N_8228,N_5669,N_5239);
and U8229 (N_8229,N_5622,N_3462);
nor U8230 (N_8230,N_4006,N_3320);
and U8231 (N_8231,N_5209,N_5762);
and U8232 (N_8232,N_5348,N_3763);
nand U8233 (N_8233,N_5180,N_3067);
or U8234 (N_8234,N_4217,N_3520);
nor U8235 (N_8235,N_4508,N_3870);
and U8236 (N_8236,N_5781,N_4833);
nand U8237 (N_8237,N_5908,N_3097);
or U8238 (N_8238,N_3931,N_4338);
nor U8239 (N_8239,N_3230,N_4220);
or U8240 (N_8240,N_3298,N_3297);
or U8241 (N_8241,N_3055,N_3859);
nand U8242 (N_8242,N_3679,N_4326);
and U8243 (N_8243,N_3589,N_5254);
or U8244 (N_8244,N_4654,N_3684);
or U8245 (N_8245,N_5194,N_4644);
nand U8246 (N_8246,N_4048,N_4339);
and U8247 (N_8247,N_3921,N_3972);
or U8248 (N_8248,N_4414,N_3401);
nor U8249 (N_8249,N_4057,N_5198);
or U8250 (N_8250,N_3552,N_5495);
and U8251 (N_8251,N_3650,N_4801);
nor U8252 (N_8252,N_4370,N_3418);
nand U8253 (N_8253,N_5431,N_5654);
nor U8254 (N_8254,N_4231,N_5798);
and U8255 (N_8255,N_4508,N_4159);
xnor U8256 (N_8256,N_3606,N_4654);
nand U8257 (N_8257,N_5369,N_3721);
nand U8258 (N_8258,N_3878,N_3359);
nand U8259 (N_8259,N_4706,N_4623);
or U8260 (N_8260,N_3902,N_4429);
and U8261 (N_8261,N_3987,N_4354);
nor U8262 (N_8262,N_4084,N_5021);
nand U8263 (N_8263,N_5898,N_3472);
nor U8264 (N_8264,N_3677,N_3578);
nand U8265 (N_8265,N_5109,N_4472);
and U8266 (N_8266,N_3823,N_5055);
nand U8267 (N_8267,N_5071,N_3946);
nor U8268 (N_8268,N_4975,N_4880);
nand U8269 (N_8269,N_4682,N_5773);
nor U8270 (N_8270,N_5237,N_5886);
and U8271 (N_8271,N_4178,N_5940);
and U8272 (N_8272,N_5199,N_5472);
nor U8273 (N_8273,N_5505,N_5506);
nor U8274 (N_8274,N_3685,N_5381);
or U8275 (N_8275,N_5899,N_3566);
nand U8276 (N_8276,N_4494,N_5340);
xor U8277 (N_8277,N_4444,N_4100);
or U8278 (N_8278,N_4227,N_3540);
or U8279 (N_8279,N_4809,N_4665);
or U8280 (N_8280,N_5898,N_5010);
nand U8281 (N_8281,N_3704,N_5997);
nand U8282 (N_8282,N_3187,N_5849);
nor U8283 (N_8283,N_5455,N_5886);
nand U8284 (N_8284,N_3573,N_5271);
nor U8285 (N_8285,N_3098,N_4845);
nand U8286 (N_8286,N_5025,N_3787);
nand U8287 (N_8287,N_3236,N_4870);
nor U8288 (N_8288,N_3945,N_3310);
and U8289 (N_8289,N_3721,N_5075);
nor U8290 (N_8290,N_3032,N_5080);
or U8291 (N_8291,N_4882,N_3891);
nand U8292 (N_8292,N_3864,N_3048);
nor U8293 (N_8293,N_4858,N_4242);
or U8294 (N_8294,N_5887,N_4265);
or U8295 (N_8295,N_5339,N_4446);
nor U8296 (N_8296,N_4832,N_4761);
or U8297 (N_8297,N_4591,N_5460);
and U8298 (N_8298,N_4005,N_5898);
and U8299 (N_8299,N_4858,N_3794);
nor U8300 (N_8300,N_5152,N_4867);
nand U8301 (N_8301,N_5731,N_4649);
nor U8302 (N_8302,N_4590,N_5494);
and U8303 (N_8303,N_5982,N_3702);
or U8304 (N_8304,N_4980,N_5770);
and U8305 (N_8305,N_3545,N_5177);
and U8306 (N_8306,N_5331,N_5397);
nor U8307 (N_8307,N_5465,N_5902);
or U8308 (N_8308,N_4247,N_3599);
nand U8309 (N_8309,N_5993,N_5828);
nor U8310 (N_8310,N_4462,N_3703);
xnor U8311 (N_8311,N_4916,N_5801);
and U8312 (N_8312,N_3058,N_3224);
and U8313 (N_8313,N_5881,N_4133);
and U8314 (N_8314,N_3744,N_5486);
nand U8315 (N_8315,N_3294,N_5434);
and U8316 (N_8316,N_3978,N_5755);
or U8317 (N_8317,N_4019,N_3017);
and U8318 (N_8318,N_5289,N_3259);
nor U8319 (N_8319,N_4180,N_3369);
nand U8320 (N_8320,N_4379,N_3017);
or U8321 (N_8321,N_5277,N_5087);
and U8322 (N_8322,N_5710,N_5548);
and U8323 (N_8323,N_5944,N_4072);
xnor U8324 (N_8324,N_5810,N_5993);
and U8325 (N_8325,N_4781,N_5628);
or U8326 (N_8326,N_4604,N_3185);
or U8327 (N_8327,N_3740,N_3617);
and U8328 (N_8328,N_3864,N_5168);
or U8329 (N_8329,N_3847,N_3399);
and U8330 (N_8330,N_3215,N_3982);
and U8331 (N_8331,N_3447,N_3850);
or U8332 (N_8332,N_5182,N_3516);
nand U8333 (N_8333,N_4864,N_3421);
and U8334 (N_8334,N_5926,N_5733);
and U8335 (N_8335,N_3089,N_3666);
nor U8336 (N_8336,N_4283,N_3071);
or U8337 (N_8337,N_5303,N_3051);
and U8338 (N_8338,N_4270,N_5780);
and U8339 (N_8339,N_5724,N_4396);
nand U8340 (N_8340,N_4279,N_3762);
and U8341 (N_8341,N_3097,N_5933);
xnor U8342 (N_8342,N_3462,N_3124);
nand U8343 (N_8343,N_4782,N_4494);
or U8344 (N_8344,N_5324,N_5684);
nand U8345 (N_8345,N_3293,N_4351);
or U8346 (N_8346,N_4766,N_3959);
or U8347 (N_8347,N_3250,N_5330);
nand U8348 (N_8348,N_5287,N_3104);
nand U8349 (N_8349,N_3935,N_5042);
nor U8350 (N_8350,N_5264,N_3426);
and U8351 (N_8351,N_4557,N_4949);
nor U8352 (N_8352,N_4571,N_4092);
nand U8353 (N_8353,N_3534,N_5585);
xnor U8354 (N_8354,N_3532,N_4412);
or U8355 (N_8355,N_4264,N_5023);
or U8356 (N_8356,N_3203,N_5823);
and U8357 (N_8357,N_4089,N_3697);
nor U8358 (N_8358,N_5339,N_4060);
nor U8359 (N_8359,N_3795,N_3744);
and U8360 (N_8360,N_3322,N_4094);
nand U8361 (N_8361,N_3766,N_4789);
nor U8362 (N_8362,N_3720,N_5881);
and U8363 (N_8363,N_5926,N_4591);
or U8364 (N_8364,N_3074,N_4353);
and U8365 (N_8365,N_3742,N_3189);
nand U8366 (N_8366,N_5750,N_3643);
and U8367 (N_8367,N_5652,N_4819);
nor U8368 (N_8368,N_4352,N_4245);
or U8369 (N_8369,N_4628,N_5082);
nor U8370 (N_8370,N_3828,N_5710);
nor U8371 (N_8371,N_4173,N_5901);
or U8372 (N_8372,N_5432,N_3367);
nand U8373 (N_8373,N_5014,N_4966);
nor U8374 (N_8374,N_5185,N_5526);
nor U8375 (N_8375,N_4181,N_5337);
nand U8376 (N_8376,N_5206,N_5683);
and U8377 (N_8377,N_4011,N_5052);
or U8378 (N_8378,N_4439,N_4496);
nand U8379 (N_8379,N_3982,N_4863);
and U8380 (N_8380,N_4729,N_4904);
or U8381 (N_8381,N_5571,N_3429);
nand U8382 (N_8382,N_4817,N_3035);
nand U8383 (N_8383,N_5905,N_3152);
and U8384 (N_8384,N_3938,N_5939);
nor U8385 (N_8385,N_4939,N_5872);
or U8386 (N_8386,N_3624,N_4220);
or U8387 (N_8387,N_5303,N_5220);
nor U8388 (N_8388,N_3174,N_3858);
and U8389 (N_8389,N_4276,N_5561);
nor U8390 (N_8390,N_4483,N_4160);
or U8391 (N_8391,N_5631,N_5915);
nand U8392 (N_8392,N_5535,N_3817);
nor U8393 (N_8393,N_5458,N_4882);
nand U8394 (N_8394,N_4201,N_3982);
nor U8395 (N_8395,N_5164,N_5855);
and U8396 (N_8396,N_4845,N_5320);
nand U8397 (N_8397,N_3991,N_3449);
nor U8398 (N_8398,N_5828,N_3863);
and U8399 (N_8399,N_5194,N_5218);
nand U8400 (N_8400,N_4103,N_4458);
or U8401 (N_8401,N_5764,N_4609);
nor U8402 (N_8402,N_4662,N_5103);
nand U8403 (N_8403,N_3153,N_4573);
nor U8404 (N_8404,N_3810,N_3253);
and U8405 (N_8405,N_5794,N_4400);
and U8406 (N_8406,N_5566,N_4425);
or U8407 (N_8407,N_4401,N_3462);
or U8408 (N_8408,N_4799,N_3038);
nand U8409 (N_8409,N_3960,N_4826);
xor U8410 (N_8410,N_5883,N_3174);
nand U8411 (N_8411,N_5966,N_4801);
and U8412 (N_8412,N_3500,N_3001);
nand U8413 (N_8413,N_4240,N_4611);
and U8414 (N_8414,N_4956,N_3329);
and U8415 (N_8415,N_4833,N_5577);
nor U8416 (N_8416,N_3881,N_4849);
and U8417 (N_8417,N_3538,N_3564);
nand U8418 (N_8418,N_3132,N_3281);
or U8419 (N_8419,N_3743,N_4950);
or U8420 (N_8420,N_3991,N_3693);
nand U8421 (N_8421,N_5765,N_3337);
xor U8422 (N_8422,N_4406,N_3696);
and U8423 (N_8423,N_3561,N_3672);
nor U8424 (N_8424,N_5560,N_3689);
nand U8425 (N_8425,N_4905,N_3554);
and U8426 (N_8426,N_3178,N_5562);
or U8427 (N_8427,N_3612,N_5227);
or U8428 (N_8428,N_4827,N_4686);
nor U8429 (N_8429,N_5500,N_5980);
and U8430 (N_8430,N_3930,N_3684);
or U8431 (N_8431,N_5445,N_3148);
or U8432 (N_8432,N_3273,N_5081);
nor U8433 (N_8433,N_3995,N_5151);
nand U8434 (N_8434,N_3408,N_4606);
nor U8435 (N_8435,N_5641,N_3183);
and U8436 (N_8436,N_4784,N_4283);
nand U8437 (N_8437,N_5043,N_3352);
or U8438 (N_8438,N_3858,N_4071);
and U8439 (N_8439,N_5057,N_5648);
or U8440 (N_8440,N_5880,N_3535);
and U8441 (N_8441,N_4032,N_4342);
and U8442 (N_8442,N_5466,N_4457);
and U8443 (N_8443,N_3066,N_3811);
nor U8444 (N_8444,N_3134,N_4714);
nand U8445 (N_8445,N_4393,N_4476);
nand U8446 (N_8446,N_3512,N_3641);
and U8447 (N_8447,N_5109,N_4874);
or U8448 (N_8448,N_3442,N_5664);
and U8449 (N_8449,N_3683,N_5259);
or U8450 (N_8450,N_3091,N_5399);
and U8451 (N_8451,N_4664,N_3346);
or U8452 (N_8452,N_3183,N_5428);
nor U8453 (N_8453,N_3095,N_5085);
or U8454 (N_8454,N_5634,N_5724);
xor U8455 (N_8455,N_3928,N_3161);
nand U8456 (N_8456,N_5405,N_4597);
and U8457 (N_8457,N_3931,N_5402);
and U8458 (N_8458,N_5186,N_4443);
nor U8459 (N_8459,N_5473,N_5509);
nand U8460 (N_8460,N_4661,N_5947);
nor U8461 (N_8461,N_5827,N_5006);
xor U8462 (N_8462,N_4296,N_4424);
nor U8463 (N_8463,N_5842,N_5555);
nor U8464 (N_8464,N_3333,N_4426);
and U8465 (N_8465,N_4070,N_3085);
nor U8466 (N_8466,N_4309,N_5327);
and U8467 (N_8467,N_4480,N_5086);
or U8468 (N_8468,N_4801,N_3802);
or U8469 (N_8469,N_4724,N_4617);
or U8470 (N_8470,N_3028,N_3302);
or U8471 (N_8471,N_5253,N_3700);
and U8472 (N_8472,N_3512,N_4267);
or U8473 (N_8473,N_3128,N_4970);
nand U8474 (N_8474,N_3573,N_4514);
and U8475 (N_8475,N_5479,N_5402);
nor U8476 (N_8476,N_4112,N_4712);
nor U8477 (N_8477,N_3533,N_3546);
nor U8478 (N_8478,N_4266,N_5534);
nand U8479 (N_8479,N_5923,N_5033);
nand U8480 (N_8480,N_5017,N_4095);
or U8481 (N_8481,N_5976,N_3978);
or U8482 (N_8482,N_5203,N_4112);
nand U8483 (N_8483,N_3927,N_5933);
or U8484 (N_8484,N_3663,N_5735);
xnor U8485 (N_8485,N_4072,N_4580);
and U8486 (N_8486,N_5955,N_3624);
or U8487 (N_8487,N_3065,N_5671);
nor U8488 (N_8488,N_5875,N_4621);
and U8489 (N_8489,N_3161,N_3057);
or U8490 (N_8490,N_5041,N_4294);
or U8491 (N_8491,N_3751,N_4958);
and U8492 (N_8492,N_3384,N_3031);
and U8493 (N_8493,N_3442,N_3478);
or U8494 (N_8494,N_4465,N_5758);
nand U8495 (N_8495,N_5591,N_5917);
and U8496 (N_8496,N_5636,N_3644);
and U8497 (N_8497,N_4767,N_4440);
nor U8498 (N_8498,N_3973,N_5038);
and U8499 (N_8499,N_5142,N_3268);
or U8500 (N_8500,N_3150,N_5677);
nand U8501 (N_8501,N_4302,N_3582);
or U8502 (N_8502,N_5103,N_5670);
nor U8503 (N_8503,N_3990,N_4410);
nand U8504 (N_8504,N_3845,N_5783);
and U8505 (N_8505,N_3179,N_3356);
nor U8506 (N_8506,N_5965,N_4516);
nor U8507 (N_8507,N_4519,N_5476);
nor U8508 (N_8508,N_5164,N_4556);
or U8509 (N_8509,N_3217,N_5246);
nor U8510 (N_8510,N_3948,N_3174);
nand U8511 (N_8511,N_5153,N_5008);
xor U8512 (N_8512,N_3975,N_5827);
or U8513 (N_8513,N_4256,N_3158);
nand U8514 (N_8514,N_3574,N_5031);
and U8515 (N_8515,N_5089,N_3091);
and U8516 (N_8516,N_3418,N_4532);
nand U8517 (N_8517,N_3833,N_3344);
nand U8518 (N_8518,N_3547,N_3763);
or U8519 (N_8519,N_5784,N_3279);
and U8520 (N_8520,N_4914,N_4416);
nand U8521 (N_8521,N_4726,N_4278);
and U8522 (N_8522,N_5523,N_4810);
nor U8523 (N_8523,N_4795,N_3058);
and U8524 (N_8524,N_5750,N_3583);
and U8525 (N_8525,N_3774,N_3478);
or U8526 (N_8526,N_5389,N_5231);
nor U8527 (N_8527,N_5612,N_3405);
nand U8528 (N_8528,N_3993,N_5816);
and U8529 (N_8529,N_5473,N_3259);
nor U8530 (N_8530,N_3495,N_5364);
nor U8531 (N_8531,N_4853,N_3097);
nand U8532 (N_8532,N_3056,N_5316);
nor U8533 (N_8533,N_3798,N_5815);
nor U8534 (N_8534,N_5828,N_5206);
and U8535 (N_8535,N_4220,N_4922);
or U8536 (N_8536,N_4333,N_3220);
and U8537 (N_8537,N_3322,N_3925);
nand U8538 (N_8538,N_3783,N_5433);
nand U8539 (N_8539,N_3644,N_4964);
or U8540 (N_8540,N_5938,N_5090);
nor U8541 (N_8541,N_3815,N_5096);
or U8542 (N_8542,N_3474,N_4467);
and U8543 (N_8543,N_4860,N_5725);
nor U8544 (N_8544,N_4373,N_3532);
nand U8545 (N_8545,N_4829,N_4889);
or U8546 (N_8546,N_4824,N_4497);
nand U8547 (N_8547,N_3813,N_5745);
nand U8548 (N_8548,N_3397,N_3151);
and U8549 (N_8549,N_4980,N_4258);
nor U8550 (N_8550,N_4430,N_5720);
and U8551 (N_8551,N_3019,N_5290);
xnor U8552 (N_8552,N_5282,N_3066);
nor U8553 (N_8553,N_4049,N_3352);
and U8554 (N_8554,N_4092,N_3609);
nand U8555 (N_8555,N_4743,N_3302);
and U8556 (N_8556,N_5636,N_3400);
nand U8557 (N_8557,N_5561,N_4791);
nand U8558 (N_8558,N_5549,N_5977);
nand U8559 (N_8559,N_4892,N_3799);
and U8560 (N_8560,N_4440,N_4601);
and U8561 (N_8561,N_3676,N_3004);
nor U8562 (N_8562,N_4319,N_4612);
nand U8563 (N_8563,N_5786,N_5151);
nor U8564 (N_8564,N_4768,N_5455);
or U8565 (N_8565,N_5616,N_3245);
nand U8566 (N_8566,N_3139,N_5525);
nor U8567 (N_8567,N_4075,N_4225);
nand U8568 (N_8568,N_5919,N_5291);
nand U8569 (N_8569,N_4402,N_4829);
and U8570 (N_8570,N_3023,N_4240);
nor U8571 (N_8571,N_5644,N_3443);
or U8572 (N_8572,N_3670,N_3803);
nand U8573 (N_8573,N_4974,N_3942);
and U8574 (N_8574,N_3305,N_3536);
nor U8575 (N_8575,N_3848,N_5683);
nor U8576 (N_8576,N_5556,N_3021);
nor U8577 (N_8577,N_3749,N_4043);
and U8578 (N_8578,N_3694,N_3610);
and U8579 (N_8579,N_4084,N_4440);
xnor U8580 (N_8580,N_5153,N_4672);
nand U8581 (N_8581,N_3174,N_5152);
or U8582 (N_8582,N_5259,N_4328);
and U8583 (N_8583,N_5656,N_4778);
nor U8584 (N_8584,N_4534,N_3414);
or U8585 (N_8585,N_5317,N_5294);
and U8586 (N_8586,N_4541,N_4124);
and U8587 (N_8587,N_4332,N_3774);
and U8588 (N_8588,N_4202,N_4210);
or U8589 (N_8589,N_3928,N_3173);
xnor U8590 (N_8590,N_3349,N_3047);
or U8591 (N_8591,N_4772,N_4802);
or U8592 (N_8592,N_4835,N_4862);
nor U8593 (N_8593,N_4992,N_4920);
or U8594 (N_8594,N_4021,N_3924);
or U8595 (N_8595,N_3816,N_5014);
and U8596 (N_8596,N_3835,N_4312);
nor U8597 (N_8597,N_4412,N_5215);
nor U8598 (N_8598,N_5240,N_3156);
or U8599 (N_8599,N_4096,N_3837);
nand U8600 (N_8600,N_5604,N_5866);
or U8601 (N_8601,N_3116,N_4428);
and U8602 (N_8602,N_3557,N_5109);
and U8603 (N_8603,N_5647,N_5500);
nor U8604 (N_8604,N_4857,N_4863);
or U8605 (N_8605,N_5279,N_4090);
and U8606 (N_8606,N_3544,N_4614);
or U8607 (N_8607,N_5824,N_5995);
nor U8608 (N_8608,N_3615,N_5460);
xor U8609 (N_8609,N_3603,N_4465);
nand U8610 (N_8610,N_3461,N_5453);
nand U8611 (N_8611,N_5170,N_5004);
nor U8612 (N_8612,N_3204,N_3933);
nand U8613 (N_8613,N_3357,N_5872);
nor U8614 (N_8614,N_5778,N_5777);
nand U8615 (N_8615,N_4017,N_3170);
and U8616 (N_8616,N_4102,N_5863);
xor U8617 (N_8617,N_5701,N_5507);
and U8618 (N_8618,N_4934,N_5432);
nand U8619 (N_8619,N_4740,N_4114);
and U8620 (N_8620,N_5507,N_3284);
nand U8621 (N_8621,N_3024,N_3223);
or U8622 (N_8622,N_5804,N_3977);
nand U8623 (N_8623,N_5395,N_4286);
nand U8624 (N_8624,N_4483,N_5858);
nand U8625 (N_8625,N_3651,N_3968);
nand U8626 (N_8626,N_5193,N_4116);
or U8627 (N_8627,N_4660,N_4698);
and U8628 (N_8628,N_5374,N_3323);
nor U8629 (N_8629,N_3912,N_5445);
and U8630 (N_8630,N_4800,N_4507);
and U8631 (N_8631,N_4420,N_3869);
nor U8632 (N_8632,N_4014,N_5985);
nand U8633 (N_8633,N_4212,N_5186);
xnor U8634 (N_8634,N_5076,N_3620);
xor U8635 (N_8635,N_3848,N_5238);
nand U8636 (N_8636,N_3621,N_3388);
and U8637 (N_8637,N_4262,N_3604);
or U8638 (N_8638,N_3926,N_5213);
nor U8639 (N_8639,N_4079,N_4078);
and U8640 (N_8640,N_3310,N_4651);
nor U8641 (N_8641,N_3696,N_5141);
nand U8642 (N_8642,N_3780,N_4501);
nand U8643 (N_8643,N_3489,N_5366);
xor U8644 (N_8644,N_5419,N_5571);
nand U8645 (N_8645,N_3277,N_5682);
and U8646 (N_8646,N_3461,N_5096);
nand U8647 (N_8647,N_4184,N_3052);
and U8648 (N_8648,N_5479,N_4737);
and U8649 (N_8649,N_5218,N_4698);
nor U8650 (N_8650,N_5961,N_4702);
and U8651 (N_8651,N_3405,N_3822);
nor U8652 (N_8652,N_4377,N_3742);
and U8653 (N_8653,N_4254,N_4030);
nor U8654 (N_8654,N_5611,N_5233);
or U8655 (N_8655,N_5633,N_5778);
nor U8656 (N_8656,N_4979,N_3919);
nor U8657 (N_8657,N_3797,N_4760);
or U8658 (N_8658,N_4130,N_5292);
or U8659 (N_8659,N_3822,N_3854);
xor U8660 (N_8660,N_5380,N_3567);
nand U8661 (N_8661,N_3519,N_5477);
nor U8662 (N_8662,N_3816,N_5082);
and U8663 (N_8663,N_3183,N_3392);
or U8664 (N_8664,N_4549,N_3471);
or U8665 (N_8665,N_5319,N_3035);
and U8666 (N_8666,N_3126,N_3464);
nor U8667 (N_8667,N_5862,N_5775);
nand U8668 (N_8668,N_5708,N_3357);
nor U8669 (N_8669,N_4773,N_3771);
nand U8670 (N_8670,N_5189,N_5592);
and U8671 (N_8671,N_5485,N_5282);
and U8672 (N_8672,N_5600,N_4022);
nand U8673 (N_8673,N_4839,N_3875);
and U8674 (N_8674,N_5254,N_3935);
or U8675 (N_8675,N_4585,N_4971);
nand U8676 (N_8676,N_5565,N_3675);
and U8677 (N_8677,N_5927,N_3678);
and U8678 (N_8678,N_4959,N_5850);
and U8679 (N_8679,N_5507,N_3436);
nand U8680 (N_8680,N_4814,N_5350);
or U8681 (N_8681,N_3590,N_3460);
nor U8682 (N_8682,N_5397,N_3470);
xnor U8683 (N_8683,N_3990,N_4199);
nor U8684 (N_8684,N_4819,N_5370);
and U8685 (N_8685,N_3770,N_5009);
or U8686 (N_8686,N_5665,N_3884);
and U8687 (N_8687,N_3000,N_3251);
or U8688 (N_8688,N_5839,N_5602);
nand U8689 (N_8689,N_5992,N_5091);
nor U8690 (N_8690,N_5908,N_4862);
or U8691 (N_8691,N_5633,N_5264);
or U8692 (N_8692,N_5775,N_3494);
nand U8693 (N_8693,N_5652,N_3337);
nand U8694 (N_8694,N_4869,N_5902);
nor U8695 (N_8695,N_5572,N_4096);
and U8696 (N_8696,N_5202,N_5321);
nand U8697 (N_8697,N_4168,N_3846);
and U8698 (N_8698,N_3028,N_4589);
and U8699 (N_8699,N_3815,N_5241);
or U8700 (N_8700,N_4712,N_3023);
and U8701 (N_8701,N_3821,N_3051);
nor U8702 (N_8702,N_5343,N_5197);
and U8703 (N_8703,N_4606,N_4316);
and U8704 (N_8704,N_4216,N_4548);
and U8705 (N_8705,N_3797,N_4684);
or U8706 (N_8706,N_4405,N_3416);
and U8707 (N_8707,N_3352,N_5388);
and U8708 (N_8708,N_5574,N_4645);
nand U8709 (N_8709,N_3432,N_3017);
nand U8710 (N_8710,N_5093,N_5413);
nor U8711 (N_8711,N_3567,N_3838);
nor U8712 (N_8712,N_5652,N_3678);
or U8713 (N_8713,N_5429,N_5921);
nand U8714 (N_8714,N_5422,N_3482);
and U8715 (N_8715,N_4046,N_3465);
and U8716 (N_8716,N_5691,N_3255);
nor U8717 (N_8717,N_3927,N_3034);
nor U8718 (N_8718,N_3548,N_4660);
or U8719 (N_8719,N_4609,N_4650);
or U8720 (N_8720,N_4345,N_4251);
or U8721 (N_8721,N_4254,N_4429);
or U8722 (N_8722,N_5558,N_4285);
or U8723 (N_8723,N_5755,N_5645);
nor U8724 (N_8724,N_5713,N_5684);
nand U8725 (N_8725,N_5977,N_5858);
or U8726 (N_8726,N_5627,N_4154);
nor U8727 (N_8727,N_3560,N_5126);
or U8728 (N_8728,N_5261,N_5327);
or U8729 (N_8729,N_4897,N_5898);
nor U8730 (N_8730,N_4396,N_4143);
and U8731 (N_8731,N_3354,N_3526);
or U8732 (N_8732,N_3486,N_3402);
nand U8733 (N_8733,N_3418,N_5093);
nor U8734 (N_8734,N_4272,N_5340);
or U8735 (N_8735,N_3413,N_4206);
or U8736 (N_8736,N_5822,N_5236);
nor U8737 (N_8737,N_5825,N_5396);
or U8738 (N_8738,N_4594,N_5701);
or U8739 (N_8739,N_5407,N_4866);
and U8740 (N_8740,N_3575,N_4055);
or U8741 (N_8741,N_3758,N_5917);
nor U8742 (N_8742,N_4353,N_5732);
nor U8743 (N_8743,N_5965,N_4609);
xor U8744 (N_8744,N_5582,N_5756);
and U8745 (N_8745,N_3378,N_4556);
nand U8746 (N_8746,N_4405,N_3258);
and U8747 (N_8747,N_4858,N_5194);
nand U8748 (N_8748,N_5670,N_5238);
nor U8749 (N_8749,N_5371,N_4651);
nand U8750 (N_8750,N_5685,N_3409);
nand U8751 (N_8751,N_4897,N_3331);
nand U8752 (N_8752,N_3279,N_4392);
nor U8753 (N_8753,N_4491,N_5710);
nand U8754 (N_8754,N_4260,N_5847);
nor U8755 (N_8755,N_3845,N_5628);
or U8756 (N_8756,N_4798,N_5273);
and U8757 (N_8757,N_4329,N_5864);
or U8758 (N_8758,N_3668,N_4379);
and U8759 (N_8759,N_3406,N_3671);
or U8760 (N_8760,N_3944,N_5076);
nand U8761 (N_8761,N_4415,N_3546);
or U8762 (N_8762,N_5852,N_4125);
or U8763 (N_8763,N_5973,N_3208);
nor U8764 (N_8764,N_4017,N_4508);
nor U8765 (N_8765,N_3600,N_4222);
nor U8766 (N_8766,N_4654,N_4880);
or U8767 (N_8767,N_3645,N_5602);
nor U8768 (N_8768,N_5992,N_5095);
xnor U8769 (N_8769,N_3856,N_4101);
and U8770 (N_8770,N_3699,N_5421);
nand U8771 (N_8771,N_4626,N_3291);
nand U8772 (N_8772,N_5888,N_5380);
nand U8773 (N_8773,N_3604,N_5749);
and U8774 (N_8774,N_5476,N_4580);
nand U8775 (N_8775,N_3158,N_4382);
nor U8776 (N_8776,N_5359,N_4114);
nor U8777 (N_8777,N_5570,N_3221);
nor U8778 (N_8778,N_5309,N_3181);
nor U8779 (N_8779,N_5251,N_4850);
and U8780 (N_8780,N_4263,N_4322);
and U8781 (N_8781,N_3847,N_3779);
or U8782 (N_8782,N_5917,N_3072);
or U8783 (N_8783,N_3001,N_4341);
nand U8784 (N_8784,N_4986,N_5371);
and U8785 (N_8785,N_5575,N_4604);
or U8786 (N_8786,N_3770,N_4333);
nand U8787 (N_8787,N_3151,N_5681);
nor U8788 (N_8788,N_5145,N_5718);
or U8789 (N_8789,N_4552,N_3455);
nor U8790 (N_8790,N_3346,N_4087);
or U8791 (N_8791,N_5671,N_5779);
or U8792 (N_8792,N_4483,N_4165);
nor U8793 (N_8793,N_4585,N_5588);
and U8794 (N_8794,N_3263,N_5308);
and U8795 (N_8795,N_4572,N_5182);
nor U8796 (N_8796,N_5028,N_4124);
and U8797 (N_8797,N_4099,N_3530);
xnor U8798 (N_8798,N_4801,N_3637);
and U8799 (N_8799,N_5481,N_4509);
or U8800 (N_8800,N_4724,N_4941);
and U8801 (N_8801,N_4927,N_4356);
nand U8802 (N_8802,N_5546,N_5442);
or U8803 (N_8803,N_4759,N_4997);
and U8804 (N_8804,N_4800,N_4370);
nand U8805 (N_8805,N_4295,N_3828);
nor U8806 (N_8806,N_5339,N_3952);
nor U8807 (N_8807,N_4371,N_3378);
nor U8808 (N_8808,N_4872,N_4552);
nand U8809 (N_8809,N_4175,N_4156);
nand U8810 (N_8810,N_5023,N_3006);
or U8811 (N_8811,N_4224,N_5771);
nand U8812 (N_8812,N_5159,N_3719);
or U8813 (N_8813,N_5854,N_5074);
or U8814 (N_8814,N_5895,N_3890);
nor U8815 (N_8815,N_4982,N_4829);
and U8816 (N_8816,N_5143,N_3643);
and U8817 (N_8817,N_3358,N_3012);
nor U8818 (N_8818,N_5253,N_5909);
or U8819 (N_8819,N_5974,N_3531);
nor U8820 (N_8820,N_3890,N_5612);
and U8821 (N_8821,N_5923,N_5827);
nand U8822 (N_8822,N_4173,N_5274);
and U8823 (N_8823,N_4017,N_5812);
nor U8824 (N_8824,N_4348,N_3529);
or U8825 (N_8825,N_5963,N_3981);
nand U8826 (N_8826,N_3079,N_3567);
nor U8827 (N_8827,N_3365,N_3899);
and U8828 (N_8828,N_5044,N_3214);
and U8829 (N_8829,N_4088,N_5513);
nor U8830 (N_8830,N_3008,N_4687);
xor U8831 (N_8831,N_4962,N_4467);
or U8832 (N_8832,N_5132,N_4117);
or U8833 (N_8833,N_4648,N_5261);
xnor U8834 (N_8834,N_5439,N_4562);
nand U8835 (N_8835,N_5412,N_4175);
and U8836 (N_8836,N_3667,N_3173);
nand U8837 (N_8837,N_4201,N_5735);
or U8838 (N_8838,N_5400,N_5762);
or U8839 (N_8839,N_5725,N_5659);
nand U8840 (N_8840,N_3906,N_5141);
nor U8841 (N_8841,N_5749,N_3011);
and U8842 (N_8842,N_3475,N_4184);
nor U8843 (N_8843,N_5822,N_3622);
nor U8844 (N_8844,N_5920,N_3578);
nand U8845 (N_8845,N_3587,N_5211);
and U8846 (N_8846,N_5399,N_5855);
nand U8847 (N_8847,N_3241,N_5129);
or U8848 (N_8848,N_3556,N_4142);
and U8849 (N_8849,N_3938,N_5904);
nand U8850 (N_8850,N_5030,N_4642);
nand U8851 (N_8851,N_3343,N_4013);
and U8852 (N_8852,N_4895,N_4629);
or U8853 (N_8853,N_5873,N_5181);
and U8854 (N_8854,N_5002,N_4359);
or U8855 (N_8855,N_3976,N_5704);
nand U8856 (N_8856,N_5950,N_5356);
or U8857 (N_8857,N_3346,N_4090);
or U8858 (N_8858,N_4517,N_4721);
and U8859 (N_8859,N_3797,N_5723);
nor U8860 (N_8860,N_3196,N_5712);
nor U8861 (N_8861,N_3887,N_4192);
and U8862 (N_8862,N_3046,N_5202);
nor U8863 (N_8863,N_4158,N_4312);
or U8864 (N_8864,N_3022,N_5010);
and U8865 (N_8865,N_5220,N_4568);
and U8866 (N_8866,N_4665,N_5125);
and U8867 (N_8867,N_4710,N_5309);
nor U8868 (N_8868,N_3243,N_5032);
nor U8869 (N_8869,N_3924,N_3035);
nor U8870 (N_8870,N_4567,N_3521);
or U8871 (N_8871,N_4802,N_5560);
and U8872 (N_8872,N_5901,N_3399);
nand U8873 (N_8873,N_5666,N_4514);
or U8874 (N_8874,N_5283,N_5372);
and U8875 (N_8875,N_4126,N_4346);
nand U8876 (N_8876,N_3322,N_4587);
nand U8877 (N_8877,N_5762,N_4938);
nand U8878 (N_8878,N_5244,N_3462);
nand U8879 (N_8879,N_3981,N_3502);
and U8880 (N_8880,N_4992,N_4243);
and U8881 (N_8881,N_4899,N_4585);
or U8882 (N_8882,N_5698,N_5513);
or U8883 (N_8883,N_5816,N_5595);
or U8884 (N_8884,N_5787,N_3914);
nand U8885 (N_8885,N_3362,N_4108);
nand U8886 (N_8886,N_5153,N_4238);
or U8887 (N_8887,N_5706,N_4460);
or U8888 (N_8888,N_5442,N_4904);
nand U8889 (N_8889,N_4595,N_5426);
or U8890 (N_8890,N_5693,N_4089);
nand U8891 (N_8891,N_5558,N_5140);
and U8892 (N_8892,N_4996,N_3082);
nand U8893 (N_8893,N_3625,N_5443);
or U8894 (N_8894,N_5979,N_3298);
nand U8895 (N_8895,N_5803,N_3044);
nor U8896 (N_8896,N_3558,N_3019);
nor U8897 (N_8897,N_3525,N_5958);
and U8898 (N_8898,N_5153,N_4317);
and U8899 (N_8899,N_4546,N_5332);
nor U8900 (N_8900,N_5243,N_3005);
and U8901 (N_8901,N_4613,N_5533);
nor U8902 (N_8902,N_4272,N_4678);
or U8903 (N_8903,N_4841,N_5827);
nand U8904 (N_8904,N_3360,N_5955);
xor U8905 (N_8905,N_5323,N_4448);
or U8906 (N_8906,N_5230,N_5828);
nor U8907 (N_8907,N_4305,N_5025);
and U8908 (N_8908,N_4509,N_5963);
or U8909 (N_8909,N_4237,N_3208);
nand U8910 (N_8910,N_5842,N_5708);
or U8911 (N_8911,N_3078,N_4055);
nand U8912 (N_8912,N_5854,N_3720);
or U8913 (N_8913,N_5906,N_4059);
nand U8914 (N_8914,N_3350,N_4117);
and U8915 (N_8915,N_3566,N_3986);
or U8916 (N_8916,N_4427,N_4445);
and U8917 (N_8917,N_4243,N_4102);
nand U8918 (N_8918,N_3726,N_4008);
nor U8919 (N_8919,N_5809,N_3846);
nand U8920 (N_8920,N_4302,N_3368);
or U8921 (N_8921,N_3764,N_5304);
and U8922 (N_8922,N_4408,N_4641);
or U8923 (N_8923,N_3134,N_5386);
nand U8924 (N_8924,N_4435,N_5965);
or U8925 (N_8925,N_3860,N_4928);
and U8926 (N_8926,N_5997,N_3559);
and U8927 (N_8927,N_4139,N_3523);
nand U8928 (N_8928,N_4211,N_5211);
and U8929 (N_8929,N_4757,N_5363);
nor U8930 (N_8930,N_5060,N_3820);
nor U8931 (N_8931,N_5113,N_5065);
nor U8932 (N_8932,N_5879,N_4438);
and U8933 (N_8933,N_5146,N_4024);
nor U8934 (N_8934,N_3651,N_3007);
or U8935 (N_8935,N_4963,N_5861);
nor U8936 (N_8936,N_4416,N_3434);
or U8937 (N_8937,N_3895,N_3989);
nand U8938 (N_8938,N_4767,N_4653);
or U8939 (N_8939,N_4302,N_3510);
and U8940 (N_8940,N_5272,N_5696);
nand U8941 (N_8941,N_3893,N_5614);
nor U8942 (N_8942,N_4462,N_3460);
and U8943 (N_8943,N_4271,N_5043);
xor U8944 (N_8944,N_3180,N_3101);
or U8945 (N_8945,N_5872,N_3883);
nor U8946 (N_8946,N_4524,N_3429);
nand U8947 (N_8947,N_5939,N_3053);
nor U8948 (N_8948,N_4229,N_3598);
nor U8949 (N_8949,N_5728,N_5653);
nand U8950 (N_8950,N_5749,N_5988);
or U8951 (N_8951,N_5195,N_3299);
nor U8952 (N_8952,N_3996,N_5420);
or U8953 (N_8953,N_5098,N_5355);
nor U8954 (N_8954,N_5123,N_5216);
nand U8955 (N_8955,N_3934,N_3345);
or U8956 (N_8956,N_4244,N_5205);
nand U8957 (N_8957,N_3990,N_4974);
or U8958 (N_8958,N_4163,N_5003);
nand U8959 (N_8959,N_4326,N_5285);
nand U8960 (N_8960,N_4131,N_3297);
xor U8961 (N_8961,N_5619,N_3117);
or U8962 (N_8962,N_3168,N_4494);
or U8963 (N_8963,N_5353,N_3058);
nor U8964 (N_8964,N_3035,N_3966);
and U8965 (N_8965,N_4484,N_3432);
and U8966 (N_8966,N_5315,N_4400);
or U8967 (N_8967,N_5890,N_4493);
nand U8968 (N_8968,N_3037,N_5695);
nand U8969 (N_8969,N_4597,N_5743);
nor U8970 (N_8970,N_4054,N_4802);
or U8971 (N_8971,N_4287,N_5495);
and U8972 (N_8972,N_5477,N_4837);
or U8973 (N_8973,N_3370,N_3413);
or U8974 (N_8974,N_4133,N_4231);
and U8975 (N_8975,N_5515,N_5469);
nor U8976 (N_8976,N_3678,N_3500);
or U8977 (N_8977,N_4701,N_3059);
nor U8978 (N_8978,N_5580,N_3639);
or U8979 (N_8979,N_3492,N_4802);
or U8980 (N_8980,N_5744,N_5139);
nor U8981 (N_8981,N_4676,N_4946);
and U8982 (N_8982,N_3978,N_5744);
or U8983 (N_8983,N_4583,N_5649);
and U8984 (N_8984,N_3008,N_3066);
or U8985 (N_8985,N_5671,N_5515);
nand U8986 (N_8986,N_5372,N_3109);
nor U8987 (N_8987,N_3242,N_3457);
and U8988 (N_8988,N_4761,N_4454);
nor U8989 (N_8989,N_4479,N_4113);
xor U8990 (N_8990,N_4478,N_3205);
or U8991 (N_8991,N_4530,N_4264);
or U8992 (N_8992,N_5057,N_4725);
nand U8993 (N_8993,N_5832,N_4898);
or U8994 (N_8994,N_3276,N_4369);
and U8995 (N_8995,N_4035,N_5221);
or U8996 (N_8996,N_4297,N_4615);
nor U8997 (N_8997,N_5359,N_3560);
nor U8998 (N_8998,N_4518,N_4163);
nor U8999 (N_8999,N_4096,N_5155);
or U9000 (N_9000,N_7723,N_7856);
or U9001 (N_9001,N_6321,N_8047);
or U9002 (N_9002,N_7400,N_7460);
and U9003 (N_9003,N_6507,N_6501);
or U9004 (N_9004,N_6368,N_7434);
and U9005 (N_9005,N_8884,N_6740);
xnor U9006 (N_9006,N_8715,N_8962);
xor U9007 (N_9007,N_8459,N_7002);
or U9008 (N_9008,N_6620,N_8313);
xor U9009 (N_9009,N_7672,N_6743);
nor U9010 (N_9010,N_7521,N_6908);
nor U9011 (N_9011,N_6296,N_7687);
nand U9012 (N_9012,N_7755,N_6162);
or U9013 (N_9013,N_7817,N_6253);
nor U9014 (N_9014,N_7603,N_7668);
nor U9015 (N_9015,N_6880,N_6491);
or U9016 (N_9016,N_7335,N_6544);
nor U9017 (N_9017,N_8049,N_8839);
xnor U9018 (N_9018,N_6338,N_7777);
and U9019 (N_9019,N_8833,N_8145);
or U9020 (N_9020,N_6808,N_7653);
nand U9021 (N_9021,N_8229,N_8285);
and U9022 (N_9022,N_7669,N_7609);
or U9023 (N_9023,N_8099,N_8955);
or U9024 (N_9024,N_8795,N_8353);
nand U9025 (N_9025,N_6900,N_6746);
xnor U9026 (N_9026,N_6647,N_7313);
or U9027 (N_9027,N_8944,N_8464);
or U9028 (N_9028,N_8129,N_8395);
nor U9029 (N_9029,N_6514,N_8873);
nand U9030 (N_9030,N_7916,N_8548);
and U9031 (N_9031,N_6856,N_6502);
nor U9032 (N_9032,N_6875,N_7206);
or U9033 (N_9033,N_8069,N_6371);
or U9034 (N_9034,N_6631,N_8429);
and U9035 (N_9035,N_8078,N_6707);
or U9036 (N_9036,N_7955,N_7488);
xor U9037 (N_9037,N_6166,N_8384);
nand U9038 (N_9038,N_8860,N_6086);
or U9039 (N_9039,N_6582,N_8478);
nor U9040 (N_9040,N_8294,N_7592);
nand U9041 (N_9041,N_8139,N_6661);
and U9042 (N_9042,N_8851,N_6776);
nand U9043 (N_9043,N_6285,N_6054);
xor U9044 (N_9044,N_8045,N_7052);
nand U9045 (N_9045,N_8472,N_8142);
or U9046 (N_9046,N_8607,N_8678);
nor U9047 (N_9047,N_6873,N_8787);
or U9048 (N_9048,N_6609,N_7486);
nor U9049 (N_9049,N_8956,N_6536);
xnor U9050 (N_9050,N_8874,N_6072);
nor U9051 (N_9051,N_7062,N_7977);
nand U9052 (N_9052,N_7204,N_7041);
nor U9053 (N_9053,N_7617,N_7732);
nand U9054 (N_9054,N_6018,N_8543);
nand U9055 (N_9055,N_7815,N_6734);
nand U9056 (N_9056,N_6560,N_7143);
nand U9057 (N_9057,N_6251,N_6576);
nand U9058 (N_9058,N_7138,N_7898);
or U9059 (N_9059,N_7957,N_8183);
nor U9060 (N_9060,N_7374,N_8112);
nor U9061 (N_9061,N_6630,N_8519);
nor U9062 (N_9062,N_8743,N_6598);
nand U9063 (N_9063,N_7824,N_6322);
or U9064 (N_9064,N_8714,N_8209);
nand U9065 (N_9065,N_6845,N_8578);
and U9066 (N_9066,N_8669,N_8486);
nor U9067 (N_9067,N_7993,N_8156);
or U9068 (N_9068,N_7185,N_8950);
nor U9069 (N_9069,N_6958,N_6279);
or U9070 (N_9070,N_8193,N_8257);
or U9071 (N_9071,N_7330,N_6813);
nand U9072 (N_9072,N_8273,N_8906);
or U9073 (N_9073,N_8565,N_7667);
nand U9074 (N_9074,N_8402,N_6174);
and U9075 (N_9075,N_7031,N_6624);
nand U9076 (N_9076,N_7380,N_8122);
nor U9077 (N_9077,N_7548,N_6033);
nand U9078 (N_9078,N_8485,N_7741);
nand U9079 (N_9079,N_7579,N_8992);
nand U9080 (N_9080,N_8627,N_8586);
or U9081 (N_9081,N_7432,N_6876);
nand U9082 (N_9082,N_7249,N_8428);
nor U9083 (N_9083,N_8938,N_8502);
or U9084 (N_9084,N_7889,N_6983);
or U9085 (N_9085,N_6613,N_6764);
nand U9086 (N_9086,N_8601,N_8298);
nor U9087 (N_9087,N_7446,N_8076);
nor U9088 (N_9088,N_8721,N_8290);
and U9089 (N_9089,N_6099,N_7768);
and U9090 (N_9090,N_8904,N_7226);
nor U9091 (N_9091,N_6870,N_7492);
nand U9092 (N_9092,N_8375,N_7282);
nor U9093 (N_9093,N_8660,N_6542);
nor U9094 (N_9094,N_8497,N_7244);
or U9095 (N_9095,N_7019,N_7343);
nand U9096 (N_9096,N_8687,N_8708);
or U9097 (N_9097,N_7612,N_6461);
and U9098 (N_9098,N_6556,N_7716);
or U9099 (N_9099,N_6244,N_8501);
nand U9100 (N_9100,N_8406,N_7053);
and U9101 (N_9101,N_7212,N_7149);
nand U9102 (N_9102,N_6658,N_6030);
nor U9103 (N_9103,N_7463,N_7262);
nor U9104 (N_9104,N_6653,N_8797);
and U9105 (N_9105,N_7406,N_8405);
nor U9106 (N_9106,N_6111,N_6546);
and U9107 (N_9107,N_8657,N_6710);
nand U9108 (N_9108,N_7284,N_6325);
or U9109 (N_9109,N_7046,N_8283);
nand U9110 (N_9110,N_6170,N_8576);
nand U9111 (N_9111,N_8799,N_8400);
nand U9112 (N_9112,N_7231,N_7736);
nor U9113 (N_9113,N_7674,N_6021);
or U9114 (N_9114,N_6597,N_6668);
or U9115 (N_9115,N_6747,N_7583);
nor U9116 (N_9116,N_7537,N_6574);
or U9117 (N_9117,N_6906,N_8180);
or U9118 (N_9118,N_7725,N_6646);
nand U9119 (N_9119,N_7342,N_6401);
nor U9120 (N_9120,N_7575,N_8506);
nor U9121 (N_9121,N_8677,N_8408);
and U9122 (N_9122,N_8963,N_6123);
or U9123 (N_9123,N_8132,N_8954);
or U9124 (N_9124,N_7851,N_8976);
nand U9125 (N_9125,N_7597,N_6976);
nor U9126 (N_9126,N_6588,N_6329);
xnor U9127 (N_9127,N_6423,N_8133);
and U9128 (N_9128,N_8986,N_7152);
or U9129 (N_9129,N_7742,N_8095);
nor U9130 (N_9130,N_6798,N_8568);
or U9131 (N_9131,N_7169,N_8067);
and U9132 (N_9132,N_8512,N_8218);
or U9133 (N_9133,N_8786,N_8882);
and U9134 (N_9134,N_7219,N_6636);
and U9135 (N_9135,N_8325,N_7784);
and U9136 (N_9136,N_7666,N_7357);
nand U9137 (N_9137,N_8410,N_7347);
nand U9138 (N_9138,N_6381,N_8516);
nand U9139 (N_9139,N_7100,N_6009);
nand U9140 (N_9140,N_7810,N_6896);
nor U9141 (N_9141,N_6828,N_7345);
xor U9142 (N_9142,N_7904,N_7436);
or U9143 (N_9143,N_8999,N_8965);
or U9144 (N_9144,N_8547,N_8612);
nor U9145 (N_9145,N_7264,N_8302);
xnor U9146 (N_9146,N_8811,N_8108);
and U9147 (N_9147,N_8086,N_8206);
or U9148 (N_9148,N_7141,N_7252);
and U9149 (N_9149,N_6224,N_8018);
nor U9150 (N_9150,N_7506,N_7084);
nand U9151 (N_9151,N_6012,N_6672);
nand U9152 (N_9152,N_6727,N_7442);
nand U9153 (N_9153,N_7620,N_7229);
nor U9154 (N_9154,N_8379,N_8017);
nand U9155 (N_9155,N_8979,N_8054);
or U9156 (N_9156,N_7168,N_8726);
nor U9157 (N_9157,N_6935,N_6071);
or U9158 (N_9158,N_7491,N_7936);
nand U9159 (N_9159,N_8367,N_8631);
nand U9160 (N_9160,N_7268,N_8261);
nor U9161 (N_9161,N_7361,N_6477);
nor U9162 (N_9162,N_7386,N_8028);
nor U9163 (N_9163,N_6871,N_6284);
or U9164 (N_9164,N_7108,N_6551);
nor U9165 (N_9165,N_8026,N_6185);
and U9166 (N_9166,N_8235,N_6211);
or U9167 (N_9167,N_7241,N_7847);
or U9168 (N_9168,N_8900,N_6150);
nor U9169 (N_9169,N_6708,N_7502);
or U9170 (N_9170,N_7594,N_7207);
or U9171 (N_9171,N_8037,N_7806);
nand U9172 (N_9172,N_6104,N_7140);
or U9173 (N_9173,N_8850,N_6252);
nand U9174 (N_9174,N_8838,N_7399);
nand U9175 (N_9175,N_8424,N_6226);
nand U9176 (N_9176,N_8117,N_8197);
or U9177 (N_9177,N_6290,N_6261);
and U9178 (N_9178,N_6923,N_6392);
or U9179 (N_9179,N_7863,N_8010);
nor U9180 (N_9180,N_8724,N_7376);
and U9181 (N_9181,N_8185,N_6519);
nor U9182 (N_9182,N_7327,N_7907);
or U9183 (N_9183,N_7981,N_7584);
nand U9184 (N_9184,N_8255,N_8058);
nor U9185 (N_9185,N_8236,N_8341);
or U9186 (N_9186,N_6677,N_8897);
nand U9187 (N_9187,N_6266,N_7448);
nand U9188 (N_9188,N_8899,N_6725);
nand U9189 (N_9189,N_8339,N_6336);
nand U9190 (N_9190,N_6769,N_7726);
nand U9191 (N_9191,N_7490,N_6910);
nand U9192 (N_9192,N_8659,N_7799);
or U9193 (N_9193,N_6070,N_8414);
and U9194 (N_9194,N_7180,N_8263);
or U9195 (N_9195,N_6079,N_8618);
or U9196 (N_9196,N_6402,N_8905);
and U9197 (N_9197,N_8694,N_7711);
nand U9198 (N_9198,N_7378,N_8534);
or U9199 (N_9199,N_6549,N_7004);
and U9200 (N_9200,N_6892,N_7980);
and U9201 (N_9201,N_8808,N_8286);
nand U9202 (N_9202,N_6874,N_8705);
or U9203 (N_9203,N_7297,N_6289);
or U9204 (N_9204,N_8447,N_8048);
nand U9205 (N_9205,N_8865,N_7882);
nand U9206 (N_9206,N_7155,N_6859);
nand U9207 (N_9207,N_7901,N_7960);
xnor U9208 (N_9208,N_8613,N_7025);
nand U9209 (N_9209,N_6530,N_6245);
nor U9210 (N_9210,N_6116,N_7765);
nand U9211 (N_9211,N_6890,N_8785);
nand U9212 (N_9212,N_8373,N_8239);
nand U9213 (N_9213,N_7568,N_7308);
nor U9214 (N_9214,N_8426,N_7976);
nand U9215 (N_9215,N_6554,N_6353);
nand U9216 (N_9216,N_7033,N_6787);
nand U9217 (N_9217,N_7582,N_6596);
nor U9218 (N_9218,N_6215,N_8973);
nor U9219 (N_9219,N_7929,N_6748);
and U9220 (N_9220,N_7999,N_6988);
and U9221 (N_9221,N_7091,N_7841);
and U9222 (N_9222,N_6623,N_6424);
nand U9223 (N_9223,N_8052,N_6805);
xor U9224 (N_9224,N_6411,N_7050);
and U9225 (N_9225,N_8902,N_8064);
nand U9226 (N_9226,N_6911,N_8583);
nand U9227 (N_9227,N_6573,N_6967);
and U9228 (N_9228,N_6745,N_7385);
or U9229 (N_9229,N_8883,N_6693);
nor U9230 (N_9230,N_8075,N_8598);
nand U9231 (N_9231,N_7469,N_8893);
nand U9232 (N_9232,N_8242,N_6075);
and U9233 (N_9233,N_8019,N_8822);
or U9234 (N_9234,N_7626,N_6173);
nor U9235 (N_9235,N_7278,N_6818);
nand U9236 (N_9236,N_7555,N_6248);
or U9237 (N_9237,N_8179,N_7748);
and U9238 (N_9238,N_8836,N_6991);
nor U9239 (N_9239,N_6102,N_8317);
nand U9240 (N_9240,N_7382,N_8396);
nor U9241 (N_9241,N_7767,N_7074);
and U9242 (N_9242,N_8378,N_7466);
and U9243 (N_9243,N_6893,N_6201);
nor U9244 (N_9244,N_7018,N_8166);
nor U9245 (N_9245,N_8957,N_6840);
and U9246 (N_9246,N_8605,N_7228);
nor U9247 (N_9247,N_8066,N_6548);
or U9248 (N_9248,N_6050,N_7247);
nand U9249 (N_9249,N_7415,N_6816);
nor U9250 (N_9250,N_6295,N_6699);
nor U9251 (N_9251,N_7833,N_6789);
nand U9252 (N_9252,N_7402,N_8796);
or U9253 (N_9253,N_8352,N_8932);
nand U9254 (N_9254,N_6420,N_8127);
or U9255 (N_9255,N_8903,N_8024);
nor U9256 (N_9256,N_6704,N_6815);
and U9257 (N_9257,N_6056,N_6168);
nand U9258 (N_9258,N_6685,N_8668);
or U9259 (N_9259,N_8460,N_7187);
and U9260 (N_9260,N_6367,N_7699);
nor U9261 (N_9261,N_6339,N_7360);
nand U9262 (N_9262,N_7321,N_6124);
or U9263 (N_9263,N_8461,N_7828);
and U9264 (N_9264,N_6024,N_6651);
and U9265 (N_9265,N_6333,N_7042);
or U9266 (N_9266,N_7937,N_6243);
xor U9267 (N_9267,N_8182,N_7307);
or U9268 (N_9268,N_7472,N_6905);
nand U9269 (N_9269,N_8879,N_7899);
and U9270 (N_9270,N_6087,N_7288);
and U9271 (N_9271,N_6872,N_7704);
and U9272 (N_9272,N_7158,N_8602);
and U9273 (N_9273,N_7835,N_8432);
and U9274 (N_9274,N_7776,N_7362);
nand U9275 (N_9275,N_7494,N_8374);
and U9276 (N_9276,N_8187,N_7334);
or U9277 (N_9277,N_6853,N_7498);
nor U9278 (N_9278,N_7997,N_6852);
or U9279 (N_9279,N_7163,N_7484);
and U9280 (N_9280,N_7632,N_8642);
and U9281 (N_9281,N_8764,N_8157);
and U9282 (N_9282,N_8274,N_6493);
nand U9283 (N_9283,N_6943,N_7173);
nor U9284 (N_9284,N_7263,N_6221);
or U9285 (N_9285,N_7786,N_7596);
nand U9286 (N_9286,N_8720,N_8337);
or U9287 (N_9287,N_6616,N_6092);
nor U9288 (N_9288,N_8380,N_7410);
nor U9289 (N_9289,N_8713,N_7827);
and U9290 (N_9290,N_8362,N_7026);
nor U9291 (N_9291,N_8262,N_7565);
nor U9292 (N_9292,N_8253,N_6006);
nand U9293 (N_9293,N_8890,N_6214);
nand U9294 (N_9294,N_6254,N_7005);
or U9295 (N_9295,N_6378,N_7554);
xor U9296 (N_9296,N_6755,N_8923);
or U9297 (N_9297,N_6825,N_8173);
nand U9298 (N_9298,N_8710,N_8589);
nor U9299 (N_9299,N_8991,N_8043);
nand U9300 (N_9300,N_8469,N_8087);
and U9301 (N_9301,N_7785,N_7805);
and U9302 (N_9302,N_6439,N_6532);
nand U9303 (N_9303,N_6343,N_6965);
nor U9304 (N_9304,N_8441,N_6361);
or U9305 (N_9305,N_7395,N_8935);
xnor U9306 (N_9306,N_6912,N_7633);
and U9307 (N_9307,N_6529,N_8840);
and U9308 (N_9308,N_6823,N_8933);
and U9309 (N_9309,N_8105,N_7202);
or U9310 (N_9310,N_8587,N_7932);
nand U9311 (N_9311,N_6144,N_6063);
or U9312 (N_9312,N_8719,N_7057);
and U9313 (N_9313,N_7465,N_7266);
or U9314 (N_9314,N_8161,N_7645);
nand U9315 (N_9315,N_7095,N_7496);
nand U9316 (N_9316,N_7552,N_6806);
nand U9317 (N_9317,N_8824,N_7728);
and U9318 (N_9318,N_8969,N_7192);
nor U9319 (N_9319,N_7707,N_6637);
nand U9320 (N_9320,N_7538,N_7855);
nor U9321 (N_9321,N_8224,N_6267);
and U9322 (N_9322,N_7299,N_6213);
nor U9323 (N_9323,N_8617,N_7607);
nand U9324 (N_9324,N_8059,N_8031);
xor U9325 (N_9325,N_6971,N_8513);
or U9326 (N_9326,N_6652,N_7341);
nor U9327 (N_9327,N_6895,N_8967);
nand U9328 (N_9328,N_8919,N_8503);
nand U9329 (N_9329,N_6257,N_7943);
or U9330 (N_9330,N_7700,N_7822);
and U9331 (N_9331,N_6639,N_7069);
and U9332 (N_9332,N_8011,N_6113);
nand U9333 (N_9333,N_6085,N_6278);
nor U9334 (N_9334,N_6434,N_6899);
nand U9335 (N_9335,N_7339,N_8296);
nor U9336 (N_9336,N_8388,N_7706);
nor U9337 (N_9337,N_7877,N_8149);
nand U9338 (N_9338,N_6671,N_6472);
and U9339 (N_9339,N_8843,N_6418);
or U9340 (N_9340,N_8141,N_8080);
nor U9341 (N_9341,N_6946,N_7780);
nor U9342 (N_9342,N_6930,N_7920);
and U9343 (N_9343,N_8763,N_6122);
nor U9344 (N_9344,N_8901,N_8636);
and U9345 (N_9345,N_7639,N_7227);
nor U9346 (N_9346,N_6632,N_8403);
and U9347 (N_9347,N_6467,N_8434);
nand U9348 (N_9348,N_6781,N_8837);
nor U9349 (N_9349,N_7998,N_6719);
or U9350 (N_9350,N_6494,N_7523);
or U9351 (N_9351,N_7778,N_8077);
or U9352 (N_9352,N_7517,N_7974);
and U9353 (N_9353,N_8091,N_6002);
or U9354 (N_9354,N_7203,N_8155);
and U9355 (N_9355,N_7516,N_7329);
nand U9356 (N_9356,N_6810,N_6476);
nor U9357 (N_9357,N_7946,N_8752);
nor U9358 (N_9358,N_7935,N_6028);
nor U9359 (N_9359,N_7979,N_8409);
nor U9360 (N_9360,N_8742,N_6388);
nand U9361 (N_9361,N_6058,N_8347);
or U9362 (N_9362,N_8744,N_7606);
nand U9363 (N_9363,N_6604,N_7894);
nor U9364 (N_9364,N_6008,N_8126);
or U9365 (N_9365,N_6280,N_8344);
and U9366 (N_9366,N_6005,N_6688);
nor U9367 (N_9367,N_8765,N_7846);
and U9368 (N_9368,N_7743,N_6406);
or U9369 (N_9369,N_8623,N_6212);
nor U9370 (N_9370,N_8243,N_6512);
xnor U9371 (N_9371,N_8207,N_6939);
and U9372 (N_9372,N_7353,N_6015);
or U9373 (N_9373,N_7326,N_8648);
or U9374 (N_9374,N_6089,N_7589);
and U9375 (N_9375,N_8237,N_7255);
and U9376 (N_9376,N_6511,N_6200);
or U9377 (N_9377,N_7075,N_6068);
xor U9378 (N_9378,N_8371,N_8098);
and U9379 (N_9379,N_8934,N_7232);
nand U9380 (N_9380,N_7066,N_6902);
nor U9381 (N_9381,N_7838,N_8297);
nor U9382 (N_9382,N_7131,N_8951);
or U9383 (N_9383,N_7948,N_8524);
or U9384 (N_9384,N_8466,N_6394);
and U9385 (N_9385,N_7477,N_6795);
and U9386 (N_9386,N_7428,N_7634);
or U9387 (N_9387,N_6565,N_7029);
nor U9388 (N_9388,N_6679,N_6247);
nand U9389 (N_9389,N_6274,N_7280);
or U9390 (N_9390,N_8171,N_8707);
or U9391 (N_9391,N_7934,N_8119);
or U9392 (N_9392,N_6230,N_7105);
nand U9393 (N_9393,N_7144,N_6959);
nor U9394 (N_9394,N_8684,N_6995);
and U9395 (N_9395,N_8300,N_7099);
or U9396 (N_9396,N_8416,N_6822);
nor U9397 (N_9397,N_6481,N_8540);
nor U9398 (N_9398,N_7349,N_6438);
or U9399 (N_9399,N_7135,N_6466);
nor U9400 (N_9400,N_6383,N_8093);
or U9401 (N_9401,N_8579,N_6114);
nor U9402 (N_9402,N_7971,N_7094);
xnor U9403 (N_9403,N_7735,N_7965);
nor U9404 (N_9404,N_8258,N_6149);
nand U9405 (N_9405,N_6994,N_6429);
and U9406 (N_9406,N_7858,N_7873);
nor U9407 (N_9407,N_7883,N_6419);
nand U9408 (N_9408,N_6619,N_7483);
nor U9409 (N_9409,N_7118,N_6614);
or U9410 (N_9410,N_7174,N_8215);
nor U9411 (N_9411,N_6404,N_6602);
nand U9412 (N_9412,N_6572,N_7081);
and U9413 (N_9413,N_8147,N_6794);
and U9414 (N_9414,N_6240,N_7162);
or U9415 (N_9415,N_8510,N_6134);
xnor U9416 (N_9416,N_6770,N_7549);
nand U9417 (N_9417,N_6633,N_6192);
or U9418 (N_9418,N_7079,N_8681);
or U9419 (N_9419,N_6654,N_6249);
xnor U9420 (N_9420,N_6412,N_8909);
nor U9421 (N_9421,N_8654,N_8329);
nand U9422 (N_9422,N_8174,N_7133);
or U9423 (N_9423,N_7504,N_7709);
and U9424 (N_9424,N_7865,N_8604);
nand U9425 (N_9425,N_6250,N_7664);
or U9426 (N_9426,N_6335,N_7830);
nor U9427 (N_9427,N_7060,N_6276);
nor U9428 (N_9428,N_7273,N_7468);
and U9429 (N_9429,N_8463,N_7317);
or U9430 (N_9430,N_6425,N_7544);
or U9431 (N_9431,N_6780,N_6081);
nor U9432 (N_9432,N_6416,N_8252);
nor U9433 (N_9433,N_8827,N_8495);
and U9434 (N_9434,N_7623,N_8250);
nor U9435 (N_9435,N_6022,N_6327);
nand U9436 (N_9436,N_6158,N_7570);
nor U9437 (N_9437,N_6791,N_7316);
nand U9438 (N_9438,N_6750,N_6753);
nor U9439 (N_9439,N_8413,N_6972);
nor U9440 (N_9440,N_8995,N_8008);
or U9441 (N_9441,N_6506,N_8751);
or U9442 (N_9442,N_7734,N_8556);
and U9443 (N_9443,N_7324,N_7694);
and U9444 (N_9444,N_7323,N_7082);
or U9445 (N_9445,N_6309,N_6666);
or U9446 (N_9446,N_7927,N_6389);
nor U9447 (N_9447,N_7416,N_6348);
and U9448 (N_9448,N_7547,N_8383);
nor U9449 (N_9449,N_8619,N_7186);
nor U9450 (N_9450,N_7121,N_6453);
and U9451 (N_9451,N_7220,N_6038);
or U9452 (N_9452,N_6821,N_6034);
nor U9453 (N_9453,N_6445,N_8136);
xor U9454 (N_9454,N_6978,N_7836);
nand U9455 (N_9455,N_8566,N_8452);
and U9456 (N_9456,N_8729,N_8716);
nor U9457 (N_9457,N_6921,N_8291);
nand U9458 (N_9458,N_6317,N_7104);
nand U9459 (N_9459,N_7677,N_7954);
and U9460 (N_9460,N_8980,N_7119);
nand U9461 (N_9461,N_7610,N_6233);
or U9462 (N_9462,N_7630,N_8662);
nor U9463 (N_9463,N_8104,N_6754);
and U9464 (N_9464,N_8574,N_7783);
nor U9465 (N_9465,N_7514,N_6496);
or U9466 (N_9466,N_8887,N_6711);
or U9467 (N_9467,N_8661,N_8465);
nor U9468 (N_9468,N_8393,N_7950);
and U9469 (N_9469,N_8289,N_6138);
or U9470 (N_9470,N_8153,N_7389);
and U9471 (N_9471,N_7127,N_8399);
nand U9472 (N_9472,N_6964,N_6115);
or U9473 (N_9473,N_8181,N_7720);
nand U9474 (N_9474,N_8816,N_6738);
nor U9475 (N_9475,N_7962,N_6898);
nor U9476 (N_9476,N_6869,N_8738);
nand U9477 (N_9477,N_7921,N_7021);
nand U9478 (N_9478,N_8445,N_6046);
and U9479 (N_9479,N_7276,N_6206);
nor U9480 (N_9480,N_8369,N_8723);
nand U9481 (N_9481,N_8220,N_6771);
nor U9482 (N_9482,N_8484,N_8528);
nand U9483 (N_9483,N_6953,N_7214);
or U9484 (N_9484,N_6013,N_8652);
and U9485 (N_9485,N_8419,N_6128);
nand U9486 (N_9486,N_8682,N_6098);
xor U9487 (N_9487,N_6583,N_6363);
nand U9488 (N_9488,N_7793,N_7283);
or U9489 (N_9489,N_6223,N_8065);
nor U9490 (N_9490,N_7112,N_7065);
nor U9491 (N_9491,N_6760,N_6475);
and U9492 (N_9492,N_6109,N_8312);
or U9493 (N_9493,N_7753,N_6723);
nand U9494 (N_9494,N_8754,N_6205);
nor U9495 (N_9495,N_6273,N_7267);
nand U9496 (N_9496,N_8014,N_6282);
nor U9497 (N_9497,N_7782,N_6497);
xnor U9498 (N_9498,N_6775,N_6178);
or U9499 (N_9499,N_6819,N_8885);
and U9500 (N_9500,N_8522,N_8693);
nor U9501 (N_9501,N_7546,N_6801);
nor U9502 (N_9502,N_8834,N_7642);
and U9503 (N_9503,N_7235,N_7294);
xor U9504 (N_9504,N_8769,N_6431);
and U9505 (N_9505,N_8767,N_6667);
nor U9506 (N_9506,N_7471,N_8022);
and U9507 (N_9507,N_6449,N_6047);
nor U9508 (N_9508,N_7890,N_6696);
and U9509 (N_9509,N_8888,N_8641);
and U9510 (N_9510,N_7184,N_6684);
nor U9511 (N_9511,N_7114,N_6364);
nand U9512 (N_9512,N_6617,N_6426);
or U9513 (N_9513,N_8356,N_6757);
or U9514 (N_9514,N_8404,N_8781);
nand U9515 (N_9515,N_8745,N_8750);
nor U9516 (N_9516,N_6796,N_6868);
nand U9517 (N_9517,N_7256,N_7933);
nand U9518 (N_9518,N_6349,N_7556);
nand U9519 (N_9519,N_8176,N_8167);
or U9520 (N_9520,N_6904,N_6628);
nand U9521 (N_9521,N_8109,N_8348);
and U9522 (N_9522,N_7844,N_6487);
nor U9523 (N_9523,N_8222,N_8386);
or U9524 (N_9524,N_6307,N_7425);
nand U9525 (N_9525,N_7651,N_8740);
and U9526 (N_9526,N_7090,N_8368);
nor U9527 (N_9527,N_7663,N_7985);
nand U9528 (N_9528,N_7132,N_6458);
or U9529 (N_9529,N_7464,N_8223);
nor U9530 (N_9530,N_6175,N_7377);
or U9531 (N_9531,N_6884,N_7422);
nor U9532 (N_9532,N_6713,N_8637);
nand U9533 (N_9533,N_7318,N_6722);
nand U9534 (N_9534,N_7426,N_6809);
and U9535 (N_9535,N_6154,N_7635);
and U9536 (N_9536,N_7172,N_7230);
nor U9537 (N_9537,N_8756,N_6758);
or U9538 (N_9538,N_8895,N_7064);
nand U9539 (N_9539,N_6432,N_8407);
nor U9540 (N_9540,N_6306,N_8162);
xor U9541 (N_9541,N_7745,N_8696);
and U9542 (N_9542,N_8621,N_6025);
nand U9543 (N_9543,N_7569,N_7281);
nand U9544 (N_9544,N_7061,N_6380);
or U9545 (N_9545,N_7246,N_8088);
nand U9546 (N_9546,N_7359,N_6675);
nand U9547 (N_9547,N_8916,N_6059);
or U9548 (N_9548,N_8927,N_8036);
or U9549 (N_9549,N_6398,N_6941);
nor U9550 (N_9550,N_6351,N_8541);
nor U9551 (N_9551,N_8685,N_8354);
and U9552 (N_9552,N_6824,N_8128);
and U9553 (N_9553,N_7242,N_6315);
nand U9554 (N_9554,N_6067,N_8082);
nand U9555 (N_9555,N_7182,N_6379);
or U9556 (N_9556,N_7658,N_6669);
nor U9557 (N_9557,N_8259,N_7224);
nand U9558 (N_9558,N_7608,N_7562);
nand U9559 (N_9559,N_7724,N_6301);
nor U9560 (N_9560,N_6027,N_7271);
nand U9561 (N_9561,N_7915,N_7054);
nand U9562 (N_9562,N_8577,N_8314);
or U9563 (N_9563,N_6594,N_7947);
nand U9564 (N_9564,N_8835,N_6793);
or U9565 (N_9565,N_8195,N_6929);
or U9566 (N_9566,N_7604,N_6026);
and U9567 (N_9567,N_6377,N_6073);
nand U9568 (N_9568,N_7148,N_8913);
or U9569 (N_9569,N_8449,N_8775);
nor U9570 (N_9570,N_8761,N_6485);
and U9571 (N_9571,N_7676,N_7072);
nand U9572 (N_9572,N_7870,N_6462);
nand U9573 (N_9573,N_6907,N_6562);
nand U9574 (N_9574,N_6837,N_6662);
nand U9575 (N_9575,N_7973,N_8034);
or U9576 (N_9576,N_7338,N_8706);
nand U9577 (N_9577,N_8175,N_6914);
nor U9578 (N_9578,N_8757,N_7691);
or U9579 (N_9579,N_8689,N_7431);
or U9580 (N_9580,N_6041,N_7628);
nand U9581 (N_9581,N_7692,N_8355);
nand U9582 (N_9582,N_6897,N_7433);
nand U9583 (N_9583,N_7715,N_7403);
and U9584 (N_9584,N_7394,N_8005);
nand U9585 (N_9585,N_6761,N_6304);
and U9586 (N_9586,N_7150,N_7461);
or U9587 (N_9587,N_7629,N_6762);
or U9588 (N_9588,N_8172,N_8188);
nor U9589 (N_9589,N_7093,N_7411);
nand U9590 (N_9590,N_8338,N_6095);
nor U9591 (N_9591,N_6298,N_6700);
or U9592 (N_9592,N_7098,N_8443);
or U9593 (N_9593,N_8125,N_7011);
and U9594 (N_9594,N_7303,N_7840);
and U9595 (N_9595,N_7578,N_6108);
or U9596 (N_9596,N_8572,N_6706);
and U9597 (N_9597,N_8365,N_8361);
and U9598 (N_9598,N_7908,N_6066);
nor U9599 (N_9599,N_6665,N_7476);
or U9600 (N_9600,N_6016,N_6133);
and U9601 (N_9601,N_6732,N_8514);
nor U9602 (N_9602,N_6865,N_7305);
and U9603 (N_9603,N_6846,N_7982);
xor U9604 (N_9604,N_6934,N_7366);
nand U9605 (N_9605,N_6673,N_8199);
nand U9606 (N_9606,N_6407,N_8411);
nand U9607 (N_9607,N_6839,N_8730);
nand U9608 (N_9608,N_6949,N_6164);
nand U9609 (N_9609,N_8483,N_7087);
nor U9610 (N_9610,N_7986,N_8861);
or U9611 (N_9611,N_7200,N_6830);
or U9612 (N_9612,N_6569,N_7270);
nor U9613 (N_9613,N_7823,N_6470);
and U9614 (N_9614,N_6877,N_8457);
nor U9615 (N_9615,N_6262,N_6397);
nand U9616 (N_9616,N_6374,N_7388);
nor U9617 (N_9617,N_7926,N_6951);
and U9618 (N_9618,N_6563,N_8227);
nor U9619 (N_9619,N_7145,N_8671);
nand U9620 (N_9620,N_6422,N_8309);
nand U9621 (N_9621,N_6169,N_8608);
nor U9622 (N_9622,N_8481,N_8722);
nand U9623 (N_9623,N_6640,N_8658);
nor U9624 (N_9624,N_8479,N_6375);
xor U9625 (N_9625,N_6954,N_7686);
nand U9626 (N_9626,N_7577,N_8326);
nor U9627 (N_9627,N_7938,N_6649);
nor U9628 (N_9628,N_6702,N_6603);
nand U9629 (N_9629,N_7387,N_6850);
nand U9630 (N_9630,N_7287,N_8322);
nand U9631 (N_9631,N_7543,N_8610);
xor U9632 (N_9632,N_7346,N_6468);
or U9633 (N_9633,N_7567,N_8625);
and U9634 (N_9634,N_7797,N_7697);
and U9635 (N_9635,N_7787,N_8530);
nor U9636 (N_9636,N_8869,N_6228);
or U9637 (N_9637,N_6735,N_8591);
nor U9638 (N_9638,N_6324,N_6061);
or U9639 (N_9639,N_8553,N_7038);
xor U9640 (N_9640,N_6650,N_7857);
or U9641 (N_9641,N_6683,N_6681);
or U9642 (N_9642,N_8266,N_6763);
or U9643 (N_9643,N_7146,N_8688);
or U9644 (N_9644,N_8702,N_7627);
and U9645 (N_9645,N_7746,N_8332);
and U9646 (N_9646,N_7447,N_6480);
nand U9647 (N_9647,N_8584,N_8753);
or U9648 (N_9648,N_7237,N_7304);
nand U9649 (N_9649,N_7397,N_8582);
nand U9650 (N_9650,N_6346,N_6945);
nand U9651 (N_9651,N_8462,N_7893);
and U9652 (N_9652,N_7602,N_8168);
nor U9653 (N_9653,N_7801,N_7437);
nor U9654 (N_9654,N_7662,N_8697);
or U9655 (N_9655,N_6557,N_7510);
and U9656 (N_9656,N_6117,N_8287);
and U9657 (N_9657,N_6341,N_8143);
nand U9658 (N_9658,N_7027,N_7319);
nor U9659 (N_9659,N_6355,N_6944);
and U9660 (N_9660,N_6332,N_7153);
or U9661 (N_9661,N_6437,N_7831);
and U9662 (N_9662,N_6608,N_8603);
or U9663 (N_9663,N_7872,N_7111);
and U9664 (N_9664,N_7000,N_6924);
and U9665 (N_9665,N_8918,N_6524);
or U9666 (N_9666,N_8948,N_6302);
nand U9667 (N_9667,N_8831,N_6999);
nor U9668 (N_9668,N_8870,N_8651);
or U9669 (N_9669,N_6405,N_6690);
nand U9670 (N_9670,N_6570,N_6300);
nand U9671 (N_9671,N_7195,N_7218);
nor U9672 (N_9672,N_6832,N_8430);
and U9673 (N_9673,N_7020,N_8985);
nor U9674 (N_9674,N_8438,N_8360);
or U9675 (N_9675,N_6435,N_6990);
nand U9676 (N_9676,N_7798,N_6854);
nor U9677 (N_9677,N_6660,N_8421);
nand U9678 (N_9678,N_6107,N_6834);
nor U9679 (N_9679,N_8952,N_6564);
or U9680 (N_9680,N_6219,N_7449);
or U9681 (N_9681,N_7842,N_6347);
and U9682 (N_9682,N_6486,N_6356);
and U9683 (N_9683,N_7788,N_7265);
nand U9684 (N_9684,N_7680,N_7097);
nor U9685 (N_9685,N_8363,N_7404);
nand U9686 (N_9686,N_7254,N_8439);
nand U9687 (N_9687,N_8268,N_8092);
nand U9688 (N_9688,N_6855,N_7164);
xnor U9689 (N_9689,N_8993,N_7808);
and U9690 (N_9690,N_8789,N_6043);
nand U9691 (N_9691,N_7722,N_8191);
and U9692 (N_9692,N_7564,N_8376);
or U9693 (N_9693,N_7945,N_7102);
or U9694 (N_9694,N_8594,N_7401);
nand U9695 (N_9695,N_8219,N_7429);
nand U9696 (N_9696,N_7541,N_8959);
nor U9697 (N_9697,N_6626,N_7685);
and U9698 (N_9698,N_6091,N_8978);
and U9699 (N_9699,N_7876,N_6227);
nand U9700 (N_9700,N_8390,N_6465);
or U9701 (N_9701,N_7424,N_7931);
and U9702 (N_9702,N_8381,N_8844);
or U9703 (N_9703,N_6790,N_6716);
nor U9704 (N_9704,N_7240,N_7497);
nor U9705 (N_9705,N_6291,N_7679);
nor U9706 (N_9706,N_8046,N_8599);
nor U9707 (N_9707,N_6365,N_7834);
nand U9708 (N_9708,N_6265,N_8813);
nand U9709 (N_9709,N_7994,N_7358);
nand U9710 (N_9710,N_8926,N_8732);
nor U9711 (N_9711,N_8892,N_7532);
or U9712 (N_9712,N_8254,N_6408);
nand U9713 (N_9713,N_8035,N_6436);
nand U9714 (N_9714,N_8025,N_7048);
and U9715 (N_9715,N_6237,N_7275);
or U9716 (N_9716,N_6414,N_7969);
nor U9717 (N_9717,N_6966,N_6137);
and U9718 (N_9718,N_7420,N_8336);
or U9719 (N_9719,N_6430,N_8925);
or U9720 (N_9720,N_7886,N_8232);
and U9721 (N_9721,N_6541,N_8178);
and U9722 (N_9722,N_8002,N_6312);
nand U9723 (N_9723,N_6523,N_6417);
nand U9724 (N_9724,N_8931,N_8392);
nor U9725 (N_9725,N_8009,N_6928);
or U9726 (N_9726,N_6566,N_6578);
nor U9727 (N_9727,N_8943,N_7487);
nand U9728 (N_9728,N_7233,N_7867);
nor U9729 (N_9729,N_8941,N_7209);
and U9730 (N_9730,N_6049,N_6817);
nor U9731 (N_9731,N_8569,N_8056);
nand U9732 (N_9732,N_8759,N_6518);
nor U9733 (N_9733,N_6323,N_7518);
nand U9734 (N_9734,N_8679,N_7729);
nor U9735 (N_9735,N_7712,N_7733);
nor U9736 (N_9736,N_6698,N_8717);
nand U9737 (N_9737,N_7306,N_7191);
and U9738 (N_9738,N_7599,N_7528);
or U9739 (N_9739,N_7816,N_7740);
nor U9740 (N_9740,N_6482,N_7222);
and U9741 (N_9741,N_7440,N_8490);
or U9742 (N_9742,N_6575,N_7077);
and U9743 (N_9743,N_7751,N_7992);
and U9744 (N_9744,N_8271,N_7619);
or U9745 (N_9745,N_8489,N_8804);
nand U9746 (N_9746,N_7804,N_6527);
and U9747 (N_9747,N_8666,N_8690);
nand U9748 (N_9748,N_8946,N_7911);
and U9749 (N_9749,N_8455,N_6313);
nor U9750 (N_9750,N_7078,N_8315);
and U9751 (N_9751,N_8930,N_6064);
nand U9752 (N_9752,N_6386,N_7587);
nand U9753 (N_9753,N_7525,N_8975);
nand U9754 (N_9754,N_8692,N_8864);
nand U9755 (N_9755,N_6866,N_6516);
nor U9756 (N_9756,N_7298,N_6768);
and U9757 (N_9757,N_6993,N_8779);
or U9758 (N_9758,N_6011,N_7479);
nand U9759 (N_9759,N_7453,N_7509);
or U9760 (N_9760,N_7730,N_7441);
nor U9761 (N_9761,N_6894,N_6678);
nor U9762 (N_9762,N_6691,N_7485);
nor U9763 (N_9763,N_7407,N_6784);
xnor U9764 (N_9764,N_8120,N_8225);
and U9765 (N_9765,N_8389,N_6118);
and U9766 (N_9766,N_8012,N_8580);
nand U9767 (N_9767,N_8398,N_8060);
nor U9768 (N_9768,N_6258,N_6093);
nand U9769 (N_9769,N_8545,N_6933);
and U9770 (N_9770,N_8152,N_8282);
nor U9771 (N_9771,N_6318,N_7040);
or U9772 (N_9772,N_8196,N_7561);
and U9773 (N_9773,N_7508,N_8190);
and U9774 (N_9774,N_7325,N_7037);
or U9775 (N_9775,N_7515,N_7930);
or U9776 (N_9776,N_6528,N_8807);
nor U9777 (N_9777,N_7058,N_8101);
or U9778 (N_9778,N_6181,N_7279);
or U9779 (N_9779,N_8845,N_6882);
and U9780 (N_9780,N_6499,N_8032);
nand U9781 (N_9781,N_8245,N_6369);
or U9782 (N_9782,N_6399,N_7665);
nor U9783 (N_9783,N_6590,N_7792);
or U9784 (N_9784,N_6641,N_6997);
nor U9785 (N_9785,N_8343,N_7126);
nand U9786 (N_9786,N_6045,N_8529);
or U9787 (N_9787,N_8907,N_8234);
nand U9788 (N_9788,N_7371,N_8829);
or U9789 (N_9789,N_8819,N_6135);
and U9790 (N_9790,N_6973,N_7731);
nand U9791 (N_9791,N_6326,N_8908);
nand U9792 (N_9792,N_6094,N_7239);
nand U9793 (N_9793,N_8575,N_6826);
nor U9794 (N_9794,N_6709,N_7705);
nor U9795 (N_9795,N_7438,N_8670);
nand U9796 (N_9796,N_8665,N_7968);
or U9797 (N_9797,N_6097,N_8269);
and U9798 (N_9798,N_8358,N_7560);
nand U9799 (N_9799,N_8739,N_6555);
and U9800 (N_9800,N_6695,N_7600);
and U9801 (N_9801,N_6783,N_7533);
nor U9802 (N_9802,N_8015,N_8113);
or U9803 (N_9803,N_7055,N_6889);
nor U9804 (N_9804,N_6052,N_7482);
xor U9805 (N_9805,N_6055,N_7975);
nor U9806 (N_9806,N_8737,N_6558);
xnor U9807 (N_9807,N_6539,N_7194);
nor U9808 (N_9808,N_7795,N_8044);
nand U9809 (N_9809,N_8964,N_6225);
or U9810 (N_9810,N_8782,N_8278);
nand U9811 (N_9811,N_8996,N_6987);
or U9812 (N_9812,N_6161,N_6858);
or U9813 (N_9813,N_8573,N_7673);
or U9814 (N_9814,N_6504,N_7310);
or U9815 (N_9815,N_7320,N_7274);
nand U9816 (N_9816,N_8544,N_7819);
nor U9817 (N_9817,N_7333,N_8345);
nand U9818 (N_9818,N_7176,N_7624);
nand U9819 (N_9819,N_7818,N_7566);
and U9820 (N_9820,N_8020,N_8698);
nor U9821 (N_9821,N_8647,N_7375);
or U9822 (N_9822,N_8562,N_7766);
or U9823 (N_9823,N_8768,N_7085);
nand U9824 (N_9824,N_7124,N_8437);
nor U9825 (N_9825,N_7396,N_8346);
nor U9826 (N_9826,N_7888,N_7843);
nand U9827 (N_9827,N_6644,N_8170);
xnor U9828 (N_9828,N_7875,N_7940);
and U9829 (N_9829,N_6413,N_6292);
nor U9830 (N_9830,N_7861,N_8894);
and U9831 (N_9831,N_6919,N_8492);
nand U9832 (N_9832,N_8815,N_7161);
nor U9833 (N_9833,N_7919,N_7878);
nand U9834 (N_9834,N_8316,N_7719);
nor U9835 (N_9835,N_8803,N_8505);
nand U9836 (N_9836,N_6088,N_7197);
or U9837 (N_9837,N_8448,N_8928);
nor U9838 (N_9838,N_8212,N_8318);
nor U9839 (N_9839,N_7043,N_7573);
and U9840 (N_9840,N_6148,N_8511);
nor U9841 (N_9841,N_7443,N_7703);
nor U9842 (N_9842,N_8794,N_6232);
xnor U9843 (N_9843,N_8792,N_8571);
nor U9844 (N_9844,N_7928,N_6153);
or U9845 (N_9845,N_8971,N_8221);
nand U9846 (N_9846,N_6600,N_7535);
or U9847 (N_9847,N_8791,N_6051);
and U9848 (N_9848,N_6180,N_7571);
or U9849 (N_9849,N_7452,N_7749);
nand U9850 (N_9850,N_8961,N_6177);
and U9851 (N_9851,N_7130,N_6752);
nand U9852 (N_9852,N_7849,N_6172);
nor U9853 (N_9853,N_8814,N_6359);
and U9854 (N_9854,N_6577,N_8736);
nor U9855 (N_9855,N_7590,N_7690);
and U9856 (N_9856,N_8868,N_7638);
or U9857 (N_9857,N_7045,N_7580);
and U9858 (N_9858,N_7614,N_8328);
and U9859 (N_9859,N_6125,N_7201);
and U9860 (N_9860,N_8331,N_7063);
nand U9861 (N_9861,N_7332,N_6131);
and U9862 (N_9862,N_7059,N_7211);
and U9863 (N_9863,N_8867,N_6328);
nand U9864 (N_9864,N_6160,N_8050);
nor U9865 (N_9865,N_8700,N_7737);
or U9866 (N_9866,N_8982,N_7892);
nor U9867 (N_9867,N_8755,N_7671);
nor U9868 (N_9868,N_7277,N_8458);
nand U9869 (N_9869,N_6686,N_8163);
or U9870 (N_9870,N_7134,N_6017);
or U9871 (N_9871,N_8532,N_7171);
or U9872 (N_9872,N_6756,N_7681);
nand U9873 (N_9873,N_6726,N_6974);
nand U9874 (N_9874,N_6042,N_7860);
nor U9875 (N_9875,N_7383,N_8561);
or U9876 (N_9876,N_6982,N_8192);
nor U9877 (N_9877,N_6345,N_6020);
and U9878 (N_9878,N_7880,N_7650);
and U9879 (N_9879,N_6927,N_8981);
nand U9880 (N_9880,N_8100,N_7754);
nand U9881 (N_9881,N_8527,N_7906);
or U9882 (N_9882,N_8194,N_6718);
or U9883 (N_9883,N_7958,N_6152);
or U9884 (N_9884,N_8570,N_7215);
nor U9885 (N_9885,N_8536,N_6851);
nor U9886 (N_9886,N_6729,N_8442);
nor U9887 (N_9887,N_7193,N_6984);
and U9888 (N_9888,N_7129,N_8953);
or U9889 (N_9889,N_8842,N_6663);
or U9890 (N_9890,N_8292,N_8418);
nor U9891 (N_9891,N_8357,N_8788);
and U9892 (N_9892,N_7539,N_8281);
or U9893 (N_9893,N_7103,N_6857);
nand U9894 (N_9894,N_7092,N_8733);
nand U9895 (N_9895,N_7070,N_7221);
nor U9896 (N_9896,N_6489,N_8896);
nor U9897 (N_9897,N_7756,N_6454);
nand U9898 (N_9898,N_6294,N_7874);
nand U9899 (N_9899,N_8453,N_8650);
nor U9900 (N_9900,N_6676,N_6310);
and U9901 (N_9901,N_6080,N_7559);
nand U9902 (N_9902,N_7147,N_7073);
or U9903 (N_9903,N_7372,N_7178);
nand U9904 (N_9904,N_6960,N_7689);
nor U9905 (N_9905,N_6901,N_7588);
xnor U9906 (N_9906,N_7047,N_7991);
nand U9907 (N_9907,N_6004,N_7419);
nor U9908 (N_9908,N_8427,N_6581);
nor U9909 (N_9909,N_7315,N_7845);
nand U9910 (N_9910,N_8284,N_8451);
nand U9911 (N_9911,N_8004,N_6199);
nand U9912 (N_9912,N_6136,N_8686);
nor U9913 (N_9913,N_8310,N_6255);
nand U9914 (N_9914,N_7959,N_6065);
nand U9915 (N_9915,N_8535,N_7285);
and U9916 (N_9916,N_8394,N_8863);
and U9917 (N_9917,N_7478,N_8488);
or U9918 (N_9918,N_6881,N_7949);
nand U9919 (N_9919,N_8085,N_6433);
nand U9920 (N_9920,N_6000,N_6393);
nor U9921 (N_9921,N_7217,N_7450);
nand U9922 (N_9922,N_6035,N_6618);
nand U9923 (N_9923,N_8914,N_7542);
nor U9924 (N_9924,N_6231,N_8123);
or U9925 (N_9925,N_8436,N_7811);
or U9926 (N_9926,N_7576,N_8862);
nand U9927 (N_9927,N_8630,N_6885);
nor U9928 (N_9928,N_6490,N_7897);
or U9929 (N_9929,N_6023,N_7534);
or U9930 (N_9930,N_8810,N_6936);
nand U9931 (N_9931,N_8749,N_8184);
nand U9932 (N_9932,N_7122,N_6084);
nand U9933 (N_9933,N_8244,N_7774);
or U9934 (N_9934,N_6559,N_8859);
nand U9935 (N_9935,N_8683,N_7972);
or U9936 (N_9936,N_6187,N_7340);
or U9937 (N_9937,N_8033,N_6774);
and U9938 (N_9938,N_7368,N_7503);
nand U9939 (N_9939,N_6415,N_8053);
or U9940 (N_9940,N_7839,N_8809);
and U9941 (N_9941,N_6766,N_7825);
and U9942 (N_9942,N_8801,N_7942);
xor U9943 (N_9943,N_7909,N_7154);
nand U9944 (N_9944,N_8307,N_6867);
nor U9945 (N_9945,N_6543,N_8211);
nor U9946 (N_9946,N_6533,N_6299);
xnor U9947 (N_9947,N_7427,N_6344);
or U9948 (N_9948,N_7761,N_6112);
or U9949 (N_9949,N_6330,N_7853);
or U9950 (N_9950,N_6611,N_6440);
or U9951 (N_9951,N_6932,N_6163);
nor U9952 (N_9952,N_7714,N_8997);
nor U9953 (N_9953,N_7044,N_7763);
and U9954 (N_9954,N_8039,N_8475);
and U9955 (N_9955,N_6820,N_7160);
nand U9956 (N_9956,N_6692,N_7136);
and U9957 (N_9957,N_6522,N_7269);
nor U9958 (N_9958,N_6785,N_7762);
nor U9959 (N_9959,N_6105,N_6387);
nand U9960 (N_9960,N_8094,N_7923);
or U9961 (N_9961,N_6337,N_6799);
and U9962 (N_9962,N_6457,N_6442);
nand U9963 (N_9963,N_8597,N_8154);
and U9964 (N_9964,N_7647,N_7128);
nor U9965 (N_9965,N_6772,N_6495);
nor U9966 (N_9966,N_7952,N_7636);
and U9967 (N_9967,N_6441,N_8130);
nor U9968 (N_9968,N_8821,N_6448);
and U9969 (N_9969,N_6395,N_6567);
nor U9970 (N_9970,N_7312,N_7120);
or U9971 (N_9971,N_6447,N_6680);
or U9972 (N_9972,N_6090,N_8301);
and U9973 (N_9973,N_6879,N_6129);
nor U9974 (N_9974,N_7364,N_6985);
and U9975 (N_9975,N_7862,N_8728);
nor U9976 (N_9976,N_7455,N_8063);
nand U9977 (N_9977,N_6931,N_7713);
nand U9978 (N_9978,N_6916,N_8214);
or U9979 (N_9979,N_6587,N_7659);
or U9980 (N_9980,N_7421,N_7314);
nor U9981 (N_9981,N_8111,N_6484);
nor U9982 (N_9982,N_7067,N_6132);
and U9983 (N_9983,N_8264,N_6229);
nor U9984 (N_9984,N_8189,N_6259);
xor U9985 (N_9985,N_7944,N_6271);
nand U9986 (N_9986,N_6372,N_8006);
and U9987 (N_9987,N_8415,N_8872);
nand U9988 (N_9988,N_7675,N_6443);
nor U9989 (N_9989,N_6778,N_6635);
or U9990 (N_9990,N_7641,N_6077);
nor U9991 (N_9991,N_7868,N_6400);
or U9992 (N_9992,N_7536,N_6183);
or U9993 (N_9993,N_8521,N_6209);
and U9994 (N_9994,N_8672,N_7354);
nor U9995 (N_9995,N_7649,N_8013);
or U9996 (N_9996,N_7001,N_7550);
xnor U9997 (N_9997,N_7881,N_7871);
and U9998 (N_9998,N_8027,N_8832);
and U9999 (N_9999,N_8335,N_7190);
nand U10000 (N_10000,N_7922,N_8124);
or U10001 (N_10001,N_8977,N_8910);
nor U10002 (N_10002,N_7682,N_7989);
nor U10003 (N_10003,N_8802,N_6767);
nor U10004 (N_10004,N_7289,N_6540);
or U10005 (N_10005,N_7322,N_7526);
nand U10006 (N_10006,N_8217,N_6208);
nor U10007 (N_10007,N_6926,N_8226);
xnor U10008 (N_10008,N_6842,N_6157);
nand U10009 (N_10009,N_7253,N_7086);
and U10010 (N_10010,N_6739,N_6593);
and U10011 (N_10011,N_8330,N_8062);
or U10012 (N_10012,N_7234,N_7076);
or U10013 (N_10013,N_6110,N_8260);
and U10014 (N_10014,N_6220,N_6744);
and U10015 (N_10015,N_6186,N_8704);
nand U10016 (N_10016,N_7165,N_8551);
nand U10017 (N_10017,N_7336,N_7661);
nand U10018 (N_10018,N_8061,N_8474);
or U10019 (N_10019,N_7771,N_6456);
nand U10020 (N_10020,N_6915,N_7684);
nor U10021 (N_10021,N_6350,N_8151);
nor U10022 (N_10022,N_6642,N_6515);
nand U10023 (N_10023,N_7137,N_8889);
nand U10024 (N_10024,N_8256,N_8135);
nand U10025 (N_10025,N_7261,N_6913);
or U10026 (N_10026,N_6831,N_6525);
nor U10027 (N_10027,N_8071,N_7088);
and U10028 (N_10028,N_8051,N_8320);
nand U10029 (N_10029,N_6342,N_8929);
nor U10030 (N_10030,N_7693,N_6311);
nand U10031 (N_10031,N_7291,N_8615);
or U10032 (N_10032,N_7964,N_6390);
nand U10033 (N_10033,N_7196,N_8366);
and U10034 (N_10034,N_6638,N_6195);
or U10035 (N_10035,N_8148,N_7545);
or U10036 (N_10036,N_7301,N_6384);
nor U10037 (N_10037,N_8968,N_6334);
nand U10038 (N_10038,N_7866,N_8444);
or U10039 (N_10039,N_7530,N_8972);
nand U10040 (N_10040,N_6039,N_7481);
nand U10041 (N_10041,N_6645,N_7413);
nor U10042 (N_10042,N_8097,N_8000);
or U10043 (N_10043,N_7913,N_8766);
or U10044 (N_10044,N_6155,N_6526);
nand U10045 (N_10045,N_7459,N_7758);
nor U10046 (N_10046,N_8518,N_7759);
or U10047 (N_10047,N_8635,N_8638);
nand U10048 (N_10048,N_7251,N_6862);
nand U10049 (N_10049,N_6952,N_6625);
nor U10050 (N_10050,N_6803,N_6721);
nor U10051 (N_10051,N_7702,N_8096);
nor U10052 (N_10052,N_7925,N_6606);
nor U10053 (N_10053,N_7198,N_6001);
nor U10054 (N_10054,N_6352,N_6838);
nand U10055 (N_10055,N_7351,N_7344);
or U10056 (N_10056,N_8238,N_6451);
or U10057 (N_10057,N_6156,N_8372);
and U10058 (N_10058,N_7363,N_6277);
or U10059 (N_10059,N_6586,N_7008);
nor U10060 (N_10060,N_8068,N_6469);
nand U10061 (N_10061,N_6479,N_7003);
nor U10062 (N_10062,N_6036,N_7807);
or U10063 (N_10063,N_7752,N_7373);
and U10064 (N_10064,N_6802,N_8231);
nand U10065 (N_10065,N_7924,N_6505);
and U10066 (N_10066,N_6303,N_6076);
or U10067 (N_10067,N_8940,N_7258);
nor U10068 (N_10068,N_7772,N_8131);
nand U10069 (N_10069,N_8160,N_6741);
nor U10070 (N_10070,N_6286,N_8942);
or U10071 (N_10071,N_8855,N_8911);
nor U10072 (N_10072,N_7199,N_7769);
and U10073 (N_10073,N_6584,N_6376);
nor U10074 (N_10074,N_8735,N_7912);
nor U10075 (N_10075,N_8040,N_8653);
or U10076 (N_10076,N_6552,N_7367);
xor U10077 (N_10077,N_7854,N_7644);
and U10078 (N_10078,N_7142,N_6909);
or U10079 (N_10079,N_6980,N_8106);
nand U10080 (N_10080,N_6664,N_8546);
or U10081 (N_10081,N_7049,N_8646);
nor U10082 (N_10082,N_8116,N_6358);
or U10083 (N_10083,N_6474,N_7770);
nor U10084 (N_10084,N_8470,N_6082);
nor U10085 (N_10085,N_6782,N_6786);
nand U10086 (N_10086,N_7670,N_7939);
nand U10087 (N_10087,N_6044,N_6629);
or U10088 (N_10088,N_8847,N_8198);
or U10089 (N_10089,N_7910,N_8272);
and U10090 (N_10090,N_6607,N_8525);
and U10091 (N_10091,N_6127,N_8563);
or U10092 (N_10092,N_6961,N_8823);
and U10093 (N_10093,N_8675,N_8494);
xor U10094 (N_10094,N_7646,N_6410);
and U10095 (N_10095,N_7213,N_6218);
or U10096 (N_10096,N_6239,N_7302);
nor U10097 (N_10097,N_8279,N_7850);
nor U10098 (N_10098,N_8293,N_8140);
and U10099 (N_10099,N_7080,N_6354);
or U10100 (N_10100,N_6100,N_8989);
nor U10101 (N_10101,N_6057,N_7328);
nand U10102 (N_10102,N_6120,N_8323);
or U10103 (N_10103,N_7439,N_8555);
or U10104 (N_10104,N_7356,N_6242);
nand U10105 (N_10105,N_7820,N_8030);
or U10106 (N_10106,N_7010,N_6446);
nor U10107 (N_10107,N_8110,N_8083);
nor U10108 (N_10108,N_6836,N_8041);
or U10109 (N_10109,N_8467,N_8655);
and U10110 (N_10110,N_8533,N_6643);
nand U10111 (N_10111,N_8560,N_6060);
nand U10112 (N_10112,N_7505,N_8866);
and U10113 (N_10113,N_7030,N_8709);
nand U10114 (N_10114,N_7405,N_8711);
or U10115 (N_10115,N_7640,N_7809);
or U10116 (N_10116,N_8758,N_8878);
nand U10117 (N_10117,N_8295,N_7701);
or U10118 (N_10118,N_6521,N_6844);
nor U10119 (N_10119,N_8021,N_7189);
nor U10120 (N_10120,N_8385,N_6373);
nand U10121 (N_10121,N_6687,N_7051);
or U10122 (N_10122,N_6579,N_7995);
nor U10123 (N_10123,N_6561,N_6062);
nand U10124 (N_10124,N_6891,N_7295);
nor U10125 (N_10125,N_6083,N_8771);
nor U10126 (N_10126,N_7520,N_8493);
nor U10127 (N_10127,N_8165,N_6599);
or U10128 (N_10128,N_7022,N_7290);
nand U10129 (N_10129,N_7272,N_6621);
or U10130 (N_10130,N_8643,N_6888);
and U10131 (N_10131,N_8267,N_7885);
nand U10132 (N_10132,N_7012,N_8350);
nor U10133 (N_10133,N_7695,N_6589);
xnor U10134 (N_10134,N_8144,N_7660);
and U10135 (N_10135,N_8777,N_8007);
nor U10136 (N_10136,N_6788,N_8158);
or U10137 (N_10137,N_8805,N_8609);
nor U10138 (N_10138,N_6331,N_7531);
nand U10139 (N_10139,N_6955,N_8880);
and U10140 (N_10140,N_6391,N_6370);
or U10141 (N_10141,N_6238,N_6714);
nand U10142 (N_10142,N_8499,N_8324);
nor U10143 (N_10143,N_7553,N_6471);
nand U10144 (N_10144,N_8150,N_6053);
and U10145 (N_10145,N_8988,N_8554);
and U10146 (N_10146,N_7529,N_6179);
nand U10147 (N_10147,N_8169,N_6749);
nand U10148 (N_10148,N_8349,N_8230);
nor U10149 (N_10149,N_8539,N_8498);
nor U10150 (N_10150,N_8038,N_6014);
nand U10151 (N_10151,N_7586,N_7683);
nor U10152 (N_10152,N_7480,N_6235);
or U10153 (N_10153,N_7293,N_7089);
or U10154 (N_10154,N_7370,N_7409);
nand U10155 (N_10155,N_7527,N_8270);
or U10156 (N_10156,N_6106,N_7557);
nand U10157 (N_10157,N_7837,N_6736);
or U10158 (N_10158,N_7348,N_7595);
and U10159 (N_10159,N_8857,N_8593);
nand U10160 (N_10160,N_7852,N_8526);
or U10161 (N_10161,N_8138,N_7773);
or U10162 (N_10162,N_6167,N_7984);
and U10163 (N_10163,N_7398,N_7859);
and U10164 (N_10164,N_6612,N_8778);
nand U10165 (N_10165,N_7156,N_6382);
nand U10166 (N_10166,N_7507,N_6500);
and U10167 (N_10167,N_8773,N_8431);
and U10168 (N_10168,N_7175,N_8204);
or U10169 (N_10169,N_8691,N_7116);
nand U10170 (N_10170,N_8425,N_8731);
and U10171 (N_10171,N_8633,N_7068);
nor U10172 (N_10172,N_8216,N_6797);
nand U10173 (N_10173,N_6427,N_6182);
or U10174 (N_10174,N_7903,N_8588);
nor U10175 (N_10175,N_7655,N_8377);
and U10176 (N_10176,N_6316,N_7500);
nor U10177 (N_10177,N_8001,N_8939);
or U10178 (N_10178,N_6835,N_6938);
nand U10179 (N_10179,N_8590,N_8473);
nand U10180 (N_10180,N_7918,N_6992);
nand U10181 (N_10181,N_8089,N_8990);
and U10182 (N_10182,N_6759,N_8606);
nand U10183 (N_10183,N_6956,N_6829);
nor U10184 (N_10184,N_6287,N_8622);
and U10185 (N_10185,N_8074,N_7418);
nand U10186 (N_10186,N_6130,N_7470);
or U10187 (N_10187,N_8276,N_6981);
nand U10188 (N_10188,N_8667,N_8770);
or U10189 (N_10189,N_6580,N_8277);
or U10190 (N_10190,N_7941,N_6147);
or U10191 (N_10191,N_8023,N_6078);
or U10192 (N_10192,N_7643,N_7259);
nor U10193 (N_10193,N_8960,N_7238);
nor U10194 (N_10194,N_7435,N_6701);
nor U10195 (N_10195,N_6887,N_7574);
nand U10196 (N_10196,N_7024,N_6103);
or U10197 (N_10197,N_6260,N_7430);
xnor U10198 (N_10198,N_7166,N_7961);
and U10199 (N_10199,N_6171,N_6659);
and U10200 (N_10200,N_8090,N_6728);
nor U10201 (N_10201,N_7654,N_8626);
nor U10202 (N_10202,N_7581,N_8600);
and U10203 (N_10203,N_7747,N_8858);
nand U10204 (N_10204,N_6886,N_6459);
or U10205 (N_10205,N_7355,N_8504);
nand U10206 (N_10206,N_7598,N_8820);
nor U10207 (N_10207,N_8382,N_6942);
and U10208 (N_10208,N_7879,N_7781);
nand U10209 (N_10209,N_8508,N_7458);
and U10210 (N_10210,N_7110,N_8886);
nor U10211 (N_10211,N_8616,N_6792);
nor U10212 (N_10212,N_7369,N_8334);
or U10213 (N_10213,N_6737,N_8520);
nand U10214 (N_10214,N_8849,N_6319);
nor U10215 (N_10215,N_6550,N_6814);
nor U10216 (N_10216,N_8592,N_6595);
nand U10217 (N_10217,N_6478,N_6293);
or U10218 (N_10218,N_8596,N_6007);
and U10219 (N_10219,N_8983,N_6779);
xor U10220 (N_10220,N_8776,N_8275);
or U10221 (N_10221,N_6610,N_8359);
nor U10222 (N_10222,N_7721,N_6142);
nor U10223 (N_10223,N_7983,N_8800);
and U10224 (N_10224,N_8634,N_6190);
nand U10225 (N_10225,N_6450,N_8387);
nor U10226 (N_10226,N_8818,N_8042);
nand U10227 (N_10227,N_6297,N_7572);
nor U10228 (N_10228,N_7177,N_8695);
nor U10229 (N_10229,N_8984,N_8118);
and U10230 (N_10230,N_7007,N_8798);
and U10231 (N_10231,N_6705,N_8828);
or U10232 (N_10232,N_7563,N_7414);
nand U10233 (N_10233,N_6216,N_7696);
and U10234 (N_10234,N_7917,N_8205);
nor U10235 (N_10235,N_7864,N_6979);
and U10236 (N_10236,N_7585,N_6986);
and U10237 (N_10237,N_8057,N_7390);
nand U10238 (N_10238,N_8581,N_6145);
or U10239 (N_10239,N_6194,N_7113);
or U10240 (N_10240,N_6731,N_8558);
and U10241 (N_10241,N_8712,N_7615);
nor U10242 (N_10242,N_8557,N_6281);
xnor U10243 (N_10243,N_7953,N_6503);
nand U10244 (N_10244,N_7757,N_8240);
or U10245 (N_10245,N_6308,N_7869);
nor U10246 (N_10246,N_8806,N_8793);
nor U10247 (N_10247,N_8727,N_6615);
nor U10248 (N_10248,N_8177,N_7896);
and U10249 (N_10249,N_8915,N_6765);
and U10250 (N_10250,N_8247,N_8055);
nand U10251 (N_10251,N_6553,N_7139);
nor U10252 (N_10252,N_8644,N_7622);
nand U10253 (N_10253,N_7035,N_6488);
and U10254 (N_10254,N_8538,N_6141);
and U10255 (N_10255,N_8812,N_6627);
and U10256 (N_10256,N_6256,N_7764);
or U10257 (N_10257,N_8482,N_8898);
and U10258 (N_10258,N_8311,N_6403);
nand U10259 (N_10259,N_8210,N_6510);
and U10260 (N_10260,N_7393,N_7216);
and U10261 (N_10261,N_7621,N_8783);
or U10262 (N_10262,N_8249,N_7117);
or U10263 (N_10263,N_6031,N_7474);
or U10264 (N_10264,N_8734,N_6989);
nand U10265 (N_10265,N_7966,N_6800);
nand U10266 (N_10266,N_7540,N_7512);
nor U10267 (N_10267,N_7718,N_6452);
nand U10268 (N_10268,N_6622,N_8891);
nand U10269 (N_10269,N_6812,N_7826);
nor U10270 (N_10270,N_7456,N_7593);
and U10271 (N_10271,N_7900,N_6139);
nor U10272 (N_10272,N_8620,N_8784);
or U10273 (N_10273,N_6396,N_8454);
xor U10274 (N_10274,N_8871,N_8917);
and U10275 (N_10275,N_7744,N_8246);
nand U10276 (N_10276,N_7016,N_6270);
nand U10277 (N_10277,N_6196,N_6962);
nand U10278 (N_10278,N_7417,N_8718);
and U10279 (N_10279,N_8760,N_7513);
and U10280 (N_10280,N_7978,N_7551);
or U10281 (N_10281,N_8134,N_8480);
and U10282 (N_10282,N_8611,N_7159);
nand U10283 (N_10283,N_8121,N_6048);
nor U10284 (N_10284,N_8115,N_6037);
or U10285 (N_10285,N_8852,N_7522);
nor U10286 (N_10286,N_7350,N_7106);
nor U10287 (N_10287,N_6320,N_8412);
xor U10288 (N_10288,N_7475,N_7558);
nor U10289 (N_10289,N_7775,N_6804);
nand U10290 (N_10290,N_7408,N_6682);
and U10291 (N_10291,N_8746,N_6003);
nor U10292 (N_10292,N_6827,N_7708);
nor U10293 (N_10293,N_8825,N_8741);
nor U10294 (N_10294,N_8559,N_6473);
or U10295 (N_10295,N_8830,N_8649);
nand U10296 (N_10296,N_6203,N_6648);
and U10297 (N_10297,N_7379,N_7791);
or U10298 (N_10298,N_6937,N_6531);
nand U10299 (N_10299,N_6537,N_6096);
and U10300 (N_10300,N_6366,N_8509);
nand U10301 (N_10301,N_8321,N_8772);
nand U10302 (N_10302,N_6217,N_8391);
and U10303 (N_10303,N_6234,N_7796);
or U10304 (N_10304,N_6483,N_8233);
and U10305 (N_10305,N_7151,N_6029);
and U10306 (N_10306,N_7071,N_8446);
or U10307 (N_10307,N_8072,N_8762);
and U10308 (N_10308,N_7813,N_7963);
nand U10309 (N_10309,N_8998,N_8016);
nand U10310 (N_10310,N_6601,N_8552);
and U10311 (N_10311,N_6360,N_6689);
and U10312 (N_10312,N_6917,N_8319);
and U10313 (N_10313,N_6977,N_8213);
nand U10314 (N_10314,N_6074,N_8841);
and U10315 (N_10315,N_7391,N_6210);
nand U10316 (N_10316,N_6674,N_7260);
nor U10317 (N_10317,N_8137,N_6409);
nor U10318 (N_10318,N_7887,N_6283);
nor U10319 (N_10319,N_6362,N_8703);
nor U10320 (N_10320,N_7017,N_6184);
and U10321 (N_10321,N_8202,N_6712);
nand U10322 (N_10322,N_8073,N_7039);
nor U10323 (N_10323,N_6513,N_7812);
or U10324 (N_10324,N_6968,N_7631);
or U10325 (N_10325,N_7309,N_6998);
nor U10326 (N_10326,N_6634,N_6724);
or U10327 (N_10327,N_8970,N_7006);
nand U10328 (N_10328,N_8656,N_7423);
nand U10329 (N_10329,N_6197,N_7698);
and U10330 (N_10330,N_7739,N_6421);
or U10331 (N_10331,N_6878,N_7015);
and U10332 (N_10332,N_8920,N_8029);
and U10333 (N_10333,N_8994,N_8471);
and U10334 (N_10334,N_7245,N_8477);
nor U10335 (N_10335,N_8241,N_7760);
nor U10336 (N_10336,N_8304,N_6571);
and U10337 (N_10337,N_8550,N_6545);
and U10338 (N_10338,N_8370,N_6146);
nand U10339 (N_10339,N_7648,N_6151);
nand U10340 (N_10340,N_7188,N_7257);
nor U10341 (N_10341,N_7286,N_7101);
or U10342 (N_10342,N_7895,N_8201);
or U10343 (N_10343,N_6655,N_8435);
nor U10344 (N_10344,N_8081,N_7167);
or U10345 (N_10345,N_7292,N_7657);
or U10346 (N_10346,N_7243,N_7028);
and U10347 (N_10347,N_8305,N_6694);
nand U10348 (N_10348,N_8103,N_6207);
or U10349 (N_10349,N_7717,N_6585);
and U10350 (N_10350,N_6444,N_8397);
nor U10351 (N_10351,N_8070,N_7618);
and U10352 (N_10352,N_6849,N_6861);
nor U10353 (N_10353,N_6697,N_6263);
and U10354 (N_10354,N_7170,N_7970);
and U10355 (N_10355,N_7392,N_8881);
or U10356 (N_10356,N_8614,N_7996);
nand U10357 (N_10357,N_7848,N_7331);
and U10358 (N_10358,N_8423,N_6264);
nand U10359 (N_10359,N_7790,N_6202);
and U10360 (N_10360,N_7123,N_7616);
nand U10361 (N_10361,N_8780,N_7524);
nor U10362 (N_10362,N_6717,N_6193);
and U10363 (N_10363,N_6920,N_6751);
or U10364 (N_10364,N_7688,N_6357);
and U10365 (N_10365,N_6188,N_8585);
and U10366 (N_10366,N_6143,N_6119);
and U10367 (N_10367,N_8440,N_8639);
nor U10368 (N_10368,N_6198,N_6019);
xor U10369 (N_10369,N_7814,N_6010);
and U10370 (N_10370,N_8875,N_8921);
nand U10371 (N_10371,N_6040,N_6460);
nor U10372 (N_10372,N_6777,N_7891);
nand U10373 (N_10373,N_6534,N_6204);
nand U10374 (N_10374,N_8476,N_6269);
nand U10375 (N_10375,N_6591,N_8680);
and U10376 (N_10376,N_7821,N_8663);
nand U10377 (N_10377,N_8856,N_6236);
or U10378 (N_10378,N_8595,N_8673);
and U10379 (N_10379,N_7181,N_8342);
nand U10380 (N_10380,N_8422,N_6101);
nor U10381 (N_10381,N_8523,N_8846);
or U10382 (N_10382,N_7779,N_8487);
and U10383 (N_10383,N_6833,N_8203);
nor U10384 (N_10384,N_7495,N_6742);
nor U10385 (N_10385,N_7445,N_8564);
or U10386 (N_10386,N_8936,N_8200);
and U10387 (N_10387,N_6715,N_7205);
nand U10388 (N_10388,N_6159,N_8491);
or U10389 (N_10389,N_6428,N_8674);
and U10390 (N_10390,N_8628,N_7311);
nand U10391 (N_10391,N_7115,N_8327);
nor U10392 (N_10392,N_7014,N_8401);
nand U10393 (N_10393,N_6568,N_6508);
or U10394 (N_10394,N_6191,N_8537);
nor U10395 (N_10395,N_8876,N_6069);
and U10396 (N_10396,N_6957,N_8725);
nor U10397 (N_10397,N_7987,N_7083);
and U10398 (N_10398,N_7605,N_6922);
and U10399 (N_10399,N_8640,N_7107);
or U10400 (N_10400,N_6492,N_7467);
nor U10401 (N_10401,N_8079,N_7462);
nand U10402 (N_10402,N_6517,N_6860);
nor U10403 (N_10403,N_8208,N_8306);
or U10404 (N_10404,N_6657,N_7738);
and U10405 (N_10405,N_6126,N_7884);
xor U10406 (N_10406,N_7601,N_6841);
nor U10407 (N_10407,N_7489,N_6903);
and U10408 (N_10408,N_8748,N_6656);
nor U10409 (N_10409,N_8186,N_8947);
or U10410 (N_10410,N_6305,N_8848);
and U10411 (N_10411,N_7956,N_7727);
nand U10412 (N_10412,N_8280,N_8102);
nor U10413 (N_10413,N_6463,N_8949);
nor U10414 (N_10414,N_8974,N_8164);
nand U10415 (N_10415,N_6275,N_7611);
nand U10416 (N_10416,N_8420,N_7493);
nand U10417 (N_10417,N_7444,N_8146);
and U10418 (N_10418,N_7794,N_6847);
or U10419 (N_10419,N_6455,N_7457);
nor U10420 (N_10420,N_6848,N_8340);
nor U10421 (N_10421,N_8958,N_7905);
nand U10422 (N_10422,N_6032,N_7902);
or U10423 (N_10423,N_8826,N_8922);
nor U10424 (N_10424,N_6950,N_8364);
nand U10425 (N_10425,N_8084,N_8645);
nand U10426 (N_10426,N_6520,N_8248);
or U10427 (N_10427,N_8987,N_8629);
or U10428 (N_10428,N_6720,N_7501);
nand U10429 (N_10429,N_7208,N_6730);
and U10430 (N_10430,N_7352,N_6811);
nand U10431 (N_10431,N_6605,N_7125);
or U10432 (N_10432,N_6940,N_6464);
nand U10433 (N_10433,N_7009,N_7056);
and U10434 (N_10434,N_6121,N_7802);
or U10435 (N_10435,N_6272,N_6807);
nor U10436 (N_10436,N_6703,N_6140);
and U10437 (N_10437,N_8945,N_6970);
nand U10438 (N_10438,N_7519,N_8251);
nor U10439 (N_10439,N_8624,N_7032);
or U10440 (N_10440,N_6547,N_7023);
and U10441 (N_10441,N_6947,N_7034);
xnor U10442 (N_10442,N_8701,N_8303);
nor U10443 (N_10443,N_7157,N_7967);
nor U10444 (N_10444,N_7096,N_6509);
and U10445 (N_10445,N_8632,N_8228);
or U10446 (N_10446,N_8496,N_7250);
and U10447 (N_10447,N_8450,N_8817);
nand U10448 (N_10448,N_7914,N_8676);
or U10449 (N_10449,N_8664,N_8288);
nor U10450 (N_10450,N_8531,N_8265);
nand U10451 (N_10451,N_6843,N_7412);
and U10452 (N_10452,N_6975,N_7591);
nor U10453 (N_10453,N_8699,N_8107);
nor U10454 (N_10454,N_7013,N_7988);
and U10455 (N_10455,N_6288,N_8747);
or U10456 (N_10456,N_7832,N_6222);
nor U10457 (N_10457,N_6883,N_7365);
and U10458 (N_10458,N_7225,N_7637);
and U10459 (N_10459,N_6996,N_7300);
nand U10460 (N_10460,N_8351,N_8433);
or U10461 (N_10461,N_8308,N_6969);
xnor U10462 (N_10462,N_6773,N_8500);
nor U10463 (N_10463,N_8417,N_7454);
nor U10464 (N_10464,N_7511,N_8877);
nor U10465 (N_10465,N_6733,N_6592);
or U10466 (N_10466,N_8299,N_8854);
nor U10467 (N_10467,N_8924,N_6948);
nor U10468 (N_10468,N_8456,N_7656);
nand U10469 (N_10469,N_7678,N_6538);
nor U10470 (N_10470,N_6165,N_8853);
nand U10471 (N_10471,N_8159,N_8517);
and U10472 (N_10472,N_6314,N_8937);
and U10473 (N_10473,N_8966,N_8507);
or U10474 (N_10474,N_8774,N_8114);
nand U10475 (N_10475,N_7183,N_7800);
or U10476 (N_10476,N_7710,N_6246);
or U10477 (N_10477,N_7990,N_6498);
xnor U10478 (N_10478,N_7210,N_6189);
nor U10479 (N_10479,N_8549,N_7789);
and U10480 (N_10480,N_7381,N_6864);
and U10481 (N_10481,N_7803,N_8790);
nor U10482 (N_10482,N_7248,N_7109);
or U10483 (N_10483,N_6918,N_6176);
and U10484 (N_10484,N_7451,N_7223);
xnor U10485 (N_10485,N_6385,N_7652);
nand U10486 (N_10486,N_7625,N_6340);
nor U10487 (N_10487,N_8515,N_8468);
nand U10488 (N_10488,N_7036,N_6268);
or U10489 (N_10489,N_7750,N_7829);
nor U10490 (N_10490,N_7473,N_6963);
and U10491 (N_10491,N_7499,N_8542);
nor U10492 (N_10492,N_7337,N_7236);
and U10493 (N_10493,N_6535,N_7384);
nor U10494 (N_10494,N_6670,N_8567);
nand U10495 (N_10495,N_6863,N_7179);
xor U10496 (N_10496,N_7296,N_6241);
nor U10497 (N_10497,N_6925,N_8003);
xor U10498 (N_10498,N_8912,N_8333);
or U10499 (N_10499,N_7613,N_7951);
nand U10500 (N_10500,N_8646,N_7125);
and U10501 (N_10501,N_7602,N_7037);
nand U10502 (N_10502,N_6487,N_8802);
and U10503 (N_10503,N_7883,N_8196);
nand U10504 (N_10504,N_6752,N_7683);
nand U10505 (N_10505,N_6054,N_7829);
nor U10506 (N_10506,N_7655,N_7652);
or U10507 (N_10507,N_7582,N_8340);
nor U10508 (N_10508,N_7561,N_8614);
nor U10509 (N_10509,N_6843,N_6436);
or U10510 (N_10510,N_6422,N_6688);
and U10511 (N_10511,N_6351,N_7292);
nor U10512 (N_10512,N_7744,N_7845);
nand U10513 (N_10513,N_7412,N_6369);
and U10514 (N_10514,N_6255,N_7728);
nand U10515 (N_10515,N_7036,N_6004);
nand U10516 (N_10516,N_8394,N_8139);
nand U10517 (N_10517,N_7157,N_6805);
nor U10518 (N_10518,N_8370,N_7401);
nand U10519 (N_10519,N_8919,N_6522);
and U10520 (N_10520,N_6328,N_8386);
xnor U10521 (N_10521,N_7516,N_8203);
xor U10522 (N_10522,N_8043,N_8324);
nand U10523 (N_10523,N_6555,N_6649);
and U10524 (N_10524,N_6675,N_6250);
or U10525 (N_10525,N_8896,N_8324);
and U10526 (N_10526,N_6177,N_6672);
nor U10527 (N_10527,N_6002,N_6917);
nand U10528 (N_10528,N_7039,N_8722);
and U10529 (N_10529,N_6294,N_7408);
nand U10530 (N_10530,N_8717,N_6433);
or U10531 (N_10531,N_6260,N_6096);
and U10532 (N_10532,N_6472,N_7207);
nand U10533 (N_10533,N_6849,N_7111);
nor U10534 (N_10534,N_7182,N_7576);
and U10535 (N_10535,N_7232,N_8447);
and U10536 (N_10536,N_8120,N_7143);
nor U10537 (N_10537,N_8493,N_6436);
nor U10538 (N_10538,N_8107,N_6304);
and U10539 (N_10539,N_7527,N_6578);
nor U10540 (N_10540,N_7060,N_8391);
and U10541 (N_10541,N_7751,N_6817);
and U10542 (N_10542,N_6180,N_8597);
nand U10543 (N_10543,N_6718,N_7819);
xor U10544 (N_10544,N_6249,N_7428);
nor U10545 (N_10545,N_7064,N_6752);
nor U10546 (N_10546,N_7670,N_8243);
or U10547 (N_10547,N_7315,N_8534);
and U10548 (N_10548,N_6656,N_8623);
nor U10549 (N_10549,N_6827,N_6765);
nor U10550 (N_10550,N_6375,N_8722);
or U10551 (N_10551,N_8487,N_8962);
nor U10552 (N_10552,N_8687,N_8438);
and U10553 (N_10553,N_8052,N_7467);
nand U10554 (N_10554,N_6536,N_8507);
and U10555 (N_10555,N_7329,N_6451);
or U10556 (N_10556,N_6955,N_8049);
or U10557 (N_10557,N_6728,N_8787);
or U10558 (N_10558,N_7067,N_8849);
or U10559 (N_10559,N_8660,N_8395);
xor U10560 (N_10560,N_8331,N_6301);
and U10561 (N_10561,N_8755,N_7070);
or U10562 (N_10562,N_8830,N_8934);
nor U10563 (N_10563,N_6639,N_8943);
nand U10564 (N_10564,N_6864,N_8339);
nor U10565 (N_10565,N_6124,N_8923);
nor U10566 (N_10566,N_8875,N_8216);
or U10567 (N_10567,N_8553,N_7917);
nand U10568 (N_10568,N_8155,N_8673);
nand U10569 (N_10569,N_7979,N_8079);
and U10570 (N_10570,N_8434,N_8736);
and U10571 (N_10571,N_6554,N_7326);
nand U10572 (N_10572,N_7523,N_7556);
and U10573 (N_10573,N_6449,N_8162);
nand U10574 (N_10574,N_8486,N_6580);
and U10575 (N_10575,N_6655,N_7386);
and U10576 (N_10576,N_7816,N_7451);
nor U10577 (N_10577,N_8412,N_6022);
nand U10578 (N_10578,N_6035,N_8553);
and U10579 (N_10579,N_6646,N_8072);
and U10580 (N_10580,N_8161,N_8583);
or U10581 (N_10581,N_6868,N_8245);
nor U10582 (N_10582,N_6339,N_6836);
nor U10583 (N_10583,N_6817,N_6604);
nand U10584 (N_10584,N_8188,N_6290);
and U10585 (N_10585,N_8823,N_8483);
or U10586 (N_10586,N_8239,N_8894);
and U10587 (N_10587,N_7884,N_7544);
and U10588 (N_10588,N_8869,N_7451);
or U10589 (N_10589,N_6005,N_8424);
and U10590 (N_10590,N_6275,N_7307);
and U10591 (N_10591,N_7217,N_8141);
and U10592 (N_10592,N_8611,N_6781);
and U10593 (N_10593,N_7933,N_8247);
and U10594 (N_10594,N_7028,N_6114);
nor U10595 (N_10595,N_6409,N_7645);
xnor U10596 (N_10596,N_6963,N_6789);
and U10597 (N_10597,N_6115,N_6828);
nand U10598 (N_10598,N_7521,N_8223);
and U10599 (N_10599,N_8780,N_6140);
or U10600 (N_10600,N_6412,N_8720);
or U10601 (N_10601,N_8813,N_8951);
nand U10602 (N_10602,N_7598,N_6996);
or U10603 (N_10603,N_6295,N_7171);
or U10604 (N_10604,N_6542,N_8512);
nor U10605 (N_10605,N_6784,N_7325);
nor U10606 (N_10606,N_7723,N_8380);
nand U10607 (N_10607,N_6925,N_7585);
and U10608 (N_10608,N_6913,N_7055);
and U10609 (N_10609,N_7637,N_6094);
or U10610 (N_10610,N_7601,N_6390);
or U10611 (N_10611,N_7324,N_7723);
or U10612 (N_10612,N_7385,N_8474);
and U10613 (N_10613,N_6660,N_6424);
or U10614 (N_10614,N_7681,N_7443);
or U10615 (N_10615,N_8976,N_6144);
nand U10616 (N_10616,N_8637,N_8951);
and U10617 (N_10617,N_6023,N_7183);
nor U10618 (N_10618,N_6301,N_8721);
nor U10619 (N_10619,N_7975,N_6177);
or U10620 (N_10620,N_6424,N_7401);
or U10621 (N_10621,N_8276,N_8251);
or U10622 (N_10622,N_6332,N_7744);
nand U10623 (N_10623,N_6617,N_6397);
nor U10624 (N_10624,N_7533,N_6944);
nand U10625 (N_10625,N_8261,N_6077);
and U10626 (N_10626,N_7360,N_7071);
or U10627 (N_10627,N_6871,N_7259);
or U10628 (N_10628,N_6968,N_7305);
nor U10629 (N_10629,N_7536,N_7016);
or U10630 (N_10630,N_6160,N_6015);
and U10631 (N_10631,N_8026,N_6882);
nand U10632 (N_10632,N_8215,N_7035);
or U10633 (N_10633,N_8383,N_8830);
nand U10634 (N_10634,N_6871,N_6593);
xnor U10635 (N_10635,N_8402,N_8722);
or U10636 (N_10636,N_7574,N_8234);
nand U10637 (N_10637,N_7668,N_8477);
and U10638 (N_10638,N_7391,N_7415);
and U10639 (N_10639,N_7349,N_6593);
and U10640 (N_10640,N_7315,N_8152);
xor U10641 (N_10641,N_6569,N_8547);
nor U10642 (N_10642,N_6327,N_8293);
and U10643 (N_10643,N_7895,N_8578);
nor U10644 (N_10644,N_6676,N_8074);
nand U10645 (N_10645,N_8707,N_7176);
nor U10646 (N_10646,N_8397,N_6716);
nand U10647 (N_10647,N_6302,N_8181);
nor U10648 (N_10648,N_7849,N_6534);
or U10649 (N_10649,N_8806,N_6201);
nand U10650 (N_10650,N_7813,N_6578);
and U10651 (N_10651,N_6738,N_6520);
or U10652 (N_10652,N_7707,N_7466);
nand U10653 (N_10653,N_8393,N_7813);
nor U10654 (N_10654,N_8253,N_6541);
nand U10655 (N_10655,N_7664,N_7386);
and U10656 (N_10656,N_8670,N_6847);
nor U10657 (N_10657,N_6830,N_7653);
xnor U10658 (N_10658,N_7010,N_6352);
or U10659 (N_10659,N_6597,N_7719);
or U10660 (N_10660,N_8008,N_6783);
or U10661 (N_10661,N_7520,N_6987);
nor U10662 (N_10662,N_7800,N_7719);
and U10663 (N_10663,N_6630,N_8023);
and U10664 (N_10664,N_8802,N_6470);
nor U10665 (N_10665,N_7398,N_6432);
nand U10666 (N_10666,N_7251,N_7885);
nand U10667 (N_10667,N_8104,N_7480);
xor U10668 (N_10668,N_8181,N_6541);
or U10669 (N_10669,N_6688,N_6823);
nand U10670 (N_10670,N_6213,N_6167);
nand U10671 (N_10671,N_6301,N_8690);
xnor U10672 (N_10672,N_8520,N_7913);
and U10673 (N_10673,N_7537,N_7389);
nor U10674 (N_10674,N_7522,N_6265);
and U10675 (N_10675,N_8928,N_6369);
nand U10676 (N_10676,N_6677,N_7280);
xor U10677 (N_10677,N_6655,N_6703);
nand U10678 (N_10678,N_8041,N_6206);
nand U10679 (N_10679,N_6819,N_8548);
or U10680 (N_10680,N_7357,N_7916);
nand U10681 (N_10681,N_7502,N_8407);
or U10682 (N_10682,N_6872,N_6206);
and U10683 (N_10683,N_7345,N_7657);
and U10684 (N_10684,N_7474,N_7280);
or U10685 (N_10685,N_7999,N_8066);
nor U10686 (N_10686,N_6970,N_6342);
xor U10687 (N_10687,N_8360,N_7875);
nand U10688 (N_10688,N_6018,N_7791);
or U10689 (N_10689,N_6450,N_7684);
nand U10690 (N_10690,N_8189,N_7779);
nand U10691 (N_10691,N_8083,N_7124);
or U10692 (N_10692,N_8238,N_7213);
nand U10693 (N_10693,N_7638,N_7881);
nand U10694 (N_10694,N_7726,N_6590);
or U10695 (N_10695,N_6269,N_6162);
or U10696 (N_10696,N_8930,N_6182);
and U10697 (N_10697,N_6159,N_8372);
and U10698 (N_10698,N_6190,N_8221);
and U10699 (N_10699,N_6659,N_8138);
nand U10700 (N_10700,N_8102,N_8277);
and U10701 (N_10701,N_8096,N_6297);
and U10702 (N_10702,N_6560,N_7648);
and U10703 (N_10703,N_8377,N_8212);
nor U10704 (N_10704,N_7066,N_8442);
or U10705 (N_10705,N_7479,N_6552);
nor U10706 (N_10706,N_7816,N_8806);
nor U10707 (N_10707,N_7864,N_6259);
nand U10708 (N_10708,N_6788,N_7476);
or U10709 (N_10709,N_6533,N_8420);
and U10710 (N_10710,N_7814,N_8558);
or U10711 (N_10711,N_6890,N_8897);
or U10712 (N_10712,N_8899,N_8015);
nand U10713 (N_10713,N_7109,N_7409);
and U10714 (N_10714,N_7129,N_6406);
and U10715 (N_10715,N_6404,N_6703);
nand U10716 (N_10716,N_7360,N_6451);
or U10717 (N_10717,N_8381,N_6263);
and U10718 (N_10718,N_6648,N_6129);
nand U10719 (N_10719,N_6289,N_6918);
xnor U10720 (N_10720,N_6065,N_7548);
nor U10721 (N_10721,N_7986,N_6782);
nand U10722 (N_10722,N_7993,N_6502);
xor U10723 (N_10723,N_7789,N_6024);
nor U10724 (N_10724,N_7470,N_7178);
nand U10725 (N_10725,N_8296,N_7202);
and U10726 (N_10726,N_8991,N_6119);
nand U10727 (N_10727,N_7319,N_7053);
and U10728 (N_10728,N_6951,N_7785);
nor U10729 (N_10729,N_6531,N_7507);
or U10730 (N_10730,N_6951,N_7906);
nor U10731 (N_10731,N_7293,N_6616);
nand U10732 (N_10732,N_8275,N_7254);
and U10733 (N_10733,N_6439,N_8659);
nor U10734 (N_10734,N_6846,N_8438);
or U10735 (N_10735,N_6721,N_8995);
nand U10736 (N_10736,N_6903,N_6481);
or U10737 (N_10737,N_6636,N_6661);
nand U10738 (N_10738,N_6766,N_6084);
xor U10739 (N_10739,N_7841,N_7807);
nand U10740 (N_10740,N_7275,N_6377);
or U10741 (N_10741,N_8917,N_6052);
or U10742 (N_10742,N_8356,N_7095);
and U10743 (N_10743,N_7268,N_7696);
nand U10744 (N_10744,N_6885,N_6991);
and U10745 (N_10745,N_6576,N_8656);
and U10746 (N_10746,N_6280,N_7550);
nor U10747 (N_10747,N_6418,N_6575);
nor U10748 (N_10748,N_6572,N_6475);
nor U10749 (N_10749,N_6464,N_8948);
nor U10750 (N_10750,N_8465,N_8179);
or U10751 (N_10751,N_6459,N_6028);
nor U10752 (N_10752,N_6974,N_6287);
nor U10753 (N_10753,N_6877,N_8122);
nor U10754 (N_10754,N_6884,N_7759);
nor U10755 (N_10755,N_6929,N_6224);
or U10756 (N_10756,N_8674,N_8109);
or U10757 (N_10757,N_6446,N_7464);
nand U10758 (N_10758,N_8317,N_7354);
nand U10759 (N_10759,N_6422,N_6784);
or U10760 (N_10760,N_6337,N_8594);
nor U10761 (N_10761,N_7729,N_7157);
nor U10762 (N_10762,N_7854,N_7498);
nor U10763 (N_10763,N_7707,N_8713);
nand U10764 (N_10764,N_6979,N_7909);
nand U10765 (N_10765,N_6089,N_7999);
nand U10766 (N_10766,N_8293,N_8562);
or U10767 (N_10767,N_7649,N_7183);
and U10768 (N_10768,N_7720,N_7987);
and U10769 (N_10769,N_7749,N_6137);
nand U10770 (N_10770,N_8936,N_6716);
xor U10771 (N_10771,N_7131,N_8739);
or U10772 (N_10772,N_7326,N_6758);
nor U10773 (N_10773,N_7589,N_8904);
and U10774 (N_10774,N_8315,N_6794);
xnor U10775 (N_10775,N_7169,N_7601);
nor U10776 (N_10776,N_6342,N_7282);
or U10777 (N_10777,N_6480,N_7971);
or U10778 (N_10778,N_8320,N_8327);
nor U10779 (N_10779,N_8977,N_8622);
and U10780 (N_10780,N_8886,N_7165);
nor U10781 (N_10781,N_8773,N_6428);
nand U10782 (N_10782,N_8463,N_6291);
or U10783 (N_10783,N_6980,N_7276);
and U10784 (N_10784,N_8562,N_6014);
or U10785 (N_10785,N_6227,N_6360);
and U10786 (N_10786,N_8283,N_6318);
nor U10787 (N_10787,N_7831,N_8131);
nand U10788 (N_10788,N_6235,N_7855);
nand U10789 (N_10789,N_7069,N_7876);
and U10790 (N_10790,N_7675,N_6842);
or U10791 (N_10791,N_7808,N_8838);
or U10792 (N_10792,N_7621,N_7356);
nand U10793 (N_10793,N_6549,N_6431);
or U10794 (N_10794,N_6232,N_7386);
and U10795 (N_10795,N_7514,N_6933);
nand U10796 (N_10796,N_7319,N_6121);
and U10797 (N_10797,N_8371,N_7298);
nand U10798 (N_10798,N_6103,N_7566);
or U10799 (N_10799,N_8047,N_7549);
nor U10800 (N_10800,N_6997,N_7216);
and U10801 (N_10801,N_8437,N_8617);
nand U10802 (N_10802,N_7735,N_7730);
nor U10803 (N_10803,N_6062,N_6119);
or U10804 (N_10804,N_8004,N_6321);
or U10805 (N_10805,N_7702,N_7353);
nor U10806 (N_10806,N_8396,N_6006);
and U10807 (N_10807,N_7754,N_6161);
and U10808 (N_10808,N_7380,N_6556);
nor U10809 (N_10809,N_7552,N_7211);
or U10810 (N_10810,N_8268,N_7274);
and U10811 (N_10811,N_6758,N_7553);
and U10812 (N_10812,N_6786,N_7182);
xnor U10813 (N_10813,N_7262,N_6432);
nand U10814 (N_10814,N_6051,N_8395);
nor U10815 (N_10815,N_8108,N_8158);
and U10816 (N_10816,N_7984,N_6445);
and U10817 (N_10817,N_8152,N_7873);
nor U10818 (N_10818,N_6900,N_7140);
nand U10819 (N_10819,N_7879,N_7402);
and U10820 (N_10820,N_8211,N_8816);
nand U10821 (N_10821,N_7186,N_7484);
or U10822 (N_10822,N_8234,N_8928);
or U10823 (N_10823,N_7479,N_7227);
nor U10824 (N_10824,N_7800,N_8141);
or U10825 (N_10825,N_7168,N_6963);
xor U10826 (N_10826,N_8647,N_8662);
or U10827 (N_10827,N_8333,N_6822);
and U10828 (N_10828,N_6382,N_7374);
or U10829 (N_10829,N_8393,N_7782);
nor U10830 (N_10830,N_8039,N_7404);
and U10831 (N_10831,N_6979,N_7907);
xnor U10832 (N_10832,N_6308,N_6607);
or U10833 (N_10833,N_7059,N_7026);
and U10834 (N_10834,N_8739,N_6744);
nor U10835 (N_10835,N_6009,N_8646);
or U10836 (N_10836,N_6890,N_8609);
nand U10837 (N_10837,N_6614,N_8807);
or U10838 (N_10838,N_6820,N_7557);
nand U10839 (N_10839,N_8820,N_7550);
nor U10840 (N_10840,N_6764,N_6183);
nor U10841 (N_10841,N_8678,N_8566);
and U10842 (N_10842,N_7433,N_8177);
and U10843 (N_10843,N_6566,N_6616);
and U10844 (N_10844,N_6220,N_8429);
nor U10845 (N_10845,N_7949,N_7951);
nand U10846 (N_10846,N_6463,N_8654);
and U10847 (N_10847,N_8360,N_7614);
and U10848 (N_10848,N_6798,N_7256);
nand U10849 (N_10849,N_8424,N_8872);
or U10850 (N_10850,N_7941,N_7348);
nor U10851 (N_10851,N_8624,N_8918);
and U10852 (N_10852,N_7015,N_8875);
nand U10853 (N_10853,N_7755,N_6124);
nor U10854 (N_10854,N_6046,N_7237);
nor U10855 (N_10855,N_6821,N_8134);
or U10856 (N_10856,N_7485,N_6779);
or U10857 (N_10857,N_7340,N_8287);
and U10858 (N_10858,N_6314,N_7534);
or U10859 (N_10859,N_6623,N_8873);
or U10860 (N_10860,N_8915,N_6007);
and U10861 (N_10861,N_8179,N_6219);
nor U10862 (N_10862,N_6001,N_8124);
and U10863 (N_10863,N_7579,N_6295);
nand U10864 (N_10864,N_7402,N_6368);
nor U10865 (N_10865,N_7886,N_6799);
or U10866 (N_10866,N_8978,N_7914);
or U10867 (N_10867,N_6322,N_7277);
or U10868 (N_10868,N_7276,N_8889);
nand U10869 (N_10869,N_7542,N_8909);
and U10870 (N_10870,N_6232,N_8765);
nor U10871 (N_10871,N_6187,N_6442);
nand U10872 (N_10872,N_8652,N_8913);
nand U10873 (N_10873,N_6948,N_6904);
or U10874 (N_10874,N_6563,N_6159);
and U10875 (N_10875,N_6037,N_8434);
nor U10876 (N_10876,N_6089,N_6977);
nand U10877 (N_10877,N_7941,N_6952);
nand U10878 (N_10878,N_6636,N_6431);
nand U10879 (N_10879,N_6393,N_8985);
nor U10880 (N_10880,N_8873,N_7427);
or U10881 (N_10881,N_7383,N_8781);
or U10882 (N_10882,N_7264,N_8087);
xnor U10883 (N_10883,N_6336,N_8347);
and U10884 (N_10884,N_6103,N_8578);
and U10885 (N_10885,N_6744,N_6319);
nor U10886 (N_10886,N_7188,N_6313);
or U10887 (N_10887,N_7486,N_8468);
and U10888 (N_10888,N_8663,N_6281);
or U10889 (N_10889,N_8252,N_7848);
or U10890 (N_10890,N_7859,N_7625);
and U10891 (N_10891,N_6369,N_8744);
or U10892 (N_10892,N_8834,N_8855);
and U10893 (N_10893,N_7262,N_8485);
nand U10894 (N_10894,N_6680,N_7554);
or U10895 (N_10895,N_7803,N_8792);
and U10896 (N_10896,N_6976,N_6696);
or U10897 (N_10897,N_8809,N_8952);
and U10898 (N_10898,N_7870,N_8875);
nand U10899 (N_10899,N_6427,N_7663);
or U10900 (N_10900,N_6150,N_8529);
and U10901 (N_10901,N_7322,N_7121);
nand U10902 (N_10902,N_6716,N_7792);
nand U10903 (N_10903,N_7766,N_8937);
nand U10904 (N_10904,N_8651,N_8099);
nor U10905 (N_10905,N_6828,N_6784);
nand U10906 (N_10906,N_6119,N_8527);
and U10907 (N_10907,N_6799,N_7336);
nor U10908 (N_10908,N_8296,N_8913);
nand U10909 (N_10909,N_6174,N_6318);
nor U10910 (N_10910,N_6628,N_6560);
and U10911 (N_10911,N_8439,N_8158);
or U10912 (N_10912,N_7019,N_8112);
or U10913 (N_10913,N_8259,N_6391);
nor U10914 (N_10914,N_6434,N_8845);
nand U10915 (N_10915,N_8175,N_6440);
or U10916 (N_10916,N_8101,N_8050);
nand U10917 (N_10917,N_8163,N_7145);
and U10918 (N_10918,N_6483,N_8971);
nor U10919 (N_10919,N_7634,N_8926);
nand U10920 (N_10920,N_7540,N_6672);
nand U10921 (N_10921,N_8290,N_8922);
nand U10922 (N_10922,N_6373,N_6430);
xor U10923 (N_10923,N_7070,N_8588);
and U10924 (N_10924,N_8021,N_7133);
or U10925 (N_10925,N_6582,N_8095);
and U10926 (N_10926,N_6981,N_6446);
and U10927 (N_10927,N_7583,N_7803);
xnor U10928 (N_10928,N_8185,N_8828);
and U10929 (N_10929,N_6457,N_6425);
and U10930 (N_10930,N_7147,N_6376);
nor U10931 (N_10931,N_6346,N_6207);
nand U10932 (N_10932,N_8273,N_6027);
or U10933 (N_10933,N_8882,N_7415);
nand U10934 (N_10934,N_6910,N_8377);
nor U10935 (N_10935,N_6006,N_8862);
nand U10936 (N_10936,N_8494,N_6086);
and U10937 (N_10937,N_6877,N_6591);
or U10938 (N_10938,N_6468,N_6488);
nor U10939 (N_10939,N_7475,N_8472);
or U10940 (N_10940,N_8371,N_8247);
nor U10941 (N_10941,N_8760,N_7224);
or U10942 (N_10942,N_6337,N_7333);
nor U10943 (N_10943,N_8421,N_7864);
nand U10944 (N_10944,N_8174,N_8353);
and U10945 (N_10945,N_7256,N_6782);
and U10946 (N_10946,N_8728,N_7975);
or U10947 (N_10947,N_8842,N_8319);
or U10948 (N_10948,N_6475,N_7387);
or U10949 (N_10949,N_8527,N_8687);
nor U10950 (N_10950,N_6771,N_8266);
nor U10951 (N_10951,N_7858,N_7399);
and U10952 (N_10952,N_8174,N_6507);
nor U10953 (N_10953,N_7573,N_7393);
or U10954 (N_10954,N_8719,N_7846);
or U10955 (N_10955,N_7003,N_8288);
nor U10956 (N_10956,N_7247,N_6220);
nand U10957 (N_10957,N_7640,N_6073);
nor U10958 (N_10958,N_8531,N_8970);
nand U10959 (N_10959,N_8679,N_7233);
and U10960 (N_10960,N_7803,N_8986);
or U10961 (N_10961,N_7382,N_7970);
nand U10962 (N_10962,N_6639,N_6282);
and U10963 (N_10963,N_6279,N_6889);
nand U10964 (N_10964,N_8115,N_7484);
nand U10965 (N_10965,N_8779,N_7501);
nand U10966 (N_10966,N_6248,N_6874);
or U10967 (N_10967,N_6933,N_6595);
and U10968 (N_10968,N_7489,N_8880);
nor U10969 (N_10969,N_8024,N_8896);
or U10970 (N_10970,N_7129,N_7530);
nor U10971 (N_10971,N_7473,N_8484);
nand U10972 (N_10972,N_6493,N_8718);
and U10973 (N_10973,N_7900,N_8575);
or U10974 (N_10974,N_7479,N_8934);
nor U10975 (N_10975,N_6641,N_7995);
nand U10976 (N_10976,N_7557,N_8146);
nand U10977 (N_10977,N_8664,N_8132);
or U10978 (N_10978,N_6546,N_7377);
nor U10979 (N_10979,N_8618,N_6342);
nand U10980 (N_10980,N_7962,N_7226);
xor U10981 (N_10981,N_8208,N_8126);
nand U10982 (N_10982,N_6835,N_7354);
nor U10983 (N_10983,N_7201,N_8040);
nor U10984 (N_10984,N_7754,N_7625);
nand U10985 (N_10985,N_7315,N_6867);
nand U10986 (N_10986,N_8231,N_8781);
and U10987 (N_10987,N_8475,N_6702);
or U10988 (N_10988,N_6232,N_8820);
nand U10989 (N_10989,N_7927,N_8485);
nand U10990 (N_10990,N_8543,N_7659);
or U10991 (N_10991,N_6192,N_6603);
nor U10992 (N_10992,N_8926,N_8863);
nor U10993 (N_10993,N_8979,N_8525);
nor U10994 (N_10994,N_7553,N_6820);
nand U10995 (N_10995,N_8791,N_8367);
and U10996 (N_10996,N_7102,N_8398);
nand U10997 (N_10997,N_8448,N_7523);
and U10998 (N_10998,N_6658,N_8771);
or U10999 (N_10999,N_6305,N_8504);
and U11000 (N_11000,N_6848,N_8025);
nand U11001 (N_11001,N_7341,N_6724);
or U11002 (N_11002,N_8681,N_8118);
nand U11003 (N_11003,N_8225,N_6384);
or U11004 (N_11004,N_6199,N_8576);
or U11005 (N_11005,N_6840,N_7283);
and U11006 (N_11006,N_8845,N_6748);
and U11007 (N_11007,N_8675,N_6771);
or U11008 (N_11008,N_6603,N_6938);
or U11009 (N_11009,N_8666,N_7253);
nor U11010 (N_11010,N_6032,N_7150);
and U11011 (N_11011,N_6924,N_7202);
and U11012 (N_11012,N_7870,N_6651);
and U11013 (N_11013,N_6243,N_8084);
and U11014 (N_11014,N_7705,N_8642);
and U11015 (N_11015,N_7542,N_7497);
nor U11016 (N_11016,N_8886,N_7589);
and U11017 (N_11017,N_8748,N_8972);
and U11018 (N_11018,N_8156,N_6608);
nand U11019 (N_11019,N_6880,N_6370);
nand U11020 (N_11020,N_7867,N_8308);
nor U11021 (N_11021,N_8560,N_6139);
nand U11022 (N_11022,N_7033,N_7593);
and U11023 (N_11023,N_6650,N_6312);
nand U11024 (N_11024,N_7066,N_8622);
or U11025 (N_11025,N_7826,N_6668);
nand U11026 (N_11026,N_8320,N_8247);
nor U11027 (N_11027,N_8207,N_7566);
and U11028 (N_11028,N_7022,N_7212);
nor U11029 (N_11029,N_7382,N_8259);
nand U11030 (N_11030,N_8998,N_6905);
nor U11031 (N_11031,N_6478,N_7420);
or U11032 (N_11032,N_7638,N_6008);
nand U11033 (N_11033,N_8817,N_7202);
and U11034 (N_11034,N_7569,N_7597);
nor U11035 (N_11035,N_7616,N_7318);
nor U11036 (N_11036,N_8241,N_6743);
or U11037 (N_11037,N_8006,N_7431);
or U11038 (N_11038,N_7224,N_6107);
nand U11039 (N_11039,N_7733,N_8209);
nand U11040 (N_11040,N_8362,N_6992);
and U11041 (N_11041,N_8319,N_8331);
nand U11042 (N_11042,N_6027,N_6608);
or U11043 (N_11043,N_8079,N_6641);
nand U11044 (N_11044,N_7546,N_8812);
nor U11045 (N_11045,N_8045,N_7521);
and U11046 (N_11046,N_8982,N_6612);
nand U11047 (N_11047,N_6001,N_8353);
nand U11048 (N_11048,N_6890,N_8754);
or U11049 (N_11049,N_6827,N_8734);
nand U11050 (N_11050,N_8655,N_7134);
and U11051 (N_11051,N_8040,N_8494);
and U11052 (N_11052,N_6616,N_7464);
nor U11053 (N_11053,N_6852,N_8446);
and U11054 (N_11054,N_7903,N_6389);
or U11055 (N_11055,N_6197,N_8667);
nand U11056 (N_11056,N_6007,N_7604);
nand U11057 (N_11057,N_8588,N_8412);
nor U11058 (N_11058,N_6141,N_7527);
nand U11059 (N_11059,N_7399,N_8758);
nand U11060 (N_11060,N_8623,N_7381);
and U11061 (N_11061,N_6557,N_7294);
and U11062 (N_11062,N_8230,N_7275);
nor U11063 (N_11063,N_7996,N_8492);
and U11064 (N_11064,N_7196,N_8430);
nor U11065 (N_11065,N_6793,N_6277);
xor U11066 (N_11066,N_7174,N_7632);
and U11067 (N_11067,N_7278,N_6307);
nor U11068 (N_11068,N_8021,N_6405);
or U11069 (N_11069,N_8896,N_8657);
nor U11070 (N_11070,N_6838,N_6457);
or U11071 (N_11071,N_7110,N_7199);
nand U11072 (N_11072,N_8175,N_7865);
nor U11073 (N_11073,N_7183,N_7912);
nand U11074 (N_11074,N_7502,N_6526);
or U11075 (N_11075,N_7191,N_7484);
nor U11076 (N_11076,N_6495,N_6209);
or U11077 (N_11077,N_8721,N_8570);
nand U11078 (N_11078,N_8859,N_7824);
or U11079 (N_11079,N_7680,N_7059);
or U11080 (N_11080,N_6139,N_7873);
nand U11081 (N_11081,N_8047,N_7356);
or U11082 (N_11082,N_6688,N_6997);
nor U11083 (N_11083,N_7559,N_6195);
nor U11084 (N_11084,N_8021,N_7642);
and U11085 (N_11085,N_8008,N_7422);
or U11086 (N_11086,N_6012,N_7899);
or U11087 (N_11087,N_8137,N_6367);
nand U11088 (N_11088,N_6213,N_7598);
nand U11089 (N_11089,N_7952,N_7489);
and U11090 (N_11090,N_6532,N_7755);
xnor U11091 (N_11091,N_7347,N_7646);
and U11092 (N_11092,N_7571,N_7164);
nor U11093 (N_11093,N_8515,N_6657);
nand U11094 (N_11094,N_7251,N_6851);
nor U11095 (N_11095,N_7947,N_6426);
or U11096 (N_11096,N_6221,N_7546);
and U11097 (N_11097,N_8747,N_6237);
nor U11098 (N_11098,N_8421,N_6281);
or U11099 (N_11099,N_8841,N_6331);
nor U11100 (N_11100,N_6451,N_7486);
or U11101 (N_11101,N_6712,N_8092);
nand U11102 (N_11102,N_6255,N_7444);
and U11103 (N_11103,N_8608,N_8114);
nand U11104 (N_11104,N_7830,N_6034);
and U11105 (N_11105,N_8599,N_6544);
and U11106 (N_11106,N_7758,N_8277);
nand U11107 (N_11107,N_6246,N_6003);
and U11108 (N_11108,N_7188,N_7679);
or U11109 (N_11109,N_7304,N_6545);
and U11110 (N_11110,N_8418,N_7367);
nand U11111 (N_11111,N_6132,N_8426);
and U11112 (N_11112,N_7243,N_6037);
and U11113 (N_11113,N_8297,N_6185);
and U11114 (N_11114,N_7288,N_8489);
xnor U11115 (N_11115,N_8561,N_8462);
nand U11116 (N_11116,N_8905,N_6410);
nor U11117 (N_11117,N_6068,N_6184);
nand U11118 (N_11118,N_8755,N_8842);
nand U11119 (N_11119,N_6546,N_7494);
nand U11120 (N_11120,N_8191,N_7152);
nor U11121 (N_11121,N_6416,N_8362);
and U11122 (N_11122,N_8267,N_6478);
or U11123 (N_11123,N_8211,N_6833);
nand U11124 (N_11124,N_8273,N_8124);
nor U11125 (N_11125,N_7805,N_8916);
or U11126 (N_11126,N_7442,N_6665);
and U11127 (N_11127,N_6395,N_6953);
nand U11128 (N_11128,N_7623,N_7261);
xor U11129 (N_11129,N_8084,N_6892);
nor U11130 (N_11130,N_8010,N_6201);
and U11131 (N_11131,N_8870,N_7654);
and U11132 (N_11132,N_7174,N_7048);
and U11133 (N_11133,N_7236,N_8878);
or U11134 (N_11134,N_7938,N_8783);
and U11135 (N_11135,N_6067,N_7345);
nand U11136 (N_11136,N_6143,N_6190);
nor U11137 (N_11137,N_8675,N_7723);
nand U11138 (N_11138,N_6507,N_7205);
nand U11139 (N_11139,N_8292,N_6263);
nand U11140 (N_11140,N_7858,N_7324);
or U11141 (N_11141,N_8930,N_8213);
nand U11142 (N_11142,N_6171,N_8946);
nand U11143 (N_11143,N_8669,N_7731);
nand U11144 (N_11144,N_6195,N_6351);
nor U11145 (N_11145,N_8859,N_6934);
or U11146 (N_11146,N_8831,N_8463);
xnor U11147 (N_11147,N_6271,N_6549);
or U11148 (N_11148,N_6986,N_7714);
and U11149 (N_11149,N_6961,N_6295);
and U11150 (N_11150,N_8866,N_6870);
or U11151 (N_11151,N_7125,N_8418);
nor U11152 (N_11152,N_8808,N_6889);
nand U11153 (N_11153,N_6909,N_7026);
nand U11154 (N_11154,N_7949,N_7446);
and U11155 (N_11155,N_8659,N_8729);
nor U11156 (N_11156,N_7879,N_7189);
or U11157 (N_11157,N_7840,N_6150);
nand U11158 (N_11158,N_8137,N_8949);
nor U11159 (N_11159,N_7086,N_8351);
nand U11160 (N_11160,N_6233,N_8946);
or U11161 (N_11161,N_8187,N_8020);
and U11162 (N_11162,N_7748,N_6043);
nand U11163 (N_11163,N_8795,N_8425);
and U11164 (N_11164,N_6208,N_8390);
and U11165 (N_11165,N_8224,N_7649);
nor U11166 (N_11166,N_6479,N_7436);
nor U11167 (N_11167,N_6738,N_7675);
and U11168 (N_11168,N_7569,N_6290);
or U11169 (N_11169,N_8035,N_7599);
and U11170 (N_11170,N_6493,N_6626);
and U11171 (N_11171,N_8845,N_8345);
nor U11172 (N_11172,N_7663,N_6403);
nand U11173 (N_11173,N_6163,N_8793);
or U11174 (N_11174,N_7504,N_8634);
or U11175 (N_11175,N_7784,N_6925);
nor U11176 (N_11176,N_8783,N_7273);
nor U11177 (N_11177,N_6650,N_8018);
and U11178 (N_11178,N_8887,N_7431);
nand U11179 (N_11179,N_7947,N_7463);
and U11180 (N_11180,N_6424,N_8891);
nor U11181 (N_11181,N_8098,N_8639);
and U11182 (N_11182,N_6138,N_6169);
nor U11183 (N_11183,N_7216,N_8280);
nor U11184 (N_11184,N_8183,N_8765);
and U11185 (N_11185,N_7227,N_6807);
and U11186 (N_11186,N_6019,N_7689);
nand U11187 (N_11187,N_8642,N_7655);
or U11188 (N_11188,N_6983,N_8328);
or U11189 (N_11189,N_7305,N_6631);
nand U11190 (N_11190,N_7099,N_6361);
nand U11191 (N_11191,N_7040,N_7512);
nand U11192 (N_11192,N_8052,N_6474);
nor U11193 (N_11193,N_7391,N_7696);
nand U11194 (N_11194,N_8562,N_7858);
nand U11195 (N_11195,N_6953,N_6116);
or U11196 (N_11196,N_8584,N_8706);
nor U11197 (N_11197,N_7929,N_8241);
nor U11198 (N_11198,N_6729,N_6063);
nor U11199 (N_11199,N_6570,N_8544);
nand U11200 (N_11200,N_6951,N_6330);
or U11201 (N_11201,N_8811,N_8830);
and U11202 (N_11202,N_7389,N_8075);
nand U11203 (N_11203,N_8078,N_6136);
or U11204 (N_11204,N_7746,N_6041);
or U11205 (N_11205,N_7466,N_6948);
nand U11206 (N_11206,N_6842,N_7279);
nor U11207 (N_11207,N_7757,N_8604);
or U11208 (N_11208,N_6410,N_7736);
and U11209 (N_11209,N_8826,N_6882);
nor U11210 (N_11210,N_8762,N_6340);
or U11211 (N_11211,N_8367,N_6068);
nor U11212 (N_11212,N_7309,N_7829);
nand U11213 (N_11213,N_8150,N_7922);
or U11214 (N_11214,N_8614,N_6936);
nor U11215 (N_11215,N_8571,N_7351);
nand U11216 (N_11216,N_6167,N_7328);
and U11217 (N_11217,N_6953,N_8379);
or U11218 (N_11218,N_6057,N_7411);
or U11219 (N_11219,N_7242,N_7541);
nor U11220 (N_11220,N_7407,N_8040);
nand U11221 (N_11221,N_7036,N_8961);
or U11222 (N_11222,N_6219,N_8655);
nor U11223 (N_11223,N_6316,N_7025);
and U11224 (N_11224,N_7236,N_6909);
nand U11225 (N_11225,N_8193,N_8649);
or U11226 (N_11226,N_7709,N_6950);
nor U11227 (N_11227,N_8175,N_6060);
nand U11228 (N_11228,N_7985,N_6054);
nand U11229 (N_11229,N_8373,N_6257);
nor U11230 (N_11230,N_6307,N_6483);
or U11231 (N_11231,N_7389,N_8925);
nor U11232 (N_11232,N_6313,N_6188);
xnor U11233 (N_11233,N_7002,N_8144);
or U11234 (N_11234,N_6266,N_7931);
and U11235 (N_11235,N_7651,N_7184);
and U11236 (N_11236,N_6548,N_8197);
nand U11237 (N_11237,N_6531,N_8468);
nor U11238 (N_11238,N_8140,N_7835);
or U11239 (N_11239,N_8029,N_8008);
nor U11240 (N_11240,N_8851,N_8424);
or U11241 (N_11241,N_6418,N_8477);
and U11242 (N_11242,N_6137,N_8872);
and U11243 (N_11243,N_8252,N_7058);
or U11244 (N_11244,N_7809,N_8893);
nand U11245 (N_11245,N_8992,N_8701);
or U11246 (N_11246,N_7437,N_6088);
nand U11247 (N_11247,N_6669,N_8923);
nor U11248 (N_11248,N_8372,N_8221);
or U11249 (N_11249,N_8881,N_8523);
and U11250 (N_11250,N_8896,N_8153);
nand U11251 (N_11251,N_6056,N_6405);
nand U11252 (N_11252,N_8720,N_7857);
nand U11253 (N_11253,N_7734,N_8808);
and U11254 (N_11254,N_6962,N_8730);
nand U11255 (N_11255,N_8184,N_6760);
and U11256 (N_11256,N_6476,N_6415);
or U11257 (N_11257,N_7616,N_8825);
or U11258 (N_11258,N_7839,N_8807);
and U11259 (N_11259,N_6984,N_6437);
xor U11260 (N_11260,N_6158,N_6769);
nor U11261 (N_11261,N_6921,N_6355);
nor U11262 (N_11262,N_7662,N_6378);
and U11263 (N_11263,N_7679,N_7347);
nor U11264 (N_11264,N_7589,N_8020);
nor U11265 (N_11265,N_7806,N_8723);
and U11266 (N_11266,N_7331,N_8528);
or U11267 (N_11267,N_7056,N_6235);
nand U11268 (N_11268,N_6306,N_7031);
nand U11269 (N_11269,N_7309,N_6530);
or U11270 (N_11270,N_7897,N_8612);
xnor U11271 (N_11271,N_8100,N_6601);
or U11272 (N_11272,N_6918,N_6646);
nor U11273 (N_11273,N_8463,N_8079);
nor U11274 (N_11274,N_7818,N_8902);
and U11275 (N_11275,N_6025,N_6710);
or U11276 (N_11276,N_7775,N_8548);
and U11277 (N_11277,N_7181,N_8740);
nor U11278 (N_11278,N_6523,N_7469);
nor U11279 (N_11279,N_7993,N_8010);
nand U11280 (N_11280,N_7677,N_6683);
nor U11281 (N_11281,N_7039,N_8971);
and U11282 (N_11282,N_6261,N_8276);
nor U11283 (N_11283,N_7576,N_8639);
and U11284 (N_11284,N_7149,N_6705);
and U11285 (N_11285,N_8797,N_8679);
nor U11286 (N_11286,N_6805,N_6495);
nand U11287 (N_11287,N_8605,N_6039);
or U11288 (N_11288,N_8367,N_8355);
nor U11289 (N_11289,N_7216,N_8761);
nor U11290 (N_11290,N_8601,N_6514);
and U11291 (N_11291,N_8112,N_8786);
and U11292 (N_11292,N_7692,N_7044);
nor U11293 (N_11293,N_7088,N_6036);
nor U11294 (N_11294,N_7552,N_8633);
and U11295 (N_11295,N_6116,N_7924);
nor U11296 (N_11296,N_7605,N_8312);
and U11297 (N_11297,N_8066,N_6728);
or U11298 (N_11298,N_8357,N_6398);
and U11299 (N_11299,N_8069,N_6925);
nand U11300 (N_11300,N_7468,N_7610);
nand U11301 (N_11301,N_8348,N_8304);
nor U11302 (N_11302,N_7872,N_6223);
and U11303 (N_11303,N_7706,N_6666);
nor U11304 (N_11304,N_7600,N_7197);
nand U11305 (N_11305,N_7689,N_6118);
xnor U11306 (N_11306,N_7228,N_7256);
nand U11307 (N_11307,N_7975,N_8530);
and U11308 (N_11308,N_6076,N_8436);
nand U11309 (N_11309,N_6599,N_8338);
nor U11310 (N_11310,N_8829,N_8379);
or U11311 (N_11311,N_7778,N_8825);
nor U11312 (N_11312,N_6721,N_7143);
nor U11313 (N_11313,N_7617,N_8759);
and U11314 (N_11314,N_7476,N_8998);
nand U11315 (N_11315,N_7834,N_6952);
nor U11316 (N_11316,N_8558,N_8307);
nor U11317 (N_11317,N_6113,N_8380);
or U11318 (N_11318,N_8169,N_6638);
nand U11319 (N_11319,N_8162,N_7954);
and U11320 (N_11320,N_6375,N_7372);
nor U11321 (N_11321,N_7089,N_8610);
and U11322 (N_11322,N_8829,N_7465);
and U11323 (N_11323,N_8656,N_8194);
xor U11324 (N_11324,N_8706,N_7584);
or U11325 (N_11325,N_8210,N_7360);
nor U11326 (N_11326,N_8886,N_6755);
xnor U11327 (N_11327,N_6614,N_6705);
or U11328 (N_11328,N_8323,N_8038);
nand U11329 (N_11329,N_6185,N_8779);
nand U11330 (N_11330,N_8732,N_6175);
or U11331 (N_11331,N_6164,N_7505);
or U11332 (N_11332,N_6312,N_8805);
nand U11333 (N_11333,N_6030,N_8888);
nand U11334 (N_11334,N_8100,N_7653);
or U11335 (N_11335,N_8412,N_6498);
nor U11336 (N_11336,N_7543,N_8981);
nor U11337 (N_11337,N_6940,N_6983);
nand U11338 (N_11338,N_7797,N_6309);
nor U11339 (N_11339,N_8344,N_6866);
and U11340 (N_11340,N_7019,N_8045);
nand U11341 (N_11341,N_8078,N_6404);
nor U11342 (N_11342,N_7151,N_7473);
nor U11343 (N_11343,N_8970,N_7342);
and U11344 (N_11344,N_8178,N_7236);
nand U11345 (N_11345,N_8039,N_6974);
nor U11346 (N_11346,N_7489,N_6312);
nand U11347 (N_11347,N_6674,N_8919);
nand U11348 (N_11348,N_6612,N_7366);
nor U11349 (N_11349,N_7442,N_8145);
or U11350 (N_11350,N_6439,N_8495);
nand U11351 (N_11351,N_6157,N_8157);
nor U11352 (N_11352,N_8015,N_8235);
nor U11353 (N_11353,N_8900,N_8721);
and U11354 (N_11354,N_6484,N_8228);
and U11355 (N_11355,N_8207,N_7122);
nand U11356 (N_11356,N_6009,N_7834);
and U11357 (N_11357,N_7281,N_6064);
nor U11358 (N_11358,N_6404,N_8235);
and U11359 (N_11359,N_8007,N_7566);
nor U11360 (N_11360,N_8691,N_6682);
nor U11361 (N_11361,N_7549,N_6783);
or U11362 (N_11362,N_6941,N_7958);
xor U11363 (N_11363,N_6360,N_6466);
and U11364 (N_11364,N_8071,N_7353);
or U11365 (N_11365,N_7712,N_6475);
nand U11366 (N_11366,N_7974,N_7357);
nor U11367 (N_11367,N_6034,N_7645);
nand U11368 (N_11368,N_8610,N_8512);
nand U11369 (N_11369,N_7163,N_7170);
or U11370 (N_11370,N_6816,N_7019);
nor U11371 (N_11371,N_8319,N_7466);
nor U11372 (N_11372,N_8868,N_7763);
and U11373 (N_11373,N_8400,N_7474);
and U11374 (N_11374,N_7601,N_7859);
nand U11375 (N_11375,N_6224,N_7869);
nor U11376 (N_11376,N_6783,N_7632);
nand U11377 (N_11377,N_7721,N_7431);
or U11378 (N_11378,N_6802,N_8719);
and U11379 (N_11379,N_6883,N_7612);
nand U11380 (N_11380,N_8142,N_8439);
nand U11381 (N_11381,N_8202,N_7850);
nand U11382 (N_11382,N_7972,N_7797);
nor U11383 (N_11383,N_8268,N_7278);
nor U11384 (N_11384,N_6095,N_6535);
or U11385 (N_11385,N_6095,N_7536);
xnor U11386 (N_11386,N_6624,N_8250);
nor U11387 (N_11387,N_7370,N_6821);
and U11388 (N_11388,N_7735,N_6783);
nor U11389 (N_11389,N_8581,N_6977);
and U11390 (N_11390,N_7517,N_6631);
and U11391 (N_11391,N_8227,N_6501);
nand U11392 (N_11392,N_7316,N_7573);
nand U11393 (N_11393,N_7751,N_8479);
nand U11394 (N_11394,N_6622,N_8422);
nand U11395 (N_11395,N_7200,N_8344);
nor U11396 (N_11396,N_7516,N_7169);
nand U11397 (N_11397,N_6643,N_7590);
and U11398 (N_11398,N_8912,N_7478);
nor U11399 (N_11399,N_8637,N_6901);
nor U11400 (N_11400,N_6648,N_7320);
and U11401 (N_11401,N_7142,N_7732);
or U11402 (N_11402,N_6523,N_6170);
or U11403 (N_11403,N_7152,N_7674);
and U11404 (N_11404,N_8062,N_6477);
nor U11405 (N_11405,N_7942,N_8208);
and U11406 (N_11406,N_6641,N_7931);
or U11407 (N_11407,N_7422,N_7469);
and U11408 (N_11408,N_7044,N_7294);
and U11409 (N_11409,N_7165,N_7850);
nor U11410 (N_11410,N_7558,N_6782);
or U11411 (N_11411,N_6614,N_8265);
and U11412 (N_11412,N_7372,N_8490);
nor U11413 (N_11413,N_8705,N_6578);
and U11414 (N_11414,N_7592,N_6625);
nor U11415 (N_11415,N_8593,N_8534);
nor U11416 (N_11416,N_8805,N_8015);
or U11417 (N_11417,N_8245,N_7192);
nand U11418 (N_11418,N_7163,N_8360);
and U11419 (N_11419,N_6977,N_7181);
and U11420 (N_11420,N_7225,N_6727);
nand U11421 (N_11421,N_6545,N_7198);
xnor U11422 (N_11422,N_7364,N_8496);
nand U11423 (N_11423,N_6629,N_6585);
or U11424 (N_11424,N_8571,N_6088);
nand U11425 (N_11425,N_7792,N_7769);
nor U11426 (N_11426,N_6929,N_6295);
and U11427 (N_11427,N_8964,N_7499);
nor U11428 (N_11428,N_7706,N_7760);
or U11429 (N_11429,N_8801,N_7962);
nand U11430 (N_11430,N_6290,N_6305);
or U11431 (N_11431,N_7151,N_8023);
and U11432 (N_11432,N_7646,N_8017);
and U11433 (N_11433,N_6107,N_7492);
or U11434 (N_11434,N_8250,N_8912);
nand U11435 (N_11435,N_8429,N_8989);
nor U11436 (N_11436,N_8303,N_7372);
nand U11437 (N_11437,N_7072,N_7746);
nand U11438 (N_11438,N_7318,N_8402);
or U11439 (N_11439,N_6977,N_7853);
or U11440 (N_11440,N_6205,N_7922);
or U11441 (N_11441,N_6183,N_6449);
nor U11442 (N_11442,N_6709,N_8217);
nor U11443 (N_11443,N_7566,N_7934);
and U11444 (N_11444,N_6892,N_7081);
xnor U11445 (N_11445,N_6854,N_7601);
nand U11446 (N_11446,N_6139,N_8137);
or U11447 (N_11447,N_6275,N_6495);
or U11448 (N_11448,N_6310,N_8914);
nor U11449 (N_11449,N_6611,N_6787);
or U11450 (N_11450,N_6482,N_8006);
nand U11451 (N_11451,N_6179,N_6994);
nor U11452 (N_11452,N_7627,N_6370);
or U11453 (N_11453,N_7112,N_6719);
nand U11454 (N_11454,N_8962,N_8845);
nor U11455 (N_11455,N_8652,N_6639);
nor U11456 (N_11456,N_6407,N_6855);
nand U11457 (N_11457,N_8675,N_7621);
nand U11458 (N_11458,N_8377,N_7741);
nor U11459 (N_11459,N_8755,N_7201);
nor U11460 (N_11460,N_7184,N_8373);
and U11461 (N_11461,N_8127,N_6572);
nor U11462 (N_11462,N_8215,N_8824);
nor U11463 (N_11463,N_6785,N_6012);
or U11464 (N_11464,N_8873,N_8704);
or U11465 (N_11465,N_7731,N_6557);
or U11466 (N_11466,N_6969,N_8198);
nor U11467 (N_11467,N_6793,N_6232);
or U11468 (N_11468,N_8851,N_7702);
xnor U11469 (N_11469,N_7777,N_6870);
nor U11470 (N_11470,N_6740,N_6495);
nand U11471 (N_11471,N_7693,N_6729);
nand U11472 (N_11472,N_6002,N_8556);
and U11473 (N_11473,N_6179,N_7510);
nand U11474 (N_11474,N_8585,N_7760);
or U11475 (N_11475,N_7709,N_7970);
and U11476 (N_11476,N_7318,N_8633);
nor U11477 (N_11477,N_8462,N_6925);
or U11478 (N_11478,N_6961,N_8676);
nor U11479 (N_11479,N_8174,N_6982);
nand U11480 (N_11480,N_8550,N_8937);
or U11481 (N_11481,N_6293,N_7816);
or U11482 (N_11482,N_8607,N_6714);
nand U11483 (N_11483,N_7665,N_6556);
or U11484 (N_11484,N_6109,N_8675);
and U11485 (N_11485,N_8553,N_6149);
or U11486 (N_11486,N_6012,N_6392);
nor U11487 (N_11487,N_7939,N_6806);
xnor U11488 (N_11488,N_8003,N_6441);
nor U11489 (N_11489,N_7930,N_7213);
and U11490 (N_11490,N_7035,N_8125);
nand U11491 (N_11491,N_6972,N_6788);
or U11492 (N_11492,N_6749,N_6289);
nor U11493 (N_11493,N_8210,N_7581);
or U11494 (N_11494,N_6170,N_8994);
nor U11495 (N_11495,N_7911,N_7197);
and U11496 (N_11496,N_7514,N_8007);
nand U11497 (N_11497,N_6697,N_8124);
or U11498 (N_11498,N_6610,N_8164);
xnor U11499 (N_11499,N_6895,N_8023);
nand U11500 (N_11500,N_7404,N_8771);
and U11501 (N_11501,N_8777,N_7003);
or U11502 (N_11502,N_7111,N_7863);
or U11503 (N_11503,N_7207,N_8351);
or U11504 (N_11504,N_8710,N_8060);
or U11505 (N_11505,N_8388,N_6189);
and U11506 (N_11506,N_7349,N_6460);
nor U11507 (N_11507,N_6554,N_6000);
nor U11508 (N_11508,N_8364,N_8979);
and U11509 (N_11509,N_8847,N_7866);
or U11510 (N_11510,N_7801,N_8112);
and U11511 (N_11511,N_6808,N_7226);
and U11512 (N_11512,N_8407,N_8415);
nand U11513 (N_11513,N_6117,N_6542);
and U11514 (N_11514,N_6064,N_8648);
or U11515 (N_11515,N_6997,N_7999);
and U11516 (N_11516,N_8198,N_6713);
nor U11517 (N_11517,N_6507,N_7778);
and U11518 (N_11518,N_6315,N_7104);
or U11519 (N_11519,N_7650,N_6523);
and U11520 (N_11520,N_7406,N_7510);
nand U11521 (N_11521,N_7836,N_7715);
nand U11522 (N_11522,N_7658,N_7545);
and U11523 (N_11523,N_8290,N_6771);
or U11524 (N_11524,N_6869,N_6592);
nor U11525 (N_11525,N_6855,N_8053);
nor U11526 (N_11526,N_8443,N_6012);
and U11527 (N_11527,N_8977,N_8505);
xnor U11528 (N_11528,N_6483,N_6192);
nand U11529 (N_11529,N_7480,N_8823);
nand U11530 (N_11530,N_7835,N_7443);
nor U11531 (N_11531,N_8006,N_6388);
and U11532 (N_11532,N_6371,N_8019);
nor U11533 (N_11533,N_8736,N_8799);
or U11534 (N_11534,N_8662,N_7601);
nor U11535 (N_11535,N_7860,N_6763);
and U11536 (N_11536,N_6858,N_8419);
or U11537 (N_11537,N_8943,N_6949);
or U11538 (N_11538,N_7054,N_6855);
or U11539 (N_11539,N_6937,N_6931);
nor U11540 (N_11540,N_6678,N_8260);
and U11541 (N_11541,N_7425,N_7217);
or U11542 (N_11542,N_6878,N_8629);
nand U11543 (N_11543,N_6494,N_8243);
or U11544 (N_11544,N_6772,N_8257);
nand U11545 (N_11545,N_8206,N_6781);
and U11546 (N_11546,N_6105,N_7537);
nand U11547 (N_11547,N_8622,N_6883);
or U11548 (N_11548,N_7239,N_8255);
nand U11549 (N_11549,N_7901,N_6992);
nand U11550 (N_11550,N_8648,N_6902);
nand U11551 (N_11551,N_8365,N_7350);
or U11552 (N_11552,N_7103,N_7100);
nor U11553 (N_11553,N_8369,N_6796);
or U11554 (N_11554,N_7852,N_7881);
and U11555 (N_11555,N_7671,N_8616);
and U11556 (N_11556,N_6508,N_7198);
nand U11557 (N_11557,N_7750,N_8495);
or U11558 (N_11558,N_6990,N_6928);
nand U11559 (N_11559,N_6921,N_8509);
or U11560 (N_11560,N_6222,N_8186);
nor U11561 (N_11561,N_8861,N_8363);
nor U11562 (N_11562,N_6632,N_8245);
or U11563 (N_11563,N_7556,N_6093);
and U11564 (N_11564,N_6951,N_6031);
nand U11565 (N_11565,N_8156,N_8766);
and U11566 (N_11566,N_8814,N_8703);
and U11567 (N_11567,N_7896,N_6901);
nor U11568 (N_11568,N_7900,N_8464);
or U11569 (N_11569,N_7575,N_6494);
nor U11570 (N_11570,N_8562,N_6101);
nand U11571 (N_11571,N_8665,N_7246);
and U11572 (N_11572,N_6524,N_8853);
and U11573 (N_11573,N_7383,N_8530);
nand U11574 (N_11574,N_6903,N_6932);
nor U11575 (N_11575,N_7710,N_6630);
and U11576 (N_11576,N_8528,N_6227);
nand U11577 (N_11577,N_8935,N_7355);
and U11578 (N_11578,N_6116,N_7630);
and U11579 (N_11579,N_7586,N_7945);
nand U11580 (N_11580,N_7218,N_8881);
nor U11581 (N_11581,N_8461,N_7609);
and U11582 (N_11582,N_7561,N_7855);
or U11583 (N_11583,N_7338,N_7954);
nor U11584 (N_11584,N_8393,N_6895);
or U11585 (N_11585,N_7155,N_8337);
and U11586 (N_11586,N_8924,N_7559);
and U11587 (N_11587,N_8839,N_6000);
or U11588 (N_11588,N_7813,N_8591);
nor U11589 (N_11589,N_6747,N_6416);
or U11590 (N_11590,N_8666,N_6189);
nor U11591 (N_11591,N_6395,N_8741);
nor U11592 (N_11592,N_7506,N_7005);
nand U11593 (N_11593,N_8314,N_8240);
and U11594 (N_11594,N_6515,N_6879);
nor U11595 (N_11595,N_6974,N_8599);
nor U11596 (N_11596,N_6256,N_8819);
and U11597 (N_11597,N_6613,N_7135);
nor U11598 (N_11598,N_7575,N_8964);
nor U11599 (N_11599,N_6489,N_6728);
and U11600 (N_11600,N_8167,N_6305);
nor U11601 (N_11601,N_6530,N_7094);
nor U11602 (N_11602,N_6943,N_6008);
or U11603 (N_11603,N_6088,N_6055);
nor U11604 (N_11604,N_7808,N_7303);
and U11605 (N_11605,N_7782,N_6961);
and U11606 (N_11606,N_8478,N_7002);
and U11607 (N_11607,N_8771,N_8113);
nand U11608 (N_11608,N_6659,N_7999);
nand U11609 (N_11609,N_6278,N_6329);
or U11610 (N_11610,N_8443,N_8719);
nand U11611 (N_11611,N_7476,N_6042);
and U11612 (N_11612,N_8183,N_7380);
or U11613 (N_11613,N_6462,N_6381);
or U11614 (N_11614,N_6565,N_7310);
nor U11615 (N_11615,N_7533,N_6046);
nor U11616 (N_11616,N_7716,N_8856);
nand U11617 (N_11617,N_7748,N_7848);
nand U11618 (N_11618,N_7784,N_7321);
nor U11619 (N_11619,N_8541,N_6000);
and U11620 (N_11620,N_8156,N_6599);
or U11621 (N_11621,N_6496,N_8592);
or U11622 (N_11622,N_6833,N_7534);
nand U11623 (N_11623,N_7695,N_7861);
or U11624 (N_11624,N_8772,N_7923);
nand U11625 (N_11625,N_8973,N_8889);
nor U11626 (N_11626,N_7563,N_8654);
and U11627 (N_11627,N_8282,N_6305);
xor U11628 (N_11628,N_6267,N_6834);
and U11629 (N_11629,N_6819,N_6692);
and U11630 (N_11630,N_8950,N_8447);
nor U11631 (N_11631,N_7732,N_7939);
or U11632 (N_11632,N_8953,N_8161);
or U11633 (N_11633,N_6474,N_7929);
nor U11634 (N_11634,N_8549,N_6352);
or U11635 (N_11635,N_7323,N_6950);
nor U11636 (N_11636,N_6201,N_8505);
nor U11637 (N_11637,N_8751,N_7107);
and U11638 (N_11638,N_8504,N_7492);
nor U11639 (N_11639,N_6403,N_7135);
and U11640 (N_11640,N_8873,N_7945);
or U11641 (N_11641,N_6030,N_6432);
nand U11642 (N_11642,N_6128,N_8480);
nand U11643 (N_11643,N_8648,N_6482);
or U11644 (N_11644,N_6347,N_7939);
nand U11645 (N_11645,N_7418,N_7145);
nor U11646 (N_11646,N_8138,N_6288);
nor U11647 (N_11647,N_7936,N_8630);
nand U11648 (N_11648,N_8669,N_8058);
and U11649 (N_11649,N_6441,N_6915);
or U11650 (N_11650,N_6779,N_8301);
or U11651 (N_11651,N_7170,N_8201);
and U11652 (N_11652,N_7344,N_7506);
or U11653 (N_11653,N_6283,N_8587);
nor U11654 (N_11654,N_8839,N_7147);
nand U11655 (N_11655,N_7908,N_6273);
or U11656 (N_11656,N_7650,N_6517);
nor U11657 (N_11657,N_8520,N_7135);
nor U11658 (N_11658,N_8224,N_7459);
and U11659 (N_11659,N_7303,N_7088);
nand U11660 (N_11660,N_8621,N_8142);
and U11661 (N_11661,N_6098,N_6442);
nand U11662 (N_11662,N_8598,N_8048);
nor U11663 (N_11663,N_7829,N_6634);
or U11664 (N_11664,N_8581,N_8217);
nand U11665 (N_11665,N_7281,N_8157);
nor U11666 (N_11666,N_8707,N_6839);
or U11667 (N_11667,N_8263,N_6990);
nor U11668 (N_11668,N_8660,N_7643);
nor U11669 (N_11669,N_8280,N_7432);
and U11670 (N_11670,N_6023,N_8017);
and U11671 (N_11671,N_8074,N_6454);
nand U11672 (N_11672,N_8030,N_8752);
or U11673 (N_11673,N_8698,N_7908);
nor U11674 (N_11674,N_8091,N_7115);
nor U11675 (N_11675,N_6480,N_8860);
nand U11676 (N_11676,N_8077,N_6826);
nor U11677 (N_11677,N_7868,N_8574);
and U11678 (N_11678,N_8706,N_7559);
and U11679 (N_11679,N_6650,N_7300);
and U11680 (N_11680,N_6953,N_7910);
nand U11681 (N_11681,N_8117,N_6411);
nand U11682 (N_11682,N_8932,N_7040);
nor U11683 (N_11683,N_6971,N_7695);
nor U11684 (N_11684,N_6489,N_8086);
or U11685 (N_11685,N_6606,N_7148);
nor U11686 (N_11686,N_6182,N_6716);
nand U11687 (N_11687,N_6612,N_6989);
or U11688 (N_11688,N_8409,N_7375);
nand U11689 (N_11689,N_6447,N_7683);
and U11690 (N_11690,N_6635,N_7920);
and U11691 (N_11691,N_6138,N_8235);
or U11692 (N_11692,N_6727,N_8764);
nand U11693 (N_11693,N_7139,N_6308);
nand U11694 (N_11694,N_8510,N_6228);
and U11695 (N_11695,N_8988,N_7757);
nor U11696 (N_11696,N_7183,N_6659);
nand U11697 (N_11697,N_6849,N_7151);
and U11698 (N_11698,N_7704,N_8407);
or U11699 (N_11699,N_7906,N_7585);
or U11700 (N_11700,N_7637,N_8183);
or U11701 (N_11701,N_6428,N_8083);
and U11702 (N_11702,N_7623,N_8178);
or U11703 (N_11703,N_6719,N_8987);
and U11704 (N_11704,N_6532,N_8923);
or U11705 (N_11705,N_8479,N_6953);
nand U11706 (N_11706,N_8694,N_6013);
nor U11707 (N_11707,N_7426,N_8905);
nand U11708 (N_11708,N_7937,N_6180);
and U11709 (N_11709,N_6793,N_8015);
nand U11710 (N_11710,N_6881,N_6175);
nand U11711 (N_11711,N_8434,N_6862);
nor U11712 (N_11712,N_8373,N_8224);
and U11713 (N_11713,N_6778,N_8020);
or U11714 (N_11714,N_6014,N_6407);
or U11715 (N_11715,N_8621,N_7228);
nand U11716 (N_11716,N_8657,N_6511);
and U11717 (N_11717,N_6795,N_8126);
or U11718 (N_11718,N_6409,N_6098);
xnor U11719 (N_11719,N_7145,N_8690);
nor U11720 (N_11720,N_6874,N_8895);
or U11721 (N_11721,N_6575,N_8445);
or U11722 (N_11722,N_8964,N_8506);
and U11723 (N_11723,N_6430,N_6429);
and U11724 (N_11724,N_6453,N_6467);
and U11725 (N_11725,N_7460,N_8786);
and U11726 (N_11726,N_6441,N_6734);
or U11727 (N_11727,N_8339,N_7361);
and U11728 (N_11728,N_8804,N_7260);
nand U11729 (N_11729,N_6320,N_8330);
or U11730 (N_11730,N_6925,N_6405);
nor U11731 (N_11731,N_7435,N_7874);
and U11732 (N_11732,N_7600,N_7792);
nor U11733 (N_11733,N_6460,N_6849);
nand U11734 (N_11734,N_7620,N_8874);
nand U11735 (N_11735,N_6423,N_7978);
or U11736 (N_11736,N_6111,N_6687);
nand U11737 (N_11737,N_8129,N_8064);
xor U11738 (N_11738,N_8902,N_6544);
and U11739 (N_11739,N_8460,N_6902);
nand U11740 (N_11740,N_6513,N_7640);
nand U11741 (N_11741,N_7251,N_7380);
or U11742 (N_11742,N_8288,N_6577);
nand U11743 (N_11743,N_8123,N_8211);
nand U11744 (N_11744,N_8023,N_6553);
or U11745 (N_11745,N_7565,N_8841);
or U11746 (N_11746,N_7195,N_7700);
nor U11747 (N_11747,N_8237,N_8661);
and U11748 (N_11748,N_7441,N_6708);
or U11749 (N_11749,N_8566,N_7711);
nand U11750 (N_11750,N_6326,N_7310);
nand U11751 (N_11751,N_8156,N_8157);
and U11752 (N_11752,N_6763,N_7241);
xnor U11753 (N_11753,N_6253,N_7868);
nand U11754 (N_11754,N_6396,N_8809);
nor U11755 (N_11755,N_7927,N_7910);
and U11756 (N_11756,N_6177,N_7079);
nor U11757 (N_11757,N_7206,N_8857);
nor U11758 (N_11758,N_8036,N_6709);
and U11759 (N_11759,N_7198,N_8774);
nand U11760 (N_11760,N_6418,N_7944);
or U11761 (N_11761,N_8128,N_6854);
nand U11762 (N_11762,N_6341,N_6168);
nor U11763 (N_11763,N_7208,N_7808);
nand U11764 (N_11764,N_8971,N_6919);
and U11765 (N_11765,N_6309,N_7881);
or U11766 (N_11766,N_7566,N_6949);
nand U11767 (N_11767,N_6768,N_6615);
nor U11768 (N_11768,N_6106,N_6607);
nor U11769 (N_11769,N_7545,N_7187);
or U11770 (N_11770,N_6670,N_6159);
nor U11771 (N_11771,N_6739,N_8938);
nand U11772 (N_11772,N_6099,N_8786);
nand U11773 (N_11773,N_8980,N_6030);
or U11774 (N_11774,N_7392,N_7538);
nor U11775 (N_11775,N_8356,N_7029);
nand U11776 (N_11776,N_7825,N_6162);
or U11777 (N_11777,N_6125,N_7374);
and U11778 (N_11778,N_6997,N_8524);
or U11779 (N_11779,N_7644,N_8302);
or U11780 (N_11780,N_7451,N_8264);
nand U11781 (N_11781,N_8161,N_7460);
or U11782 (N_11782,N_8870,N_7831);
nor U11783 (N_11783,N_7962,N_6675);
and U11784 (N_11784,N_7150,N_7771);
nor U11785 (N_11785,N_6141,N_8630);
and U11786 (N_11786,N_8849,N_6124);
and U11787 (N_11787,N_8280,N_7586);
nor U11788 (N_11788,N_6226,N_7280);
nand U11789 (N_11789,N_7527,N_6730);
nor U11790 (N_11790,N_7090,N_7043);
xnor U11791 (N_11791,N_6841,N_6160);
nor U11792 (N_11792,N_8381,N_6583);
or U11793 (N_11793,N_7702,N_6575);
or U11794 (N_11794,N_8684,N_7740);
nand U11795 (N_11795,N_8010,N_8441);
nor U11796 (N_11796,N_8859,N_7221);
nor U11797 (N_11797,N_7041,N_8964);
nor U11798 (N_11798,N_7979,N_6790);
nand U11799 (N_11799,N_7821,N_8925);
nand U11800 (N_11800,N_7238,N_7307);
nor U11801 (N_11801,N_7319,N_7800);
xnor U11802 (N_11802,N_8844,N_6586);
and U11803 (N_11803,N_7171,N_6663);
and U11804 (N_11804,N_6027,N_6319);
and U11805 (N_11805,N_7395,N_6099);
or U11806 (N_11806,N_6608,N_7511);
and U11807 (N_11807,N_8652,N_8425);
nor U11808 (N_11808,N_7537,N_8241);
and U11809 (N_11809,N_8451,N_8749);
or U11810 (N_11810,N_8968,N_7381);
or U11811 (N_11811,N_6381,N_7262);
and U11812 (N_11812,N_8144,N_7279);
nor U11813 (N_11813,N_7172,N_7024);
or U11814 (N_11814,N_6559,N_7028);
or U11815 (N_11815,N_6916,N_8851);
nor U11816 (N_11816,N_7849,N_7069);
nand U11817 (N_11817,N_6404,N_8368);
and U11818 (N_11818,N_7154,N_8958);
xnor U11819 (N_11819,N_6217,N_8311);
nor U11820 (N_11820,N_8571,N_8488);
nor U11821 (N_11821,N_7047,N_7760);
nor U11822 (N_11822,N_6883,N_6182);
or U11823 (N_11823,N_8313,N_6721);
and U11824 (N_11824,N_6688,N_6090);
and U11825 (N_11825,N_8712,N_8869);
nand U11826 (N_11826,N_8136,N_6194);
xnor U11827 (N_11827,N_8734,N_8458);
and U11828 (N_11828,N_7990,N_6107);
or U11829 (N_11829,N_6688,N_8580);
and U11830 (N_11830,N_8863,N_8322);
and U11831 (N_11831,N_6045,N_7477);
or U11832 (N_11832,N_6896,N_6713);
or U11833 (N_11833,N_8962,N_7629);
nand U11834 (N_11834,N_6818,N_6283);
nor U11835 (N_11835,N_6072,N_8554);
and U11836 (N_11836,N_8403,N_7289);
or U11837 (N_11837,N_6493,N_8402);
and U11838 (N_11838,N_7504,N_8707);
and U11839 (N_11839,N_8039,N_8926);
nor U11840 (N_11840,N_6644,N_7329);
nor U11841 (N_11841,N_7275,N_6796);
nand U11842 (N_11842,N_6053,N_7294);
nor U11843 (N_11843,N_8574,N_7498);
nand U11844 (N_11844,N_7142,N_7025);
xnor U11845 (N_11845,N_8635,N_7828);
nor U11846 (N_11846,N_8126,N_7582);
nand U11847 (N_11847,N_7393,N_6213);
and U11848 (N_11848,N_7920,N_6745);
nand U11849 (N_11849,N_6161,N_7370);
or U11850 (N_11850,N_7708,N_7961);
nor U11851 (N_11851,N_6568,N_8679);
nor U11852 (N_11852,N_6651,N_6661);
and U11853 (N_11853,N_7307,N_8233);
and U11854 (N_11854,N_7492,N_6627);
nor U11855 (N_11855,N_8359,N_6250);
or U11856 (N_11856,N_6706,N_6998);
nor U11857 (N_11857,N_6151,N_8118);
nor U11858 (N_11858,N_7246,N_6357);
nand U11859 (N_11859,N_6216,N_8347);
and U11860 (N_11860,N_7477,N_8629);
or U11861 (N_11861,N_7305,N_6134);
and U11862 (N_11862,N_7440,N_7216);
and U11863 (N_11863,N_6289,N_6666);
nand U11864 (N_11864,N_6821,N_8489);
nand U11865 (N_11865,N_7277,N_6555);
or U11866 (N_11866,N_7573,N_6814);
or U11867 (N_11867,N_7676,N_6125);
nand U11868 (N_11868,N_6445,N_7943);
nand U11869 (N_11869,N_7559,N_7468);
nand U11870 (N_11870,N_8983,N_6814);
and U11871 (N_11871,N_8248,N_7767);
or U11872 (N_11872,N_8999,N_8642);
nor U11873 (N_11873,N_8366,N_6277);
and U11874 (N_11874,N_8773,N_7050);
nand U11875 (N_11875,N_6287,N_8464);
and U11876 (N_11876,N_6859,N_7522);
nand U11877 (N_11877,N_8915,N_7636);
nand U11878 (N_11878,N_8762,N_8788);
and U11879 (N_11879,N_7917,N_7482);
or U11880 (N_11880,N_6346,N_6712);
nor U11881 (N_11881,N_8255,N_6845);
and U11882 (N_11882,N_8246,N_6370);
and U11883 (N_11883,N_8191,N_8309);
nor U11884 (N_11884,N_6678,N_6398);
and U11885 (N_11885,N_8212,N_6735);
or U11886 (N_11886,N_6654,N_8132);
nor U11887 (N_11887,N_8109,N_6588);
and U11888 (N_11888,N_6484,N_7300);
and U11889 (N_11889,N_8720,N_6700);
and U11890 (N_11890,N_8320,N_7504);
and U11891 (N_11891,N_8915,N_7189);
nand U11892 (N_11892,N_8014,N_6857);
or U11893 (N_11893,N_7832,N_8709);
and U11894 (N_11894,N_8276,N_8469);
or U11895 (N_11895,N_8721,N_7976);
and U11896 (N_11896,N_8150,N_6106);
and U11897 (N_11897,N_7905,N_8387);
nand U11898 (N_11898,N_8116,N_8561);
nor U11899 (N_11899,N_7539,N_8331);
and U11900 (N_11900,N_7189,N_7176);
nor U11901 (N_11901,N_7936,N_7973);
nor U11902 (N_11902,N_7088,N_6714);
nand U11903 (N_11903,N_8513,N_7373);
nor U11904 (N_11904,N_7159,N_7780);
xor U11905 (N_11905,N_7260,N_7196);
or U11906 (N_11906,N_6568,N_7423);
nand U11907 (N_11907,N_6354,N_7082);
nor U11908 (N_11908,N_7759,N_8057);
nor U11909 (N_11909,N_7190,N_6677);
nor U11910 (N_11910,N_6572,N_7969);
nand U11911 (N_11911,N_8410,N_8053);
and U11912 (N_11912,N_8882,N_8552);
and U11913 (N_11913,N_7434,N_7234);
and U11914 (N_11914,N_6269,N_6294);
nor U11915 (N_11915,N_6716,N_6729);
nor U11916 (N_11916,N_7510,N_8300);
nand U11917 (N_11917,N_6435,N_8340);
nand U11918 (N_11918,N_7140,N_6923);
nor U11919 (N_11919,N_6552,N_7234);
nor U11920 (N_11920,N_7900,N_6619);
or U11921 (N_11921,N_8164,N_7204);
nor U11922 (N_11922,N_7689,N_8496);
and U11923 (N_11923,N_7373,N_7478);
and U11924 (N_11924,N_8736,N_8487);
or U11925 (N_11925,N_7142,N_7996);
and U11926 (N_11926,N_6991,N_8809);
or U11927 (N_11927,N_8705,N_8924);
and U11928 (N_11928,N_6713,N_6102);
and U11929 (N_11929,N_8930,N_7596);
and U11930 (N_11930,N_6132,N_6628);
nor U11931 (N_11931,N_6752,N_7281);
nor U11932 (N_11932,N_7427,N_8569);
nand U11933 (N_11933,N_6044,N_6457);
and U11934 (N_11934,N_7062,N_6694);
nor U11935 (N_11935,N_8738,N_8623);
nor U11936 (N_11936,N_6309,N_7476);
nor U11937 (N_11937,N_8247,N_8721);
nor U11938 (N_11938,N_7389,N_7952);
nor U11939 (N_11939,N_8384,N_7641);
and U11940 (N_11940,N_8751,N_7637);
or U11941 (N_11941,N_7968,N_8306);
nor U11942 (N_11942,N_6093,N_7986);
or U11943 (N_11943,N_7869,N_7036);
nor U11944 (N_11944,N_8100,N_6648);
nand U11945 (N_11945,N_7641,N_8698);
or U11946 (N_11946,N_7039,N_7995);
xnor U11947 (N_11947,N_7690,N_7785);
and U11948 (N_11948,N_8127,N_7554);
nor U11949 (N_11949,N_7600,N_7562);
and U11950 (N_11950,N_7769,N_6987);
nor U11951 (N_11951,N_8858,N_7168);
nor U11952 (N_11952,N_8164,N_7281);
nand U11953 (N_11953,N_7344,N_7146);
or U11954 (N_11954,N_6223,N_8713);
or U11955 (N_11955,N_8342,N_7275);
nor U11956 (N_11956,N_7904,N_8283);
and U11957 (N_11957,N_8658,N_6179);
or U11958 (N_11958,N_8371,N_6015);
or U11959 (N_11959,N_8351,N_7314);
nor U11960 (N_11960,N_8100,N_8392);
nand U11961 (N_11961,N_7898,N_6427);
and U11962 (N_11962,N_6231,N_7522);
nand U11963 (N_11963,N_6683,N_8772);
nand U11964 (N_11964,N_7444,N_8428);
nand U11965 (N_11965,N_8160,N_8382);
or U11966 (N_11966,N_8061,N_7777);
and U11967 (N_11967,N_8214,N_8875);
nor U11968 (N_11968,N_6932,N_7081);
and U11969 (N_11969,N_6495,N_6873);
nor U11970 (N_11970,N_7842,N_6483);
nor U11971 (N_11971,N_7760,N_6008);
and U11972 (N_11972,N_7513,N_6186);
nand U11973 (N_11973,N_8096,N_7214);
nor U11974 (N_11974,N_6326,N_7302);
nor U11975 (N_11975,N_6604,N_7812);
nor U11976 (N_11976,N_6370,N_8769);
or U11977 (N_11977,N_7880,N_7240);
or U11978 (N_11978,N_8798,N_7236);
or U11979 (N_11979,N_7365,N_8351);
and U11980 (N_11980,N_8085,N_7415);
nor U11981 (N_11981,N_7806,N_7900);
and U11982 (N_11982,N_7005,N_6811);
nor U11983 (N_11983,N_7042,N_8947);
and U11984 (N_11984,N_6616,N_7417);
nand U11985 (N_11985,N_7964,N_6582);
xnor U11986 (N_11986,N_8997,N_8487);
nor U11987 (N_11987,N_6847,N_8351);
and U11988 (N_11988,N_8589,N_7976);
and U11989 (N_11989,N_7704,N_7528);
nand U11990 (N_11990,N_6823,N_6767);
or U11991 (N_11991,N_7043,N_6377);
and U11992 (N_11992,N_7209,N_6685);
nor U11993 (N_11993,N_7990,N_8343);
nand U11994 (N_11994,N_6587,N_7162);
nor U11995 (N_11995,N_7523,N_8020);
nor U11996 (N_11996,N_6315,N_6622);
and U11997 (N_11997,N_6991,N_6767);
and U11998 (N_11998,N_7615,N_6020);
nand U11999 (N_11999,N_6687,N_8167);
xor U12000 (N_12000,N_10201,N_11207);
nor U12001 (N_12001,N_11572,N_11045);
nand U12002 (N_12002,N_11694,N_10436);
nor U12003 (N_12003,N_9993,N_9525);
nand U12004 (N_12004,N_9391,N_10129);
and U12005 (N_12005,N_9953,N_11157);
or U12006 (N_12006,N_11283,N_10065);
nor U12007 (N_12007,N_11054,N_11604);
nor U12008 (N_12008,N_11715,N_9755);
nand U12009 (N_12009,N_9902,N_11146);
nor U12010 (N_12010,N_10170,N_9783);
nand U12011 (N_12011,N_10137,N_11427);
or U12012 (N_12012,N_10697,N_9785);
nand U12013 (N_12013,N_11131,N_9269);
or U12014 (N_12014,N_10670,N_11184);
nor U12015 (N_12015,N_9750,N_9363);
nor U12016 (N_12016,N_9157,N_11527);
or U12017 (N_12017,N_9610,N_11060);
nand U12018 (N_12018,N_10557,N_10844);
or U12019 (N_12019,N_10875,N_9367);
and U12020 (N_12020,N_9218,N_10612);
or U12021 (N_12021,N_11410,N_9686);
and U12022 (N_12022,N_9480,N_10410);
or U12023 (N_12023,N_11957,N_11798);
or U12024 (N_12024,N_9105,N_9547);
nor U12025 (N_12025,N_11423,N_11325);
nor U12026 (N_12026,N_11387,N_10125);
nor U12027 (N_12027,N_9456,N_11154);
or U12028 (N_12028,N_11679,N_10099);
or U12029 (N_12029,N_9256,N_9650);
nand U12030 (N_12030,N_9912,N_11964);
xnor U12031 (N_12031,N_9703,N_11804);
or U12032 (N_12032,N_11087,N_9243);
nand U12033 (N_12033,N_10668,N_10925);
nand U12034 (N_12034,N_9837,N_11021);
nand U12035 (N_12035,N_11809,N_11185);
nand U12036 (N_12036,N_10705,N_10495);
nor U12037 (N_12037,N_11823,N_9466);
or U12038 (N_12038,N_11240,N_9962);
nor U12039 (N_12039,N_11033,N_11611);
nand U12040 (N_12040,N_10744,N_11269);
and U12041 (N_12041,N_9581,N_11379);
nand U12042 (N_12042,N_9145,N_11331);
nor U12043 (N_12043,N_10823,N_10822);
and U12044 (N_12044,N_11908,N_10117);
or U12045 (N_12045,N_11554,N_10837);
nand U12046 (N_12046,N_10763,N_10360);
nand U12047 (N_12047,N_9676,N_11357);
and U12048 (N_12048,N_11195,N_11663);
and U12049 (N_12049,N_11291,N_11987);
nor U12050 (N_12050,N_10511,N_9245);
nor U12051 (N_12051,N_9146,N_11512);
and U12052 (N_12052,N_9536,N_11229);
or U12053 (N_12053,N_11392,N_11210);
or U12054 (N_12054,N_10838,N_10419);
nor U12055 (N_12055,N_9098,N_11655);
nor U12056 (N_12056,N_10832,N_10627);
and U12057 (N_12057,N_10813,N_10055);
xor U12058 (N_12058,N_10874,N_11876);
xnor U12059 (N_12059,N_9784,N_11488);
or U12060 (N_12060,N_9636,N_10082);
nor U12061 (N_12061,N_11874,N_9955);
nand U12062 (N_12062,N_10262,N_11298);
nor U12063 (N_12063,N_10275,N_11647);
nor U12064 (N_12064,N_9726,N_11485);
nand U12065 (N_12065,N_11413,N_11481);
or U12066 (N_12066,N_10255,N_9501);
or U12067 (N_12067,N_10302,N_9317);
nor U12068 (N_12068,N_9402,N_11913);
nand U12069 (N_12069,N_10138,N_10184);
and U12070 (N_12070,N_11993,N_11175);
nand U12071 (N_12071,N_9896,N_10250);
and U12072 (N_12072,N_11729,N_11539);
or U12073 (N_12073,N_9596,N_9436);
and U12074 (N_12074,N_10634,N_9021);
nor U12075 (N_12075,N_9043,N_11634);
nor U12076 (N_12076,N_11955,N_10672);
and U12077 (N_12077,N_9879,N_9813);
and U12078 (N_12078,N_10206,N_9980);
nand U12079 (N_12079,N_9376,N_9476);
nor U12080 (N_12080,N_11199,N_10268);
or U12081 (N_12081,N_10828,N_9081);
or U12082 (N_12082,N_11119,N_10260);
nand U12083 (N_12083,N_10816,N_10377);
nor U12084 (N_12084,N_11305,N_11954);
nand U12085 (N_12085,N_11447,N_9004);
nand U12086 (N_12086,N_11575,N_9624);
nand U12087 (N_12087,N_11228,N_9121);
nand U12088 (N_12088,N_11275,N_10328);
and U12089 (N_12089,N_10873,N_11577);
and U12090 (N_12090,N_11100,N_11134);
nor U12091 (N_12091,N_10718,N_11330);
or U12092 (N_12092,N_9926,N_11368);
or U12093 (N_12093,N_11123,N_10251);
nor U12094 (N_12094,N_11998,N_11983);
or U12095 (N_12095,N_9278,N_11311);
nor U12096 (N_12096,N_9803,N_10113);
or U12097 (N_12097,N_11942,N_9116);
nand U12098 (N_12098,N_9080,N_10247);
or U12099 (N_12099,N_9205,N_11280);
nor U12100 (N_12100,N_10717,N_9776);
and U12101 (N_12101,N_9297,N_10437);
and U12102 (N_12102,N_9066,N_11419);
nand U12103 (N_12103,N_11276,N_10076);
or U12104 (N_12104,N_9621,N_9568);
or U12105 (N_12105,N_10997,N_9746);
and U12106 (N_12106,N_10870,N_10062);
and U12107 (N_12107,N_9756,N_11989);
or U12108 (N_12108,N_11927,N_9348);
nor U12109 (N_12109,N_10265,N_11069);
nor U12110 (N_12110,N_10485,N_9869);
nor U12111 (N_12111,N_10347,N_10330);
or U12112 (N_12112,N_9576,N_10343);
nand U12113 (N_12113,N_11500,N_11863);
nand U12114 (N_12114,N_9469,N_10001);
and U12115 (N_12115,N_9370,N_10010);
nor U12116 (N_12116,N_9625,N_9031);
and U12117 (N_12117,N_10514,N_9129);
or U12118 (N_12118,N_11828,N_10590);
nor U12119 (N_12119,N_10415,N_9407);
nor U12120 (N_12120,N_11141,N_11439);
and U12121 (N_12121,N_10715,N_11264);
nor U12122 (N_12122,N_10094,N_11681);
or U12123 (N_12123,N_10887,N_9194);
xnor U12124 (N_12124,N_10968,N_10957);
nor U12125 (N_12125,N_9384,N_9274);
nand U12126 (N_12126,N_11349,N_11560);
and U12127 (N_12127,N_9214,N_10522);
nand U12128 (N_12128,N_11643,N_10596);
nor U12129 (N_12129,N_9488,N_9207);
nor U12130 (N_12130,N_9174,N_11053);
or U12131 (N_12131,N_11181,N_9571);
or U12132 (N_12132,N_11990,N_9800);
nand U12133 (N_12133,N_11599,N_9575);
and U12134 (N_12134,N_10509,N_10897);
or U12135 (N_12135,N_10123,N_9110);
or U12136 (N_12136,N_11347,N_11108);
or U12137 (N_12137,N_10981,N_9851);
or U12138 (N_12138,N_9286,N_9362);
or U12139 (N_12139,N_10329,N_11630);
nor U12140 (N_12140,N_9343,N_9818);
and U12141 (N_12141,N_10257,N_11057);
xor U12142 (N_12142,N_11846,N_11056);
nand U12143 (N_12143,N_10909,N_10673);
and U12144 (N_12144,N_9169,N_10043);
nor U12145 (N_12145,N_11180,N_10620);
nand U12146 (N_12146,N_11139,N_10190);
nor U12147 (N_12147,N_11718,N_11683);
nor U12148 (N_12148,N_10573,N_11084);
nor U12149 (N_12149,N_10397,N_9615);
or U12150 (N_12150,N_11140,N_11462);
nand U12151 (N_12151,N_11487,N_10176);
and U12152 (N_12152,N_10479,N_10526);
or U12153 (N_12153,N_11548,N_9210);
and U12154 (N_12154,N_10594,N_9984);
nor U12155 (N_12155,N_11509,N_10417);
nor U12156 (N_12156,N_9016,N_11710);
or U12157 (N_12157,N_9695,N_10505);
nand U12158 (N_12158,N_9874,N_10142);
or U12159 (N_12159,N_11104,N_10621);
and U12160 (N_12160,N_9112,N_10578);
nand U12161 (N_12161,N_10466,N_9234);
or U12162 (N_12162,N_9607,N_9449);
nand U12163 (N_12163,N_11594,N_9414);
and U12164 (N_12164,N_10233,N_11915);
or U12165 (N_12165,N_10795,N_11922);
or U12166 (N_12166,N_10236,N_9171);
nor U12167 (N_12167,N_11428,N_9713);
nand U12168 (N_12168,N_9345,N_10779);
and U12169 (N_12169,N_11531,N_9462);
or U12170 (N_12170,N_11564,N_10753);
and U12171 (N_12171,N_9061,N_11832);
nor U12172 (N_12172,N_11351,N_10973);
nor U12173 (N_12173,N_11274,N_9415);
nor U12174 (N_12174,N_10216,N_9511);
nand U12175 (N_12175,N_11969,N_10711);
and U12176 (N_12176,N_11083,N_11189);
or U12177 (N_12177,N_11711,N_10311);
and U12178 (N_12178,N_11085,N_10426);
xor U12179 (N_12179,N_9251,N_11742);
nor U12180 (N_12180,N_9564,N_9059);
or U12181 (N_12181,N_9326,N_10323);
or U12182 (N_12182,N_10198,N_9058);
and U12183 (N_12183,N_9117,N_10563);
nand U12184 (N_12184,N_11415,N_11639);
nor U12185 (N_12185,N_10295,N_11565);
nand U12186 (N_12186,N_10308,N_11511);
or U12187 (N_12187,N_10631,N_9339);
nor U12188 (N_12188,N_10508,N_9073);
nand U12189 (N_12189,N_9288,N_10034);
nand U12190 (N_12190,N_11338,N_10224);
nor U12191 (N_12191,N_10127,N_10011);
and U12192 (N_12192,N_11938,N_11029);
nand U12193 (N_12193,N_11994,N_11297);
nor U12194 (N_12194,N_9669,N_9114);
nor U12195 (N_12195,N_9573,N_11177);
nand U12196 (N_12196,N_9196,N_9787);
and U12197 (N_12197,N_9316,N_9392);
nor U12198 (N_12198,N_10455,N_11573);
nand U12199 (N_12199,N_10244,N_10588);
and U12200 (N_12200,N_11595,N_11707);
nor U12201 (N_12201,N_11656,N_10685);
nand U12202 (N_12202,N_9753,N_10222);
and U12203 (N_12203,N_9313,N_10956);
nand U12204 (N_12204,N_10133,N_10856);
and U12205 (N_12205,N_9089,N_11748);
nand U12206 (N_12206,N_10452,N_9730);
nand U12207 (N_12207,N_11765,N_11926);
xor U12208 (N_12208,N_11609,N_9029);
nor U12209 (N_12209,N_10263,N_10453);
and U12210 (N_12210,N_11225,N_10183);
and U12211 (N_12211,N_9211,N_9855);
nand U12212 (N_12212,N_10618,N_9594);
or U12213 (N_12213,N_10387,N_11321);
or U12214 (N_12214,N_9050,N_9794);
nand U12215 (N_12215,N_9007,N_11557);
or U12216 (N_12216,N_11975,N_10205);
nand U12217 (N_12217,N_9190,N_11695);
or U12218 (N_12218,N_9802,N_9508);
nand U12219 (N_12219,N_9053,N_11925);
nand U12220 (N_12220,N_9033,N_11246);
nor U12221 (N_12221,N_10691,N_11992);
nand U12222 (N_12222,N_11991,N_10248);
nand U12223 (N_12223,N_9679,N_10995);
and U12224 (N_12224,N_10615,N_11310);
nor U12225 (N_12225,N_10309,N_11206);
and U12226 (N_12226,N_10507,N_11224);
or U12227 (N_12227,N_9118,N_11179);
or U12228 (N_12228,N_10282,N_9170);
nand U12229 (N_12229,N_11783,N_10407);
nand U12230 (N_12230,N_10405,N_9461);
nand U12231 (N_12231,N_9934,N_11380);
and U12232 (N_12232,N_11172,N_9412);
and U12233 (N_12233,N_11543,N_10904);
nor U12234 (N_12234,N_10154,N_9947);
nor U12235 (N_12235,N_10338,N_11799);
or U12236 (N_12236,N_10824,N_10100);
and U12237 (N_12237,N_11308,N_9270);
and U12238 (N_12238,N_10081,N_10132);
and U12239 (N_12239,N_9123,N_10105);
or U12240 (N_12240,N_9433,N_9260);
or U12241 (N_12241,N_9035,N_10911);
nor U12242 (N_12242,N_11109,N_11807);
nor U12243 (N_12243,N_10759,N_10177);
nor U12244 (N_12244,N_9705,N_10079);
and U12245 (N_12245,N_9077,N_11735);
and U12246 (N_12246,N_9520,N_10470);
nand U12247 (N_12247,N_9913,N_11793);
and U12248 (N_12248,N_11219,N_10441);
and U12249 (N_12249,N_11587,N_11528);
nand U12250 (N_12250,N_9846,N_9324);
and U12251 (N_12251,N_11149,N_9972);
nand U12252 (N_12252,N_9272,N_9852);
or U12253 (N_12253,N_9888,N_10287);
and U12254 (N_12254,N_11558,N_9092);
and U12255 (N_12255,N_9394,N_11884);
nor U12256 (N_12256,N_10357,N_10708);
nand U12257 (N_12257,N_9532,N_11168);
or U12258 (N_12258,N_9975,N_11037);
nand U12259 (N_12259,N_10848,N_11345);
nand U12260 (N_12260,N_11961,N_9789);
nand U12261 (N_12261,N_11796,N_9743);
and U12262 (N_12262,N_11820,N_11064);
xnor U12263 (N_12263,N_11535,N_11336);
and U12264 (N_12264,N_9064,N_10944);
or U12265 (N_12265,N_9687,N_10547);
nand U12266 (N_12266,N_10752,N_11887);
nand U12267 (N_12267,N_9159,N_10380);
or U12268 (N_12268,N_9009,N_10799);
nor U12269 (N_12269,N_11965,N_11260);
or U12270 (N_12270,N_11120,N_10093);
and U12271 (N_12271,N_9323,N_11111);
nand U12272 (N_12272,N_9044,N_9566);
nor U12273 (N_12273,N_10286,N_10732);
nand U12274 (N_12274,N_11529,N_10274);
nand U12275 (N_12275,N_9078,N_11862);
nor U12276 (N_12276,N_10074,N_10068);
or U12277 (N_12277,N_11165,N_9823);
or U12278 (N_12278,N_9475,N_9151);
or U12279 (N_12279,N_10690,N_9609);
nand U12280 (N_12280,N_10543,N_9528);
or U12281 (N_12281,N_11480,N_9700);
xnor U12282 (N_12282,N_10382,N_9900);
or U12283 (N_12283,N_9526,N_10789);
or U12284 (N_12284,N_9149,N_11190);
nand U12285 (N_12285,N_11040,N_9965);
nor U12286 (N_12286,N_11188,N_11125);
xor U12287 (N_12287,N_9804,N_10513);
and U12288 (N_12288,N_11034,N_11337);
xor U12289 (N_12289,N_9329,N_9864);
and U12290 (N_12290,N_9641,N_11589);
nand U12291 (N_12291,N_9217,N_11289);
nand U12292 (N_12292,N_11466,N_10230);
xnor U12293 (N_12293,N_9423,N_9749);
and U12294 (N_12294,N_10106,N_9527);
nand U12295 (N_12295,N_10755,N_10345);
xor U12296 (N_12296,N_11002,N_9390);
nand U12297 (N_12297,N_10280,N_11088);
nor U12298 (N_12298,N_9835,N_9982);
nand U12299 (N_12299,N_10073,N_10375);
nand U12300 (N_12300,N_10312,N_10734);
and U12301 (N_12301,N_10006,N_10242);
or U12302 (N_12302,N_10908,N_11317);
nand U12303 (N_12303,N_10821,N_9328);
nand U12304 (N_12304,N_11038,N_10019);
or U12305 (N_12305,N_10934,N_11353);
nor U12306 (N_12306,N_9322,N_9393);
and U12307 (N_12307,N_9472,N_10991);
nor U12308 (N_12308,N_10396,N_10228);
nor U12309 (N_12309,N_10237,N_11516);
nand U12310 (N_12310,N_10090,N_11135);
nor U12311 (N_12311,N_10818,N_10126);
and U12312 (N_12312,N_9276,N_11143);
or U12313 (N_12313,N_11923,N_10253);
and U12314 (N_12314,N_9284,N_9312);
nand U12315 (N_12315,N_11436,N_9538);
or U12316 (N_12316,N_10564,N_11648);
and U12317 (N_12317,N_9420,N_10931);
and U12318 (N_12318,N_10862,N_11314);
nand U12319 (N_12319,N_10801,N_10331);
nand U12320 (N_12320,N_9046,N_11364);
nor U12321 (N_12321,N_9303,N_9946);
nand U12322 (N_12322,N_9264,N_9150);
or U12323 (N_12323,N_9949,N_11896);
nor U12324 (N_12324,N_9337,N_11006);
xnor U12325 (N_12325,N_10439,N_10524);
nand U12326 (N_12326,N_9361,N_9878);
or U12327 (N_12327,N_9503,N_11785);
and U12328 (N_12328,N_10423,N_9386);
nor U12329 (N_12329,N_11518,N_10881);
and U12330 (N_12330,N_11027,N_10726);
and U12331 (N_12331,N_9163,N_9179);
and U12332 (N_12332,N_10959,N_9350);
or U12333 (N_12333,N_9781,N_11477);
or U12334 (N_12334,N_11354,N_10276);
nor U12335 (N_12335,N_10042,N_9465);
nor U12336 (N_12336,N_10088,N_10624);
nor U12337 (N_12337,N_11580,N_11183);
nor U12338 (N_12338,N_9529,N_9748);
nand U12339 (N_12339,N_11430,N_9165);
nor U12340 (N_12340,N_10463,N_9240);
nor U12341 (N_12341,N_10865,N_9100);
and U12342 (N_12342,N_10688,N_9585);
and U12343 (N_12343,N_11881,N_10027);
nand U12344 (N_12344,N_11903,N_11450);
or U12345 (N_12345,N_11526,N_11075);
or U12346 (N_12346,N_11327,N_11373);
and U12347 (N_12347,N_9780,N_11369);
nand U12348 (N_12348,N_10156,N_10401);
nand U12349 (N_12349,N_10383,N_11794);
or U12350 (N_12350,N_10782,N_9176);
and U12351 (N_12351,N_10561,N_10078);
or U12352 (N_12352,N_11024,N_11719);
nand U12353 (N_12353,N_10409,N_9192);
and U12354 (N_12354,N_9850,N_10545);
or U12355 (N_12355,N_11764,N_11644);
nor U12356 (N_12356,N_10971,N_11401);
nand U12357 (N_12357,N_9389,N_9691);
nand U12358 (N_12358,N_10515,N_10735);
nand U12359 (N_12359,N_9973,N_11095);
and U12360 (N_12360,N_11323,N_9647);
or U12361 (N_12361,N_11920,N_11272);
nand U12362 (N_12362,N_11028,N_11534);
nor U12363 (N_12363,N_11740,N_10936);
nor U12364 (N_12364,N_10684,N_9427);
nor U12365 (N_12365,N_10339,N_11949);
and U12366 (N_12366,N_10445,N_11137);
or U12367 (N_12367,N_10730,N_10359);
or U12368 (N_12368,N_9023,N_9054);
nand U12369 (N_12369,N_11370,N_10102);
or U12370 (N_12370,N_10471,N_10135);
or U12371 (N_12371,N_11051,N_10830);
nor U12372 (N_12372,N_10566,N_11399);
nor U12373 (N_12373,N_9000,N_10424);
xor U12374 (N_12374,N_9249,N_11475);
nand U12375 (N_12375,N_11671,N_11590);
nand U12376 (N_12376,N_11928,N_11407);
nand U12377 (N_12377,N_10760,N_9366);
nor U12378 (N_12378,N_9195,N_11727);
nor U12379 (N_12379,N_9408,N_10698);
nor U12380 (N_12380,N_10214,N_10450);
xor U12381 (N_12381,N_11468,N_11464);
nor U12382 (N_12382,N_10787,N_9599);
and U12383 (N_12383,N_10028,N_11821);
or U12384 (N_12384,N_11916,N_9690);
or U12385 (N_12385,N_10576,N_11503);
nand U12386 (N_12386,N_10358,N_9617);
nor U12387 (N_12387,N_11725,N_11909);
and U12388 (N_12388,N_11842,N_11974);
or U12389 (N_12389,N_10836,N_9216);
nor U12390 (N_12390,N_9981,N_11956);
nand U12391 (N_12391,N_11667,N_10587);
nand U12392 (N_12392,N_11932,N_10071);
or U12393 (N_12393,N_11152,N_11736);
nor U12394 (N_12394,N_11576,N_11878);
nor U12395 (N_12395,N_9831,N_10872);
nand U12396 (N_12396,N_11046,N_10970);
nand U12397 (N_12397,N_11588,N_11016);
nor U12398 (N_12398,N_9153,N_10155);
nand U12399 (N_12399,N_10894,N_10187);
and U12400 (N_12400,N_10695,N_11929);
nor U12401 (N_12401,N_11843,N_10111);
nand U12402 (N_12402,N_11815,N_11733);
nand U12403 (N_12403,N_9140,N_11601);
nor U12404 (N_12404,N_10993,N_11192);
and U12405 (N_12405,N_11687,N_10542);
nand U12406 (N_12406,N_9758,N_9006);
nor U12407 (N_12407,N_11233,N_11497);
or U12408 (N_12408,N_11282,N_9235);
nand U12409 (N_12409,N_10713,N_10194);
nor U12410 (N_12410,N_11700,N_9883);
or U12411 (N_12411,N_11457,N_11101);
nor U12412 (N_12412,N_9719,N_11365);
nand U12413 (N_12413,N_10171,N_10846);
nand U12414 (N_12414,N_10585,N_9586);
or U12415 (N_12415,N_9908,N_11514);
nand U12416 (N_12416,N_11344,N_11888);
and U12417 (N_12417,N_11525,N_10412);
and U12418 (N_12418,N_9744,N_9139);
nor U12419 (N_12419,N_11126,N_10577);
or U12420 (N_12420,N_11238,N_10281);
or U12421 (N_12421,N_10966,N_11092);
and U12422 (N_12422,N_11052,N_11921);
and U12423 (N_12423,N_11962,N_11902);
or U12424 (N_12424,N_11726,N_11661);
or U12425 (N_12425,N_9246,N_9535);
nor U12426 (N_12426,N_9238,N_11950);
nand U12427 (N_12427,N_11833,N_11768);
nor U12428 (N_12428,N_10924,N_9796);
nor U12429 (N_12429,N_10694,N_10912);
nand U12430 (N_12430,N_11629,N_11632);
and U12431 (N_12431,N_11886,N_11673);
and U12432 (N_12432,N_9259,N_9255);
nor U12433 (N_12433,N_11872,N_11483);
nor U12434 (N_12434,N_9651,N_9544);
nand U12435 (N_12435,N_11704,N_9654);
nand U12436 (N_12436,N_9996,N_10617);
nand U12437 (N_12437,N_11507,N_9907);
nor U12438 (N_12438,N_10352,N_9819);
nand U12439 (N_12439,N_10707,N_10092);
and U12440 (N_12440,N_11194,N_10662);
or U12441 (N_12441,N_11571,N_9325);
nand U12442 (N_12442,N_9226,N_9262);
or U12443 (N_12443,N_9964,N_11355);
and U12444 (N_12444,N_10659,N_10211);
and U12445 (N_12445,N_9019,N_9849);
and U12446 (N_12446,N_9791,N_11556);
nand U12447 (N_12447,N_10845,N_9664);
nor U12448 (N_12448,N_9998,N_9997);
or U12449 (N_12449,N_11906,N_11844);
nand U12450 (N_12450,N_10116,N_11118);
and U12451 (N_12451,N_11019,N_9740);
nor U12452 (N_12452,N_11221,N_11692);
nor U12453 (N_12453,N_9416,N_9952);
or U12454 (N_12454,N_9113,N_9771);
nand U12455 (N_12455,N_9786,N_11658);
nor U12456 (N_12456,N_11247,N_9228);
xor U12457 (N_12457,N_9518,N_11003);
or U12458 (N_12458,N_9937,N_11096);
nand U12459 (N_12459,N_10941,N_9574);
and U12460 (N_12460,N_9459,N_11536);
nand U12461 (N_12461,N_9765,N_10080);
nor U12462 (N_12462,N_11852,N_9882);
and U12463 (N_12463,N_11493,N_9070);
nand U12464 (N_12464,N_11972,N_11760);
nand U12465 (N_12465,N_10645,N_11128);
nor U12466 (N_12466,N_10880,N_9237);
nand U12467 (N_12467,N_11698,N_10774);
or U12468 (N_12468,N_11012,N_11677);
nand U12469 (N_12469,N_10085,N_9628);
xor U12470 (N_12470,N_10609,N_9342);
nor U12471 (N_12471,N_10007,N_11586);
nor U12472 (N_12472,N_9652,N_10546);
nand U12473 (N_12473,N_10657,N_9332);
or U12474 (N_12474,N_10797,N_11216);
nand U12475 (N_12475,N_10850,N_9301);
or U12476 (N_12476,N_11486,N_9107);
and U12477 (N_12477,N_11777,N_10861);
and U12478 (N_12478,N_11787,N_11786);
or U12479 (N_12479,N_10773,N_9848);
nor U12480 (N_12480,N_10413,N_10781);
or U12481 (N_12481,N_10398,N_10878);
and U12482 (N_12482,N_9156,N_10696);
and U12483 (N_12483,N_10605,N_11814);
nor U12484 (N_12484,N_9735,N_10000);
and U12485 (N_12485,N_10525,N_10667);
nand U12486 (N_12486,N_9481,N_10044);
nand U12487 (N_12487,N_10905,N_9542);
nor U12488 (N_12488,N_9168,N_9801);
nor U12489 (N_12489,N_9109,N_9497);
nand U12490 (N_12490,N_11262,N_9045);
and U12491 (N_12491,N_9788,N_11446);
nand U12492 (N_12492,N_9533,N_10679);
nand U12493 (N_12493,N_10958,N_9757);
nand U12494 (N_12494,N_11159,N_10178);
or U12495 (N_12495,N_9132,N_9643);
nand U12496 (N_12496,N_9760,N_11592);
and U12497 (N_12497,N_10899,N_10984);
and U12498 (N_12498,N_10291,N_9842);
nand U12499 (N_12499,N_9658,N_11890);
and U12500 (N_12500,N_9693,N_9162);
nor U12501 (N_12501,N_10807,N_10809);
nor U12502 (N_12502,N_9969,N_9111);
or U12503 (N_12503,N_9613,N_9057);
xor U12504 (N_12504,N_9920,N_11593);
or U12505 (N_12505,N_11970,N_11148);
and U12506 (N_12506,N_9152,N_10256);
nor U12507 (N_12507,N_11617,N_10603);
nor U12508 (N_12508,N_11315,N_10179);
nand U12509 (N_12509,N_11086,N_9185);
nor U12510 (N_12510,N_11541,N_11800);
nor U12511 (N_12511,N_10227,N_10504);
nand U12512 (N_12512,N_9824,N_9901);
nor U12513 (N_12513,N_10420,N_11495);
or U12514 (N_12514,N_11530,N_11854);
or U12515 (N_12515,N_11699,N_9495);
nand U12516 (N_12516,N_10907,N_11633);
nand U12517 (N_12517,N_10721,N_10553);
nor U12518 (N_12518,N_10058,N_11967);
nor U12519 (N_12519,N_11849,N_10724);
nor U12520 (N_12520,N_10884,N_11400);
nor U12521 (N_12521,N_11741,N_10049);
and U12522 (N_12522,N_9261,N_11625);
or U12523 (N_12523,N_10091,N_10606);
nand U12524 (N_12524,N_10539,N_9305);
and U12525 (N_12525,N_10108,N_10070);
nand U12526 (N_12526,N_11860,N_11014);
xor U12527 (N_12527,N_10186,N_10468);
nand U12528 (N_12528,N_9841,N_10363);
nor U12529 (N_12529,N_10601,N_9634);
nor U12530 (N_12530,N_10740,N_10095);
nand U12531 (N_12531,N_11640,N_10960);
nor U12532 (N_12532,N_11816,N_9942);
and U12533 (N_12533,N_10520,N_11205);
nor U12534 (N_12534,N_10544,N_9677);
nand U12535 (N_12535,N_10395,N_11422);
nor U12536 (N_12536,N_11931,N_11999);
nand U12537 (N_12537,N_10197,N_9263);
and U12538 (N_12538,N_10786,N_9790);
or U12539 (N_12539,N_9860,N_11251);
and U12540 (N_12540,N_9960,N_9924);
or U12541 (N_12541,N_11822,N_9941);
nand U12542 (N_12542,N_11015,N_11650);
and U12543 (N_12543,N_9933,N_11324);
nor U12544 (N_12544,N_11752,N_9030);
and U12545 (N_12545,N_11653,N_9844);
nor U12546 (N_12546,N_9716,N_10537);
or U12547 (N_12547,N_9768,N_10185);
nand U12548 (N_12548,N_11073,N_9834);
nor U12549 (N_12549,N_9619,N_10267);
nand U12550 (N_12550,N_9173,N_10521);
xnor U12551 (N_12551,N_11829,N_9918);
nand U12552 (N_12552,N_9293,N_9659);
and U12553 (N_12553,N_11971,N_9919);
and U12554 (N_12554,N_9554,N_10192);
nor U12555 (N_12555,N_10474,N_9991);
nand U12556 (N_12556,N_9181,N_11859);
nand U12557 (N_12557,N_9722,N_11009);
and U12558 (N_12558,N_9556,N_9069);
or U12559 (N_12559,N_11537,N_10075);
nand U12560 (N_12560,N_10460,N_10084);
and U12561 (N_12561,N_11602,N_11182);
or U12562 (N_12562,N_11013,N_11304);
nor U12563 (N_12563,N_11236,N_9727);
or U12564 (N_12564,N_10540,N_10240);
and U12565 (N_12565,N_10834,N_11979);
or U12566 (N_12566,N_10810,N_9377);
xor U12567 (N_12567,N_11892,N_10703);
nand U12568 (N_12568,N_10868,N_9220);
nand U12569 (N_12569,N_9136,N_10145);
nand U12570 (N_12570,N_9346,N_9611);
nor U12571 (N_12571,N_10635,N_11883);
nand U12572 (N_12572,N_10089,N_11581);
nand U12573 (N_12573,N_9562,N_10528);
nor U12574 (N_12574,N_11065,N_9374);
or U12575 (N_12575,N_9202,N_9766);
and U12576 (N_12576,N_10313,N_11359);
or U12577 (N_12577,N_10571,N_9017);
nor U12578 (N_12578,N_10994,N_9287);
and U12579 (N_12579,N_9898,N_10462);
or U12580 (N_12580,N_9032,N_10776);
and U12581 (N_12581,N_10582,N_9347);
or U12582 (N_12582,N_10051,N_9537);
or U12583 (N_12583,N_9158,N_10866);
and U12584 (N_12584,N_11361,N_11910);
nand U12585 (N_12585,N_10325,N_10769);
nor U12586 (N_12586,N_9553,N_11377);
and U12587 (N_12587,N_11550,N_9160);
and U12588 (N_12588,N_9108,N_9310);
nor U12589 (N_12589,N_9640,N_9213);
nor U12590 (N_12590,N_10805,N_9838);
and U12591 (N_12591,N_11067,N_9457);
and U12592 (N_12592,N_11730,N_10431);
nand U12593 (N_12593,N_10580,N_10867);
and U12594 (N_12594,N_11905,N_9966);
nand U12595 (N_12595,N_11082,N_9411);
nand U12596 (N_12596,N_9012,N_10929);
nand U12597 (N_12597,N_9704,N_10661);
and U12598 (N_12598,N_9774,N_9479);
and U12599 (N_12599,N_9198,N_11519);
and U12600 (N_12600,N_11708,N_11214);
and U12601 (N_12601,N_10751,N_11107);
nor U12602 (N_12602,N_10775,N_10604);
nor U12603 (N_12603,N_10989,N_9612);
xnor U12604 (N_12604,N_9365,N_10764);
or U12605 (N_12605,N_11734,N_9206);
and U12606 (N_12606,N_9015,N_11218);
or U12607 (N_12607,N_9752,N_10614);
or U12608 (N_12608,N_9502,N_10464);
or U12609 (N_12609,N_11510,N_9616);
nand U12610 (N_12610,N_11063,N_10906);
nand U12611 (N_12611,N_10640,N_10608);
or U12612 (N_12612,N_10935,N_11731);
or U12613 (N_12613,N_9137,N_9828);
nor U12614 (N_12614,N_11758,N_10519);
nand U12615 (N_12615,N_11074,N_9661);
nor U12616 (N_12616,N_11339,N_11036);
or U12617 (N_12617,N_10890,N_10990);
or U12618 (N_12618,N_10146,N_11812);
nand U12619 (N_12619,N_9935,N_11712);
or U12620 (N_12620,N_9747,N_9463);
nand U12621 (N_12621,N_10344,N_11682);
or U12622 (N_12622,N_10992,N_10366);
nand U12623 (N_12623,N_9025,N_11117);
nor U12624 (N_12624,N_10921,N_11122);
nor U12625 (N_12625,N_10165,N_9627);
nor U12626 (N_12626,N_11607,N_11566);
nand U12627 (N_12627,N_10843,N_10849);
nor U12628 (N_12628,N_11319,N_10663);
nor U12629 (N_12629,N_11039,N_11898);
or U12630 (N_12630,N_11772,N_10920);
nand U12631 (N_12631,N_9147,N_9453);
or U12632 (N_12632,N_11235,N_11948);
or U12633 (N_12633,N_10693,N_11986);
or U12634 (N_12634,N_9927,N_11781);
nand U12635 (N_12635,N_9349,N_11098);
or U12636 (N_12636,N_11406,N_9431);
nor U12637 (N_12637,N_10077,N_10565);
or U12638 (N_12638,N_9892,N_10871);
or U12639 (N_12639,N_10949,N_9222);
nor U12640 (N_12640,N_9968,N_10916);
xnor U12641 (N_12641,N_11603,N_9779);
nand U12642 (N_12642,N_11138,N_9055);
nand U12643 (N_12643,N_10879,N_9369);
nand U12644 (N_12644,N_11416,N_9273);
and U12645 (N_12645,N_11478,N_9709);
or U12646 (N_12646,N_11133,N_11506);
or U12647 (N_12647,N_9351,N_11211);
or U12648 (N_12648,N_9827,N_9588);
and U12649 (N_12649,N_9373,N_9632);
nand U12650 (N_12650,N_11440,N_9872);
nor U12651 (N_12651,N_9437,N_9432);
and U12652 (N_12652,N_10675,N_10656);
nor U12653 (N_12653,N_9130,N_11936);
and U12654 (N_12654,N_9091,N_10736);
nor U12655 (N_12655,N_11867,N_10112);
and U12656 (N_12656,N_9088,N_11567);
or U12657 (N_12657,N_10324,N_10969);
nor U12658 (N_12658,N_11934,N_10434);
and U12659 (N_12659,N_10628,N_9507);
or U12660 (N_12660,N_9540,N_9655);
and U12661 (N_12661,N_10246,N_11288);
and U12662 (N_12662,N_11505,N_11724);
or U12663 (N_12663,N_11811,N_11499);
or U12664 (N_12664,N_11420,N_10341);
nand U12665 (N_12665,N_10266,N_10589);
or U12666 (N_12666,N_11452,N_11522);
nor U12667 (N_12667,N_11212,N_11810);
and U12668 (N_12668,N_10611,N_9405);
and U12669 (N_12669,N_11329,N_9858);
or U12670 (N_12670,N_11797,N_9296);
nor U12671 (N_12671,N_10210,N_10549);
and U12672 (N_12672,N_9388,N_11121);
nor U12673 (N_12673,N_9254,N_11381);
nor U12674 (N_12674,N_11638,N_11007);
nor U12675 (N_12675,N_11102,N_9289);
and U12676 (N_12676,N_11066,N_9494);
or U12677 (N_12677,N_10249,N_10290);
nand U12678 (N_12678,N_9971,N_9642);
nor U12679 (N_12679,N_9983,N_11309);
and U12680 (N_12680,N_10493,N_9618);
or U12681 (N_12681,N_11252,N_11737);
xor U12682 (N_12682,N_10637,N_9489);
or U12683 (N_12683,N_10927,N_10699);
nor U12684 (N_12684,N_10784,N_10298);
and U12685 (N_12685,N_11723,N_10538);
xor U12686 (N_12686,N_11424,N_9714);
and U12687 (N_12687,N_10655,N_10131);
nor U12688 (N_12688,N_11011,N_11579);
and U12689 (N_12689,N_11431,N_9001);
nor U12690 (N_12690,N_10683,N_11944);
or U12691 (N_12691,N_10766,N_9555);
or U12692 (N_12692,N_10342,N_11552);
nand U12693 (N_12693,N_10207,N_11105);
and U12694 (N_12694,N_10160,N_10167);
or U12695 (N_12695,N_10643,N_10649);
nor U12696 (N_12696,N_9204,N_9825);
and U12697 (N_12697,N_11847,N_10057);
nor U12698 (N_12698,N_9557,N_10586);
or U12699 (N_12699,N_9485,N_10842);
nand U12700 (N_12700,N_11472,N_9104);
or U12701 (N_12701,N_11237,N_11933);
and U12702 (N_12702,N_11030,N_10238);
nand U12703 (N_12703,N_10500,N_11875);
or U12704 (N_12704,N_9957,N_10134);
or U12705 (N_12705,N_10013,N_10098);
nand U12706 (N_12706,N_10285,N_11079);
and U12707 (N_12707,N_11562,N_10340);
nor U12708 (N_12708,N_11914,N_11953);
or U12709 (N_12709,N_9496,N_10166);
nor U12710 (N_12710,N_9491,N_9398);
and U12711 (N_12711,N_11453,N_11597);
nand U12712 (N_12712,N_10658,N_10599);
or U12713 (N_12713,N_10530,N_9899);
and U12714 (N_12714,N_10945,N_9352);
or U12715 (N_12715,N_10534,N_11343);
nor U12716 (N_12716,N_10272,N_11978);
nand U12717 (N_12717,N_9995,N_9189);
nand U12718 (N_12718,N_9778,N_9606);
nor U12719 (N_12719,N_10444,N_9720);
nand U12720 (N_12720,N_10385,N_10750);
nor U12721 (N_12721,N_10532,N_11396);
and U12722 (N_12722,N_10316,N_9863);
and U12723 (N_12723,N_11071,N_11145);
or U12724 (N_12724,N_10743,N_9005);
xnor U12725 (N_12725,N_9548,N_10491);
nand U12726 (N_12726,N_10045,N_9215);
nor U12727 (N_12727,N_9762,N_11750);
and U12728 (N_12728,N_9840,N_10982);
or U12729 (N_12729,N_11720,N_11467);
xnor U12730 (N_12730,N_11090,N_11267);
nor U12731 (N_12731,N_11390,N_11153);
nor U12732 (N_12732,N_11674,N_9821);
and U12733 (N_12733,N_9306,N_11209);
nor U12734 (N_12734,N_11714,N_9144);
nor U12735 (N_12735,N_9331,N_9884);
or U12736 (N_12736,N_11851,N_10478);
or U12737 (N_12737,N_9701,N_11091);
nand U12738 (N_12738,N_11598,N_9887);
nor U12739 (N_12739,N_10475,N_11386);
nand U12740 (N_12740,N_10650,N_10680);
and U12741 (N_12741,N_9134,N_10456);
nor U12742 (N_12742,N_10953,N_11551);
and U12743 (N_12743,N_9200,N_9429);
or U12744 (N_12744,N_9208,N_11688);
nor U12745 (N_12745,N_10021,N_11041);
or U12746 (N_12746,N_10368,N_9311);
nor U12747 (N_12747,N_10144,N_11418);
or U12748 (N_12748,N_11479,N_11819);
and U12749 (N_12749,N_9083,N_9967);
nand U12750 (N_12750,N_9685,N_9717);
or U12751 (N_12751,N_9552,N_9068);
and U12752 (N_12752,N_9589,N_9441);
and U12753 (N_12753,N_9076,N_11470);
and U12754 (N_12754,N_11635,N_9510);
and U12755 (N_12755,N_11290,N_9364);
and U12756 (N_12756,N_9745,N_9775);
nand U12757 (N_12757,N_10002,N_11524);
nor U12758 (N_12758,N_9381,N_10440);
nand U12759 (N_12759,N_11563,N_10646);
and U12760 (N_12760,N_9662,N_10017);
and U12761 (N_12761,N_11937,N_9197);
nor U12762 (N_12762,N_10320,N_9961);
nor U12763 (N_12763,N_10428,N_10258);
and U12764 (N_12764,N_9487,N_11162);
nor U12765 (N_12765,N_10742,N_11332);
nor U12766 (N_12766,N_10768,N_9645);
nand U12767 (N_12767,N_10942,N_9354);
or U12768 (N_12768,N_9440,N_9379);
nor U12769 (N_12769,N_11193,N_11806);
and U12770 (N_12770,N_11284,N_11281);
nor U12771 (N_12771,N_10182,N_11904);
or U12772 (N_12772,N_9101,N_9584);
nor U12773 (N_12773,N_10234,N_10296);
nor U12774 (N_12774,N_11766,N_11831);
nor U12775 (N_12775,N_10148,N_10859);
nor U12776 (N_12776,N_9605,N_10804);
or U12777 (N_12777,N_10213,N_9187);
nor U12778 (N_12778,N_9253,N_10512);
nand U12779 (N_12779,N_9252,N_10269);
and U12780 (N_12780,N_9292,N_11023);
nand U12781 (N_12781,N_10482,N_9490);
nor U12782 (N_12782,N_11619,N_9582);
or U12783 (N_12783,N_11129,N_9321);
or U12784 (N_12784,N_11826,N_9635);
nand U12785 (N_12785,N_11945,N_11360);
nand U12786 (N_12786,N_10008,N_9928);
or U12787 (N_12787,N_11348,N_10030);
or U12788 (N_12788,N_11335,N_9396);
nor U12789 (N_12789,N_11201,N_11721);
nand U12790 (N_12790,N_9099,N_11665);
nand U12791 (N_12791,N_10638,N_10882);
and U12792 (N_12792,N_9577,N_9521);
nand U12793 (N_12793,N_10901,N_9014);
or U12794 (N_12794,N_9166,N_9298);
nand U12795 (N_12795,N_10304,N_11476);
nand U12796 (N_12796,N_11231,N_11081);
nor U12797 (N_12797,N_10196,N_11802);
xnor U12798 (N_12798,N_9843,N_9895);
nand U12799 (N_12799,N_11871,N_10432);
and U12800 (N_12800,N_11411,N_9128);
or U12801 (N_12801,N_9764,N_10188);
nor U12802 (N_12802,N_9318,N_11858);
and U12803 (N_12803,N_10056,N_10480);
and U12804 (N_12804,N_9120,N_10327);
or U12805 (N_12805,N_10622,N_11520);
nor U12806 (N_12806,N_11855,N_9523);
nor U12807 (N_12807,N_10794,N_11924);
nand U12808 (N_12808,N_9723,N_10097);
nand U12809 (N_12809,N_11106,N_10448);
and U12810 (N_12810,N_10965,N_9814);
xnor U12811 (N_12811,N_9067,N_10372);
nand U12812 (N_12812,N_9279,N_11968);
or U12813 (N_12813,N_10279,N_11613);
nor U12814 (N_12814,N_9122,N_9079);
and U12815 (N_12815,N_11542,N_10164);
and U12816 (N_12816,N_11697,N_9141);
xor U12817 (N_12817,N_10983,N_9986);
and U12818 (N_12818,N_9680,N_11055);
and U12819 (N_12819,N_10139,N_10812);
nand U12820 (N_12820,N_11367,N_9177);
and U12821 (N_12821,N_10738,N_10288);
and U12822 (N_12822,N_9283,N_10371);
nor U12823 (N_12823,N_10416,N_11561);
nand U12824 (N_12824,N_10506,N_10217);
and U12825 (N_12825,N_10647,N_11248);
nand U12826 (N_12826,N_9622,N_11286);
or U12827 (N_12827,N_10852,N_10114);
or U12828 (N_12828,N_11747,N_11443);
and U12829 (N_12829,N_9266,N_11239);
nor U12830 (N_12830,N_10831,N_9224);
nor U12831 (N_12831,N_9644,N_10888);
nor U12832 (N_12832,N_9155,N_10972);
or U12833 (N_12833,N_10035,N_10446);
or U12834 (N_12834,N_9666,N_11841);
and U12835 (N_12835,N_11623,N_9493);
nor U12836 (N_12836,N_11384,N_10406);
and U12837 (N_12837,N_9335,N_10985);
nand U12838 (N_12838,N_11825,N_11559);
xnor U12839 (N_12839,N_10050,N_9439);
nand U12840 (N_12840,N_9380,N_9909);
and U12841 (N_12841,N_11685,N_10319);
and U12842 (N_12842,N_9742,N_9868);
nand U12843 (N_12843,N_9295,N_10583);
nand U12844 (N_12844,N_10009,N_10061);
nor U12845 (N_12845,N_11328,N_9890);
nand U12846 (N_12846,N_11917,N_10665);
and U12847 (N_12847,N_9334,N_9561);
nor U12848 (N_12848,N_9737,N_10592);
nor U12849 (N_12849,N_10261,N_10737);
or U12850 (N_12850,N_9767,N_10826);
nor U12851 (N_12851,N_9678,N_10548);
nand U12852 (N_12852,N_10152,N_9219);
nand U12853 (N_12853,N_9569,N_9881);
and U12854 (N_12854,N_10632,N_10447);
or U12855 (N_12855,N_9383,N_10676);
and U12856 (N_12856,N_11803,N_10259);
and U12857 (N_12857,N_11743,N_10430);
or U12858 (N_12858,N_10026,N_9022);
or U12859 (N_12859,N_11334,N_9733);
and U12860 (N_12860,N_11616,N_10555);
nor U12861 (N_12861,N_9943,N_11062);
nand U12862 (N_12862,N_11204,N_9281);
and U12863 (N_12863,N_9473,N_9877);
or U12864 (N_12864,N_11717,N_10531);
nand U12865 (N_12865,N_9567,N_10922);
and U12866 (N_12866,N_11191,N_9455);
or U12867 (N_12867,N_11788,N_11402);
or U12868 (N_12868,N_9633,N_10817);
nor U12869 (N_12869,N_9649,N_10457);
or U12870 (N_12870,N_9340,N_10303);
or U12871 (N_12871,N_10686,N_11350);
nor U12872 (N_12872,N_10674,N_9699);
and U12873 (N_12873,N_10788,N_11911);
or U12874 (N_12874,N_10354,N_11523);
and U12875 (N_12875,N_11678,N_10399);
nor U12876 (N_12876,N_9832,N_9812);
nor U12877 (N_12877,N_9232,N_11547);
nor U12878 (N_12878,N_9387,N_11089);
xnor U12879 (N_12879,N_10584,N_11278);
or U12880 (N_12880,N_9319,N_11371);
and U12881 (N_12881,N_9904,N_9876);
and U12882 (N_12882,N_11186,N_9484);
nor U12883 (N_12883,N_11022,N_9950);
or U12884 (N_12884,N_11068,N_11779);
or U12885 (N_12885,N_10811,N_10783);
nor U12886 (N_12886,N_11836,N_9992);
nand U12887 (N_12887,N_9458,N_10337);
or U12888 (N_12888,N_10064,N_9773);
or U12889 (N_12889,N_11076,N_11894);
and U12890 (N_12890,N_9148,N_9925);
nand U12891 (N_12891,N_9857,N_10681);
or U12892 (N_12892,N_11362,N_11448);
nand U12893 (N_12893,N_9072,N_11515);
nor U12894 (N_12894,N_10793,N_9715);
nor U12895 (N_12895,N_10630,N_10476);
nor U12896 (N_12896,N_10716,N_11458);
or U12897 (N_12897,N_10719,N_9534);
nor U12898 (N_12898,N_9668,N_10086);
nand U12899 (N_12899,N_9444,N_10118);
or U12900 (N_12900,N_10317,N_10814);
or U12901 (N_12901,N_9551,N_11378);
nor U12902 (N_12902,N_9707,N_9770);
and U12903 (N_12903,N_11754,N_10517);
nor U12904 (N_12904,N_10806,N_10031);
nand U12905 (N_12905,N_9570,N_11918);
and U12906 (N_12906,N_10168,N_9974);
nand U12907 (N_12907,N_10130,N_10015);
or U12908 (N_12908,N_10791,N_10277);
nor U12909 (N_12909,N_10231,N_9034);
nor U12910 (N_12910,N_11397,N_9115);
or U12911 (N_12911,N_10151,N_9759);
and U12912 (N_12912,N_11097,N_9280);
nand U12913 (N_12913,N_10792,N_10270);
or U12914 (N_12914,N_9060,N_10923);
nor U12915 (N_12915,N_10193,N_11217);
nor U12916 (N_12916,N_10404,N_11417);
nor U12917 (N_12917,N_11706,N_9531);
or U12918 (N_12918,N_9880,N_11268);
nor U12919 (N_12919,N_9071,N_11958);
and U12920 (N_12920,N_11094,N_10978);
and U12921 (N_12921,N_9314,N_9209);
nand U12922 (N_12922,N_9330,N_10018);
nor U12923 (N_12923,N_11412,N_9754);
or U12924 (N_12924,N_11801,N_10728);
or U12925 (N_12925,N_11919,N_9718);
nor U12926 (N_12926,N_10712,N_11299);
nand U12927 (N_12927,N_11375,N_11709);
nor U12928 (N_12928,N_9977,N_9558);
or U12929 (N_12929,N_10762,N_9483);
or U12930 (N_12930,N_10727,N_10568);
nand U12931 (N_12931,N_9397,N_11988);
nand U12932 (N_12932,N_10314,N_9327);
nand U12933 (N_12933,N_9698,N_9833);
nand U12934 (N_12934,N_11870,N_10741);
nand U12935 (N_12935,N_11771,N_9268);
or U12936 (N_12936,N_10494,N_11110);
nor U12937 (N_12937,N_9178,N_9434);
or U12938 (N_12938,N_11657,N_9836);
nor U12939 (N_12939,N_9811,N_10418);
nand U12940 (N_12940,N_10278,N_11103);
nor U12941 (N_12941,N_10349,N_10772);
nand U12942 (N_12942,N_9522,N_11652);
nor U12943 (N_12943,N_9563,N_11845);
nor U12944 (N_12944,N_9167,N_9265);
nor U12945 (N_12945,N_10939,N_9509);
or U12946 (N_12946,N_11490,N_9516);
nor U12947 (N_12947,N_11047,N_10839);
or U12948 (N_12948,N_9241,N_10858);
nor U12949 (N_12949,N_10025,N_10765);
and U12950 (N_12950,N_10529,N_11352);
and U12951 (N_12951,N_10189,N_10745);
nand U12952 (N_12952,N_11144,N_10054);
nor U12953 (N_12953,N_9018,N_10602);
nand U12954 (N_12954,N_11169,N_9871);
nor U12955 (N_12955,N_10486,N_9371);
nor U12956 (N_12956,N_11342,N_11322);
or U12957 (N_12957,N_10161,N_9359);
nand U12958 (N_12958,N_11533,N_11882);
or U12959 (N_12959,N_11223,N_10289);
nor U12960 (N_12960,N_10575,N_9183);
nand U12961 (N_12961,N_10533,N_11271);
nand U12962 (N_12962,N_10642,N_9184);
and U12963 (N_12963,N_10722,N_9450);
nor U12964 (N_12964,N_9199,N_9500);
xor U12965 (N_12965,N_10963,N_10353);
nand U12966 (N_12966,N_11770,N_9039);
xnor U12967 (N_12967,N_9639,N_10226);
and U12968 (N_12968,N_9082,N_9539);
and U12969 (N_12969,N_11025,N_10860);
nor U12970 (N_12970,N_10913,N_11070);
nor U12971 (N_12971,N_10536,N_11261);
nand U12972 (N_12972,N_10829,N_10254);
and U12973 (N_12973,N_10046,N_10332);
nor U12974 (N_12974,N_9447,N_11808);
nor U12975 (N_12975,N_10864,N_10598);
xnor U12976 (N_12976,N_10496,N_10729);
or U12977 (N_12977,N_11624,N_10110);
and U12978 (N_12978,N_11301,N_11202);
nor U12979 (N_12979,N_11912,N_9646);
nand U12980 (N_12980,N_11259,N_9894);
nand U12981 (N_12981,N_11891,N_11570);
nand U12982 (N_12982,N_10771,N_11163);
nor U12983 (N_12983,N_11382,N_10204);
or U12984 (N_12984,N_10910,N_9103);
nor U12985 (N_12985,N_10610,N_10403);
or U12986 (N_12986,N_10195,N_9936);
nor U12987 (N_12987,N_10370,N_9445);
nor U12988 (N_12988,N_9404,N_11226);
nor U12989 (N_12989,N_9267,N_11778);
and U12990 (N_12990,N_9671,N_10851);
nand U12991 (N_12991,N_9692,N_10666);
nand U12992 (N_12992,N_10149,N_10173);
or U12993 (N_12993,N_9512,N_9093);
nand U12994 (N_12994,N_10040,N_10115);
nor U12995 (N_12995,N_10389,N_11705);
nand U12996 (N_12996,N_10820,N_9320);
or U12997 (N_12997,N_10701,N_10039);
nand U12998 (N_12998,N_10550,N_10574);
and U12999 (N_12999,N_10322,N_10636);
xnor U13000 (N_13000,N_11631,N_9830);
and U13001 (N_13001,N_10451,N_10488);
or U13002 (N_13002,N_11600,N_10800);
or U13003 (N_13003,N_9037,N_10710);
and U13004 (N_13004,N_11496,N_10069);
xnor U13005 (N_13005,N_11745,N_11115);
xnor U13006 (N_13006,N_10307,N_10692);
nand U13007 (N_13007,N_11615,N_9873);
or U13008 (N_13008,N_10919,N_11753);
and U13009 (N_13009,N_11279,N_9826);
and U13010 (N_13010,N_9125,N_11158);
nor U13011 (N_13011,N_11995,N_9999);
nand U13012 (N_13012,N_11208,N_9688);
and U13013 (N_13013,N_11277,N_9729);
and U13014 (N_13014,N_11213,N_10928);
nor U13015 (N_13015,N_10467,N_10454);
or U13016 (N_13016,N_10689,N_9954);
or U13017 (N_13017,N_10052,N_11393);
nand U13018 (N_13018,N_9672,N_11877);
or U13019 (N_13019,N_9382,N_11250);
nand U13020 (N_13020,N_9591,N_10770);
and U13021 (N_13021,N_9805,N_10301);
nor U13022 (N_13022,N_10053,N_9084);
or U13023 (N_13023,N_9915,N_11963);
and U13024 (N_13024,N_9428,N_10104);
nand U13025 (N_13025,N_11482,N_9702);
nand U13026 (N_13026,N_11254,N_10933);
nand U13027 (N_13027,N_9711,N_11020);
nand U13028 (N_13028,N_11451,N_10175);
or U13029 (N_13029,N_11702,N_10169);
nand U13030 (N_13030,N_11686,N_10306);
nor U13031 (N_13031,N_10029,N_10980);
or U13032 (N_13032,N_11660,N_9188);
nand U13033 (N_13033,N_11469,N_10489);
or U13034 (N_13034,N_9806,N_10239);
or U13035 (N_13035,N_9761,N_11614);
and U13036 (N_13036,N_11018,N_9499);
and U13037 (N_13037,N_11976,N_10391);
and U13038 (N_13038,N_9236,N_11873);
and U13039 (N_13039,N_11257,N_11243);
or U13040 (N_13040,N_10898,N_9923);
or U13041 (N_13041,N_10487,N_10458);
and U13042 (N_13042,N_11318,N_9478);
nor U13043 (N_13043,N_9603,N_9002);
nor U13044 (N_13044,N_11161,N_9911);
nand U13045 (N_13045,N_11553,N_11465);
or U13046 (N_13046,N_11864,N_11232);
or U13047 (N_13047,N_11637,N_11130);
nand U13048 (N_13048,N_11404,N_11265);
or U13049 (N_13049,N_10283,N_11893);
nor U13050 (N_13050,N_10180,N_10374);
xnor U13051 (N_13051,N_9931,N_9653);
and U13052 (N_13052,N_9438,N_11606);
and U13053 (N_13053,N_10633,N_10367);
nand U13054 (N_13054,N_10150,N_9917);
nand U13055 (N_13055,N_9660,N_9875);
and U13056 (N_13056,N_11866,N_9963);
or U13057 (N_13057,N_11200,N_9315);
nor U13058 (N_13058,N_10559,N_9486);
nor U13059 (N_13059,N_10318,N_9138);
or U13060 (N_13060,N_9451,N_11651);
and U13061 (N_13061,N_9665,N_9706);
and U13062 (N_13062,N_10815,N_10365);
or U13063 (N_13063,N_10999,N_10623);
nor U13064 (N_13064,N_10181,N_11273);
or U13065 (N_13065,N_10499,N_10503);
and U13066 (N_13066,N_9307,N_9353);
and U13067 (N_13067,N_9355,N_10037);
nor U13068 (N_13068,N_9602,N_10335);
and U13069 (N_13069,N_9856,N_9889);
and U13070 (N_13070,N_11147,N_11675);
or U13071 (N_13071,N_9897,N_9543);
nand U13072 (N_13072,N_9452,N_10527);
nor U13073 (N_13073,N_11739,N_10947);
nand U13074 (N_13074,N_11010,N_11093);
nor U13075 (N_13075,N_10747,N_9598);
nand U13076 (N_13076,N_11077,N_9741);
nand U13077 (N_13077,N_10200,N_9565);
or U13078 (N_13078,N_9799,N_9938);
nand U13079 (N_13079,N_11376,N_11669);
nor U13080 (N_13080,N_11837,N_9186);
or U13081 (N_13081,N_9656,N_9623);
and U13082 (N_13082,N_11985,N_11585);
or U13083 (N_13083,N_9549,N_11256);
nand U13084 (N_13084,N_11043,N_11521);
or U13085 (N_13085,N_9932,N_11432);
nand U13086 (N_13086,N_9126,N_11441);
nand U13087 (N_13087,N_10819,N_10648);
xnor U13088 (N_13088,N_11340,N_10326);
xnor U13089 (N_13089,N_11049,N_11173);
nand U13090 (N_13090,N_9385,N_9180);
and U13091 (N_13091,N_10825,N_11127);
and U13092 (N_13092,N_11245,N_10016);
nand U13093 (N_13093,N_10886,N_10096);
nor U13094 (N_13094,N_9201,N_10651);
or U13095 (N_13095,N_10087,N_11689);
nor U13096 (N_13096,N_10996,N_9721);
and U13097 (N_13097,N_10523,N_11513);
nor U13098 (N_13098,N_10569,N_9242);
nor U13099 (N_13099,N_10038,N_11728);
and U13100 (N_13100,N_10364,N_10932);
and U13101 (N_13101,N_11366,N_9867);
nor U13102 (N_13102,N_10955,N_10767);
and U13103 (N_13103,N_9797,N_11608);
nand U13104 (N_13104,N_9530,N_10961);
nand U13105 (N_13105,N_10896,N_9285);
nor U13106 (N_13106,N_11947,N_9230);
and U13107 (N_13107,N_11984,N_10757);
nand U13108 (N_13108,N_10552,N_10654);
and U13109 (N_13109,N_11628,N_11473);
xnor U13110 (N_13110,N_9223,N_9914);
and U13111 (N_13111,N_11198,N_9985);
nand U13112 (N_13112,N_11946,N_9614);
and U13113 (N_13113,N_10964,N_11940);
and U13114 (N_13114,N_9517,N_11164);
nand U13115 (N_13115,N_11666,N_11696);
or U13116 (N_13116,N_9417,N_10895);
or U13117 (N_13117,N_10060,N_9074);
nand U13118 (N_13118,N_9085,N_9257);
or U13119 (N_13119,N_10591,N_11885);
and U13120 (N_13120,N_11792,N_10101);
and U13121 (N_13121,N_9294,N_10172);
nor U13122 (N_13122,N_10671,N_11939);
or U13123 (N_13123,N_9626,N_10107);
nand U13124 (N_13124,N_9689,N_9042);
or U13125 (N_13125,N_9193,N_9135);
and U13126 (N_13126,N_9793,N_10252);
or U13127 (N_13127,N_11307,N_9592);
nor U13128 (N_13128,N_9231,N_11626);
nand U13129 (N_13129,N_11234,N_11449);
or U13130 (N_13130,N_10218,N_11294);
nand U13131 (N_13131,N_11838,N_10629);
nand U13132 (N_13132,N_9090,N_11196);
and U13133 (N_13133,N_9866,N_9048);
or U13134 (N_13134,N_9839,N_10421);
nand U13135 (N_13135,N_11649,N_9027);
nor U13136 (N_13136,N_10020,N_11517);
and U13137 (N_13137,N_10891,N_10607);
nor U13138 (N_13138,N_11713,N_10954);
or U13139 (N_13139,N_10986,N_10472);
or U13140 (N_13140,N_10033,N_10918);
nor U13141 (N_13141,N_10616,N_10223);
xnor U13142 (N_13142,N_9482,N_11982);
and U13143 (N_13143,N_11395,N_9271);
or U13144 (N_13144,N_9970,N_9579);
nor U13145 (N_13145,N_10003,N_9906);
and U13146 (N_13146,N_11099,N_10067);
nor U13147 (N_13147,N_11242,N_11058);
or U13148 (N_13148,N_11761,N_10297);
nand U13149 (N_13149,N_9413,N_11255);
and U13150 (N_13150,N_11426,N_10687);
and U13151 (N_13151,N_10930,N_10390);
nor U13152 (N_13152,N_9468,N_11385);
and U13153 (N_13153,N_9505,N_11455);
and U13154 (N_13154,N_11759,N_10987);
nand U13155 (N_13155,N_11817,N_11504);
and U13156 (N_13156,N_9008,N_11680);
or U13157 (N_13157,N_9154,N_9820);
and U13158 (N_13158,N_11582,N_10023);
nand U13159 (N_13159,N_11952,N_10979);
and U13160 (N_13160,N_9862,N_9258);
nor U13161 (N_13161,N_11959,N_9815);
or U13162 (N_13162,N_9951,N_9696);
nor U13163 (N_13163,N_11442,N_10394);
or U13164 (N_13164,N_11437,N_11341);
or U13165 (N_13165,N_11757,N_10438);
nor U13166 (N_13166,N_10024,N_11374);
nand U13167 (N_13167,N_9559,N_10273);
or U13168 (N_13168,N_11546,N_10948);
or U13169 (N_13169,N_11429,N_9597);
or U13170 (N_13170,N_10232,N_11574);
nand U13171 (N_13171,N_11502,N_10600);
and U13172 (N_13172,N_9400,N_10305);
nor U13173 (N_13173,N_10664,N_10778);
nand U13174 (N_13174,N_9299,N_9905);
nor U13175 (N_13175,N_9419,N_11749);
and U13176 (N_13176,N_11150,N_11805);
nand U13177 (N_13177,N_11356,N_9247);
nor U13178 (N_13178,N_10012,N_11498);
nand U13179 (N_13179,N_11061,N_10411);
nand U13180 (N_13180,N_9052,N_9498);
or U13181 (N_13181,N_11645,N_9038);
nand U13182 (N_13182,N_9684,N_9360);
or U13183 (N_13183,N_11032,N_9086);
and U13184 (N_13184,N_10749,N_10706);
or U13185 (N_13185,N_9578,N_11230);
or U13186 (N_13186,N_10163,N_9989);
or U13187 (N_13187,N_10477,N_9378);
nor U13188 (N_13188,N_9409,N_11642);
nor U13189 (N_13189,N_11664,N_10835);
or U13190 (N_13190,N_9403,N_10974);
nand U13191 (N_13191,N_11383,N_9637);
nand U13192 (N_13192,N_9886,N_10619);
nand U13193 (N_13193,N_10720,N_9865);
nand U13194 (N_13194,N_10443,N_11461);
and U13195 (N_13195,N_11670,N_10376);
nand U13196 (N_13196,N_9513,N_10857);
or U13197 (N_13197,N_11981,N_11296);
nand U13198 (N_13198,N_10346,N_10461);
and U13199 (N_13199,N_11610,N_10036);
and U13200 (N_13200,N_9474,N_9763);
and U13201 (N_13201,N_11258,N_9638);
and U13202 (N_13202,N_9399,N_11303);
nor U13203 (N_13203,N_10063,N_9065);
or U13204 (N_13204,N_10120,N_11951);
or U13205 (N_13205,N_9124,N_10334);
or U13206 (N_13206,N_10041,N_11722);
nor U13207 (N_13207,N_9095,N_10348);
nand U13208 (N_13208,N_9024,N_9959);
nand U13209 (N_13209,N_10780,N_10535);
nand U13210 (N_13210,N_10005,N_10388);
or U13211 (N_13211,N_9910,N_9976);
nor U13212 (N_13212,N_9227,N_11880);
nor U13213 (N_13213,N_10422,N_10066);
nand U13214 (N_13214,N_10235,N_10951);
or U13215 (N_13215,N_10863,N_9308);
nand U13216 (N_13216,N_10299,N_10950);
nor U13217 (N_13217,N_11789,N_9401);
nand U13218 (N_13218,N_9683,N_10501);
nor U13219 (N_13219,N_10350,N_11861);
nor U13220 (N_13220,N_10373,N_9041);
and U13221 (N_13221,N_10725,N_11155);
nand U13222 (N_13222,N_9739,N_9344);
nand U13223 (N_13223,N_10433,N_11716);
or U13224 (N_13224,N_11197,N_9541);
and U13225 (N_13225,N_11114,N_9161);
or U13226 (N_13226,N_9629,N_11484);
and U13227 (N_13227,N_10203,N_11996);
and U13228 (N_13228,N_10136,N_11621);
and U13229 (N_13229,N_9182,N_9290);
nor U13230 (N_13230,N_10893,N_10157);
or U13231 (N_13231,N_9916,N_10977);
nor U13232 (N_13232,N_9595,N_10159);
nor U13233 (N_13233,N_11166,N_11285);
and U13234 (N_13234,N_10229,N_10938);
nand U13235 (N_13235,N_11295,N_11782);
nor U13236 (N_13236,N_11848,N_9736);
or U13237 (N_13237,N_11583,N_10854);
nor U13238 (N_13238,N_10481,N_11684);
xor U13239 (N_13239,N_10153,N_9250);
xnor U13240 (N_13240,N_11856,N_9460);
or U13241 (N_13241,N_11943,N_10381);
nand U13242 (N_13242,N_9047,N_9515);
nand U13243 (N_13243,N_11775,N_10386);
nor U13244 (N_13244,N_11080,N_10199);
nand U13245 (N_13245,N_10704,N_10803);
nand U13246 (N_13246,N_9300,N_11124);
nand U13247 (N_13247,N_10678,N_10510);
nand U13248 (N_13248,N_11612,N_10551);
and U13249 (N_13249,N_9275,N_9891);
nor U13250 (N_13250,N_11738,N_9172);
nor U13251 (N_13251,N_9410,N_9769);
and U13252 (N_13252,N_11403,N_10682);
or U13253 (N_13253,N_11438,N_11203);
and U13254 (N_13254,N_11474,N_9930);
or U13255 (N_13255,N_11050,N_9795);
and U13256 (N_13256,N_10877,N_9028);
or U13257 (N_13257,N_10109,N_11869);
or U13258 (N_13258,N_9175,N_9675);
xnor U13259 (N_13259,N_9302,N_11471);
or U13260 (N_13260,N_11568,N_10915);
or U13261 (N_13261,N_9470,N_11767);
nor U13262 (N_13262,N_11042,N_11492);
and U13263 (N_13263,N_10702,N_11596);
or U13264 (N_13264,N_9847,N_9020);
or U13265 (N_13265,N_11835,N_10798);
xnor U13266 (N_13266,N_9212,N_9580);
nand U13267 (N_13267,N_9694,N_11501);
and U13268 (N_13268,N_9133,N_10264);
and U13269 (N_13269,N_10315,N_9127);
nor U13270 (N_13270,N_9506,N_9772);
or U13271 (N_13271,N_11935,N_9421);
and U13272 (N_13272,N_11538,N_11780);
nor U13273 (N_13273,N_11790,N_11300);
or U13274 (N_13274,N_9810,N_9422);
and U13275 (N_13275,N_9164,N_11641);
nand U13276 (N_13276,N_11755,N_11142);
nor U13277 (N_13277,N_11662,N_9119);
nand U13278 (N_13278,N_9809,N_9939);
nand U13279 (N_13279,N_11113,N_11227);
nand U13280 (N_13280,N_9010,N_9094);
and U13281 (N_13281,N_10723,N_9893);
nand U13282 (N_13282,N_11306,N_10429);
or U13283 (N_13283,N_9056,N_9356);
nand U13284 (N_13284,N_11287,N_11414);
nand U13285 (N_13285,N_9051,N_10595);
nor U13286 (N_13286,N_9418,N_11899);
nand U13287 (N_13287,N_9751,N_9956);
nor U13288 (N_13288,N_11997,N_9102);
or U13289 (N_13289,N_11751,N_11756);
and U13290 (N_13290,N_10333,N_11834);
or U13291 (N_13291,N_9191,N_9425);
nor U13292 (N_13292,N_9708,N_9225);
nor U13293 (N_13293,N_11857,N_11508);
nand U13294 (N_13294,N_10709,N_9244);
nand U13295 (N_13295,N_9467,N_9854);
or U13296 (N_13296,N_11668,N_9291);
and U13297 (N_13297,N_11578,N_10356);
nand U13298 (N_13298,N_9341,N_10174);
and U13299 (N_13299,N_10083,N_10483);
xnor U13300 (N_13300,N_9630,N_9143);
and U13301 (N_13301,N_10946,N_10516);
nand U13302 (N_13302,N_11850,N_10733);
and U13303 (N_13303,N_11316,N_10351);
nor U13304 (N_13304,N_9657,N_10885);
nor U13305 (N_13305,N_9229,N_10321);
or U13306 (N_13306,N_11879,N_9648);
and U13307 (N_13307,N_10490,N_11072);
nand U13308 (N_13308,N_11389,N_9601);
nand U13309 (N_13309,N_9464,N_11454);
and U13310 (N_13310,N_10414,N_11263);
nor U13311 (N_13311,N_9859,N_10103);
and U13312 (N_13312,N_9430,N_10808);
and U13313 (N_13313,N_9724,N_11818);
nand U13314 (N_13314,N_11690,N_9477);
and U13315 (N_13315,N_10032,N_10128);
nor U13316 (N_13316,N_9063,N_11622);
nand U13317 (N_13317,N_11791,N_11358);
nand U13318 (N_13318,N_11977,N_9448);
nand U13319 (N_13319,N_10572,N_10777);
nand U13320 (N_13320,N_11241,N_9620);
nor U13321 (N_13321,N_9248,N_11605);
or U13322 (N_13322,N_9682,N_11215);
xor U13323 (N_13323,N_10943,N_11773);
nor U13324 (N_13324,N_10581,N_9861);
and U13325 (N_13325,N_9471,N_11398);
nand U13326 (N_13326,N_11408,N_11889);
nor U13327 (N_13327,N_10677,N_10215);
nand U13328 (N_13328,N_9903,N_9944);
nand U13329 (N_13329,N_11008,N_10162);
nand U13330 (N_13330,N_10392,N_10435);
and U13331 (N_13331,N_11646,N_9782);
or U13332 (N_13332,N_10570,N_10293);
nand U13333 (N_13333,N_9929,N_11433);
or U13334 (N_13334,N_9426,N_9492);
or U13335 (N_13335,N_10484,N_10976);
and U13336 (N_13336,N_10903,N_10141);
or U13337 (N_13337,N_9994,N_9442);
nor U13338 (N_13338,N_9106,N_11839);
nor U13339 (N_13339,N_10790,N_10937);
or U13340 (N_13340,N_9504,N_10597);
nor U13341 (N_13341,N_11732,N_10158);
or U13342 (N_13342,N_10212,N_9406);
and U13343 (N_13343,N_11491,N_9036);
and U13344 (N_13344,N_10469,N_10855);
and U13345 (N_13345,N_9663,N_11363);
or U13346 (N_13346,N_9590,N_9845);
and U13347 (N_13347,N_11346,N_11703);
nor U13348 (N_13348,N_11421,N_9233);
and U13349 (N_13349,N_10355,N_10988);
or U13350 (N_13350,N_10892,N_10271);
nor U13351 (N_13351,N_10827,N_11017);
or U13352 (N_13352,N_11960,N_11827);
and U13353 (N_13353,N_11584,N_10121);
or U13354 (N_13354,N_9583,N_10756);
or U13355 (N_13355,N_11569,N_9990);
xor U13356 (N_13356,N_11941,N_9807);
and U13357 (N_13357,N_11784,N_10644);
nand U13358 (N_13358,N_9560,N_10562);
nor U13359 (N_13359,N_10220,N_9062);
nor U13360 (N_13360,N_9978,N_10883);
nor U13361 (N_13361,N_11701,N_11312);
and U13362 (N_13362,N_10802,N_11676);
nor U13363 (N_13363,N_10660,N_9631);
and U13364 (N_13364,N_11253,N_11372);
or U13365 (N_13365,N_10225,N_11000);
or U13366 (N_13366,N_11048,N_11132);
and U13367 (N_13367,N_11691,N_11897);
nand U13368 (N_13368,N_11795,N_11489);
nand U13369 (N_13369,N_11636,N_10004);
and U13370 (N_13370,N_9697,N_10497);
nand U13371 (N_13371,N_10758,N_10914);
nand U13372 (N_13372,N_9336,N_11266);
nand U13373 (N_13373,N_11244,N_10442);
nand U13374 (N_13374,N_10408,N_11160);
and U13375 (N_13375,N_10379,N_9282);
or U13376 (N_13376,N_9732,N_9798);
nor U13377 (N_13377,N_10294,N_9738);
or U13378 (N_13378,N_9572,N_9454);
or U13379 (N_13379,N_10221,N_9979);
nor U13380 (N_13380,N_9712,N_11549);
and U13381 (N_13381,N_11249,N_10917);
nor U13382 (N_13382,N_10393,N_9026);
and U13383 (N_13383,N_10554,N_11618);
and U13384 (N_13384,N_11405,N_11555);
nor U13385 (N_13385,N_11320,N_10748);
nand U13386 (N_13386,N_10310,N_10653);
and U13387 (N_13387,N_11813,N_10124);
and U13388 (N_13388,N_10459,N_10014);
nand U13389 (N_13389,N_9987,N_11762);
nor U13390 (N_13390,N_10425,N_10498);
and U13391 (N_13391,N_9395,N_9958);
nor U13392 (N_13392,N_9710,N_11171);
and U13393 (N_13393,N_10579,N_10761);
nor U13394 (N_13394,N_10122,N_11460);
nor U13395 (N_13395,N_10652,N_9357);
nor U13396 (N_13396,N_9728,N_11744);
or U13397 (N_13397,N_11620,N_9519);
nor U13398 (N_13398,N_9817,N_11167);
and U13399 (N_13399,N_10560,N_10362);
or U13400 (N_13400,N_10926,N_9075);
nor U13401 (N_13401,N_11544,N_9988);
nor U13402 (N_13402,N_9203,N_9816);
and U13403 (N_13403,N_11178,N_10558);
nor U13404 (N_13404,N_11292,N_9514);
xnor U13405 (N_13405,N_9545,N_10022);
and U13406 (N_13406,N_10626,N_11187);
and U13407 (N_13407,N_11824,N_9822);
nand U13408 (N_13408,N_11293,N_10465);
nand U13409 (N_13409,N_9524,N_11156);
and U13410 (N_13410,N_9550,N_10902);
and U13411 (N_13411,N_9372,N_9674);
nor U13412 (N_13412,N_11302,N_10669);
nand U13413 (N_13413,N_9011,N_10336);
nand U13414 (N_13414,N_11776,N_10841);
and U13415 (N_13415,N_11980,N_11059);
nor U13416 (N_13416,N_11220,N_11591);
or U13417 (N_13417,N_10492,N_9096);
nand U13418 (N_13418,N_11901,N_11174);
and U13419 (N_13419,N_9309,N_9870);
or U13420 (N_13420,N_10243,N_10556);
and U13421 (N_13421,N_9922,N_10714);
and U13422 (N_13422,N_9333,N_10840);
nand U13423 (N_13423,N_11112,N_11865);
nand U13424 (N_13424,N_11494,N_9667);
nand U13425 (N_13425,N_11001,N_10378);
or U13426 (N_13426,N_9600,N_11532);
and U13427 (N_13427,N_9734,N_10072);
nor U13428 (N_13428,N_9853,N_11270);
nand U13429 (N_13429,N_9424,N_10143);
or U13430 (N_13430,N_10384,N_9670);
or U13431 (N_13431,N_11222,N_10975);
nor U13432 (N_13432,N_10292,N_11459);
and U13433 (N_13433,N_11388,N_10952);
and U13434 (N_13434,N_10641,N_11830);
nand U13435 (N_13435,N_10541,N_9142);
or U13436 (N_13436,N_9948,N_11840);
nand U13437 (N_13437,N_9593,N_11769);
and U13438 (N_13438,N_10119,N_10284);
nand U13439 (N_13439,N_11868,N_11966);
and U13440 (N_13440,N_10361,N_10047);
and U13441 (N_13441,N_9013,N_11170);
and U13442 (N_13442,N_11930,N_11031);
or U13443 (N_13443,N_10998,N_10833);
and U13444 (N_13444,N_9131,N_9087);
nand U13445 (N_13445,N_9587,N_9049);
or U13446 (N_13446,N_9608,N_9731);
nand U13447 (N_13447,N_9829,N_11973);
nor U13448 (N_13448,N_9446,N_10639);
or U13449 (N_13449,N_11444,N_9808);
nor U13450 (N_13450,N_11627,N_11853);
or U13451 (N_13451,N_10967,N_10473);
and U13452 (N_13452,N_10785,N_9304);
nand U13453 (N_13453,N_9443,N_9921);
nand U13454 (N_13454,N_9277,N_9725);
nor U13455 (N_13455,N_11540,N_10731);
nor U13456 (N_13456,N_10900,N_10147);
and U13457 (N_13457,N_9040,N_10593);
and U13458 (N_13458,N_9681,N_11434);
and U13459 (N_13459,N_9945,N_10625);
or U13460 (N_13460,N_11900,N_9375);
nor U13461 (N_13461,N_10739,N_11044);
nand U13462 (N_13462,N_11004,N_11326);
nand U13463 (N_13463,N_10567,N_10245);
nor U13464 (N_13464,N_10962,N_10208);
or U13465 (N_13465,N_11026,N_11078);
and U13466 (N_13466,N_10796,N_9940);
and U13467 (N_13467,N_9435,N_9358);
nand U13468 (N_13468,N_10427,N_9097);
or U13469 (N_13469,N_11659,N_9673);
nor U13470 (N_13470,N_11391,N_11313);
or U13471 (N_13471,N_10449,N_10400);
nand U13472 (N_13472,N_11394,N_10502);
and U13473 (N_13473,N_10847,N_11763);
nor U13474 (N_13474,N_9546,N_9777);
and U13475 (N_13475,N_11463,N_11693);
or U13476 (N_13476,N_11545,N_11005);
nand U13477 (N_13477,N_10402,N_10876);
and U13478 (N_13478,N_9604,N_9239);
or U13479 (N_13479,N_11445,N_10869);
nand U13480 (N_13480,N_9003,N_11746);
nand U13481 (N_13481,N_10059,N_10853);
nand U13482 (N_13482,N_10300,N_10613);
nand U13483 (N_13483,N_9792,N_10209);
nor U13484 (N_13484,N_11907,N_11333);
or U13485 (N_13485,N_9221,N_10746);
or U13486 (N_13486,N_11672,N_11136);
and U13487 (N_13487,N_11116,N_11409);
or U13488 (N_13488,N_11895,N_10048);
nor U13489 (N_13489,N_10219,N_11151);
nand U13490 (N_13490,N_11654,N_11425);
nand U13491 (N_13491,N_11435,N_10940);
and U13492 (N_13492,N_10202,N_10754);
nand U13493 (N_13493,N_10369,N_10140);
or U13494 (N_13494,N_9338,N_9368);
and U13495 (N_13495,N_10518,N_11774);
or U13496 (N_13496,N_9885,N_10700);
or U13497 (N_13497,N_11456,N_10241);
nand U13498 (N_13498,N_10191,N_10889);
or U13499 (N_13499,N_11035,N_11176);
nand U13500 (N_13500,N_10071,N_10595);
or U13501 (N_13501,N_11414,N_11806);
or U13502 (N_13502,N_9072,N_10541);
nor U13503 (N_13503,N_11408,N_10641);
nand U13504 (N_13504,N_11982,N_10472);
nand U13505 (N_13505,N_11517,N_9737);
nand U13506 (N_13506,N_11187,N_10368);
and U13507 (N_13507,N_11181,N_11921);
nand U13508 (N_13508,N_10608,N_10837);
nor U13509 (N_13509,N_9062,N_10234);
and U13510 (N_13510,N_11075,N_11704);
and U13511 (N_13511,N_10980,N_10462);
nand U13512 (N_13512,N_10251,N_10523);
nand U13513 (N_13513,N_9865,N_11557);
and U13514 (N_13514,N_11082,N_11420);
xor U13515 (N_13515,N_9320,N_10188);
and U13516 (N_13516,N_11455,N_11444);
and U13517 (N_13517,N_9818,N_9405);
and U13518 (N_13518,N_9139,N_9670);
or U13519 (N_13519,N_9024,N_11032);
or U13520 (N_13520,N_9167,N_9036);
nor U13521 (N_13521,N_11693,N_9464);
nor U13522 (N_13522,N_9337,N_9292);
or U13523 (N_13523,N_9333,N_9151);
nor U13524 (N_13524,N_10674,N_10665);
or U13525 (N_13525,N_10968,N_10879);
and U13526 (N_13526,N_9550,N_10027);
or U13527 (N_13527,N_9425,N_11336);
nor U13528 (N_13528,N_11947,N_10768);
nor U13529 (N_13529,N_9764,N_10070);
or U13530 (N_13530,N_9357,N_9762);
nand U13531 (N_13531,N_10606,N_10170);
or U13532 (N_13532,N_9303,N_10531);
and U13533 (N_13533,N_11769,N_11299);
or U13534 (N_13534,N_9647,N_11681);
nor U13535 (N_13535,N_11869,N_9776);
nand U13536 (N_13536,N_11293,N_10244);
nand U13537 (N_13537,N_11981,N_11468);
and U13538 (N_13538,N_11187,N_11991);
nand U13539 (N_13539,N_11385,N_9364);
nor U13540 (N_13540,N_10485,N_10446);
and U13541 (N_13541,N_9681,N_10279);
nand U13542 (N_13542,N_11402,N_11634);
nand U13543 (N_13543,N_11568,N_11550);
nand U13544 (N_13544,N_9038,N_10912);
and U13545 (N_13545,N_10304,N_10081);
and U13546 (N_13546,N_11110,N_11393);
nand U13547 (N_13547,N_9355,N_11425);
nand U13548 (N_13548,N_11780,N_9238);
or U13549 (N_13549,N_11146,N_11256);
nor U13550 (N_13550,N_11012,N_11145);
nand U13551 (N_13551,N_10565,N_9702);
nor U13552 (N_13552,N_11117,N_9727);
nor U13553 (N_13553,N_10733,N_10551);
or U13554 (N_13554,N_10957,N_10908);
and U13555 (N_13555,N_11792,N_11648);
or U13556 (N_13556,N_11146,N_11000);
nand U13557 (N_13557,N_10571,N_10966);
nand U13558 (N_13558,N_10525,N_9800);
or U13559 (N_13559,N_11443,N_11319);
and U13560 (N_13560,N_9589,N_11224);
xor U13561 (N_13561,N_11368,N_9955);
nand U13562 (N_13562,N_10178,N_11401);
nand U13563 (N_13563,N_9452,N_9351);
and U13564 (N_13564,N_9754,N_11395);
nand U13565 (N_13565,N_10131,N_10411);
or U13566 (N_13566,N_11948,N_10282);
nand U13567 (N_13567,N_10919,N_11679);
nand U13568 (N_13568,N_9575,N_11102);
nor U13569 (N_13569,N_11478,N_9986);
or U13570 (N_13570,N_9326,N_9644);
nand U13571 (N_13571,N_9384,N_11127);
or U13572 (N_13572,N_9367,N_9530);
nand U13573 (N_13573,N_11441,N_9046);
nand U13574 (N_13574,N_11968,N_11769);
or U13575 (N_13575,N_11227,N_10591);
or U13576 (N_13576,N_9521,N_11296);
nor U13577 (N_13577,N_9812,N_9463);
and U13578 (N_13578,N_9906,N_9136);
or U13579 (N_13579,N_11338,N_10234);
nand U13580 (N_13580,N_10691,N_11035);
nand U13581 (N_13581,N_9067,N_9777);
nand U13582 (N_13582,N_10618,N_11299);
nor U13583 (N_13583,N_10139,N_9566);
or U13584 (N_13584,N_9589,N_11197);
nor U13585 (N_13585,N_9989,N_9661);
nand U13586 (N_13586,N_11506,N_9779);
or U13587 (N_13587,N_11689,N_10745);
or U13588 (N_13588,N_11263,N_11493);
nand U13589 (N_13589,N_9037,N_9494);
nand U13590 (N_13590,N_10593,N_11589);
or U13591 (N_13591,N_10313,N_9053);
nand U13592 (N_13592,N_9603,N_9520);
nor U13593 (N_13593,N_11428,N_9153);
nand U13594 (N_13594,N_10360,N_11636);
nand U13595 (N_13595,N_10181,N_10554);
and U13596 (N_13596,N_10475,N_9659);
or U13597 (N_13597,N_9496,N_9444);
and U13598 (N_13598,N_9074,N_11608);
nor U13599 (N_13599,N_11088,N_11856);
and U13600 (N_13600,N_11756,N_10038);
and U13601 (N_13601,N_10553,N_10942);
and U13602 (N_13602,N_10278,N_10476);
nand U13603 (N_13603,N_9243,N_11287);
nand U13604 (N_13604,N_11182,N_11580);
or U13605 (N_13605,N_11562,N_11810);
and U13606 (N_13606,N_11836,N_9685);
and U13607 (N_13607,N_11402,N_10093);
or U13608 (N_13608,N_11907,N_9285);
or U13609 (N_13609,N_10583,N_10987);
and U13610 (N_13610,N_9120,N_10502);
or U13611 (N_13611,N_10108,N_9716);
nand U13612 (N_13612,N_10620,N_10230);
nor U13613 (N_13613,N_10256,N_10636);
nor U13614 (N_13614,N_9770,N_9438);
nor U13615 (N_13615,N_10177,N_11719);
and U13616 (N_13616,N_11162,N_9168);
nor U13617 (N_13617,N_9287,N_11748);
or U13618 (N_13618,N_9995,N_11144);
and U13619 (N_13619,N_11144,N_9074);
nand U13620 (N_13620,N_9055,N_10960);
or U13621 (N_13621,N_11125,N_11214);
or U13622 (N_13622,N_9487,N_10614);
and U13623 (N_13623,N_11421,N_11949);
and U13624 (N_13624,N_9475,N_9961);
or U13625 (N_13625,N_11348,N_11238);
and U13626 (N_13626,N_11354,N_9796);
and U13627 (N_13627,N_11106,N_11953);
nand U13628 (N_13628,N_10616,N_9016);
and U13629 (N_13629,N_9898,N_9057);
or U13630 (N_13630,N_9280,N_11133);
or U13631 (N_13631,N_9121,N_9165);
nand U13632 (N_13632,N_11608,N_9716);
nand U13633 (N_13633,N_11273,N_11994);
or U13634 (N_13634,N_10883,N_9894);
and U13635 (N_13635,N_9914,N_11346);
nor U13636 (N_13636,N_9651,N_10576);
and U13637 (N_13637,N_11711,N_11814);
nor U13638 (N_13638,N_11119,N_9718);
or U13639 (N_13639,N_10051,N_10391);
or U13640 (N_13640,N_10572,N_10897);
or U13641 (N_13641,N_9229,N_11173);
or U13642 (N_13642,N_10502,N_9216);
nor U13643 (N_13643,N_9872,N_10282);
and U13644 (N_13644,N_10294,N_10187);
and U13645 (N_13645,N_11089,N_11250);
nor U13646 (N_13646,N_10356,N_10875);
xor U13647 (N_13647,N_10059,N_11928);
nand U13648 (N_13648,N_10464,N_11630);
nor U13649 (N_13649,N_11341,N_9815);
nor U13650 (N_13650,N_10733,N_10269);
or U13651 (N_13651,N_10161,N_9602);
nor U13652 (N_13652,N_11792,N_11624);
nor U13653 (N_13653,N_11394,N_10638);
nand U13654 (N_13654,N_9780,N_10638);
nor U13655 (N_13655,N_9710,N_11475);
and U13656 (N_13656,N_9937,N_9415);
nand U13657 (N_13657,N_10766,N_11327);
or U13658 (N_13658,N_9284,N_9042);
nor U13659 (N_13659,N_9031,N_9808);
nand U13660 (N_13660,N_9349,N_11635);
nand U13661 (N_13661,N_9767,N_11942);
nand U13662 (N_13662,N_11951,N_10422);
or U13663 (N_13663,N_9222,N_11688);
or U13664 (N_13664,N_11468,N_11629);
nor U13665 (N_13665,N_10475,N_10846);
nor U13666 (N_13666,N_11491,N_11039);
nand U13667 (N_13667,N_10935,N_10257);
or U13668 (N_13668,N_10203,N_9642);
and U13669 (N_13669,N_10581,N_9072);
nand U13670 (N_13670,N_10732,N_11262);
nor U13671 (N_13671,N_10261,N_10064);
and U13672 (N_13672,N_11450,N_10983);
and U13673 (N_13673,N_10307,N_9687);
and U13674 (N_13674,N_9257,N_10500);
or U13675 (N_13675,N_9702,N_10482);
nand U13676 (N_13676,N_11662,N_11221);
nand U13677 (N_13677,N_9754,N_11417);
nor U13678 (N_13678,N_11273,N_11656);
and U13679 (N_13679,N_9851,N_11838);
nor U13680 (N_13680,N_9661,N_10432);
and U13681 (N_13681,N_11622,N_9859);
nor U13682 (N_13682,N_9309,N_9818);
nand U13683 (N_13683,N_10685,N_10583);
or U13684 (N_13684,N_9974,N_11402);
nand U13685 (N_13685,N_11525,N_11243);
nor U13686 (N_13686,N_10374,N_10253);
or U13687 (N_13687,N_11938,N_9327);
nor U13688 (N_13688,N_10722,N_10759);
nand U13689 (N_13689,N_9729,N_9769);
and U13690 (N_13690,N_10745,N_11651);
and U13691 (N_13691,N_11466,N_9674);
nor U13692 (N_13692,N_10938,N_10860);
nand U13693 (N_13693,N_9848,N_11641);
nand U13694 (N_13694,N_9547,N_10178);
nand U13695 (N_13695,N_11459,N_10483);
and U13696 (N_13696,N_9224,N_10468);
nand U13697 (N_13697,N_10210,N_10288);
or U13698 (N_13698,N_9557,N_11845);
nand U13699 (N_13699,N_11581,N_11689);
and U13700 (N_13700,N_11841,N_11174);
nand U13701 (N_13701,N_11409,N_11237);
and U13702 (N_13702,N_10619,N_10116);
and U13703 (N_13703,N_9357,N_9034);
or U13704 (N_13704,N_9369,N_11352);
and U13705 (N_13705,N_10704,N_9219);
and U13706 (N_13706,N_11764,N_9761);
and U13707 (N_13707,N_10528,N_11880);
nor U13708 (N_13708,N_10039,N_9312);
and U13709 (N_13709,N_10335,N_9427);
and U13710 (N_13710,N_11755,N_11480);
and U13711 (N_13711,N_9461,N_10163);
and U13712 (N_13712,N_10154,N_10707);
or U13713 (N_13713,N_9665,N_10695);
nand U13714 (N_13714,N_10223,N_11633);
nor U13715 (N_13715,N_11320,N_10247);
nand U13716 (N_13716,N_10315,N_10924);
xnor U13717 (N_13717,N_10928,N_11745);
and U13718 (N_13718,N_10382,N_9842);
nand U13719 (N_13719,N_10764,N_10128);
or U13720 (N_13720,N_11888,N_11069);
or U13721 (N_13721,N_10006,N_10193);
nand U13722 (N_13722,N_11845,N_10826);
or U13723 (N_13723,N_10779,N_11532);
and U13724 (N_13724,N_9697,N_9220);
and U13725 (N_13725,N_10395,N_10504);
or U13726 (N_13726,N_9472,N_10758);
nand U13727 (N_13727,N_9113,N_10490);
nand U13728 (N_13728,N_11781,N_9422);
and U13729 (N_13729,N_9324,N_10181);
nand U13730 (N_13730,N_11270,N_10225);
or U13731 (N_13731,N_10873,N_10615);
and U13732 (N_13732,N_10792,N_9278);
and U13733 (N_13733,N_9519,N_11094);
or U13734 (N_13734,N_11629,N_10527);
or U13735 (N_13735,N_10820,N_11693);
or U13736 (N_13736,N_9797,N_9427);
nand U13737 (N_13737,N_9817,N_10010);
xnor U13738 (N_13738,N_10670,N_10835);
and U13739 (N_13739,N_11682,N_11994);
nand U13740 (N_13740,N_11716,N_10578);
nor U13741 (N_13741,N_9791,N_11677);
and U13742 (N_13742,N_10018,N_11192);
nor U13743 (N_13743,N_11609,N_11116);
or U13744 (N_13744,N_9281,N_10747);
nor U13745 (N_13745,N_9115,N_10730);
or U13746 (N_13746,N_10595,N_11137);
and U13747 (N_13747,N_10994,N_9035);
nor U13748 (N_13748,N_9787,N_9564);
or U13749 (N_13749,N_11670,N_11486);
and U13750 (N_13750,N_10699,N_9572);
and U13751 (N_13751,N_9071,N_10945);
or U13752 (N_13752,N_11412,N_11328);
nand U13753 (N_13753,N_11773,N_10443);
xnor U13754 (N_13754,N_10051,N_10671);
nor U13755 (N_13755,N_10924,N_11362);
and U13756 (N_13756,N_11280,N_9595);
nand U13757 (N_13757,N_9368,N_10561);
nor U13758 (N_13758,N_10428,N_10717);
or U13759 (N_13759,N_9319,N_10987);
and U13760 (N_13760,N_11872,N_11855);
or U13761 (N_13761,N_11508,N_10886);
or U13762 (N_13762,N_9131,N_9297);
and U13763 (N_13763,N_10881,N_10469);
nand U13764 (N_13764,N_10969,N_11644);
nor U13765 (N_13765,N_9158,N_11467);
nor U13766 (N_13766,N_9865,N_9742);
or U13767 (N_13767,N_9459,N_9435);
nor U13768 (N_13768,N_11321,N_11795);
nor U13769 (N_13769,N_10132,N_10892);
and U13770 (N_13770,N_9605,N_11620);
nand U13771 (N_13771,N_9023,N_10019);
and U13772 (N_13772,N_10961,N_10100);
nand U13773 (N_13773,N_9312,N_10607);
nand U13774 (N_13774,N_11799,N_11022);
and U13775 (N_13775,N_11291,N_10790);
nor U13776 (N_13776,N_9614,N_10232);
or U13777 (N_13777,N_9928,N_11393);
and U13778 (N_13778,N_10740,N_10867);
and U13779 (N_13779,N_10476,N_9382);
or U13780 (N_13780,N_11331,N_9154);
nand U13781 (N_13781,N_9570,N_10107);
nor U13782 (N_13782,N_10813,N_11884);
and U13783 (N_13783,N_11038,N_10135);
nand U13784 (N_13784,N_10721,N_9564);
or U13785 (N_13785,N_11572,N_9502);
nor U13786 (N_13786,N_9665,N_9457);
nor U13787 (N_13787,N_11733,N_10209);
nor U13788 (N_13788,N_10853,N_9049);
nor U13789 (N_13789,N_11207,N_10907);
nand U13790 (N_13790,N_11531,N_10332);
and U13791 (N_13791,N_9198,N_10355);
or U13792 (N_13792,N_11414,N_11063);
nor U13793 (N_13793,N_10079,N_10267);
nor U13794 (N_13794,N_11216,N_11651);
nor U13795 (N_13795,N_10454,N_10326);
nor U13796 (N_13796,N_9738,N_11186);
nor U13797 (N_13797,N_10742,N_9170);
nand U13798 (N_13798,N_10455,N_9705);
nor U13799 (N_13799,N_9569,N_9800);
or U13800 (N_13800,N_11928,N_9857);
and U13801 (N_13801,N_10273,N_10724);
and U13802 (N_13802,N_10034,N_10747);
and U13803 (N_13803,N_9551,N_9978);
or U13804 (N_13804,N_11730,N_9588);
nand U13805 (N_13805,N_10778,N_10587);
nand U13806 (N_13806,N_10648,N_9291);
and U13807 (N_13807,N_10413,N_10075);
nand U13808 (N_13808,N_10959,N_9634);
or U13809 (N_13809,N_10310,N_11095);
and U13810 (N_13810,N_9737,N_11339);
and U13811 (N_13811,N_9846,N_10119);
or U13812 (N_13812,N_9168,N_11138);
or U13813 (N_13813,N_9945,N_10980);
and U13814 (N_13814,N_10611,N_11223);
nor U13815 (N_13815,N_11051,N_10344);
and U13816 (N_13816,N_11805,N_9069);
nor U13817 (N_13817,N_9552,N_10405);
nor U13818 (N_13818,N_9697,N_9503);
nor U13819 (N_13819,N_9311,N_9453);
nand U13820 (N_13820,N_9529,N_10005);
or U13821 (N_13821,N_9205,N_10280);
or U13822 (N_13822,N_11461,N_9838);
and U13823 (N_13823,N_10884,N_11652);
and U13824 (N_13824,N_10404,N_9294);
and U13825 (N_13825,N_10967,N_9419);
or U13826 (N_13826,N_9430,N_10075);
or U13827 (N_13827,N_9742,N_9389);
nor U13828 (N_13828,N_11895,N_11685);
and U13829 (N_13829,N_11565,N_10082);
nand U13830 (N_13830,N_11866,N_11587);
or U13831 (N_13831,N_11675,N_10828);
and U13832 (N_13832,N_10331,N_10816);
and U13833 (N_13833,N_11848,N_9742);
or U13834 (N_13834,N_10460,N_9985);
xnor U13835 (N_13835,N_10939,N_10437);
and U13836 (N_13836,N_11834,N_9670);
nor U13837 (N_13837,N_9084,N_11993);
and U13838 (N_13838,N_11701,N_10738);
nand U13839 (N_13839,N_11413,N_11787);
nor U13840 (N_13840,N_9010,N_11497);
or U13841 (N_13841,N_9647,N_9620);
or U13842 (N_13842,N_11633,N_9276);
nand U13843 (N_13843,N_10617,N_10512);
nand U13844 (N_13844,N_10558,N_10261);
and U13845 (N_13845,N_11430,N_10539);
nor U13846 (N_13846,N_11338,N_11421);
or U13847 (N_13847,N_10433,N_10781);
nand U13848 (N_13848,N_10511,N_11057);
or U13849 (N_13849,N_11804,N_11862);
nor U13850 (N_13850,N_10255,N_10034);
and U13851 (N_13851,N_10825,N_11334);
nor U13852 (N_13852,N_10375,N_11358);
and U13853 (N_13853,N_10380,N_9977);
nor U13854 (N_13854,N_11172,N_11878);
nor U13855 (N_13855,N_10677,N_9780);
nand U13856 (N_13856,N_11767,N_11580);
or U13857 (N_13857,N_11932,N_9963);
nor U13858 (N_13858,N_11978,N_9324);
and U13859 (N_13859,N_9816,N_9445);
nand U13860 (N_13860,N_11749,N_10350);
nor U13861 (N_13861,N_9259,N_10938);
or U13862 (N_13862,N_10358,N_11994);
and U13863 (N_13863,N_11580,N_10847);
and U13864 (N_13864,N_10123,N_10813);
and U13865 (N_13865,N_11688,N_11955);
nor U13866 (N_13866,N_10521,N_9716);
and U13867 (N_13867,N_9267,N_9232);
nand U13868 (N_13868,N_11015,N_9691);
and U13869 (N_13869,N_10399,N_9101);
and U13870 (N_13870,N_10210,N_10382);
and U13871 (N_13871,N_10176,N_11768);
nand U13872 (N_13872,N_9906,N_11110);
and U13873 (N_13873,N_10057,N_9572);
or U13874 (N_13874,N_11002,N_11811);
nor U13875 (N_13875,N_11655,N_10637);
nor U13876 (N_13876,N_9025,N_9727);
and U13877 (N_13877,N_10060,N_9983);
nor U13878 (N_13878,N_9383,N_11997);
nand U13879 (N_13879,N_11836,N_10915);
and U13880 (N_13880,N_10347,N_10164);
nor U13881 (N_13881,N_11935,N_11686);
xnor U13882 (N_13882,N_9064,N_11454);
nand U13883 (N_13883,N_9114,N_9148);
or U13884 (N_13884,N_10151,N_11996);
nand U13885 (N_13885,N_11491,N_9180);
or U13886 (N_13886,N_11747,N_10358);
nand U13887 (N_13887,N_10617,N_9588);
xnor U13888 (N_13888,N_9239,N_10242);
nand U13889 (N_13889,N_10499,N_10073);
xor U13890 (N_13890,N_10013,N_11717);
nor U13891 (N_13891,N_9284,N_11037);
or U13892 (N_13892,N_11205,N_10973);
nor U13893 (N_13893,N_9881,N_11266);
nand U13894 (N_13894,N_9923,N_10342);
or U13895 (N_13895,N_10117,N_9504);
nor U13896 (N_13896,N_9348,N_9795);
nor U13897 (N_13897,N_11470,N_10075);
nor U13898 (N_13898,N_10979,N_10061);
or U13899 (N_13899,N_10242,N_11315);
or U13900 (N_13900,N_10987,N_11025);
nand U13901 (N_13901,N_11979,N_9384);
nand U13902 (N_13902,N_10884,N_9067);
and U13903 (N_13903,N_10810,N_10787);
nor U13904 (N_13904,N_11989,N_9163);
nand U13905 (N_13905,N_10206,N_11970);
and U13906 (N_13906,N_11160,N_9749);
nor U13907 (N_13907,N_9930,N_10693);
nor U13908 (N_13908,N_11651,N_11685);
and U13909 (N_13909,N_11545,N_10021);
nand U13910 (N_13910,N_11952,N_10734);
or U13911 (N_13911,N_11425,N_10416);
nor U13912 (N_13912,N_11756,N_11820);
or U13913 (N_13913,N_9771,N_10935);
and U13914 (N_13914,N_10217,N_11720);
or U13915 (N_13915,N_10908,N_10412);
nor U13916 (N_13916,N_10274,N_9070);
nor U13917 (N_13917,N_9938,N_9285);
nand U13918 (N_13918,N_11105,N_11711);
nor U13919 (N_13919,N_9073,N_10089);
nor U13920 (N_13920,N_11337,N_11164);
nor U13921 (N_13921,N_10207,N_10650);
or U13922 (N_13922,N_9240,N_9638);
xor U13923 (N_13923,N_9018,N_11244);
nand U13924 (N_13924,N_10396,N_11031);
or U13925 (N_13925,N_10483,N_11556);
nor U13926 (N_13926,N_10598,N_9333);
xor U13927 (N_13927,N_9565,N_11368);
or U13928 (N_13928,N_9559,N_11411);
nand U13929 (N_13929,N_10040,N_10770);
and U13930 (N_13930,N_11943,N_9353);
nand U13931 (N_13931,N_10259,N_11701);
nor U13932 (N_13932,N_11963,N_9348);
and U13933 (N_13933,N_11538,N_10638);
nand U13934 (N_13934,N_9082,N_11462);
nand U13935 (N_13935,N_11284,N_10850);
or U13936 (N_13936,N_9850,N_10052);
and U13937 (N_13937,N_9822,N_10217);
nand U13938 (N_13938,N_11568,N_10075);
nor U13939 (N_13939,N_10443,N_9586);
nand U13940 (N_13940,N_11832,N_11664);
or U13941 (N_13941,N_9238,N_10418);
or U13942 (N_13942,N_9214,N_11817);
nand U13943 (N_13943,N_9501,N_10790);
and U13944 (N_13944,N_10846,N_10918);
and U13945 (N_13945,N_9663,N_11870);
and U13946 (N_13946,N_10888,N_9758);
or U13947 (N_13947,N_10663,N_9112);
nand U13948 (N_13948,N_11344,N_11201);
and U13949 (N_13949,N_11808,N_11817);
or U13950 (N_13950,N_9644,N_9006);
or U13951 (N_13951,N_9940,N_10446);
and U13952 (N_13952,N_10463,N_11128);
and U13953 (N_13953,N_11836,N_10388);
or U13954 (N_13954,N_9935,N_11018);
xnor U13955 (N_13955,N_9107,N_11812);
nor U13956 (N_13956,N_9640,N_11960);
or U13957 (N_13957,N_9692,N_10896);
and U13958 (N_13958,N_11990,N_9832);
and U13959 (N_13959,N_9631,N_10312);
or U13960 (N_13960,N_10222,N_11723);
nand U13961 (N_13961,N_10175,N_10723);
nor U13962 (N_13962,N_9965,N_10896);
and U13963 (N_13963,N_11783,N_9140);
nand U13964 (N_13964,N_10704,N_9774);
or U13965 (N_13965,N_9873,N_11713);
or U13966 (N_13966,N_10425,N_10476);
nor U13967 (N_13967,N_9000,N_10540);
xor U13968 (N_13968,N_11842,N_9223);
and U13969 (N_13969,N_11205,N_10635);
or U13970 (N_13970,N_9854,N_9134);
or U13971 (N_13971,N_11564,N_9839);
and U13972 (N_13972,N_10609,N_9500);
and U13973 (N_13973,N_9861,N_11727);
or U13974 (N_13974,N_9642,N_9449);
xor U13975 (N_13975,N_11685,N_11928);
and U13976 (N_13976,N_10842,N_11381);
or U13977 (N_13977,N_10486,N_11551);
xor U13978 (N_13978,N_11467,N_9622);
or U13979 (N_13979,N_10373,N_11072);
nor U13980 (N_13980,N_9323,N_10523);
or U13981 (N_13981,N_11729,N_9214);
or U13982 (N_13982,N_10936,N_10290);
nand U13983 (N_13983,N_9358,N_10881);
nor U13984 (N_13984,N_10726,N_9259);
and U13985 (N_13985,N_10143,N_10020);
nand U13986 (N_13986,N_9241,N_11375);
or U13987 (N_13987,N_10092,N_9441);
nand U13988 (N_13988,N_9932,N_11054);
and U13989 (N_13989,N_9149,N_10105);
and U13990 (N_13990,N_9449,N_11754);
nand U13991 (N_13991,N_10944,N_9240);
nand U13992 (N_13992,N_9404,N_9084);
nand U13993 (N_13993,N_11758,N_10927);
nand U13994 (N_13994,N_9813,N_9686);
nand U13995 (N_13995,N_10587,N_11423);
or U13996 (N_13996,N_9222,N_11697);
nor U13997 (N_13997,N_10294,N_11225);
nand U13998 (N_13998,N_9422,N_11161);
or U13999 (N_13999,N_10176,N_11697);
nand U14000 (N_14000,N_11451,N_11426);
and U14001 (N_14001,N_11417,N_9409);
nor U14002 (N_14002,N_11728,N_11654);
or U14003 (N_14003,N_9644,N_10226);
nand U14004 (N_14004,N_10798,N_11120);
nand U14005 (N_14005,N_9777,N_10694);
or U14006 (N_14006,N_11675,N_11914);
nand U14007 (N_14007,N_10577,N_10630);
or U14008 (N_14008,N_11273,N_11723);
and U14009 (N_14009,N_11839,N_9553);
nand U14010 (N_14010,N_10674,N_9576);
nand U14011 (N_14011,N_9484,N_10673);
nor U14012 (N_14012,N_11850,N_11370);
nor U14013 (N_14013,N_11753,N_9365);
and U14014 (N_14014,N_10221,N_9494);
or U14015 (N_14015,N_9437,N_9479);
nand U14016 (N_14016,N_11146,N_9562);
and U14017 (N_14017,N_11787,N_11329);
nor U14018 (N_14018,N_9532,N_9704);
xor U14019 (N_14019,N_10169,N_11963);
nor U14020 (N_14020,N_10749,N_9144);
nand U14021 (N_14021,N_9563,N_11593);
nor U14022 (N_14022,N_9672,N_10488);
xor U14023 (N_14023,N_11008,N_11997);
nor U14024 (N_14024,N_11314,N_9104);
and U14025 (N_14025,N_9186,N_10183);
nand U14026 (N_14026,N_10225,N_9758);
and U14027 (N_14027,N_11148,N_10881);
or U14028 (N_14028,N_10463,N_9479);
nor U14029 (N_14029,N_11562,N_11649);
and U14030 (N_14030,N_9891,N_11816);
xor U14031 (N_14031,N_11216,N_9604);
and U14032 (N_14032,N_11315,N_9870);
and U14033 (N_14033,N_11658,N_11694);
or U14034 (N_14034,N_11955,N_10179);
nor U14035 (N_14035,N_9748,N_9311);
nor U14036 (N_14036,N_9335,N_9403);
nor U14037 (N_14037,N_11529,N_9155);
nor U14038 (N_14038,N_11545,N_11027);
or U14039 (N_14039,N_9205,N_11055);
or U14040 (N_14040,N_9706,N_9218);
nand U14041 (N_14041,N_10893,N_9177);
and U14042 (N_14042,N_9127,N_9160);
nor U14043 (N_14043,N_10741,N_11282);
and U14044 (N_14044,N_10170,N_9708);
and U14045 (N_14045,N_10324,N_11955);
or U14046 (N_14046,N_10720,N_11451);
nor U14047 (N_14047,N_10121,N_10813);
xor U14048 (N_14048,N_11262,N_9022);
or U14049 (N_14049,N_11005,N_11145);
or U14050 (N_14050,N_11242,N_9689);
and U14051 (N_14051,N_9152,N_11599);
and U14052 (N_14052,N_11948,N_9802);
xnor U14053 (N_14053,N_11222,N_9536);
or U14054 (N_14054,N_11146,N_10712);
nor U14055 (N_14055,N_9781,N_11507);
or U14056 (N_14056,N_9573,N_10508);
nand U14057 (N_14057,N_9843,N_10350);
nor U14058 (N_14058,N_9827,N_11267);
or U14059 (N_14059,N_10635,N_11387);
nor U14060 (N_14060,N_11970,N_9711);
xnor U14061 (N_14061,N_10769,N_10794);
or U14062 (N_14062,N_10073,N_9419);
nand U14063 (N_14063,N_11419,N_9217);
nor U14064 (N_14064,N_11723,N_9239);
and U14065 (N_14065,N_11987,N_9383);
nand U14066 (N_14066,N_11477,N_11960);
or U14067 (N_14067,N_10598,N_11946);
xor U14068 (N_14068,N_10796,N_9704);
nor U14069 (N_14069,N_11461,N_10403);
or U14070 (N_14070,N_10796,N_10683);
or U14071 (N_14071,N_10876,N_11030);
or U14072 (N_14072,N_9607,N_11697);
and U14073 (N_14073,N_9311,N_11211);
and U14074 (N_14074,N_9744,N_10633);
or U14075 (N_14075,N_11564,N_11234);
nand U14076 (N_14076,N_11966,N_10895);
nand U14077 (N_14077,N_9402,N_11314);
nand U14078 (N_14078,N_9262,N_9780);
or U14079 (N_14079,N_11246,N_10451);
nand U14080 (N_14080,N_11494,N_9470);
nor U14081 (N_14081,N_10805,N_10172);
or U14082 (N_14082,N_11837,N_9673);
and U14083 (N_14083,N_9376,N_11799);
or U14084 (N_14084,N_10535,N_11657);
or U14085 (N_14085,N_10620,N_10471);
nand U14086 (N_14086,N_10515,N_9731);
nor U14087 (N_14087,N_9022,N_9256);
nor U14088 (N_14088,N_11332,N_9110);
nor U14089 (N_14089,N_9933,N_11057);
nor U14090 (N_14090,N_9970,N_10706);
and U14091 (N_14091,N_9744,N_11087);
nor U14092 (N_14092,N_9517,N_11746);
nand U14093 (N_14093,N_11422,N_11660);
xor U14094 (N_14094,N_11649,N_9617);
nand U14095 (N_14095,N_10751,N_10619);
and U14096 (N_14096,N_11720,N_11576);
nand U14097 (N_14097,N_10022,N_9992);
nand U14098 (N_14098,N_11999,N_11210);
and U14099 (N_14099,N_10614,N_11408);
nand U14100 (N_14100,N_9609,N_9051);
nor U14101 (N_14101,N_11739,N_11459);
or U14102 (N_14102,N_9722,N_11147);
nor U14103 (N_14103,N_10414,N_11075);
nand U14104 (N_14104,N_11773,N_11306);
and U14105 (N_14105,N_11496,N_11193);
and U14106 (N_14106,N_10980,N_10207);
nand U14107 (N_14107,N_9390,N_11530);
nor U14108 (N_14108,N_11693,N_11316);
nand U14109 (N_14109,N_11500,N_11924);
and U14110 (N_14110,N_9455,N_9541);
or U14111 (N_14111,N_9605,N_9313);
nor U14112 (N_14112,N_10191,N_11897);
nand U14113 (N_14113,N_11263,N_9404);
nand U14114 (N_14114,N_10075,N_10563);
or U14115 (N_14115,N_9803,N_11600);
xor U14116 (N_14116,N_11296,N_11735);
and U14117 (N_14117,N_11646,N_11569);
xor U14118 (N_14118,N_10466,N_9080);
nand U14119 (N_14119,N_11961,N_9257);
and U14120 (N_14120,N_9610,N_9571);
nand U14121 (N_14121,N_9799,N_11711);
nand U14122 (N_14122,N_11526,N_9910);
nand U14123 (N_14123,N_9706,N_10847);
or U14124 (N_14124,N_11270,N_9460);
and U14125 (N_14125,N_9184,N_11009);
and U14126 (N_14126,N_9852,N_10174);
nor U14127 (N_14127,N_11986,N_11923);
nand U14128 (N_14128,N_11217,N_11483);
nor U14129 (N_14129,N_9606,N_9267);
nand U14130 (N_14130,N_10046,N_11986);
xor U14131 (N_14131,N_11375,N_11700);
nand U14132 (N_14132,N_10293,N_10838);
and U14133 (N_14133,N_9159,N_10336);
and U14134 (N_14134,N_10125,N_9406);
and U14135 (N_14135,N_10300,N_10269);
nor U14136 (N_14136,N_10421,N_11439);
nor U14137 (N_14137,N_9751,N_9759);
and U14138 (N_14138,N_10172,N_11297);
nor U14139 (N_14139,N_11809,N_11049);
nand U14140 (N_14140,N_11327,N_11968);
and U14141 (N_14141,N_11388,N_10465);
nor U14142 (N_14142,N_11447,N_9013);
nand U14143 (N_14143,N_10891,N_10875);
nand U14144 (N_14144,N_11357,N_11293);
nand U14145 (N_14145,N_10950,N_10327);
or U14146 (N_14146,N_11205,N_10600);
nand U14147 (N_14147,N_9834,N_10388);
nor U14148 (N_14148,N_11895,N_9600);
nor U14149 (N_14149,N_11769,N_10776);
and U14150 (N_14150,N_10605,N_10046);
and U14151 (N_14151,N_11293,N_9678);
and U14152 (N_14152,N_10200,N_9459);
nor U14153 (N_14153,N_9429,N_10435);
and U14154 (N_14154,N_11166,N_10744);
nor U14155 (N_14155,N_9894,N_10807);
or U14156 (N_14156,N_10503,N_10383);
and U14157 (N_14157,N_10537,N_9836);
or U14158 (N_14158,N_11059,N_9694);
and U14159 (N_14159,N_10413,N_9269);
or U14160 (N_14160,N_11131,N_9198);
nand U14161 (N_14161,N_10472,N_10207);
or U14162 (N_14162,N_11009,N_11097);
and U14163 (N_14163,N_11305,N_11778);
nand U14164 (N_14164,N_10708,N_11184);
nand U14165 (N_14165,N_11263,N_10678);
nor U14166 (N_14166,N_9802,N_9148);
xnor U14167 (N_14167,N_11493,N_9870);
or U14168 (N_14168,N_10955,N_9358);
or U14169 (N_14169,N_9594,N_11549);
nor U14170 (N_14170,N_11825,N_9459);
or U14171 (N_14171,N_11197,N_9508);
or U14172 (N_14172,N_10035,N_9855);
nand U14173 (N_14173,N_11135,N_10890);
and U14174 (N_14174,N_9221,N_10941);
nand U14175 (N_14175,N_9872,N_10543);
nor U14176 (N_14176,N_9627,N_10266);
or U14177 (N_14177,N_11820,N_9943);
nand U14178 (N_14178,N_11559,N_9049);
or U14179 (N_14179,N_9369,N_10779);
nor U14180 (N_14180,N_11582,N_10621);
or U14181 (N_14181,N_11203,N_9440);
nand U14182 (N_14182,N_9345,N_9771);
nor U14183 (N_14183,N_10874,N_11903);
or U14184 (N_14184,N_11182,N_10055);
and U14185 (N_14185,N_10911,N_9946);
nand U14186 (N_14186,N_10634,N_10027);
and U14187 (N_14187,N_11001,N_11817);
nor U14188 (N_14188,N_11695,N_11264);
nand U14189 (N_14189,N_10006,N_10518);
nor U14190 (N_14190,N_9612,N_9140);
nand U14191 (N_14191,N_10400,N_10955);
or U14192 (N_14192,N_9857,N_10648);
or U14193 (N_14193,N_10762,N_9373);
nand U14194 (N_14194,N_10440,N_11843);
nor U14195 (N_14195,N_9739,N_9504);
or U14196 (N_14196,N_9901,N_10939);
or U14197 (N_14197,N_10065,N_10539);
nand U14198 (N_14198,N_11483,N_10443);
or U14199 (N_14199,N_9680,N_11828);
and U14200 (N_14200,N_11354,N_10606);
and U14201 (N_14201,N_11342,N_11943);
and U14202 (N_14202,N_11252,N_9819);
and U14203 (N_14203,N_9947,N_11516);
nor U14204 (N_14204,N_9577,N_9168);
nand U14205 (N_14205,N_11861,N_9153);
and U14206 (N_14206,N_11235,N_11030);
or U14207 (N_14207,N_9850,N_10423);
nor U14208 (N_14208,N_9193,N_11907);
nand U14209 (N_14209,N_10896,N_9809);
nand U14210 (N_14210,N_11504,N_11975);
nor U14211 (N_14211,N_10887,N_9066);
nor U14212 (N_14212,N_10479,N_9290);
nand U14213 (N_14213,N_9176,N_11926);
xor U14214 (N_14214,N_9402,N_9434);
nand U14215 (N_14215,N_10678,N_10843);
nor U14216 (N_14216,N_11561,N_9609);
and U14217 (N_14217,N_11529,N_11921);
nor U14218 (N_14218,N_11556,N_10014);
nand U14219 (N_14219,N_10441,N_11643);
or U14220 (N_14220,N_10044,N_9782);
nor U14221 (N_14221,N_11907,N_11394);
nand U14222 (N_14222,N_11901,N_11978);
or U14223 (N_14223,N_11138,N_9530);
nand U14224 (N_14224,N_11808,N_9492);
and U14225 (N_14225,N_10458,N_11511);
and U14226 (N_14226,N_10379,N_10092);
or U14227 (N_14227,N_9547,N_9662);
or U14228 (N_14228,N_10601,N_10621);
nor U14229 (N_14229,N_9000,N_10895);
or U14230 (N_14230,N_11746,N_11693);
nor U14231 (N_14231,N_11593,N_11461);
nor U14232 (N_14232,N_10114,N_9362);
and U14233 (N_14233,N_9799,N_11798);
or U14234 (N_14234,N_9081,N_9448);
nor U14235 (N_14235,N_11668,N_9640);
or U14236 (N_14236,N_11781,N_9843);
and U14237 (N_14237,N_11094,N_10060);
or U14238 (N_14238,N_10121,N_9969);
nor U14239 (N_14239,N_9120,N_11581);
nand U14240 (N_14240,N_11539,N_10940);
nor U14241 (N_14241,N_11225,N_11528);
nor U14242 (N_14242,N_9347,N_11430);
or U14243 (N_14243,N_11493,N_11722);
nand U14244 (N_14244,N_9872,N_10295);
nor U14245 (N_14245,N_10491,N_9252);
or U14246 (N_14246,N_9664,N_9956);
xor U14247 (N_14247,N_11043,N_9056);
or U14248 (N_14248,N_11114,N_9195);
and U14249 (N_14249,N_9552,N_11815);
xnor U14250 (N_14250,N_11110,N_9971);
nand U14251 (N_14251,N_11672,N_9221);
or U14252 (N_14252,N_10126,N_9862);
nand U14253 (N_14253,N_11115,N_9098);
nor U14254 (N_14254,N_11105,N_9320);
nor U14255 (N_14255,N_9722,N_10058);
or U14256 (N_14256,N_9598,N_9308);
nor U14257 (N_14257,N_11867,N_10920);
nand U14258 (N_14258,N_9361,N_11791);
nor U14259 (N_14259,N_9060,N_10127);
or U14260 (N_14260,N_9607,N_9141);
or U14261 (N_14261,N_11024,N_11707);
or U14262 (N_14262,N_11778,N_9237);
or U14263 (N_14263,N_9455,N_11941);
xnor U14264 (N_14264,N_11347,N_9077);
nor U14265 (N_14265,N_11184,N_10974);
and U14266 (N_14266,N_11071,N_10884);
and U14267 (N_14267,N_11098,N_10716);
nor U14268 (N_14268,N_9455,N_9593);
nand U14269 (N_14269,N_9935,N_11442);
nor U14270 (N_14270,N_10462,N_9237);
or U14271 (N_14271,N_9321,N_9578);
or U14272 (N_14272,N_9294,N_11468);
nand U14273 (N_14273,N_10253,N_9128);
nor U14274 (N_14274,N_9869,N_11058);
and U14275 (N_14275,N_11463,N_11382);
and U14276 (N_14276,N_10589,N_10214);
or U14277 (N_14277,N_9219,N_9399);
nand U14278 (N_14278,N_10823,N_11907);
or U14279 (N_14279,N_11820,N_9693);
and U14280 (N_14280,N_10958,N_9991);
nor U14281 (N_14281,N_10242,N_11618);
and U14282 (N_14282,N_11150,N_10567);
nand U14283 (N_14283,N_9160,N_10525);
nand U14284 (N_14284,N_10923,N_11109);
nor U14285 (N_14285,N_9153,N_11681);
nor U14286 (N_14286,N_10506,N_11967);
or U14287 (N_14287,N_11892,N_10789);
or U14288 (N_14288,N_11437,N_11516);
and U14289 (N_14289,N_10744,N_10249);
or U14290 (N_14290,N_11516,N_9790);
nor U14291 (N_14291,N_9583,N_9654);
and U14292 (N_14292,N_9673,N_9761);
nor U14293 (N_14293,N_10829,N_9983);
nand U14294 (N_14294,N_9986,N_10472);
nor U14295 (N_14295,N_10764,N_10942);
or U14296 (N_14296,N_9450,N_11982);
and U14297 (N_14297,N_10357,N_10202);
and U14298 (N_14298,N_9568,N_9945);
nor U14299 (N_14299,N_9280,N_10326);
and U14300 (N_14300,N_11816,N_9053);
xnor U14301 (N_14301,N_11520,N_9280);
or U14302 (N_14302,N_9736,N_9390);
nand U14303 (N_14303,N_10610,N_11467);
and U14304 (N_14304,N_10099,N_9742);
or U14305 (N_14305,N_9112,N_10377);
nor U14306 (N_14306,N_11035,N_10695);
nor U14307 (N_14307,N_9167,N_9534);
or U14308 (N_14308,N_11957,N_9467);
nor U14309 (N_14309,N_9432,N_10638);
and U14310 (N_14310,N_9402,N_11886);
nor U14311 (N_14311,N_9097,N_10684);
nand U14312 (N_14312,N_11712,N_9584);
or U14313 (N_14313,N_10162,N_10385);
and U14314 (N_14314,N_11335,N_9595);
and U14315 (N_14315,N_10113,N_9489);
or U14316 (N_14316,N_9163,N_9990);
nor U14317 (N_14317,N_9488,N_11349);
nand U14318 (N_14318,N_10556,N_9728);
nor U14319 (N_14319,N_9535,N_11172);
or U14320 (N_14320,N_11532,N_10313);
and U14321 (N_14321,N_11276,N_10422);
nor U14322 (N_14322,N_9426,N_9039);
nor U14323 (N_14323,N_10628,N_9786);
nor U14324 (N_14324,N_11042,N_9658);
or U14325 (N_14325,N_10341,N_11999);
and U14326 (N_14326,N_9574,N_9339);
and U14327 (N_14327,N_11858,N_10374);
nand U14328 (N_14328,N_10712,N_10074);
nor U14329 (N_14329,N_11315,N_9857);
and U14330 (N_14330,N_9202,N_9299);
nor U14331 (N_14331,N_9735,N_11047);
xnor U14332 (N_14332,N_11849,N_10753);
nand U14333 (N_14333,N_10416,N_9265);
and U14334 (N_14334,N_10763,N_11400);
and U14335 (N_14335,N_11113,N_11184);
and U14336 (N_14336,N_9105,N_11065);
xor U14337 (N_14337,N_9861,N_9234);
xor U14338 (N_14338,N_10717,N_10921);
and U14339 (N_14339,N_9030,N_10829);
nor U14340 (N_14340,N_11686,N_9275);
xor U14341 (N_14341,N_11092,N_9698);
or U14342 (N_14342,N_11149,N_11719);
or U14343 (N_14343,N_9151,N_11734);
nor U14344 (N_14344,N_10518,N_10484);
nor U14345 (N_14345,N_11114,N_10622);
nand U14346 (N_14346,N_10876,N_11840);
nand U14347 (N_14347,N_9883,N_11301);
and U14348 (N_14348,N_10907,N_11909);
nor U14349 (N_14349,N_10652,N_11427);
nand U14350 (N_14350,N_10573,N_11063);
or U14351 (N_14351,N_9669,N_11310);
or U14352 (N_14352,N_9764,N_9426);
or U14353 (N_14353,N_10280,N_11365);
nor U14354 (N_14354,N_10444,N_10532);
nor U14355 (N_14355,N_11709,N_9201);
nor U14356 (N_14356,N_11873,N_9056);
and U14357 (N_14357,N_11168,N_11856);
and U14358 (N_14358,N_11113,N_11226);
nand U14359 (N_14359,N_11937,N_9771);
or U14360 (N_14360,N_10077,N_10720);
and U14361 (N_14361,N_11409,N_10448);
and U14362 (N_14362,N_11211,N_11238);
nand U14363 (N_14363,N_9376,N_10677);
nand U14364 (N_14364,N_10181,N_11338);
nand U14365 (N_14365,N_9669,N_10164);
and U14366 (N_14366,N_10520,N_9217);
and U14367 (N_14367,N_11797,N_9983);
nand U14368 (N_14368,N_11461,N_11898);
nor U14369 (N_14369,N_10740,N_10194);
nor U14370 (N_14370,N_10644,N_11138);
and U14371 (N_14371,N_10063,N_11927);
nand U14372 (N_14372,N_10364,N_11042);
and U14373 (N_14373,N_10139,N_9259);
and U14374 (N_14374,N_9598,N_11652);
nand U14375 (N_14375,N_10131,N_9828);
and U14376 (N_14376,N_9489,N_10466);
and U14377 (N_14377,N_9119,N_9044);
or U14378 (N_14378,N_10204,N_9398);
nor U14379 (N_14379,N_11021,N_10233);
or U14380 (N_14380,N_9867,N_11281);
and U14381 (N_14381,N_9034,N_11055);
or U14382 (N_14382,N_9924,N_11306);
or U14383 (N_14383,N_9072,N_11946);
and U14384 (N_14384,N_9677,N_10731);
or U14385 (N_14385,N_9836,N_10660);
or U14386 (N_14386,N_10484,N_10666);
and U14387 (N_14387,N_10589,N_9335);
nor U14388 (N_14388,N_11292,N_11191);
and U14389 (N_14389,N_11365,N_11364);
and U14390 (N_14390,N_9999,N_9921);
nand U14391 (N_14391,N_9528,N_11534);
nor U14392 (N_14392,N_11786,N_9033);
nor U14393 (N_14393,N_11316,N_9548);
or U14394 (N_14394,N_11389,N_9583);
and U14395 (N_14395,N_9420,N_10374);
and U14396 (N_14396,N_9294,N_10866);
nor U14397 (N_14397,N_10291,N_10714);
or U14398 (N_14398,N_10046,N_9858);
or U14399 (N_14399,N_9008,N_10792);
or U14400 (N_14400,N_9730,N_9633);
or U14401 (N_14401,N_10396,N_10506);
nand U14402 (N_14402,N_10296,N_9388);
nand U14403 (N_14403,N_10659,N_9466);
or U14404 (N_14404,N_11483,N_10180);
nand U14405 (N_14405,N_9125,N_9185);
nor U14406 (N_14406,N_11920,N_10925);
nor U14407 (N_14407,N_10067,N_10198);
or U14408 (N_14408,N_11748,N_10957);
nand U14409 (N_14409,N_9597,N_10510);
nand U14410 (N_14410,N_9559,N_10467);
and U14411 (N_14411,N_10438,N_11478);
nand U14412 (N_14412,N_10192,N_11841);
nand U14413 (N_14413,N_10704,N_11286);
or U14414 (N_14414,N_11507,N_11900);
nor U14415 (N_14415,N_9614,N_11927);
and U14416 (N_14416,N_10146,N_11624);
and U14417 (N_14417,N_11995,N_9516);
nand U14418 (N_14418,N_10201,N_10190);
or U14419 (N_14419,N_9546,N_11742);
or U14420 (N_14420,N_10937,N_11292);
and U14421 (N_14421,N_11993,N_9072);
nand U14422 (N_14422,N_9628,N_10951);
nand U14423 (N_14423,N_9159,N_11509);
nor U14424 (N_14424,N_10301,N_9987);
and U14425 (N_14425,N_11992,N_10095);
or U14426 (N_14426,N_9312,N_9283);
or U14427 (N_14427,N_9439,N_11966);
nor U14428 (N_14428,N_11285,N_10960);
nor U14429 (N_14429,N_11561,N_11589);
and U14430 (N_14430,N_10945,N_11921);
or U14431 (N_14431,N_11765,N_11100);
nor U14432 (N_14432,N_10474,N_11837);
nor U14433 (N_14433,N_11533,N_10072);
nor U14434 (N_14434,N_11707,N_11621);
and U14435 (N_14435,N_9121,N_11738);
nor U14436 (N_14436,N_11303,N_9826);
xnor U14437 (N_14437,N_10285,N_9813);
nand U14438 (N_14438,N_9147,N_11354);
nand U14439 (N_14439,N_10202,N_9469);
or U14440 (N_14440,N_11721,N_9899);
or U14441 (N_14441,N_9044,N_11410);
or U14442 (N_14442,N_11105,N_9366);
and U14443 (N_14443,N_10365,N_10347);
and U14444 (N_14444,N_11751,N_10151);
or U14445 (N_14445,N_11771,N_9243);
nor U14446 (N_14446,N_11072,N_10319);
nand U14447 (N_14447,N_9588,N_10529);
nand U14448 (N_14448,N_10059,N_11166);
or U14449 (N_14449,N_9910,N_10368);
or U14450 (N_14450,N_9566,N_11177);
nor U14451 (N_14451,N_10218,N_10314);
and U14452 (N_14452,N_11746,N_11259);
nand U14453 (N_14453,N_10684,N_10579);
or U14454 (N_14454,N_11272,N_9140);
nand U14455 (N_14455,N_10420,N_11346);
and U14456 (N_14456,N_10756,N_10857);
nand U14457 (N_14457,N_11255,N_10248);
nor U14458 (N_14458,N_10822,N_11123);
and U14459 (N_14459,N_10598,N_11116);
or U14460 (N_14460,N_11552,N_11231);
nor U14461 (N_14461,N_11789,N_9154);
nand U14462 (N_14462,N_10860,N_9317);
nor U14463 (N_14463,N_10060,N_11965);
or U14464 (N_14464,N_11207,N_10051);
nand U14465 (N_14465,N_9651,N_9098);
nor U14466 (N_14466,N_9325,N_11624);
nor U14467 (N_14467,N_11044,N_9234);
or U14468 (N_14468,N_9055,N_11259);
nor U14469 (N_14469,N_11378,N_9073);
nand U14470 (N_14470,N_11315,N_10715);
or U14471 (N_14471,N_11741,N_9965);
nand U14472 (N_14472,N_10409,N_10998);
and U14473 (N_14473,N_9952,N_10614);
and U14474 (N_14474,N_10069,N_9843);
nand U14475 (N_14475,N_11999,N_10116);
xor U14476 (N_14476,N_11673,N_10635);
or U14477 (N_14477,N_9928,N_11087);
and U14478 (N_14478,N_11792,N_10460);
and U14479 (N_14479,N_10005,N_9972);
or U14480 (N_14480,N_11288,N_10329);
nor U14481 (N_14481,N_11055,N_11392);
nand U14482 (N_14482,N_9875,N_10601);
nand U14483 (N_14483,N_10516,N_10457);
nand U14484 (N_14484,N_10745,N_11985);
nor U14485 (N_14485,N_10350,N_10283);
nand U14486 (N_14486,N_9637,N_9738);
and U14487 (N_14487,N_10371,N_10511);
and U14488 (N_14488,N_10528,N_11923);
nand U14489 (N_14489,N_10654,N_11959);
and U14490 (N_14490,N_11589,N_9951);
nand U14491 (N_14491,N_10448,N_11843);
or U14492 (N_14492,N_9533,N_9617);
or U14493 (N_14493,N_9290,N_9022);
nor U14494 (N_14494,N_9201,N_9127);
or U14495 (N_14495,N_9571,N_10421);
nor U14496 (N_14496,N_9808,N_10153);
nand U14497 (N_14497,N_9973,N_11344);
and U14498 (N_14498,N_9006,N_10358);
nor U14499 (N_14499,N_10000,N_11349);
nor U14500 (N_14500,N_9194,N_10510);
nor U14501 (N_14501,N_11677,N_11597);
nor U14502 (N_14502,N_11505,N_11406);
nor U14503 (N_14503,N_9792,N_9451);
and U14504 (N_14504,N_11754,N_9773);
nand U14505 (N_14505,N_9886,N_10835);
nand U14506 (N_14506,N_10093,N_11244);
nor U14507 (N_14507,N_9768,N_10781);
nor U14508 (N_14508,N_10666,N_11914);
or U14509 (N_14509,N_11542,N_11148);
and U14510 (N_14510,N_10183,N_11280);
and U14511 (N_14511,N_11713,N_11780);
nand U14512 (N_14512,N_10978,N_10750);
and U14513 (N_14513,N_9550,N_10046);
nand U14514 (N_14514,N_9491,N_9483);
and U14515 (N_14515,N_11087,N_11959);
nor U14516 (N_14516,N_10172,N_11892);
or U14517 (N_14517,N_11747,N_10058);
nor U14518 (N_14518,N_11482,N_10416);
and U14519 (N_14519,N_10493,N_10688);
or U14520 (N_14520,N_11114,N_11563);
or U14521 (N_14521,N_9768,N_9656);
nor U14522 (N_14522,N_9714,N_10932);
or U14523 (N_14523,N_11802,N_10116);
nand U14524 (N_14524,N_11487,N_9120);
or U14525 (N_14525,N_9113,N_10688);
and U14526 (N_14526,N_10435,N_11661);
nand U14527 (N_14527,N_10523,N_10991);
nand U14528 (N_14528,N_11696,N_9014);
and U14529 (N_14529,N_11773,N_11953);
and U14530 (N_14530,N_10414,N_10521);
nand U14531 (N_14531,N_10752,N_11032);
nor U14532 (N_14532,N_11736,N_10729);
and U14533 (N_14533,N_11328,N_10413);
nor U14534 (N_14534,N_10013,N_11110);
nor U14535 (N_14535,N_10424,N_10309);
and U14536 (N_14536,N_10799,N_9132);
nand U14537 (N_14537,N_10490,N_11557);
and U14538 (N_14538,N_9178,N_11846);
nand U14539 (N_14539,N_9448,N_9607);
nor U14540 (N_14540,N_11004,N_10850);
nor U14541 (N_14541,N_11241,N_9324);
nor U14542 (N_14542,N_11976,N_10602);
or U14543 (N_14543,N_10291,N_9990);
and U14544 (N_14544,N_11968,N_10450);
and U14545 (N_14545,N_11435,N_9010);
and U14546 (N_14546,N_11271,N_11122);
and U14547 (N_14547,N_10819,N_9424);
and U14548 (N_14548,N_11310,N_9676);
or U14549 (N_14549,N_10271,N_11034);
nor U14550 (N_14550,N_11954,N_11555);
nor U14551 (N_14551,N_11636,N_11525);
nor U14552 (N_14552,N_11127,N_9659);
nand U14553 (N_14553,N_11651,N_11041);
and U14554 (N_14554,N_11448,N_10225);
nor U14555 (N_14555,N_10492,N_11049);
nor U14556 (N_14556,N_10207,N_9140);
nor U14557 (N_14557,N_10683,N_10454);
or U14558 (N_14558,N_10867,N_10346);
nor U14559 (N_14559,N_9389,N_11163);
nand U14560 (N_14560,N_9375,N_11404);
xnor U14561 (N_14561,N_9378,N_11909);
and U14562 (N_14562,N_10427,N_11072);
xnor U14563 (N_14563,N_10320,N_10022);
or U14564 (N_14564,N_11231,N_11095);
nor U14565 (N_14565,N_11286,N_10928);
xnor U14566 (N_14566,N_11645,N_11687);
nor U14567 (N_14567,N_10378,N_11453);
or U14568 (N_14568,N_11675,N_11558);
or U14569 (N_14569,N_11100,N_9883);
and U14570 (N_14570,N_11806,N_10994);
nor U14571 (N_14571,N_10843,N_10975);
and U14572 (N_14572,N_9736,N_9459);
nand U14573 (N_14573,N_11621,N_9048);
and U14574 (N_14574,N_11388,N_11483);
nand U14575 (N_14575,N_9968,N_10419);
or U14576 (N_14576,N_10328,N_9303);
nand U14577 (N_14577,N_9799,N_11406);
or U14578 (N_14578,N_9023,N_9191);
and U14579 (N_14579,N_11322,N_11331);
nand U14580 (N_14580,N_11805,N_9369);
and U14581 (N_14581,N_9699,N_11982);
or U14582 (N_14582,N_10277,N_9314);
and U14583 (N_14583,N_11136,N_10722);
or U14584 (N_14584,N_10565,N_10146);
nand U14585 (N_14585,N_10680,N_11283);
or U14586 (N_14586,N_9016,N_9138);
and U14587 (N_14587,N_9583,N_10345);
nor U14588 (N_14588,N_9375,N_9535);
nor U14589 (N_14589,N_9842,N_9895);
nor U14590 (N_14590,N_11458,N_10099);
or U14591 (N_14591,N_10968,N_10679);
or U14592 (N_14592,N_10101,N_11173);
nor U14593 (N_14593,N_10184,N_10235);
and U14594 (N_14594,N_11397,N_9111);
and U14595 (N_14595,N_9528,N_11741);
nand U14596 (N_14596,N_11564,N_10007);
and U14597 (N_14597,N_9035,N_10145);
or U14598 (N_14598,N_11333,N_9046);
nand U14599 (N_14599,N_11622,N_11326);
or U14600 (N_14600,N_11199,N_10327);
and U14601 (N_14601,N_10610,N_10079);
nand U14602 (N_14602,N_9635,N_11548);
or U14603 (N_14603,N_10105,N_9422);
and U14604 (N_14604,N_10863,N_9392);
nor U14605 (N_14605,N_10527,N_10463);
nor U14606 (N_14606,N_10325,N_10125);
or U14607 (N_14607,N_10948,N_10568);
or U14608 (N_14608,N_9387,N_9517);
and U14609 (N_14609,N_10068,N_10419);
nand U14610 (N_14610,N_11224,N_9464);
nor U14611 (N_14611,N_9991,N_10669);
or U14612 (N_14612,N_10372,N_10544);
nand U14613 (N_14613,N_11287,N_10216);
or U14614 (N_14614,N_10377,N_10302);
nor U14615 (N_14615,N_11000,N_9794);
nor U14616 (N_14616,N_11826,N_9841);
and U14617 (N_14617,N_9282,N_9030);
and U14618 (N_14618,N_10127,N_11139);
nor U14619 (N_14619,N_11146,N_10568);
nand U14620 (N_14620,N_11745,N_10870);
or U14621 (N_14621,N_9230,N_10928);
nor U14622 (N_14622,N_10632,N_11680);
nand U14623 (N_14623,N_9807,N_9635);
and U14624 (N_14624,N_10874,N_10391);
or U14625 (N_14625,N_9416,N_11496);
nand U14626 (N_14626,N_11401,N_10817);
or U14627 (N_14627,N_9555,N_10818);
nor U14628 (N_14628,N_11823,N_11928);
and U14629 (N_14629,N_9593,N_11542);
and U14630 (N_14630,N_10726,N_9825);
and U14631 (N_14631,N_11552,N_9427);
nand U14632 (N_14632,N_11667,N_10983);
nand U14633 (N_14633,N_9590,N_11992);
nor U14634 (N_14634,N_9761,N_10578);
nand U14635 (N_14635,N_9955,N_11857);
nor U14636 (N_14636,N_9118,N_11990);
and U14637 (N_14637,N_10174,N_10276);
nand U14638 (N_14638,N_11770,N_11633);
nand U14639 (N_14639,N_9269,N_11256);
nor U14640 (N_14640,N_9242,N_9058);
nor U14641 (N_14641,N_9087,N_10608);
nor U14642 (N_14642,N_9559,N_9585);
nand U14643 (N_14643,N_11219,N_9888);
and U14644 (N_14644,N_9846,N_9401);
nand U14645 (N_14645,N_10896,N_11069);
or U14646 (N_14646,N_9957,N_9091);
nand U14647 (N_14647,N_9695,N_10209);
nor U14648 (N_14648,N_11959,N_10899);
or U14649 (N_14649,N_11372,N_9386);
xor U14650 (N_14650,N_10680,N_10082);
nand U14651 (N_14651,N_10881,N_9006);
and U14652 (N_14652,N_11633,N_11738);
nor U14653 (N_14653,N_11005,N_10333);
or U14654 (N_14654,N_10132,N_10015);
and U14655 (N_14655,N_11741,N_10371);
and U14656 (N_14656,N_9701,N_10674);
or U14657 (N_14657,N_11841,N_11270);
nor U14658 (N_14658,N_10078,N_9581);
and U14659 (N_14659,N_10490,N_11135);
and U14660 (N_14660,N_9107,N_9043);
or U14661 (N_14661,N_11747,N_9350);
nor U14662 (N_14662,N_11252,N_9749);
and U14663 (N_14663,N_10624,N_11761);
or U14664 (N_14664,N_11684,N_11127);
and U14665 (N_14665,N_11750,N_11141);
and U14666 (N_14666,N_11369,N_11484);
nand U14667 (N_14667,N_10390,N_10662);
or U14668 (N_14668,N_11957,N_9753);
nor U14669 (N_14669,N_10501,N_10585);
nand U14670 (N_14670,N_9701,N_10976);
nand U14671 (N_14671,N_9550,N_11634);
nand U14672 (N_14672,N_11562,N_11849);
and U14673 (N_14673,N_10977,N_9385);
xnor U14674 (N_14674,N_11403,N_10538);
nand U14675 (N_14675,N_9642,N_11284);
or U14676 (N_14676,N_10869,N_9049);
and U14677 (N_14677,N_11306,N_9421);
or U14678 (N_14678,N_9821,N_9230);
nor U14679 (N_14679,N_10290,N_9058);
nand U14680 (N_14680,N_9878,N_11554);
or U14681 (N_14681,N_11369,N_11522);
nor U14682 (N_14682,N_10921,N_11549);
nor U14683 (N_14683,N_9040,N_11614);
and U14684 (N_14684,N_9806,N_11156);
xnor U14685 (N_14685,N_9257,N_11885);
and U14686 (N_14686,N_11435,N_10373);
and U14687 (N_14687,N_9480,N_9342);
nand U14688 (N_14688,N_11136,N_9638);
nor U14689 (N_14689,N_9438,N_11773);
nor U14690 (N_14690,N_9139,N_11343);
nand U14691 (N_14691,N_10763,N_11612);
nand U14692 (N_14692,N_9069,N_10629);
and U14693 (N_14693,N_10375,N_10760);
nor U14694 (N_14694,N_9463,N_10939);
or U14695 (N_14695,N_11160,N_11741);
and U14696 (N_14696,N_9947,N_11097);
nor U14697 (N_14697,N_10497,N_11856);
nor U14698 (N_14698,N_9137,N_11843);
and U14699 (N_14699,N_10562,N_10979);
or U14700 (N_14700,N_9009,N_10263);
nor U14701 (N_14701,N_10590,N_9854);
and U14702 (N_14702,N_11098,N_11344);
nor U14703 (N_14703,N_9982,N_11093);
and U14704 (N_14704,N_9677,N_9039);
xor U14705 (N_14705,N_11167,N_11068);
and U14706 (N_14706,N_11602,N_10118);
nor U14707 (N_14707,N_11225,N_11837);
nor U14708 (N_14708,N_11336,N_10894);
or U14709 (N_14709,N_10118,N_11545);
and U14710 (N_14710,N_9061,N_10966);
and U14711 (N_14711,N_11239,N_9623);
or U14712 (N_14712,N_10822,N_11763);
and U14713 (N_14713,N_9007,N_9806);
and U14714 (N_14714,N_11730,N_9010);
nand U14715 (N_14715,N_10461,N_10128);
nor U14716 (N_14716,N_9428,N_11611);
nor U14717 (N_14717,N_9405,N_10691);
and U14718 (N_14718,N_11542,N_11152);
and U14719 (N_14719,N_10237,N_11764);
nand U14720 (N_14720,N_9481,N_9801);
and U14721 (N_14721,N_9795,N_9902);
nand U14722 (N_14722,N_11943,N_9826);
nor U14723 (N_14723,N_10568,N_9637);
nor U14724 (N_14724,N_11643,N_11895);
nor U14725 (N_14725,N_11171,N_10565);
nand U14726 (N_14726,N_11798,N_10214);
nand U14727 (N_14727,N_10982,N_9905);
or U14728 (N_14728,N_11272,N_11531);
nand U14729 (N_14729,N_10668,N_9858);
or U14730 (N_14730,N_9664,N_11149);
nand U14731 (N_14731,N_9816,N_11369);
or U14732 (N_14732,N_10343,N_9387);
nor U14733 (N_14733,N_10518,N_9087);
nor U14734 (N_14734,N_10467,N_9678);
xor U14735 (N_14735,N_10659,N_10726);
nor U14736 (N_14736,N_11733,N_10646);
and U14737 (N_14737,N_11790,N_9299);
nand U14738 (N_14738,N_11406,N_10802);
or U14739 (N_14739,N_11817,N_11039);
nor U14740 (N_14740,N_11582,N_9109);
or U14741 (N_14741,N_11803,N_10721);
or U14742 (N_14742,N_11883,N_10570);
or U14743 (N_14743,N_9800,N_11671);
nor U14744 (N_14744,N_11690,N_10876);
nand U14745 (N_14745,N_11985,N_11260);
nor U14746 (N_14746,N_10454,N_9700);
nand U14747 (N_14747,N_11922,N_10873);
xnor U14748 (N_14748,N_11263,N_10602);
nor U14749 (N_14749,N_11633,N_11397);
or U14750 (N_14750,N_11589,N_9826);
or U14751 (N_14751,N_11198,N_9016);
nand U14752 (N_14752,N_10921,N_9121);
or U14753 (N_14753,N_10157,N_11406);
and U14754 (N_14754,N_11756,N_11716);
and U14755 (N_14755,N_9958,N_11584);
or U14756 (N_14756,N_11270,N_10888);
nor U14757 (N_14757,N_11819,N_9267);
and U14758 (N_14758,N_11999,N_9077);
and U14759 (N_14759,N_11137,N_10540);
nand U14760 (N_14760,N_11558,N_11505);
nor U14761 (N_14761,N_10766,N_11769);
nand U14762 (N_14762,N_9255,N_9298);
or U14763 (N_14763,N_9529,N_9278);
or U14764 (N_14764,N_11497,N_11601);
and U14765 (N_14765,N_10097,N_9677);
nand U14766 (N_14766,N_11441,N_11218);
nor U14767 (N_14767,N_10396,N_11669);
or U14768 (N_14768,N_11620,N_11613);
and U14769 (N_14769,N_10747,N_10623);
nand U14770 (N_14770,N_9932,N_11354);
or U14771 (N_14771,N_11532,N_9855);
and U14772 (N_14772,N_10443,N_10631);
and U14773 (N_14773,N_9207,N_11662);
or U14774 (N_14774,N_10452,N_11716);
xor U14775 (N_14775,N_11636,N_10230);
or U14776 (N_14776,N_9118,N_10387);
or U14777 (N_14777,N_9860,N_9949);
or U14778 (N_14778,N_11950,N_9032);
nand U14779 (N_14779,N_9299,N_10987);
or U14780 (N_14780,N_9167,N_10176);
or U14781 (N_14781,N_10477,N_9510);
nand U14782 (N_14782,N_10357,N_9538);
or U14783 (N_14783,N_11253,N_10269);
nor U14784 (N_14784,N_10381,N_9923);
nor U14785 (N_14785,N_11871,N_11268);
nor U14786 (N_14786,N_11339,N_10658);
or U14787 (N_14787,N_10957,N_11308);
and U14788 (N_14788,N_11211,N_11409);
and U14789 (N_14789,N_9625,N_11133);
nand U14790 (N_14790,N_10194,N_9076);
nor U14791 (N_14791,N_11827,N_10416);
nor U14792 (N_14792,N_11630,N_9177);
nor U14793 (N_14793,N_9242,N_11892);
nor U14794 (N_14794,N_10925,N_11654);
nand U14795 (N_14795,N_9180,N_9764);
or U14796 (N_14796,N_10852,N_11021);
or U14797 (N_14797,N_10991,N_10872);
nand U14798 (N_14798,N_11881,N_11028);
nand U14799 (N_14799,N_11624,N_9533);
or U14800 (N_14800,N_11325,N_11082);
nand U14801 (N_14801,N_10500,N_10425);
and U14802 (N_14802,N_9391,N_9853);
nor U14803 (N_14803,N_11801,N_9416);
or U14804 (N_14804,N_10067,N_9337);
nor U14805 (N_14805,N_10817,N_10197);
and U14806 (N_14806,N_9116,N_10529);
and U14807 (N_14807,N_9667,N_11642);
nand U14808 (N_14808,N_11108,N_11934);
nand U14809 (N_14809,N_10272,N_9881);
nor U14810 (N_14810,N_9005,N_9900);
nand U14811 (N_14811,N_11561,N_10362);
and U14812 (N_14812,N_9492,N_11847);
and U14813 (N_14813,N_11903,N_9368);
nor U14814 (N_14814,N_10913,N_9533);
or U14815 (N_14815,N_10770,N_9118);
nor U14816 (N_14816,N_9737,N_10634);
or U14817 (N_14817,N_11448,N_10617);
or U14818 (N_14818,N_10635,N_11356);
and U14819 (N_14819,N_11775,N_9174);
nor U14820 (N_14820,N_10184,N_9370);
or U14821 (N_14821,N_11278,N_9586);
and U14822 (N_14822,N_11601,N_11349);
or U14823 (N_14823,N_11581,N_10101);
nand U14824 (N_14824,N_10946,N_9246);
nand U14825 (N_14825,N_10174,N_10738);
xnor U14826 (N_14826,N_10265,N_11830);
or U14827 (N_14827,N_9034,N_11016);
or U14828 (N_14828,N_9732,N_11785);
nand U14829 (N_14829,N_11735,N_11950);
or U14830 (N_14830,N_11710,N_11691);
nor U14831 (N_14831,N_10071,N_10574);
nand U14832 (N_14832,N_11916,N_11376);
nand U14833 (N_14833,N_10895,N_11449);
nor U14834 (N_14834,N_9095,N_9312);
nand U14835 (N_14835,N_11979,N_9325);
or U14836 (N_14836,N_10058,N_10439);
or U14837 (N_14837,N_11403,N_11822);
xor U14838 (N_14838,N_10012,N_10345);
or U14839 (N_14839,N_11651,N_9348);
or U14840 (N_14840,N_9891,N_9373);
and U14841 (N_14841,N_10511,N_11464);
nor U14842 (N_14842,N_9864,N_9236);
nand U14843 (N_14843,N_10319,N_10354);
nand U14844 (N_14844,N_10841,N_10872);
and U14845 (N_14845,N_10671,N_11987);
or U14846 (N_14846,N_11412,N_11719);
or U14847 (N_14847,N_9366,N_10467);
nand U14848 (N_14848,N_10335,N_10103);
nor U14849 (N_14849,N_9875,N_9027);
nand U14850 (N_14850,N_11704,N_10600);
and U14851 (N_14851,N_11462,N_11108);
and U14852 (N_14852,N_9408,N_10409);
or U14853 (N_14853,N_10663,N_10066);
nand U14854 (N_14854,N_11162,N_10445);
nand U14855 (N_14855,N_9380,N_10906);
nor U14856 (N_14856,N_11711,N_11537);
nor U14857 (N_14857,N_10139,N_10245);
and U14858 (N_14858,N_11957,N_10975);
and U14859 (N_14859,N_9130,N_11694);
or U14860 (N_14860,N_10364,N_11847);
or U14861 (N_14861,N_10442,N_10907);
or U14862 (N_14862,N_10348,N_10319);
nor U14863 (N_14863,N_10035,N_10790);
nor U14864 (N_14864,N_11511,N_9222);
and U14865 (N_14865,N_9027,N_10927);
nand U14866 (N_14866,N_11630,N_9540);
and U14867 (N_14867,N_11434,N_11800);
nand U14868 (N_14868,N_11362,N_11496);
nor U14869 (N_14869,N_9908,N_11568);
nand U14870 (N_14870,N_11698,N_9393);
nand U14871 (N_14871,N_10620,N_9636);
and U14872 (N_14872,N_10694,N_11374);
nor U14873 (N_14873,N_11804,N_9531);
nand U14874 (N_14874,N_10765,N_10426);
nand U14875 (N_14875,N_9602,N_10818);
and U14876 (N_14876,N_10790,N_10689);
nor U14877 (N_14877,N_9871,N_11568);
nand U14878 (N_14878,N_11860,N_9947);
and U14879 (N_14879,N_10718,N_9468);
and U14880 (N_14880,N_10945,N_10160);
and U14881 (N_14881,N_10582,N_10750);
nand U14882 (N_14882,N_11583,N_10285);
nand U14883 (N_14883,N_11970,N_9014);
and U14884 (N_14884,N_9561,N_11413);
nor U14885 (N_14885,N_9314,N_11821);
nor U14886 (N_14886,N_9271,N_11790);
and U14887 (N_14887,N_11061,N_9183);
nand U14888 (N_14888,N_10792,N_11907);
and U14889 (N_14889,N_10197,N_10902);
or U14890 (N_14890,N_9406,N_9388);
and U14891 (N_14891,N_11195,N_10340);
and U14892 (N_14892,N_9637,N_11609);
and U14893 (N_14893,N_9958,N_9917);
nand U14894 (N_14894,N_11139,N_10056);
or U14895 (N_14895,N_10729,N_9942);
nand U14896 (N_14896,N_10123,N_10218);
and U14897 (N_14897,N_11085,N_11160);
or U14898 (N_14898,N_9938,N_9543);
nand U14899 (N_14899,N_11488,N_11150);
nand U14900 (N_14900,N_11484,N_9090);
nand U14901 (N_14901,N_10719,N_11819);
nand U14902 (N_14902,N_10426,N_10586);
and U14903 (N_14903,N_10065,N_11987);
or U14904 (N_14904,N_10454,N_10338);
nor U14905 (N_14905,N_9119,N_10040);
or U14906 (N_14906,N_10473,N_10109);
nor U14907 (N_14907,N_10713,N_10923);
or U14908 (N_14908,N_9969,N_11677);
or U14909 (N_14909,N_9759,N_11792);
and U14910 (N_14910,N_10683,N_10993);
xor U14911 (N_14911,N_9319,N_9096);
nand U14912 (N_14912,N_10804,N_10359);
or U14913 (N_14913,N_11744,N_10683);
nand U14914 (N_14914,N_9937,N_10471);
nand U14915 (N_14915,N_10917,N_11950);
and U14916 (N_14916,N_9474,N_10101);
nand U14917 (N_14917,N_10084,N_9551);
nand U14918 (N_14918,N_9883,N_11084);
and U14919 (N_14919,N_10754,N_10504);
nand U14920 (N_14920,N_10035,N_10558);
and U14921 (N_14921,N_10373,N_10399);
nor U14922 (N_14922,N_9546,N_10562);
and U14923 (N_14923,N_10541,N_9583);
or U14924 (N_14924,N_11015,N_11201);
nor U14925 (N_14925,N_10040,N_10857);
and U14926 (N_14926,N_11658,N_9992);
and U14927 (N_14927,N_11429,N_11028);
nand U14928 (N_14928,N_9954,N_10622);
or U14929 (N_14929,N_9847,N_9158);
or U14930 (N_14930,N_10891,N_11445);
and U14931 (N_14931,N_11072,N_9996);
nand U14932 (N_14932,N_10169,N_11826);
nor U14933 (N_14933,N_10231,N_10758);
nand U14934 (N_14934,N_9901,N_10313);
and U14935 (N_14935,N_10385,N_9698);
nor U14936 (N_14936,N_9292,N_10917);
nand U14937 (N_14937,N_11243,N_9498);
or U14938 (N_14938,N_11688,N_10592);
or U14939 (N_14939,N_11735,N_11643);
nor U14940 (N_14940,N_9334,N_9374);
and U14941 (N_14941,N_10494,N_10264);
xor U14942 (N_14942,N_9607,N_11831);
nand U14943 (N_14943,N_10185,N_11073);
and U14944 (N_14944,N_11112,N_10033);
and U14945 (N_14945,N_10374,N_10609);
or U14946 (N_14946,N_10993,N_10544);
nor U14947 (N_14947,N_11912,N_11966);
nor U14948 (N_14948,N_9559,N_10034);
nor U14949 (N_14949,N_9057,N_11682);
nand U14950 (N_14950,N_10027,N_9747);
nor U14951 (N_14951,N_11230,N_11701);
and U14952 (N_14952,N_9198,N_10233);
nor U14953 (N_14953,N_11397,N_10167);
or U14954 (N_14954,N_11198,N_10481);
and U14955 (N_14955,N_9515,N_11715);
nand U14956 (N_14956,N_11450,N_9203);
nand U14957 (N_14957,N_10616,N_10875);
or U14958 (N_14958,N_10617,N_11783);
nor U14959 (N_14959,N_10495,N_11179);
or U14960 (N_14960,N_9341,N_11312);
nand U14961 (N_14961,N_9020,N_11128);
and U14962 (N_14962,N_11983,N_9949);
or U14963 (N_14963,N_9653,N_10549);
nand U14964 (N_14964,N_11328,N_11751);
and U14965 (N_14965,N_9458,N_11763);
or U14966 (N_14966,N_9919,N_10359);
nand U14967 (N_14967,N_11406,N_10911);
and U14968 (N_14968,N_11258,N_10668);
nor U14969 (N_14969,N_11106,N_11631);
and U14970 (N_14970,N_9488,N_11510);
nor U14971 (N_14971,N_9520,N_11527);
nand U14972 (N_14972,N_11481,N_11068);
and U14973 (N_14973,N_9160,N_10978);
nand U14974 (N_14974,N_9116,N_10283);
and U14975 (N_14975,N_9092,N_11945);
nor U14976 (N_14976,N_10002,N_11402);
or U14977 (N_14977,N_11473,N_9135);
nor U14978 (N_14978,N_10552,N_11699);
nor U14979 (N_14979,N_11553,N_11815);
nor U14980 (N_14980,N_11736,N_11053);
nor U14981 (N_14981,N_10354,N_10078);
and U14982 (N_14982,N_11510,N_9533);
and U14983 (N_14983,N_11307,N_10425);
xor U14984 (N_14984,N_10097,N_10415);
xnor U14985 (N_14985,N_10259,N_9169);
and U14986 (N_14986,N_11966,N_10690);
nand U14987 (N_14987,N_10127,N_9678);
nand U14988 (N_14988,N_10284,N_11019);
nor U14989 (N_14989,N_10272,N_9628);
nor U14990 (N_14990,N_11927,N_10605);
or U14991 (N_14991,N_9729,N_11881);
or U14992 (N_14992,N_9227,N_10044);
or U14993 (N_14993,N_10617,N_9720);
nor U14994 (N_14994,N_9863,N_11755);
and U14995 (N_14995,N_9835,N_11532);
or U14996 (N_14996,N_11254,N_9730);
nor U14997 (N_14997,N_11849,N_9817);
nand U14998 (N_14998,N_10928,N_9452);
nor U14999 (N_14999,N_10712,N_11218);
and UO_0 (O_0,N_13531,N_13502);
nand UO_1 (O_1,N_12710,N_14457);
nand UO_2 (O_2,N_14598,N_13981);
nand UO_3 (O_3,N_12397,N_13869);
nand UO_4 (O_4,N_13999,N_12265);
and UO_5 (O_5,N_12105,N_13404);
nand UO_6 (O_6,N_14699,N_13949);
nand UO_7 (O_7,N_14201,N_12109);
nor UO_8 (O_8,N_14348,N_12232);
or UO_9 (O_9,N_14291,N_13405);
nand UO_10 (O_10,N_14051,N_12590);
nand UO_11 (O_11,N_12243,N_14825);
and UO_12 (O_12,N_12474,N_12306);
or UO_13 (O_13,N_14976,N_13825);
nand UO_14 (O_14,N_12159,N_13448);
and UO_15 (O_15,N_12624,N_13560);
or UO_16 (O_16,N_12227,N_12356);
nor UO_17 (O_17,N_13051,N_13879);
nor UO_18 (O_18,N_12438,N_13896);
and UO_19 (O_19,N_14687,N_14685);
xor UO_20 (O_20,N_13602,N_12766);
or UO_21 (O_21,N_14220,N_14127);
or UO_22 (O_22,N_13307,N_13222);
nand UO_23 (O_23,N_13342,N_14152);
nand UO_24 (O_24,N_13826,N_13056);
nand UO_25 (O_25,N_13696,N_14069);
xnor UO_26 (O_26,N_12118,N_14091);
nand UO_27 (O_27,N_14904,N_12421);
or UO_28 (O_28,N_14740,N_13295);
nor UO_29 (O_29,N_12389,N_12514);
nand UO_30 (O_30,N_13365,N_12807);
xnor UO_31 (O_31,N_12504,N_12603);
or UO_32 (O_32,N_12130,N_12772);
and UO_33 (O_33,N_12354,N_13645);
and UO_34 (O_34,N_13532,N_14301);
and UO_35 (O_35,N_12775,N_14359);
nand UO_36 (O_36,N_12900,N_12281);
nand UO_37 (O_37,N_12594,N_13475);
nand UO_38 (O_38,N_14979,N_12789);
or UO_39 (O_39,N_14721,N_13741);
nand UO_40 (O_40,N_12406,N_12086);
nand UO_41 (O_41,N_14345,N_12932);
nand UO_42 (O_42,N_13478,N_14112);
nor UO_43 (O_43,N_13422,N_13918);
nor UO_44 (O_44,N_13193,N_14946);
and UO_45 (O_45,N_12595,N_13830);
nand UO_46 (O_46,N_14562,N_14060);
nor UO_47 (O_47,N_14443,N_13732);
or UO_48 (O_48,N_13855,N_12025);
or UO_49 (O_49,N_14128,N_13940);
and UO_50 (O_50,N_13240,N_12926);
and UO_51 (O_51,N_13761,N_14821);
and UO_52 (O_52,N_14912,N_14219);
and UO_53 (O_53,N_12097,N_13287);
nand UO_54 (O_54,N_13873,N_12705);
or UO_55 (O_55,N_12393,N_14545);
or UO_56 (O_56,N_13921,N_12158);
or UO_57 (O_57,N_14894,N_13088);
and UO_58 (O_58,N_12058,N_13194);
nand UO_59 (O_59,N_14185,N_13627);
xor UO_60 (O_60,N_12920,N_12446);
nand UO_61 (O_61,N_13774,N_12587);
or UO_62 (O_62,N_14897,N_13523);
or UO_63 (O_63,N_13119,N_14939);
nand UO_64 (O_64,N_14196,N_12852);
nand UO_65 (O_65,N_13450,N_13902);
nor UO_66 (O_66,N_12656,N_12103);
nand UO_67 (O_67,N_13655,N_12170);
nand UO_68 (O_68,N_12890,N_14563);
or UO_69 (O_69,N_14993,N_12480);
nor UO_70 (O_70,N_14115,N_12795);
and UO_71 (O_71,N_14782,N_12568);
or UO_72 (O_72,N_14949,N_13614);
nand UO_73 (O_73,N_13571,N_14271);
nand UO_74 (O_74,N_14144,N_13785);
nor UO_75 (O_75,N_14674,N_12867);
and UO_76 (O_76,N_12950,N_13149);
nor UO_77 (O_77,N_13617,N_13250);
xnor UO_78 (O_78,N_13148,N_14851);
or UO_79 (O_79,N_12378,N_14458);
nor UO_80 (O_80,N_13062,N_14257);
and UO_81 (O_81,N_13700,N_12748);
and UO_82 (O_82,N_14288,N_13917);
and UO_83 (O_83,N_13214,N_12847);
nand UO_84 (O_84,N_13884,N_14722);
nor UO_85 (O_85,N_14159,N_14354);
and UO_86 (O_86,N_14202,N_13800);
or UO_87 (O_87,N_12813,N_13990);
and UO_88 (O_88,N_12558,N_12889);
nand UO_89 (O_89,N_12304,N_12197);
xor UO_90 (O_90,N_13901,N_13457);
and UO_91 (O_91,N_12543,N_13637);
and UO_92 (O_92,N_14815,N_12317);
and UO_93 (O_93,N_12429,N_13485);
nor UO_94 (O_94,N_12075,N_13745);
or UO_95 (O_95,N_12314,N_14497);
nand UO_96 (O_96,N_12173,N_13216);
nor UO_97 (O_97,N_14566,N_12200);
nand UO_98 (O_98,N_14819,N_13041);
or UO_99 (O_99,N_14072,N_14396);
xnor UO_100 (O_100,N_14372,N_14393);
xor UO_101 (O_101,N_13052,N_14567);
and UO_102 (O_102,N_12231,N_12277);
and UO_103 (O_103,N_12776,N_13244);
nor UO_104 (O_104,N_14436,N_13187);
or UO_105 (O_105,N_12387,N_13043);
nor UO_106 (O_106,N_14863,N_13408);
or UO_107 (O_107,N_14120,N_14840);
nand UO_108 (O_108,N_12946,N_14056);
or UO_109 (O_109,N_13402,N_12468);
and UO_110 (O_110,N_13663,N_13456);
or UO_111 (O_111,N_13740,N_12141);
or UO_112 (O_112,N_13013,N_12817);
nand UO_113 (O_113,N_12648,N_12757);
or UO_114 (O_114,N_14356,N_13492);
nor UO_115 (O_115,N_14285,N_13958);
and UO_116 (O_116,N_12997,N_12038);
or UO_117 (O_117,N_14216,N_13762);
nand UO_118 (O_118,N_13874,N_14337);
nor UO_119 (O_119,N_14872,N_14045);
xnor UO_120 (O_120,N_13097,N_13372);
nor UO_121 (O_121,N_13561,N_12207);
or UO_122 (O_122,N_12791,N_14832);
and UO_123 (O_123,N_13181,N_12691);
or UO_124 (O_124,N_12916,N_12567);
nor UO_125 (O_125,N_14125,N_13369);
nor UO_126 (O_126,N_13131,N_12608);
nand UO_127 (O_127,N_14113,N_13929);
nand UO_128 (O_128,N_12683,N_13754);
nand UO_129 (O_129,N_12961,N_14690);
and UO_130 (O_130,N_14384,N_14542);
or UO_131 (O_131,N_12576,N_12477);
or UO_132 (O_132,N_14004,N_14631);
xor UO_133 (O_133,N_12904,N_13154);
nand UO_134 (O_134,N_13652,N_13567);
nand UO_135 (O_135,N_12614,N_14119);
xnor UO_136 (O_136,N_14943,N_13195);
and UO_137 (O_137,N_12879,N_12280);
and UO_138 (O_138,N_14561,N_12257);
or UO_139 (O_139,N_12760,N_12827);
nand UO_140 (O_140,N_12746,N_14106);
and UO_141 (O_141,N_13789,N_12942);
nor UO_142 (O_142,N_14244,N_14247);
and UO_143 (O_143,N_13775,N_13517);
nand UO_144 (O_144,N_12484,N_12230);
nor UO_145 (O_145,N_13474,N_13458);
nand UO_146 (O_146,N_12975,N_13207);
nand UO_147 (O_147,N_12466,N_13590);
or UO_148 (O_148,N_12095,N_13853);
nand UO_149 (O_149,N_14734,N_12859);
nand UO_150 (O_150,N_13178,N_14491);
nand UO_151 (O_151,N_13246,N_13773);
and UO_152 (O_152,N_12600,N_13234);
nor UO_153 (O_153,N_14030,N_13199);
and UO_154 (O_154,N_12869,N_12687);
nand UO_155 (O_155,N_14837,N_13280);
nor UO_156 (O_156,N_13599,N_13054);
and UO_157 (O_157,N_13329,N_14657);
nand UO_158 (O_158,N_12810,N_13160);
nand UO_159 (O_159,N_13805,N_12270);
nand UO_160 (O_160,N_14710,N_13048);
nor UO_161 (O_161,N_12897,N_12903);
xor UO_162 (O_162,N_12353,N_13488);
or UO_163 (O_163,N_13138,N_14527);
or UO_164 (O_164,N_12470,N_12360);
and UO_165 (O_165,N_12625,N_12008);
nor UO_166 (O_166,N_14813,N_12617);
or UO_167 (O_167,N_13336,N_14223);
nor UO_168 (O_168,N_13758,N_14370);
nand UO_169 (O_169,N_12166,N_13339);
nand UO_170 (O_170,N_12552,N_13955);
nor UO_171 (O_171,N_14558,N_12915);
nand UO_172 (O_172,N_12398,N_13166);
nor UO_173 (O_173,N_13049,N_14360);
nand UO_174 (O_174,N_13114,N_14531);
or UO_175 (O_175,N_12137,N_12195);
nor UO_176 (O_176,N_12053,N_13586);
and UO_177 (O_177,N_14237,N_14585);
and UO_178 (O_178,N_12366,N_14937);
nor UO_179 (O_179,N_12606,N_13379);
nor UO_180 (O_180,N_12156,N_13911);
or UO_181 (O_181,N_14541,N_12924);
or UO_182 (O_182,N_13093,N_12189);
nor UO_183 (O_183,N_14015,N_13155);
xor UO_184 (O_184,N_14958,N_12411);
and UO_185 (O_185,N_14422,N_13084);
or UO_186 (O_186,N_12161,N_12163);
nand UO_187 (O_187,N_14555,N_12634);
nand UO_188 (O_188,N_13993,N_12068);
and UO_189 (O_189,N_12702,N_12806);
nor UO_190 (O_190,N_13351,N_14686);
and UO_191 (O_191,N_14640,N_14700);
or UO_192 (O_192,N_14807,N_14811);
xor UO_193 (O_193,N_13931,N_12071);
nand UO_194 (O_194,N_12093,N_14586);
and UO_195 (O_195,N_14974,N_12826);
and UO_196 (O_196,N_14834,N_13197);
and UO_197 (O_197,N_12209,N_14100);
or UO_198 (O_198,N_12001,N_13248);
nand UO_199 (O_199,N_13833,N_14252);
nor UO_200 (O_200,N_14057,N_14519);
or UO_201 (O_201,N_13476,N_12251);
nor UO_202 (O_202,N_12525,N_13871);
or UO_203 (O_203,N_14075,N_13629);
nor UO_204 (O_204,N_14684,N_12738);
or UO_205 (O_205,N_14856,N_13804);
or UO_206 (O_206,N_13156,N_13941);
nand UO_207 (O_207,N_13439,N_12340);
or UO_208 (O_208,N_12017,N_13684);
nand UO_209 (O_209,N_13421,N_13712);
nand UO_210 (O_210,N_12420,N_14298);
or UO_211 (O_211,N_14080,N_12267);
or UO_212 (O_212,N_12367,N_14772);
or UO_213 (O_213,N_14565,N_14178);
and UO_214 (O_214,N_13098,N_12147);
nor UO_215 (O_215,N_13861,N_13649);
nor UO_216 (O_216,N_12296,N_12499);
and UO_217 (O_217,N_14875,N_12963);
nand UO_218 (O_218,N_13814,N_13064);
nor UO_219 (O_219,N_12220,N_12711);
xor UO_220 (O_220,N_14316,N_12927);
and UO_221 (O_221,N_12899,N_12191);
or UO_222 (O_222,N_13289,N_13514);
or UO_223 (O_223,N_14675,N_14866);
and UO_224 (O_224,N_12733,N_14568);
nand UO_225 (O_225,N_12744,N_12016);
nand UO_226 (O_226,N_13172,N_14046);
nand UO_227 (O_227,N_12066,N_14629);
and UO_228 (O_228,N_14190,N_13101);
nor UO_229 (O_229,N_14084,N_14751);
or UO_230 (O_230,N_14149,N_14307);
or UO_231 (O_231,N_13415,N_12821);
nand UO_232 (O_232,N_14229,N_13963);
xor UO_233 (O_233,N_13109,N_13664);
or UO_234 (O_234,N_13736,N_13524);
or UO_235 (O_235,N_14973,N_12873);
nor UO_236 (O_236,N_13624,N_12184);
or UO_237 (O_237,N_12699,N_13647);
and UO_238 (O_238,N_14377,N_14992);
and UO_239 (O_239,N_14203,N_13923);
nand UO_240 (O_240,N_14707,N_12553);
nand UO_241 (O_241,N_13140,N_13660);
or UO_242 (O_242,N_13445,N_14537);
nand UO_243 (O_243,N_14501,N_12672);
nand UO_244 (O_244,N_12096,N_12258);
or UO_245 (O_245,N_12784,N_13787);
nor UO_246 (O_246,N_12682,N_12059);
and UO_247 (O_247,N_12960,N_12723);
nor UO_248 (O_248,N_14472,N_12235);
and UO_249 (O_249,N_12464,N_13755);
or UO_250 (O_250,N_13936,N_13724);
nor UO_251 (O_251,N_13121,N_14961);
nor UO_252 (O_252,N_14070,N_14999);
or UO_253 (O_253,N_12607,N_13580);
nor UO_254 (O_254,N_12721,N_12012);
and UO_255 (O_255,N_14513,N_14151);
nor UO_256 (O_256,N_14131,N_12433);
nor UO_257 (O_257,N_13867,N_13959);
nand UO_258 (O_258,N_12749,N_13832);
and UO_259 (O_259,N_14179,N_14156);
or UO_260 (O_260,N_14169,N_13841);
nand UO_261 (O_261,N_13520,N_13933);
nand UO_262 (O_262,N_13127,N_13033);
or UO_263 (O_263,N_14704,N_14320);
or UO_264 (O_264,N_14475,N_13889);
nand UO_265 (O_265,N_12021,N_12459);
nand UO_266 (O_266,N_12117,N_14087);
or UO_267 (O_267,N_12526,N_12039);
nand UO_268 (O_268,N_12048,N_12593);
or UO_269 (O_269,N_14088,N_13147);
nor UO_270 (O_270,N_13799,N_14717);
or UO_271 (O_271,N_14085,N_14380);
nor UO_272 (O_272,N_13390,N_14990);
nand UO_273 (O_273,N_14867,N_13134);
and UO_274 (O_274,N_12125,N_14495);
or UO_275 (O_275,N_14293,N_13899);
nand UO_276 (O_276,N_12734,N_14663);
nor UO_277 (O_277,N_13263,N_13528);
xor UO_278 (O_278,N_13730,N_12883);
or UO_279 (O_279,N_13648,N_13912);
and UO_280 (O_280,N_12269,N_12335);
nor UO_281 (O_281,N_14998,N_12246);
and UO_282 (O_282,N_13209,N_14887);
nor UO_283 (O_283,N_13793,N_14269);
nor UO_284 (O_284,N_13768,N_12042);
and UO_285 (O_285,N_14189,N_12385);
nand UO_286 (O_286,N_13926,N_13538);
nand UO_287 (O_287,N_12388,N_13068);
nor UO_288 (O_288,N_12994,N_13596);
and UO_289 (O_289,N_14754,N_12516);
nor UO_290 (O_290,N_14646,N_13085);
nand UO_291 (O_291,N_12700,N_12218);
and UO_292 (O_292,N_13983,N_12217);
and UO_293 (O_293,N_13023,N_12461);
nand UO_294 (O_294,N_12094,N_14652);
or UO_295 (O_295,N_12693,N_12285);
or UO_296 (O_296,N_12886,N_13837);
nand UO_297 (O_297,N_14095,N_12236);
nor UO_298 (O_298,N_12718,N_14464);
or UO_299 (O_299,N_14427,N_14615);
nand UO_300 (O_300,N_14789,N_12101);
and UO_301 (O_301,N_12077,N_12386);
and UO_302 (O_302,N_14705,N_13757);
nand UO_303 (O_303,N_13419,N_13734);
and UO_304 (O_304,N_12626,N_12968);
nand UO_305 (O_305,N_12004,N_13245);
or UO_306 (O_306,N_13219,N_14636);
nor UO_307 (O_307,N_14608,N_13190);
xor UO_308 (O_308,N_14232,N_13255);
or UO_309 (O_309,N_14135,N_13984);
nor UO_310 (O_310,N_14383,N_14275);
nor UO_311 (O_311,N_12768,N_14854);
nand UO_312 (O_312,N_12376,N_12554);
nand UO_313 (O_313,N_13495,N_14000);
nand UO_314 (O_314,N_12610,N_13689);
nand UO_315 (O_315,N_12108,N_13847);
nor UO_316 (O_316,N_14597,N_14035);
nand UO_317 (O_317,N_14651,N_12344);
nor UO_318 (O_318,N_12331,N_14877);
nand UO_319 (O_319,N_13735,N_12792);
or UO_320 (O_320,N_12957,N_14516);
and UO_321 (O_321,N_12891,N_13878);
nand UO_322 (O_322,N_13508,N_14506);
and UO_323 (O_323,N_14708,N_12977);
and UO_324 (O_324,N_12011,N_14076);
or UO_325 (O_325,N_12698,N_13872);
nor UO_326 (O_326,N_12872,N_12666);
or UO_327 (O_327,N_12692,N_12602);
nor UO_328 (O_328,N_13704,N_13987);
nand UO_329 (O_329,N_13236,N_13835);
and UO_330 (O_330,N_13020,N_14682);
and UO_331 (O_331,N_13845,N_14816);
or UO_332 (O_332,N_14575,N_12057);
or UO_333 (O_333,N_13136,N_13001);
nand UO_334 (O_334,N_13946,N_13242);
nand UO_335 (O_335,N_12882,N_13551);
or UO_336 (O_336,N_12190,N_14243);
nor UO_337 (O_337,N_13469,N_13081);
or UO_338 (O_338,N_12884,N_13040);
nor UO_339 (O_339,N_12831,N_13893);
nor UO_340 (O_340,N_12545,N_13201);
and UO_341 (O_341,N_12260,N_14019);
nor UO_342 (O_342,N_13985,N_13094);
or UO_343 (O_343,N_14445,N_14342);
nand UO_344 (O_344,N_14148,N_12570);
nand UO_345 (O_345,N_14385,N_14549);
and UO_346 (O_346,N_13191,N_13438);
nor UO_347 (O_347,N_12501,N_13529);
nor UO_348 (O_348,N_12364,N_13585);
and UO_349 (O_349,N_14101,N_13314);
and UO_350 (O_350,N_14326,N_14227);
and UO_351 (O_351,N_13996,N_14677);
and UO_352 (O_352,N_14376,N_13678);
and UO_353 (O_353,N_14023,N_12134);
or UO_354 (O_354,N_12481,N_13862);
and UO_355 (O_355,N_12384,N_12178);
nand UO_356 (O_356,N_13759,N_13838);
and UO_357 (O_357,N_12193,N_14638);
or UO_358 (O_358,N_12870,N_14467);
nand UO_359 (O_359,N_14312,N_12546);
nor UO_360 (O_360,N_12457,N_13534);
nor UO_361 (O_361,N_13332,N_12361);
xor UO_362 (O_362,N_13151,N_13815);
nand UO_363 (O_363,N_14648,N_13129);
or UO_364 (O_364,N_13516,N_12573);
or UO_365 (O_365,N_14324,N_12860);
nand UO_366 (O_366,N_14769,N_13706);
nor UO_367 (O_367,N_13739,N_12755);
nand UO_368 (O_368,N_13213,N_14669);
nand UO_369 (O_369,N_12876,N_12253);
nor UO_370 (O_370,N_14104,N_13843);
nand UO_371 (O_371,N_12483,N_14560);
nor UO_372 (O_372,N_14471,N_13840);
or UO_373 (O_373,N_13000,N_14212);
or UO_374 (O_374,N_14617,N_13353);
and UO_375 (O_375,N_13327,N_12469);
nand UO_376 (O_376,N_14985,N_13908);
nor UO_377 (O_377,N_14231,N_13371);
nor UO_378 (O_378,N_12833,N_13919);
nand UO_379 (O_379,N_14081,N_12984);
or UO_380 (O_380,N_14254,N_14957);
nand UO_381 (O_381,N_13611,N_13142);
nor UO_382 (O_382,N_13819,N_13965);
and UO_383 (O_383,N_14871,N_13325);
and UO_384 (O_384,N_13047,N_14067);
or UO_385 (O_385,N_12352,N_12530);
nand UO_386 (O_386,N_12974,N_12049);
or UO_387 (O_387,N_12151,N_14373);
and UO_388 (O_388,N_12585,N_12365);
or UO_389 (O_389,N_12013,N_14805);
or UO_390 (O_390,N_14843,N_13096);
nor UO_391 (O_391,N_13133,N_12348);
nand UO_392 (O_392,N_12023,N_12864);
or UO_393 (O_393,N_14820,N_13009);
or UO_394 (O_394,N_14077,N_13932);
nand UO_395 (O_395,N_12653,N_12781);
nor UO_396 (O_396,N_13685,N_13135);
nor UO_397 (O_397,N_12002,N_13794);
or UO_398 (O_398,N_14800,N_14655);
and UO_399 (O_399,N_12560,N_14409);
or UO_400 (O_400,N_13066,N_12986);
nand UO_401 (O_401,N_13232,N_12688);
and UO_402 (O_402,N_14770,N_14032);
or UO_403 (O_403,N_14919,N_13481);
nor UO_404 (O_404,N_14909,N_13018);
and UO_405 (O_405,N_13954,N_12814);
nand UO_406 (O_406,N_14042,N_12695);
nand UO_407 (O_407,N_13829,N_14804);
nor UO_408 (O_408,N_12237,N_13393);
and UO_409 (O_409,N_12127,N_12858);
nand UO_410 (O_410,N_14142,N_14073);
and UO_411 (O_411,N_13890,N_14021);
nor UO_412 (O_412,N_14234,N_12455);
or UO_413 (O_413,N_12912,N_13429);
nor UO_414 (O_414,N_13957,N_13077);
or UO_415 (O_415,N_14415,N_14079);
and UO_416 (O_416,N_13271,N_12153);
or UO_417 (O_417,N_14771,N_13642);
or UO_418 (O_418,N_12985,N_13603);
and UO_419 (O_419,N_12563,N_14176);
and UO_420 (O_420,N_14273,N_14791);
nand UO_421 (O_421,N_13661,N_12719);
or UO_422 (O_422,N_12533,N_14204);
nor UO_423 (O_423,N_12319,N_12550);
nand UO_424 (O_424,N_12965,N_12060);
and UO_425 (O_425,N_13716,N_14451);
or UO_426 (O_426,N_12850,N_12907);
or UO_427 (O_427,N_12322,N_12701);
nand UO_428 (O_428,N_14323,N_13012);
or UO_429 (O_429,N_12419,N_13349);
nand UO_430 (O_430,N_13673,N_14177);
nand UO_431 (O_431,N_14551,N_13281);
nand UO_432 (O_432,N_14743,N_14881);
nand UO_433 (O_433,N_12432,N_13279);
nand UO_434 (O_434,N_14818,N_13221);
and UO_435 (O_435,N_12382,N_14941);
nand UO_436 (O_436,N_12707,N_13489);
nand UO_437 (O_437,N_14005,N_13261);
nand UO_438 (O_438,N_12223,N_12853);
nor UO_439 (O_439,N_13719,N_14355);
or UO_440 (O_440,N_12660,N_13947);
nand UO_441 (O_441,N_14366,N_13784);
nor UO_442 (O_442,N_12294,N_14857);
nand UO_443 (O_443,N_14040,N_13776);
nand UO_444 (O_444,N_12787,N_14476);
and UO_445 (O_445,N_14022,N_12287);
nand UO_446 (O_446,N_13709,N_13749);
nand UO_447 (O_447,N_13466,N_13462);
and UO_448 (O_448,N_14145,N_13075);
nand UO_449 (O_449,N_14846,N_13834);
xor UO_450 (O_450,N_14773,N_14140);
nand UO_451 (O_451,N_13334,N_12917);
nor UO_452 (O_452,N_13612,N_13937);
nor UO_453 (O_453,N_14795,N_14158);
nand UO_454 (O_454,N_13072,N_13764);
nand UO_455 (O_455,N_12152,N_12289);
and UO_456 (O_456,N_13161,N_14053);
xor UO_457 (O_457,N_13416,N_12136);
nor UO_458 (O_458,N_14173,N_14327);
and UO_459 (O_459,N_13891,N_12621);
or UO_460 (O_460,N_13500,N_14465);
nor UO_461 (O_461,N_12471,N_12678);
nand UO_462 (O_462,N_12896,N_12239);
and UO_463 (O_463,N_13657,N_14971);
or UO_464 (O_464,N_14074,N_14485);
nor UO_465 (O_465,N_14061,N_14386);
nor UO_466 (O_466,N_12041,N_12798);
or UO_467 (O_467,N_14037,N_14191);
nand UO_468 (O_468,N_14888,N_12473);
or UO_469 (O_469,N_12282,N_12399);
nand UO_470 (O_470,N_13491,N_12548);
nand UO_471 (O_471,N_14062,N_14645);
and UO_472 (O_472,N_14164,N_13267);
nor UO_473 (O_473,N_12262,N_14268);
nor UO_474 (O_474,N_14259,N_13582);
nand UO_475 (O_475,N_13818,N_13887);
nand UO_476 (O_476,N_12871,N_13039);
and UO_477 (O_477,N_14460,N_13515);
or UO_478 (O_478,N_13381,N_13727);
xnor UO_479 (O_479,N_13144,N_12009);
or UO_480 (O_480,N_13208,N_12636);
nand UO_481 (O_481,N_12754,N_14146);
nand UO_482 (O_482,N_14865,N_14421);
nor UO_483 (O_483,N_13278,N_13010);
or UO_484 (O_484,N_12334,N_14838);
xor UO_485 (O_485,N_12456,N_12709);
or UO_486 (O_486,N_12036,N_13167);
nand UO_487 (O_487,N_12706,N_14253);
and UO_488 (O_488,N_12845,N_13882);
nor UO_489 (O_489,N_12072,N_12264);
nor UO_490 (O_490,N_12497,N_14785);
and UO_491 (O_491,N_13548,N_13374);
or UO_492 (O_492,N_13915,N_13934);
or UO_493 (O_493,N_12283,N_13539);
or UO_494 (O_494,N_14256,N_12332);
nand UO_495 (O_495,N_13956,N_14777);
nand UO_496 (O_496,N_14947,N_12741);
and UO_497 (O_497,N_13535,N_12198);
nand UO_498 (O_498,N_13587,N_14803);
nand UO_499 (O_499,N_12203,N_14858);
and UO_500 (O_500,N_14727,N_12291);
or UO_501 (O_501,N_12392,N_14403);
nand UO_502 (O_502,N_12940,N_13468);
nand UO_503 (O_503,N_12442,N_13309);
and UO_504 (O_504,N_12508,N_13061);
and UO_505 (O_505,N_13668,N_12085);
nor UO_506 (O_506,N_14952,N_14869);
nand UO_507 (O_507,N_14914,N_12679);
and UO_508 (O_508,N_12362,N_12310);
nor UO_509 (O_509,N_13226,N_14956);
nand UO_510 (O_510,N_14267,N_12449);
and UO_511 (O_511,N_13751,N_12210);
nor UO_512 (O_512,N_14016,N_12839);
and UO_513 (O_513,N_13518,N_13397);
nor UO_514 (O_514,N_13527,N_14311);
and UO_515 (O_515,N_13104,N_13153);
or UO_516 (O_516,N_14400,N_13783);
nand UO_517 (O_517,N_13123,N_12520);
xor UO_518 (O_518,N_13598,N_12342);
xnor UO_519 (O_519,N_13433,N_12980);
nand UO_520 (O_520,N_12030,N_14862);
or UO_521 (O_521,N_12186,N_13067);
or UO_522 (O_522,N_12969,N_14930);
or UO_523 (O_523,N_14538,N_13441);
nand UO_524 (O_524,N_13270,N_14199);
nor UO_525 (O_525,N_12122,N_13569);
nor UO_526 (O_526,N_12911,N_13961);
or UO_527 (O_527,N_13615,N_13152);
nor UO_528 (O_528,N_13558,N_14063);
or UO_529 (O_529,N_14860,N_14759);
nor UO_530 (O_530,N_13589,N_12846);
nor UO_531 (O_531,N_13171,N_14300);
nand UO_532 (O_532,N_13224,N_14296);
or UO_533 (O_533,N_14371,N_13235);
nor UO_534 (O_534,N_14429,N_12547);
and UO_535 (O_535,N_12836,N_14616);
nor UO_536 (O_536,N_14978,N_14052);
nand UO_537 (O_537,N_14123,N_12460);
and UO_538 (O_538,N_12668,N_14049);
nor UO_539 (O_539,N_12110,N_14043);
nand UO_540 (O_540,N_13467,N_13945);
and UO_541 (O_541,N_12292,N_13640);
or UO_542 (O_542,N_12000,N_12215);
or UO_543 (O_543,N_12349,N_14792);
nand UO_544 (O_544,N_14509,N_13102);
and UO_545 (O_545,N_13053,N_12339);
nand UO_546 (O_546,N_13063,N_13272);
or UO_547 (O_547,N_13691,N_13105);
and UO_548 (O_548,N_12064,N_13694);
and UO_549 (O_549,N_12179,N_12555);
or UO_550 (O_550,N_12715,N_13431);
or UO_551 (O_551,N_13525,N_12783);
nor UO_552 (O_552,N_13400,N_14603);
and UO_553 (O_553,N_12931,N_12949);
and UO_554 (O_554,N_14121,N_13916);
and UO_555 (O_555,N_14633,N_14662);
nand UO_556 (O_556,N_14407,N_12123);
xnor UO_557 (O_557,N_12033,N_13169);
nor UO_558 (O_558,N_13857,N_14484);
or UO_559 (O_559,N_13099,N_14263);
or UO_560 (O_560,N_12144,N_13731);
nand UO_561 (O_561,N_12437,N_13252);
nor UO_562 (O_562,N_14186,N_14090);
or UO_563 (O_563,N_13382,N_14014);
xor UO_564 (O_564,N_13669,N_14432);
nand UO_565 (O_565,N_12569,N_13995);
and UO_566 (O_566,N_12412,N_14510);
or UO_567 (O_567,N_14557,N_12835);
nor UO_568 (O_568,N_14222,N_12737);
and UO_569 (O_569,N_12987,N_14059);
and UO_570 (O_570,N_12252,N_13076);
or UO_571 (O_571,N_14447,N_14200);
nand UO_572 (O_572,N_14097,N_12745);
nor UO_573 (O_573,N_14533,N_12972);
and UO_574 (O_574,N_13581,N_13070);
and UO_575 (O_575,N_14632,N_13974);
xnor UO_576 (O_576,N_14781,N_14277);
nand UO_577 (O_577,N_12333,N_14001);
or UO_578 (O_578,N_14518,N_12275);
and UO_579 (O_579,N_12478,N_14969);
nor UO_580 (O_580,N_12233,N_14855);
nand UO_581 (O_581,N_14913,N_13497);
nor UO_582 (O_582,N_14983,N_14889);
or UO_583 (O_583,N_14822,N_12371);
nor UO_584 (O_584,N_12454,N_12740);
nand UO_585 (O_585,N_12541,N_12630);
nand UO_586 (O_586,N_13482,N_13227);
nand UO_587 (O_587,N_14262,N_13865);
nand UO_588 (O_588,N_12417,N_12486);
and UO_589 (O_589,N_14927,N_13772);
or UO_590 (O_590,N_13338,N_14228);
nand UO_591 (O_591,N_13412,N_12489);
nor UO_592 (O_592,N_12578,N_13836);
and UO_593 (O_593,N_14321,N_14261);
nor UO_594 (O_594,N_12574,N_12659);
and UO_595 (O_595,N_12726,N_12080);
nor UO_596 (O_596,N_14797,N_13322);
nand UO_597 (O_597,N_14038,N_14765);
nor UO_598 (O_598,N_13301,N_13998);
nand UO_599 (O_599,N_13549,N_13780);
nor UO_600 (O_600,N_13705,N_12114);
and UO_601 (O_601,N_14096,N_13202);
xnor UO_602 (O_602,N_13718,N_12724);
nand UO_603 (O_603,N_13982,N_14500);
or UO_604 (O_604,N_14539,N_14942);
nor UO_605 (O_605,N_12586,N_12407);
nand UO_606 (O_606,N_13786,N_14488);
nand UO_607 (O_607,N_12893,N_12185);
nor UO_608 (O_608,N_14459,N_14344);
xor UO_609 (O_609,N_14489,N_14801);
nand UO_610 (O_610,N_13028,N_12770);
and UO_611 (O_611,N_12490,N_14900);
nor UO_612 (O_612,N_12148,N_12312);
nand UO_613 (O_613,N_14276,N_13976);
nor UO_614 (O_614,N_12579,N_13437);
or UO_615 (O_615,N_12971,N_12910);
nand UO_616 (O_616,N_12805,N_14830);
or UO_617 (O_617,N_13257,N_13566);
and UO_618 (O_618,N_14681,N_13417);
or UO_619 (O_619,N_12423,N_12729);
nand UO_620 (O_620,N_12843,N_14911);
nand UO_621 (O_621,N_12201,N_12528);
and UO_622 (O_622,N_13239,N_12622);
and UO_623 (O_623,N_13312,N_12712);
nor UO_624 (O_624,N_13432,N_14335);
or UO_625 (O_625,N_12180,N_13656);
nor UO_626 (O_626,N_12758,N_14006);
or UO_627 (O_627,N_14147,N_14017);
or UO_628 (O_628,N_14008,N_12811);
nand UO_629 (O_629,N_14255,N_13032);
or UO_630 (O_630,N_14712,N_14762);
nor UO_631 (O_631,N_12956,N_14977);
nand UO_632 (O_632,N_12652,N_12261);
or UO_633 (O_633,N_14398,N_13036);
and UO_634 (O_634,N_13449,N_12714);
nand UO_635 (O_635,N_14350,N_14569);
nand UO_636 (O_636,N_13343,N_13858);
and UO_637 (O_637,N_14523,N_14689);
and UO_638 (O_638,N_13435,N_14667);
or UO_639 (O_639,N_12325,N_13082);
and UO_640 (O_640,N_14987,N_13750);
nand UO_641 (O_641,N_13436,N_14692);
nand UO_642 (O_642,N_13290,N_12825);
nor UO_643 (O_643,N_12435,N_13315);
or UO_644 (O_644,N_13424,N_12696);
and UO_645 (O_645,N_14213,N_13407);
or UO_646 (O_646,N_14031,N_12259);
xnor UO_647 (O_647,N_14011,N_13714);
xnor UO_648 (O_648,N_13175,N_13403);
and UO_649 (O_649,N_13771,N_14339);
and UO_650 (O_650,N_13319,N_12557);
nand UO_651 (O_651,N_14827,N_13282);
and UO_652 (O_652,N_14905,N_12549);
and UO_653 (O_653,N_12092,N_14641);
and UO_654 (O_654,N_12034,N_13472);
nor UO_655 (O_655,N_13233,N_14233);
nand UO_656 (O_656,N_13442,N_14572);
nand UO_657 (O_657,N_13035,N_13748);
nor UO_658 (O_658,N_14526,N_13973);
nor UO_659 (O_659,N_12808,N_14410);
nand UO_660 (O_660,N_12081,N_13797);
and UO_661 (O_661,N_12898,N_12771);
or UO_662 (O_662,N_13396,N_12323);
and UO_663 (O_663,N_13821,N_14329);
and UO_664 (O_664,N_12138,N_13002);
and UO_665 (O_665,N_14482,N_13556);
or UO_666 (O_666,N_12063,N_13173);
nand UO_667 (O_667,N_13687,N_13881);
and UO_668 (O_668,N_12667,N_13864);
nor UO_669 (O_669,N_13543,N_13179);
or UO_670 (O_670,N_12192,N_12676);
and UO_671 (O_671,N_14556,N_13675);
nor UO_672 (O_672,N_12538,N_12255);
nand UO_673 (O_673,N_14003,N_14133);
or UO_674 (O_674,N_12324,N_12441);
xnor UO_675 (O_675,N_12575,N_14314);
nor UO_676 (O_676,N_14582,N_14143);
or UO_677 (O_677,N_13352,N_14988);
or UO_678 (O_678,N_14020,N_13848);
and UO_679 (O_679,N_13285,N_14806);
xor UO_680 (O_680,N_14581,N_13262);
and UO_681 (O_681,N_13302,N_13326);
and UO_682 (O_682,N_13798,N_13817);
or UO_683 (O_683,N_12299,N_13316);
nand UO_684 (O_684,N_13710,N_12165);
nor UO_685 (O_685,N_14955,N_14137);
nand UO_686 (O_686,N_13086,N_14922);
and UO_687 (O_687,N_14435,N_14605);
nor UO_688 (O_688,N_14221,N_13765);
nand UO_689 (O_689,N_14374,N_12027);
and UO_690 (O_690,N_14353,N_14908);
or UO_691 (O_691,N_13266,N_13790);
nor UO_692 (O_692,N_14920,N_13484);
xor UO_693 (O_693,N_13610,N_13570);
nor UO_694 (O_694,N_14473,N_12452);
and UO_695 (O_695,N_14265,N_13414);
and UO_696 (O_696,N_13042,N_12440);
or UO_697 (O_697,N_12273,N_14150);
xnor UO_698 (O_698,N_13625,N_14744);
and UO_699 (O_699,N_14578,N_12326);
and UO_700 (O_700,N_12309,N_13788);
nor UO_701 (O_701,N_14452,N_14995);
and UO_702 (O_702,N_14390,N_12119);
nand UO_703 (O_703,N_12303,N_13505);
nand UO_704 (O_704,N_14160,N_12357);
or UO_705 (O_705,N_12539,N_13243);
and UO_706 (O_706,N_13621,N_13641);
nor UO_707 (O_707,N_13050,N_12581);
xnor UO_708 (O_708,N_13994,N_14136);
nor UO_709 (O_709,N_13447,N_12644);
and UO_710 (O_710,N_13677,N_12677);
nor UO_711 (O_711,N_12014,N_14209);
nand UO_712 (O_712,N_14416,N_12941);
and UO_713 (O_713,N_14725,N_14964);
or UO_714 (O_714,N_14752,N_12820);
nand UO_715 (O_715,N_12051,N_14571);
or UO_716 (O_716,N_14266,N_12359);
and UO_717 (O_717,N_13897,N_14102);
nor UO_718 (O_718,N_14543,N_14917);
and UO_719 (O_719,N_14614,N_14315);
nand UO_720 (O_720,N_12923,N_14089);
or UO_721 (O_721,N_13605,N_13522);
nor UO_722 (O_722,N_12954,N_14530);
nand UO_723 (O_723,N_14250,N_12822);
nor UO_724 (O_724,N_14361,N_13177);
and UO_725 (O_725,N_14716,N_13952);
nor UO_726 (O_726,N_13894,N_13540);
and UO_727 (O_727,N_14453,N_14368);
nor UO_728 (O_728,N_13130,N_12556);
or UO_729 (O_729,N_12043,N_14980);
xor UO_730 (O_730,N_14736,N_13205);
and UO_731 (O_731,N_13576,N_14718);
or UO_732 (O_732,N_13997,N_13275);
nor UO_733 (O_733,N_14661,N_14047);
or UO_734 (O_734,N_12671,N_14719);
nor UO_735 (O_735,N_12849,N_13746);
and UO_736 (O_736,N_13311,N_13651);
nor UO_737 (O_737,N_12790,N_14466);
or UO_738 (O_738,N_12919,N_14498);
nor UO_739 (O_739,N_14165,N_13546);
and UO_740 (O_740,N_14696,N_13383);
or UO_741 (O_741,N_14331,N_12115);
nor UO_742 (O_742,N_12518,N_12887);
nand UO_743 (O_743,N_14444,N_14656);
and UO_744 (O_744,N_13440,N_13163);
nor UO_745 (O_745,N_14162,N_12316);
or UO_746 (O_746,N_12288,N_12824);
or UO_747 (O_747,N_12226,N_12750);
nand UO_748 (O_748,N_14673,N_12409);
or UO_749 (O_749,N_13037,N_13452);
nor UO_750 (O_750,N_14287,N_14493);
or UO_751 (O_751,N_13183,N_12172);
or UO_752 (O_752,N_13410,N_13591);
nand UO_753 (O_753,N_12727,N_12513);
or UO_754 (O_754,N_13386,N_12221);
nand UO_755 (O_755,N_14668,N_12052);
nand UO_756 (O_756,N_13145,N_14492);
and UO_757 (O_757,N_13839,N_14885);
xor UO_758 (O_758,N_14732,N_13006);
nand UO_759 (O_759,N_14644,N_13291);
or UO_760 (O_760,N_12534,N_14428);
nor UO_761 (O_761,N_12479,N_13526);
and UO_762 (O_762,N_12589,N_12542);
or UO_763 (O_763,N_12088,N_12658);
nor UO_764 (O_764,N_13454,N_12690);
nand UO_765 (O_765,N_13486,N_14666);
and UO_766 (O_766,N_12229,N_13256);
nor UO_767 (O_767,N_12320,N_14068);
nand UO_768 (O_768,N_12327,N_14525);
nand UO_769 (O_769,N_14654,N_12990);
or UO_770 (O_770,N_13446,N_12797);
nand UO_771 (O_771,N_13846,N_14033);
nand UO_772 (O_772,N_12674,N_13483);
nand UO_773 (O_773,N_13357,N_14729);
or UO_774 (O_774,N_13477,N_13851);
nor UO_775 (O_775,N_14375,N_13512);
nand UO_776 (O_776,N_12788,N_14607);
nor UO_777 (O_777,N_14188,N_13722);
and UO_778 (O_778,N_13276,N_14831);
or UO_779 (O_779,N_14505,N_13143);
and UO_780 (O_780,N_12983,N_12408);
nor UO_781 (O_781,N_12861,N_13220);
nor UO_782 (O_782,N_13509,N_12673);
and UO_783 (O_783,N_14982,N_13654);
and UO_784 (O_784,N_14665,N_12139);
nand UO_785 (O_785,N_14066,N_13810);
nand UO_786 (O_786,N_12003,N_14901);
nand UO_787 (O_787,N_14589,N_12828);
nor UO_788 (O_788,N_14397,N_13579);
or UO_789 (O_789,N_13003,N_12769);
nand UO_790 (O_790,N_14071,N_12565);
nor UO_791 (O_791,N_12493,N_13927);
nand UO_792 (O_792,N_12996,N_12966);
or UO_793 (O_793,N_14713,N_14009);
and UO_794 (O_794,N_14778,N_14094);
or UO_795 (O_795,N_14864,N_14278);
nor UO_796 (O_796,N_12112,N_13139);
nor UO_797 (O_797,N_14029,N_14967);
nor UO_798 (O_798,N_14761,N_12529);
and UO_799 (O_799,N_12681,N_14933);
or UO_800 (O_800,N_13935,N_14225);
and UO_801 (O_801,N_12571,N_12402);
and UO_802 (O_802,N_12040,N_14328);
and UO_803 (O_803,N_14715,N_13078);
nand UO_804 (O_804,N_14970,N_13490);
or UO_805 (O_805,N_13630,N_12596);
and UO_806 (O_806,N_12321,N_13643);
nand UO_807 (O_807,N_13286,N_13212);
or UO_808 (O_808,N_13723,N_13399);
or UO_809 (O_809,N_13016,N_14332);
nand UO_810 (O_810,N_14286,N_13575);
xnor UO_811 (O_811,N_14241,N_14248);
nor UO_812 (O_812,N_12204,N_12862);
nor UO_813 (O_813,N_12623,N_14013);
and UO_814 (O_814,N_12559,N_14798);
nand UO_815 (O_815,N_14739,N_12881);
nand UO_816 (O_816,N_12844,N_13802);
nor UO_817 (O_817,N_14903,N_12290);
or UO_818 (O_818,N_12720,N_12535);
or UO_819 (O_819,N_12584,N_13350);
and UO_820 (O_820,N_13715,N_12866);
nor UO_821 (O_821,N_12369,N_12503);
nand UO_822 (O_822,N_13141,N_14161);
and UO_823 (O_823,N_13679,N_13972);
nand UO_824 (O_824,N_14490,N_13398);
nor UO_825 (O_825,N_13713,N_12592);
and UO_826 (O_826,N_14695,N_12970);
nand UO_827 (O_827,N_14604,N_12804);
or UO_828 (O_828,N_12609,N_12874);
nor UO_829 (O_829,N_14167,N_13960);
and UO_830 (O_830,N_12196,N_14620);
and UO_831 (O_831,N_12047,N_14208);
xor UO_832 (O_832,N_13451,N_13886);
and UO_833 (O_833,N_12580,N_12208);
or UO_834 (O_834,N_14317,N_13007);
or UO_835 (O_835,N_13363,N_14215);
nand UO_836 (O_836,N_13434,N_12958);
nand UO_837 (O_837,N_14334,N_13328);
or UO_838 (O_838,N_14902,N_14214);
nor UO_839 (O_839,N_14780,N_14679);
and UO_840 (O_840,N_13967,N_14086);
and UO_841 (O_841,N_13110,N_12336);
nor UO_842 (O_842,N_12395,N_14779);
or UO_843 (O_843,N_12597,N_12345);
nor UO_844 (O_844,N_12146,N_14155);
nand UO_845 (O_845,N_12202,N_13938);
nand UO_846 (O_846,N_12078,N_14405);
or UO_847 (O_847,N_13672,N_12351);
and UO_848 (O_848,N_13283,N_14157);
and UO_849 (O_849,N_14621,N_13692);
or UO_850 (O_850,N_13807,N_12976);
nor UO_851 (O_851,N_12517,N_13251);
nor UO_852 (O_852,N_12300,N_14760);
nand UO_853 (O_853,N_13203,N_13898);
nand UO_854 (O_854,N_14776,N_13210);
nor UO_855 (O_855,N_14098,N_13126);
or UO_856 (O_856,N_14392,N_12120);
nor UO_857 (O_857,N_12168,N_13292);
or UO_858 (O_858,N_13480,N_13015);
or UO_859 (O_859,N_12271,N_12591);
or UO_860 (O_860,N_12308,N_12240);
and UO_861 (O_861,N_14691,N_12015);
nor UO_862 (O_862,N_13425,N_14512);
nor UO_863 (O_863,N_13646,N_13308);
and UO_864 (O_864,N_14547,N_12007);
or UO_865 (O_865,N_14294,N_14842);
and UO_866 (O_866,N_14433,N_12162);
nor UO_867 (O_867,N_12444,N_13095);
and UO_868 (O_868,N_13760,N_12074);
or UO_869 (O_869,N_14570,N_14783);
nor UO_870 (O_870,N_14742,N_14630);
and UO_871 (O_871,N_12651,N_14319);
and UO_872 (O_872,N_14637,N_12665);
or UO_873 (O_873,N_13717,N_14627);
and UO_874 (O_874,N_12145,N_14139);
or UO_875 (O_875,N_12400,N_12430);
or UO_876 (O_876,N_12981,N_12854);
nand UO_877 (O_877,N_12967,N_12664);
and UO_878 (O_878,N_13376,N_13026);
nand UO_879 (O_879,N_12857,N_14876);
nor UO_880 (O_880,N_14918,N_14698);
or UO_881 (O_881,N_12026,N_14336);
nor UO_882 (O_882,N_12646,N_12082);
nand UO_883 (O_883,N_12801,N_12973);
nor UO_884 (O_884,N_14193,N_12612);
and UO_885 (O_885,N_13079,N_14833);
or UO_886 (O_886,N_12759,N_13620);
nor UO_887 (O_887,N_12263,N_12355);
nor UO_888 (O_888,N_13046,N_13310);
or UO_889 (O_889,N_14891,N_14217);
or UO_890 (O_890,N_12129,N_14893);
nor UO_891 (O_891,N_12154,N_14936);
nand UO_892 (O_892,N_12779,N_14520);
or UO_893 (O_893,N_13029,N_12902);
nand UO_894 (O_894,N_13264,N_14341);
nand UO_895 (O_895,N_13752,N_13860);
and UO_896 (O_896,N_12952,N_12631);
xor UO_897 (O_897,N_13159,N_13639);
or UO_898 (O_898,N_14924,N_12279);
nor UO_899 (O_899,N_14309,N_12453);
nor UO_900 (O_900,N_12913,N_12167);
or UO_901 (O_901,N_13866,N_13394);
and UO_902 (O_902,N_12885,N_14249);
nor UO_903 (O_903,N_12829,N_14879);
and UO_904 (O_904,N_14910,N_12087);
or UO_905 (O_905,N_14448,N_12383);
and UO_906 (O_906,N_12065,N_12418);
nand UO_907 (O_907,N_13330,N_12583);
or UO_908 (O_908,N_14163,N_14274);
nand UO_909 (O_909,N_12742,N_14758);
or UO_910 (O_910,N_12527,N_13388);
or UO_911 (O_911,N_14587,N_14240);
and UO_912 (O_912,N_12375,N_12018);
nand UO_913 (O_913,N_14757,N_14730);
nor UO_914 (O_914,N_14844,N_12716);
nand UO_915 (O_915,N_13459,N_14197);
nor UO_916 (O_916,N_12368,N_13019);
or UO_917 (O_917,N_13813,N_13550);
nand UO_918 (O_918,N_12268,N_13298);
and UO_919 (O_919,N_13681,N_14065);
and UO_920 (O_920,N_14548,N_12878);
nand UO_921 (O_921,N_12374,N_12381);
nor UO_922 (O_922,N_13089,N_14601);
nor UO_923 (O_923,N_12169,N_13782);
and UO_924 (O_924,N_12511,N_13989);
or UO_925 (O_925,N_14154,N_13300);
nand UO_926 (O_926,N_12328,N_14676);
or UO_927 (O_927,N_14579,N_14442);
nand UO_928 (O_928,N_14944,N_14584);
nand UO_929 (O_929,N_13618,N_14649);
or UO_930 (O_930,N_13323,N_14552);
nor UO_931 (O_931,N_13658,N_12598);
nand UO_932 (O_932,N_13176,N_12182);
and UO_933 (O_933,N_14122,N_14438);
or UO_934 (O_934,N_14206,N_14330);
or UO_935 (O_935,N_13593,N_14230);
and UO_936 (O_936,N_13552,N_14236);
xor UO_937 (O_937,N_12448,N_14039);
or UO_938 (O_938,N_13345,N_12436);
nand UO_939 (O_939,N_13418,N_13977);
nor UO_940 (O_940,N_13479,N_13562);
or UO_941 (O_941,N_14166,N_12832);
nor UO_942 (O_942,N_12343,N_14886);
and UO_943 (O_943,N_12416,N_13461);
and UO_944 (O_944,N_12491,N_14083);
nand UO_945 (O_945,N_12988,N_14680);
or UO_946 (O_946,N_13544,N_13389);
and UO_947 (O_947,N_12424,N_13619);
or UO_948 (O_948,N_13254,N_14873);
nand UO_949 (O_949,N_14388,N_13384);
or UO_950 (O_950,N_13638,N_13697);
and UO_951 (O_951,N_12877,N_14693);
nand UO_952 (O_952,N_13331,N_12149);
nand UO_953 (O_953,N_14625,N_14790);
nand UO_954 (O_954,N_13707,N_14446);
or UO_955 (O_955,N_14413,N_12126);
nor UO_956 (O_956,N_13055,N_14768);
or UO_957 (O_957,N_12735,N_13572);
nor UO_958 (O_958,N_13626,N_12561);
and UO_959 (O_959,N_13636,N_14746);
or UO_960 (O_960,N_14404,N_12451);
nor UO_961 (O_961,N_13948,N_13305);
or UO_962 (O_962,N_12616,N_14823);
or UO_963 (O_963,N_13682,N_14224);
xor UO_964 (O_964,N_13460,N_14508);
and UO_965 (O_965,N_12953,N_12044);
nand UO_966 (O_966,N_12618,N_13803);
or UO_967 (O_967,N_12856,N_12054);
nor UO_968 (O_968,N_14347,N_14845);
or UO_969 (O_969,N_14289,N_14109);
and UO_970 (O_970,N_14826,N_13111);
or UO_971 (O_971,N_14456,N_13913);
nor UO_972 (O_972,N_14418,N_14599);
or UO_973 (O_973,N_13907,N_13116);
xnor UO_974 (O_974,N_13831,N_12938);
nor UO_975 (O_975,N_13113,N_13444);
nor UO_976 (O_976,N_14997,N_14767);
nor UO_977 (O_977,N_12684,N_12662);
and UO_978 (O_978,N_14634,N_13038);
nand UO_979 (O_979,N_13487,N_12892);
nand UO_980 (O_980,N_14153,N_14401);
nand UO_981 (O_981,N_14671,N_12964);
and UO_982 (O_982,N_12629,N_12635);
or UO_983 (O_983,N_14026,N_13966);
nand UO_984 (O_984,N_12241,N_12006);
and UO_985 (O_985,N_13344,N_12669);
nand UO_986 (O_986,N_14349,N_12305);
nor UO_987 (O_987,N_13229,N_14441);
nand UO_988 (O_988,N_14594,N_14697);
or UO_989 (O_989,N_13777,N_12084);
and UO_990 (O_990,N_12763,N_14251);
or UO_991 (O_991,N_13080,N_12099);
nor UO_992 (O_992,N_13728,N_14808);
or UO_993 (O_993,N_13914,N_13686);
and UO_994 (O_994,N_14479,N_13738);
nand UO_995 (O_995,N_13733,N_12834);
nand UO_996 (O_996,N_14411,N_13943);
or UO_997 (O_997,N_14018,N_14511);
or UO_998 (O_998,N_14012,N_13609);
and UO_999 (O_999,N_13968,N_12183);
nand UO_1000 (O_1000,N_12143,N_14559);
nor UO_1001 (O_1001,N_14172,N_14481);
and UO_1002 (O_1002,N_12930,N_12512);
and UO_1003 (O_1003,N_12809,N_12642);
and UO_1004 (O_1004,N_14282,N_12680);
and UO_1005 (O_1005,N_13100,N_12020);
nand UO_1006 (O_1006,N_12177,N_12005);
or UO_1007 (O_1007,N_13870,N_13430);
nor UO_1008 (O_1008,N_12090,N_13695);
nand UO_1009 (O_1009,N_12841,N_14297);
nor UO_1010 (O_1010,N_13925,N_12450);
and UO_1011 (O_1011,N_14602,N_14399);
nor UO_1012 (O_1012,N_13910,N_12643);
nand UO_1013 (O_1013,N_13494,N_13763);
xnor UO_1014 (O_1014,N_14678,N_14940);
and UO_1015 (O_1015,N_14406,N_13753);
or UO_1016 (O_1016,N_14882,N_13970);
or UO_1017 (O_1017,N_13547,N_14351);
nor UO_1018 (O_1018,N_12925,N_12079);
nor UO_1019 (O_1019,N_14618,N_14938);
and UO_1020 (O_1020,N_14766,N_13536);
and UO_1021 (O_1021,N_12091,N_13511);
and UO_1022 (O_1022,N_13025,N_13574);
nand UO_1023 (O_1023,N_12507,N_12029);
and UO_1024 (O_1024,N_12076,N_14794);
and UO_1025 (O_1025,N_12106,N_14325);
nand UO_1026 (O_1026,N_14890,N_13674);
and UO_1027 (O_1027,N_12301,N_13406);
nor UO_1028 (O_1028,N_13297,N_14367);
or UO_1029 (O_1029,N_13670,N_14852);
and UO_1030 (O_1030,N_12024,N_14733);
nor UO_1031 (O_1031,N_13065,N_12428);
xnor UO_1032 (O_1032,N_13132,N_13939);
and UO_1033 (O_1033,N_14381,N_12194);
and UO_1034 (O_1034,N_12815,N_12638);
nor UO_1035 (O_1035,N_13317,N_13465);
nor UO_1036 (O_1036,N_12510,N_12318);
nand UO_1037 (O_1037,N_13106,N_14929);
nor UO_1038 (O_1038,N_14626,N_13294);
and UO_1039 (O_1039,N_13362,N_13721);
or UO_1040 (O_1040,N_12908,N_14099);
or UO_1041 (O_1041,N_14963,N_12888);
or UO_1042 (O_1042,N_14141,N_12045);
or UO_1043 (O_1043,N_13346,N_13702);
xnor UO_1044 (O_1044,N_14382,N_13162);
nor UO_1045 (O_1045,N_14198,N_14487);
or UO_1046 (O_1046,N_12337,N_12786);
nor UO_1047 (O_1047,N_12050,N_12751);
and UO_1048 (O_1048,N_13553,N_12494);
nor UO_1049 (O_1049,N_12111,N_12936);
and UO_1050 (O_1050,N_14305,N_12121);
nor UO_1051 (O_1051,N_14932,N_14809);
nor UO_1052 (O_1052,N_12993,N_13530);
and UO_1053 (O_1053,N_13247,N_13249);
nor UO_1054 (O_1054,N_14745,N_14836);
nor UO_1055 (O_1055,N_13217,N_13324);
nor UO_1056 (O_1056,N_12945,N_12722);
nand UO_1057 (O_1057,N_13368,N_12242);
nor UO_1058 (O_1058,N_13228,N_12816);
nand UO_1059 (O_1059,N_13904,N_13354);
and UO_1060 (O_1060,N_13711,N_12415);
nand UO_1061 (O_1061,N_12500,N_13827);
and UO_1062 (O_1062,N_14870,N_13842);
nand UO_1063 (O_1063,N_14606,N_12485);
nand UO_1064 (O_1064,N_14439,N_14402);
and UO_1065 (O_1065,N_13391,N_12868);
nand UO_1066 (O_1066,N_13200,N_12131);
or UO_1067 (O_1067,N_13969,N_14036);
and UO_1068 (O_1068,N_12413,N_13504);
nor UO_1069 (O_1069,N_13348,N_12731);
nor UO_1070 (O_1070,N_14714,N_12488);
nor UO_1071 (O_1071,N_13124,N_14580);
or UO_1072 (O_1072,N_12372,N_13071);
nor UO_1073 (O_1073,N_13268,N_12639);
nand UO_1074 (O_1074,N_13455,N_12214);
nor UO_1075 (O_1075,N_14907,N_12293);
nand UO_1076 (O_1076,N_12905,N_12394);
or UO_1077 (O_1077,N_14302,N_14284);
nand UO_1078 (O_1078,N_12725,N_13856);
nor UO_1079 (O_1079,N_12551,N_13616);
xnor UO_1080 (O_1080,N_14828,N_12605);
nor UO_1081 (O_1081,N_14420,N_13378);
and UO_1082 (O_1082,N_14802,N_13274);
or UO_1083 (O_1083,N_14536,N_12073);
nor UO_1084 (O_1084,N_12708,N_14896);
nand UO_1085 (O_1085,N_14194,N_12645);
nor UO_1086 (O_1086,N_14183,N_12982);
nand UO_1087 (O_1087,N_12472,N_12803);
or UO_1088 (O_1088,N_13573,N_14108);
nand UO_1089 (O_1089,N_14295,N_12761);
xor UO_1090 (O_1090,N_12895,N_12401);
or UO_1091 (O_1091,N_12046,N_14494);
or UO_1092 (O_1092,N_14103,N_14468);
nand UO_1093 (O_1093,N_14544,N_14044);
nand UO_1094 (O_1094,N_14470,N_12601);
xor UO_1095 (O_1095,N_13951,N_13186);
nor UO_1096 (O_1096,N_14853,N_13796);
or UO_1097 (O_1097,N_14728,N_14753);
nor UO_1098 (O_1098,N_13577,N_13868);
xnor UO_1099 (O_1099,N_12730,N_13471);
nor UO_1100 (O_1100,N_13992,N_14034);
and UO_1101 (O_1101,N_12176,N_13876);
or UO_1102 (O_1102,N_13688,N_12224);
nor UO_1103 (O_1103,N_12475,N_12509);
nand UO_1104 (O_1104,N_14622,N_13259);
or UO_1105 (O_1105,N_14546,N_13980);
or UO_1106 (O_1106,N_13950,N_13729);
nor UO_1107 (O_1107,N_14389,N_14218);
xnor UO_1108 (O_1108,N_13632,N_13122);
nand UO_1109 (O_1109,N_13370,N_14588);
nor UO_1110 (O_1110,N_14793,N_12506);
nor UO_1111 (O_1111,N_14996,N_12330);
nand UO_1112 (O_1112,N_14660,N_12764);
nand UO_1113 (O_1113,N_13698,N_13470);
and UO_1114 (O_1114,N_13364,N_13766);
nor UO_1115 (O_1115,N_13211,N_12842);
nor UO_1116 (O_1116,N_14540,N_13653);
nor UO_1117 (O_1117,N_13671,N_12150);
and UO_1118 (O_1118,N_14187,N_14111);
and UO_1119 (O_1119,N_14357,N_14010);
and UO_1120 (O_1120,N_12978,N_13008);
nand UO_1121 (O_1121,N_12641,N_14895);
and UO_1122 (O_1122,N_14923,N_13823);
nand UO_1123 (O_1123,N_14504,N_14849);
and UO_1124 (O_1124,N_13903,N_13634);
nor UO_1125 (O_1125,N_12901,N_13608);
nand UO_1126 (O_1126,N_12174,N_14709);
nand UO_1127 (O_1127,N_12447,N_14424);
nand UO_1128 (O_1128,N_12694,N_12181);
xor UO_1129 (O_1129,N_13496,N_14503);
or UO_1130 (O_1130,N_14306,N_13554);
or UO_1131 (O_1131,N_12069,N_13340);
and UO_1132 (O_1132,N_12661,N_13366);
nand UO_1133 (O_1133,N_12777,N_13375);
or UO_1134 (O_1134,N_14639,N_12245);
nor UO_1135 (O_1135,N_13241,N_14928);
nand UO_1136 (O_1136,N_13850,N_13215);
and UO_1137 (O_1137,N_13087,N_12955);
nand UO_1138 (O_1138,N_12055,N_13650);
and UO_1139 (O_1139,N_14861,N_14292);
or UO_1140 (O_1140,N_12663,N_12089);
and UO_1141 (O_1141,N_14609,N_12588);
or UO_1142 (O_1142,N_13321,N_14246);
and UO_1143 (O_1143,N_12022,N_13924);
or UO_1144 (O_1144,N_13024,N_12572);
nand UO_1145 (O_1145,N_14711,N_13756);
nor UO_1146 (O_1146,N_12061,N_14528);
or UO_1147 (O_1147,N_13659,N_12921);
nor UO_1148 (O_1148,N_14573,N_13304);
nand UO_1149 (O_1149,N_12171,N_14735);
or UO_1150 (O_1150,N_13808,N_12767);
xnor UO_1151 (O_1151,N_12918,N_12244);
nand UO_1152 (O_1152,N_14878,N_14515);
nor UO_1153 (O_1153,N_12947,N_13103);
nand UO_1154 (O_1154,N_12796,N_12238);
and UO_1155 (O_1155,N_13701,N_13781);
nor UO_1156 (O_1156,N_13320,N_14483);
nand UO_1157 (O_1157,N_14688,N_12102);
or UO_1158 (O_1158,N_13360,N_13034);
or UO_1159 (O_1159,N_13563,N_13021);
nand UO_1160 (O_1160,N_13537,N_13377);
or UO_1161 (O_1161,N_13057,N_14114);
nand UO_1162 (O_1162,N_13165,N_13742);
or UO_1163 (O_1163,N_13513,N_12228);
or UO_1164 (O_1164,N_13004,N_13206);
or UO_1165 (O_1165,N_12254,N_14984);
nor UO_1166 (O_1166,N_14412,N_14378);
or UO_1167 (O_1167,N_12404,N_14304);
nor UO_1168 (O_1168,N_12840,N_12284);
nand UO_1169 (O_1169,N_13303,N_12396);
and UO_1170 (O_1170,N_13770,N_12628);
nand UO_1171 (O_1171,N_12035,N_12132);
nand UO_1172 (O_1172,N_14596,N_12462);
nor UO_1173 (O_1173,N_14425,N_13192);
nand UO_1174 (O_1174,N_14170,N_13880);
nor UO_1175 (O_1175,N_12544,N_14463);
nand UO_1176 (O_1176,N_12989,N_12028);
or UO_1177 (O_1177,N_13743,N_13083);
or UO_1178 (O_1178,N_14050,N_12752);
nor UO_1179 (O_1179,N_13644,N_14535);
nor UO_1180 (O_1180,N_13600,N_12713);
or UO_1181 (O_1181,N_12274,N_12704);
and UO_1182 (O_1182,N_13146,N_12812);
and UO_1183 (O_1183,N_12934,N_13769);
and UO_1184 (O_1184,N_13778,N_12979);
xnor UO_1185 (O_1185,N_13568,N_12929);
nand UO_1186 (O_1186,N_13622,N_14426);
and UO_1187 (O_1187,N_13164,N_13683);
and UO_1188 (O_1188,N_13387,N_12819);
and UO_1189 (O_1189,N_13533,N_13069);
nor UO_1190 (O_1190,N_13060,N_14701);
and UO_1191 (O_1191,N_14449,N_13816);
nand UO_1192 (O_1192,N_13335,N_12732);
nor UO_1193 (O_1193,N_12346,N_13542);
nand UO_1194 (O_1194,N_12582,N_13225);
and UO_1195 (O_1195,N_13699,N_14210);
or UO_1196 (O_1196,N_14975,N_13812);
nand UO_1197 (O_1197,N_13852,N_12689);
nand UO_1198 (O_1198,N_12225,N_12523);
and UO_1199 (O_1199,N_14280,N_13809);
nand UO_1200 (O_1200,N_12697,N_14279);
and UO_1201 (O_1201,N_12999,N_12604);
nor UO_1202 (O_1202,N_13559,N_12315);
or UO_1203 (O_1203,N_12995,N_12164);
nand UO_1204 (O_1204,N_12505,N_14706);
or UO_1205 (O_1205,N_14576,N_12113);
or UO_1206 (O_1206,N_14817,N_12939);
xnor UO_1207 (O_1207,N_13269,N_13604);
and UO_1208 (O_1208,N_13184,N_13595);
nor UO_1209 (O_1209,N_12951,N_13395);
and UO_1210 (O_1210,N_14117,N_13895);
or UO_1211 (O_1211,N_13306,N_14960);
nor UO_1212 (O_1212,N_12286,N_14529);
nand UO_1213 (O_1213,N_12142,N_13258);
nor UO_1214 (O_1214,N_12157,N_14968);
nand UO_1215 (O_1215,N_12358,N_14264);
nor UO_1216 (O_1216,N_12650,N_13885);
and UO_1217 (O_1217,N_14784,N_12250);
nor UO_1218 (O_1218,N_13820,N_12426);
or UO_1219 (O_1219,N_14577,N_12410);
nand UO_1220 (O_1220,N_13849,N_12031);
nand UO_1221 (O_1221,N_13108,N_14702);
nor UO_1222 (O_1222,N_13877,N_14521);
or UO_1223 (O_1223,N_14258,N_14694);
and UO_1224 (O_1224,N_12363,N_14829);
and UO_1225 (O_1225,N_12298,N_13011);
or UO_1226 (O_1226,N_14951,N_12302);
nor UO_1227 (O_1227,N_14884,N_12524);
or UO_1228 (O_1228,N_13906,N_14517);
or UO_1229 (O_1229,N_12037,N_13613);
nor UO_1230 (O_1230,N_13359,N_14058);
nor UO_1231 (O_1231,N_13801,N_12272);
nand UO_1232 (O_1232,N_12620,N_14591);
or UO_1233 (O_1233,N_14514,N_12943);
or UO_1234 (O_1234,N_13204,N_14379);
nor UO_1235 (O_1235,N_14659,N_12307);
or UO_1236 (O_1236,N_14299,N_12632);
or UO_1237 (O_1237,N_12762,N_14270);
and UO_1238 (O_1238,N_13017,N_14181);
xnor UO_1239 (O_1239,N_12703,N_14749);
or UO_1240 (O_1240,N_14281,N_14524);
and UO_1241 (O_1241,N_14590,N_13427);
nor UO_1242 (O_1242,N_12128,N_14124);
or UO_1243 (O_1243,N_14774,N_13168);
and UO_1244 (O_1244,N_14238,N_14107);
and UO_1245 (O_1245,N_13564,N_12615);
and UO_1246 (O_1246,N_12124,N_13022);
nand UO_1247 (O_1247,N_12187,N_13928);
or UO_1248 (O_1248,N_13555,N_13583);
and UO_1249 (O_1249,N_14391,N_12959);
and UO_1250 (O_1250,N_14239,N_13367);
nand UO_1251 (O_1251,N_13058,N_14756);
nor UO_1252 (O_1252,N_12496,N_13112);
nor UO_1253 (O_1253,N_12519,N_12206);
nand UO_1254 (O_1254,N_12403,N_12637);
nor UO_1255 (O_1255,N_13944,N_14192);
or UO_1256 (O_1256,N_14430,N_13288);
or UO_1257 (O_1257,N_13198,N_13180);
nor UO_1258 (O_1258,N_12799,N_14116);
nor UO_1259 (O_1259,N_13411,N_12613);
nand UO_1260 (O_1260,N_12083,N_13107);
and UO_1261 (O_1261,N_13333,N_14600);
nor UO_1262 (O_1262,N_12498,N_13464);
nand UO_1263 (O_1263,N_14812,N_14318);
nor UO_1264 (O_1264,N_12515,N_13667);
or UO_1265 (O_1265,N_14824,N_12778);
or UO_1266 (O_1266,N_13463,N_14423);
and UO_1267 (O_1267,N_12992,N_12933);
nor UO_1268 (O_1268,N_12522,N_14835);
or UO_1269 (O_1269,N_14959,N_14763);
and UO_1270 (O_1270,N_13737,N_12753);
nand UO_1271 (O_1271,N_12863,N_14611);
nor UO_1272 (O_1272,N_13811,N_14670);
or UO_1273 (O_1273,N_14810,N_14628);
or UO_1274 (O_1274,N_14658,N_12531);
and UO_1275 (O_1275,N_12056,N_12104);
nand UO_1276 (O_1276,N_14921,N_14954);
nand UO_1277 (O_1277,N_14664,N_13806);
and UO_1278 (O_1278,N_13883,N_12377);
and UO_1279 (O_1279,N_12991,N_13218);
nand UO_1280 (O_1280,N_12785,N_12341);
nor UO_1281 (O_1281,N_12463,N_12313);
or UO_1282 (O_1282,N_12685,N_13979);
or UO_1283 (O_1283,N_13014,N_12562);
or UO_1284 (O_1284,N_14553,N_14175);
nand UO_1285 (O_1285,N_12837,N_14775);
or UO_1286 (O_1286,N_12838,N_14522);
and UO_1287 (O_1287,N_14205,N_14747);
nand UO_1288 (O_1288,N_13356,N_12937);
nand UO_1289 (O_1289,N_12851,N_14007);
nand UO_1290 (O_1290,N_12736,N_13594);
and UO_1291 (O_1291,N_13260,N_12894);
nand UO_1292 (O_1292,N_12649,N_14093);
nand UO_1293 (O_1293,N_12329,N_14724);
or UO_1294 (O_1294,N_13703,N_14859);
nand UO_1295 (O_1295,N_12278,N_12476);
or UO_1296 (O_1296,N_13635,N_14338);
nor UO_1297 (O_1297,N_13726,N_14395);
and UO_1298 (O_1298,N_12830,N_14847);
or UO_1299 (O_1299,N_14972,N_14310);
nand UO_1300 (O_1300,N_13503,N_14874);
or UO_1301 (O_1301,N_13584,N_13128);
and UO_1302 (O_1302,N_14365,N_13662);
nand UO_1303 (O_1303,N_14245,N_13909);
or UO_1304 (O_1304,N_14364,N_13380);
nor UO_1305 (O_1305,N_13565,N_13273);
nand UO_1306 (O_1306,N_14469,N_14024);
nand UO_1307 (O_1307,N_13501,N_14064);
and UO_1308 (O_1308,N_13182,N_13373);
and UO_1309 (O_1309,N_14168,N_12848);
or UO_1310 (O_1310,N_13005,N_14496);
and UO_1311 (O_1311,N_14369,N_12338);
xor UO_1312 (O_1312,N_14290,N_13779);
nand UO_1313 (O_1313,N_12928,N_13237);
nor UO_1314 (O_1314,N_14635,N_14129);
nand UO_1315 (O_1315,N_14612,N_14672);
nand UO_1316 (O_1316,N_12199,N_12627);
nor UO_1317 (O_1317,N_12458,N_13073);
or UO_1318 (O_1318,N_14132,N_13892);
nor UO_1319 (O_1319,N_12062,N_14437);
nand UO_1320 (O_1320,N_12425,N_12793);
and UO_1321 (O_1321,N_12465,N_14786);
and UO_1322 (O_1322,N_12794,N_14799);
nand UO_1323 (O_1323,N_12633,N_12654);
and UO_1324 (O_1324,N_13953,N_12577);
nand UO_1325 (O_1325,N_13499,N_12686);
or UO_1326 (O_1326,N_14358,N_14650);
or UO_1327 (O_1327,N_13828,N_14741);
or UO_1328 (O_1328,N_14925,N_12492);
nor UO_1329 (O_1329,N_13942,N_13341);
nand UO_1330 (O_1330,N_12482,N_13519);
nand UO_1331 (O_1331,N_14171,N_14363);
nor UO_1332 (O_1332,N_13744,N_14027);
or UO_1333 (O_1333,N_13725,N_14814);
nand UO_1334 (O_1334,N_13188,N_12747);
and UO_1335 (O_1335,N_14994,N_13392);
nor UO_1336 (O_1336,N_13507,N_14440);
and UO_1337 (O_1337,N_14726,N_13117);
nand UO_1338 (O_1338,N_13150,N_14532);
or UO_1339 (O_1339,N_12495,N_14574);
and UO_1340 (O_1340,N_13964,N_14848);
nand UO_1341 (O_1341,N_14055,N_13189);
or UO_1342 (O_1342,N_14105,N_12347);
and UO_1343 (O_1343,N_12962,N_13597);
nand UO_1344 (O_1344,N_12248,N_14184);
nand UO_1345 (O_1345,N_14283,N_12276);
nand UO_1346 (O_1346,N_13385,N_13426);
nor UO_1347 (O_1347,N_12774,N_13031);
or UO_1348 (O_1348,N_14041,N_12914);
nor UO_1349 (O_1349,N_14394,N_12670);
or UO_1350 (O_1350,N_14174,N_14926);
or UO_1351 (O_1351,N_14564,N_12948);
and UO_1352 (O_1352,N_12773,N_14499);
and UO_1353 (O_1353,N_14534,N_12032);
nand UO_1354 (O_1354,N_13361,N_14703);
or UO_1355 (O_1355,N_14333,N_14748);
and UO_1356 (O_1356,N_12765,N_13971);
or UO_1357 (O_1357,N_14118,N_13920);
nand UO_1358 (O_1358,N_14953,N_12800);
or UO_1359 (O_1359,N_12070,N_12234);
or UO_1360 (O_1360,N_14126,N_14583);
and UO_1361 (O_1361,N_14054,N_12379);
and UO_1362 (O_1362,N_14643,N_12802);
or UO_1363 (O_1363,N_14653,N_13299);
or UO_1364 (O_1364,N_14989,N_14272);
nor UO_1365 (O_1365,N_12213,N_12414);
nand UO_1366 (O_1366,N_13293,N_14965);
or UO_1367 (O_1367,N_14991,N_12297);
nor UO_1368 (O_1368,N_12944,N_13253);
nand UO_1369 (O_1369,N_13708,N_14898);
or UO_1370 (O_1370,N_13473,N_12443);
nand UO_1371 (O_1371,N_13601,N_14419);
or UO_1372 (O_1372,N_12135,N_13318);
or UO_1373 (O_1373,N_14787,N_12998);
or UO_1374 (O_1374,N_12909,N_14138);
nor UO_1375 (O_1375,N_12391,N_14945);
and UO_1376 (O_1376,N_12431,N_13185);
or UO_1377 (O_1377,N_12205,N_13693);
or UO_1378 (O_1378,N_14322,N_14226);
or UO_1379 (O_1379,N_14892,N_14764);
nor UO_1380 (O_1380,N_13922,N_13623);
and UO_1381 (O_1381,N_13578,N_14610);
nand UO_1382 (O_1382,N_13521,N_14738);
and UO_1383 (O_1383,N_13059,N_12717);
and UO_1384 (O_1384,N_12222,N_13115);
nand UO_1385 (O_1385,N_13690,N_14455);
nor UO_1386 (O_1386,N_12487,N_14308);
nor UO_1387 (O_1387,N_14130,N_12818);
nor UO_1388 (O_1388,N_14624,N_14134);
or UO_1389 (O_1389,N_12140,N_13120);
nor UO_1390 (O_1390,N_12311,N_13854);
or UO_1391 (O_1391,N_13238,N_12599);
nor UO_1392 (O_1392,N_12439,N_13443);
nand UO_1393 (O_1393,N_12906,N_13720);
and UO_1394 (O_1394,N_12188,N_12219);
xnor UO_1395 (O_1395,N_12675,N_14434);
or UO_1396 (O_1396,N_12247,N_14486);
or UO_1397 (O_1397,N_13991,N_12855);
and UO_1398 (O_1398,N_12373,N_14841);
nor UO_1399 (O_1399,N_13347,N_14554);
nor UO_1400 (O_1400,N_13118,N_12266);
nor UO_1401 (O_1401,N_13633,N_14387);
and UO_1402 (O_1402,N_13157,N_13676);
nand UO_1403 (O_1403,N_13498,N_14182);
or UO_1404 (O_1404,N_13628,N_13541);
nor UO_1405 (O_1405,N_12922,N_14915);
and UO_1406 (O_1406,N_13767,N_13137);
nand UO_1407 (O_1407,N_13355,N_12370);
nor UO_1408 (O_1408,N_13962,N_12502);
and UO_1409 (O_1409,N_12249,N_14478);
nor UO_1410 (O_1410,N_13863,N_12880);
nand UO_1411 (O_1411,N_14647,N_14507);
and UO_1412 (O_1412,N_12743,N_14935);
nand UO_1413 (O_1413,N_12160,N_14002);
or UO_1414 (O_1414,N_12212,N_14207);
nor UO_1415 (O_1415,N_12521,N_14737);
and UO_1416 (O_1416,N_14454,N_14723);
or UO_1417 (O_1417,N_13044,N_14868);
nand UO_1418 (O_1418,N_13265,N_12875);
xor UO_1419 (O_1419,N_12067,N_13401);
xnor UO_1420 (O_1420,N_14966,N_14414);
and UO_1421 (O_1421,N_13844,N_13125);
or UO_1422 (O_1422,N_14450,N_12427);
nand UO_1423 (O_1423,N_12782,N_14906);
or UO_1424 (O_1424,N_14619,N_12619);
nor UO_1425 (O_1425,N_14362,N_13158);
nand UO_1426 (O_1426,N_12019,N_14755);
nor UO_1427 (O_1427,N_14796,N_13313);
nand UO_1428 (O_1428,N_14408,N_14731);
nand UO_1429 (O_1429,N_13196,N_14883);
and UO_1430 (O_1430,N_14480,N_13792);
nand UO_1431 (O_1431,N_14899,N_12350);
and UO_1432 (O_1432,N_12647,N_12116);
nor UO_1433 (O_1433,N_14623,N_13930);
and UO_1434 (O_1434,N_12564,N_14110);
or UO_1435 (O_1435,N_14750,N_14950);
or UO_1436 (O_1436,N_13413,N_12175);
nor UO_1437 (O_1437,N_13747,N_13409);
and UO_1438 (O_1438,N_14180,N_14461);
nor UO_1439 (O_1439,N_13859,N_14048);
or UO_1440 (O_1440,N_13631,N_14260);
nand UO_1441 (O_1441,N_12540,N_14082);
nor UO_1442 (O_1442,N_14592,N_14474);
xnor UO_1443 (O_1443,N_13666,N_13092);
nor UO_1444 (O_1444,N_14934,N_13296);
or UO_1445 (O_1445,N_14839,N_13975);
or UO_1446 (O_1446,N_13824,N_12640);
and UO_1447 (O_1447,N_13027,N_13170);
and UO_1448 (O_1448,N_12728,N_13665);
nand UO_1449 (O_1449,N_13091,N_12434);
nor UO_1450 (O_1450,N_14195,N_14078);
and UO_1451 (O_1451,N_12756,N_14242);
nor UO_1452 (O_1452,N_13875,N_12422);
nor UO_1453 (O_1453,N_13506,N_14417);
or UO_1454 (O_1454,N_13423,N_14303);
and UO_1455 (O_1455,N_12445,N_12216);
nor UO_1456 (O_1456,N_12155,N_13030);
or UO_1457 (O_1457,N_13223,N_13822);
nand UO_1458 (O_1458,N_14092,N_12256);
and UO_1459 (O_1459,N_13557,N_14477);
nand UO_1460 (O_1460,N_12566,N_12935);
nand UO_1461 (O_1461,N_14340,N_13045);
and UO_1462 (O_1462,N_14352,N_12532);
or UO_1463 (O_1463,N_13174,N_12537);
or UO_1464 (O_1464,N_12780,N_13791);
or UO_1465 (O_1465,N_12211,N_14642);
or UO_1466 (O_1466,N_14211,N_14343);
nor UO_1467 (O_1467,N_14502,N_12467);
nor UO_1468 (O_1468,N_14683,N_13607);
or UO_1469 (O_1469,N_13986,N_12133);
xnor UO_1470 (O_1470,N_13074,N_13680);
nor UO_1471 (O_1471,N_12390,N_12405);
or UO_1472 (O_1472,N_13795,N_12611);
nor UO_1473 (O_1473,N_13978,N_14981);
nor UO_1474 (O_1474,N_13231,N_14313);
and UO_1475 (O_1475,N_12100,N_12010);
nor UO_1476 (O_1476,N_13284,N_13090);
nor UO_1477 (O_1477,N_13428,N_14025);
nor UO_1478 (O_1478,N_12107,N_14595);
or UO_1479 (O_1479,N_12739,N_13988);
nand UO_1480 (O_1480,N_12295,N_12865);
or UO_1481 (O_1481,N_14880,N_13420);
or UO_1482 (O_1482,N_12098,N_14613);
nor UO_1483 (O_1483,N_12655,N_14916);
nand UO_1484 (O_1484,N_12823,N_13277);
or UO_1485 (O_1485,N_14986,N_13230);
xnor UO_1486 (O_1486,N_14593,N_14850);
nand UO_1487 (O_1487,N_13493,N_13510);
nor UO_1488 (O_1488,N_14431,N_13606);
nand UO_1489 (O_1489,N_14931,N_13358);
and UO_1490 (O_1490,N_14028,N_13337);
and UO_1491 (O_1491,N_13900,N_14346);
nand UO_1492 (O_1492,N_14948,N_13545);
nor UO_1493 (O_1493,N_12536,N_14788);
or UO_1494 (O_1494,N_14720,N_12657);
nor UO_1495 (O_1495,N_12380,N_13453);
or UO_1496 (O_1496,N_13592,N_13905);
nand UO_1497 (O_1497,N_14962,N_14550);
nor UO_1498 (O_1498,N_14462,N_13588);
nand UO_1499 (O_1499,N_14235,N_13888);
and UO_1500 (O_1500,N_13788,N_12516);
and UO_1501 (O_1501,N_12307,N_14690);
or UO_1502 (O_1502,N_14211,N_12266);
and UO_1503 (O_1503,N_13934,N_12146);
and UO_1504 (O_1504,N_13971,N_13803);
or UO_1505 (O_1505,N_14545,N_14633);
nor UO_1506 (O_1506,N_13536,N_14274);
and UO_1507 (O_1507,N_12285,N_12924);
xnor UO_1508 (O_1508,N_12681,N_12550);
nand UO_1509 (O_1509,N_14485,N_13309);
and UO_1510 (O_1510,N_14457,N_13757);
xnor UO_1511 (O_1511,N_12186,N_13542);
nor UO_1512 (O_1512,N_14984,N_14369);
nand UO_1513 (O_1513,N_13194,N_12140);
nand UO_1514 (O_1514,N_14959,N_13233);
or UO_1515 (O_1515,N_14689,N_13773);
or UO_1516 (O_1516,N_13605,N_12597);
nand UO_1517 (O_1517,N_13668,N_12117);
nand UO_1518 (O_1518,N_12821,N_13391);
nand UO_1519 (O_1519,N_14568,N_14874);
nor UO_1520 (O_1520,N_13231,N_13125);
and UO_1521 (O_1521,N_12505,N_14780);
nand UO_1522 (O_1522,N_13656,N_14184);
or UO_1523 (O_1523,N_13356,N_14475);
nand UO_1524 (O_1524,N_14276,N_14079);
or UO_1525 (O_1525,N_13078,N_12331);
or UO_1526 (O_1526,N_14188,N_13635);
xnor UO_1527 (O_1527,N_12009,N_13954);
nor UO_1528 (O_1528,N_12156,N_12026);
and UO_1529 (O_1529,N_13252,N_13963);
nand UO_1530 (O_1530,N_14976,N_12083);
nand UO_1531 (O_1531,N_13417,N_13554);
nand UO_1532 (O_1532,N_14942,N_14485);
nand UO_1533 (O_1533,N_13103,N_12186);
nor UO_1534 (O_1534,N_13363,N_13985);
nand UO_1535 (O_1535,N_13741,N_14898);
and UO_1536 (O_1536,N_14626,N_14855);
or UO_1537 (O_1537,N_13081,N_12720);
and UO_1538 (O_1538,N_13629,N_14322);
and UO_1539 (O_1539,N_12451,N_13682);
nand UO_1540 (O_1540,N_12250,N_14453);
nor UO_1541 (O_1541,N_13615,N_12086);
and UO_1542 (O_1542,N_12153,N_13953);
nor UO_1543 (O_1543,N_14606,N_14585);
and UO_1544 (O_1544,N_12978,N_14433);
or UO_1545 (O_1545,N_13808,N_13378);
nor UO_1546 (O_1546,N_12224,N_13535);
nor UO_1547 (O_1547,N_13604,N_12787);
nand UO_1548 (O_1548,N_14184,N_14629);
nand UO_1549 (O_1549,N_12137,N_14917);
xnor UO_1550 (O_1550,N_12843,N_14971);
nor UO_1551 (O_1551,N_13619,N_14634);
nand UO_1552 (O_1552,N_14174,N_12405);
nand UO_1553 (O_1553,N_12758,N_13091);
nand UO_1554 (O_1554,N_14516,N_12290);
nor UO_1555 (O_1555,N_13181,N_13241);
and UO_1556 (O_1556,N_13973,N_12779);
xnor UO_1557 (O_1557,N_13592,N_14347);
nor UO_1558 (O_1558,N_13851,N_13509);
xor UO_1559 (O_1559,N_12263,N_13332);
or UO_1560 (O_1560,N_13605,N_13932);
nor UO_1561 (O_1561,N_14111,N_14541);
nor UO_1562 (O_1562,N_13454,N_13316);
nand UO_1563 (O_1563,N_13522,N_12897);
nor UO_1564 (O_1564,N_14767,N_14008);
and UO_1565 (O_1565,N_13285,N_14166);
and UO_1566 (O_1566,N_14845,N_12084);
and UO_1567 (O_1567,N_13761,N_13347);
or UO_1568 (O_1568,N_12270,N_12852);
nor UO_1569 (O_1569,N_12401,N_12619);
and UO_1570 (O_1570,N_13383,N_14436);
and UO_1571 (O_1571,N_14606,N_12657);
nand UO_1572 (O_1572,N_12180,N_14327);
nor UO_1573 (O_1573,N_13530,N_13796);
and UO_1574 (O_1574,N_14998,N_13575);
or UO_1575 (O_1575,N_12537,N_13938);
or UO_1576 (O_1576,N_14848,N_12357);
or UO_1577 (O_1577,N_13827,N_14224);
nand UO_1578 (O_1578,N_14113,N_14404);
and UO_1579 (O_1579,N_12817,N_12703);
and UO_1580 (O_1580,N_13479,N_14425);
nor UO_1581 (O_1581,N_12446,N_14819);
nor UO_1582 (O_1582,N_12293,N_12891);
and UO_1583 (O_1583,N_12197,N_14681);
and UO_1584 (O_1584,N_12439,N_12028);
or UO_1585 (O_1585,N_12568,N_12777);
or UO_1586 (O_1586,N_13274,N_13335);
or UO_1587 (O_1587,N_14098,N_14730);
nor UO_1588 (O_1588,N_13118,N_12272);
or UO_1589 (O_1589,N_14216,N_13466);
nor UO_1590 (O_1590,N_12682,N_13467);
nor UO_1591 (O_1591,N_14026,N_12523);
nor UO_1592 (O_1592,N_14955,N_13860);
xor UO_1593 (O_1593,N_12676,N_14941);
nor UO_1594 (O_1594,N_14793,N_13517);
nand UO_1595 (O_1595,N_12914,N_14057);
or UO_1596 (O_1596,N_14770,N_14703);
nand UO_1597 (O_1597,N_12541,N_13153);
nor UO_1598 (O_1598,N_14991,N_14911);
or UO_1599 (O_1599,N_13212,N_13142);
or UO_1600 (O_1600,N_12401,N_13572);
nor UO_1601 (O_1601,N_13641,N_14718);
and UO_1602 (O_1602,N_14947,N_13131);
nand UO_1603 (O_1603,N_12124,N_13179);
or UO_1604 (O_1604,N_12703,N_12416);
nor UO_1605 (O_1605,N_13315,N_12647);
and UO_1606 (O_1606,N_13636,N_12720);
and UO_1607 (O_1607,N_14892,N_13683);
or UO_1608 (O_1608,N_13608,N_13271);
nand UO_1609 (O_1609,N_14518,N_13472);
and UO_1610 (O_1610,N_14917,N_12630);
xnor UO_1611 (O_1611,N_12671,N_12660);
and UO_1612 (O_1612,N_12782,N_12814);
nand UO_1613 (O_1613,N_13721,N_13633);
and UO_1614 (O_1614,N_13439,N_13476);
nor UO_1615 (O_1615,N_12606,N_13442);
or UO_1616 (O_1616,N_13303,N_12156);
nand UO_1617 (O_1617,N_12170,N_14629);
and UO_1618 (O_1618,N_13728,N_13165);
nand UO_1619 (O_1619,N_14571,N_13555);
and UO_1620 (O_1620,N_12391,N_12777);
and UO_1621 (O_1621,N_12363,N_13030);
nand UO_1622 (O_1622,N_13435,N_12614);
and UO_1623 (O_1623,N_14105,N_14283);
nand UO_1624 (O_1624,N_12675,N_13779);
nor UO_1625 (O_1625,N_14350,N_12457);
nand UO_1626 (O_1626,N_14822,N_12976);
nor UO_1627 (O_1627,N_14539,N_13851);
and UO_1628 (O_1628,N_12801,N_13332);
and UO_1629 (O_1629,N_13730,N_13234);
nand UO_1630 (O_1630,N_14600,N_14716);
and UO_1631 (O_1631,N_13036,N_14697);
nor UO_1632 (O_1632,N_14639,N_13986);
nor UO_1633 (O_1633,N_14423,N_12067);
nor UO_1634 (O_1634,N_14014,N_12740);
nand UO_1635 (O_1635,N_13541,N_14464);
and UO_1636 (O_1636,N_12857,N_13695);
and UO_1637 (O_1637,N_13505,N_13148);
or UO_1638 (O_1638,N_14364,N_13040);
or UO_1639 (O_1639,N_13004,N_12992);
nand UO_1640 (O_1640,N_13902,N_12357);
nand UO_1641 (O_1641,N_13867,N_14400);
nand UO_1642 (O_1642,N_12294,N_13512);
and UO_1643 (O_1643,N_13587,N_14290);
nor UO_1644 (O_1644,N_14122,N_13314);
or UO_1645 (O_1645,N_14332,N_12567);
nor UO_1646 (O_1646,N_12625,N_13770);
and UO_1647 (O_1647,N_12429,N_13769);
nor UO_1648 (O_1648,N_13311,N_14913);
nand UO_1649 (O_1649,N_13942,N_12791);
and UO_1650 (O_1650,N_12098,N_12132);
nor UO_1651 (O_1651,N_12407,N_14349);
and UO_1652 (O_1652,N_12641,N_12175);
nor UO_1653 (O_1653,N_12706,N_13751);
nor UO_1654 (O_1654,N_12722,N_12091);
nor UO_1655 (O_1655,N_14841,N_12604);
nor UO_1656 (O_1656,N_12756,N_14691);
or UO_1657 (O_1657,N_14372,N_12104);
and UO_1658 (O_1658,N_14825,N_14881);
and UO_1659 (O_1659,N_12995,N_12796);
and UO_1660 (O_1660,N_13571,N_12011);
and UO_1661 (O_1661,N_12622,N_14109);
nand UO_1662 (O_1662,N_13452,N_14176);
and UO_1663 (O_1663,N_12331,N_13414);
or UO_1664 (O_1664,N_12433,N_14769);
or UO_1665 (O_1665,N_13126,N_12369);
nand UO_1666 (O_1666,N_14543,N_12681);
nand UO_1667 (O_1667,N_12549,N_13916);
nand UO_1668 (O_1668,N_12480,N_12577);
nor UO_1669 (O_1669,N_12132,N_13023);
nand UO_1670 (O_1670,N_13137,N_14154);
nand UO_1671 (O_1671,N_13554,N_12791);
and UO_1672 (O_1672,N_14217,N_12276);
nand UO_1673 (O_1673,N_13258,N_13519);
nor UO_1674 (O_1674,N_14586,N_13215);
and UO_1675 (O_1675,N_14568,N_14505);
nor UO_1676 (O_1676,N_12322,N_14511);
and UO_1677 (O_1677,N_12087,N_13734);
or UO_1678 (O_1678,N_12112,N_14914);
nor UO_1679 (O_1679,N_12440,N_12694);
and UO_1680 (O_1680,N_14949,N_13456);
nand UO_1681 (O_1681,N_12597,N_13165);
nor UO_1682 (O_1682,N_14662,N_13237);
nand UO_1683 (O_1683,N_13405,N_12297);
and UO_1684 (O_1684,N_14427,N_14056);
and UO_1685 (O_1685,N_13677,N_14659);
nor UO_1686 (O_1686,N_14231,N_14995);
and UO_1687 (O_1687,N_13559,N_14002);
and UO_1688 (O_1688,N_13121,N_12151);
and UO_1689 (O_1689,N_12902,N_14238);
and UO_1690 (O_1690,N_14020,N_14500);
nand UO_1691 (O_1691,N_12323,N_13678);
nor UO_1692 (O_1692,N_13223,N_14282);
or UO_1693 (O_1693,N_14095,N_13249);
xor UO_1694 (O_1694,N_13429,N_13027);
or UO_1695 (O_1695,N_13461,N_13701);
and UO_1696 (O_1696,N_12152,N_14295);
nor UO_1697 (O_1697,N_14832,N_13196);
nor UO_1698 (O_1698,N_14913,N_14559);
and UO_1699 (O_1699,N_14883,N_12304);
and UO_1700 (O_1700,N_13274,N_13961);
and UO_1701 (O_1701,N_12615,N_14738);
and UO_1702 (O_1702,N_13586,N_14723);
and UO_1703 (O_1703,N_14750,N_13661);
or UO_1704 (O_1704,N_14510,N_12967);
and UO_1705 (O_1705,N_13325,N_12844);
or UO_1706 (O_1706,N_12694,N_12483);
and UO_1707 (O_1707,N_14961,N_13064);
nor UO_1708 (O_1708,N_13738,N_13483);
nand UO_1709 (O_1709,N_14451,N_13420);
and UO_1710 (O_1710,N_13529,N_13219);
nor UO_1711 (O_1711,N_12469,N_13995);
and UO_1712 (O_1712,N_14082,N_12164);
or UO_1713 (O_1713,N_13619,N_12654);
or UO_1714 (O_1714,N_13895,N_12925);
nand UO_1715 (O_1715,N_14666,N_12579);
and UO_1716 (O_1716,N_14907,N_12747);
and UO_1717 (O_1717,N_14909,N_14233);
or UO_1718 (O_1718,N_14716,N_13557);
nor UO_1719 (O_1719,N_12766,N_14290);
or UO_1720 (O_1720,N_12441,N_12130);
and UO_1721 (O_1721,N_13228,N_13099);
or UO_1722 (O_1722,N_14797,N_14364);
nor UO_1723 (O_1723,N_14576,N_12294);
nand UO_1724 (O_1724,N_13776,N_14214);
nand UO_1725 (O_1725,N_12769,N_14616);
nand UO_1726 (O_1726,N_12247,N_14730);
nor UO_1727 (O_1727,N_12894,N_14552);
nand UO_1728 (O_1728,N_12379,N_13781);
nand UO_1729 (O_1729,N_13525,N_13422);
or UO_1730 (O_1730,N_12673,N_12808);
or UO_1731 (O_1731,N_12828,N_12815);
nor UO_1732 (O_1732,N_13863,N_12425);
and UO_1733 (O_1733,N_13037,N_13212);
and UO_1734 (O_1734,N_14816,N_14448);
nand UO_1735 (O_1735,N_12828,N_13392);
nor UO_1736 (O_1736,N_13754,N_12018);
nand UO_1737 (O_1737,N_14135,N_13901);
or UO_1738 (O_1738,N_13257,N_14339);
and UO_1739 (O_1739,N_12102,N_13043);
nand UO_1740 (O_1740,N_14880,N_13374);
nor UO_1741 (O_1741,N_13908,N_13646);
or UO_1742 (O_1742,N_12628,N_14538);
nor UO_1743 (O_1743,N_14964,N_12704);
or UO_1744 (O_1744,N_12320,N_12125);
nand UO_1745 (O_1745,N_13631,N_12393);
and UO_1746 (O_1746,N_14076,N_12744);
nor UO_1747 (O_1747,N_13626,N_13321);
nand UO_1748 (O_1748,N_12087,N_12655);
or UO_1749 (O_1749,N_12361,N_13855);
or UO_1750 (O_1750,N_13408,N_12799);
or UO_1751 (O_1751,N_14819,N_13480);
nor UO_1752 (O_1752,N_14095,N_14535);
xnor UO_1753 (O_1753,N_12192,N_13001);
or UO_1754 (O_1754,N_12111,N_13997);
nand UO_1755 (O_1755,N_12199,N_12310);
nor UO_1756 (O_1756,N_12561,N_13400);
or UO_1757 (O_1757,N_12170,N_13882);
nand UO_1758 (O_1758,N_12182,N_14924);
and UO_1759 (O_1759,N_13105,N_12842);
or UO_1760 (O_1760,N_14055,N_12881);
and UO_1761 (O_1761,N_13483,N_12357);
and UO_1762 (O_1762,N_14687,N_12703);
and UO_1763 (O_1763,N_13937,N_14294);
nor UO_1764 (O_1764,N_13010,N_13948);
and UO_1765 (O_1765,N_12515,N_14213);
nor UO_1766 (O_1766,N_13141,N_14163);
or UO_1767 (O_1767,N_14446,N_12409);
nor UO_1768 (O_1768,N_12066,N_13377);
and UO_1769 (O_1769,N_12566,N_14168);
nor UO_1770 (O_1770,N_12021,N_14606);
nor UO_1771 (O_1771,N_13845,N_12468);
or UO_1772 (O_1772,N_13370,N_14734);
nor UO_1773 (O_1773,N_13876,N_12737);
and UO_1774 (O_1774,N_14655,N_14729);
or UO_1775 (O_1775,N_12656,N_12403);
or UO_1776 (O_1776,N_13307,N_13643);
and UO_1777 (O_1777,N_13483,N_13539);
and UO_1778 (O_1778,N_13697,N_14661);
xor UO_1779 (O_1779,N_12972,N_13753);
nor UO_1780 (O_1780,N_12213,N_13765);
nand UO_1781 (O_1781,N_14081,N_14697);
nor UO_1782 (O_1782,N_14899,N_14825);
and UO_1783 (O_1783,N_12671,N_12254);
nand UO_1784 (O_1784,N_12930,N_14267);
xor UO_1785 (O_1785,N_13479,N_12988);
or UO_1786 (O_1786,N_14558,N_13924);
nor UO_1787 (O_1787,N_13325,N_12189);
nand UO_1788 (O_1788,N_14353,N_14117);
nor UO_1789 (O_1789,N_12958,N_12936);
nor UO_1790 (O_1790,N_12760,N_12362);
nor UO_1791 (O_1791,N_14378,N_14898);
and UO_1792 (O_1792,N_13645,N_12795);
nand UO_1793 (O_1793,N_12612,N_12743);
and UO_1794 (O_1794,N_12598,N_13770);
or UO_1795 (O_1795,N_12652,N_13449);
nand UO_1796 (O_1796,N_13926,N_12882);
and UO_1797 (O_1797,N_14028,N_14933);
nor UO_1798 (O_1798,N_14952,N_14600);
or UO_1799 (O_1799,N_12118,N_13552);
or UO_1800 (O_1800,N_14908,N_13436);
nor UO_1801 (O_1801,N_12945,N_14531);
and UO_1802 (O_1802,N_14408,N_12605);
nand UO_1803 (O_1803,N_13563,N_13133);
and UO_1804 (O_1804,N_12501,N_12935);
nand UO_1805 (O_1805,N_14752,N_13477);
nand UO_1806 (O_1806,N_14720,N_13094);
xor UO_1807 (O_1807,N_14050,N_13577);
nand UO_1808 (O_1808,N_12497,N_13634);
nand UO_1809 (O_1809,N_14731,N_13377);
or UO_1810 (O_1810,N_13197,N_13643);
and UO_1811 (O_1811,N_13854,N_13565);
or UO_1812 (O_1812,N_12207,N_12750);
nand UO_1813 (O_1813,N_12121,N_13301);
or UO_1814 (O_1814,N_14738,N_13927);
nand UO_1815 (O_1815,N_14832,N_13107);
and UO_1816 (O_1816,N_12242,N_14273);
or UO_1817 (O_1817,N_14638,N_12889);
and UO_1818 (O_1818,N_13455,N_12709);
nand UO_1819 (O_1819,N_13924,N_14239);
nor UO_1820 (O_1820,N_13861,N_13367);
and UO_1821 (O_1821,N_12983,N_13164);
or UO_1822 (O_1822,N_13489,N_13431);
nor UO_1823 (O_1823,N_14481,N_13113);
and UO_1824 (O_1824,N_14168,N_14268);
or UO_1825 (O_1825,N_13581,N_14725);
or UO_1826 (O_1826,N_12226,N_12165);
nand UO_1827 (O_1827,N_12995,N_14012);
nand UO_1828 (O_1828,N_14715,N_14493);
and UO_1829 (O_1829,N_14254,N_13008);
and UO_1830 (O_1830,N_14749,N_12767);
and UO_1831 (O_1831,N_13587,N_14466);
nand UO_1832 (O_1832,N_13870,N_14140);
or UO_1833 (O_1833,N_13626,N_12783);
nand UO_1834 (O_1834,N_12322,N_14084);
and UO_1835 (O_1835,N_14147,N_14642);
or UO_1836 (O_1836,N_14891,N_13819);
nor UO_1837 (O_1837,N_13018,N_12578);
nand UO_1838 (O_1838,N_13868,N_14447);
or UO_1839 (O_1839,N_12831,N_14334);
xor UO_1840 (O_1840,N_12674,N_13492);
nand UO_1841 (O_1841,N_14218,N_14873);
and UO_1842 (O_1842,N_14425,N_13413);
or UO_1843 (O_1843,N_14385,N_14703);
or UO_1844 (O_1844,N_14166,N_14635);
xnor UO_1845 (O_1845,N_12460,N_12259);
and UO_1846 (O_1846,N_14203,N_12348);
nand UO_1847 (O_1847,N_14375,N_12858);
nand UO_1848 (O_1848,N_12954,N_12530);
and UO_1849 (O_1849,N_14215,N_14912);
nand UO_1850 (O_1850,N_13061,N_12634);
nor UO_1851 (O_1851,N_14337,N_13825);
nand UO_1852 (O_1852,N_14895,N_12200);
nand UO_1853 (O_1853,N_14297,N_13901);
or UO_1854 (O_1854,N_13967,N_12525);
and UO_1855 (O_1855,N_13868,N_12335);
nand UO_1856 (O_1856,N_12103,N_14766);
and UO_1857 (O_1857,N_13271,N_14246);
and UO_1858 (O_1858,N_13014,N_14086);
and UO_1859 (O_1859,N_13470,N_13650);
and UO_1860 (O_1860,N_13092,N_12797);
or UO_1861 (O_1861,N_14113,N_12844);
nor UO_1862 (O_1862,N_12129,N_12654);
and UO_1863 (O_1863,N_13665,N_13624);
nor UO_1864 (O_1864,N_12355,N_14478);
or UO_1865 (O_1865,N_12931,N_14622);
or UO_1866 (O_1866,N_12134,N_13810);
and UO_1867 (O_1867,N_12167,N_14806);
and UO_1868 (O_1868,N_14183,N_12892);
nand UO_1869 (O_1869,N_14687,N_13646);
and UO_1870 (O_1870,N_12467,N_14573);
nor UO_1871 (O_1871,N_12895,N_13364);
and UO_1872 (O_1872,N_12168,N_12888);
and UO_1873 (O_1873,N_13207,N_14929);
and UO_1874 (O_1874,N_13721,N_12378);
nor UO_1875 (O_1875,N_14634,N_13859);
nor UO_1876 (O_1876,N_12791,N_13581);
and UO_1877 (O_1877,N_13874,N_12244);
and UO_1878 (O_1878,N_12941,N_14656);
and UO_1879 (O_1879,N_14599,N_14875);
xor UO_1880 (O_1880,N_14932,N_13269);
xor UO_1881 (O_1881,N_12452,N_14306);
nand UO_1882 (O_1882,N_13074,N_14254);
nand UO_1883 (O_1883,N_12441,N_12979);
and UO_1884 (O_1884,N_12957,N_12508);
nand UO_1885 (O_1885,N_12273,N_13871);
nor UO_1886 (O_1886,N_13365,N_13524);
nand UO_1887 (O_1887,N_13227,N_13443);
nand UO_1888 (O_1888,N_12628,N_13578);
or UO_1889 (O_1889,N_13988,N_13545);
nand UO_1890 (O_1890,N_14677,N_14905);
or UO_1891 (O_1891,N_12896,N_14062);
and UO_1892 (O_1892,N_14304,N_14058);
or UO_1893 (O_1893,N_14294,N_12664);
or UO_1894 (O_1894,N_13523,N_12347);
nor UO_1895 (O_1895,N_13769,N_14609);
xor UO_1896 (O_1896,N_14377,N_12687);
or UO_1897 (O_1897,N_14294,N_13308);
and UO_1898 (O_1898,N_14352,N_12884);
and UO_1899 (O_1899,N_13860,N_14962);
and UO_1900 (O_1900,N_13767,N_12402);
and UO_1901 (O_1901,N_12446,N_14505);
and UO_1902 (O_1902,N_12972,N_13188);
or UO_1903 (O_1903,N_13051,N_14770);
nand UO_1904 (O_1904,N_12750,N_14756);
or UO_1905 (O_1905,N_12410,N_13099);
nor UO_1906 (O_1906,N_14848,N_14590);
or UO_1907 (O_1907,N_14603,N_14899);
nand UO_1908 (O_1908,N_14341,N_12656);
and UO_1909 (O_1909,N_12311,N_13543);
nor UO_1910 (O_1910,N_13099,N_12859);
nand UO_1911 (O_1911,N_14583,N_13803);
and UO_1912 (O_1912,N_14807,N_13376);
or UO_1913 (O_1913,N_14947,N_13062);
or UO_1914 (O_1914,N_12462,N_12255);
or UO_1915 (O_1915,N_14086,N_13671);
xor UO_1916 (O_1916,N_14634,N_12259);
nand UO_1917 (O_1917,N_13852,N_13121);
nor UO_1918 (O_1918,N_13386,N_14830);
nor UO_1919 (O_1919,N_12314,N_12129);
and UO_1920 (O_1920,N_12049,N_12480);
nand UO_1921 (O_1921,N_12100,N_12687);
nor UO_1922 (O_1922,N_14578,N_12755);
nand UO_1923 (O_1923,N_12940,N_13340);
or UO_1924 (O_1924,N_13060,N_14876);
or UO_1925 (O_1925,N_12358,N_14844);
nand UO_1926 (O_1926,N_13604,N_14904);
or UO_1927 (O_1927,N_12913,N_14385);
and UO_1928 (O_1928,N_12310,N_13154);
and UO_1929 (O_1929,N_14019,N_14513);
or UO_1930 (O_1930,N_12436,N_12708);
and UO_1931 (O_1931,N_13572,N_13579);
nand UO_1932 (O_1932,N_13430,N_14185);
nor UO_1933 (O_1933,N_14827,N_14724);
or UO_1934 (O_1934,N_13648,N_14608);
nor UO_1935 (O_1935,N_13298,N_14088);
nor UO_1936 (O_1936,N_12078,N_13948);
nor UO_1937 (O_1937,N_12048,N_14050);
or UO_1938 (O_1938,N_12313,N_12525);
nor UO_1939 (O_1939,N_13143,N_12969);
or UO_1940 (O_1940,N_14089,N_14002);
and UO_1941 (O_1941,N_14394,N_14686);
nand UO_1942 (O_1942,N_14679,N_13556);
nor UO_1943 (O_1943,N_14161,N_13794);
or UO_1944 (O_1944,N_13821,N_12677);
nand UO_1945 (O_1945,N_13127,N_13340);
nand UO_1946 (O_1946,N_13127,N_14776);
nand UO_1947 (O_1947,N_13745,N_13857);
or UO_1948 (O_1948,N_12867,N_13417);
nand UO_1949 (O_1949,N_14348,N_14037);
or UO_1950 (O_1950,N_13128,N_14240);
nand UO_1951 (O_1951,N_14151,N_13465);
nand UO_1952 (O_1952,N_13445,N_12479);
nand UO_1953 (O_1953,N_14494,N_12800);
nor UO_1954 (O_1954,N_12103,N_14121);
nor UO_1955 (O_1955,N_14972,N_12758);
and UO_1956 (O_1956,N_14723,N_14830);
nor UO_1957 (O_1957,N_14926,N_12921);
and UO_1958 (O_1958,N_12633,N_12775);
nand UO_1959 (O_1959,N_13729,N_12702);
and UO_1960 (O_1960,N_14214,N_14789);
and UO_1961 (O_1961,N_12770,N_13440);
nand UO_1962 (O_1962,N_13853,N_13129);
and UO_1963 (O_1963,N_14343,N_12907);
nor UO_1964 (O_1964,N_13962,N_13935);
nand UO_1965 (O_1965,N_14449,N_12337);
or UO_1966 (O_1966,N_12363,N_14885);
or UO_1967 (O_1967,N_12688,N_12268);
nand UO_1968 (O_1968,N_14448,N_14169);
or UO_1969 (O_1969,N_12633,N_13968);
nand UO_1970 (O_1970,N_13342,N_13732);
nor UO_1971 (O_1971,N_13868,N_14708);
and UO_1972 (O_1972,N_13012,N_12055);
nor UO_1973 (O_1973,N_13888,N_14054);
or UO_1974 (O_1974,N_14018,N_12286);
or UO_1975 (O_1975,N_14570,N_14214);
nor UO_1976 (O_1976,N_14445,N_12848);
nor UO_1977 (O_1977,N_12727,N_12189);
xor UO_1978 (O_1978,N_14884,N_14784);
nand UO_1979 (O_1979,N_12106,N_14743);
and UO_1980 (O_1980,N_13596,N_12640);
or UO_1981 (O_1981,N_13294,N_12179);
nor UO_1982 (O_1982,N_12531,N_13945);
or UO_1983 (O_1983,N_12394,N_14467);
and UO_1984 (O_1984,N_12929,N_13093);
and UO_1985 (O_1985,N_12618,N_12686);
or UO_1986 (O_1986,N_14291,N_14861);
or UO_1987 (O_1987,N_12444,N_13671);
and UO_1988 (O_1988,N_12448,N_14390);
or UO_1989 (O_1989,N_14289,N_13534);
nand UO_1990 (O_1990,N_13625,N_12582);
nor UO_1991 (O_1991,N_12275,N_14996);
or UO_1992 (O_1992,N_13169,N_12778);
nor UO_1993 (O_1993,N_13661,N_13411);
and UO_1994 (O_1994,N_13729,N_12575);
and UO_1995 (O_1995,N_12012,N_12510);
or UO_1996 (O_1996,N_13399,N_14725);
and UO_1997 (O_1997,N_12760,N_14112);
nor UO_1998 (O_1998,N_13095,N_13392);
and UO_1999 (O_1999,N_14581,N_13542);
endmodule