module basic_3000_30000_3500_5_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_1812,In_525);
xnor U1 (N_1,In_2790,In_1822);
nand U2 (N_2,In_287,In_309);
or U3 (N_3,In_2962,In_1730);
nand U4 (N_4,In_268,In_2779);
xnor U5 (N_5,In_200,In_385);
and U6 (N_6,In_2320,In_214);
nand U7 (N_7,In_2625,In_2671);
xor U8 (N_8,In_247,In_1663);
and U9 (N_9,In_705,In_985);
nand U10 (N_10,In_1450,In_1736);
nand U11 (N_11,In_2987,In_2799);
nand U12 (N_12,In_1479,In_2984);
nor U13 (N_13,In_2111,In_1472);
xor U14 (N_14,In_2896,In_1901);
or U15 (N_15,In_1742,In_277);
nand U16 (N_16,In_645,In_205);
and U17 (N_17,In_414,In_2570);
nor U18 (N_18,In_1449,In_2433);
and U19 (N_19,In_2794,In_180);
xnor U20 (N_20,In_699,In_536);
or U21 (N_21,In_1635,In_1185);
and U22 (N_22,In_439,In_1747);
and U23 (N_23,In_1991,In_2481);
nor U24 (N_24,In_2319,In_692);
and U25 (N_25,In_2050,In_1188);
nor U26 (N_26,In_1287,In_1361);
or U27 (N_27,In_2894,In_556);
xor U28 (N_28,In_1580,In_2740);
xnor U29 (N_29,In_2933,In_2332);
and U30 (N_30,In_2659,In_1519);
nand U31 (N_31,In_339,In_592);
or U32 (N_32,In_388,In_738);
nor U33 (N_33,In_377,In_1197);
xnor U34 (N_34,In_1928,In_2759);
and U35 (N_35,In_955,In_1825);
xnor U36 (N_36,In_248,In_954);
nand U37 (N_37,In_1165,In_516);
or U38 (N_38,In_2104,In_917);
nor U39 (N_39,In_2158,In_1204);
xor U40 (N_40,In_1946,In_1958);
or U41 (N_41,In_1856,In_843);
nor U42 (N_42,In_882,In_1801);
nor U43 (N_43,In_453,In_1269);
and U44 (N_44,In_2792,In_2172);
nor U45 (N_45,In_1778,In_2170);
or U46 (N_46,In_1786,In_575);
or U47 (N_47,In_749,In_2943);
and U48 (N_48,In_623,In_1555);
or U49 (N_49,In_294,In_463);
nor U50 (N_50,In_282,In_179);
nand U51 (N_51,In_1485,In_2087);
xor U52 (N_52,In_2919,In_1978);
nand U53 (N_53,In_2995,In_1054);
xor U54 (N_54,In_259,In_291);
and U55 (N_55,In_2168,In_203);
nand U56 (N_56,In_2054,In_2819);
or U57 (N_57,In_2491,In_182);
nand U58 (N_58,In_1021,In_2692);
and U59 (N_59,In_1608,In_523);
xor U60 (N_60,In_2100,In_2365);
xor U61 (N_61,In_1163,In_2338);
and U62 (N_62,In_1029,In_142);
and U63 (N_63,In_506,In_1175);
nor U64 (N_64,In_1324,In_1317);
and U65 (N_65,In_1937,In_2525);
nand U66 (N_66,In_2895,In_1619);
nor U67 (N_67,In_1275,In_434);
nand U68 (N_68,In_1283,In_2150);
nor U69 (N_69,In_1629,In_119);
nor U70 (N_70,In_584,In_1233);
or U71 (N_71,In_56,In_588);
nand U72 (N_72,In_418,In_1504);
nor U73 (N_73,In_758,In_361);
or U74 (N_74,In_1068,In_2574);
nor U75 (N_75,In_2367,In_2245);
nand U76 (N_76,In_2994,In_780);
nor U77 (N_77,In_286,In_2745);
nor U78 (N_78,In_2078,In_2364);
xor U79 (N_79,In_109,In_2500);
nor U80 (N_80,In_1183,In_1086);
and U81 (N_81,In_1423,In_1848);
and U82 (N_82,In_2567,In_2556);
nand U83 (N_83,In_980,In_1025);
or U84 (N_84,In_338,In_1913);
xor U85 (N_85,In_17,In_986);
or U86 (N_86,In_1403,In_1173);
xor U87 (N_87,In_2515,In_940);
and U88 (N_88,In_1473,In_1988);
nor U89 (N_89,In_1834,In_2484);
xnor U90 (N_90,In_2932,In_684);
xor U91 (N_91,In_2923,In_2107);
nand U92 (N_92,In_2566,In_2086);
or U93 (N_93,In_124,In_2611);
nand U94 (N_94,In_832,In_387);
xor U95 (N_95,In_1126,In_1070);
xnor U96 (N_96,In_130,In_1613);
nor U97 (N_97,In_1690,In_1544);
and U98 (N_98,In_368,In_1105);
nand U99 (N_99,In_530,In_1350);
or U100 (N_100,In_406,In_881);
and U101 (N_101,In_932,In_1740);
or U102 (N_102,In_31,In_2108);
nand U103 (N_103,In_1203,In_381);
nor U104 (N_104,In_640,In_880);
nor U105 (N_105,In_1119,In_2471);
xnor U106 (N_106,In_643,In_2804);
and U107 (N_107,In_1929,In_84);
nand U108 (N_108,In_1157,In_718);
nor U109 (N_109,In_1898,In_1732);
xor U110 (N_110,In_1721,In_238);
nor U111 (N_111,In_1408,In_2483);
nor U112 (N_112,In_2475,In_9);
or U113 (N_113,In_145,In_2972);
nor U114 (N_114,In_234,In_1092);
or U115 (N_115,In_1514,In_2463);
or U116 (N_116,In_1083,In_469);
and U117 (N_117,In_1191,In_577);
nor U118 (N_118,In_2391,In_2957);
xor U119 (N_119,In_1813,In_2315);
nand U120 (N_120,In_1713,In_2612);
xnor U121 (N_121,In_266,In_1873);
xor U122 (N_122,In_2494,In_671);
and U123 (N_123,In_598,In_1093);
nor U124 (N_124,In_793,In_425);
or U125 (N_125,In_2029,In_1964);
nand U126 (N_126,In_1139,In_1493);
or U127 (N_127,In_2699,In_805);
and U128 (N_128,In_107,In_342);
nor U129 (N_129,In_468,In_1272);
nor U130 (N_130,In_1523,In_1917);
and U131 (N_131,In_2527,In_2660);
xnor U132 (N_132,In_208,In_801);
and U133 (N_133,In_112,In_1760);
nor U134 (N_134,In_628,In_1411);
or U135 (N_135,In_2241,In_1809);
or U136 (N_136,In_987,In_1155);
xor U137 (N_137,In_1775,In_1915);
nor U138 (N_138,In_1541,In_593);
xor U139 (N_139,In_736,In_2891);
nor U140 (N_140,In_1642,In_977);
nand U141 (N_141,In_672,In_1986);
nor U142 (N_142,In_918,In_2129);
or U143 (N_143,In_2493,In_2911);
xnor U144 (N_144,In_379,In_1246);
and U145 (N_145,In_1985,In_1285);
and U146 (N_146,In_2872,In_1885);
nor U147 (N_147,In_2650,In_1217);
and U148 (N_148,In_2325,In_1823);
and U149 (N_149,In_1075,In_622);
xor U150 (N_150,In_2024,In_1346);
or U151 (N_151,In_779,In_2835);
and U152 (N_152,In_1067,In_1062);
nand U153 (N_153,In_301,In_2003);
and U154 (N_154,In_26,In_1765);
xor U155 (N_155,In_1551,In_1871);
nor U156 (N_156,In_1118,In_2595);
nand U157 (N_157,In_2591,In_2064);
and U158 (N_158,In_1797,In_2198);
or U159 (N_159,In_1242,In_108);
nor U160 (N_160,In_73,In_2066);
nor U161 (N_161,In_2865,In_150);
nand U162 (N_162,In_2429,In_1431);
nand U163 (N_163,In_2431,In_243);
nand U164 (N_164,In_365,In_1647);
xnor U165 (N_165,In_1766,In_2856);
and U166 (N_166,In_2942,In_298);
nand U167 (N_167,In_289,In_1824);
xnor U168 (N_168,In_895,In_1558);
xor U169 (N_169,In_1798,In_1464);
and U170 (N_170,In_1112,In_2459);
nand U171 (N_171,In_2509,In_2452);
nand U172 (N_172,In_589,In_1664);
nor U173 (N_173,In_710,In_2934);
and U174 (N_174,In_2251,In_135);
and U175 (N_175,In_120,In_2353);
and U176 (N_176,In_1933,In_436);
nand U177 (N_177,In_1547,In_483);
xnor U178 (N_178,In_1889,In_2828);
nor U179 (N_179,In_2123,In_1792);
xnor U180 (N_180,In_2867,In_1421);
xor U181 (N_181,In_2091,In_1435);
nor U182 (N_182,In_2753,In_1733);
xnor U183 (N_183,In_1627,In_1677);
nand U184 (N_184,In_2148,In_1926);
or U185 (N_185,In_1772,In_902);
nor U186 (N_186,In_1193,In_2128);
nor U187 (N_187,In_373,In_224);
nor U188 (N_188,In_1425,In_1405);
nor U189 (N_189,In_2210,In_702);
or U190 (N_190,In_2990,In_1465);
nor U191 (N_191,In_2035,In_2358);
and U192 (N_192,In_2284,In_147);
xnor U193 (N_193,In_251,In_2613);
nor U194 (N_194,In_2547,In_2427);
or U195 (N_195,In_1113,In_423);
nor U196 (N_196,In_567,In_320);
nand U197 (N_197,In_747,In_1187);
xor U198 (N_198,In_315,In_2827);
or U199 (N_199,In_1320,In_1845);
nand U200 (N_200,In_1130,In_2512);
nor U201 (N_201,In_2157,In_2592);
nor U202 (N_202,In_155,In_1655);
xor U203 (N_203,In_2420,In_1327);
nor U204 (N_204,In_1018,In_1562);
nor U205 (N_205,In_92,In_229);
nand U206 (N_206,In_1074,In_1910);
nand U207 (N_207,In_118,In_494);
xnor U208 (N_208,In_2536,In_1417);
and U209 (N_209,In_1162,In_1347);
nand U210 (N_210,In_1050,In_2618);
xor U211 (N_211,In_2232,In_2034);
nor U212 (N_212,In_1553,In_544);
or U213 (N_213,In_1695,In_824);
nand U214 (N_214,In_2434,In_106);
xnor U215 (N_215,In_761,In_2290);
and U216 (N_216,In_1752,In_2057);
and U217 (N_217,In_834,In_1416);
or U218 (N_218,In_2614,In_1643);
xor U219 (N_219,In_1303,In_2996);
and U220 (N_220,In_897,In_2821);
and U221 (N_221,In_2372,In_2321);
or U222 (N_222,In_785,In_2263);
nand U223 (N_223,In_420,In_2246);
and U224 (N_224,In_2022,In_1728);
and U225 (N_225,In_856,In_2221);
or U226 (N_226,In_2514,In_1480);
or U227 (N_227,In_1355,In_2240);
and U228 (N_228,In_1774,In_460);
or U229 (N_229,In_808,In_249);
or U230 (N_230,In_85,In_1424);
or U231 (N_231,In_1266,In_825);
nor U232 (N_232,In_1329,In_926);
nand U233 (N_233,In_2698,In_1314);
and U234 (N_234,In_1058,In_1604);
nor U235 (N_235,In_1458,In_1996);
nor U236 (N_236,In_127,In_1605);
and U237 (N_237,In_1190,In_100);
and U238 (N_238,In_1141,In_609);
or U239 (N_239,In_1459,In_1279);
nor U240 (N_240,In_1152,In_1282);
or U241 (N_241,In_2324,In_2876);
nor U242 (N_242,In_1218,In_1236);
nor U243 (N_243,In_2897,In_2925);
nand U244 (N_244,In_111,In_1396);
nor U245 (N_245,In_1699,In_2092);
xnor U246 (N_246,In_1618,In_1082);
nor U247 (N_247,In_1484,In_1267);
xor U248 (N_248,In_1051,In_1154);
xnor U249 (N_249,In_2880,In_22);
and U250 (N_250,In_1364,In_1973);
nor U251 (N_251,In_966,In_1005);
or U252 (N_252,In_2354,In_891);
nor U253 (N_253,In_1345,In_1953);
nand U254 (N_254,In_2838,In_1631);
xnor U255 (N_255,In_1371,In_1791);
or U256 (N_256,In_809,In_2079);
xor U257 (N_257,In_2346,In_308);
and U258 (N_258,In_547,In_1637);
nand U259 (N_259,In_1867,In_393);
nor U260 (N_260,In_576,In_32);
nand U261 (N_261,In_1835,In_281);
and U262 (N_262,In_1507,In_680);
or U263 (N_263,In_2098,In_1697);
xnor U264 (N_264,In_51,In_161);
nor U265 (N_265,In_139,In_1881);
and U266 (N_266,In_2380,In_1446);
and U267 (N_267,In_1448,In_2147);
nor U268 (N_268,In_839,In_800);
and U269 (N_269,In_413,In_1516);
xor U270 (N_270,In_273,In_2033);
or U271 (N_271,In_629,In_1936);
and U272 (N_272,In_6,In_1970);
and U273 (N_273,In_2610,In_1753);
and U274 (N_274,In_1646,In_852);
and U275 (N_275,In_2732,In_1993);
nand U276 (N_276,In_305,In_213);
nor U277 (N_277,In_211,In_662);
nand U278 (N_278,In_2978,In_121);
and U279 (N_279,In_204,In_1998);
nor U280 (N_280,In_686,In_2317);
xnor U281 (N_281,In_1701,In_1461);
nor U282 (N_282,In_2710,In_2741);
or U283 (N_283,In_2018,In_919);
and U284 (N_284,In_2490,In_2080);
or U285 (N_285,In_2118,In_1100);
xor U286 (N_286,In_363,In_1120);
nor U287 (N_287,In_1633,In_86);
or U288 (N_288,In_1145,In_642);
xnor U289 (N_289,In_790,In_2960);
nand U290 (N_290,In_1056,In_1243);
nor U291 (N_291,In_2765,In_1496);
nor U292 (N_292,In_2849,In_716);
xor U293 (N_293,In_1960,In_1076);
xnor U294 (N_294,In_2814,In_1665);
nor U295 (N_295,In_2674,In_715);
nor U296 (N_296,In_1549,In_590);
and U297 (N_297,In_2629,In_2385);
or U298 (N_298,In_2016,In_2820);
or U299 (N_299,In_1526,In_1223);
nor U300 (N_300,In_845,In_2219);
xor U301 (N_301,In_1088,In_10);
nand U302 (N_302,In_242,In_2407);
nand U303 (N_303,In_2460,In_1574);
xnor U304 (N_304,In_730,In_1815);
nand U305 (N_305,In_49,In_535);
or U306 (N_306,In_2090,In_2025);
nor U307 (N_307,In_430,In_2900);
xor U308 (N_308,In_2936,In_113);
and U309 (N_309,In_930,In_956);
nor U310 (N_310,In_1925,In_689);
or U311 (N_311,In_1821,In_771);
xor U312 (N_312,In_2023,In_2907);
xor U313 (N_313,In_2575,In_98);
and U314 (N_314,In_2983,In_562);
nor U315 (N_315,In_2802,In_2883);
nor U316 (N_316,In_1622,In_2748);
or U317 (N_317,In_2853,In_781);
and U318 (N_318,In_2126,In_1156);
or U319 (N_319,In_646,In_2470);
or U320 (N_320,In_1768,In_2539);
or U321 (N_321,In_1950,In_2998);
nor U322 (N_322,In_1597,In_831);
xnor U323 (N_323,In_492,In_1048);
nand U324 (N_324,In_2510,In_2307);
nor U325 (N_325,In_725,In_74);
and U326 (N_326,In_39,In_2626);
xnor U327 (N_327,In_464,In_1342);
and U328 (N_328,In_1683,In_1718);
or U329 (N_329,In_274,In_1238);
xnor U330 (N_330,In_2289,In_1257);
and U331 (N_331,In_669,In_1447);
xnor U332 (N_332,In_2476,In_417);
nand U333 (N_333,In_201,In_1490);
nand U334 (N_334,In_1340,In_1300);
xnor U335 (N_335,In_743,In_768);
xor U336 (N_336,In_2194,In_165);
xor U337 (N_337,In_2106,In_531);
nor U338 (N_338,In_355,In_2019);
and U339 (N_339,In_431,In_1575);
and U340 (N_340,In_2884,In_157);
nor U341 (N_341,In_2337,In_404);
xor U342 (N_342,In_2077,In_2436);
xnor U343 (N_343,In_850,In_2946);
nand U344 (N_344,In_246,In_1146);
and U345 (N_345,In_1625,In_1767);
nand U346 (N_346,In_132,In_2330);
xor U347 (N_347,In_2679,In_602);
or U348 (N_348,In_2127,In_451);
nor U349 (N_349,In_647,In_2482);
nand U350 (N_350,In_2027,In_2557);
or U351 (N_351,In_1194,In_1626);
nor U352 (N_352,In_1965,In_1556);
or U353 (N_353,In_1291,In_1307);
or U354 (N_354,In_466,In_1440);
and U355 (N_355,In_1529,In_2860);
xnor U356 (N_356,In_1984,In_677);
or U357 (N_357,In_1044,In_1153);
and U358 (N_358,In_2384,In_685);
nand U359 (N_359,In_216,In_487);
or U360 (N_360,In_569,In_2653);
nor U361 (N_361,In_2938,In_2136);
or U362 (N_362,In_521,In_2747);
or U363 (N_363,In_664,In_1133);
xnor U364 (N_364,In_901,In_866);
nor U365 (N_365,In_2043,In_345);
xnor U366 (N_366,In_2248,In_2052);
nor U367 (N_367,In_864,In_482);
nand U368 (N_368,In_2915,In_1084);
nand U369 (N_369,In_1680,In_704);
nand U370 (N_370,In_411,In_2600);
or U371 (N_371,In_2405,In_2160);
and U372 (N_372,In_1542,In_1253);
xnor U373 (N_373,In_1035,In_44);
nand U374 (N_374,In_963,In_2146);
or U375 (N_375,In_2193,In_2787);
nand U376 (N_376,In_353,In_1482);
nor U377 (N_377,In_1564,In_2639);
nand U378 (N_378,In_81,In_1814);
nor U379 (N_379,In_2037,In_724);
or U380 (N_380,In_1395,In_457);
or U381 (N_381,In_1981,In_2334);
nand U382 (N_382,In_821,In_1462);
or U383 (N_383,In_2524,In_637);
nand U384 (N_384,In_389,In_1334);
xor U385 (N_385,In_2760,In_1802);
and U386 (N_386,In_2065,In_285);
nor U387 (N_387,In_606,In_2914);
and U388 (N_388,In_978,In_1393);
nand U389 (N_389,In_2901,In_1181);
xnor U390 (N_390,In_2737,In_2072);
or U391 (N_391,In_278,In_2700);
or U392 (N_392,In_1623,In_2563);
or U393 (N_393,In_220,In_2440);
xnor U394 (N_394,In_250,In_2784);
nor U395 (N_395,In_2212,In_1366);
nor U396 (N_396,In_1632,In_2530);
or U397 (N_397,In_2597,In_2229);
nor U398 (N_398,In_2882,In_1932);
or U399 (N_399,In_2793,In_811);
and U400 (N_400,In_925,In_1271);
xor U401 (N_401,In_674,In_803);
nor U402 (N_402,In_1080,In_504);
nor U403 (N_403,In_1148,In_2795);
nand U404 (N_404,In_495,In_2950);
and U405 (N_405,In_2579,In_1169);
nand U406 (N_406,In_2685,In_1795);
nand U407 (N_407,In_424,In_2339);
xor U408 (N_408,In_1045,In_916);
and U409 (N_409,In_2561,In_2889);
xor U410 (N_410,In_2124,In_546);
nor U411 (N_411,In_1091,In_83);
and U412 (N_412,In_2392,In_708);
nor U413 (N_413,In_2125,In_1963);
xor U414 (N_414,In_879,In_2988);
or U415 (N_415,In_1333,In_2654);
nor U416 (N_416,In_2084,In_2190);
and U417 (N_417,In_2417,In_968);
nor U418 (N_418,In_2013,In_538);
xor U419 (N_419,In_1134,In_1476);
nor U420 (N_420,In_2428,In_756);
and U421 (N_421,In_2885,In_1968);
nor U422 (N_422,In_2492,In_2267);
and U423 (N_423,In_826,In_2408);
or U424 (N_424,In_2062,In_1323);
or U425 (N_425,In_711,In_2116);
nand U426 (N_426,In_1586,In_2719);
and U427 (N_427,In_2414,In_126);
nand U428 (N_428,In_378,In_1225);
and U429 (N_429,In_1702,In_1397);
or U430 (N_430,In_920,In_2068);
or U431 (N_431,In_841,In_2442);
or U432 (N_432,In_415,In_2419);
nor U433 (N_433,In_860,In_1443);
xor U434 (N_434,In_144,In_855);
xor U435 (N_435,In_618,In_2448);
nand U436 (N_436,In_2155,In_1277);
or U437 (N_437,In_1337,In_799);
nand U438 (N_438,In_75,In_2931);
or U439 (N_439,In_358,In_2991);
xnor U440 (N_440,In_750,In_1755);
or U441 (N_441,In_2707,In_1987);
nand U442 (N_442,In_868,In_2049);
xnor U443 (N_443,In_1128,In_1612);
or U444 (N_444,In_2056,In_2426);
nor U445 (N_445,In_1794,In_2581);
nand U446 (N_446,In_1077,In_2299);
xor U447 (N_447,In_2902,In_35);
nor U448 (N_448,In_64,In_1908);
nand U449 (N_449,In_312,In_1666);
xnor U450 (N_450,In_231,In_1170);
and U451 (N_451,In_971,In_1262);
and U452 (N_452,In_1260,In_905);
xnor U453 (N_453,In_1897,In_196);
nor U454 (N_454,In_2242,In_2989);
nand U455 (N_455,In_734,In_2133);
nor U456 (N_456,In_2560,In_2866);
or U457 (N_457,In_773,In_2350);
and U458 (N_458,In_2006,In_1956);
nor U459 (N_459,In_2306,In_1621);
nor U460 (N_460,In_1330,In_1382);
nand U461 (N_461,In_1178,In_2585);
nand U462 (N_462,In_2153,In_763);
nand U463 (N_463,In_2046,In_691);
or U464 (N_464,In_513,In_138);
and U465 (N_465,In_193,In_2316);
or U466 (N_466,In_2209,In_2389);
or U467 (N_467,In_2472,In_311);
nand U468 (N_468,In_2498,In_459);
and U469 (N_469,In_2236,In_2410);
nor U470 (N_470,In_2163,In_333);
nand U471 (N_471,In_921,In_2397);
and U472 (N_472,In_2196,In_1228);
and U473 (N_473,In_1326,In_1995);
or U474 (N_474,In_1543,In_2047);
and U475 (N_475,In_1979,In_1247);
and U476 (N_476,In_1388,In_1365);
nand U477 (N_477,In_2668,In_346);
nor U478 (N_478,In_2576,In_1512);
nor U479 (N_479,In_2189,In_1356);
or U480 (N_480,In_853,In_957);
xor U481 (N_481,In_1634,In_2113);
and U482 (N_482,In_2461,In_380);
xnor U483 (N_483,In_1101,In_1833);
xor U484 (N_484,In_280,In_731);
nor U485 (N_485,In_1692,In_1418);
nor U486 (N_486,In_448,In_2038);
nor U487 (N_487,In_2051,In_1488);
xor U488 (N_488,In_1237,In_507);
or U489 (N_489,In_1433,In_1511);
and U490 (N_490,In_2873,In_2278);
nor U491 (N_491,In_260,In_2616);
and U492 (N_492,In_2675,In_1895);
nor U493 (N_493,In_1308,In_549);
or U494 (N_494,In_1325,In_398);
nor U495 (N_495,In_2094,In_360);
nor U496 (N_496,In_2763,In_953);
xnor U497 (N_497,In_2542,In_1135);
nand U498 (N_498,In_2298,In_115);
and U499 (N_499,In_2800,In_70);
xor U500 (N_500,In_480,In_458);
nand U501 (N_501,In_1955,In_117);
xnor U502 (N_502,In_2252,In_2844);
nor U503 (N_503,In_2980,In_712);
xor U504 (N_504,In_631,In_1280);
nand U505 (N_505,In_1869,In_2269);
and U506 (N_506,In_2261,In_136);
or U507 (N_507,In_875,In_561);
nand U508 (N_508,In_522,In_2836);
xor U509 (N_509,In_2726,In_2850);
or U510 (N_510,In_2222,In_2352);
nand U511 (N_511,In_488,In_192);
and U512 (N_512,In_2396,In_2965);
and U513 (N_513,In_2818,In_306);
nand U514 (N_514,In_2467,In_23);
or U515 (N_515,In_2048,In_181);
nand U516 (N_516,In_2905,In_141);
xnor U517 (N_517,In_348,In_2383);
and U518 (N_518,In_2709,In_1301);
or U519 (N_519,In_1617,In_1527);
nand U520 (N_520,In_176,In_240);
nand U521 (N_521,In_1457,In_543);
nor U522 (N_522,In_2855,In_898);
nand U523 (N_523,In_2226,In_2845);
and U524 (N_524,In_2015,In_326);
and U525 (N_525,In_2690,In_2439);
xnor U526 (N_526,In_962,In_1295);
nand U527 (N_527,In_1147,In_1799);
or U528 (N_528,In_2258,In_1299);
or U529 (N_529,In_1536,In_1358);
nand U530 (N_530,In_746,In_2893);
or U531 (N_531,In_2070,In_2357);
xnor U532 (N_532,In_597,In_2739);
nand U533 (N_533,In_1391,In_1131);
and U534 (N_534,In_976,In_2132);
and U535 (N_535,In_444,In_1585);
xor U536 (N_536,In_2227,In_2620);
nor U537 (N_537,In_2403,In_1827);
and U538 (N_538,In_2206,In_1592);
or U539 (N_539,In_765,In_1037);
or U540 (N_540,In_1079,In_1264);
or U541 (N_541,In_2135,In_965);
xor U542 (N_542,In_1894,In_2971);
xnor U543 (N_543,In_1107,In_2039);
nor U544 (N_544,In_1316,In_739);
or U545 (N_545,In_2295,In_2430);
xnor U546 (N_546,In_2120,In_1769);
nor U547 (N_547,In_71,In_1843);
nand U548 (N_548,In_1255,In_996);
nand U549 (N_549,In_1180,In_2117);
and U550 (N_550,In_1353,In_792);
nand U551 (N_551,In_1557,In_1031);
xnor U552 (N_552,In_471,In_131);
nor U553 (N_553,In_599,In_1649);
or U554 (N_554,In_2255,In_226);
and U555 (N_555,In_518,In_2568);
nor U556 (N_556,In_2412,In_1495);
and U557 (N_557,In_427,In_390);
or U558 (N_558,In_343,In_665);
nor U559 (N_559,In_2159,In_2647);
nand U560 (N_560,In_770,In_2947);
nand U561 (N_561,In_636,In_798);
and U562 (N_562,In_1302,In_2340);
or U563 (N_563,In_551,In_183);
xnor U564 (N_564,In_1352,In_2553);
or U565 (N_565,In_1422,In_1278);
or U566 (N_566,In_1103,In_1057);
nand U567 (N_567,In_2264,In_892);
xnor U568 (N_568,In_1601,In_2406);
nand U569 (N_569,In_1854,In_2924);
nand U570 (N_570,In_814,In_604);
xnor U571 (N_571,In_1254,In_2165);
and U572 (N_572,In_842,In_329);
nor U573 (N_573,In_2959,In_2555);
xnor U574 (N_574,In_1890,In_776);
and U575 (N_575,In_20,In_1492);
nand U576 (N_576,In_2823,In_137);
and U577 (N_577,In_1059,In_456);
xor U578 (N_578,In_1687,In_2270);
or U579 (N_579,In_1875,In_1452);
nand U580 (N_580,In_2462,In_1997);
and U581 (N_581,In_2223,In_103);
or U582 (N_582,In_215,In_2564);
and U583 (N_583,In_1453,In_1566);
and U584 (N_584,In_1383,In_648);
xor U585 (N_585,In_2704,In_2341);
nand U586 (N_586,In_2489,In_2722);
xnor U587 (N_587,In_133,In_2776);
xor U588 (N_588,In_876,In_651);
nor U589 (N_589,In_336,In_1989);
nand U590 (N_590,In_2580,In_2749);
xnor U591 (N_591,In_797,In_514);
nor U592 (N_592,In_2259,In_582);
nor U593 (N_593,In_2031,In_2502);
nor U594 (N_594,In_936,In_681);
nand U595 (N_595,In_581,In_89);
and U596 (N_596,In_299,In_1012);
xor U597 (N_597,In_1099,In_1974);
xnor U598 (N_598,In_397,In_1842);
and U599 (N_599,In_914,In_969);
nor U600 (N_600,In_344,In_2458);
and U601 (N_601,In_1888,In_2218);
xnor U602 (N_602,In_2968,In_318);
or U603 (N_603,In_2953,In_2394);
nor U604 (N_604,In_2249,In_666);
and U605 (N_605,In_327,In_719);
xor U606 (N_606,In_1349,In_2966);
nor U607 (N_607,In_1381,In_2067);
nand U608 (N_608,In_2211,In_1132);
or U609 (N_609,In_1708,In_2785);
or U610 (N_610,In_300,In_1176);
nand U611 (N_611,In_595,In_2605);
xnor U612 (N_612,In_2393,In_910);
or U613 (N_613,In_1415,In_1803);
or U614 (N_614,In_2273,In_579);
xnor U615 (N_615,In_586,In_1678);
nor U616 (N_616,In_893,In_1682);
and U617 (N_617,In_591,In_1335);
nand U618 (N_618,In_668,In_696);
nor U619 (N_619,In_2930,In_2326);
and U620 (N_620,In_2643,In_1943);
nand U621 (N_621,In_2724,In_2617);
xor U622 (N_622,In_1859,In_129);
nor U623 (N_623,In_2712,In_2161);
nor U624 (N_624,In_869,In_1876);
xor U625 (N_625,In_1106,In_1610);
and U626 (N_626,In_255,In_2488);
nor U627 (N_627,In_1905,In_1377);
nand U628 (N_628,In_1069,In_1214);
and U629 (N_629,In_911,In_236);
nand U630 (N_630,In_1456,In_1331);
nand U631 (N_631,In_1883,In_2738);
nand U632 (N_632,In_973,In_2345);
nand U633 (N_633,In_1033,In_2008);
and U634 (N_634,In_2552,In_2277);
and U635 (N_635,In_2411,In_2045);
or U636 (N_636,In_1782,In_499);
xor U637 (N_637,In_2310,In_102);
nor U638 (N_638,In_1,In_2742);
nand U639 (N_639,In_2234,In_1581);
or U640 (N_640,In_2485,In_1952);
and U641 (N_641,In_959,In_2641);
nand U642 (N_642,In_2314,In_1081);
nor U643 (N_643,In_2680,In_1042);
xnor U644 (N_644,In_2926,In_2002);
xnor U645 (N_645,In_922,In_2026);
and U646 (N_646,In_2829,In_1866);
xor U647 (N_647,In_2669,In_1222);
or U648 (N_648,In_1837,In_2982);
or U649 (N_649,In_2810,In_1734);
nor U650 (N_650,In_1055,In_465);
and U651 (N_651,In_1852,In_1359);
nor U652 (N_652,In_1990,In_1136);
and U653 (N_653,In_2171,In_836);
nand U654 (N_654,In_1019,In_2812);
and U655 (N_655,In_2961,In_2767);
and U656 (N_656,In_2997,In_1104);
or U657 (N_657,In_1249,In_2074);
nand U658 (N_658,In_830,In_2766);
xor U659 (N_659,In_1182,In_1641);
xnor U660 (N_660,In_1310,In_1942);
xor U661 (N_661,In_2422,In_225);
xnor U662 (N_662,In_1537,In_1780);
and U663 (N_663,In_654,In_449);
nor U664 (N_664,In_1640,In_2651);
or U665 (N_665,In_2627,In_1644);
nand U666 (N_666,In_2571,In_509);
xor U667 (N_667,In_25,In_1007);
nand U668 (N_668,In_635,In_1705);
xor U669 (N_669,In_2468,In_616);
nand U670 (N_670,In_1491,In_2009);
nor U671 (N_671,In_1589,In_396);
xnor U672 (N_672,In_638,In_657);
xor U673 (N_673,In_1502,In_1087);
or U674 (N_674,In_497,In_1673);
nor U675 (N_675,In_1380,In_822);
and U676 (N_676,In_2725,In_1032);
nor U677 (N_677,In_1669,In_2729);
and U678 (N_678,In_854,In_1052);
nor U679 (N_679,In_1561,In_1851);
and U680 (N_680,In_899,In_1967);
or U681 (N_681,In_2085,In_1606);
or U682 (N_682,In_2890,In_2409);
nor U683 (N_683,In_2318,In_158);
or U684 (N_684,In_2142,In_772);
nor U685 (N_685,In_580,In_149);
nor U686 (N_686,In_1659,In_620);
nor U687 (N_687,In_2005,In_619);
and U688 (N_688,In_1312,In_1209);
and U689 (N_689,In_1602,In_2138);
nand U690 (N_690,In_906,In_1745);
or U691 (N_691,In_2940,In_2305);
xnor U692 (N_692,In_2435,In_1144);
nand U693 (N_693,In_2139,In_1836);
or U694 (N_694,In_319,In_783);
nand U695 (N_695,In_438,In_2847);
nand U696 (N_696,In_2182,In_356);
or U697 (N_697,In_261,In_2333);
and U698 (N_698,In_2801,In_695);
xor U699 (N_699,In_2344,In_362);
or U700 (N_700,In_510,In_1703);
nand U701 (N_701,In_1013,In_2474);
and U702 (N_702,In_1857,In_258);
or U703 (N_703,In_2811,In_2271);
nor U704 (N_704,In_697,In_894);
nor U705 (N_705,In_2286,In_2505);
nand U706 (N_706,In_2681,In_1645);
nor U707 (N_707,In_1611,In_2775);
or U708 (N_708,In_804,In_2606);
xor U709 (N_709,In_1129,In_1252);
or U710 (N_710,In_807,In_55);
and U711 (N_711,In_2642,In_1234);
and U712 (N_712,In_740,In_627);
nor U713 (N_713,In_313,In_195);
xor U714 (N_714,In_663,In_1438);
nand U715 (N_715,In_1861,In_2447);
xor U716 (N_716,In_239,In_477);
or U717 (N_717,In_1097,In_2816);
nor U718 (N_718,In_1700,In_1918);
nand U719 (N_719,In_2870,In_2879);
xnor U720 (N_720,In_767,In_367);
xnor U721 (N_721,In_566,In_1008);
nor U722 (N_722,In_2727,In_1027);
or U723 (N_723,In_1717,In_1737);
nand U724 (N_724,In_1348,In_884);
and U725 (N_725,In_1000,In_2373);
or U726 (N_726,In_981,In_1878);
xnor U727 (N_727,In_1198,In_944);
xor U728 (N_728,In_1662,In_2293);
nand U729 (N_729,In_1977,In_2673);
xnor U730 (N_730,In_419,In_1220);
xor U731 (N_731,In_303,In_775);
nor U732 (N_732,In_670,In_2554);
and U733 (N_733,In_2368,In_1039);
and U734 (N_734,In_1800,In_2705);
or U735 (N_735,In_2773,In_1923);
xor U736 (N_736,In_194,In_1781);
or U737 (N_737,In_874,In_958);
and U738 (N_738,In_2162,In_2511);
and U739 (N_739,In_256,In_1587);
nor U740 (N_740,In_2369,In_1921);
nand U741 (N_741,In_173,In_1951);
nand U742 (N_742,In_1143,In_601);
and U743 (N_743,In_479,In_96);
nand U744 (N_744,In_1213,In_578);
and U745 (N_745,In_2308,In_2688);
xor U746 (N_746,In_1290,In_2010);
and U747 (N_747,In_2970,In_2881);
nor U748 (N_748,In_573,In_952);
xnor U749 (N_749,In_1534,In_1743);
xor U750 (N_750,In_1614,In_1167);
and U751 (N_751,In_2858,In_2756);
xnor U752 (N_752,In_2347,In_766);
nor U753 (N_753,In_79,In_2846);
nor U754 (N_754,In_1922,In_1847);
xnor U755 (N_755,In_1763,In_199);
nand U756 (N_756,In_1525,In_1115);
nand U757 (N_757,In_2551,In_1508);
xor U758 (N_758,In_1796,In_1714);
and U759 (N_759,In_481,In_2287);
or U760 (N_760,In_1521,In_2154);
xnor U761 (N_761,In_502,In_2275);
xor U762 (N_762,In_762,In_2663);
xor U763 (N_763,In_270,In_2283);
nor U764 (N_764,In_244,In_653);
or U765 (N_765,In_617,In_1817);
nor U766 (N_766,In_82,In_16);
or U767 (N_767,In_2473,In_304);
and U768 (N_768,In_198,In_587);
nand U769 (N_769,In_1095,In_2529);
nand U770 (N_770,In_2207,In_1014);
or U771 (N_771,In_1432,In_1785);
and U772 (N_772,In_401,In_2466);
nand U773 (N_773,In_729,In_1201);
nand U774 (N_774,In_57,In_1899);
xor U775 (N_775,In_27,In_778);
nor U776 (N_776,In_887,In_2061);
and U777 (N_777,In_1487,In_2956);
or U778 (N_778,In_995,In_227);
or U779 (N_779,In_1064,In_532);
nor U780 (N_780,In_2543,In_1838);
xnor U781 (N_781,In_230,In_2399);
nor U782 (N_782,In_1594,In_1387);
nor U783 (N_783,In_2706,In_5);
nand U784 (N_784,In_827,In_2497);
nand U785 (N_785,In_632,In_1931);
and U786 (N_786,In_386,In_2593);
or U787 (N_787,In_2963,In_1463);
and U788 (N_788,In_1919,In_2053);
and U789 (N_789,In_2913,In_1616);
nor U790 (N_790,In_2220,In_2291);
nor U791 (N_791,In_1400,In_872);
or U792 (N_792,In_2910,In_2666);
nor U793 (N_793,In_2017,In_384);
or U794 (N_794,In_269,In_175);
nor U795 (N_795,In_1517,In_42);
nor U796 (N_796,In_2922,In_1124);
xnor U797 (N_797,In_63,In_2202);
nand U798 (N_798,In_253,In_994);
or U799 (N_799,In_1927,In_1628);
xor U800 (N_800,In_66,In_1009);
nand U801 (N_801,In_2081,In_2586);
or U802 (N_802,In_1509,In_693);
nand U803 (N_803,In_2423,In_2780);
and U804 (N_804,In_2021,In_1938);
and U805 (N_805,In_416,In_2114);
xor U806 (N_806,In_1043,In_596);
or U807 (N_807,In_493,In_2619);
and U808 (N_808,In_1651,In_806);
nand U809 (N_809,In_1961,In_1127);
or U810 (N_810,In_2723,In_1379);
xor U811 (N_811,In_2020,In_2175);
xor U812 (N_812,In_1428,In_2030);
and U813 (N_813,In_999,In_1288);
or U814 (N_814,In_2603,In_1351);
nand U815 (N_815,In_683,In_717);
nand U816 (N_816,In_1189,In_1406);
xor U817 (N_817,In_2296,In_1399);
and U818 (N_818,In_2204,In_2059);
or U819 (N_819,In_2174,In_2912);
or U820 (N_820,In_1579,In_2327);
nor U821 (N_821,In_38,In_2119);
and U822 (N_822,In_1657,In_2103);
and U823 (N_823,In_741,In_2588);
or U824 (N_824,In_2041,In_1293);
and U825 (N_825,In_1980,In_541);
or U826 (N_826,In_931,In_782);
and U827 (N_827,In_2381,In_2469);
nor U828 (N_828,In_2355,In_908);
xnor U829 (N_829,In_732,In_54);
and U830 (N_830,In_2646,In_1211);
xor U831 (N_831,In_537,In_505);
nor U832 (N_832,In_435,In_322);
nand U833 (N_833,In_1945,In_688);
and U834 (N_834,In_2569,In_2063);
nor U835 (N_835,In_1595,In_1966);
and U836 (N_836,In_2717,In_2262);
xor U837 (N_837,In_1286,In_1466);
nand U838 (N_838,In_186,In_2239);
and U839 (N_839,In_2878,In_53);
xnor U840 (N_840,In_1546,In_151);
or U841 (N_841,In_934,In_2796);
nor U842 (N_842,In_2060,In_2071);
nor U843 (N_843,In_1200,In_633);
nand U844 (N_844,In_209,In_302);
and U845 (N_845,In_764,In_2243);
or U846 (N_846,In_1149,In_1481);
xnor U847 (N_847,In_2214,In_1685);
or U848 (N_848,In_330,In_2589);
and U849 (N_849,In_432,In_655);
xor U850 (N_850,In_2149,In_2892);
and U851 (N_851,In_1609,In_706);
xnor U852 (N_852,In_1389,In_2655);
or U853 (N_853,In_1992,In_340);
nand U854 (N_854,In_2540,In_1554);
nor U855 (N_855,In_788,In_1550);
nand U856 (N_856,In_1034,In_2645);
nor U857 (N_857,In_1741,In_1367);
nor U858 (N_858,In_1221,In_1924);
xnor U859 (N_859,In_909,In_1868);
or U860 (N_860,In_1321,In_99);
or U861 (N_861,In_2007,In_2215);
and U862 (N_862,In_612,In_2122);
nand U863 (N_863,In_2519,In_2716);
nand U864 (N_864,In_292,In_796);
nor U865 (N_865,In_116,In_152);
xor U866 (N_866,In_169,In_759);
or U867 (N_867,In_1771,In_2387);
and U868 (N_868,In_2178,In_737);
nor U869 (N_869,In_1896,In_1846);
or U870 (N_870,In_1232,In_2105);
or U871 (N_871,In_2920,In_2208);
nand U872 (N_872,In_844,In_1123);
or U873 (N_873,In_948,In_2714);
nand U874 (N_874,In_1172,In_1761);
and U875 (N_875,In_913,In_1322);
nor U876 (N_876,In_1339,In_838);
or U877 (N_877,In_1831,In_2253);
and U878 (N_878,In_787,In_405);
and U879 (N_879,In_585,In_422);
nand U880 (N_880,In_374,In_2501);
and U881 (N_881,In_550,In_87);
nand U882 (N_882,In_1137,In_166);
nand U883 (N_883,In_553,In_613);
xnor U884 (N_884,In_1715,In_950);
nor U885 (N_885,In_36,In_2359);
xor U886 (N_886,In_2783,In_837);
or U887 (N_887,In_2032,In_988);
xor U888 (N_888,In_937,In_1343);
nand U889 (N_889,In_170,In_2001);
xnor U890 (N_890,In_2791,In_1368);
or U891 (N_891,In_2521,In_1332);
nand U892 (N_892,In_1679,In_1684);
or U893 (N_893,In_2213,In_2887);
nor U894 (N_894,In_658,In_1948);
nand U895 (N_895,In_219,In_337);
or U896 (N_896,In_2701,In_2302);
and U897 (N_897,In_1419,In_990);
xnor U898 (N_898,In_2328,In_2096);
nor U899 (N_899,In_2083,In_1522);
or U900 (N_900,In_904,In_395);
nor U901 (N_901,In_1313,In_1259);
nor U902 (N_902,In_1208,In_974);
or U903 (N_903,In_2728,In_2322);
xnor U904 (N_904,In_2888,In_2102);
nor U905 (N_905,In_1670,In_1731);
or U906 (N_906,In_212,In_2134);
nor U907 (N_907,In_2825,In_1195);
nor U908 (N_908,In_794,In_870);
or U909 (N_909,In_1455,In_2832);
and U910 (N_910,In_1940,In_189);
nor U911 (N_911,In_1319,In_2266);
nand U912 (N_912,In_1196,In_2624);
or U913 (N_913,In_1693,In_1475);
nand U914 (N_914,In_1026,In_2181);
nand U915 (N_915,In_383,In_2842);
and U916 (N_916,In_1578,In_2145);
xnor U917 (N_917,In_271,In_392);
nand U918 (N_918,In_2301,In_2762);
and U919 (N_919,In_1844,In_1567);
or U920 (N_920,In_2798,In_1036);
nor U921 (N_921,In_237,In_134);
nor U922 (N_922,In_2904,In_610);
or U923 (N_923,In_153,In_2441);
and U924 (N_924,In_2203,In_1344);
xor U925 (N_925,In_1230,In_1434);
xnor U926 (N_926,In_2948,In_2830);
nand U927 (N_927,In_2418,In_2375);
and U928 (N_928,In_1826,In_2069);
or U929 (N_929,In_2750,In_2192);
and U930 (N_930,In_2455,In_933);
nor U931 (N_931,In_1274,In_1954);
nor U932 (N_932,In_467,In_1298);
and U933 (N_933,In_2371,In_1654);
nor U934 (N_934,In_997,In_1660);
nor U935 (N_935,In_1624,In_533);
or U936 (N_936,In_450,In_2374);
and U937 (N_937,In_222,In_19);
or U938 (N_938,In_473,In_1756);
nor U939 (N_939,In_2831,In_2803);
or U940 (N_940,In_2854,In_223);
or U941 (N_941,In_2323,In_2686);
xnor U942 (N_942,In_375,In_2443);
or U943 (N_943,In_753,In_218);
nor U944 (N_944,In_701,In_1179);
and U945 (N_945,In_2993,In_1240);
or U946 (N_946,In_961,In_1607);
xnor U947 (N_947,In_2628,In_1583);
or U948 (N_948,In_2630,In_2981);
nor U949 (N_949,In_350,In_2577);
xnor U950 (N_950,In_1863,In_818);
nand U951 (N_951,In_447,In_2735);
nand U952 (N_952,In_1751,In_2044);
nand U953 (N_953,In_123,In_2752);
nand U954 (N_954,In_335,In_927);
xor U955 (N_955,In_433,In_2986);
xnor U956 (N_956,In_1268,In_903);
nand U957 (N_957,In_1392,In_1117);
or U958 (N_958,In_1674,In_2974);
or U959 (N_959,In_1891,In_1572);
nor U960 (N_960,In_2187,In_1591);
nor U961 (N_961,In_1486,In_2583);
nor U962 (N_962,In_1906,In_1328);
xnor U963 (N_963,In_1650,In_2444);
xor U964 (N_964,In_1378,In_1227);
nand U965 (N_965,In_426,In_1442);
and U966 (N_966,In_2388,In_50);
nor U967 (N_967,In_1858,In_1046);
xnor U968 (N_968,In_733,In_1808);
or U969 (N_969,In_2903,In_88);
xor U970 (N_970,In_2309,In_1882);
and U971 (N_971,In_288,In_1532);
nand U972 (N_972,In_1372,In_428);
and U973 (N_973,In_548,In_69);
xnor U974 (N_974,In_1724,In_1711);
or U975 (N_975,In_429,In_1251);
xnor U976 (N_976,In_1828,In_1427);
nor U977 (N_977,In_2144,In_979);
and U978 (N_978,In_2538,In_2076);
xnor U979 (N_979,In_2404,In_1704);
and U980 (N_980,In_2596,In_1520);
xnor U981 (N_981,In_496,In_529);
and U982 (N_982,In_500,In_2928);
nand U983 (N_983,In_162,In_1880);
nand U984 (N_984,In_290,In_2097);
xor U985 (N_985,In_2004,In_2667);
nand U986 (N_986,In_829,In_2416);
and U987 (N_987,In_534,In_245);
or U988 (N_988,In_1892,In_2058);
and U989 (N_989,In_2734,In_886);
nor U990 (N_990,In_2755,In_1011);
nor U991 (N_991,In_2141,In_2143);
xnor U992 (N_992,In_262,In_2110);
xnor U993 (N_993,In_1498,In_2693);
nand U994 (N_994,In_594,In_1874);
or U995 (N_995,In_721,In_1318);
nor U996 (N_996,In_1494,In_1451);
xnor U997 (N_997,In_1436,In_858);
nand U998 (N_998,In_1681,In_1513);
nor U999 (N_999,In_900,In_700);
nand U1000 (N_1000,In_2425,In_1870);
nand U1001 (N_1001,In_2546,In_2185);
nor U1002 (N_1002,In_2992,In_284);
xnor U1003 (N_1003,In_1315,In_1903);
and U1004 (N_1004,In_2806,In_1265);
nand U1005 (N_1005,In_2312,In_2661);
and U1006 (N_1006,In_2486,In_2609);
xor U1007 (N_1007,In_1754,In_1584);
or U1008 (N_1008,In_2808,In_1573);
nand U1009 (N_1009,In_1256,In_1620);
nand U1010 (N_1010,In_2532,In_442);
or U1011 (N_1011,In_812,In_2311);
xnor U1012 (N_1012,In_2637,In_352);
nor U1013 (N_1013,In_2508,In_2935);
or U1014 (N_1014,In_45,In_2520);
nor U1015 (N_1015,In_557,In_1108);
xor U1016 (N_1016,In_817,In_90);
and U1017 (N_1017,In_1390,In_2402);
and U1018 (N_1018,In_1577,In_726);
xnor U1019 (N_1019,In_2073,In_2973);
and U1020 (N_1020,In_2826,In_2012);
xor U1021 (N_1021,In_2014,In_989);
xnor U1022 (N_1022,In_992,In_774);
xor U1023 (N_1023,In_2817,In_2840);
and U1024 (N_1024,In_58,In_2861);
xor U1025 (N_1025,In_2622,In_2349);
nor U1026 (N_1026,In_1096,In_97);
nand U1027 (N_1027,In_2684,In_1709);
and U1028 (N_1028,In_2356,In_2256);
or U1029 (N_1029,In_399,In_1720);
nor U1030 (N_1030,In_634,In_652);
nor U1031 (N_1031,In_1528,In_849);
or U1032 (N_1032,In_2112,In_2770);
and U1033 (N_1033,In_1855,In_324);
or U1034 (N_1034,In_2774,In_1174);
or U1035 (N_1035,In_2777,In_929);
and U1036 (N_1036,In_2632,In_354);
nand U1037 (N_1037,In_1750,In_470);
nand U1038 (N_1038,In_486,In_1832);
nor U1039 (N_1039,In_15,In_848);
nor U1040 (N_1040,In_1078,In_2869);
xor U1041 (N_1041,In_1540,In_2451);
nand U1042 (N_1042,In_283,In_2781);
and U1043 (N_1043,In_65,In_1689);
xnor U1044 (N_1044,In_2534,In_2558);
xor U1045 (N_1045,In_2082,In_1239);
or U1046 (N_1046,In_1281,In_1710);
nor U1047 (N_1047,In_2758,In_2805);
xnor U1048 (N_1048,In_2746,In_177);
nand U1049 (N_1049,In_1944,In_2664);
or U1050 (N_1050,In_2424,In_95);
nor U1051 (N_1051,In_2954,In_2225);
or U1052 (N_1052,In_1603,In_520);
nor U1053 (N_1053,In_1811,In_2678);
nor U1054 (N_1054,In_2565,In_174);
and U1055 (N_1055,In_552,In_1864);
xor U1056 (N_1056,In_641,In_1538);
nor U1057 (N_1057,In_2395,In_2782);
nor U1058 (N_1058,In_37,In_515);
and U1059 (N_1059,In_1477,In_924);
xnor U1060 (N_1060,In_2851,In_752);
nor U1061 (N_1061,In_265,In_1072);
nand U1062 (N_1062,In_511,In_2545);
xnor U1063 (N_1063,In_29,In_607);
xor U1064 (N_1064,In_1818,In_11);
or U1065 (N_1065,In_890,In_1049);
xnor U1066 (N_1066,In_2363,In_1370);
and U1067 (N_1067,In_810,In_1675);
and U1068 (N_1068,In_187,In_2254);
xor U1069 (N_1069,In_676,In_2398);
nor U1070 (N_1070,In_2244,In_2797);
or U1071 (N_1071,In_2453,In_1949);
nand U1072 (N_1072,In_1779,In_476);
or U1073 (N_1073,In_745,In_2351);
nand U1074 (N_1074,In_659,In_760);
nor U1075 (N_1075,In_2868,In_1235);
nor U1076 (N_1076,In_1653,In_2691);
xnor U1077 (N_1077,In_2281,In_371);
nand U1078 (N_1078,In_2496,In_366);
xor U1079 (N_1079,In_2944,In_349);
nor U1080 (N_1080,In_939,In_264);
nor U1081 (N_1081,In_2413,In_941);
or U1082 (N_1082,In_1028,In_2839);
nor U1083 (N_1083,In_1615,In_2949);
and U1084 (N_1084,In_2623,In_2179);
and U1085 (N_1085,In_1468,In_156);
nand U1086 (N_1086,In_1971,In_815);
nor U1087 (N_1087,In_735,In_2342);
xor U1088 (N_1088,In_154,In_2415);
and U1089 (N_1089,In_2513,In_1111);
or U1090 (N_1090,In_60,In_2528);
or U1091 (N_1091,In_1524,In_2672);
and U1092 (N_1092,In_519,In_382);
or U1093 (N_1093,In_1306,In_408);
nor U1094 (N_1094,In_1444,In_2109);
xor U1095 (N_1095,In_2292,In_1671);
nand U1096 (N_1096,In_871,In_2535);
nand U1097 (N_1097,In_172,In_2272);
or U1098 (N_1098,In_1999,In_1276);
nand U1099 (N_1099,In_2772,In_2297);
xnor U1100 (N_1100,In_2644,In_571);
xor U1101 (N_1101,In_114,In_370);
or U1102 (N_1102,In_885,In_2506);
and U1103 (N_1103,In_2279,In_2590);
or U1104 (N_1104,In_1229,In_754);
nor U1105 (N_1105,In_1789,In_1959);
xnor U1106 (N_1106,In_656,In_110);
xor U1107 (N_1107,In_2195,In_347);
nor U1108 (N_1108,In_539,In_1916);
xor U1109 (N_1109,In_2843,In_190);
xor U1110 (N_1110,In_649,In_851);
and U1111 (N_1111,In_1939,In_440);
or U1112 (N_1112,In_1219,In_351);
and U1113 (N_1113,In_1727,In_1764);
nor U1114 (N_1114,In_861,In_923);
and U1115 (N_1115,In_2744,In_2480);
xnor U1116 (N_1116,In_445,In_1930);
nand U1117 (N_1117,In_2205,In_21);
nand U1118 (N_1118,In_2769,In_1506);
and U1119 (N_1119,In_1725,In_407);
nor U1120 (N_1120,In_1820,In_263);
xor U1121 (N_1121,In_2656,In_2584);
and U1122 (N_1122,In_455,In_210);
nand U1123 (N_1123,In_1688,In_1094);
nand U1124 (N_1124,In_1402,In_568);
xnor U1125 (N_1125,In_960,In_1887);
xor U1126 (N_1126,In_30,In_2633);
and U1127 (N_1127,In_1909,In_667);
or U1128 (N_1128,In_1893,In_2200);
nor U1129 (N_1129,In_2898,In_1160);
nor U1130 (N_1130,In_2761,In_1505);
and U1131 (N_1131,In_517,In_1159);
nor U1132 (N_1132,In_2101,In_2857);
nand U1133 (N_1133,In_2694,In_605);
and U1134 (N_1134,In_563,In_2465);
or U1135 (N_1135,In_296,In_2683);
nand U1136 (N_1136,In_2733,In_2999);
nand U1137 (N_1137,In_835,In_94);
nor U1138 (N_1138,In_2631,In_1304);
nor U1139 (N_1139,In_2449,In_1499);
nor U1140 (N_1140,In_1016,In_2604);
or U1141 (N_1141,In_1309,In_1003);
or U1142 (N_1142,In_1510,In_935);
nand U1143 (N_1143,In_1503,In_624);
nand U1144 (N_1144,In_2516,In_2864);
nand U1145 (N_1145,In_1972,In_1063);
nand U1146 (N_1146,In_2335,In_1166);
xor U1147 (N_1147,In_1454,In_2863);
nand U1148 (N_1148,In_2437,In_1570);
or U1149 (N_1149,In_2598,In_503);
xor U1150 (N_1150,In_1362,In_2587);
and U1151 (N_1151,In_1245,In_2541);
xnor U1152 (N_1152,In_1250,In_2788);
or U1153 (N_1153,In_1205,In_2233);
nand U1154 (N_1154,In_2975,In_1593);
nor U1155 (N_1155,In_528,In_639);
nand U1156 (N_1156,In_2602,In_2937);
or U1157 (N_1157,In_40,In_217);
or U1158 (N_1158,In_947,In_1138);
or U1159 (N_1159,In_1518,In_2361);
nor U1160 (N_1160,In_865,In_2390);
nor U1161 (N_1161,In_1047,In_1489);
xor U1162 (N_1162,In_1412,In_2638);
nand U1163 (N_1163,In_2055,In_2478);
or U1164 (N_1164,In_1338,In_2379);
nand U1165 (N_1165,In_912,In_77);
and U1166 (N_1166,In_2230,In_1150);
nor U1167 (N_1167,In_2697,In_877);
nand U1168 (N_1168,In_1114,In_1017);
nor U1169 (N_1169,In_2495,In_421);
and U1170 (N_1170,In_714,In_1004);
and U1171 (N_1171,In_2824,In_1053);
xor U1172 (N_1172,In_328,In_2730);
nand U1173 (N_1173,In_751,In_2176);
nor U1174 (N_1174,In_889,In_2615);
xnor U1175 (N_1175,In_679,In_185);
xor U1176 (N_1176,In_2703,In_2115);
and U1177 (N_1177,In_1474,In_2751);
nand U1178 (N_1178,In_1914,In_122);
and U1179 (N_1179,In_982,In_2036);
and U1180 (N_1180,In_2702,In_626);
nor U1181 (N_1181,In_1386,In_252);
and U1182 (N_1182,In_1002,In_2531);
nor U1183 (N_1183,In_1426,In_2432);
nand U1184 (N_1184,In_475,In_777);
and U1185 (N_1185,In_678,In_1941);
nand U1186 (N_1186,In_2874,In_1841);
xnor U1187 (N_1187,In_501,In_1122);
nor U1188 (N_1188,In_1186,In_608);
or U1189 (N_1189,In_1161,In_2979);
nor U1190 (N_1190,In_819,In_1793);
xnor U1191 (N_1191,In_2964,In_276);
xnor U1192 (N_1192,In_2445,In_235);
xnor U1193 (N_1193,In_1957,In_2268);
or U1194 (N_1194,In_441,In_221);
nor U1195 (N_1195,In_2303,In_437);
xor U1196 (N_1196,In_1559,In_603);
nand U1197 (N_1197,In_359,In_873);
nor U1198 (N_1198,In_484,In_630);
and U1199 (N_1199,In_2833,In_1533);
nand U1200 (N_1200,In_2562,In_2362);
and U1201 (N_1201,In_2164,In_2677);
xor U1202 (N_1202,In_742,In_1401);
nand U1203 (N_1203,In_2421,In_325);
and U1204 (N_1204,In_2657,In_478);
nand U1205 (N_1205,In_93,In_2370);
and U1206 (N_1206,In_412,In_1719);
nor U1207 (N_1207,In_946,In_24);
or U1208 (N_1208,In_1142,In_33);
nand U1209 (N_1209,In_1648,In_2093);
nor U1210 (N_1210,In_41,In_2533);
nand U1211 (N_1211,In_1015,In_279);
xnor U1212 (N_1212,In_1471,In_1212);
or U1213 (N_1213,In_1409,In_72);
and U1214 (N_1214,In_2875,In_188);
and U1215 (N_1215,In_1171,In_143);
nand U1216 (N_1216,In_275,In_2294);
nand U1217 (N_1217,In_896,In_784);
nand U1218 (N_1218,In_1210,In_295);
nand U1219 (N_1219,In_1588,In_661);
nand U1220 (N_1220,In_1912,In_1776);
and U1221 (N_1221,In_687,In_2809);
nand U1222 (N_1222,In_802,In_2523);
nand U1223 (N_1223,In_1787,In_1065);
and U1224 (N_1224,In_1911,In_2768);
xnor U1225 (N_1225,In_1483,In_1788);
nand U1226 (N_1226,In_1385,In_2649);
and U1227 (N_1227,In_2599,In_364);
or U1228 (N_1228,In_2754,In_512);
xor U1229 (N_1229,In_1816,In_1289);
or U1230 (N_1230,In_68,In_2877);
or U1231 (N_1231,In_2377,In_314);
or U1232 (N_1232,In_1073,In_1773);
nand U1233 (N_1233,In_1038,In_682);
nor U1234 (N_1234,In_1040,In_795);
or U1235 (N_1235,In_28,In_2621);
or U1236 (N_1236,In_1982,In_709);
nor U1237 (N_1237,In_1983,In_823);
or U1238 (N_1238,In_2862,In_228);
and U1239 (N_1239,In_332,In_555);
and U1240 (N_1240,In_2789,In_2695);
nand U1241 (N_1241,In_698,In_14);
xor U1242 (N_1242,In_1840,In_2304);
or U1243 (N_1243,In_1006,In_2969);
and U1244 (N_1244,In_394,In_524);
nor U1245 (N_1245,In_2662,In_2985);
nor U1246 (N_1246,In_2257,In_1041);
nand U1247 (N_1247,In_1758,In_2689);
nand U1248 (N_1248,In_2152,In_820);
nor U1249 (N_1249,In_2088,In_2658);
and U1250 (N_1250,In_1630,In_621);
nor U1251 (N_1251,In_970,In_1430);
and U1252 (N_1252,In_310,In_1829);
or U1253 (N_1253,In_2952,In_297);
xor U1254 (N_1254,In_2186,In_232);
and U1255 (N_1255,In_1294,In_1865);
xnor U1256 (N_1256,In_2871,In_1394);
or U1257 (N_1257,In_2859,In_1739);
xnor U1258 (N_1258,In_2916,In_1749);
nor U1259 (N_1259,In_1636,In_2336);
nor U1260 (N_1260,In_472,In_2238);
nand U1261 (N_1261,In_2582,In_1723);
nor U1262 (N_1262,In_2977,In_1548);
or U1263 (N_1263,In_1224,In_1902);
and U1264 (N_1264,In_625,In_0);
nor U1265 (N_1265,In_2228,In_1886);
and U1266 (N_1266,In_59,In_307);
and U1267 (N_1267,In_1360,In_600);
xnor U1268 (N_1268,In_558,In_1226);
or U1269 (N_1269,In_2216,In_1691);
xor U1270 (N_1270,In_1296,In_1907);
xor U1271 (N_1271,In_2000,In_148);
xnor U1272 (N_1272,In_1429,In_1746);
nor U1273 (N_1273,In_813,In_1877);
nor U1274 (N_1274,In_1469,In_984);
nor U1275 (N_1275,In_140,In_341);
and U1276 (N_1276,In_2939,In_1969);
and U1277 (N_1277,In_2499,In_2918);
nand U1278 (N_1278,In_2217,In_2197);
nand U1279 (N_1279,In_2121,In_1261);
nand U1280 (N_1280,In_722,In_2288);
nand U1281 (N_1281,In_2955,In_1672);
nand U1282 (N_1282,In_2075,In_1121);
nor U1283 (N_1283,In_1373,In_2366);
nor U1284 (N_1284,In_2343,In_1661);
xor U1285 (N_1285,In_1676,In_2265);
xnor U1286 (N_1286,In_1470,In_727);
nor U1287 (N_1287,In_1374,In_391);
nand U1288 (N_1288,In_2507,In_1668);
nand U1289 (N_1289,In_1839,In_572);
or U1290 (N_1290,In_1460,In_1023);
and U1291 (N_1291,In_907,In_1060);
nand U1292 (N_1292,In_67,In_1140);
xnor U1293 (N_1293,In_2300,In_403);
or U1294 (N_1294,In_452,In_1500);
xor U1295 (N_1295,In_2457,In_1576);
and U1296 (N_1296,In_2450,In_48);
nand U1297 (N_1297,In_2648,In_2464);
and U1298 (N_1298,In_1098,In_1777);
or U1299 (N_1299,In_1860,In_206);
nand U1300 (N_1300,In_660,In_184);
xor U1301 (N_1301,In_241,In_833);
nor U1302 (N_1302,In_1357,In_1192);
xnor U1303 (N_1303,In_2607,In_410);
or U1304 (N_1304,In_2518,In_527);
nor U1305 (N_1305,In_4,In_1010);
nor U1306 (N_1306,In_1810,In_443);
xor U1307 (N_1307,In_1202,In_554);
or U1308 (N_1308,In_560,In_2608);
nor U1309 (N_1309,In_2169,In_164);
and U1310 (N_1310,In_1270,In_1638);
nor U1311 (N_1311,In_1770,In_1501);
nand U1312 (N_1312,In_125,In_2095);
and U1313 (N_1313,In_2191,In_2477);
or U1314 (N_1314,In_964,In_545);
and U1315 (N_1315,In_402,In_76);
xor U1316 (N_1316,In_2522,In_2682);
or U1317 (N_1317,In_1441,In_207);
xnor U1318 (N_1318,In_748,In_2771);
or U1319 (N_1319,In_2479,In_1407);
nor U1320 (N_1320,In_2360,In_357);
or U1321 (N_1321,In_2601,In_46);
nor U1322 (N_1322,In_915,In_2274);
or U1323 (N_1323,In_1102,In_2670);
and U1324 (N_1324,In_2718,In_1071);
or U1325 (N_1325,In_720,In_728);
and U1326 (N_1326,In_1884,In_2526);
and U1327 (N_1327,In_723,In_1904);
xnor U1328 (N_1328,In_975,In_1748);
xnor U1329 (N_1329,In_1652,In_1375);
nor U1330 (N_1330,In_1738,In_2348);
xor U1331 (N_1331,In_2183,In_564);
nor U1332 (N_1332,In_1248,In_943);
nor U1333 (N_1333,In_2696,In_1024);
nand U1334 (N_1334,In_707,In_828);
and U1335 (N_1335,In_1116,In_1759);
or U1336 (N_1336,In_1437,In_1872);
and U1337 (N_1337,In_454,In_2537);
or U1338 (N_1338,In_1439,In_317);
and U1339 (N_1339,In_2958,In_2927);
nor U1340 (N_1340,In_1284,In_1258);
nand U1341 (N_1341,In_2578,In_293);
or U1342 (N_1342,In_2040,In_1694);
xor U1343 (N_1343,In_485,In_1698);
nand U1344 (N_1344,In_1109,In_1849);
and U1345 (N_1345,In_34,In_769);
nand U1346 (N_1346,In_1151,In_1735);
and U1347 (N_1347,In_1231,In_1110);
and U1348 (N_1348,In_1976,In_2635);
and U1349 (N_1349,In_2929,In_3);
nor U1350 (N_1350,In_1061,In_2559);
nand U1351 (N_1351,In_1292,In_1596);
nor U1352 (N_1352,In_526,In_2676);
or U1353 (N_1353,In_1020,In_400);
xor U1354 (N_1354,In_2549,In_1263);
nand U1355 (N_1355,In_1363,In_12);
or U1356 (N_1356,In_2042,In_1125);
and U1357 (N_1357,In_786,In_2708);
nor U1358 (N_1358,In_816,In_2834);
nand U1359 (N_1359,In_2813,In_1729);
and U1360 (N_1360,In_2634,In_1420);
xnor U1361 (N_1361,In_2166,In_878);
or U1362 (N_1362,In_2837,In_2378);
or U1363 (N_1363,In_1369,In_565);
nand U1364 (N_1364,In_2247,In_1706);
or U1365 (N_1365,In_972,In_867);
or U1366 (N_1366,In_1582,In_2573);
xor U1367 (N_1367,In_1515,In_1560);
nand U1368 (N_1368,In_2548,In_2487);
nand U1369 (N_1369,In_2456,In_2313);
xor U1370 (N_1370,In_372,In_2899);
nor U1371 (N_1371,In_1639,In_1085);
nand U1372 (N_1372,In_650,In_2177);
or U1373 (N_1373,In_755,In_857);
or U1374 (N_1374,In_1656,In_2276);
and U1375 (N_1375,In_2594,In_1445);
or U1376 (N_1376,In_570,In_508);
xor U1377 (N_1377,In_1497,In_1467);
xnor U1378 (N_1378,In_840,In_2967);
or U1379 (N_1379,In_1590,In_1001);
xor U1380 (N_1380,In_2151,In_1598);
and U1381 (N_1381,In_52,In_1686);
or U1382 (N_1382,In_2285,In_938);
xnor U1383 (N_1383,In_2917,In_1478);
nor U1384 (N_1384,In_2282,In_2386);
and U1385 (N_1385,In_789,In_171);
and U1386 (N_1386,In_1531,In_2237);
and U1387 (N_1387,In_1862,In_2550);
and U1388 (N_1388,In_2945,In_945);
xor U1389 (N_1389,In_160,In_167);
and U1390 (N_1390,In_1819,In_43);
nand U1391 (N_1391,In_1600,In_80);
nor U1392 (N_1392,In_574,In_2572);
xor U1393 (N_1393,In_1806,In_1030);
nor U1394 (N_1394,In_1879,In_316);
or U1395 (N_1395,In_1757,In_446);
xor U1396 (N_1396,In_1535,In_2184);
nor U1397 (N_1397,In_1667,In_2224);
nor U1398 (N_1398,In_2713,In_1563);
and U1399 (N_1399,In_2454,In_191);
or U1400 (N_1400,In_1696,In_2400);
nand U1401 (N_1401,In_2822,In_104);
xor U1402 (N_1402,In_644,In_1712);
nand U1403 (N_1403,In_7,In_1305);
nand U1404 (N_1404,In_847,In_159);
or U1405 (N_1405,In_254,In_2807);
nand U1406 (N_1406,In_1241,In_2180);
and U1407 (N_1407,In_1273,In_257);
nor U1408 (N_1408,In_1022,In_1565);
xor U1409 (N_1409,In_1297,In_2721);
xor U1410 (N_1410,In_998,In_2201);
or U1411 (N_1411,In_2640,In_1900);
or U1412 (N_1412,In_2446,In_791);
and U1413 (N_1413,In_1920,In_2235);
nand U1414 (N_1414,In_1658,In_690);
xnor U1415 (N_1415,In_1090,In_267);
nor U1416 (N_1416,In_1726,In_321);
nand U1417 (N_1417,In_1850,In_983);
or U1418 (N_1418,In_331,In_18);
nand U1419 (N_1419,In_1790,In_1716);
xnor U1420 (N_1420,In_1089,In_2260);
nand U1421 (N_1421,In_2099,In_163);
xor U1422 (N_1422,In_489,In_1962);
and U1423 (N_1423,In_2652,In_2401);
xor U1424 (N_1424,In_1184,In_1158);
xnor U1425 (N_1425,In_1216,In_1398);
nand U1426 (N_1426,In_2848,In_1215);
or U1427 (N_1427,In_1066,In_462);
nor U1428 (N_1428,In_2786,In_2976);
nor U1429 (N_1429,In_498,In_1376);
and U1430 (N_1430,In_2909,In_1404);
nand U1431 (N_1431,In_233,In_491);
or U1432 (N_1432,In_2331,In_1807);
and U1433 (N_1433,In_146,In_2736);
or U1434 (N_1434,In_2250,In_2438);
xor U1435 (N_1435,In_1530,In_703);
nand U1436 (N_1436,In_2011,In_2711);
nor U1437 (N_1437,In_1569,In_928);
nand U1438 (N_1438,In_673,In_2906);
nor U1439 (N_1439,In_1762,In_967);
nor U1440 (N_1440,In_2687,In_675);
or U1441 (N_1441,In_1571,In_2376);
and U1442 (N_1442,In_542,In_376);
nor U1443 (N_1443,In_2280,In_1744);
xor U1444 (N_1444,In_1783,In_2715);
or U1445 (N_1445,In_951,In_2731);
or U1446 (N_1446,In_2028,In_1384);
nor U1447 (N_1447,In_1539,In_2140);
nand U1448 (N_1448,In_91,In_13);
nand U1449 (N_1449,In_1994,In_178);
and U1450 (N_1450,In_2329,In_2173);
nor U1451 (N_1451,In_846,In_2089);
xor U1452 (N_1452,In_1545,In_409);
or U1453 (N_1453,In_1207,In_101);
nand U1454 (N_1454,In_1830,In_559);
nor U1455 (N_1455,In_2886,In_859);
and U1456 (N_1456,In_1804,In_1552);
or U1457 (N_1457,In_1805,In_2167);
xor U1458 (N_1458,In_949,In_1414);
nor U1459 (N_1459,In_2764,In_2130);
nor U1460 (N_1460,In_1853,In_105);
nor U1461 (N_1461,In_694,In_2231);
xnor U1462 (N_1462,In_1168,In_1975);
nor U1463 (N_1463,In_757,In_2815);
nor U1464 (N_1464,In_1341,In_713);
nor U1465 (N_1465,In_2504,In_888);
and U1466 (N_1466,In_540,In_1935);
or U1467 (N_1467,In_1599,In_1311);
and U1468 (N_1468,In_991,In_2720);
nor U1469 (N_1469,In_2665,In_1410);
and U1470 (N_1470,In_883,In_197);
xnor U1471 (N_1471,In_2636,In_369);
and U1472 (N_1472,In_2131,In_461);
nand U1473 (N_1473,In_1244,In_615);
xor U1474 (N_1474,In_1707,In_8);
or U1475 (N_1475,In_862,In_2);
nand U1476 (N_1476,In_62,In_168);
and U1477 (N_1477,In_2852,In_2544);
or U1478 (N_1478,In_323,In_1934);
and U1479 (N_1479,In_611,In_2757);
xor U1480 (N_1480,In_1199,In_863);
and U1481 (N_1481,In_2156,In_1164);
or U1482 (N_1482,In_2199,In_2743);
nand U1483 (N_1483,In_1336,In_993);
and U1484 (N_1484,In_1784,In_2503);
nor U1485 (N_1485,In_2137,In_2382);
nor U1486 (N_1486,In_1177,In_2941);
or U1487 (N_1487,In_61,In_128);
nor U1488 (N_1488,In_1568,In_47);
or U1489 (N_1489,In_744,In_2517);
xnor U1490 (N_1490,In_490,In_2908);
and U1491 (N_1491,In_1722,In_1354);
and U1492 (N_1492,In_2841,In_942);
or U1493 (N_1493,In_2921,In_2951);
nand U1494 (N_1494,In_2778,In_614);
nand U1495 (N_1495,In_474,In_334);
and U1496 (N_1496,In_1206,In_272);
nor U1497 (N_1497,In_2188,In_78);
and U1498 (N_1498,In_583,In_202);
or U1499 (N_1499,In_1413,In_1947);
or U1500 (N_1500,In_1734,In_2563);
or U1501 (N_1501,In_1547,In_1535);
nor U1502 (N_1502,In_2536,In_2587);
or U1503 (N_1503,In_2415,In_2066);
nor U1504 (N_1504,In_1951,In_1330);
nor U1505 (N_1505,In_2668,In_498);
nand U1506 (N_1506,In_2643,In_2201);
xnor U1507 (N_1507,In_1975,In_2698);
or U1508 (N_1508,In_423,In_2160);
or U1509 (N_1509,In_1140,In_1258);
or U1510 (N_1510,In_2576,In_2855);
nor U1511 (N_1511,In_1961,In_2220);
nand U1512 (N_1512,In_2545,In_1559);
xnor U1513 (N_1513,In_1653,In_2943);
nor U1514 (N_1514,In_64,In_629);
or U1515 (N_1515,In_2154,In_1309);
xnor U1516 (N_1516,In_2494,In_1454);
and U1517 (N_1517,In_958,In_1037);
xnor U1518 (N_1518,In_1125,In_2129);
nor U1519 (N_1519,In_743,In_2781);
nor U1520 (N_1520,In_2060,In_2914);
xnor U1521 (N_1521,In_2591,In_1903);
or U1522 (N_1522,In_1519,In_2460);
nor U1523 (N_1523,In_1418,In_2822);
xor U1524 (N_1524,In_2787,In_2047);
xor U1525 (N_1525,In_2552,In_1762);
and U1526 (N_1526,In_1992,In_389);
nand U1527 (N_1527,In_829,In_429);
and U1528 (N_1528,In_2171,In_2215);
xor U1529 (N_1529,In_674,In_1056);
and U1530 (N_1530,In_1999,In_2975);
xor U1531 (N_1531,In_703,In_2948);
nand U1532 (N_1532,In_1519,In_1195);
and U1533 (N_1533,In_2880,In_61);
and U1534 (N_1534,In_2014,In_1299);
or U1535 (N_1535,In_1563,In_1800);
and U1536 (N_1536,In_1516,In_2035);
nand U1537 (N_1537,In_364,In_2330);
or U1538 (N_1538,In_1360,In_58);
nor U1539 (N_1539,In_1124,In_348);
xor U1540 (N_1540,In_1147,In_2328);
and U1541 (N_1541,In_1047,In_2853);
or U1542 (N_1542,In_472,In_2353);
nor U1543 (N_1543,In_1062,In_918);
xnor U1544 (N_1544,In_2185,In_1384);
and U1545 (N_1545,In_897,In_2941);
nor U1546 (N_1546,In_2652,In_1473);
nand U1547 (N_1547,In_2908,In_87);
nand U1548 (N_1548,In_2418,In_2995);
nand U1549 (N_1549,In_1741,In_117);
or U1550 (N_1550,In_339,In_2267);
or U1551 (N_1551,In_1990,In_1631);
nand U1552 (N_1552,In_2326,In_1307);
nand U1553 (N_1553,In_1644,In_736);
and U1554 (N_1554,In_2099,In_2254);
and U1555 (N_1555,In_493,In_2879);
nand U1556 (N_1556,In_442,In_1278);
or U1557 (N_1557,In_1532,In_2346);
nand U1558 (N_1558,In_1594,In_1343);
xnor U1559 (N_1559,In_1870,In_2249);
nor U1560 (N_1560,In_2693,In_876);
nor U1561 (N_1561,In_2909,In_1705);
nor U1562 (N_1562,In_1924,In_1663);
or U1563 (N_1563,In_369,In_1644);
nor U1564 (N_1564,In_1545,In_2644);
and U1565 (N_1565,In_86,In_1536);
and U1566 (N_1566,In_2838,In_1981);
and U1567 (N_1567,In_2152,In_306);
xnor U1568 (N_1568,In_1648,In_2633);
and U1569 (N_1569,In_374,In_417);
or U1570 (N_1570,In_2951,In_1820);
and U1571 (N_1571,In_2619,In_1334);
nor U1572 (N_1572,In_1508,In_2025);
or U1573 (N_1573,In_2346,In_1677);
nand U1574 (N_1574,In_1839,In_401);
and U1575 (N_1575,In_1304,In_2180);
xor U1576 (N_1576,In_315,In_2758);
and U1577 (N_1577,In_2470,In_1319);
nor U1578 (N_1578,In_1298,In_1552);
or U1579 (N_1579,In_2120,In_1834);
nor U1580 (N_1580,In_2120,In_1539);
nor U1581 (N_1581,In_745,In_797);
or U1582 (N_1582,In_1456,In_2739);
nand U1583 (N_1583,In_470,In_1189);
or U1584 (N_1584,In_391,In_1405);
nand U1585 (N_1585,In_0,In_109);
or U1586 (N_1586,In_2217,In_894);
or U1587 (N_1587,In_1365,In_722);
or U1588 (N_1588,In_2146,In_1860);
xor U1589 (N_1589,In_1389,In_216);
and U1590 (N_1590,In_454,In_2438);
xnor U1591 (N_1591,In_2419,In_743);
nand U1592 (N_1592,In_2301,In_2971);
or U1593 (N_1593,In_441,In_2029);
and U1594 (N_1594,In_1445,In_1759);
xnor U1595 (N_1595,In_2938,In_2007);
nand U1596 (N_1596,In_436,In_720);
or U1597 (N_1597,In_2724,In_80);
xor U1598 (N_1598,In_476,In_114);
and U1599 (N_1599,In_2589,In_2696);
and U1600 (N_1600,In_2158,In_242);
and U1601 (N_1601,In_1068,In_1481);
and U1602 (N_1602,In_980,In_2637);
or U1603 (N_1603,In_2173,In_634);
nand U1604 (N_1604,In_48,In_600);
or U1605 (N_1605,In_2339,In_660);
or U1606 (N_1606,In_2024,In_736);
nand U1607 (N_1607,In_410,In_870);
nor U1608 (N_1608,In_784,In_398);
xnor U1609 (N_1609,In_2730,In_2587);
or U1610 (N_1610,In_379,In_2032);
nand U1611 (N_1611,In_855,In_664);
nand U1612 (N_1612,In_2474,In_1696);
or U1613 (N_1613,In_2560,In_2786);
nand U1614 (N_1614,In_1421,In_2255);
nand U1615 (N_1615,In_2874,In_446);
nor U1616 (N_1616,In_1394,In_547);
xor U1617 (N_1617,In_240,In_698);
nor U1618 (N_1618,In_488,In_1878);
xor U1619 (N_1619,In_2094,In_1135);
xnor U1620 (N_1620,In_2321,In_2346);
or U1621 (N_1621,In_665,In_2025);
and U1622 (N_1622,In_282,In_607);
and U1623 (N_1623,In_1733,In_2809);
nand U1624 (N_1624,In_1855,In_2294);
nor U1625 (N_1625,In_2172,In_1457);
and U1626 (N_1626,In_2461,In_2596);
nor U1627 (N_1627,In_1244,In_1615);
nor U1628 (N_1628,In_2167,In_1683);
xor U1629 (N_1629,In_744,In_2824);
and U1630 (N_1630,In_2728,In_2855);
nand U1631 (N_1631,In_2848,In_1374);
xnor U1632 (N_1632,In_1258,In_1868);
and U1633 (N_1633,In_2722,In_2348);
nand U1634 (N_1634,In_2413,In_2868);
xnor U1635 (N_1635,In_2846,In_1476);
nor U1636 (N_1636,In_2458,In_1616);
nor U1637 (N_1637,In_2821,In_647);
xnor U1638 (N_1638,In_1736,In_2917);
or U1639 (N_1639,In_2437,In_1214);
and U1640 (N_1640,In_424,In_2073);
xnor U1641 (N_1641,In_325,In_1389);
xnor U1642 (N_1642,In_1454,In_1784);
and U1643 (N_1643,In_38,In_2536);
or U1644 (N_1644,In_2241,In_489);
and U1645 (N_1645,In_2841,In_351);
nor U1646 (N_1646,In_1020,In_246);
nor U1647 (N_1647,In_1433,In_1895);
or U1648 (N_1648,In_2884,In_1285);
nor U1649 (N_1649,In_1299,In_1317);
or U1650 (N_1650,In_2285,In_2056);
xnor U1651 (N_1651,In_448,In_1236);
and U1652 (N_1652,In_2304,In_2795);
nand U1653 (N_1653,In_2995,In_2662);
xor U1654 (N_1654,In_2803,In_1569);
nand U1655 (N_1655,In_2971,In_34);
or U1656 (N_1656,In_2891,In_889);
or U1657 (N_1657,In_383,In_2710);
nand U1658 (N_1658,In_1429,In_498);
nor U1659 (N_1659,In_1055,In_583);
and U1660 (N_1660,In_285,In_2448);
xnor U1661 (N_1661,In_1446,In_121);
and U1662 (N_1662,In_1381,In_2894);
or U1663 (N_1663,In_2081,In_870);
nor U1664 (N_1664,In_402,In_1743);
nand U1665 (N_1665,In_66,In_231);
and U1666 (N_1666,In_561,In_862);
and U1667 (N_1667,In_266,In_796);
nor U1668 (N_1668,In_2211,In_821);
or U1669 (N_1669,In_1728,In_1881);
nor U1670 (N_1670,In_771,In_2354);
nor U1671 (N_1671,In_95,In_1277);
and U1672 (N_1672,In_970,In_445);
nand U1673 (N_1673,In_7,In_2832);
xor U1674 (N_1674,In_1277,In_919);
xor U1675 (N_1675,In_181,In_2900);
or U1676 (N_1676,In_1287,In_1717);
nor U1677 (N_1677,In_396,In_1810);
nor U1678 (N_1678,In_1294,In_2867);
xor U1679 (N_1679,In_0,In_1334);
xor U1680 (N_1680,In_2914,In_2242);
nor U1681 (N_1681,In_1191,In_1308);
xor U1682 (N_1682,In_2200,In_2495);
or U1683 (N_1683,In_2247,In_1462);
xor U1684 (N_1684,In_1811,In_1038);
nor U1685 (N_1685,In_1401,In_1391);
and U1686 (N_1686,In_149,In_1778);
and U1687 (N_1687,In_2520,In_723);
xor U1688 (N_1688,In_1226,In_2299);
nand U1689 (N_1689,In_2891,In_722);
nand U1690 (N_1690,In_234,In_2250);
or U1691 (N_1691,In_1443,In_2002);
nand U1692 (N_1692,In_27,In_2391);
nor U1693 (N_1693,In_1526,In_1098);
or U1694 (N_1694,In_859,In_607);
and U1695 (N_1695,In_963,In_1967);
and U1696 (N_1696,In_1593,In_2702);
and U1697 (N_1697,In_663,In_2024);
and U1698 (N_1698,In_2305,In_2788);
and U1699 (N_1699,In_2633,In_1044);
nand U1700 (N_1700,In_1025,In_1575);
and U1701 (N_1701,In_826,In_2319);
nor U1702 (N_1702,In_1558,In_2362);
nor U1703 (N_1703,In_2518,In_289);
nor U1704 (N_1704,In_2137,In_86);
xnor U1705 (N_1705,In_1486,In_1699);
xor U1706 (N_1706,In_1609,In_2400);
and U1707 (N_1707,In_2852,In_1012);
nor U1708 (N_1708,In_366,In_1372);
or U1709 (N_1709,In_1600,In_2397);
nand U1710 (N_1710,In_654,In_403);
and U1711 (N_1711,In_1455,In_774);
nor U1712 (N_1712,In_506,In_308);
nand U1713 (N_1713,In_406,In_630);
nor U1714 (N_1714,In_1668,In_535);
nand U1715 (N_1715,In_1385,In_1421);
nor U1716 (N_1716,In_1233,In_1017);
or U1717 (N_1717,In_493,In_2945);
and U1718 (N_1718,In_1943,In_125);
nand U1719 (N_1719,In_134,In_1151);
xor U1720 (N_1720,In_2116,In_546);
nor U1721 (N_1721,In_1604,In_1270);
nand U1722 (N_1722,In_2537,In_2160);
or U1723 (N_1723,In_1350,In_2880);
and U1724 (N_1724,In_804,In_1419);
xnor U1725 (N_1725,In_2308,In_2624);
xnor U1726 (N_1726,In_919,In_348);
nor U1727 (N_1727,In_25,In_2440);
nand U1728 (N_1728,In_480,In_1585);
nand U1729 (N_1729,In_351,In_2571);
nand U1730 (N_1730,In_1600,In_455);
and U1731 (N_1731,In_1806,In_2452);
nand U1732 (N_1732,In_954,In_661);
or U1733 (N_1733,In_2012,In_1035);
nor U1734 (N_1734,In_2963,In_46);
or U1735 (N_1735,In_381,In_1400);
and U1736 (N_1736,In_2123,In_2259);
xnor U1737 (N_1737,In_1952,In_2139);
or U1738 (N_1738,In_332,In_0);
and U1739 (N_1739,In_1275,In_2253);
xor U1740 (N_1740,In_1867,In_441);
nor U1741 (N_1741,In_1183,In_694);
or U1742 (N_1742,In_2761,In_1363);
or U1743 (N_1743,In_1334,In_2405);
or U1744 (N_1744,In_1395,In_2430);
nand U1745 (N_1745,In_1619,In_539);
nand U1746 (N_1746,In_1344,In_2028);
or U1747 (N_1747,In_2026,In_191);
and U1748 (N_1748,In_1770,In_1560);
nor U1749 (N_1749,In_910,In_1065);
xor U1750 (N_1750,In_25,In_586);
nand U1751 (N_1751,In_1753,In_860);
and U1752 (N_1752,In_2484,In_2792);
and U1753 (N_1753,In_902,In_1071);
nor U1754 (N_1754,In_2456,In_2472);
nand U1755 (N_1755,In_1506,In_893);
nor U1756 (N_1756,In_447,In_285);
nand U1757 (N_1757,In_2833,In_519);
nor U1758 (N_1758,In_2535,In_958);
nand U1759 (N_1759,In_1493,In_933);
xnor U1760 (N_1760,In_754,In_1396);
and U1761 (N_1761,In_2569,In_1831);
and U1762 (N_1762,In_1249,In_645);
nor U1763 (N_1763,In_410,In_350);
or U1764 (N_1764,In_685,In_2578);
xnor U1765 (N_1765,In_2834,In_550);
nand U1766 (N_1766,In_654,In_2175);
and U1767 (N_1767,In_736,In_1107);
nor U1768 (N_1768,In_340,In_301);
or U1769 (N_1769,In_2942,In_2375);
nor U1770 (N_1770,In_2611,In_1841);
nand U1771 (N_1771,In_1001,In_1532);
xor U1772 (N_1772,In_1955,In_527);
and U1773 (N_1773,In_1502,In_1043);
or U1774 (N_1774,In_1050,In_1015);
nor U1775 (N_1775,In_2635,In_626);
and U1776 (N_1776,In_1982,In_866);
xor U1777 (N_1777,In_1148,In_173);
nor U1778 (N_1778,In_2414,In_272);
xor U1779 (N_1779,In_1612,In_191);
or U1780 (N_1780,In_999,In_2294);
nor U1781 (N_1781,In_323,In_1675);
or U1782 (N_1782,In_2073,In_2328);
nor U1783 (N_1783,In_2712,In_234);
nor U1784 (N_1784,In_1554,In_547);
and U1785 (N_1785,In_1427,In_1414);
and U1786 (N_1786,In_1321,In_815);
nor U1787 (N_1787,In_2068,In_1865);
xor U1788 (N_1788,In_1974,In_254);
or U1789 (N_1789,In_2304,In_560);
xor U1790 (N_1790,In_548,In_791);
nand U1791 (N_1791,In_884,In_2623);
or U1792 (N_1792,In_1713,In_2879);
nand U1793 (N_1793,In_1870,In_2875);
nand U1794 (N_1794,In_2764,In_2708);
nor U1795 (N_1795,In_1503,In_2536);
xnor U1796 (N_1796,In_1102,In_1917);
or U1797 (N_1797,In_1889,In_2074);
xnor U1798 (N_1798,In_1244,In_546);
and U1799 (N_1799,In_2764,In_2811);
or U1800 (N_1800,In_2530,In_1508);
or U1801 (N_1801,In_2453,In_2860);
nand U1802 (N_1802,In_1470,In_1071);
xnor U1803 (N_1803,In_248,In_1713);
xor U1804 (N_1804,In_514,In_763);
xor U1805 (N_1805,In_20,In_210);
and U1806 (N_1806,In_568,In_640);
and U1807 (N_1807,In_2384,In_2700);
nor U1808 (N_1808,In_798,In_88);
nand U1809 (N_1809,In_1927,In_674);
nor U1810 (N_1810,In_142,In_247);
xor U1811 (N_1811,In_2030,In_2473);
and U1812 (N_1812,In_1525,In_2746);
nand U1813 (N_1813,In_399,In_769);
nor U1814 (N_1814,In_1212,In_2719);
nor U1815 (N_1815,In_668,In_2749);
and U1816 (N_1816,In_2546,In_2718);
nand U1817 (N_1817,In_1748,In_2222);
and U1818 (N_1818,In_2496,In_155);
nand U1819 (N_1819,In_2560,In_1456);
xor U1820 (N_1820,In_421,In_1833);
nand U1821 (N_1821,In_2918,In_1942);
and U1822 (N_1822,In_94,In_1388);
nor U1823 (N_1823,In_1865,In_234);
nand U1824 (N_1824,In_2787,In_2667);
nor U1825 (N_1825,In_463,In_1071);
nand U1826 (N_1826,In_1220,In_2131);
nor U1827 (N_1827,In_6,In_103);
nand U1828 (N_1828,In_1325,In_2883);
nor U1829 (N_1829,In_100,In_1833);
nor U1830 (N_1830,In_98,In_869);
xnor U1831 (N_1831,In_788,In_973);
xnor U1832 (N_1832,In_851,In_2726);
and U1833 (N_1833,In_1657,In_2354);
xnor U1834 (N_1834,In_2264,In_2196);
and U1835 (N_1835,In_2196,In_1881);
xor U1836 (N_1836,In_2761,In_56);
nand U1837 (N_1837,In_1497,In_1056);
and U1838 (N_1838,In_518,In_2382);
and U1839 (N_1839,In_2922,In_2825);
or U1840 (N_1840,In_2586,In_1729);
or U1841 (N_1841,In_314,In_1791);
nor U1842 (N_1842,In_1227,In_2282);
and U1843 (N_1843,In_2119,In_2246);
nand U1844 (N_1844,In_552,In_2916);
nor U1845 (N_1845,In_2725,In_1288);
or U1846 (N_1846,In_1126,In_2041);
xnor U1847 (N_1847,In_2685,In_1211);
and U1848 (N_1848,In_2140,In_2991);
nand U1849 (N_1849,In_1095,In_1077);
nor U1850 (N_1850,In_1123,In_1980);
or U1851 (N_1851,In_2692,In_152);
nor U1852 (N_1852,In_2093,In_1042);
nand U1853 (N_1853,In_2887,In_707);
nand U1854 (N_1854,In_1890,In_2802);
or U1855 (N_1855,In_49,In_1848);
and U1856 (N_1856,In_2394,In_1005);
and U1857 (N_1857,In_1874,In_2709);
and U1858 (N_1858,In_247,In_1098);
and U1859 (N_1859,In_2471,In_1327);
xnor U1860 (N_1860,In_2588,In_603);
and U1861 (N_1861,In_776,In_2501);
nand U1862 (N_1862,In_148,In_2768);
nor U1863 (N_1863,In_1093,In_795);
nand U1864 (N_1864,In_1202,In_525);
or U1865 (N_1865,In_2511,In_1320);
and U1866 (N_1866,In_1023,In_54);
nand U1867 (N_1867,In_2065,In_1317);
and U1868 (N_1868,In_2256,In_2497);
nor U1869 (N_1869,In_942,In_445);
nor U1870 (N_1870,In_2483,In_400);
and U1871 (N_1871,In_114,In_2386);
nor U1872 (N_1872,In_2323,In_2374);
or U1873 (N_1873,In_1816,In_2589);
and U1874 (N_1874,In_1177,In_395);
xor U1875 (N_1875,In_501,In_1776);
nor U1876 (N_1876,In_1263,In_365);
or U1877 (N_1877,In_2006,In_1874);
nor U1878 (N_1878,In_1795,In_2278);
and U1879 (N_1879,In_2521,In_1854);
nand U1880 (N_1880,In_714,In_495);
and U1881 (N_1881,In_429,In_2293);
nand U1882 (N_1882,In_2088,In_2296);
nor U1883 (N_1883,In_1780,In_779);
and U1884 (N_1884,In_1037,In_1222);
nor U1885 (N_1885,In_378,In_1507);
or U1886 (N_1886,In_98,In_277);
nand U1887 (N_1887,In_2492,In_2073);
and U1888 (N_1888,In_566,In_1596);
and U1889 (N_1889,In_2393,In_1183);
xnor U1890 (N_1890,In_1896,In_1378);
nand U1891 (N_1891,In_707,In_711);
or U1892 (N_1892,In_2412,In_2485);
nor U1893 (N_1893,In_1125,In_823);
or U1894 (N_1894,In_2439,In_1486);
nand U1895 (N_1895,In_2381,In_100);
nor U1896 (N_1896,In_225,In_560);
and U1897 (N_1897,In_649,In_1024);
nor U1898 (N_1898,In_1269,In_2274);
nand U1899 (N_1899,In_629,In_2580);
and U1900 (N_1900,In_1853,In_16);
xnor U1901 (N_1901,In_123,In_693);
nand U1902 (N_1902,In_1986,In_1963);
nor U1903 (N_1903,In_736,In_2686);
xnor U1904 (N_1904,In_1062,In_945);
nor U1905 (N_1905,In_1051,In_861);
or U1906 (N_1906,In_2217,In_2565);
and U1907 (N_1907,In_1152,In_2467);
nor U1908 (N_1908,In_1237,In_2138);
nor U1909 (N_1909,In_2922,In_353);
nand U1910 (N_1910,In_2436,In_1415);
nor U1911 (N_1911,In_1756,In_1034);
and U1912 (N_1912,In_437,In_1259);
nor U1913 (N_1913,In_2030,In_689);
nor U1914 (N_1914,In_2103,In_31);
xor U1915 (N_1915,In_2951,In_1455);
or U1916 (N_1916,In_428,In_1222);
or U1917 (N_1917,In_322,In_2645);
nor U1918 (N_1918,In_2853,In_2204);
or U1919 (N_1919,In_1699,In_1394);
and U1920 (N_1920,In_155,In_474);
nand U1921 (N_1921,In_2186,In_2644);
xnor U1922 (N_1922,In_323,In_1950);
or U1923 (N_1923,In_1219,In_2713);
nor U1924 (N_1924,In_1409,In_1275);
nand U1925 (N_1925,In_435,In_2548);
nor U1926 (N_1926,In_810,In_151);
and U1927 (N_1927,In_2206,In_2222);
nor U1928 (N_1928,In_2659,In_789);
and U1929 (N_1929,In_450,In_247);
xor U1930 (N_1930,In_1243,In_118);
nor U1931 (N_1931,In_2605,In_522);
and U1932 (N_1932,In_346,In_2680);
xor U1933 (N_1933,In_692,In_2061);
nor U1934 (N_1934,In_2406,In_2777);
nor U1935 (N_1935,In_719,In_1297);
xor U1936 (N_1936,In_293,In_1595);
and U1937 (N_1937,In_1422,In_1295);
and U1938 (N_1938,In_4,In_2891);
and U1939 (N_1939,In_58,In_1060);
xor U1940 (N_1940,In_2112,In_161);
xor U1941 (N_1941,In_328,In_1511);
or U1942 (N_1942,In_2301,In_506);
xnor U1943 (N_1943,In_2448,In_1658);
or U1944 (N_1944,In_2721,In_123);
or U1945 (N_1945,In_1455,In_2956);
or U1946 (N_1946,In_1700,In_1758);
xor U1947 (N_1947,In_2509,In_638);
or U1948 (N_1948,In_2353,In_1675);
and U1949 (N_1949,In_1990,In_2579);
or U1950 (N_1950,In_1268,In_975);
nand U1951 (N_1951,In_2180,In_1331);
xnor U1952 (N_1952,In_2915,In_2476);
nor U1953 (N_1953,In_1670,In_1480);
nand U1954 (N_1954,In_1393,In_1953);
xor U1955 (N_1955,In_1602,In_165);
and U1956 (N_1956,In_2419,In_1258);
and U1957 (N_1957,In_1117,In_2578);
nor U1958 (N_1958,In_35,In_1729);
xor U1959 (N_1959,In_1208,In_1600);
nand U1960 (N_1960,In_1765,In_1553);
or U1961 (N_1961,In_2593,In_1246);
and U1962 (N_1962,In_81,In_972);
xnor U1963 (N_1963,In_1673,In_458);
or U1964 (N_1964,In_523,In_2096);
nor U1965 (N_1965,In_114,In_218);
or U1966 (N_1966,In_1520,In_2965);
nand U1967 (N_1967,In_2722,In_402);
xor U1968 (N_1968,In_943,In_1650);
or U1969 (N_1969,In_574,In_2391);
and U1970 (N_1970,In_1226,In_2512);
or U1971 (N_1971,In_288,In_2221);
and U1972 (N_1972,In_2968,In_996);
or U1973 (N_1973,In_270,In_2238);
or U1974 (N_1974,In_1008,In_636);
nand U1975 (N_1975,In_1072,In_1592);
and U1976 (N_1976,In_1368,In_1149);
nand U1977 (N_1977,In_1694,In_2851);
nand U1978 (N_1978,In_1768,In_2159);
xnor U1979 (N_1979,In_2835,In_2435);
nor U1980 (N_1980,In_1797,In_272);
nor U1981 (N_1981,In_201,In_649);
nand U1982 (N_1982,In_317,In_2981);
xor U1983 (N_1983,In_1638,In_1899);
nand U1984 (N_1984,In_1082,In_906);
nor U1985 (N_1985,In_1702,In_1011);
or U1986 (N_1986,In_509,In_65);
nor U1987 (N_1987,In_132,In_979);
and U1988 (N_1988,In_2917,In_408);
xor U1989 (N_1989,In_502,In_662);
and U1990 (N_1990,In_786,In_21);
or U1991 (N_1991,In_1823,In_2561);
and U1992 (N_1992,In_157,In_738);
or U1993 (N_1993,In_725,In_1435);
xnor U1994 (N_1994,In_1223,In_2213);
xor U1995 (N_1995,In_1535,In_722);
nor U1996 (N_1996,In_1999,In_1761);
xor U1997 (N_1997,In_1072,In_2675);
xor U1998 (N_1998,In_1039,In_757);
nand U1999 (N_1999,In_2528,In_1881);
or U2000 (N_2000,In_1718,In_572);
nor U2001 (N_2001,In_51,In_530);
nor U2002 (N_2002,In_1605,In_1796);
and U2003 (N_2003,In_265,In_2469);
and U2004 (N_2004,In_2436,In_2412);
nor U2005 (N_2005,In_493,In_1409);
xnor U2006 (N_2006,In_875,In_1666);
xor U2007 (N_2007,In_884,In_2934);
nand U2008 (N_2008,In_2206,In_473);
nor U2009 (N_2009,In_459,In_2464);
nor U2010 (N_2010,In_2671,In_255);
nand U2011 (N_2011,In_1283,In_831);
or U2012 (N_2012,In_997,In_529);
nand U2013 (N_2013,In_1381,In_1610);
xnor U2014 (N_2014,In_2782,In_2719);
and U2015 (N_2015,In_2864,In_1642);
and U2016 (N_2016,In_169,In_1132);
nand U2017 (N_2017,In_1384,In_2191);
nor U2018 (N_2018,In_1804,In_154);
nor U2019 (N_2019,In_831,In_781);
and U2020 (N_2020,In_17,In_1945);
nor U2021 (N_2021,In_1370,In_1215);
xnor U2022 (N_2022,In_2715,In_1395);
nand U2023 (N_2023,In_836,In_1624);
nand U2024 (N_2024,In_1688,In_503);
nor U2025 (N_2025,In_684,In_1799);
nor U2026 (N_2026,In_999,In_1984);
or U2027 (N_2027,In_1604,In_1331);
or U2028 (N_2028,In_2381,In_925);
xor U2029 (N_2029,In_750,In_375);
nand U2030 (N_2030,In_1169,In_1261);
nor U2031 (N_2031,In_2441,In_1972);
xnor U2032 (N_2032,In_820,In_1148);
nand U2033 (N_2033,In_188,In_1098);
xor U2034 (N_2034,In_809,In_114);
nor U2035 (N_2035,In_2340,In_2631);
and U2036 (N_2036,In_551,In_588);
and U2037 (N_2037,In_455,In_1322);
xor U2038 (N_2038,In_71,In_85);
xor U2039 (N_2039,In_612,In_1140);
nand U2040 (N_2040,In_1387,In_2715);
nor U2041 (N_2041,In_1952,In_1035);
or U2042 (N_2042,In_1542,In_1467);
xnor U2043 (N_2043,In_1124,In_1451);
nand U2044 (N_2044,In_1812,In_2752);
and U2045 (N_2045,In_42,In_1528);
xnor U2046 (N_2046,In_78,In_2711);
and U2047 (N_2047,In_1063,In_662);
and U2048 (N_2048,In_2217,In_1167);
xnor U2049 (N_2049,In_2274,In_1129);
and U2050 (N_2050,In_2340,In_1213);
and U2051 (N_2051,In_2233,In_509);
or U2052 (N_2052,In_1431,In_1006);
or U2053 (N_2053,In_107,In_1797);
xnor U2054 (N_2054,In_1687,In_926);
nor U2055 (N_2055,In_533,In_2238);
nand U2056 (N_2056,In_1644,In_894);
nand U2057 (N_2057,In_2691,In_1948);
and U2058 (N_2058,In_2660,In_2590);
nand U2059 (N_2059,In_1208,In_2405);
xnor U2060 (N_2060,In_239,In_984);
xor U2061 (N_2061,In_2519,In_1956);
or U2062 (N_2062,In_2976,In_1225);
and U2063 (N_2063,In_2380,In_546);
nand U2064 (N_2064,In_2590,In_1152);
or U2065 (N_2065,In_1115,In_1611);
or U2066 (N_2066,In_611,In_2096);
or U2067 (N_2067,In_86,In_879);
nor U2068 (N_2068,In_1897,In_804);
xor U2069 (N_2069,In_2975,In_2424);
xnor U2070 (N_2070,In_1209,In_2957);
xor U2071 (N_2071,In_1319,In_1938);
or U2072 (N_2072,In_1627,In_2615);
nand U2073 (N_2073,In_705,In_1924);
xnor U2074 (N_2074,In_1015,In_1478);
nor U2075 (N_2075,In_2996,In_1253);
nor U2076 (N_2076,In_1876,In_2722);
nor U2077 (N_2077,In_1469,In_2829);
nor U2078 (N_2078,In_1866,In_2299);
and U2079 (N_2079,In_55,In_1169);
xor U2080 (N_2080,In_2836,In_2609);
and U2081 (N_2081,In_2212,In_1099);
nand U2082 (N_2082,In_2548,In_2645);
nand U2083 (N_2083,In_1465,In_2435);
and U2084 (N_2084,In_2213,In_432);
or U2085 (N_2085,In_2132,In_2790);
nand U2086 (N_2086,In_444,In_451);
nand U2087 (N_2087,In_2244,In_2488);
and U2088 (N_2088,In_1250,In_133);
nor U2089 (N_2089,In_1668,In_1877);
or U2090 (N_2090,In_204,In_1661);
nand U2091 (N_2091,In_1616,In_748);
xor U2092 (N_2092,In_293,In_1806);
nand U2093 (N_2093,In_1518,In_671);
or U2094 (N_2094,In_2284,In_1089);
xnor U2095 (N_2095,In_1057,In_2605);
xor U2096 (N_2096,In_779,In_2627);
xnor U2097 (N_2097,In_1260,In_1973);
and U2098 (N_2098,In_2328,In_1081);
nor U2099 (N_2099,In_917,In_582);
or U2100 (N_2100,In_432,In_797);
and U2101 (N_2101,In_38,In_1837);
and U2102 (N_2102,In_585,In_979);
and U2103 (N_2103,In_2747,In_2109);
nand U2104 (N_2104,In_2257,In_2696);
or U2105 (N_2105,In_2443,In_614);
or U2106 (N_2106,In_803,In_578);
or U2107 (N_2107,In_1781,In_1429);
xor U2108 (N_2108,In_635,In_1893);
nor U2109 (N_2109,In_2335,In_2712);
or U2110 (N_2110,In_1802,In_1923);
or U2111 (N_2111,In_1282,In_912);
nand U2112 (N_2112,In_60,In_1985);
nand U2113 (N_2113,In_2741,In_2531);
xor U2114 (N_2114,In_369,In_1149);
xor U2115 (N_2115,In_2094,In_2475);
nor U2116 (N_2116,In_503,In_541);
xnor U2117 (N_2117,In_1154,In_1572);
or U2118 (N_2118,In_925,In_47);
nand U2119 (N_2119,In_1742,In_2778);
or U2120 (N_2120,In_633,In_2534);
or U2121 (N_2121,In_1465,In_320);
and U2122 (N_2122,In_1747,In_1959);
or U2123 (N_2123,In_61,In_179);
nor U2124 (N_2124,In_859,In_147);
or U2125 (N_2125,In_70,In_596);
nor U2126 (N_2126,In_1597,In_1629);
or U2127 (N_2127,In_321,In_117);
xnor U2128 (N_2128,In_1943,In_1702);
and U2129 (N_2129,In_1,In_2073);
and U2130 (N_2130,In_2917,In_2065);
xnor U2131 (N_2131,In_72,In_1177);
or U2132 (N_2132,In_2206,In_614);
nand U2133 (N_2133,In_93,In_562);
and U2134 (N_2134,In_2007,In_2311);
or U2135 (N_2135,In_2300,In_1031);
or U2136 (N_2136,In_172,In_2978);
nand U2137 (N_2137,In_2649,In_108);
nand U2138 (N_2138,In_1561,In_2775);
and U2139 (N_2139,In_276,In_1322);
nor U2140 (N_2140,In_996,In_238);
nor U2141 (N_2141,In_157,In_1869);
nor U2142 (N_2142,In_383,In_1583);
nor U2143 (N_2143,In_2179,In_1484);
and U2144 (N_2144,In_1915,In_233);
and U2145 (N_2145,In_1615,In_547);
xnor U2146 (N_2146,In_2211,In_583);
or U2147 (N_2147,In_2143,In_488);
or U2148 (N_2148,In_1303,In_526);
nand U2149 (N_2149,In_1875,In_2547);
nor U2150 (N_2150,In_561,In_840);
or U2151 (N_2151,In_2770,In_2948);
or U2152 (N_2152,In_2449,In_1427);
or U2153 (N_2153,In_1360,In_1072);
nor U2154 (N_2154,In_399,In_44);
nand U2155 (N_2155,In_1222,In_997);
and U2156 (N_2156,In_662,In_705);
xor U2157 (N_2157,In_359,In_2461);
xnor U2158 (N_2158,In_500,In_50);
and U2159 (N_2159,In_697,In_1748);
nand U2160 (N_2160,In_1999,In_369);
and U2161 (N_2161,In_597,In_2454);
xor U2162 (N_2162,In_740,In_429);
nand U2163 (N_2163,In_1302,In_387);
nor U2164 (N_2164,In_717,In_16);
and U2165 (N_2165,In_822,In_955);
and U2166 (N_2166,In_2021,In_1543);
or U2167 (N_2167,In_2055,In_1096);
and U2168 (N_2168,In_522,In_2675);
xnor U2169 (N_2169,In_496,In_1904);
or U2170 (N_2170,In_562,In_2929);
and U2171 (N_2171,In_1502,In_1090);
and U2172 (N_2172,In_472,In_1639);
xnor U2173 (N_2173,In_2794,In_2218);
and U2174 (N_2174,In_882,In_1421);
nand U2175 (N_2175,In_1897,In_34);
xor U2176 (N_2176,In_1419,In_319);
or U2177 (N_2177,In_418,In_272);
and U2178 (N_2178,In_1781,In_198);
and U2179 (N_2179,In_2484,In_2566);
xnor U2180 (N_2180,In_2798,In_2566);
or U2181 (N_2181,In_2247,In_2893);
nand U2182 (N_2182,In_997,In_735);
xnor U2183 (N_2183,In_414,In_1015);
nor U2184 (N_2184,In_1694,In_540);
xnor U2185 (N_2185,In_1508,In_1315);
xnor U2186 (N_2186,In_126,In_2352);
nand U2187 (N_2187,In_751,In_1921);
or U2188 (N_2188,In_1187,In_546);
or U2189 (N_2189,In_2513,In_90);
nand U2190 (N_2190,In_2567,In_1431);
or U2191 (N_2191,In_2321,In_410);
and U2192 (N_2192,In_2250,In_2492);
xor U2193 (N_2193,In_2341,In_124);
or U2194 (N_2194,In_1947,In_2079);
xor U2195 (N_2195,In_265,In_2657);
nor U2196 (N_2196,In_670,In_1099);
xor U2197 (N_2197,In_2492,In_1315);
and U2198 (N_2198,In_732,In_2138);
or U2199 (N_2199,In_2913,In_332);
and U2200 (N_2200,In_2936,In_1875);
nor U2201 (N_2201,In_2185,In_795);
xor U2202 (N_2202,In_861,In_407);
xor U2203 (N_2203,In_637,In_1965);
nand U2204 (N_2204,In_2392,In_920);
xnor U2205 (N_2205,In_373,In_134);
nor U2206 (N_2206,In_196,In_832);
or U2207 (N_2207,In_2533,In_756);
nand U2208 (N_2208,In_531,In_1517);
nand U2209 (N_2209,In_53,In_2811);
nor U2210 (N_2210,In_36,In_1007);
and U2211 (N_2211,In_496,In_1299);
or U2212 (N_2212,In_946,In_2043);
or U2213 (N_2213,In_2312,In_370);
nor U2214 (N_2214,In_640,In_1005);
and U2215 (N_2215,In_1843,In_1195);
xor U2216 (N_2216,In_529,In_1802);
or U2217 (N_2217,In_1745,In_1101);
nand U2218 (N_2218,In_758,In_761);
xnor U2219 (N_2219,In_595,In_1681);
or U2220 (N_2220,In_2068,In_1493);
xnor U2221 (N_2221,In_845,In_1683);
nand U2222 (N_2222,In_932,In_1583);
xor U2223 (N_2223,In_1577,In_1188);
nor U2224 (N_2224,In_1962,In_414);
nand U2225 (N_2225,In_930,In_936);
nand U2226 (N_2226,In_1724,In_2083);
or U2227 (N_2227,In_552,In_1972);
xor U2228 (N_2228,In_539,In_555);
or U2229 (N_2229,In_1866,In_110);
nor U2230 (N_2230,In_1307,In_2828);
or U2231 (N_2231,In_1724,In_2237);
nand U2232 (N_2232,In_2473,In_897);
or U2233 (N_2233,In_2135,In_2778);
nand U2234 (N_2234,In_1858,In_1905);
nor U2235 (N_2235,In_2432,In_2163);
nand U2236 (N_2236,In_856,In_2122);
and U2237 (N_2237,In_2154,In_1099);
or U2238 (N_2238,In_1611,In_2714);
xor U2239 (N_2239,In_2004,In_1315);
nor U2240 (N_2240,In_2961,In_432);
or U2241 (N_2241,In_849,In_1816);
or U2242 (N_2242,In_659,In_2395);
or U2243 (N_2243,In_2167,In_60);
nor U2244 (N_2244,In_1475,In_1315);
and U2245 (N_2245,In_2077,In_179);
and U2246 (N_2246,In_111,In_1410);
or U2247 (N_2247,In_362,In_1213);
or U2248 (N_2248,In_999,In_51);
or U2249 (N_2249,In_2967,In_602);
or U2250 (N_2250,In_1042,In_1594);
nand U2251 (N_2251,In_1476,In_1580);
nor U2252 (N_2252,In_2599,In_1559);
nor U2253 (N_2253,In_2168,In_547);
nand U2254 (N_2254,In_1564,In_1582);
xnor U2255 (N_2255,In_1304,In_165);
and U2256 (N_2256,In_1421,In_1607);
nand U2257 (N_2257,In_2030,In_40);
xor U2258 (N_2258,In_486,In_1054);
and U2259 (N_2259,In_1918,In_1341);
nor U2260 (N_2260,In_1256,In_2317);
nand U2261 (N_2261,In_1159,In_1635);
xor U2262 (N_2262,In_43,In_153);
or U2263 (N_2263,In_1222,In_2307);
or U2264 (N_2264,In_1998,In_1267);
xnor U2265 (N_2265,In_789,In_1291);
and U2266 (N_2266,In_2791,In_1444);
nand U2267 (N_2267,In_1484,In_707);
and U2268 (N_2268,In_1945,In_2895);
or U2269 (N_2269,In_2621,In_1599);
nor U2270 (N_2270,In_2938,In_504);
nor U2271 (N_2271,In_1681,In_1642);
nor U2272 (N_2272,In_1363,In_1193);
xor U2273 (N_2273,In_368,In_2442);
and U2274 (N_2274,In_1504,In_2897);
nand U2275 (N_2275,In_1963,In_832);
and U2276 (N_2276,In_1827,In_561);
xnor U2277 (N_2277,In_824,In_1997);
or U2278 (N_2278,In_1622,In_1175);
nor U2279 (N_2279,In_500,In_1394);
or U2280 (N_2280,In_2048,In_2663);
nor U2281 (N_2281,In_1616,In_2070);
nor U2282 (N_2282,In_1023,In_974);
xor U2283 (N_2283,In_81,In_551);
nand U2284 (N_2284,In_1955,In_183);
and U2285 (N_2285,In_2455,In_201);
xor U2286 (N_2286,In_667,In_1117);
nor U2287 (N_2287,In_2630,In_928);
nor U2288 (N_2288,In_2152,In_2971);
or U2289 (N_2289,In_2520,In_2949);
and U2290 (N_2290,In_1833,In_796);
or U2291 (N_2291,In_1985,In_822);
xor U2292 (N_2292,In_2277,In_2933);
or U2293 (N_2293,In_2354,In_154);
nor U2294 (N_2294,In_2380,In_785);
nand U2295 (N_2295,In_1316,In_2036);
nor U2296 (N_2296,In_712,In_1688);
nand U2297 (N_2297,In_62,In_1643);
nand U2298 (N_2298,In_1415,In_1452);
and U2299 (N_2299,In_235,In_2553);
and U2300 (N_2300,In_21,In_1570);
nand U2301 (N_2301,In_1364,In_95);
nand U2302 (N_2302,In_380,In_232);
or U2303 (N_2303,In_563,In_944);
nand U2304 (N_2304,In_2879,In_1865);
xor U2305 (N_2305,In_2909,In_2160);
and U2306 (N_2306,In_2793,In_505);
nor U2307 (N_2307,In_869,In_1188);
or U2308 (N_2308,In_1532,In_1762);
or U2309 (N_2309,In_2577,In_1067);
nor U2310 (N_2310,In_288,In_1457);
and U2311 (N_2311,In_1306,In_908);
or U2312 (N_2312,In_1268,In_1702);
nand U2313 (N_2313,In_2266,In_689);
nand U2314 (N_2314,In_619,In_2124);
or U2315 (N_2315,In_1414,In_497);
or U2316 (N_2316,In_2194,In_1568);
nor U2317 (N_2317,In_680,In_565);
and U2318 (N_2318,In_2127,In_2977);
nand U2319 (N_2319,In_2095,In_1190);
and U2320 (N_2320,In_8,In_666);
xor U2321 (N_2321,In_953,In_2304);
and U2322 (N_2322,In_297,In_1442);
nand U2323 (N_2323,In_312,In_2821);
or U2324 (N_2324,In_2505,In_2448);
nor U2325 (N_2325,In_1614,In_331);
or U2326 (N_2326,In_1997,In_758);
and U2327 (N_2327,In_832,In_2223);
xnor U2328 (N_2328,In_1984,In_2075);
nor U2329 (N_2329,In_2749,In_2143);
xor U2330 (N_2330,In_2255,In_2646);
nand U2331 (N_2331,In_1962,In_462);
nor U2332 (N_2332,In_649,In_432);
nand U2333 (N_2333,In_1191,In_2584);
and U2334 (N_2334,In_1287,In_943);
xnor U2335 (N_2335,In_1350,In_1800);
xnor U2336 (N_2336,In_772,In_1637);
or U2337 (N_2337,In_493,In_622);
nor U2338 (N_2338,In_33,In_1743);
nand U2339 (N_2339,In_31,In_769);
and U2340 (N_2340,In_978,In_2302);
nand U2341 (N_2341,In_1781,In_1881);
or U2342 (N_2342,In_240,In_2408);
xor U2343 (N_2343,In_951,In_417);
nand U2344 (N_2344,In_2108,In_374);
and U2345 (N_2345,In_1537,In_2901);
nand U2346 (N_2346,In_2376,In_1812);
and U2347 (N_2347,In_2835,In_2558);
nor U2348 (N_2348,In_1330,In_896);
xor U2349 (N_2349,In_1526,In_1137);
nand U2350 (N_2350,In_2819,In_2577);
nand U2351 (N_2351,In_2526,In_1320);
xor U2352 (N_2352,In_914,In_630);
nor U2353 (N_2353,In_2024,In_2612);
or U2354 (N_2354,In_227,In_1998);
nor U2355 (N_2355,In_1413,In_1754);
nand U2356 (N_2356,In_1140,In_2751);
or U2357 (N_2357,In_2081,In_2314);
xnor U2358 (N_2358,In_679,In_1084);
nand U2359 (N_2359,In_2314,In_2660);
xor U2360 (N_2360,In_1393,In_1649);
nand U2361 (N_2361,In_392,In_2192);
or U2362 (N_2362,In_1257,In_85);
or U2363 (N_2363,In_924,In_1721);
or U2364 (N_2364,In_1619,In_1884);
or U2365 (N_2365,In_1859,In_649);
or U2366 (N_2366,In_822,In_2752);
and U2367 (N_2367,In_596,In_1971);
and U2368 (N_2368,In_2067,In_2781);
nor U2369 (N_2369,In_1719,In_2428);
or U2370 (N_2370,In_250,In_1048);
nand U2371 (N_2371,In_637,In_33);
nor U2372 (N_2372,In_2583,In_950);
nor U2373 (N_2373,In_157,In_2516);
nand U2374 (N_2374,In_1272,In_1166);
or U2375 (N_2375,In_1948,In_1702);
or U2376 (N_2376,In_323,In_1628);
or U2377 (N_2377,In_1461,In_1365);
or U2378 (N_2378,In_1751,In_936);
xor U2379 (N_2379,In_2893,In_1379);
nand U2380 (N_2380,In_711,In_2727);
nand U2381 (N_2381,In_2718,In_2694);
nor U2382 (N_2382,In_1881,In_2333);
xor U2383 (N_2383,In_574,In_2928);
nand U2384 (N_2384,In_909,In_2310);
or U2385 (N_2385,In_843,In_2622);
or U2386 (N_2386,In_2941,In_73);
or U2387 (N_2387,In_1413,In_2813);
and U2388 (N_2388,In_1337,In_565);
nor U2389 (N_2389,In_2049,In_2241);
xor U2390 (N_2390,In_1503,In_61);
or U2391 (N_2391,In_800,In_834);
xor U2392 (N_2392,In_1339,In_2246);
or U2393 (N_2393,In_574,In_1061);
xor U2394 (N_2394,In_1903,In_1976);
and U2395 (N_2395,In_2318,In_922);
xnor U2396 (N_2396,In_40,In_1327);
nor U2397 (N_2397,In_1154,In_2835);
and U2398 (N_2398,In_1207,In_329);
xnor U2399 (N_2399,In_1620,In_1398);
xor U2400 (N_2400,In_1513,In_1508);
xnor U2401 (N_2401,In_1407,In_1231);
nand U2402 (N_2402,In_1734,In_110);
and U2403 (N_2403,In_2812,In_153);
or U2404 (N_2404,In_1463,In_224);
and U2405 (N_2405,In_972,In_813);
xnor U2406 (N_2406,In_137,In_2573);
nand U2407 (N_2407,In_1263,In_373);
and U2408 (N_2408,In_1411,In_1152);
xnor U2409 (N_2409,In_877,In_2826);
nand U2410 (N_2410,In_1569,In_62);
or U2411 (N_2411,In_2489,In_1095);
nor U2412 (N_2412,In_2552,In_1616);
nand U2413 (N_2413,In_905,In_2474);
nor U2414 (N_2414,In_984,In_190);
nor U2415 (N_2415,In_1717,In_224);
or U2416 (N_2416,In_2949,In_2010);
nand U2417 (N_2417,In_2932,In_1917);
xnor U2418 (N_2418,In_1653,In_851);
or U2419 (N_2419,In_2735,In_1944);
nor U2420 (N_2420,In_2643,In_703);
nand U2421 (N_2421,In_2642,In_503);
or U2422 (N_2422,In_1187,In_2837);
or U2423 (N_2423,In_240,In_1277);
xnor U2424 (N_2424,In_801,In_2732);
or U2425 (N_2425,In_2058,In_2921);
xnor U2426 (N_2426,In_508,In_1830);
xor U2427 (N_2427,In_673,In_1974);
xnor U2428 (N_2428,In_248,In_2146);
and U2429 (N_2429,In_1505,In_274);
and U2430 (N_2430,In_648,In_2639);
xnor U2431 (N_2431,In_1891,In_155);
xor U2432 (N_2432,In_2229,In_2140);
and U2433 (N_2433,In_186,In_1902);
and U2434 (N_2434,In_1075,In_2604);
nor U2435 (N_2435,In_2464,In_1776);
or U2436 (N_2436,In_276,In_885);
xor U2437 (N_2437,In_276,In_2309);
and U2438 (N_2438,In_202,In_2061);
or U2439 (N_2439,In_2897,In_2301);
nand U2440 (N_2440,In_97,In_1287);
and U2441 (N_2441,In_2596,In_1684);
and U2442 (N_2442,In_704,In_1528);
xor U2443 (N_2443,In_933,In_209);
xnor U2444 (N_2444,In_956,In_2539);
and U2445 (N_2445,In_828,In_1037);
or U2446 (N_2446,In_822,In_2243);
nor U2447 (N_2447,In_2206,In_2382);
and U2448 (N_2448,In_2394,In_842);
or U2449 (N_2449,In_1663,In_388);
nor U2450 (N_2450,In_1751,In_156);
nand U2451 (N_2451,In_1659,In_1442);
nor U2452 (N_2452,In_1977,In_85);
or U2453 (N_2453,In_1731,In_700);
xnor U2454 (N_2454,In_1318,In_1970);
nand U2455 (N_2455,In_2540,In_656);
nand U2456 (N_2456,In_759,In_2900);
xor U2457 (N_2457,In_1903,In_2538);
nor U2458 (N_2458,In_716,In_2020);
or U2459 (N_2459,In_943,In_1141);
or U2460 (N_2460,In_1124,In_974);
and U2461 (N_2461,In_1902,In_2613);
and U2462 (N_2462,In_400,In_928);
nand U2463 (N_2463,In_1219,In_534);
xor U2464 (N_2464,In_243,In_1855);
or U2465 (N_2465,In_943,In_2324);
nor U2466 (N_2466,In_763,In_1114);
or U2467 (N_2467,In_602,In_2334);
and U2468 (N_2468,In_373,In_1689);
or U2469 (N_2469,In_96,In_2479);
or U2470 (N_2470,In_74,In_385);
or U2471 (N_2471,In_2043,In_942);
xnor U2472 (N_2472,In_740,In_629);
nand U2473 (N_2473,In_2917,In_539);
nor U2474 (N_2474,In_1943,In_1569);
xnor U2475 (N_2475,In_976,In_1486);
nor U2476 (N_2476,In_2598,In_2917);
nor U2477 (N_2477,In_1087,In_2686);
or U2478 (N_2478,In_1022,In_1745);
and U2479 (N_2479,In_2824,In_1860);
nand U2480 (N_2480,In_1057,In_2819);
or U2481 (N_2481,In_163,In_140);
or U2482 (N_2482,In_2347,In_1100);
and U2483 (N_2483,In_1905,In_150);
nand U2484 (N_2484,In_968,In_2288);
or U2485 (N_2485,In_2533,In_1061);
and U2486 (N_2486,In_2626,In_312);
or U2487 (N_2487,In_1206,In_2552);
nor U2488 (N_2488,In_633,In_886);
nor U2489 (N_2489,In_817,In_2863);
nand U2490 (N_2490,In_534,In_231);
xor U2491 (N_2491,In_2978,In_1935);
and U2492 (N_2492,In_802,In_153);
nor U2493 (N_2493,In_730,In_453);
xnor U2494 (N_2494,In_2706,In_2452);
nor U2495 (N_2495,In_2721,In_1979);
nor U2496 (N_2496,In_879,In_2032);
xnor U2497 (N_2497,In_2997,In_2200);
nand U2498 (N_2498,In_2656,In_2271);
nor U2499 (N_2499,In_633,In_988);
and U2500 (N_2500,In_2011,In_1657);
or U2501 (N_2501,In_799,In_2506);
nand U2502 (N_2502,In_2586,In_1107);
nor U2503 (N_2503,In_1204,In_1249);
or U2504 (N_2504,In_746,In_890);
and U2505 (N_2505,In_1418,In_1309);
nor U2506 (N_2506,In_1965,In_1912);
nand U2507 (N_2507,In_944,In_2413);
xor U2508 (N_2508,In_424,In_193);
and U2509 (N_2509,In_2192,In_844);
and U2510 (N_2510,In_339,In_1294);
xor U2511 (N_2511,In_2398,In_1398);
and U2512 (N_2512,In_530,In_1658);
nand U2513 (N_2513,In_1824,In_1131);
xor U2514 (N_2514,In_453,In_215);
or U2515 (N_2515,In_2536,In_2349);
and U2516 (N_2516,In_1495,In_27);
nand U2517 (N_2517,In_1663,In_125);
or U2518 (N_2518,In_1603,In_2253);
and U2519 (N_2519,In_604,In_110);
nor U2520 (N_2520,In_2930,In_2096);
nor U2521 (N_2521,In_262,In_1041);
or U2522 (N_2522,In_1243,In_2055);
nand U2523 (N_2523,In_1567,In_2674);
nand U2524 (N_2524,In_1038,In_162);
nand U2525 (N_2525,In_475,In_921);
and U2526 (N_2526,In_1952,In_2542);
nor U2527 (N_2527,In_1672,In_2073);
xnor U2528 (N_2528,In_1764,In_2201);
xor U2529 (N_2529,In_939,In_253);
and U2530 (N_2530,In_1260,In_2033);
and U2531 (N_2531,In_1971,In_719);
nand U2532 (N_2532,In_923,In_1815);
nand U2533 (N_2533,In_1716,In_2196);
xnor U2534 (N_2534,In_681,In_836);
nand U2535 (N_2535,In_709,In_1975);
xor U2536 (N_2536,In_1677,In_1204);
nor U2537 (N_2537,In_2621,In_33);
and U2538 (N_2538,In_2892,In_993);
or U2539 (N_2539,In_2866,In_1861);
xor U2540 (N_2540,In_2239,In_2359);
xnor U2541 (N_2541,In_1369,In_393);
and U2542 (N_2542,In_2560,In_2890);
nor U2543 (N_2543,In_2084,In_151);
xnor U2544 (N_2544,In_1767,In_756);
nor U2545 (N_2545,In_1049,In_1652);
nor U2546 (N_2546,In_718,In_2435);
or U2547 (N_2547,In_141,In_2819);
nor U2548 (N_2548,In_237,In_2473);
nor U2549 (N_2549,In_42,In_2994);
nand U2550 (N_2550,In_2888,In_1885);
or U2551 (N_2551,In_324,In_1035);
or U2552 (N_2552,In_1985,In_1808);
nand U2553 (N_2553,In_1888,In_1784);
xor U2554 (N_2554,In_1845,In_2787);
nor U2555 (N_2555,In_1581,In_1764);
nor U2556 (N_2556,In_2860,In_857);
nor U2557 (N_2557,In_904,In_99);
xnor U2558 (N_2558,In_1402,In_1589);
or U2559 (N_2559,In_1354,In_292);
xor U2560 (N_2560,In_955,In_781);
nor U2561 (N_2561,In_824,In_2094);
or U2562 (N_2562,In_1390,In_2852);
or U2563 (N_2563,In_1610,In_2826);
nand U2564 (N_2564,In_2428,In_2282);
or U2565 (N_2565,In_2501,In_2969);
xor U2566 (N_2566,In_994,In_2616);
and U2567 (N_2567,In_1279,In_2380);
and U2568 (N_2568,In_540,In_1212);
nand U2569 (N_2569,In_2238,In_2388);
xor U2570 (N_2570,In_1337,In_721);
or U2571 (N_2571,In_168,In_2768);
or U2572 (N_2572,In_445,In_2933);
nor U2573 (N_2573,In_813,In_1353);
nor U2574 (N_2574,In_883,In_900);
or U2575 (N_2575,In_505,In_931);
or U2576 (N_2576,In_2130,In_1660);
nor U2577 (N_2577,In_1872,In_1043);
or U2578 (N_2578,In_1723,In_1112);
nor U2579 (N_2579,In_491,In_2194);
xor U2580 (N_2580,In_1198,In_2324);
or U2581 (N_2581,In_249,In_892);
xnor U2582 (N_2582,In_61,In_1791);
nand U2583 (N_2583,In_1648,In_1448);
nor U2584 (N_2584,In_2186,In_2739);
xnor U2585 (N_2585,In_124,In_208);
nand U2586 (N_2586,In_1212,In_326);
nor U2587 (N_2587,In_2783,In_2419);
nand U2588 (N_2588,In_855,In_521);
xnor U2589 (N_2589,In_52,In_1920);
or U2590 (N_2590,In_1086,In_389);
xor U2591 (N_2591,In_2359,In_802);
nand U2592 (N_2592,In_2049,In_1631);
and U2593 (N_2593,In_1154,In_1637);
or U2594 (N_2594,In_337,In_897);
nand U2595 (N_2595,In_2383,In_2586);
or U2596 (N_2596,In_2767,In_712);
xnor U2597 (N_2597,In_1169,In_650);
or U2598 (N_2598,In_1651,In_2004);
xor U2599 (N_2599,In_2,In_2017);
nor U2600 (N_2600,In_1111,In_1779);
nor U2601 (N_2601,In_2767,In_1936);
xor U2602 (N_2602,In_543,In_2876);
nor U2603 (N_2603,In_964,In_550);
nor U2604 (N_2604,In_2630,In_354);
xnor U2605 (N_2605,In_2631,In_1198);
nand U2606 (N_2606,In_2807,In_639);
and U2607 (N_2607,In_1131,In_2201);
nand U2608 (N_2608,In_614,In_1128);
or U2609 (N_2609,In_2935,In_622);
or U2610 (N_2610,In_2611,In_2651);
xor U2611 (N_2611,In_2346,In_73);
nand U2612 (N_2612,In_473,In_2975);
nand U2613 (N_2613,In_1521,In_1082);
and U2614 (N_2614,In_2033,In_1447);
xor U2615 (N_2615,In_1698,In_1347);
nand U2616 (N_2616,In_1109,In_2820);
xor U2617 (N_2617,In_2700,In_291);
nand U2618 (N_2618,In_1927,In_2370);
nand U2619 (N_2619,In_1017,In_1949);
nand U2620 (N_2620,In_295,In_2614);
and U2621 (N_2621,In_2641,In_433);
xor U2622 (N_2622,In_1483,In_2932);
and U2623 (N_2623,In_513,In_813);
or U2624 (N_2624,In_1803,In_432);
nand U2625 (N_2625,In_1024,In_2058);
nor U2626 (N_2626,In_1137,In_1743);
and U2627 (N_2627,In_2058,In_663);
or U2628 (N_2628,In_1061,In_1950);
or U2629 (N_2629,In_842,In_1302);
or U2630 (N_2630,In_1362,In_1263);
and U2631 (N_2631,In_936,In_1499);
or U2632 (N_2632,In_129,In_581);
nand U2633 (N_2633,In_1604,In_983);
nand U2634 (N_2634,In_2537,In_1295);
nor U2635 (N_2635,In_277,In_1088);
and U2636 (N_2636,In_2622,In_2127);
xnor U2637 (N_2637,In_955,In_1379);
or U2638 (N_2638,In_1057,In_1519);
or U2639 (N_2639,In_2944,In_1559);
or U2640 (N_2640,In_326,In_1472);
nor U2641 (N_2641,In_809,In_555);
or U2642 (N_2642,In_332,In_1012);
nand U2643 (N_2643,In_1438,In_1829);
nand U2644 (N_2644,In_1467,In_1780);
and U2645 (N_2645,In_903,In_2785);
nor U2646 (N_2646,In_1975,In_1883);
xor U2647 (N_2647,In_822,In_444);
nand U2648 (N_2648,In_2628,In_2945);
nor U2649 (N_2649,In_876,In_1163);
xnor U2650 (N_2650,In_1823,In_800);
or U2651 (N_2651,In_573,In_701);
nor U2652 (N_2652,In_660,In_1363);
and U2653 (N_2653,In_264,In_271);
xnor U2654 (N_2654,In_460,In_1431);
or U2655 (N_2655,In_1795,In_879);
or U2656 (N_2656,In_1219,In_1376);
or U2657 (N_2657,In_2349,In_2304);
and U2658 (N_2658,In_2517,In_936);
nand U2659 (N_2659,In_2350,In_784);
or U2660 (N_2660,In_1971,In_2163);
or U2661 (N_2661,In_1020,In_567);
and U2662 (N_2662,In_986,In_188);
or U2663 (N_2663,In_1746,In_1095);
or U2664 (N_2664,In_56,In_417);
xnor U2665 (N_2665,In_1073,In_1509);
nand U2666 (N_2666,In_1511,In_1534);
nor U2667 (N_2667,In_420,In_416);
or U2668 (N_2668,In_1123,In_2782);
xnor U2669 (N_2669,In_203,In_521);
xor U2670 (N_2670,In_663,In_2524);
or U2671 (N_2671,In_2866,In_1029);
nor U2672 (N_2672,In_919,In_1370);
xor U2673 (N_2673,In_383,In_1661);
xor U2674 (N_2674,In_424,In_2916);
or U2675 (N_2675,In_574,In_1788);
nor U2676 (N_2676,In_1879,In_2760);
or U2677 (N_2677,In_1255,In_747);
and U2678 (N_2678,In_1474,In_630);
or U2679 (N_2679,In_2629,In_2760);
nor U2680 (N_2680,In_1698,In_534);
or U2681 (N_2681,In_860,In_2784);
or U2682 (N_2682,In_1798,In_2339);
nand U2683 (N_2683,In_206,In_57);
xnor U2684 (N_2684,In_2463,In_67);
or U2685 (N_2685,In_911,In_1557);
or U2686 (N_2686,In_2803,In_365);
nor U2687 (N_2687,In_2526,In_410);
and U2688 (N_2688,In_1285,In_1173);
or U2689 (N_2689,In_910,In_2029);
xnor U2690 (N_2690,In_18,In_1052);
nand U2691 (N_2691,In_528,In_1971);
xnor U2692 (N_2692,In_767,In_1025);
or U2693 (N_2693,In_2951,In_1696);
xnor U2694 (N_2694,In_2470,In_604);
or U2695 (N_2695,In_423,In_1413);
and U2696 (N_2696,In_2318,In_355);
xnor U2697 (N_2697,In_2641,In_301);
xnor U2698 (N_2698,In_1783,In_557);
nand U2699 (N_2699,In_94,In_479);
nor U2700 (N_2700,In_1200,In_291);
or U2701 (N_2701,In_1260,In_1035);
xnor U2702 (N_2702,In_1739,In_1242);
or U2703 (N_2703,In_1066,In_756);
nand U2704 (N_2704,In_1283,In_1671);
nor U2705 (N_2705,In_2520,In_2866);
and U2706 (N_2706,In_611,In_2467);
nand U2707 (N_2707,In_1454,In_841);
and U2708 (N_2708,In_2731,In_495);
xor U2709 (N_2709,In_2069,In_1183);
nand U2710 (N_2710,In_329,In_2059);
and U2711 (N_2711,In_2555,In_1718);
or U2712 (N_2712,In_970,In_2671);
nor U2713 (N_2713,In_2759,In_1238);
xor U2714 (N_2714,In_2622,In_2789);
and U2715 (N_2715,In_1843,In_1753);
or U2716 (N_2716,In_2998,In_551);
or U2717 (N_2717,In_2276,In_613);
xnor U2718 (N_2718,In_1140,In_1341);
and U2719 (N_2719,In_2177,In_1843);
xor U2720 (N_2720,In_1876,In_388);
and U2721 (N_2721,In_909,In_1979);
or U2722 (N_2722,In_2985,In_868);
nand U2723 (N_2723,In_2386,In_1043);
or U2724 (N_2724,In_1096,In_643);
nand U2725 (N_2725,In_229,In_2303);
and U2726 (N_2726,In_2791,In_370);
nor U2727 (N_2727,In_1634,In_2064);
nor U2728 (N_2728,In_403,In_76);
or U2729 (N_2729,In_1520,In_1037);
nor U2730 (N_2730,In_983,In_873);
xor U2731 (N_2731,In_422,In_792);
nand U2732 (N_2732,In_1407,In_1178);
xor U2733 (N_2733,In_55,In_1789);
nor U2734 (N_2734,In_1578,In_2261);
nor U2735 (N_2735,In_232,In_595);
and U2736 (N_2736,In_678,In_1001);
nor U2737 (N_2737,In_1674,In_1247);
xor U2738 (N_2738,In_386,In_874);
nand U2739 (N_2739,In_1427,In_1370);
nor U2740 (N_2740,In_553,In_401);
or U2741 (N_2741,In_131,In_1434);
nor U2742 (N_2742,In_752,In_2623);
nand U2743 (N_2743,In_1882,In_608);
or U2744 (N_2744,In_2757,In_2916);
and U2745 (N_2745,In_555,In_2206);
xor U2746 (N_2746,In_720,In_747);
nand U2747 (N_2747,In_755,In_2203);
nand U2748 (N_2748,In_916,In_1679);
nor U2749 (N_2749,In_1237,In_2488);
xor U2750 (N_2750,In_264,In_118);
and U2751 (N_2751,In_1530,In_89);
nor U2752 (N_2752,In_91,In_699);
xnor U2753 (N_2753,In_723,In_609);
xnor U2754 (N_2754,In_2332,In_869);
or U2755 (N_2755,In_1823,In_2281);
nand U2756 (N_2756,In_2678,In_372);
and U2757 (N_2757,In_148,In_787);
and U2758 (N_2758,In_1563,In_1321);
and U2759 (N_2759,In_470,In_26);
nor U2760 (N_2760,In_2929,In_1088);
nand U2761 (N_2761,In_2917,In_1878);
or U2762 (N_2762,In_1736,In_2563);
and U2763 (N_2763,In_1266,In_1271);
or U2764 (N_2764,In_1473,In_2664);
nor U2765 (N_2765,In_2417,In_641);
nor U2766 (N_2766,In_348,In_1577);
nor U2767 (N_2767,In_76,In_2480);
nor U2768 (N_2768,In_211,In_1358);
xnor U2769 (N_2769,In_668,In_869);
xnor U2770 (N_2770,In_1666,In_1692);
xnor U2771 (N_2771,In_1392,In_2508);
nand U2772 (N_2772,In_2035,In_536);
and U2773 (N_2773,In_1337,In_442);
or U2774 (N_2774,In_1236,In_1943);
or U2775 (N_2775,In_342,In_148);
nor U2776 (N_2776,In_433,In_157);
xnor U2777 (N_2777,In_2782,In_739);
nand U2778 (N_2778,In_562,In_2488);
nor U2779 (N_2779,In_1991,In_2769);
xor U2780 (N_2780,In_2667,In_2986);
xor U2781 (N_2781,In_1419,In_1153);
nand U2782 (N_2782,In_2324,In_2816);
nand U2783 (N_2783,In_2213,In_1509);
nor U2784 (N_2784,In_1248,In_74);
xnor U2785 (N_2785,In_1307,In_1099);
nor U2786 (N_2786,In_1697,In_2748);
or U2787 (N_2787,In_1443,In_2045);
and U2788 (N_2788,In_1501,In_1484);
or U2789 (N_2789,In_2761,In_27);
xor U2790 (N_2790,In_2513,In_1266);
or U2791 (N_2791,In_2598,In_2200);
nor U2792 (N_2792,In_1540,In_374);
and U2793 (N_2793,In_2113,In_1561);
nor U2794 (N_2794,In_443,In_2412);
or U2795 (N_2795,In_2648,In_108);
or U2796 (N_2796,In_1526,In_2613);
nand U2797 (N_2797,In_2666,In_2059);
nand U2798 (N_2798,In_1875,In_1231);
nand U2799 (N_2799,In_1045,In_1708);
and U2800 (N_2800,In_726,In_2546);
nor U2801 (N_2801,In_2643,In_1872);
xnor U2802 (N_2802,In_2910,In_2991);
nor U2803 (N_2803,In_939,In_1767);
nor U2804 (N_2804,In_1156,In_1974);
xnor U2805 (N_2805,In_1107,In_528);
xor U2806 (N_2806,In_14,In_2);
nor U2807 (N_2807,In_526,In_903);
nor U2808 (N_2808,In_1008,In_1618);
nand U2809 (N_2809,In_596,In_113);
nand U2810 (N_2810,In_2055,In_2556);
or U2811 (N_2811,In_1924,In_2907);
xor U2812 (N_2812,In_788,In_1531);
xnor U2813 (N_2813,In_374,In_1510);
nand U2814 (N_2814,In_1965,In_2710);
or U2815 (N_2815,In_1326,In_1607);
and U2816 (N_2816,In_1649,In_1925);
xnor U2817 (N_2817,In_1771,In_1903);
xnor U2818 (N_2818,In_977,In_2423);
nor U2819 (N_2819,In_438,In_668);
or U2820 (N_2820,In_541,In_2573);
nand U2821 (N_2821,In_1324,In_859);
and U2822 (N_2822,In_2179,In_1924);
nand U2823 (N_2823,In_1397,In_1017);
nor U2824 (N_2824,In_604,In_2219);
nor U2825 (N_2825,In_950,In_607);
nand U2826 (N_2826,In_1395,In_1022);
nor U2827 (N_2827,In_2586,In_1460);
nor U2828 (N_2828,In_1111,In_2245);
nand U2829 (N_2829,In_228,In_1164);
xor U2830 (N_2830,In_1591,In_1159);
and U2831 (N_2831,In_1577,In_1812);
and U2832 (N_2832,In_1360,In_2202);
nor U2833 (N_2833,In_1246,In_2453);
or U2834 (N_2834,In_1406,In_1955);
and U2835 (N_2835,In_154,In_2149);
and U2836 (N_2836,In_181,In_1339);
and U2837 (N_2837,In_196,In_1276);
xor U2838 (N_2838,In_1342,In_811);
nand U2839 (N_2839,In_874,In_1991);
xnor U2840 (N_2840,In_1636,In_385);
nand U2841 (N_2841,In_2549,In_2107);
and U2842 (N_2842,In_993,In_2473);
and U2843 (N_2843,In_923,In_520);
nor U2844 (N_2844,In_1862,In_1302);
and U2845 (N_2845,In_2257,In_2080);
and U2846 (N_2846,In_306,In_2081);
nor U2847 (N_2847,In_2361,In_514);
xor U2848 (N_2848,In_2073,In_602);
xor U2849 (N_2849,In_262,In_257);
and U2850 (N_2850,In_2132,In_1695);
or U2851 (N_2851,In_2874,In_682);
and U2852 (N_2852,In_2556,In_2977);
xor U2853 (N_2853,In_1703,In_1651);
or U2854 (N_2854,In_1904,In_2257);
nand U2855 (N_2855,In_1404,In_2739);
or U2856 (N_2856,In_1210,In_2377);
or U2857 (N_2857,In_2060,In_2341);
nand U2858 (N_2858,In_2290,In_2373);
and U2859 (N_2859,In_1591,In_2861);
xnor U2860 (N_2860,In_2783,In_1637);
nor U2861 (N_2861,In_2249,In_2862);
xnor U2862 (N_2862,In_2803,In_2365);
nor U2863 (N_2863,In_602,In_1419);
or U2864 (N_2864,In_1546,In_1071);
xnor U2865 (N_2865,In_459,In_1974);
and U2866 (N_2866,In_2156,In_203);
nand U2867 (N_2867,In_93,In_2953);
nor U2868 (N_2868,In_2575,In_77);
nor U2869 (N_2869,In_2347,In_2965);
xor U2870 (N_2870,In_1549,In_196);
and U2871 (N_2871,In_2013,In_1970);
xor U2872 (N_2872,In_914,In_2843);
and U2873 (N_2873,In_2838,In_624);
xor U2874 (N_2874,In_2077,In_1511);
nor U2875 (N_2875,In_2474,In_2711);
or U2876 (N_2876,In_2235,In_1864);
or U2877 (N_2877,In_325,In_992);
nand U2878 (N_2878,In_1607,In_2276);
or U2879 (N_2879,In_1276,In_468);
nand U2880 (N_2880,In_2515,In_2330);
nand U2881 (N_2881,In_2214,In_1571);
nand U2882 (N_2882,In_1192,In_2226);
xor U2883 (N_2883,In_1850,In_726);
or U2884 (N_2884,In_722,In_1277);
or U2885 (N_2885,In_401,In_1676);
and U2886 (N_2886,In_2761,In_1035);
and U2887 (N_2887,In_308,In_244);
or U2888 (N_2888,In_1232,In_2024);
nor U2889 (N_2889,In_2398,In_309);
nor U2890 (N_2890,In_2152,In_2520);
and U2891 (N_2891,In_246,In_303);
nor U2892 (N_2892,In_1313,In_643);
or U2893 (N_2893,In_1853,In_960);
xnor U2894 (N_2894,In_1049,In_72);
xnor U2895 (N_2895,In_885,In_2105);
xor U2896 (N_2896,In_468,In_871);
nor U2897 (N_2897,In_552,In_2613);
or U2898 (N_2898,In_442,In_2604);
xor U2899 (N_2899,In_1589,In_1199);
xor U2900 (N_2900,In_906,In_1517);
and U2901 (N_2901,In_247,In_2804);
nand U2902 (N_2902,In_1940,In_2708);
and U2903 (N_2903,In_308,In_1487);
nand U2904 (N_2904,In_1903,In_1122);
and U2905 (N_2905,In_416,In_394);
xnor U2906 (N_2906,In_1246,In_276);
nand U2907 (N_2907,In_798,In_2987);
or U2908 (N_2908,In_655,In_1020);
nand U2909 (N_2909,In_77,In_671);
xor U2910 (N_2910,In_1572,In_2173);
or U2911 (N_2911,In_2982,In_1208);
or U2912 (N_2912,In_534,In_1002);
and U2913 (N_2913,In_1971,In_1801);
or U2914 (N_2914,In_2712,In_1152);
nand U2915 (N_2915,In_933,In_133);
or U2916 (N_2916,In_464,In_585);
and U2917 (N_2917,In_720,In_1582);
nor U2918 (N_2918,In_1370,In_2001);
nor U2919 (N_2919,In_787,In_2569);
or U2920 (N_2920,In_2848,In_1884);
nand U2921 (N_2921,In_2308,In_2014);
and U2922 (N_2922,In_508,In_497);
xnor U2923 (N_2923,In_769,In_2739);
nand U2924 (N_2924,In_2779,In_2072);
nor U2925 (N_2925,In_1280,In_2749);
and U2926 (N_2926,In_1002,In_953);
nand U2927 (N_2927,In_261,In_248);
xnor U2928 (N_2928,In_319,In_985);
nand U2929 (N_2929,In_2551,In_59);
nor U2930 (N_2930,In_2749,In_1303);
or U2931 (N_2931,In_2171,In_1096);
xor U2932 (N_2932,In_2075,In_2295);
or U2933 (N_2933,In_2070,In_778);
xnor U2934 (N_2934,In_1679,In_5);
nor U2935 (N_2935,In_936,In_1544);
nand U2936 (N_2936,In_2227,In_624);
and U2937 (N_2937,In_1456,In_495);
xor U2938 (N_2938,In_26,In_332);
nor U2939 (N_2939,In_1750,In_381);
or U2940 (N_2940,In_827,In_2592);
and U2941 (N_2941,In_2037,In_2463);
xnor U2942 (N_2942,In_2694,In_20);
nor U2943 (N_2943,In_2865,In_1823);
or U2944 (N_2944,In_1793,In_2693);
or U2945 (N_2945,In_2260,In_2104);
nand U2946 (N_2946,In_1803,In_2379);
xnor U2947 (N_2947,In_511,In_411);
nand U2948 (N_2948,In_295,In_1202);
xnor U2949 (N_2949,In_516,In_414);
or U2950 (N_2950,In_2761,In_2469);
xnor U2951 (N_2951,In_2611,In_1500);
nor U2952 (N_2952,In_1449,In_433);
nor U2953 (N_2953,In_2804,In_159);
or U2954 (N_2954,In_931,In_1046);
nand U2955 (N_2955,In_1312,In_1856);
nand U2956 (N_2956,In_2075,In_2024);
nand U2957 (N_2957,In_1150,In_2516);
nand U2958 (N_2958,In_366,In_1435);
nand U2959 (N_2959,In_2197,In_2);
or U2960 (N_2960,In_2269,In_165);
nor U2961 (N_2961,In_942,In_2300);
or U2962 (N_2962,In_150,In_2712);
nand U2963 (N_2963,In_1831,In_1321);
nand U2964 (N_2964,In_465,In_2734);
nand U2965 (N_2965,In_1583,In_2608);
nor U2966 (N_2966,In_1081,In_1766);
nor U2967 (N_2967,In_2149,In_885);
nor U2968 (N_2968,In_198,In_1118);
nand U2969 (N_2969,In_1331,In_1770);
xor U2970 (N_2970,In_2445,In_866);
or U2971 (N_2971,In_1774,In_986);
and U2972 (N_2972,In_9,In_929);
and U2973 (N_2973,In_1379,In_680);
nand U2974 (N_2974,In_2033,In_967);
and U2975 (N_2975,In_816,In_2077);
nor U2976 (N_2976,In_183,In_1318);
or U2977 (N_2977,In_332,In_367);
or U2978 (N_2978,In_417,In_2051);
and U2979 (N_2979,In_2466,In_2287);
nor U2980 (N_2980,In_1261,In_554);
nor U2981 (N_2981,In_1168,In_1860);
nand U2982 (N_2982,In_1670,In_1758);
or U2983 (N_2983,In_1159,In_258);
nand U2984 (N_2984,In_781,In_1578);
and U2985 (N_2985,In_1853,In_1635);
nand U2986 (N_2986,In_2922,In_2650);
nand U2987 (N_2987,In_1253,In_365);
and U2988 (N_2988,In_1082,In_1744);
nor U2989 (N_2989,In_2302,In_862);
nor U2990 (N_2990,In_1311,In_1042);
or U2991 (N_2991,In_2533,In_909);
xor U2992 (N_2992,In_752,In_1945);
and U2993 (N_2993,In_2294,In_2787);
or U2994 (N_2994,In_2759,In_2673);
and U2995 (N_2995,In_1120,In_1225);
or U2996 (N_2996,In_2236,In_2816);
xnor U2997 (N_2997,In_517,In_1217);
xnor U2998 (N_2998,In_923,In_767);
and U2999 (N_2999,In_477,In_733);
xor U3000 (N_3000,In_1215,In_1657);
xnor U3001 (N_3001,In_2245,In_1185);
nor U3002 (N_3002,In_499,In_2401);
xnor U3003 (N_3003,In_580,In_1670);
or U3004 (N_3004,In_2215,In_465);
nand U3005 (N_3005,In_2476,In_611);
nor U3006 (N_3006,In_405,In_1892);
xor U3007 (N_3007,In_1254,In_2267);
and U3008 (N_3008,In_736,In_2983);
xor U3009 (N_3009,In_2791,In_1653);
nor U3010 (N_3010,In_2370,In_149);
nand U3011 (N_3011,In_331,In_1736);
nor U3012 (N_3012,In_1803,In_2832);
nand U3013 (N_3013,In_1666,In_692);
and U3014 (N_3014,In_626,In_1650);
nor U3015 (N_3015,In_1320,In_2855);
xnor U3016 (N_3016,In_1943,In_348);
or U3017 (N_3017,In_2566,In_612);
nand U3018 (N_3018,In_1714,In_1652);
nor U3019 (N_3019,In_1647,In_2838);
nor U3020 (N_3020,In_2599,In_1477);
nand U3021 (N_3021,In_1620,In_1603);
and U3022 (N_3022,In_2275,In_1946);
and U3023 (N_3023,In_1111,In_716);
and U3024 (N_3024,In_2483,In_1201);
and U3025 (N_3025,In_1569,In_1738);
or U3026 (N_3026,In_642,In_1460);
and U3027 (N_3027,In_276,In_661);
and U3028 (N_3028,In_202,In_745);
nor U3029 (N_3029,In_1069,In_93);
nor U3030 (N_3030,In_1123,In_1395);
or U3031 (N_3031,In_1563,In_2831);
and U3032 (N_3032,In_2742,In_634);
xnor U3033 (N_3033,In_70,In_2863);
nor U3034 (N_3034,In_285,In_1425);
xor U3035 (N_3035,In_989,In_482);
or U3036 (N_3036,In_159,In_2967);
nor U3037 (N_3037,In_151,In_2432);
xor U3038 (N_3038,In_1232,In_807);
nor U3039 (N_3039,In_915,In_936);
and U3040 (N_3040,In_354,In_2719);
nand U3041 (N_3041,In_2841,In_1493);
nand U3042 (N_3042,In_1346,In_158);
nand U3043 (N_3043,In_238,In_2532);
nor U3044 (N_3044,In_356,In_2931);
xor U3045 (N_3045,In_655,In_679);
nand U3046 (N_3046,In_2390,In_1540);
or U3047 (N_3047,In_2560,In_2820);
nor U3048 (N_3048,In_1270,In_302);
nand U3049 (N_3049,In_1434,In_250);
nor U3050 (N_3050,In_2941,In_2640);
xor U3051 (N_3051,In_757,In_740);
and U3052 (N_3052,In_1666,In_2544);
nand U3053 (N_3053,In_1414,In_2536);
nor U3054 (N_3054,In_1168,In_2226);
nor U3055 (N_3055,In_2600,In_2283);
or U3056 (N_3056,In_2440,In_2613);
and U3057 (N_3057,In_2336,In_1335);
nand U3058 (N_3058,In_1240,In_909);
nand U3059 (N_3059,In_1543,In_943);
or U3060 (N_3060,In_465,In_487);
nor U3061 (N_3061,In_499,In_2442);
or U3062 (N_3062,In_2669,In_931);
and U3063 (N_3063,In_557,In_2764);
and U3064 (N_3064,In_916,In_176);
nor U3065 (N_3065,In_2,In_2534);
or U3066 (N_3066,In_2228,In_2999);
nand U3067 (N_3067,In_2648,In_83);
xnor U3068 (N_3068,In_1845,In_149);
nor U3069 (N_3069,In_2575,In_2042);
nand U3070 (N_3070,In_896,In_2229);
nand U3071 (N_3071,In_2502,In_2556);
or U3072 (N_3072,In_1871,In_1149);
and U3073 (N_3073,In_709,In_1680);
nand U3074 (N_3074,In_398,In_837);
nand U3075 (N_3075,In_67,In_1258);
nand U3076 (N_3076,In_1671,In_2177);
and U3077 (N_3077,In_2748,In_226);
and U3078 (N_3078,In_1381,In_2508);
xor U3079 (N_3079,In_1083,In_1118);
nand U3080 (N_3080,In_284,In_2353);
nand U3081 (N_3081,In_566,In_2436);
nor U3082 (N_3082,In_2024,In_1892);
and U3083 (N_3083,In_2638,In_2476);
xor U3084 (N_3084,In_2955,In_1022);
nand U3085 (N_3085,In_383,In_2948);
nor U3086 (N_3086,In_315,In_763);
nor U3087 (N_3087,In_2380,In_2901);
nor U3088 (N_3088,In_2097,In_1863);
and U3089 (N_3089,In_1899,In_2959);
xor U3090 (N_3090,In_281,In_2333);
or U3091 (N_3091,In_840,In_483);
nand U3092 (N_3092,In_788,In_2325);
and U3093 (N_3093,In_2146,In_1264);
nor U3094 (N_3094,In_937,In_1404);
nor U3095 (N_3095,In_287,In_480);
nand U3096 (N_3096,In_1624,In_1041);
nand U3097 (N_3097,In_728,In_54);
nor U3098 (N_3098,In_2245,In_593);
xor U3099 (N_3099,In_687,In_1940);
nand U3100 (N_3100,In_1998,In_2042);
nor U3101 (N_3101,In_613,In_627);
nor U3102 (N_3102,In_1145,In_991);
or U3103 (N_3103,In_2838,In_1088);
and U3104 (N_3104,In_1407,In_2231);
nand U3105 (N_3105,In_598,In_1610);
and U3106 (N_3106,In_2905,In_380);
xnor U3107 (N_3107,In_2580,In_2253);
xnor U3108 (N_3108,In_267,In_602);
nor U3109 (N_3109,In_1760,In_2907);
nand U3110 (N_3110,In_2666,In_95);
nor U3111 (N_3111,In_2703,In_2862);
xnor U3112 (N_3112,In_2107,In_632);
or U3113 (N_3113,In_1719,In_523);
and U3114 (N_3114,In_1655,In_44);
nand U3115 (N_3115,In_2337,In_2370);
xnor U3116 (N_3116,In_1223,In_673);
xor U3117 (N_3117,In_146,In_9);
and U3118 (N_3118,In_2322,In_1217);
or U3119 (N_3119,In_2775,In_1928);
and U3120 (N_3120,In_1225,In_132);
or U3121 (N_3121,In_2683,In_2903);
nand U3122 (N_3122,In_2636,In_90);
nor U3123 (N_3123,In_516,In_284);
nor U3124 (N_3124,In_985,In_29);
nor U3125 (N_3125,In_2467,In_1401);
nand U3126 (N_3126,In_607,In_1729);
or U3127 (N_3127,In_1717,In_585);
nor U3128 (N_3128,In_2759,In_1270);
or U3129 (N_3129,In_1735,In_609);
or U3130 (N_3130,In_2306,In_2076);
or U3131 (N_3131,In_463,In_2019);
nor U3132 (N_3132,In_2271,In_2800);
and U3133 (N_3133,In_800,In_248);
nor U3134 (N_3134,In_676,In_1311);
and U3135 (N_3135,In_987,In_1067);
xor U3136 (N_3136,In_2390,In_1680);
nand U3137 (N_3137,In_772,In_1968);
nand U3138 (N_3138,In_961,In_2370);
xnor U3139 (N_3139,In_332,In_737);
nand U3140 (N_3140,In_26,In_528);
and U3141 (N_3141,In_657,In_1971);
xor U3142 (N_3142,In_2364,In_1531);
nor U3143 (N_3143,In_1413,In_1775);
or U3144 (N_3144,In_2081,In_2263);
nand U3145 (N_3145,In_379,In_699);
nand U3146 (N_3146,In_318,In_756);
or U3147 (N_3147,In_24,In_1498);
nor U3148 (N_3148,In_446,In_1935);
and U3149 (N_3149,In_288,In_987);
and U3150 (N_3150,In_1269,In_591);
nand U3151 (N_3151,In_264,In_392);
nand U3152 (N_3152,In_1774,In_314);
nand U3153 (N_3153,In_1304,In_2086);
nand U3154 (N_3154,In_1449,In_1531);
nand U3155 (N_3155,In_838,In_2888);
nand U3156 (N_3156,In_1036,In_718);
nand U3157 (N_3157,In_125,In_1007);
and U3158 (N_3158,In_73,In_1402);
nand U3159 (N_3159,In_1300,In_2648);
or U3160 (N_3160,In_1790,In_304);
nand U3161 (N_3161,In_2804,In_1928);
xnor U3162 (N_3162,In_1263,In_2769);
nand U3163 (N_3163,In_1461,In_1227);
or U3164 (N_3164,In_930,In_388);
nand U3165 (N_3165,In_1698,In_1659);
nand U3166 (N_3166,In_2087,In_1443);
or U3167 (N_3167,In_2023,In_1155);
nand U3168 (N_3168,In_102,In_1590);
xnor U3169 (N_3169,In_2427,In_531);
or U3170 (N_3170,In_1507,In_2530);
xnor U3171 (N_3171,In_1900,In_1569);
and U3172 (N_3172,In_116,In_660);
nor U3173 (N_3173,In_2259,In_1797);
xor U3174 (N_3174,In_2959,In_1501);
nand U3175 (N_3175,In_1558,In_840);
nand U3176 (N_3176,In_143,In_427);
xor U3177 (N_3177,In_842,In_1414);
nand U3178 (N_3178,In_2816,In_827);
and U3179 (N_3179,In_1873,In_1372);
and U3180 (N_3180,In_1430,In_2789);
and U3181 (N_3181,In_1534,In_2607);
nand U3182 (N_3182,In_579,In_100);
nand U3183 (N_3183,In_12,In_313);
nand U3184 (N_3184,In_2692,In_1531);
and U3185 (N_3185,In_1870,In_1183);
xor U3186 (N_3186,In_2481,In_2026);
xor U3187 (N_3187,In_1589,In_2161);
and U3188 (N_3188,In_2551,In_2783);
nor U3189 (N_3189,In_2674,In_1746);
xor U3190 (N_3190,In_2719,In_407);
or U3191 (N_3191,In_548,In_756);
xnor U3192 (N_3192,In_1402,In_2994);
or U3193 (N_3193,In_124,In_2058);
xnor U3194 (N_3194,In_2441,In_1324);
nor U3195 (N_3195,In_2431,In_711);
nand U3196 (N_3196,In_2482,In_1637);
nor U3197 (N_3197,In_247,In_1257);
and U3198 (N_3198,In_1177,In_658);
nor U3199 (N_3199,In_1505,In_2395);
xnor U3200 (N_3200,In_55,In_2919);
xor U3201 (N_3201,In_2219,In_546);
nor U3202 (N_3202,In_2236,In_2614);
nor U3203 (N_3203,In_1653,In_1418);
nor U3204 (N_3204,In_618,In_649);
xor U3205 (N_3205,In_2771,In_1481);
or U3206 (N_3206,In_2256,In_2408);
and U3207 (N_3207,In_475,In_1058);
or U3208 (N_3208,In_323,In_527);
nand U3209 (N_3209,In_2336,In_191);
nor U3210 (N_3210,In_2547,In_234);
and U3211 (N_3211,In_2163,In_2280);
xnor U3212 (N_3212,In_2693,In_1342);
nand U3213 (N_3213,In_2056,In_677);
and U3214 (N_3214,In_339,In_165);
nand U3215 (N_3215,In_37,In_14);
and U3216 (N_3216,In_574,In_751);
nand U3217 (N_3217,In_803,In_136);
xnor U3218 (N_3218,In_2374,In_2544);
xor U3219 (N_3219,In_306,In_2856);
or U3220 (N_3220,In_1174,In_1247);
and U3221 (N_3221,In_109,In_1185);
nand U3222 (N_3222,In_1088,In_347);
or U3223 (N_3223,In_2275,In_2790);
and U3224 (N_3224,In_2375,In_2616);
xnor U3225 (N_3225,In_2411,In_2708);
and U3226 (N_3226,In_1112,In_1882);
nand U3227 (N_3227,In_2082,In_2834);
and U3228 (N_3228,In_779,In_2908);
or U3229 (N_3229,In_1973,In_1680);
nand U3230 (N_3230,In_1647,In_2064);
and U3231 (N_3231,In_1416,In_1127);
nor U3232 (N_3232,In_350,In_1571);
nor U3233 (N_3233,In_2162,In_85);
or U3234 (N_3234,In_1738,In_2366);
nor U3235 (N_3235,In_2886,In_2622);
or U3236 (N_3236,In_340,In_1612);
nor U3237 (N_3237,In_1754,In_2604);
and U3238 (N_3238,In_1115,In_2436);
and U3239 (N_3239,In_1656,In_652);
xnor U3240 (N_3240,In_1857,In_636);
xnor U3241 (N_3241,In_699,In_1002);
or U3242 (N_3242,In_101,In_1220);
nor U3243 (N_3243,In_723,In_2569);
or U3244 (N_3244,In_1803,In_895);
or U3245 (N_3245,In_2633,In_2328);
nand U3246 (N_3246,In_1139,In_2040);
xnor U3247 (N_3247,In_2207,In_2433);
nor U3248 (N_3248,In_2365,In_1929);
nor U3249 (N_3249,In_2474,In_695);
or U3250 (N_3250,In_2937,In_2199);
or U3251 (N_3251,In_1127,In_1694);
or U3252 (N_3252,In_2512,In_2771);
and U3253 (N_3253,In_2818,In_621);
nand U3254 (N_3254,In_2862,In_1536);
or U3255 (N_3255,In_2,In_2905);
and U3256 (N_3256,In_2754,In_1739);
and U3257 (N_3257,In_245,In_1788);
and U3258 (N_3258,In_2130,In_508);
xor U3259 (N_3259,In_1479,In_1851);
and U3260 (N_3260,In_1866,In_2525);
xnor U3261 (N_3261,In_1944,In_558);
and U3262 (N_3262,In_2793,In_2629);
nor U3263 (N_3263,In_2690,In_2796);
xor U3264 (N_3264,In_2677,In_1634);
nor U3265 (N_3265,In_2995,In_174);
nand U3266 (N_3266,In_427,In_835);
and U3267 (N_3267,In_1636,In_2083);
or U3268 (N_3268,In_1296,In_2694);
nor U3269 (N_3269,In_1386,In_2991);
and U3270 (N_3270,In_2106,In_423);
xor U3271 (N_3271,In_1554,In_2455);
or U3272 (N_3272,In_1425,In_983);
nand U3273 (N_3273,In_1560,In_1800);
and U3274 (N_3274,In_1395,In_1750);
or U3275 (N_3275,In_1850,In_766);
nor U3276 (N_3276,In_2799,In_2535);
xor U3277 (N_3277,In_1770,In_2408);
nand U3278 (N_3278,In_626,In_2347);
and U3279 (N_3279,In_1577,In_2196);
xor U3280 (N_3280,In_1527,In_605);
xnor U3281 (N_3281,In_1290,In_1510);
or U3282 (N_3282,In_792,In_2504);
nand U3283 (N_3283,In_415,In_979);
or U3284 (N_3284,In_1789,In_542);
nand U3285 (N_3285,In_2355,In_1189);
or U3286 (N_3286,In_351,In_1000);
xor U3287 (N_3287,In_2779,In_572);
nand U3288 (N_3288,In_1514,In_2601);
or U3289 (N_3289,In_548,In_2445);
nand U3290 (N_3290,In_550,In_375);
or U3291 (N_3291,In_2954,In_2314);
or U3292 (N_3292,In_1342,In_2153);
nor U3293 (N_3293,In_1972,In_1802);
nor U3294 (N_3294,In_670,In_939);
nor U3295 (N_3295,In_1981,In_2254);
nand U3296 (N_3296,In_1646,In_2581);
nand U3297 (N_3297,In_286,In_434);
xnor U3298 (N_3298,In_2078,In_2107);
or U3299 (N_3299,In_1288,In_816);
xnor U3300 (N_3300,In_754,In_922);
or U3301 (N_3301,In_2234,In_1627);
nor U3302 (N_3302,In_2797,In_1428);
nor U3303 (N_3303,In_2066,In_421);
or U3304 (N_3304,In_357,In_1088);
nand U3305 (N_3305,In_2335,In_830);
xor U3306 (N_3306,In_1666,In_717);
xor U3307 (N_3307,In_2335,In_1042);
nor U3308 (N_3308,In_1620,In_1686);
and U3309 (N_3309,In_436,In_1784);
xnor U3310 (N_3310,In_603,In_2854);
and U3311 (N_3311,In_292,In_1935);
nor U3312 (N_3312,In_1538,In_2548);
xor U3313 (N_3313,In_1069,In_2197);
xnor U3314 (N_3314,In_799,In_2221);
nor U3315 (N_3315,In_1785,In_2740);
nand U3316 (N_3316,In_2146,In_164);
nor U3317 (N_3317,In_914,In_2471);
or U3318 (N_3318,In_2166,In_1959);
xnor U3319 (N_3319,In_2065,In_810);
nand U3320 (N_3320,In_188,In_251);
or U3321 (N_3321,In_1152,In_731);
nor U3322 (N_3322,In_960,In_442);
and U3323 (N_3323,In_2683,In_2908);
and U3324 (N_3324,In_1667,In_1257);
or U3325 (N_3325,In_1586,In_495);
nand U3326 (N_3326,In_2197,In_1218);
or U3327 (N_3327,In_2139,In_915);
nand U3328 (N_3328,In_1338,In_2280);
and U3329 (N_3329,In_677,In_2391);
xor U3330 (N_3330,In_1842,In_2271);
xor U3331 (N_3331,In_2266,In_1846);
nor U3332 (N_3332,In_1873,In_2421);
xor U3333 (N_3333,In_44,In_144);
nand U3334 (N_3334,In_2063,In_2209);
nand U3335 (N_3335,In_1546,In_2472);
and U3336 (N_3336,In_1781,In_1158);
xor U3337 (N_3337,In_731,In_2498);
nor U3338 (N_3338,In_1241,In_1181);
nor U3339 (N_3339,In_2241,In_834);
nand U3340 (N_3340,In_2419,In_383);
nor U3341 (N_3341,In_1346,In_2854);
and U3342 (N_3342,In_182,In_1796);
xor U3343 (N_3343,In_2553,In_2404);
or U3344 (N_3344,In_726,In_1954);
or U3345 (N_3345,In_1650,In_450);
nand U3346 (N_3346,In_182,In_952);
nand U3347 (N_3347,In_1546,In_2532);
nand U3348 (N_3348,In_372,In_2754);
or U3349 (N_3349,In_2337,In_1025);
nor U3350 (N_3350,In_744,In_2508);
or U3351 (N_3351,In_1086,In_1371);
nor U3352 (N_3352,In_2512,In_2218);
nor U3353 (N_3353,In_1212,In_742);
nor U3354 (N_3354,In_1556,In_1163);
nor U3355 (N_3355,In_568,In_1206);
and U3356 (N_3356,In_1827,In_1331);
or U3357 (N_3357,In_2652,In_2073);
xnor U3358 (N_3358,In_268,In_1678);
nor U3359 (N_3359,In_1341,In_29);
and U3360 (N_3360,In_1546,In_2055);
and U3361 (N_3361,In_2699,In_171);
or U3362 (N_3362,In_2687,In_2383);
nor U3363 (N_3363,In_1194,In_919);
nor U3364 (N_3364,In_56,In_2785);
or U3365 (N_3365,In_685,In_1265);
or U3366 (N_3366,In_912,In_168);
xnor U3367 (N_3367,In_1686,In_825);
xor U3368 (N_3368,In_832,In_896);
or U3369 (N_3369,In_689,In_2097);
xor U3370 (N_3370,In_2831,In_262);
xor U3371 (N_3371,In_1010,In_2850);
and U3372 (N_3372,In_1548,In_295);
nor U3373 (N_3373,In_2021,In_1679);
and U3374 (N_3374,In_619,In_1026);
and U3375 (N_3375,In_90,In_195);
or U3376 (N_3376,In_120,In_70);
nand U3377 (N_3377,In_280,In_2381);
and U3378 (N_3378,In_180,In_80);
and U3379 (N_3379,In_2106,In_2108);
and U3380 (N_3380,In_1641,In_1835);
nor U3381 (N_3381,In_1153,In_2109);
xnor U3382 (N_3382,In_1229,In_2470);
or U3383 (N_3383,In_1479,In_984);
nand U3384 (N_3384,In_2609,In_728);
or U3385 (N_3385,In_2215,In_2480);
or U3386 (N_3386,In_2095,In_1544);
nor U3387 (N_3387,In_104,In_2070);
nor U3388 (N_3388,In_896,In_730);
xor U3389 (N_3389,In_1420,In_1109);
nor U3390 (N_3390,In_2921,In_2757);
or U3391 (N_3391,In_518,In_1647);
and U3392 (N_3392,In_428,In_2239);
nor U3393 (N_3393,In_2347,In_1385);
xnor U3394 (N_3394,In_2647,In_2636);
nand U3395 (N_3395,In_185,In_1087);
xnor U3396 (N_3396,In_2289,In_116);
nand U3397 (N_3397,In_2558,In_1964);
or U3398 (N_3398,In_878,In_2853);
nand U3399 (N_3399,In_1010,In_1074);
xor U3400 (N_3400,In_867,In_180);
or U3401 (N_3401,In_982,In_983);
and U3402 (N_3402,In_426,In_778);
nor U3403 (N_3403,In_1413,In_90);
and U3404 (N_3404,In_1545,In_477);
or U3405 (N_3405,In_204,In_993);
xor U3406 (N_3406,In_1771,In_593);
or U3407 (N_3407,In_815,In_2266);
and U3408 (N_3408,In_923,In_573);
and U3409 (N_3409,In_2082,In_2860);
or U3410 (N_3410,In_258,In_1467);
or U3411 (N_3411,In_2659,In_1884);
nor U3412 (N_3412,In_1739,In_2466);
or U3413 (N_3413,In_1140,In_624);
xnor U3414 (N_3414,In_2709,In_2552);
nor U3415 (N_3415,In_2701,In_2742);
and U3416 (N_3416,In_2073,In_2035);
and U3417 (N_3417,In_837,In_2895);
and U3418 (N_3418,In_1001,In_2230);
or U3419 (N_3419,In_1266,In_187);
nand U3420 (N_3420,In_712,In_286);
xnor U3421 (N_3421,In_2032,In_762);
or U3422 (N_3422,In_256,In_1062);
nand U3423 (N_3423,In_526,In_2621);
xnor U3424 (N_3424,In_2242,In_2098);
xor U3425 (N_3425,In_963,In_1745);
nand U3426 (N_3426,In_391,In_1631);
nor U3427 (N_3427,In_363,In_1261);
or U3428 (N_3428,In_2100,In_627);
nor U3429 (N_3429,In_907,In_450);
xor U3430 (N_3430,In_1983,In_2289);
and U3431 (N_3431,In_1884,In_1779);
or U3432 (N_3432,In_1822,In_614);
nor U3433 (N_3433,In_1657,In_1621);
nor U3434 (N_3434,In_2631,In_1569);
xnor U3435 (N_3435,In_481,In_299);
xnor U3436 (N_3436,In_2562,In_1258);
xor U3437 (N_3437,In_1911,In_652);
nand U3438 (N_3438,In_1849,In_57);
nand U3439 (N_3439,In_210,In_1318);
nand U3440 (N_3440,In_2996,In_154);
or U3441 (N_3441,In_149,In_1022);
and U3442 (N_3442,In_2328,In_2784);
or U3443 (N_3443,In_43,In_890);
and U3444 (N_3444,In_1332,In_1516);
nor U3445 (N_3445,In_539,In_488);
or U3446 (N_3446,In_2143,In_594);
or U3447 (N_3447,In_176,In_864);
xor U3448 (N_3448,In_814,In_1080);
nand U3449 (N_3449,In_1667,In_1411);
nand U3450 (N_3450,In_0,In_2559);
nor U3451 (N_3451,In_1749,In_1281);
and U3452 (N_3452,In_2204,In_1082);
nand U3453 (N_3453,In_763,In_2528);
and U3454 (N_3454,In_2809,In_1097);
and U3455 (N_3455,In_716,In_150);
and U3456 (N_3456,In_1744,In_1909);
or U3457 (N_3457,In_2648,In_1953);
or U3458 (N_3458,In_2157,In_144);
nand U3459 (N_3459,In_546,In_1130);
and U3460 (N_3460,In_1662,In_2023);
and U3461 (N_3461,In_840,In_1919);
or U3462 (N_3462,In_1567,In_1958);
and U3463 (N_3463,In_2299,In_1382);
nand U3464 (N_3464,In_1455,In_115);
xnor U3465 (N_3465,In_1949,In_547);
xor U3466 (N_3466,In_1209,In_187);
nor U3467 (N_3467,In_287,In_1136);
xnor U3468 (N_3468,In_594,In_1255);
nand U3469 (N_3469,In_2000,In_1929);
xnor U3470 (N_3470,In_294,In_1848);
or U3471 (N_3471,In_1757,In_475);
and U3472 (N_3472,In_1452,In_1237);
or U3473 (N_3473,In_59,In_125);
nand U3474 (N_3474,In_2010,In_702);
nand U3475 (N_3475,In_1509,In_761);
nor U3476 (N_3476,In_844,In_584);
or U3477 (N_3477,In_1960,In_1208);
or U3478 (N_3478,In_2179,In_594);
and U3479 (N_3479,In_2592,In_2073);
and U3480 (N_3480,In_2923,In_156);
nor U3481 (N_3481,In_593,In_1170);
and U3482 (N_3482,In_1455,In_2625);
xnor U3483 (N_3483,In_743,In_2477);
xor U3484 (N_3484,In_1255,In_642);
xor U3485 (N_3485,In_515,In_1264);
nor U3486 (N_3486,In_1322,In_1705);
xnor U3487 (N_3487,In_99,In_564);
xor U3488 (N_3488,In_2160,In_353);
or U3489 (N_3489,In_2551,In_1966);
and U3490 (N_3490,In_1721,In_2221);
nor U3491 (N_3491,In_2630,In_699);
and U3492 (N_3492,In_242,In_1844);
nor U3493 (N_3493,In_1,In_1828);
and U3494 (N_3494,In_448,In_2985);
nand U3495 (N_3495,In_1707,In_2959);
nor U3496 (N_3496,In_1178,In_2070);
nor U3497 (N_3497,In_927,In_59);
and U3498 (N_3498,In_365,In_645);
nand U3499 (N_3499,In_1789,In_2372);
or U3500 (N_3500,In_1172,In_1375);
nand U3501 (N_3501,In_2889,In_526);
and U3502 (N_3502,In_254,In_222);
nor U3503 (N_3503,In_2335,In_104);
or U3504 (N_3504,In_720,In_206);
and U3505 (N_3505,In_196,In_2648);
and U3506 (N_3506,In_2899,In_2913);
and U3507 (N_3507,In_2061,In_255);
or U3508 (N_3508,In_757,In_592);
and U3509 (N_3509,In_1790,In_2316);
nand U3510 (N_3510,In_1318,In_184);
nor U3511 (N_3511,In_3,In_2658);
and U3512 (N_3512,In_955,In_946);
nand U3513 (N_3513,In_2614,In_2515);
xnor U3514 (N_3514,In_1489,In_908);
xor U3515 (N_3515,In_2363,In_2146);
nor U3516 (N_3516,In_94,In_2354);
or U3517 (N_3517,In_2673,In_267);
nand U3518 (N_3518,In_404,In_1259);
xor U3519 (N_3519,In_935,In_2727);
nand U3520 (N_3520,In_983,In_28);
xnor U3521 (N_3521,In_676,In_1052);
or U3522 (N_3522,In_2398,In_1154);
nand U3523 (N_3523,In_2335,In_1922);
and U3524 (N_3524,In_1041,In_43);
or U3525 (N_3525,In_2693,In_1301);
xor U3526 (N_3526,In_2923,In_1228);
or U3527 (N_3527,In_1119,In_576);
nor U3528 (N_3528,In_1233,In_1996);
nand U3529 (N_3529,In_1606,In_1288);
nand U3530 (N_3530,In_1486,In_280);
nor U3531 (N_3531,In_1195,In_2772);
or U3532 (N_3532,In_2522,In_1378);
and U3533 (N_3533,In_1561,In_2739);
and U3534 (N_3534,In_52,In_1468);
and U3535 (N_3535,In_392,In_288);
and U3536 (N_3536,In_1607,In_1463);
and U3537 (N_3537,In_970,In_2130);
and U3538 (N_3538,In_1496,In_1087);
or U3539 (N_3539,In_1298,In_1474);
nand U3540 (N_3540,In_1373,In_908);
nor U3541 (N_3541,In_934,In_140);
xor U3542 (N_3542,In_1212,In_2459);
and U3543 (N_3543,In_956,In_442);
nand U3544 (N_3544,In_1802,In_1808);
xor U3545 (N_3545,In_776,In_1391);
or U3546 (N_3546,In_2521,In_1068);
xor U3547 (N_3547,In_1960,In_1762);
nand U3548 (N_3548,In_930,In_782);
and U3549 (N_3549,In_1796,In_224);
xor U3550 (N_3550,In_252,In_2758);
xor U3551 (N_3551,In_237,In_1086);
and U3552 (N_3552,In_2749,In_2155);
xnor U3553 (N_3553,In_2149,In_906);
nand U3554 (N_3554,In_1171,In_1250);
or U3555 (N_3555,In_229,In_1493);
and U3556 (N_3556,In_1843,In_2019);
xor U3557 (N_3557,In_1730,In_346);
xor U3558 (N_3558,In_2081,In_2524);
nor U3559 (N_3559,In_2831,In_1974);
xnor U3560 (N_3560,In_460,In_825);
xnor U3561 (N_3561,In_6,In_2197);
and U3562 (N_3562,In_1520,In_729);
nor U3563 (N_3563,In_969,In_1829);
nor U3564 (N_3564,In_160,In_928);
nor U3565 (N_3565,In_1592,In_1377);
nand U3566 (N_3566,In_512,In_1436);
nand U3567 (N_3567,In_492,In_1861);
and U3568 (N_3568,In_2836,In_1664);
nand U3569 (N_3569,In_1397,In_2605);
xor U3570 (N_3570,In_752,In_1330);
or U3571 (N_3571,In_25,In_1570);
and U3572 (N_3572,In_2660,In_802);
nor U3573 (N_3573,In_1975,In_678);
xor U3574 (N_3574,In_598,In_1042);
and U3575 (N_3575,In_152,In_1151);
nand U3576 (N_3576,In_1177,In_1180);
nor U3577 (N_3577,In_2637,In_223);
or U3578 (N_3578,In_2051,In_1655);
nor U3579 (N_3579,In_2294,In_138);
nor U3580 (N_3580,In_2937,In_1492);
xor U3581 (N_3581,In_2719,In_250);
nand U3582 (N_3582,In_1551,In_1657);
nand U3583 (N_3583,In_1269,In_2883);
nand U3584 (N_3584,In_1654,In_2500);
nor U3585 (N_3585,In_2007,In_1523);
nor U3586 (N_3586,In_1564,In_238);
xor U3587 (N_3587,In_404,In_385);
nand U3588 (N_3588,In_2528,In_43);
xnor U3589 (N_3589,In_1835,In_756);
or U3590 (N_3590,In_37,In_1810);
or U3591 (N_3591,In_1910,In_615);
nor U3592 (N_3592,In_2530,In_2988);
or U3593 (N_3593,In_2341,In_1637);
and U3594 (N_3594,In_2660,In_1678);
nand U3595 (N_3595,In_2682,In_1306);
nand U3596 (N_3596,In_71,In_2098);
or U3597 (N_3597,In_2827,In_1335);
nor U3598 (N_3598,In_565,In_1034);
nor U3599 (N_3599,In_1051,In_1303);
and U3600 (N_3600,In_2481,In_177);
and U3601 (N_3601,In_1365,In_2488);
xnor U3602 (N_3602,In_2611,In_2426);
and U3603 (N_3603,In_682,In_1271);
nand U3604 (N_3604,In_1103,In_379);
or U3605 (N_3605,In_1627,In_2484);
xnor U3606 (N_3606,In_233,In_2287);
xnor U3607 (N_3607,In_990,In_254);
and U3608 (N_3608,In_1891,In_2488);
xnor U3609 (N_3609,In_1644,In_34);
and U3610 (N_3610,In_2061,In_66);
nand U3611 (N_3611,In_725,In_788);
xor U3612 (N_3612,In_1868,In_1004);
xnor U3613 (N_3613,In_953,In_1076);
nor U3614 (N_3614,In_351,In_2626);
xor U3615 (N_3615,In_2507,In_1664);
nand U3616 (N_3616,In_1820,In_975);
nor U3617 (N_3617,In_905,In_594);
nand U3618 (N_3618,In_304,In_835);
xnor U3619 (N_3619,In_1909,In_1004);
nand U3620 (N_3620,In_1236,In_1448);
and U3621 (N_3621,In_141,In_1829);
xor U3622 (N_3622,In_1697,In_49);
nor U3623 (N_3623,In_202,In_364);
xor U3624 (N_3624,In_2997,In_103);
nor U3625 (N_3625,In_2635,In_87);
xor U3626 (N_3626,In_349,In_1217);
or U3627 (N_3627,In_241,In_274);
or U3628 (N_3628,In_1215,In_638);
nand U3629 (N_3629,In_31,In_2038);
nand U3630 (N_3630,In_2644,In_1248);
or U3631 (N_3631,In_2379,In_1262);
nand U3632 (N_3632,In_2983,In_1802);
nand U3633 (N_3633,In_1105,In_1625);
and U3634 (N_3634,In_75,In_2308);
xnor U3635 (N_3635,In_2973,In_663);
or U3636 (N_3636,In_513,In_666);
nor U3637 (N_3637,In_1929,In_473);
or U3638 (N_3638,In_292,In_2705);
or U3639 (N_3639,In_1492,In_2058);
nand U3640 (N_3640,In_1059,In_2096);
xnor U3641 (N_3641,In_377,In_2156);
nand U3642 (N_3642,In_1866,In_1508);
or U3643 (N_3643,In_2950,In_2697);
xnor U3644 (N_3644,In_183,In_2292);
and U3645 (N_3645,In_1391,In_1011);
nand U3646 (N_3646,In_2306,In_2393);
or U3647 (N_3647,In_2582,In_1023);
xnor U3648 (N_3648,In_1060,In_891);
xnor U3649 (N_3649,In_1777,In_526);
and U3650 (N_3650,In_1166,In_306);
nor U3651 (N_3651,In_641,In_622);
xnor U3652 (N_3652,In_1347,In_2406);
and U3653 (N_3653,In_1015,In_2358);
xor U3654 (N_3654,In_2679,In_348);
and U3655 (N_3655,In_259,In_2617);
or U3656 (N_3656,In_2334,In_938);
nand U3657 (N_3657,In_322,In_222);
nand U3658 (N_3658,In_1144,In_1522);
nand U3659 (N_3659,In_488,In_2710);
or U3660 (N_3660,In_449,In_1724);
xnor U3661 (N_3661,In_2684,In_2736);
and U3662 (N_3662,In_2397,In_1661);
xor U3663 (N_3663,In_2979,In_2796);
xor U3664 (N_3664,In_1114,In_2983);
or U3665 (N_3665,In_1151,In_590);
and U3666 (N_3666,In_121,In_1369);
or U3667 (N_3667,In_459,In_559);
xnor U3668 (N_3668,In_367,In_295);
nor U3669 (N_3669,In_1272,In_2622);
or U3670 (N_3670,In_1759,In_1164);
xor U3671 (N_3671,In_1792,In_402);
nor U3672 (N_3672,In_641,In_2282);
nand U3673 (N_3673,In_2044,In_2088);
nor U3674 (N_3674,In_178,In_524);
xnor U3675 (N_3675,In_2600,In_234);
and U3676 (N_3676,In_235,In_2250);
xor U3677 (N_3677,In_1970,In_2306);
and U3678 (N_3678,In_2263,In_226);
nor U3679 (N_3679,In_829,In_399);
and U3680 (N_3680,In_2564,In_1305);
or U3681 (N_3681,In_263,In_1332);
xnor U3682 (N_3682,In_494,In_1521);
xnor U3683 (N_3683,In_1472,In_2648);
nand U3684 (N_3684,In_437,In_2593);
nor U3685 (N_3685,In_1223,In_2419);
nor U3686 (N_3686,In_1958,In_2519);
nor U3687 (N_3687,In_2581,In_522);
nor U3688 (N_3688,In_769,In_245);
xnor U3689 (N_3689,In_1530,In_2360);
or U3690 (N_3690,In_608,In_1870);
or U3691 (N_3691,In_524,In_951);
xnor U3692 (N_3692,In_2701,In_2760);
xnor U3693 (N_3693,In_1710,In_51);
and U3694 (N_3694,In_559,In_1836);
nand U3695 (N_3695,In_540,In_1865);
nor U3696 (N_3696,In_2290,In_954);
nand U3697 (N_3697,In_1607,In_187);
xnor U3698 (N_3698,In_911,In_2287);
nor U3699 (N_3699,In_2557,In_1418);
xnor U3700 (N_3700,In_2059,In_1400);
nand U3701 (N_3701,In_2932,In_1754);
and U3702 (N_3702,In_1195,In_541);
nand U3703 (N_3703,In_2595,In_1782);
nor U3704 (N_3704,In_2607,In_460);
xor U3705 (N_3705,In_974,In_1394);
or U3706 (N_3706,In_1544,In_614);
or U3707 (N_3707,In_1734,In_940);
xor U3708 (N_3708,In_996,In_5);
nor U3709 (N_3709,In_1661,In_124);
xor U3710 (N_3710,In_1787,In_1115);
nor U3711 (N_3711,In_2851,In_30);
xnor U3712 (N_3712,In_2614,In_2995);
and U3713 (N_3713,In_362,In_2143);
nand U3714 (N_3714,In_1097,In_1033);
or U3715 (N_3715,In_1487,In_1704);
nor U3716 (N_3716,In_1859,In_2738);
and U3717 (N_3717,In_982,In_1744);
xor U3718 (N_3718,In_1784,In_646);
nor U3719 (N_3719,In_2633,In_666);
nor U3720 (N_3720,In_2184,In_745);
xnor U3721 (N_3721,In_623,In_1919);
or U3722 (N_3722,In_1670,In_2815);
xor U3723 (N_3723,In_39,In_2781);
nand U3724 (N_3724,In_674,In_1285);
xnor U3725 (N_3725,In_405,In_1199);
or U3726 (N_3726,In_2508,In_1557);
nand U3727 (N_3727,In_2739,In_520);
xor U3728 (N_3728,In_2465,In_1803);
xnor U3729 (N_3729,In_12,In_1938);
or U3730 (N_3730,In_722,In_743);
or U3731 (N_3731,In_601,In_2857);
and U3732 (N_3732,In_1106,In_2965);
or U3733 (N_3733,In_2305,In_1427);
nor U3734 (N_3734,In_930,In_1817);
nand U3735 (N_3735,In_2060,In_2155);
or U3736 (N_3736,In_2246,In_671);
or U3737 (N_3737,In_239,In_877);
and U3738 (N_3738,In_385,In_2389);
nor U3739 (N_3739,In_1400,In_486);
nand U3740 (N_3740,In_1907,In_116);
xnor U3741 (N_3741,In_1226,In_562);
nand U3742 (N_3742,In_636,In_1672);
or U3743 (N_3743,In_868,In_1214);
nand U3744 (N_3744,In_2403,In_2398);
and U3745 (N_3745,In_63,In_419);
nand U3746 (N_3746,In_700,In_568);
or U3747 (N_3747,In_1108,In_38);
and U3748 (N_3748,In_909,In_266);
xnor U3749 (N_3749,In_1436,In_68);
nand U3750 (N_3750,In_378,In_506);
and U3751 (N_3751,In_1852,In_1686);
and U3752 (N_3752,In_1413,In_2356);
xor U3753 (N_3753,In_2453,In_1938);
nand U3754 (N_3754,In_89,In_2693);
nor U3755 (N_3755,In_744,In_2123);
nand U3756 (N_3756,In_257,In_187);
nand U3757 (N_3757,In_2277,In_2872);
or U3758 (N_3758,In_2986,In_1185);
nor U3759 (N_3759,In_1589,In_2805);
or U3760 (N_3760,In_430,In_110);
or U3761 (N_3761,In_1791,In_1625);
and U3762 (N_3762,In_2186,In_2726);
nand U3763 (N_3763,In_119,In_667);
xor U3764 (N_3764,In_614,In_554);
or U3765 (N_3765,In_2579,In_1130);
or U3766 (N_3766,In_2923,In_2548);
and U3767 (N_3767,In_1880,In_2580);
xnor U3768 (N_3768,In_1845,In_927);
nor U3769 (N_3769,In_2144,In_1412);
xnor U3770 (N_3770,In_217,In_2890);
and U3771 (N_3771,In_1096,In_2033);
or U3772 (N_3772,In_1866,In_1016);
nand U3773 (N_3773,In_2380,In_2829);
xnor U3774 (N_3774,In_2658,In_242);
nor U3775 (N_3775,In_1989,In_257);
or U3776 (N_3776,In_1448,In_427);
and U3777 (N_3777,In_893,In_511);
nand U3778 (N_3778,In_2732,In_2893);
or U3779 (N_3779,In_680,In_608);
nand U3780 (N_3780,In_341,In_618);
nand U3781 (N_3781,In_709,In_2714);
nor U3782 (N_3782,In_1759,In_2882);
nand U3783 (N_3783,In_1371,In_1094);
xnor U3784 (N_3784,In_569,In_822);
xor U3785 (N_3785,In_508,In_2403);
and U3786 (N_3786,In_1187,In_560);
xnor U3787 (N_3787,In_1762,In_1828);
and U3788 (N_3788,In_2039,In_358);
xnor U3789 (N_3789,In_2119,In_2546);
nor U3790 (N_3790,In_1123,In_1915);
nand U3791 (N_3791,In_2076,In_1309);
nor U3792 (N_3792,In_1306,In_2376);
or U3793 (N_3793,In_166,In_509);
nand U3794 (N_3794,In_2527,In_2891);
xor U3795 (N_3795,In_2085,In_166);
xnor U3796 (N_3796,In_613,In_1849);
or U3797 (N_3797,In_99,In_221);
or U3798 (N_3798,In_2282,In_361);
or U3799 (N_3799,In_1334,In_1970);
nand U3800 (N_3800,In_2226,In_1103);
nor U3801 (N_3801,In_1118,In_311);
nand U3802 (N_3802,In_2625,In_761);
nor U3803 (N_3803,In_874,In_1470);
nor U3804 (N_3804,In_1307,In_2849);
xor U3805 (N_3805,In_2777,In_1908);
nor U3806 (N_3806,In_2500,In_2581);
nand U3807 (N_3807,In_2526,In_2224);
xor U3808 (N_3808,In_701,In_2810);
nor U3809 (N_3809,In_2672,In_1665);
nand U3810 (N_3810,In_686,In_1992);
or U3811 (N_3811,In_1519,In_1535);
nand U3812 (N_3812,In_2067,In_701);
xnor U3813 (N_3813,In_2345,In_1503);
nand U3814 (N_3814,In_201,In_1184);
and U3815 (N_3815,In_1059,In_1622);
or U3816 (N_3816,In_2075,In_2491);
xor U3817 (N_3817,In_2954,In_1179);
and U3818 (N_3818,In_1047,In_1250);
nand U3819 (N_3819,In_876,In_294);
or U3820 (N_3820,In_211,In_2057);
or U3821 (N_3821,In_2760,In_1747);
nor U3822 (N_3822,In_593,In_2537);
nand U3823 (N_3823,In_2320,In_805);
nand U3824 (N_3824,In_483,In_1840);
or U3825 (N_3825,In_1499,In_317);
and U3826 (N_3826,In_2405,In_2708);
xor U3827 (N_3827,In_1442,In_1721);
nor U3828 (N_3828,In_1479,In_1586);
and U3829 (N_3829,In_1554,In_1810);
xnor U3830 (N_3830,In_1633,In_841);
nand U3831 (N_3831,In_608,In_1163);
and U3832 (N_3832,In_1378,In_1056);
nand U3833 (N_3833,In_558,In_2512);
nor U3834 (N_3834,In_312,In_89);
xor U3835 (N_3835,In_251,In_2560);
or U3836 (N_3836,In_1784,In_1298);
nor U3837 (N_3837,In_1909,In_1395);
nor U3838 (N_3838,In_606,In_803);
nand U3839 (N_3839,In_1721,In_2130);
and U3840 (N_3840,In_2901,In_1732);
or U3841 (N_3841,In_2900,In_1468);
xnor U3842 (N_3842,In_1877,In_1882);
xor U3843 (N_3843,In_774,In_1340);
xnor U3844 (N_3844,In_2671,In_2808);
nor U3845 (N_3845,In_2726,In_1198);
xor U3846 (N_3846,In_2565,In_51);
nor U3847 (N_3847,In_1120,In_562);
and U3848 (N_3848,In_1238,In_711);
xor U3849 (N_3849,In_1475,In_94);
nand U3850 (N_3850,In_2503,In_1431);
xor U3851 (N_3851,In_2784,In_1091);
xor U3852 (N_3852,In_2900,In_155);
or U3853 (N_3853,In_2894,In_2169);
nor U3854 (N_3854,In_662,In_1092);
nor U3855 (N_3855,In_1689,In_2081);
xnor U3856 (N_3856,In_91,In_1742);
nor U3857 (N_3857,In_1350,In_2293);
and U3858 (N_3858,In_144,In_2773);
nand U3859 (N_3859,In_2005,In_546);
xnor U3860 (N_3860,In_1630,In_2327);
nor U3861 (N_3861,In_109,In_2224);
nor U3862 (N_3862,In_1862,In_1211);
and U3863 (N_3863,In_2455,In_2685);
xnor U3864 (N_3864,In_2962,In_2024);
and U3865 (N_3865,In_1663,In_2766);
and U3866 (N_3866,In_2656,In_1068);
nor U3867 (N_3867,In_253,In_2933);
nand U3868 (N_3868,In_195,In_891);
or U3869 (N_3869,In_1949,In_829);
nor U3870 (N_3870,In_984,In_944);
or U3871 (N_3871,In_1038,In_1399);
nor U3872 (N_3872,In_263,In_1486);
or U3873 (N_3873,In_1653,In_1905);
nor U3874 (N_3874,In_2741,In_2369);
and U3875 (N_3875,In_731,In_891);
nor U3876 (N_3876,In_1092,In_1436);
xnor U3877 (N_3877,In_2502,In_2660);
nor U3878 (N_3878,In_1114,In_1478);
nand U3879 (N_3879,In_1359,In_329);
xor U3880 (N_3880,In_1279,In_927);
or U3881 (N_3881,In_2929,In_1670);
xor U3882 (N_3882,In_2313,In_2123);
nor U3883 (N_3883,In_1414,In_97);
or U3884 (N_3884,In_2881,In_2185);
nor U3885 (N_3885,In_441,In_1134);
and U3886 (N_3886,In_1844,In_1508);
nor U3887 (N_3887,In_777,In_2921);
nor U3888 (N_3888,In_381,In_2449);
nand U3889 (N_3889,In_2508,In_1607);
xor U3890 (N_3890,In_4,In_1610);
nand U3891 (N_3891,In_1765,In_185);
nor U3892 (N_3892,In_2489,In_1071);
nand U3893 (N_3893,In_1075,In_2032);
and U3894 (N_3894,In_1911,In_1445);
nand U3895 (N_3895,In_1453,In_1129);
xnor U3896 (N_3896,In_1837,In_351);
nor U3897 (N_3897,In_1544,In_2962);
or U3898 (N_3898,In_149,In_2065);
xor U3899 (N_3899,In_1707,In_1745);
and U3900 (N_3900,In_1084,In_1066);
or U3901 (N_3901,In_1781,In_375);
nor U3902 (N_3902,In_517,In_539);
and U3903 (N_3903,In_2038,In_1841);
and U3904 (N_3904,In_710,In_1129);
xnor U3905 (N_3905,In_780,In_1097);
or U3906 (N_3906,In_58,In_2646);
and U3907 (N_3907,In_650,In_105);
and U3908 (N_3908,In_661,In_2675);
nor U3909 (N_3909,In_593,In_1948);
or U3910 (N_3910,In_1334,In_2601);
xor U3911 (N_3911,In_1646,In_2406);
or U3912 (N_3912,In_2585,In_976);
or U3913 (N_3913,In_1335,In_2983);
xnor U3914 (N_3914,In_878,In_2450);
nor U3915 (N_3915,In_1113,In_555);
nand U3916 (N_3916,In_2790,In_1360);
or U3917 (N_3917,In_2653,In_631);
or U3918 (N_3918,In_2632,In_2915);
nand U3919 (N_3919,In_699,In_1852);
and U3920 (N_3920,In_2264,In_1334);
or U3921 (N_3921,In_2778,In_1046);
and U3922 (N_3922,In_1400,In_159);
nand U3923 (N_3923,In_1508,In_943);
xnor U3924 (N_3924,In_2555,In_255);
xor U3925 (N_3925,In_1015,In_2979);
xnor U3926 (N_3926,In_607,In_941);
nor U3927 (N_3927,In_1239,In_567);
xor U3928 (N_3928,In_1016,In_891);
xnor U3929 (N_3929,In_1358,In_2403);
nand U3930 (N_3930,In_219,In_2660);
nor U3931 (N_3931,In_1699,In_1617);
and U3932 (N_3932,In_3,In_27);
or U3933 (N_3933,In_240,In_923);
nor U3934 (N_3934,In_508,In_1470);
nor U3935 (N_3935,In_597,In_142);
xnor U3936 (N_3936,In_2453,In_784);
or U3937 (N_3937,In_237,In_2230);
or U3938 (N_3938,In_2598,In_436);
xnor U3939 (N_3939,In_2647,In_449);
or U3940 (N_3940,In_1604,In_672);
xnor U3941 (N_3941,In_2107,In_2557);
and U3942 (N_3942,In_2617,In_2370);
or U3943 (N_3943,In_2904,In_2111);
xnor U3944 (N_3944,In_327,In_388);
and U3945 (N_3945,In_1648,In_2198);
xnor U3946 (N_3946,In_1781,In_341);
or U3947 (N_3947,In_2484,In_1757);
or U3948 (N_3948,In_2418,In_978);
nor U3949 (N_3949,In_1561,In_1242);
nand U3950 (N_3950,In_18,In_602);
xnor U3951 (N_3951,In_2970,In_2044);
or U3952 (N_3952,In_420,In_2404);
nand U3953 (N_3953,In_1785,In_425);
or U3954 (N_3954,In_1136,In_1545);
and U3955 (N_3955,In_2440,In_657);
or U3956 (N_3956,In_1847,In_493);
or U3957 (N_3957,In_1288,In_2082);
nor U3958 (N_3958,In_2938,In_2033);
xor U3959 (N_3959,In_2281,In_1647);
xnor U3960 (N_3960,In_2591,In_2236);
and U3961 (N_3961,In_431,In_1920);
nand U3962 (N_3962,In_2717,In_297);
or U3963 (N_3963,In_466,In_1438);
nand U3964 (N_3964,In_2825,In_1892);
and U3965 (N_3965,In_270,In_726);
xnor U3966 (N_3966,In_1940,In_941);
or U3967 (N_3967,In_1838,In_2561);
xnor U3968 (N_3968,In_2826,In_71);
nor U3969 (N_3969,In_1811,In_2554);
and U3970 (N_3970,In_2459,In_1388);
nor U3971 (N_3971,In_2175,In_1412);
nand U3972 (N_3972,In_2537,In_2439);
xor U3973 (N_3973,In_2298,In_75);
nor U3974 (N_3974,In_68,In_1856);
xor U3975 (N_3975,In_1489,In_906);
or U3976 (N_3976,In_1719,In_812);
or U3977 (N_3977,In_10,In_1360);
nand U3978 (N_3978,In_2747,In_1854);
and U3979 (N_3979,In_1160,In_1945);
or U3980 (N_3980,In_1205,In_1257);
or U3981 (N_3981,In_1482,In_231);
xor U3982 (N_3982,In_274,In_1936);
or U3983 (N_3983,In_183,In_1184);
nand U3984 (N_3984,In_2468,In_988);
xnor U3985 (N_3985,In_706,In_2821);
and U3986 (N_3986,In_762,In_791);
xor U3987 (N_3987,In_1769,In_18);
and U3988 (N_3988,In_2505,In_1713);
nor U3989 (N_3989,In_884,In_2741);
nand U3990 (N_3990,In_2224,In_2312);
xnor U3991 (N_3991,In_2630,In_1636);
and U3992 (N_3992,In_1364,In_2196);
nor U3993 (N_3993,In_1701,In_2395);
xnor U3994 (N_3994,In_229,In_164);
and U3995 (N_3995,In_974,In_1680);
nor U3996 (N_3996,In_2482,In_865);
and U3997 (N_3997,In_2006,In_861);
xnor U3998 (N_3998,In_1065,In_43);
nand U3999 (N_3999,In_145,In_210);
nand U4000 (N_4000,In_1668,In_277);
nand U4001 (N_4001,In_2716,In_2155);
nor U4002 (N_4002,In_2197,In_84);
xnor U4003 (N_4003,In_1765,In_751);
or U4004 (N_4004,In_1020,In_1927);
or U4005 (N_4005,In_2067,In_2470);
nand U4006 (N_4006,In_2735,In_1686);
and U4007 (N_4007,In_281,In_2733);
xnor U4008 (N_4008,In_1110,In_428);
or U4009 (N_4009,In_2884,In_1955);
xnor U4010 (N_4010,In_2279,In_2476);
nor U4011 (N_4011,In_2685,In_493);
xnor U4012 (N_4012,In_2626,In_2159);
nand U4013 (N_4013,In_2977,In_2782);
or U4014 (N_4014,In_2956,In_2158);
or U4015 (N_4015,In_1410,In_855);
or U4016 (N_4016,In_717,In_1433);
nor U4017 (N_4017,In_968,In_296);
nand U4018 (N_4018,In_1622,In_2847);
nor U4019 (N_4019,In_96,In_794);
nor U4020 (N_4020,In_46,In_204);
nand U4021 (N_4021,In_2122,In_864);
xor U4022 (N_4022,In_674,In_1075);
and U4023 (N_4023,In_1670,In_2988);
nand U4024 (N_4024,In_2523,In_631);
nand U4025 (N_4025,In_1686,In_2128);
or U4026 (N_4026,In_178,In_1518);
or U4027 (N_4027,In_2055,In_579);
xor U4028 (N_4028,In_2611,In_25);
and U4029 (N_4029,In_2180,In_1940);
xor U4030 (N_4030,In_1433,In_1298);
xor U4031 (N_4031,In_2747,In_368);
xnor U4032 (N_4032,In_1987,In_395);
nand U4033 (N_4033,In_701,In_2213);
xor U4034 (N_4034,In_2005,In_896);
nand U4035 (N_4035,In_376,In_1523);
xnor U4036 (N_4036,In_2740,In_1993);
nor U4037 (N_4037,In_1538,In_2100);
and U4038 (N_4038,In_599,In_22);
or U4039 (N_4039,In_435,In_373);
nor U4040 (N_4040,In_410,In_590);
nand U4041 (N_4041,In_2765,In_2547);
nor U4042 (N_4042,In_1177,In_1784);
xnor U4043 (N_4043,In_1398,In_2118);
xnor U4044 (N_4044,In_2687,In_781);
nor U4045 (N_4045,In_97,In_920);
xnor U4046 (N_4046,In_1265,In_470);
and U4047 (N_4047,In_1028,In_2880);
nand U4048 (N_4048,In_1084,In_515);
and U4049 (N_4049,In_1660,In_611);
xnor U4050 (N_4050,In_949,In_2799);
and U4051 (N_4051,In_177,In_2621);
or U4052 (N_4052,In_543,In_1253);
and U4053 (N_4053,In_1359,In_1773);
and U4054 (N_4054,In_993,In_1110);
nor U4055 (N_4055,In_1611,In_1371);
and U4056 (N_4056,In_2133,In_1498);
nand U4057 (N_4057,In_2270,In_2430);
or U4058 (N_4058,In_1288,In_113);
and U4059 (N_4059,In_891,In_2365);
xnor U4060 (N_4060,In_210,In_280);
xnor U4061 (N_4061,In_2581,In_1989);
or U4062 (N_4062,In_1876,In_2121);
nor U4063 (N_4063,In_1771,In_526);
nand U4064 (N_4064,In_434,In_1368);
and U4065 (N_4065,In_2027,In_190);
or U4066 (N_4066,In_1709,In_1739);
nand U4067 (N_4067,In_198,In_2490);
or U4068 (N_4068,In_1109,In_1588);
and U4069 (N_4069,In_835,In_1385);
and U4070 (N_4070,In_2352,In_842);
and U4071 (N_4071,In_619,In_45);
and U4072 (N_4072,In_1357,In_2057);
and U4073 (N_4073,In_713,In_1602);
xnor U4074 (N_4074,In_2787,In_971);
nor U4075 (N_4075,In_737,In_1214);
nand U4076 (N_4076,In_1463,In_382);
or U4077 (N_4077,In_213,In_1573);
nand U4078 (N_4078,In_25,In_2338);
and U4079 (N_4079,In_2518,In_1273);
xor U4080 (N_4080,In_2352,In_710);
and U4081 (N_4081,In_1439,In_966);
and U4082 (N_4082,In_949,In_349);
and U4083 (N_4083,In_2200,In_1048);
nand U4084 (N_4084,In_882,In_1573);
nand U4085 (N_4085,In_1886,In_1376);
nand U4086 (N_4086,In_1101,In_2045);
nor U4087 (N_4087,In_1831,In_652);
xor U4088 (N_4088,In_1140,In_547);
or U4089 (N_4089,In_1521,In_154);
nand U4090 (N_4090,In_323,In_1497);
and U4091 (N_4091,In_476,In_726);
and U4092 (N_4092,In_1336,In_1793);
or U4093 (N_4093,In_1435,In_660);
and U4094 (N_4094,In_221,In_415);
and U4095 (N_4095,In_110,In_611);
nor U4096 (N_4096,In_1029,In_1940);
nand U4097 (N_4097,In_710,In_1595);
xnor U4098 (N_4098,In_2875,In_1266);
xor U4099 (N_4099,In_1823,In_547);
or U4100 (N_4100,In_955,In_2561);
or U4101 (N_4101,In_1855,In_1411);
or U4102 (N_4102,In_2259,In_554);
and U4103 (N_4103,In_217,In_65);
and U4104 (N_4104,In_1973,In_2108);
xor U4105 (N_4105,In_1865,In_2561);
nor U4106 (N_4106,In_1262,In_2475);
and U4107 (N_4107,In_1299,In_745);
nor U4108 (N_4108,In_858,In_2126);
nor U4109 (N_4109,In_682,In_1814);
and U4110 (N_4110,In_2282,In_1294);
and U4111 (N_4111,In_2719,In_1473);
nor U4112 (N_4112,In_902,In_2401);
or U4113 (N_4113,In_1775,In_1467);
or U4114 (N_4114,In_1761,In_531);
and U4115 (N_4115,In_2216,In_628);
and U4116 (N_4116,In_1717,In_1251);
nor U4117 (N_4117,In_1773,In_1286);
xor U4118 (N_4118,In_2205,In_2637);
nand U4119 (N_4119,In_253,In_2067);
xor U4120 (N_4120,In_2998,In_995);
xor U4121 (N_4121,In_2146,In_1457);
and U4122 (N_4122,In_1431,In_2689);
and U4123 (N_4123,In_593,In_113);
or U4124 (N_4124,In_180,In_1003);
nand U4125 (N_4125,In_1232,In_2743);
or U4126 (N_4126,In_1391,In_2931);
or U4127 (N_4127,In_219,In_2748);
xnor U4128 (N_4128,In_768,In_2190);
and U4129 (N_4129,In_2195,In_2152);
xnor U4130 (N_4130,In_2174,In_1480);
and U4131 (N_4131,In_1017,In_6);
xor U4132 (N_4132,In_853,In_2987);
nor U4133 (N_4133,In_1975,In_2891);
or U4134 (N_4134,In_1561,In_1353);
or U4135 (N_4135,In_781,In_2589);
and U4136 (N_4136,In_2893,In_1532);
or U4137 (N_4137,In_1165,In_831);
nand U4138 (N_4138,In_1812,In_1569);
nand U4139 (N_4139,In_2458,In_1358);
and U4140 (N_4140,In_782,In_532);
xnor U4141 (N_4141,In_2991,In_295);
nand U4142 (N_4142,In_2719,In_796);
nor U4143 (N_4143,In_759,In_1812);
and U4144 (N_4144,In_1789,In_1897);
or U4145 (N_4145,In_2737,In_1328);
nor U4146 (N_4146,In_2851,In_772);
and U4147 (N_4147,In_1781,In_470);
or U4148 (N_4148,In_507,In_763);
or U4149 (N_4149,In_2697,In_43);
nor U4150 (N_4150,In_1578,In_1744);
nand U4151 (N_4151,In_228,In_2436);
xor U4152 (N_4152,In_2657,In_646);
or U4153 (N_4153,In_2045,In_2993);
or U4154 (N_4154,In_2360,In_2939);
and U4155 (N_4155,In_1144,In_916);
nand U4156 (N_4156,In_2871,In_625);
nor U4157 (N_4157,In_1346,In_2484);
or U4158 (N_4158,In_911,In_888);
nor U4159 (N_4159,In_2059,In_2734);
and U4160 (N_4160,In_331,In_609);
and U4161 (N_4161,In_1718,In_763);
nand U4162 (N_4162,In_572,In_48);
and U4163 (N_4163,In_1176,In_684);
or U4164 (N_4164,In_2071,In_531);
nor U4165 (N_4165,In_2052,In_2283);
xor U4166 (N_4166,In_1285,In_690);
and U4167 (N_4167,In_486,In_2975);
and U4168 (N_4168,In_1464,In_6);
nand U4169 (N_4169,In_435,In_903);
nor U4170 (N_4170,In_1265,In_1962);
nor U4171 (N_4171,In_2267,In_39);
or U4172 (N_4172,In_1188,In_1991);
xor U4173 (N_4173,In_1444,In_2334);
nand U4174 (N_4174,In_2993,In_275);
or U4175 (N_4175,In_1824,In_296);
xor U4176 (N_4176,In_1485,In_2329);
nor U4177 (N_4177,In_2003,In_516);
and U4178 (N_4178,In_2207,In_1169);
xnor U4179 (N_4179,In_1648,In_844);
xnor U4180 (N_4180,In_1457,In_346);
xor U4181 (N_4181,In_1640,In_2176);
xor U4182 (N_4182,In_1856,In_410);
and U4183 (N_4183,In_2803,In_2477);
and U4184 (N_4184,In_2571,In_228);
and U4185 (N_4185,In_2258,In_2005);
xor U4186 (N_4186,In_216,In_737);
or U4187 (N_4187,In_187,In_2349);
and U4188 (N_4188,In_400,In_2287);
or U4189 (N_4189,In_1812,In_2181);
xnor U4190 (N_4190,In_2908,In_215);
nand U4191 (N_4191,In_1774,In_870);
nand U4192 (N_4192,In_110,In_1925);
xor U4193 (N_4193,In_617,In_126);
xnor U4194 (N_4194,In_379,In_1454);
and U4195 (N_4195,In_959,In_2075);
and U4196 (N_4196,In_289,In_2376);
and U4197 (N_4197,In_2111,In_803);
nor U4198 (N_4198,In_2451,In_1482);
nand U4199 (N_4199,In_1701,In_1402);
or U4200 (N_4200,In_1495,In_437);
and U4201 (N_4201,In_92,In_313);
and U4202 (N_4202,In_2158,In_1477);
nor U4203 (N_4203,In_1706,In_528);
and U4204 (N_4204,In_2089,In_2949);
nor U4205 (N_4205,In_128,In_1466);
nand U4206 (N_4206,In_1297,In_151);
nor U4207 (N_4207,In_752,In_1659);
xnor U4208 (N_4208,In_46,In_662);
xor U4209 (N_4209,In_115,In_234);
nand U4210 (N_4210,In_909,In_1481);
xnor U4211 (N_4211,In_437,In_671);
and U4212 (N_4212,In_1168,In_1044);
xor U4213 (N_4213,In_2718,In_520);
xnor U4214 (N_4214,In_1419,In_1951);
xor U4215 (N_4215,In_2075,In_2850);
nand U4216 (N_4216,In_2581,In_972);
and U4217 (N_4217,In_2509,In_1895);
xnor U4218 (N_4218,In_2483,In_1527);
nand U4219 (N_4219,In_972,In_2512);
nor U4220 (N_4220,In_627,In_1532);
xnor U4221 (N_4221,In_2239,In_2690);
or U4222 (N_4222,In_219,In_653);
and U4223 (N_4223,In_192,In_2418);
nand U4224 (N_4224,In_2690,In_2108);
nand U4225 (N_4225,In_2844,In_2180);
or U4226 (N_4226,In_2367,In_2514);
nor U4227 (N_4227,In_1694,In_2087);
xnor U4228 (N_4228,In_672,In_525);
or U4229 (N_4229,In_413,In_2090);
nor U4230 (N_4230,In_1768,In_1670);
or U4231 (N_4231,In_1958,In_2402);
nand U4232 (N_4232,In_1389,In_1381);
nor U4233 (N_4233,In_1800,In_1510);
and U4234 (N_4234,In_72,In_1507);
or U4235 (N_4235,In_2503,In_357);
and U4236 (N_4236,In_1710,In_2162);
and U4237 (N_4237,In_1380,In_2095);
and U4238 (N_4238,In_2957,In_837);
or U4239 (N_4239,In_1991,In_1383);
nand U4240 (N_4240,In_408,In_594);
xor U4241 (N_4241,In_1767,In_2723);
or U4242 (N_4242,In_791,In_1572);
nand U4243 (N_4243,In_2301,In_1566);
or U4244 (N_4244,In_1137,In_1033);
nor U4245 (N_4245,In_1415,In_984);
nand U4246 (N_4246,In_2476,In_2900);
or U4247 (N_4247,In_1735,In_1878);
nor U4248 (N_4248,In_553,In_608);
and U4249 (N_4249,In_998,In_968);
nor U4250 (N_4250,In_1272,In_5);
nand U4251 (N_4251,In_128,In_593);
xor U4252 (N_4252,In_789,In_742);
nand U4253 (N_4253,In_1806,In_881);
nor U4254 (N_4254,In_981,In_2632);
xor U4255 (N_4255,In_2989,In_689);
or U4256 (N_4256,In_880,In_1283);
nand U4257 (N_4257,In_2404,In_1213);
nand U4258 (N_4258,In_229,In_2254);
nor U4259 (N_4259,In_91,In_992);
and U4260 (N_4260,In_1142,In_2225);
or U4261 (N_4261,In_101,In_2835);
or U4262 (N_4262,In_147,In_2453);
nand U4263 (N_4263,In_976,In_610);
xnor U4264 (N_4264,In_1492,In_924);
or U4265 (N_4265,In_1705,In_2142);
nor U4266 (N_4266,In_1031,In_1835);
or U4267 (N_4267,In_157,In_2240);
nor U4268 (N_4268,In_317,In_1750);
and U4269 (N_4269,In_307,In_2224);
nor U4270 (N_4270,In_2046,In_1018);
xor U4271 (N_4271,In_26,In_1658);
or U4272 (N_4272,In_141,In_1648);
nand U4273 (N_4273,In_432,In_2528);
nor U4274 (N_4274,In_2673,In_233);
nand U4275 (N_4275,In_2147,In_2369);
and U4276 (N_4276,In_1617,In_1543);
or U4277 (N_4277,In_273,In_1451);
nand U4278 (N_4278,In_66,In_2438);
or U4279 (N_4279,In_397,In_2572);
nor U4280 (N_4280,In_884,In_896);
nor U4281 (N_4281,In_820,In_2146);
nand U4282 (N_4282,In_2030,In_214);
nand U4283 (N_4283,In_2783,In_594);
nor U4284 (N_4284,In_2079,In_2261);
nand U4285 (N_4285,In_1151,In_1469);
nand U4286 (N_4286,In_1736,In_740);
nor U4287 (N_4287,In_36,In_1278);
nor U4288 (N_4288,In_2757,In_645);
nor U4289 (N_4289,In_1135,In_1346);
and U4290 (N_4290,In_2286,In_2112);
nand U4291 (N_4291,In_928,In_2739);
nor U4292 (N_4292,In_679,In_1437);
xor U4293 (N_4293,In_2816,In_1385);
or U4294 (N_4294,In_806,In_535);
nor U4295 (N_4295,In_2916,In_2287);
nor U4296 (N_4296,In_654,In_143);
nor U4297 (N_4297,In_658,In_1277);
xor U4298 (N_4298,In_2898,In_2490);
nor U4299 (N_4299,In_1721,In_200);
nor U4300 (N_4300,In_798,In_1251);
or U4301 (N_4301,In_1387,In_1044);
xor U4302 (N_4302,In_2958,In_922);
xor U4303 (N_4303,In_2310,In_2372);
nand U4304 (N_4304,In_36,In_153);
nor U4305 (N_4305,In_783,In_2055);
xor U4306 (N_4306,In_1734,In_2924);
and U4307 (N_4307,In_14,In_1953);
or U4308 (N_4308,In_56,In_2937);
nand U4309 (N_4309,In_2005,In_1856);
xnor U4310 (N_4310,In_1002,In_1011);
nand U4311 (N_4311,In_853,In_894);
and U4312 (N_4312,In_2110,In_1990);
or U4313 (N_4313,In_338,In_664);
xor U4314 (N_4314,In_2448,In_982);
and U4315 (N_4315,In_1654,In_1376);
nand U4316 (N_4316,In_1621,In_2843);
and U4317 (N_4317,In_1781,In_2747);
nor U4318 (N_4318,In_1848,In_2309);
or U4319 (N_4319,In_2264,In_856);
and U4320 (N_4320,In_2886,In_1129);
and U4321 (N_4321,In_1636,In_1919);
and U4322 (N_4322,In_1409,In_173);
nor U4323 (N_4323,In_57,In_852);
xor U4324 (N_4324,In_2671,In_1877);
and U4325 (N_4325,In_2955,In_509);
nand U4326 (N_4326,In_2897,In_1623);
xor U4327 (N_4327,In_2991,In_207);
nand U4328 (N_4328,In_2269,In_109);
or U4329 (N_4329,In_1290,In_1452);
xnor U4330 (N_4330,In_2446,In_2117);
nand U4331 (N_4331,In_2931,In_1846);
nor U4332 (N_4332,In_154,In_302);
and U4333 (N_4333,In_2235,In_2265);
and U4334 (N_4334,In_579,In_2894);
nor U4335 (N_4335,In_25,In_1246);
or U4336 (N_4336,In_451,In_1975);
xor U4337 (N_4337,In_1340,In_35);
xor U4338 (N_4338,In_712,In_1276);
xnor U4339 (N_4339,In_296,In_1056);
xor U4340 (N_4340,In_2638,In_2995);
nand U4341 (N_4341,In_536,In_2957);
or U4342 (N_4342,In_2615,In_442);
xnor U4343 (N_4343,In_1012,In_301);
nand U4344 (N_4344,In_13,In_667);
or U4345 (N_4345,In_1892,In_2165);
nand U4346 (N_4346,In_2964,In_2589);
and U4347 (N_4347,In_1820,In_1288);
xnor U4348 (N_4348,In_1632,In_2881);
nor U4349 (N_4349,In_2198,In_1087);
or U4350 (N_4350,In_1892,In_696);
nor U4351 (N_4351,In_2943,In_1772);
nand U4352 (N_4352,In_2043,In_421);
nand U4353 (N_4353,In_905,In_2692);
xnor U4354 (N_4354,In_1234,In_160);
and U4355 (N_4355,In_553,In_1211);
nor U4356 (N_4356,In_1463,In_373);
and U4357 (N_4357,In_2782,In_1184);
nor U4358 (N_4358,In_1110,In_135);
and U4359 (N_4359,In_1431,In_1671);
nand U4360 (N_4360,In_783,In_715);
xnor U4361 (N_4361,In_2481,In_2117);
and U4362 (N_4362,In_1774,In_2728);
nor U4363 (N_4363,In_57,In_479);
nand U4364 (N_4364,In_2979,In_1634);
xor U4365 (N_4365,In_2444,In_1718);
xor U4366 (N_4366,In_1904,In_1441);
nor U4367 (N_4367,In_674,In_1198);
xnor U4368 (N_4368,In_1882,In_2044);
nand U4369 (N_4369,In_2192,In_2742);
nor U4370 (N_4370,In_625,In_624);
nor U4371 (N_4371,In_1215,In_1021);
and U4372 (N_4372,In_2695,In_1417);
nand U4373 (N_4373,In_2980,In_2187);
nand U4374 (N_4374,In_2615,In_2559);
nand U4375 (N_4375,In_521,In_2494);
nand U4376 (N_4376,In_2682,In_2129);
nand U4377 (N_4377,In_2279,In_2428);
nand U4378 (N_4378,In_2045,In_1992);
or U4379 (N_4379,In_340,In_946);
nand U4380 (N_4380,In_2441,In_2271);
or U4381 (N_4381,In_120,In_747);
and U4382 (N_4382,In_1709,In_1649);
xnor U4383 (N_4383,In_1241,In_766);
and U4384 (N_4384,In_1581,In_2645);
xnor U4385 (N_4385,In_1392,In_619);
or U4386 (N_4386,In_2448,In_470);
xor U4387 (N_4387,In_2101,In_2353);
nand U4388 (N_4388,In_1947,In_883);
nor U4389 (N_4389,In_1714,In_2279);
xor U4390 (N_4390,In_1756,In_2872);
or U4391 (N_4391,In_1754,In_283);
nand U4392 (N_4392,In_1204,In_1199);
nand U4393 (N_4393,In_274,In_2212);
and U4394 (N_4394,In_2517,In_1414);
and U4395 (N_4395,In_253,In_64);
xor U4396 (N_4396,In_875,In_754);
or U4397 (N_4397,In_2064,In_2526);
and U4398 (N_4398,In_1867,In_2668);
nor U4399 (N_4399,In_2269,In_2044);
xor U4400 (N_4400,In_220,In_125);
nor U4401 (N_4401,In_2808,In_2017);
nor U4402 (N_4402,In_2606,In_2822);
nand U4403 (N_4403,In_1134,In_2992);
and U4404 (N_4404,In_690,In_2499);
and U4405 (N_4405,In_230,In_1492);
and U4406 (N_4406,In_2321,In_2281);
or U4407 (N_4407,In_2850,In_2123);
and U4408 (N_4408,In_2375,In_155);
nand U4409 (N_4409,In_42,In_587);
and U4410 (N_4410,In_2686,In_562);
xor U4411 (N_4411,In_2000,In_390);
nor U4412 (N_4412,In_1326,In_2006);
and U4413 (N_4413,In_1372,In_71);
xor U4414 (N_4414,In_188,In_2308);
nor U4415 (N_4415,In_2201,In_762);
nor U4416 (N_4416,In_1621,In_2701);
or U4417 (N_4417,In_587,In_1319);
and U4418 (N_4418,In_1740,In_1470);
xor U4419 (N_4419,In_2458,In_1088);
nand U4420 (N_4420,In_784,In_2440);
nand U4421 (N_4421,In_246,In_1762);
nand U4422 (N_4422,In_1954,In_7);
and U4423 (N_4423,In_1056,In_2442);
and U4424 (N_4424,In_1562,In_2263);
xor U4425 (N_4425,In_23,In_1242);
nand U4426 (N_4426,In_2722,In_443);
and U4427 (N_4427,In_2013,In_2004);
xor U4428 (N_4428,In_470,In_1371);
or U4429 (N_4429,In_1231,In_1766);
nand U4430 (N_4430,In_2254,In_1822);
or U4431 (N_4431,In_343,In_828);
xor U4432 (N_4432,In_1608,In_717);
or U4433 (N_4433,In_1880,In_1215);
and U4434 (N_4434,In_1741,In_14);
nand U4435 (N_4435,In_55,In_2805);
nor U4436 (N_4436,In_1787,In_2182);
xor U4437 (N_4437,In_1410,In_869);
and U4438 (N_4438,In_1973,In_1542);
and U4439 (N_4439,In_2029,In_1992);
xor U4440 (N_4440,In_532,In_2843);
nand U4441 (N_4441,In_1968,In_2594);
and U4442 (N_4442,In_1162,In_447);
nor U4443 (N_4443,In_348,In_506);
or U4444 (N_4444,In_508,In_2660);
nand U4445 (N_4445,In_843,In_2909);
or U4446 (N_4446,In_949,In_896);
and U4447 (N_4447,In_2623,In_109);
nand U4448 (N_4448,In_841,In_470);
nor U4449 (N_4449,In_2838,In_709);
or U4450 (N_4450,In_2535,In_90);
and U4451 (N_4451,In_2685,In_2436);
nor U4452 (N_4452,In_916,In_2460);
xor U4453 (N_4453,In_1051,In_341);
or U4454 (N_4454,In_403,In_2977);
or U4455 (N_4455,In_1936,In_896);
xor U4456 (N_4456,In_2515,In_1210);
nand U4457 (N_4457,In_487,In_649);
or U4458 (N_4458,In_1410,In_696);
xnor U4459 (N_4459,In_2660,In_2001);
nor U4460 (N_4460,In_109,In_2582);
xnor U4461 (N_4461,In_736,In_1088);
xor U4462 (N_4462,In_2484,In_1339);
nand U4463 (N_4463,In_2868,In_1304);
nand U4464 (N_4464,In_2277,In_2423);
nor U4465 (N_4465,In_2373,In_1536);
or U4466 (N_4466,In_2058,In_2282);
xnor U4467 (N_4467,In_2799,In_582);
xnor U4468 (N_4468,In_2353,In_1882);
nor U4469 (N_4469,In_167,In_1628);
nand U4470 (N_4470,In_2801,In_2588);
nand U4471 (N_4471,In_557,In_439);
nor U4472 (N_4472,In_273,In_1676);
nor U4473 (N_4473,In_1670,In_2007);
nor U4474 (N_4474,In_1569,In_2689);
nor U4475 (N_4475,In_894,In_1078);
nor U4476 (N_4476,In_821,In_829);
xor U4477 (N_4477,In_2854,In_1064);
and U4478 (N_4478,In_1216,In_1002);
nor U4479 (N_4479,In_281,In_2047);
nand U4480 (N_4480,In_2261,In_2041);
or U4481 (N_4481,In_1906,In_2681);
and U4482 (N_4482,In_758,In_1067);
nor U4483 (N_4483,In_1150,In_1952);
nor U4484 (N_4484,In_1275,In_2604);
and U4485 (N_4485,In_319,In_1077);
nand U4486 (N_4486,In_2766,In_2059);
xnor U4487 (N_4487,In_118,In_2825);
and U4488 (N_4488,In_856,In_710);
and U4489 (N_4489,In_105,In_2134);
and U4490 (N_4490,In_195,In_1848);
and U4491 (N_4491,In_1054,In_1784);
nor U4492 (N_4492,In_1833,In_2103);
nor U4493 (N_4493,In_950,In_302);
and U4494 (N_4494,In_922,In_2169);
nand U4495 (N_4495,In_2017,In_1593);
nand U4496 (N_4496,In_1574,In_738);
nor U4497 (N_4497,In_824,In_2278);
nand U4498 (N_4498,In_79,In_105);
and U4499 (N_4499,In_1880,In_164);
and U4500 (N_4500,In_755,In_878);
and U4501 (N_4501,In_1126,In_1761);
nor U4502 (N_4502,In_1244,In_825);
or U4503 (N_4503,In_2980,In_925);
and U4504 (N_4504,In_2955,In_2011);
nand U4505 (N_4505,In_1753,In_2859);
xnor U4506 (N_4506,In_517,In_1913);
nor U4507 (N_4507,In_659,In_2032);
nand U4508 (N_4508,In_1969,In_313);
and U4509 (N_4509,In_476,In_1161);
and U4510 (N_4510,In_798,In_2836);
nor U4511 (N_4511,In_855,In_1433);
or U4512 (N_4512,In_928,In_2468);
and U4513 (N_4513,In_900,In_1586);
xor U4514 (N_4514,In_423,In_897);
nand U4515 (N_4515,In_5,In_1583);
nor U4516 (N_4516,In_2546,In_394);
xnor U4517 (N_4517,In_1537,In_1965);
nand U4518 (N_4518,In_1831,In_2367);
nor U4519 (N_4519,In_2074,In_1608);
xnor U4520 (N_4520,In_142,In_545);
nor U4521 (N_4521,In_1607,In_171);
and U4522 (N_4522,In_2550,In_2337);
and U4523 (N_4523,In_1830,In_2857);
xnor U4524 (N_4524,In_642,In_1077);
nor U4525 (N_4525,In_2690,In_2896);
nand U4526 (N_4526,In_1624,In_2299);
and U4527 (N_4527,In_770,In_2850);
or U4528 (N_4528,In_2774,In_1830);
xnor U4529 (N_4529,In_1639,In_2004);
or U4530 (N_4530,In_326,In_574);
xnor U4531 (N_4531,In_2199,In_1802);
or U4532 (N_4532,In_2738,In_1441);
or U4533 (N_4533,In_493,In_1760);
and U4534 (N_4534,In_1313,In_2427);
nand U4535 (N_4535,In_1277,In_50);
and U4536 (N_4536,In_1505,In_450);
or U4537 (N_4537,In_645,In_464);
xor U4538 (N_4538,In_61,In_820);
or U4539 (N_4539,In_2659,In_223);
nand U4540 (N_4540,In_1940,In_1410);
and U4541 (N_4541,In_443,In_2447);
xor U4542 (N_4542,In_36,In_2980);
xor U4543 (N_4543,In_720,In_642);
or U4544 (N_4544,In_2292,In_2163);
nor U4545 (N_4545,In_2497,In_2762);
xnor U4546 (N_4546,In_1867,In_2932);
xor U4547 (N_4547,In_2533,In_2841);
and U4548 (N_4548,In_1059,In_991);
nor U4549 (N_4549,In_2381,In_422);
nand U4550 (N_4550,In_1678,In_206);
xnor U4551 (N_4551,In_2008,In_2778);
and U4552 (N_4552,In_1724,In_1575);
nor U4553 (N_4553,In_2334,In_172);
nor U4554 (N_4554,In_211,In_1606);
nand U4555 (N_4555,In_391,In_1855);
and U4556 (N_4556,In_63,In_1338);
and U4557 (N_4557,In_419,In_2468);
xnor U4558 (N_4558,In_526,In_1798);
or U4559 (N_4559,In_853,In_1907);
xor U4560 (N_4560,In_524,In_1607);
nor U4561 (N_4561,In_1581,In_2995);
and U4562 (N_4562,In_1821,In_2842);
and U4563 (N_4563,In_1578,In_1550);
nand U4564 (N_4564,In_1131,In_1073);
nor U4565 (N_4565,In_1466,In_432);
nor U4566 (N_4566,In_2687,In_1112);
or U4567 (N_4567,In_395,In_459);
nand U4568 (N_4568,In_407,In_880);
nand U4569 (N_4569,In_1491,In_2652);
and U4570 (N_4570,In_2621,In_1514);
nor U4571 (N_4571,In_1933,In_2623);
xor U4572 (N_4572,In_2763,In_1083);
or U4573 (N_4573,In_2012,In_2713);
xnor U4574 (N_4574,In_109,In_246);
nand U4575 (N_4575,In_1449,In_253);
nand U4576 (N_4576,In_2865,In_378);
xnor U4577 (N_4577,In_2287,In_2091);
or U4578 (N_4578,In_790,In_1699);
or U4579 (N_4579,In_1535,In_1838);
nand U4580 (N_4580,In_95,In_579);
nor U4581 (N_4581,In_898,In_785);
or U4582 (N_4582,In_1709,In_2776);
xor U4583 (N_4583,In_642,In_710);
nand U4584 (N_4584,In_2302,In_2634);
or U4585 (N_4585,In_2316,In_551);
and U4586 (N_4586,In_2859,In_1856);
nand U4587 (N_4587,In_2137,In_263);
nand U4588 (N_4588,In_957,In_2771);
or U4589 (N_4589,In_2233,In_898);
xnor U4590 (N_4590,In_598,In_2626);
and U4591 (N_4591,In_2890,In_575);
and U4592 (N_4592,In_1412,In_1006);
and U4593 (N_4593,In_1033,In_1636);
xnor U4594 (N_4594,In_1250,In_81);
and U4595 (N_4595,In_1054,In_1899);
and U4596 (N_4596,In_1172,In_469);
nor U4597 (N_4597,In_2027,In_1642);
nand U4598 (N_4598,In_2008,In_1743);
and U4599 (N_4599,In_527,In_1580);
xnor U4600 (N_4600,In_2179,In_1671);
xor U4601 (N_4601,In_1445,In_2779);
and U4602 (N_4602,In_1486,In_2374);
xor U4603 (N_4603,In_2695,In_9);
nand U4604 (N_4604,In_2531,In_2987);
and U4605 (N_4605,In_1609,In_1422);
and U4606 (N_4606,In_367,In_571);
nand U4607 (N_4607,In_1699,In_1720);
and U4608 (N_4608,In_117,In_2170);
nor U4609 (N_4609,In_1428,In_2543);
and U4610 (N_4610,In_2672,In_687);
nand U4611 (N_4611,In_599,In_227);
nor U4612 (N_4612,In_2416,In_1529);
xor U4613 (N_4613,In_1396,In_1531);
xnor U4614 (N_4614,In_1022,In_2683);
and U4615 (N_4615,In_1677,In_1851);
xor U4616 (N_4616,In_1071,In_2020);
nor U4617 (N_4617,In_1108,In_2196);
or U4618 (N_4618,In_1827,In_1338);
nand U4619 (N_4619,In_1363,In_1184);
or U4620 (N_4620,In_2083,In_1013);
and U4621 (N_4621,In_2882,In_2032);
xor U4622 (N_4622,In_2433,In_2286);
nand U4623 (N_4623,In_592,In_8);
nand U4624 (N_4624,In_1631,In_1935);
or U4625 (N_4625,In_1838,In_693);
xnor U4626 (N_4626,In_108,In_2151);
xor U4627 (N_4627,In_2391,In_22);
nor U4628 (N_4628,In_2192,In_1703);
xnor U4629 (N_4629,In_2148,In_536);
or U4630 (N_4630,In_2329,In_2458);
nor U4631 (N_4631,In_1620,In_2466);
and U4632 (N_4632,In_1848,In_1169);
and U4633 (N_4633,In_2082,In_2548);
or U4634 (N_4634,In_1254,In_2303);
or U4635 (N_4635,In_528,In_1948);
xor U4636 (N_4636,In_1031,In_1045);
nor U4637 (N_4637,In_1355,In_26);
nor U4638 (N_4638,In_1721,In_904);
nor U4639 (N_4639,In_1516,In_941);
and U4640 (N_4640,In_767,In_1987);
or U4641 (N_4641,In_985,In_264);
or U4642 (N_4642,In_2001,In_2875);
nand U4643 (N_4643,In_2319,In_2944);
nor U4644 (N_4644,In_1151,In_1134);
xnor U4645 (N_4645,In_1868,In_1891);
xor U4646 (N_4646,In_557,In_2792);
or U4647 (N_4647,In_2662,In_882);
or U4648 (N_4648,In_697,In_955);
xnor U4649 (N_4649,In_2386,In_2198);
nor U4650 (N_4650,In_1162,In_558);
xnor U4651 (N_4651,In_122,In_1583);
nor U4652 (N_4652,In_750,In_2373);
or U4653 (N_4653,In_558,In_1242);
nand U4654 (N_4654,In_1087,In_1038);
nor U4655 (N_4655,In_409,In_2103);
nor U4656 (N_4656,In_2586,In_2731);
xor U4657 (N_4657,In_2194,In_186);
and U4658 (N_4658,In_1343,In_958);
and U4659 (N_4659,In_1909,In_2607);
or U4660 (N_4660,In_1453,In_2946);
or U4661 (N_4661,In_1761,In_1688);
and U4662 (N_4662,In_1330,In_2374);
nand U4663 (N_4663,In_2416,In_2415);
and U4664 (N_4664,In_1073,In_1536);
and U4665 (N_4665,In_2003,In_1331);
and U4666 (N_4666,In_4,In_1364);
and U4667 (N_4667,In_1169,In_135);
xnor U4668 (N_4668,In_1037,In_1357);
xor U4669 (N_4669,In_1058,In_2004);
xnor U4670 (N_4670,In_433,In_229);
and U4671 (N_4671,In_2322,In_793);
nor U4672 (N_4672,In_1062,In_152);
nand U4673 (N_4673,In_1082,In_2953);
nand U4674 (N_4674,In_2736,In_1371);
xnor U4675 (N_4675,In_751,In_2955);
nand U4676 (N_4676,In_2518,In_2032);
nor U4677 (N_4677,In_1416,In_1953);
and U4678 (N_4678,In_892,In_2544);
nand U4679 (N_4679,In_695,In_377);
or U4680 (N_4680,In_2406,In_2976);
and U4681 (N_4681,In_28,In_1557);
and U4682 (N_4682,In_411,In_2125);
xor U4683 (N_4683,In_967,In_2643);
xor U4684 (N_4684,In_1464,In_1655);
nor U4685 (N_4685,In_1624,In_1593);
nor U4686 (N_4686,In_1377,In_1772);
nor U4687 (N_4687,In_1945,In_2857);
nand U4688 (N_4688,In_2958,In_1033);
xor U4689 (N_4689,In_434,In_504);
nand U4690 (N_4690,In_197,In_917);
nor U4691 (N_4691,In_2613,In_999);
and U4692 (N_4692,In_2696,In_2111);
xnor U4693 (N_4693,In_1504,In_828);
and U4694 (N_4694,In_370,In_1084);
or U4695 (N_4695,In_2076,In_1132);
xor U4696 (N_4696,In_2978,In_2732);
or U4697 (N_4697,In_702,In_1419);
or U4698 (N_4698,In_2568,In_574);
nand U4699 (N_4699,In_1840,In_1815);
xnor U4700 (N_4700,In_1640,In_2026);
nand U4701 (N_4701,In_231,In_1578);
and U4702 (N_4702,In_347,In_937);
or U4703 (N_4703,In_300,In_109);
xor U4704 (N_4704,In_704,In_1214);
nand U4705 (N_4705,In_542,In_2046);
nand U4706 (N_4706,In_16,In_2650);
xor U4707 (N_4707,In_1681,In_1208);
xnor U4708 (N_4708,In_2277,In_1186);
nand U4709 (N_4709,In_2858,In_2532);
nand U4710 (N_4710,In_2714,In_357);
and U4711 (N_4711,In_1604,In_1301);
and U4712 (N_4712,In_1959,In_2972);
or U4713 (N_4713,In_2722,In_2205);
and U4714 (N_4714,In_1122,In_2614);
nand U4715 (N_4715,In_46,In_1622);
xor U4716 (N_4716,In_2374,In_2626);
or U4717 (N_4717,In_525,In_2604);
xnor U4718 (N_4718,In_1034,In_719);
nand U4719 (N_4719,In_682,In_128);
and U4720 (N_4720,In_481,In_2976);
xnor U4721 (N_4721,In_328,In_1989);
xnor U4722 (N_4722,In_1556,In_1297);
nor U4723 (N_4723,In_144,In_904);
and U4724 (N_4724,In_1305,In_2492);
or U4725 (N_4725,In_2858,In_1476);
nand U4726 (N_4726,In_896,In_2064);
or U4727 (N_4727,In_1451,In_508);
and U4728 (N_4728,In_2321,In_1229);
or U4729 (N_4729,In_1258,In_2445);
or U4730 (N_4730,In_1463,In_1962);
nand U4731 (N_4731,In_1790,In_2835);
and U4732 (N_4732,In_1677,In_2009);
xor U4733 (N_4733,In_366,In_1864);
nor U4734 (N_4734,In_226,In_322);
nand U4735 (N_4735,In_1882,In_1483);
or U4736 (N_4736,In_1843,In_1684);
nand U4737 (N_4737,In_2942,In_1872);
nand U4738 (N_4738,In_1863,In_2232);
xor U4739 (N_4739,In_2479,In_888);
nand U4740 (N_4740,In_1526,In_1394);
nand U4741 (N_4741,In_1730,In_710);
xnor U4742 (N_4742,In_1890,In_2177);
and U4743 (N_4743,In_341,In_2002);
xor U4744 (N_4744,In_419,In_1772);
xor U4745 (N_4745,In_362,In_1264);
or U4746 (N_4746,In_2929,In_1059);
nand U4747 (N_4747,In_135,In_1084);
xor U4748 (N_4748,In_389,In_977);
or U4749 (N_4749,In_502,In_254);
nor U4750 (N_4750,In_1357,In_1025);
nand U4751 (N_4751,In_23,In_878);
and U4752 (N_4752,In_1319,In_2849);
nand U4753 (N_4753,In_2688,In_1248);
or U4754 (N_4754,In_348,In_1402);
nor U4755 (N_4755,In_1831,In_1258);
and U4756 (N_4756,In_2298,In_1315);
and U4757 (N_4757,In_1597,In_1678);
and U4758 (N_4758,In_1004,In_242);
or U4759 (N_4759,In_2004,In_319);
xnor U4760 (N_4760,In_2370,In_1418);
xnor U4761 (N_4761,In_2573,In_1086);
or U4762 (N_4762,In_1995,In_1399);
xnor U4763 (N_4763,In_853,In_2133);
or U4764 (N_4764,In_439,In_1904);
or U4765 (N_4765,In_1966,In_1345);
or U4766 (N_4766,In_1347,In_2296);
nor U4767 (N_4767,In_751,In_1681);
nor U4768 (N_4768,In_934,In_1959);
and U4769 (N_4769,In_2082,In_1161);
or U4770 (N_4770,In_1012,In_1137);
nand U4771 (N_4771,In_2342,In_1127);
and U4772 (N_4772,In_168,In_1856);
xor U4773 (N_4773,In_2499,In_992);
or U4774 (N_4774,In_2937,In_2734);
xnor U4775 (N_4775,In_157,In_2937);
and U4776 (N_4776,In_1225,In_304);
or U4777 (N_4777,In_1886,In_975);
nand U4778 (N_4778,In_86,In_262);
or U4779 (N_4779,In_1729,In_2689);
nor U4780 (N_4780,In_1770,In_1428);
nand U4781 (N_4781,In_608,In_210);
xor U4782 (N_4782,In_1804,In_1968);
and U4783 (N_4783,In_1248,In_484);
nor U4784 (N_4784,In_20,In_559);
nor U4785 (N_4785,In_1830,In_2949);
or U4786 (N_4786,In_2774,In_1357);
nand U4787 (N_4787,In_2141,In_2168);
xor U4788 (N_4788,In_2080,In_1471);
xnor U4789 (N_4789,In_1906,In_963);
and U4790 (N_4790,In_190,In_2760);
or U4791 (N_4791,In_1930,In_208);
nand U4792 (N_4792,In_1088,In_1580);
and U4793 (N_4793,In_1929,In_2997);
nor U4794 (N_4794,In_2798,In_651);
nor U4795 (N_4795,In_1669,In_2577);
and U4796 (N_4796,In_2839,In_2507);
nor U4797 (N_4797,In_1206,In_1173);
or U4798 (N_4798,In_596,In_1601);
or U4799 (N_4799,In_2412,In_259);
nor U4800 (N_4800,In_2967,In_2189);
or U4801 (N_4801,In_886,In_2653);
nand U4802 (N_4802,In_2366,In_2702);
xnor U4803 (N_4803,In_2740,In_946);
or U4804 (N_4804,In_2479,In_1960);
nor U4805 (N_4805,In_2995,In_600);
xnor U4806 (N_4806,In_1373,In_1105);
xnor U4807 (N_4807,In_1576,In_2111);
or U4808 (N_4808,In_2014,In_592);
nand U4809 (N_4809,In_432,In_800);
or U4810 (N_4810,In_994,In_1686);
nand U4811 (N_4811,In_1344,In_404);
nor U4812 (N_4812,In_1073,In_1550);
or U4813 (N_4813,In_767,In_451);
nor U4814 (N_4814,In_931,In_1419);
or U4815 (N_4815,In_1234,In_458);
nor U4816 (N_4816,In_1853,In_29);
and U4817 (N_4817,In_2604,In_2613);
xnor U4818 (N_4818,In_812,In_545);
xnor U4819 (N_4819,In_2548,In_2866);
or U4820 (N_4820,In_1979,In_2107);
and U4821 (N_4821,In_1419,In_1767);
nand U4822 (N_4822,In_1149,In_1382);
nor U4823 (N_4823,In_1290,In_1802);
nor U4824 (N_4824,In_1404,In_1370);
or U4825 (N_4825,In_2030,In_1128);
or U4826 (N_4826,In_2472,In_1263);
nand U4827 (N_4827,In_2106,In_922);
or U4828 (N_4828,In_1674,In_1449);
xor U4829 (N_4829,In_2846,In_948);
xnor U4830 (N_4830,In_2192,In_2069);
and U4831 (N_4831,In_2802,In_1264);
nand U4832 (N_4832,In_272,In_764);
and U4833 (N_4833,In_2620,In_2054);
or U4834 (N_4834,In_656,In_645);
or U4835 (N_4835,In_1890,In_2851);
xor U4836 (N_4836,In_1071,In_916);
and U4837 (N_4837,In_316,In_9);
nor U4838 (N_4838,In_1563,In_1950);
xor U4839 (N_4839,In_113,In_2679);
xnor U4840 (N_4840,In_2660,In_1117);
and U4841 (N_4841,In_1565,In_2941);
and U4842 (N_4842,In_1244,In_384);
and U4843 (N_4843,In_1757,In_33);
and U4844 (N_4844,In_1035,In_373);
nor U4845 (N_4845,In_677,In_336);
or U4846 (N_4846,In_2492,In_2960);
nor U4847 (N_4847,In_1751,In_410);
and U4848 (N_4848,In_680,In_1717);
xnor U4849 (N_4849,In_342,In_899);
xnor U4850 (N_4850,In_876,In_2357);
xor U4851 (N_4851,In_1250,In_2176);
and U4852 (N_4852,In_2954,In_2501);
and U4853 (N_4853,In_456,In_2229);
nor U4854 (N_4854,In_2257,In_2690);
nand U4855 (N_4855,In_2168,In_2001);
and U4856 (N_4856,In_1540,In_2425);
nor U4857 (N_4857,In_2294,In_1252);
xnor U4858 (N_4858,In_1756,In_1028);
and U4859 (N_4859,In_2892,In_394);
nor U4860 (N_4860,In_774,In_2389);
xor U4861 (N_4861,In_657,In_2992);
nor U4862 (N_4862,In_853,In_2836);
and U4863 (N_4863,In_184,In_251);
xor U4864 (N_4864,In_743,In_2573);
or U4865 (N_4865,In_2834,In_2890);
xor U4866 (N_4866,In_2697,In_2348);
nand U4867 (N_4867,In_2133,In_2438);
nor U4868 (N_4868,In_1912,In_457);
xor U4869 (N_4869,In_1650,In_1752);
nor U4870 (N_4870,In_2003,In_397);
or U4871 (N_4871,In_988,In_1605);
or U4872 (N_4872,In_577,In_1002);
or U4873 (N_4873,In_204,In_2251);
nor U4874 (N_4874,In_1831,In_972);
or U4875 (N_4875,In_1821,In_2441);
and U4876 (N_4876,In_763,In_1331);
and U4877 (N_4877,In_123,In_953);
nor U4878 (N_4878,In_2738,In_2265);
nand U4879 (N_4879,In_661,In_2567);
nor U4880 (N_4880,In_556,In_808);
or U4881 (N_4881,In_583,In_302);
and U4882 (N_4882,In_556,In_2254);
nor U4883 (N_4883,In_958,In_1109);
nand U4884 (N_4884,In_1863,In_2156);
nand U4885 (N_4885,In_2946,In_2347);
nand U4886 (N_4886,In_2607,In_1404);
or U4887 (N_4887,In_2598,In_928);
nand U4888 (N_4888,In_2193,In_1440);
and U4889 (N_4889,In_2074,In_806);
xnor U4890 (N_4890,In_849,In_155);
or U4891 (N_4891,In_1684,In_1020);
or U4892 (N_4892,In_646,In_638);
nor U4893 (N_4893,In_130,In_1440);
and U4894 (N_4894,In_101,In_527);
or U4895 (N_4895,In_23,In_2812);
xor U4896 (N_4896,In_2262,In_2589);
nor U4897 (N_4897,In_955,In_2684);
xnor U4898 (N_4898,In_1371,In_334);
nand U4899 (N_4899,In_1072,In_1591);
nor U4900 (N_4900,In_1403,In_2042);
xor U4901 (N_4901,In_1172,In_1199);
nand U4902 (N_4902,In_407,In_1351);
or U4903 (N_4903,In_1432,In_748);
and U4904 (N_4904,In_155,In_2005);
nand U4905 (N_4905,In_2736,In_2940);
nor U4906 (N_4906,In_1920,In_570);
nor U4907 (N_4907,In_739,In_394);
or U4908 (N_4908,In_2250,In_1633);
nor U4909 (N_4909,In_2085,In_192);
and U4910 (N_4910,In_1592,In_1699);
nor U4911 (N_4911,In_336,In_548);
nor U4912 (N_4912,In_977,In_918);
or U4913 (N_4913,In_2032,In_1578);
and U4914 (N_4914,In_2467,In_2868);
xnor U4915 (N_4915,In_580,In_2897);
nor U4916 (N_4916,In_1402,In_2478);
or U4917 (N_4917,In_1553,In_903);
and U4918 (N_4918,In_447,In_250);
nor U4919 (N_4919,In_539,In_100);
or U4920 (N_4920,In_1086,In_1776);
xnor U4921 (N_4921,In_1768,In_79);
xor U4922 (N_4922,In_1487,In_2420);
nand U4923 (N_4923,In_2155,In_947);
or U4924 (N_4924,In_1741,In_2203);
nor U4925 (N_4925,In_433,In_2153);
nand U4926 (N_4926,In_976,In_999);
or U4927 (N_4927,In_698,In_2934);
and U4928 (N_4928,In_716,In_1085);
nand U4929 (N_4929,In_2267,In_2991);
or U4930 (N_4930,In_1923,In_1711);
nand U4931 (N_4931,In_2903,In_848);
nand U4932 (N_4932,In_589,In_1054);
or U4933 (N_4933,In_2304,In_2251);
xnor U4934 (N_4934,In_1392,In_625);
nand U4935 (N_4935,In_1091,In_604);
nand U4936 (N_4936,In_1480,In_1333);
or U4937 (N_4937,In_311,In_1274);
and U4938 (N_4938,In_2765,In_637);
or U4939 (N_4939,In_824,In_1143);
nor U4940 (N_4940,In_2970,In_1010);
nand U4941 (N_4941,In_262,In_2740);
nor U4942 (N_4942,In_1491,In_1516);
nand U4943 (N_4943,In_559,In_1528);
and U4944 (N_4944,In_1542,In_797);
and U4945 (N_4945,In_1544,In_290);
or U4946 (N_4946,In_155,In_2393);
or U4947 (N_4947,In_1928,In_643);
or U4948 (N_4948,In_1522,In_94);
nor U4949 (N_4949,In_2871,In_291);
and U4950 (N_4950,In_2434,In_2043);
or U4951 (N_4951,In_1799,In_984);
nor U4952 (N_4952,In_1849,In_1753);
and U4953 (N_4953,In_887,In_1649);
nand U4954 (N_4954,In_883,In_661);
xor U4955 (N_4955,In_1391,In_123);
nor U4956 (N_4956,In_1963,In_570);
xor U4957 (N_4957,In_2548,In_1927);
or U4958 (N_4958,In_539,In_1416);
nor U4959 (N_4959,In_2467,In_1557);
or U4960 (N_4960,In_1122,In_2827);
nand U4961 (N_4961,In_959,In_1591);
and U4962 (N_4962,In_269,In_2656);
nand U4963 (N_4963,In_1940,In_150);
or U4964 (N_4964,In_2857,In_2616);
nor U4965 (N_4965,In_298,In_2050);
xor U4966 (N_4966,In_1857,In_267);
and U4967 (N_4967,In_2103,In_1022);
nor U4968 (N_4968,In_498,In_2319);
nor U4969 (N_4969,In_1658,In_2592);
xor U4970 (N_4970,In_2881,In_2585);
nor U4971 (N_4971,In_470,In_854);
xor U4972 (N_4972,In_1672,In_2229);
nor U4973 (N_4973,In_2898,In_2969);
xnor U4974 (N_4974,In_2248,In_2420);
and U4975 (N_4975,In_1748,In_2780);
or U4976 (N_4976,In_893,In_1787);
and U4977 (N_4977,In_1821,In_397);
nor U4978 (N_4978,In_132,In_2173);
and U4979 (N_4979,In_234,In_2461);
nor U4980 (N_4980,In_304,In_787);
nor U4981 (N_4981,In_448,In_817);
and U4982 (N_4982,In_1251,In_86);
nor U4983 (N_4983,In_1431,In_484);
or U4984 (N_4984,In_2010,In_924);
nor U4985 (N_4985,In_962,In_120);
nand U4986 (N_4986,In_762,In_1152);
nor U4987 (N_4987,In_685,In_1047);
or U4988 (N_4988,In_1726,In_401);
and U4989 (N_4989,In_2519,In_931);
or U4990 (N_4990,In_175,In_499);
nor U4991 (N_4991,In_277,In_2748);
xnor U4992 (N_4992,In_653,In_2115);
nand U4993 (N_4993,In_1971,In_2946);
nand U4994 (N_4994,In_79,In_457);
nand U4995 (N_4995,In_696,In_65);
xnor U4996 (N_4996,In_1524,In_2829);
xor U4997 (N_4997,In_2094,In_1683);
nand U4998 (N_4998,In_2358,In_127);
and U4999 (N_4999,In_1874,In_472);
xor U5000 (N_5000,In_1518,In_2689);
or U5001 (N_5001,In_1684,In_1809);
xnor U5002 (N_5002,In_607,In_850);
xnor U5003 (N_5003,In_37,In_634);
and U5004 (N_5004,In_140,In_602);
xor U5005 (N_5005,In_1043,In_1366);
xor U5006 (N_5006,In_2711,In_2678);
nor U5007 (N_5007,In_973,In_1092);
xnor U5008 (N_5008,In_1669,In_1206);
nor U5009 (N_5009,In_790,In_269);
nor U5010 (N_5010,In_97,In_810);
nor U5011 (N_5011,In_2699,In_1029);
nand U5012 (N_5012,In_1961,In_1516);
xor U5013 (N_5013,In_1285,In_1268);
and U5014 (N_5014,In_1838,In_1932);
or U5015 (N_5015,In_1850,In_873);
nand U5016 (N_5016,In_2982,In_182);
and U5017 (N_5017,In_263,In_501);
nand U5018 (N_5018,In_2607,In_583);
xnor U5019 (N_5019,In_1003,In_2701);
or U5020 (N_5020,In_2537,In_385);
nand U5021 (N_5021,In_690,In_1979);
nor U5022 (N_5022,In_2325,In_1842);
or U5023 (N_5023,In_931,In_824);
or U5024 (N_5024,In_276,In_2694);
or U5025 (N_5025,In_125,In_1473);
and U5026 (N_5026,In_915,In_2515);
or U5027 (N_5027,In_1609,In_1817);
and U5028 (N_5028,In_2430,In_1077);
xnor U5029 (N_5029,In_2353,In_1668);
and U5030 (N_5030,In_2436,In_2344);
nor U5031 (N_5031,In_429,In_662);
nand U5032 (N_5032,In_2602,In_1661);
or U5033 (N_5033,In_2318,In_2684);
and U5034 (N_5034,In_925,In_2529);
nand U5035 (N_5035,In_1014,In_2910);
and U5036 (N_5036,In_184,In_206);
or U5037 (N_5037,In_991,In_1287);
nand U5038 (N_5038,In_68,In_2255);
or U5039 (N_5039,In_637,In_1698);
nor U5040 (N_5040,In_1070,In_644);
and U5041 (N_5041,In_996,In_2864);
and U5042 (N_5042,In_1680,In_2304);
or U5043 (N_5043,In_1045,In_2387);
or U5044 (N_5044,In_166,In_1051);
or U5045 (N_5045,In_1777,In_1237);
nor U5046 (N_5046,In_2334,In_972);
or U5047 (N_5047,In_1108,In_1630);
or U5048 (N_5048,In_1336,In_1026);
nand U5049 (N_5049,In_2899,In_179);
nor U5050 (N_5050,In_1528,In_255);
nor U5051 (N_5051,In_2584,In_1675);
nor U5052 (N_5052,In_680,In_1383);
xor U5053 (N_5053,In_2293,In_2163);
or U5054 (N_5054,In_1227,In_2753);
nand U5055 (N_5055,In_2925,In_1294);
nor U5056 (N_5056,In_2350,In_2985);
or U5057 (N_5057,In_2893,In_533);
nand U5058 (N_5058,In_1898,In_535);
xnor U5059 (N_5059,In_2822,In_2687);
xnor U5060 (N_5060,In_1008,In_427);
nor U5061 (N_5061,In_2811,In_2067);
or U5062 (N_5062,In_1726,In_2278);
or U5063 (N_5063,In_2063,In_1818);
xnor U5064 (N_5064,In_1359,In_1830);
nand U5065 (N_5065,In_2261,In_2004);
xor U5066 (N_5066,In_265,In_1288);
nand U5067 (N_5067,In_1040,In_998);
nor U5068 (N_5068,In_2874,In_434);
or U5069 (N_5069,In_2129,In_1422);
xnor U5070 (N_5070,In_1818,In_579);
nor U5071 (N_5071,In_2781,In_925);
nor U5072 (N_5072,In_2769,In_2470);
or U5073 (N_5073,In_1616,In_416);
xor U5074 (N_5074,In_1928,In_1886);
and U5075 (N_5075,In_936,In_2617);
xnor U5076 (N_5076,In_1453,In_2186);
or U5077 (N_5077,In_414,In_2309);
nand U5078 (N_5078,In_2126,In_2906);
or U5079 (N_5079,In_2434,In_816);
nand U5080 (N_5080,In_2646,In_1476);
and U5081 (N_5081,In_1282,In_2127);
nand U5082 (N_5082,In_1716,In_1648);
xnor U5083 (N_5083,In_2820,In_2014);
or U5084 (N_5084,In_1633,In_1884);
and U5085 (N_5085,In_2643,In_183);
and U5086 (N_5086,In_915,In_2410);
xor U5087 (N_5087,In_1693,In_1302);
and U5088 (N_5088,In_619,In_2547);
nand U5089 (N_5089,In_2450,In_860);
xnor U5090 (N_5090,In_2488,In_1185);
nor U5091 (N_5091,In_1379,In_2999);
xor U5092 (N_5092,In_2207,In_1753);
or U5093 (N_5093,In_2930,In_2151);
nor U5094 (N_5094,In_1715,In_1989);
and U5095 (N_5095,In_1178,In_834);
xnor U5096 (N_5096,In_1860,In_2513);
or U5097 (N_5097,In_1719,In_2383);
and U5098 (N_5098,In_2448,In_1760);
nor U5099 (N_5099,In_2717,In_533);
or U5100 (N_5100,In_1117,In_2947);
nor U5101 (N_5101,In_1556,In_651);
or U5102 (N_5102,In_2032,In_781);
nand U5103 (N_5103,In_1355,In_2387);
and U5104 (N_5104,In_342,In_284);
and U5105 (N_5105,In_2317,In_2444);
or U5106 (N_5106,In_1774,In_1212);
and U5107 (N_5107,In_2397,In_2748);
nor U5108 (N_5108,In_1300,In_1005);
nor U5109 (N_5109,In_578,In_2833);
nand U5110 (N_5110,In_27,In_1571);
nand U5111 (N_5111,In_1000,In_937);
nor U5112 (N_5112,In_197,In_1448);
xor U5113 (N_5113,In_2649,In_2567);
xor U5114 (N_5114,In_400,In_2624);
xnor U5115 (N_5115,In_1642,In_1562);
and U5116 (N_5116,In_2752,In_2569);
or U5117 (N_5117,In_2783,In_1472);
xor U5118 (N_5118,In_2996,In_2551);
nand U5119 (N_5119,In_971,In_2635);
or U5120 (N_5120,In_1086,In_1253);
nor U5121 (N_5121,In_2671,In_2352);
nor U5122 (N_5122,In_337,In_1907);
nor U5123 (N_5123,In_2110,In_2185);
xor U5124 (N_5124,In_2506,In_2112);
xnor U5125 (N_5125,In_945,In_496);
xor U5126 (N_5126,In_572,In_1410);
nand U5127 (N_5127,In_1069,In_1972);
or U5128 (N_5128,In_156,In_2819);
nand U5129 (N_5129,In_1158,In_1308);
nor U5130 (N_5130,In_1699,In_2251);
nor U5131 (N_5131,In_1978,In_1485);
nand U5132 (N_5132,In_670,In_2904);
nand U5133 (N_5133,In_1703,In_2097);
or U5134 (N_5134,In_2653,In_1181);
or U5135 (N_5135,In_2134,In_1645);
nand U5136 (N_5136,In_1527,In_384);
and U5137 (N_5137,In_2592,In_2711);
and U5138 (N_5138,In_2615,In_204);
xnor U5139 (N_5139,In_2923,In_1632);
or U5140 (N_5140,In_1813,In_1052);
xnor U5141 (N_5141,In_602,In_847);
and U5142 (N_5142,In_2134,In_2299);
xor U5143 (N_5143,In_1753,In_975);
and U5144 (N_5144,In_299,In_1528);
nand U5145 (N_5145,In_1215,In_1795);
nor U5146 (N_5146,In_1928,In_2901);
nor U5147 (N_5147,In_467,In_2843);
nand U5148 (N_5148,In_1030,In_1016);
or U5149 (N_5149,In_332,In_860);
or U5150 (N_5150,In_909,In_480);
or U5151 (N_5151,In_1234,In_2480);
nor U5152 (N_5152,In_604,In_2370);
or U5153 (N_5153,In_2652,In_737);
nor U5154 (N_5154,In_2580,In_1536);
xor U5155 (N_5155,In_1340,In_365);
nand U5156 (N_5156,In_642,In_1965);
and U5157 (N_5157,In_1189,In_1766);
xnor U5158 (N_5158,In_2141,In_760);
and U5159 (N_5159,In_1968,In_289);
or U5160 (N_5160,In_1525,In_1868);
or U5161 (N_5161,In_1968,In_62);
or U5162 (N_5162,In_1144,In_1085);
nor U5163 (N_5163,In_471,In_1728);
nand U5164 (N_5164,In_427,In_466);
nand U5165 (N_5165,In_1535,In_2801);
and U5166 (N_5166,In_2725,In_974);
and U5167 (N_5167,In_2175,In_586);
nand U5168 (N_5168,In_1887,In_2586);
and U5169 (N_5169,In_1899,In_1523);
or U5170 (N_5170,In_395,In_1797);
nor U5171 (N_5171,In_760,In_2880);
and U5172 (N_5172,In_2820,In_142);
xnor U5173 (N_5173,In_2533,In_2620);
xor U5174 (N_5174,In_762,In_1859);
nand U5175 (N_5175,In_1675,In_1333);
nor U5176 (N_5176,In_1654,In_1954);
nor U5177 (N_5177,In_2977,In_1136);
and U5178 (N_5178,In_1965,In_2528);
and U5179 (N_5179,In_1008,In_1453);
xnor U5180 (N_5180,In_1253,In_2935);
nand U5181 (N_5181,In_851,In_1824);
nor U5182 (N_5182,In_1077,In_2182);
nor U5183 (N_5183,In_1301,In_64);
or U5184 (N_5184,In_81,In_2113);
nor U5185 (N_5185,In_1206,In_2710);
nand U5186 (N_5186,In_2695,In_291);
or U5187 (N_5187,In_668,In_1305);
nand U5188 (N_5188,In_1007,In_2071);
nand U5189 (N_5189,In_668,In_2412);
or U5190 (N_5190,In_1988,In_2037);
and U5191 (N_5191,In_1693,In_2233);
or U5192 (N_5192,In_1298,In_779);
and U5193 (N_5193,In_895,In_1307);
nor U5194 (N_5194,In_1901,In_2727);
or U5195 (N_5195,In_2319,In_908);
nor U5196 (N_5196,In_17,In_1142);
nor U5197 (N_5197,In_98,In_1035);
nand U5198 (N_5198,In_925,In_1951);
nor U5199 (N_5199,In_687,In_1726);
nand U5200 (N_5200,In_2680,In_2922);
or U5201 (N_5201,In_2186,In_1797);
nand U5202 (N_5202,In_609,In_2450);
xnor U5203 (N_5203,In_767,In_2073);
xor U5204 (N_5204,In_1986,In_2735);
or U5205 (N_5205,In_983,In_2606);
or U5206 (N_5206,In_2257,In_170);
nor U5207 (N_5207,In_879,In_1692);
and U5208 (N_5208,In_2411,In_635);
and U5209 (N_5209,In_2624,In_808);
xor U5210 (N_5210,In_134,In_2892);
and U5211 (N_5211,In_107,In_2722);
nand U5212 (N_5212,In_937,In_286);
nor U5213 (N_5213,In_1295,In_2298);
nand U5214 (N_5214,In_1375,In_1223);
nor U5215 (N_5215,In_1107,In_2389);
or U5216 (N_5216,In_149,In_2140);
and U5217 (N_5217,In_842,In_929);
nand U5218 (N_5218,In_2502,In_513);
or U5219 (N_5219,In_1941,In_2949);
nor U5220 (N_5220,In_816,In_2236);
and U5221 (N_5221,In_1756,In_348);
and U5222 (N_5222,In_2971,In_2446);
nor U5223 (N_5223,In_260,In_1929);
and U5224 (N_5224,In_2633,In_624);
and U5225 (N_5225,In_846,In_1665);
xor U5226 (N_5226,In_707,In_2612);
nand U5227 (N_5227,In_1095,In_969);
or U5228 (N_5228,In_8,In_1438);
nor U5229 (N_5229,In_1225,In_2646);
or U5230 (N_5230,In_220,In_872);
and U5231 (N_5231,In_1210,In_811);
nor U5232 (N_5232,In_1284,In_443);
or U5233 (N_5233,In_826,In_2636);
xor U5234 (N_5234,In_1931,In_2522);
xnor U5235 (N_5235,In_1874,In_2431);
or U5236 (N_5236,In_2826,In_2391);
nand U5237 (N_5237,In_1882,In_2040);
nor U5238 (N_5238,In_2212,In_1820);
and U5239 (N_5239,In_989,In_280);
and U5240 (N_5240,In_1501,In_563);
nand U5241 (N_5241,In_2116,In_2138);
or U5242 (N_5242,In_2539,In_35);
nand U5243 (N_5243,In_1139,In_540);
nor U5244 (N_5244,In_203,In_105);
and U5245 (N_5245,In_35,In_1926);
nand U5246 (N_5246,In_511,In_2990);
xnor U5247 (N_5247,In_2374,In_779);
nor U5248 (N_5248,In_2346,In_586);
nand U5249 (N_5249,In_2002,In_1401);
or U5250 (N_5250,In_1053,In_805);
xor U5251 (N_5251,In_1083,In_1941);
nor U5252 (N_5252,In_349,In_1115);
nand U5253 (N_5253,In_1768,In_2646);
and U5254 (N_5254,In_2986,In_684);
or U5255 (N_5255,In_2452,In_102);
and U5256 (N_5256,In_23,In_373);
nand U5257 (N_5257,In_2584,In_2860);
nor U5258 (N_5258,In_818,In_1375);
nand U5259 (N_5259,In_1816,In_1702);
and U5260 (N_5260,In_432,In_1271);
and U5261 (N_5261,In_1122,In_447);
xor U5262 (N_5262,In_2497,In_1511);
xor U5263 (N_5263,In_2515,In_1765);
xor U5264 (N_5264,In_563,In_949);
or U5265 (N_5265,In_1159,In_1050);
or U5266 (N_5266,In_2542,In_2113);
and U5267 (N_5267,In_1459,In_2361);
xnor U5268 (N_5268,In_672,In_2007);
nand U5269 (N_5269,In_2982,In_1202);
or U5270 (N_5270,In_1197,In_1894);
nand U5271 (N_5271,In_17,In_1928);
xnor U5272 (N_5272,In_1684,In_1985);
nor U5273 (N_5273,In_792,In_1927);
nor U5274 (N_5274,In_638,In_351);
or U5275 (N_5275,In_1602,In_2671);
nand U5276 (N_5276,In_1241,In_2394);
nor U5277 (N_5277,In_2556,In_1812);
xor U5278 (N_5278,In_1924,In_2841);
xor U5279 (N_5279,In_2260,In_727);
xnor U5280 (N_5280,In_2138,In_1598);
and U5281 (N_5281,In_2625,In_2676);
nor U5282 (N_5282,In_575,In_89);
nor U5283 (N_5283,In_782,In_906);
or U5284 (N_5284,In_2246,In_1763);
xnor U5285 (N_5285,In_402,In_2774);
nor U5286 (N_5286,In_985,In_2534);
or U5287 (N_5287,In_1846,In_2557);
or U5288 (N_5288,In_737,In_1541);
and U5289 (N_5289,In_1408,In_2043);
or U5290 (N_5290,In_2712,In_294);
xnor U5291 (N_5291,In_529,In_798);
or U5292 (N_5292,In_968,In_704);
or U5293 (N_5293,In_1893,In_1534);
nor U5294 (N_5294,In_1595,In_1692);
or U5295 (N_5295,In_769,In_1686);
nor U5296 (N_5296,In_96,In_1409);
and U5297 (N_5297,In_327,In_878);
nand U5298 (N_5298,In_2396,In_573);
xnor U5299 (N_5299,In_181,In_1435);
xnor U5300 (N_5300,In_2370,In_2407);
nor U5301 (N_5301,In_2939,In_936);
and U5302 (N_5302,In_824,In_245);
and U5303 (N_5303,In_2488,In_1088);
or U5304 (N_5304,In_2750,In_900);
or U5305 (N_5305,In_1072,In_544);
or U5306 (N_5306,In_1077,In_2479);
nand U5307 (N_5307,In_388,In_2101);
nand U5308 (N_5308,In_2632,In_2659);
or U5309 (N_5309,In_1654,In_2278);
nor U5310 (N_5310,In_177,In_866);
xnor U5311 (N_5311,In_2648,In_1817);
nor U5312 (N_5312,In_1640,In_396);
or U5313 (N_5313,In_2305,In_504);
and U5314 (N_5314,In_2215,In_580);
and U5315 (N_5315,In_2459,In_1841);
nand U5316 (N_5316,In_1584,In_1961);
or U5317 (N_5317,In_1469,In_2764);
nor U5318 (N_5318,In_2542,In_1037);
xnor U5319 (N_5319,In_2789,In_2377);
nand U5320 (N_5320,In_507,In_2550);
nand U5321 (N_5321,In_1773,In_1254);
nand U5322 (N_5322,In_2928,In_2250);
and U5323 (N_5323,In_2905,In_2337);
xor U5324 (N_5324,In_2222,In_2239);
xnor U5325 (N_5325,In_2164,In_2778);
xor U5326 (N_5326,In_175,In_2356);
nand U5327 (N_5327,In_698,In_155);
and U5328 (N_5328,In_0,In_1368);
xor U5329 (N_5329,In_730,In_1920);
xnor U5330 (N_5330,In_1274,In_2406);
nor U5331 (N_5331,In_1647,In_1802);
nand U5332 (N_5332,In_2781,In_139);
nor U5333 (N_5333,In_1054,In_2689);
xnor U5334 (N_5334,In_2815,In_988);
nand U5335 (N_5335,In_1093,In_1711);
and U5336 (N_5336,In_1936,In_1339);
nand U5337 (N_5337,In_2131,In_2848);
nand U5338 (N_5338,In_1370,In_1025);
or U5339 (N_5339,In_1809,In_936);
nand U5340 (N_5340,In_2453,In_309);
nor U5341 (N_5341,In_1583,In_1166);
or U5342 (N_5342,In_2204,In_2408);
nor U5343 (N_5343,In_1205,In_910);
or U5344 (N_5344,In_57,In_1401);
and U5345 (N_5345,In_2154,In_2183);
nand U5346 (N_5346,In_556,In_2582);
and U5347 (N_5347,In_2316,In_2933);
nor U5348 (N_5348,In_204,In_2997);
and U5349 (N_5349,In_65,In_1922);
and U5350 (N_5350,In_566,In_306);
nor U5351 (N_5351,In_1957,In_1996);
nor U5352 (N_5352,In_161,In_2929);
nor U5353 (N_5353,In_1121,In_1608);
xnor U5354 (N_5354,In_456,In_55);
nand U5355 (N_5355,In_71,In_1578);
or U5356 (N_5356,In_684,In_45);
and U5357 (N_5357,In_1020,In_2039);
nor U5358 (N_5358,In_320,In_1030);
xnor U5359 (N_5359,In_550,In_2957);
nand U5360 (N_5360,In_233,In_2080);
xor U5361 (N_5361,In_1684,In_99);
xnor U5362 (N_5362,In_1492,In_1465);
nor U5363 (N_5363,In_1646,In_1423);
nand U5364 (N_5364,In_1834,In_2935);
nor U5365 (N_5365,In_1413,In_2547);
xor U5366 (N_5366,In_648,In_2331);
xor U5367 (N_5367,In_2389,In_688);
nand U5368 (N_5368,In_587,In_761);
nand U5369 (N_5369,In_2170,In_2251);
nor U5370 (N_5370,In_1059,In_166);
and U5371 (N_5371,In_1963,In_845);
and U5372 (N_5372,In_2213,In_1122);
nand U5373 (N_5373,In_1723,In_2979);
and U5374 (N_5374,In_1717,In_2419);
and U5375 (N_5375,In_2745,In_1257);
nand U5376 (N_5376,In_2305,In_2539);
and U5377 (N_5377,In_2427,In_207);
nor U5378 (N_5378,In_2229,In_1469);
or U5379 (N_5379,In_1126,In_762);
and U5380 (N_5380,In_316,In_2595);
and U5381 (N_5381,In_275,In_198);
or U5382 (N_5382,In_2745,In_2530);
or U5383 (N_5383,In_2461,In_1472);
or U5384 (N_5384,In_2985,In_721);
or U5385 (N_5385,In_1726,In_1229);
or U5386 (N_5386,In_2432,In_2701);
and U5387 (N_5387,In_2230,In_2916);
and U5388 (N_5388,In_597,In_723);
nor U5389 (N_5389,In_905,In_368);
xnor U5390 (N_5390,In_1897,In_881);
xor U5391 (N_5391,In_2672,In_1733);
and U5392 (N_5392,In_1372,In_1631);
and U5393 (N_5393,In_2734,In_2223);
and U5394 (N_5394,In_2052,In_1123);
and U5395 (N_5395,In_115,In_1367);
xnor U5396 (N_5396,In_2078,In_2845);
and U5397 (N_5397,In_1270,In_1356);
or U5398 (N_5398,In_2161,In_2020);
nand U5399 (N_5399,In_2462,In_1291);
xor U5400 (N_5400,In_1373,In_1060);
or U5401 (N_5401,In_2883,In_2271);
or U5402 (N_5402,In_2889,In_2630);
nor U5403 (N_5403,In_2967,In_60);
nor U5404 (N_5404,In_9,In_2184);
nand U5405 (N_5405,In_2012,In_2054);
and U5406 (N_5406,In_2215,In_2995);
xor U5407 (N_5407,In_1747,In_2690);
nand U5408 (N_5408,In_1833,In_1376);
nand U5409 (N_5409,In_378,In_1849);
or U5410 (N_5410,In_1569,In_2223);
and U5411 (N_5411,In_1394,In_457);
nor U5412 (N_5412,In_1328,In_44);
xor U5413 (N_5413,In_1174,In_659);
nand U5414 (N_5414,In_617,In_2036);
and U5415 (N_5415,In_1622,In_588);
nand U5416 (N_5416,In_224,In_2216);
xor U5417 (N_5417,In_671,In_1400);
nand U5418 (N_5418,In_552,In_296);
nand U5419 (N_5419,In_2605,In_1657);
or U5420 (N_5420,In_2785,In_531);
nand U5421 (N_5421,In_2674,In_1483);
or U5422 (N_5422,In_2689,In_853);
nand U5423 (N_5423,In_899,In_170);
xnor U5424 (N_5424,In_106,In_2869);
or U5425 (N_5425,In_166,In_2555);
xnor U5426 (N_5426,In_2017,In_1820);
xor U5427 (N_5427,In_168,In_1642);
or U5428 (N_5428,In_2689,In_2600);
nand U5429 (N_5429,In_1929,In_2205);
xnor U5430 (N_5430,In_1148,In_2215);
or U5431 (N_5431,In_690,In_962);
and U5432 (N_5432,In_225,In_1108);
and U5433 (N_5433,In_2839,In_2557);
nand U5434 (N_5434,In_2437,In_2040);
nand U5435 (N_5435,In_2905,In_1202);
nand U5436 (N_5436,In_1726,In_2205);
or U5437 (N_5437,In_2102,In_407);
nand U5438 (N_5438,In_2600,In_2086);
xnor U5439 (N_5439,In_2308,In_1618);
nand U5440 (N_5440,In_2149,In_477);
and U5441 (N_5441,In_1851,In_2847);
nand U5442 (N_5442,In_849,In_1103);
and U5443 (N_5443,In_1491,In_751);
or U5444 (N_5444,In_2752,In_2547);
nand U5445 (N_5445,In_1618,In_2194);
and U5446 (N_5446,In_716,In_2105);
or U5447 (N_5447,In_672,In_2824);
and U5448 (N_5448,In_1229,In_683);
nor U5449 (N_5449,In_2414,In_1136);
xnor U5450 (N_5450,In_1232,In_2185);
nand U5451 (N_5451,In_1412,In_562);
or U5452 (N_5452,In_1083,In_880);
nand U5453 (N_5453,In_2995,In_31);
or U5454 (N_5454,In_1501,In_1744);
nand U5455 (N_5455,In_1931,In_595);
nor U5456 (N_5456,In_582,In_1204);
nor U5457 (N_5457,In_974,In_486);
xnor U5458 (N_5458,In_1185,In_1334);
nand U5459 (N_5459,In_297,In_1026);
and U5460 (N_5460,In_2602,In_2955);
nand U5461 (N_5461,In_1129,In_1897);
and U5462 (N_5462,In_608,In_2677);
or U5463 (N_5463,In_1835,In_737);
nand U5464 (N_5464,In_1094,In_2166);
xnor U5465 (N_5465,In_803,In_2603);
nor U5466 (N_5466,In_2787,In_1813);
and U5467 (N_5467,In_2213,In_349);
xor U5468 (N_5468,In_1265,In_1089);
or U5469 (N_5469,In_1757,In_2559);
and U5470 (N_5470,In_1114,In_1640);
xor U5471 (N_5471,In_2230,In_230);
nor U5472 (N_5472,In_2208,In_1457);
nand U5473 (N_5473,In_2504,In_952);
nor U5474 (N_5474,In_598,In_128);
and U5475 (N_5475,In_2246,In_709);
xnor U5476 (N_5476,In_2598,In_1267);
nand U5477 (N_5477,In_401,In_2216);
and U5478 (N_5478,In_1138,In_2407);
or U5479 (N_5479,In_388,In_1743);
nand U5480 (N_5480,In_1633,In_2810);
nand U5481 (N_5481,In_1709,In_1097);
nor U5482 (N_5482,In_1779,In_186);
and U5483 (N_5483,In_1419,In_183);
and U5484 (N_5484,In_2275,In_2116);
nand U5485 (N_5485,In_1385,In_2910);
nor U5486 (N_5486,In_1340,In_2053);
nor U5487 (N_5487,In_1890,In_1256);
nor U5488 (N_5488,In_1713,In_2728);
nand U5489 (N_5489,In_1587,In_630);
nor U5490 (N_5490,In_22,In_203);
or U5491 (N_5491,In_1137,In_271);
nor U5492 (N_5492,In_2878,In_2916);
and U5493 (N_5493,In_1258,In_627);
nor U5494 (N_5494,In_2227,In_1578);
or U5495 (N_5495,In_1181,In_1365);
or U5496 (N_5496,In_1840,In_2624);
nand U5497 (N_5497,In_10,In_105);
xor U5498 (N_5498,In_320,In_709);
nand U5499 (N_5499,In_496,In_1912);
nand U5500 (N_5500,In_2718,In_38);
nand U5501 (N_5501,In_1001,In_2455);
nand U5502 (N_5502,In_156,In_2421);
or U5503 (N_5503,In_1738,In_1075);
xnor U5504 (N_5504,In_1571,In_780);
xor U5505 (N_5505,In_1699,In_2066);
and U5506 (N_5506,In_515,In_1399);
and U5507 (N_5507,In_2189,In_1125);
nand U5508 (N_5508,In_920,In_646);
nand U5509 (N_5509,In_2888,In_1220);
and U5510 (N_5510,In_1066,In_1773);
xor U5511 (N_5511,In_100,In_2027);
and U5512 (N_5512,In_343,In_116);
or U5513 (N_5513,In_923,In_715);
or U5514 (N_5514,In_163,In_2810);
nand U5515 (N_5515,In_1132,In_2496);
nor U5516 (N_5516,In_366,In_1761);
or U5517 (N_5517,In_2460,In_2833);
xnor U5518 (N_5518,In_2239,In_2218);
nor U5519 (N_5519,In_1273,In_2204);
or U5520 (N_5520,In_185,In_223);
nor U5521 (N_5521,In_816,In_1027);
nand U5522 (N_5522,In_1631,In_2632);
or U5523 (N_5523,In_2874,In_2706);
nand U5524 (N_5524,In_797,In_1889);
nor U5525 (N_5525,In_398,In_2459);
or U5526 (N_5526,In_1969,In_2236);
and U5527 (N_5527,In_1626,In_1095);
nor U5528 (N_5528,In_481,In_1376);
nor U5529 (N_5529,In_195,In_2005);
or U5530 (N_5530,In_621,In_1929);
or U5531 (N_5531,In_555,In_2268);
nand U5532 (N_5532,In_2657,In_2362);
and U5533 (N_5533,In_1327,In_1606);
nor U5534 (N_5534,In_2054,In_1489);
or U5535 (N_5535,In_1823,In_2256);
or U5536 (N_5536,In_1411,In_1898);
or U5537 (N_5537,In_2370,In_1739);
or U5538 (N_5538,In_14,In_2491);
nand U5539 (N_5539,In_2805,In_409);
nand U5540 (N_5540,In_766,In_711);
nand U5541 (N_5541,In_254,In_2234);
xnor U5542 (N_5542,In_207,In_1917);
xor U5543 (N_5543,In_594,In_1851);
nor U5544 (N_5544,In_1399,In_2783);
or U5545 (N_5545,In_2744,In_513);
or U5546 (N_5546,In_2660,In_2207);
or U5547 (N_5547,In_1791,In_2290);
nor U5548 (N_5548,In_86,In_1609);
or U5549 (N_5549,In_2923,In_1956);
nor U5550 (N_5550,In_1359,In_69);
xor U5551 (N_5551,In_375,In_2934);
xor U5552 (N_5552,In_509,In_1701);
and U5553 (N_5553,In_2462,In_2106);
or U5554 (N_5554,In_1039,In_2879);
nor U5555 (N_5555,In_1478,In_2065);
nor U5556 (N_5556,In_1232,In_2494);
nor U5557 (N_5557,In_349,In_223);
xor U5558 (N_5558,In_122,In_126);
xor U5559 (N_5559,In_701,In_2121);
and U5560 (N_5560,In_299,In_2799);
nand U5561 (N_5561,In_691,In_689);
or U5562 (N_5562,In_2519,In_2832);
nand U5563 (N_5563,In_83,In_2899);
nor U5564 (N_5564,In_2448,In_1012);
and U5565 (N_5565,In_1453,In_86);
nor U5566 (N_5566,In_2174,In_1392);
nor U5567 (N_5567,In_529,In_1596);
or U5568 (N_5568,In_2479,In_1632);
nand U5569 (N_5569,In_429,In_261);
nand U5570 (N_5570,In_2210,In_156);
or U5571 (N_5571,In_2104,In_1720);
nand U5572 (N_5572,In_1330,In_1468);
or U5573 (N_5573,In_2325,In_1561);
nor U5574 (N_5574,In_2871,In_487);
or U5575 (N_5575,In_2240,In_1520);
nor U5576 (N_5576,In_1793,In_1339);
and U5577 (N_5577,In_875,In_916);
nor U5578 (N_5578,In_990,In_2190);
xor U5579 (N_5579,In_1780,In_869);
nor U5580 (N_5580,In_312,In_456);
nand U5581 (N_5581,In_2655,In_1744);
xnor U5582 (N_5582,In_1822,In_1985);
and U5583 (N_5583,In_2384,In_2778);
nand U5584 (N_5584,In_837,In_1447);
nor U5585 (N_5585,In_1005,In_2626);
or U5586 (N_5586,In_845,In_927);
and U5587 (N_5587,In_733,In_1807);
or U5588 (N_5588,In_2987,In_335);
xor U5589 (N_5589,In_2402,In_634);
nand U5590 (N_5590,In_928,In_953);
xnor U5591 (N_5591,In_81,In_1692);
nand U5592 (N_5592,In_536,In_1083);
xnor U5593 (N_5593,In_1472,In_961);
or U5594 (N_5594,In_1588,In_2452);
nor U5595 (N_5595,In_2570,In_1349);
or U5596 (N_5596,In_2725,In_1823);
or U5597 (N_5597,In_606,In_2613);
xnor U5598 (N_5598,In_1903,In_1408);
xor U5599 (N_5599,In_1747,In_1594);
nand U5600 (N_5600,In_2399,In_2515);
and U5601 (N_5601,In_2755,In_1862);
or U5602 (N_5602,In_1994,In_195);
nor U5603 (N_5603,In_2772,In_2465);
and U5604 (N_5604,In_2679,In_2298);
and U5605 (N_5605,In_91,In_1049);
and U5606 (N_5606,In_1063,In_62);
nand U5607 (N_5607,In_1529,In_676);
and U5608 (N_5608,In_2878,In_46);
nor U5609 (N_5609,In_2501,In_1499);
and U5610 (N_5610,In_1916,In_72);
nand U5611 (N_5611,In_1070,In_2770);
and U5612 (N_5612,In_458,In_291);
xor U5613 (N_5613,In_237,In_2760);
xnor U5614 (N_5614,In_1638,In_782);
nor U5615 (N_5615,In_548,In_2483);
or U5616 (N_5616,In_1626,In_859);
nand U5617 (N_5617,In_496,In_1385);
nor U5618 (N_5618,In_1611,In_647);
and U5619 (N_5619,In_769,In_1828);
xnor U5620 (N_5620,In_2892,In_2526);
nand U5621 (N_5621,In_93,In_410);
nor U5622 (N_5622,In_1652,In_41);
or U5623 (N_5623,In_1370,In_1206);
xor U5624 (N_5624,In_2473,In_70);
or U5625 (N_5625,In_1617,In_2168);
nand U5626 (N_5626,In_1454,In_974);
xor U5627 (N_5627,In_1608,In_1569);
nor U5628 (N_5628,In_346,In_1488);
and U5629 (N_5629,In_357,In_1961);
or U5630 (N_5630,In_1673,In_988);
nand U5631 (N_5631,In_1832,In_223);
or U5632 (N_5632,In_357,In_2905);
and U5633 (N_5633,In_2783,In_1148);
nor U5634 (N_5634,In_2026,In_1173);
nor U5635 (N_5635,In_1966,In_2876);
or U5636 (N_5636,In_2186,In_2245);
nor U5637 (N_5637,In_327,In_231);
or U5638 (N_5638,In_328,In_479);
and U5639 (N_5639,In_2532,In_1842);
xor U5640 (N_5640,In_1510,In_1616);
or U5641 (N_5641,In_1850,In_2952);
and U5642 (N_5642,In_1613,In_2600);
nor U5643 (N_5643,In_382,In_1332);
and U5644 (N_5644,In_127,In_2805);
nand U5645 (N_5645,In_207,In_2211);
xnor U5646 (N_5646,In_2269,In_2001);
nor U5647 (N_5647,In_2031,In_1722);
nand U5648 (N_5648,In_1308,In_2794);
xor U5649 (N_5649,In_301,In_2334);
nor U5650 (N_5650,In_945,In_2580);
nor U5651 (N_5651,In_1414,In_290);
nand U5652 (N_5652,In_2221,In_2262);
nand U5653 (N_5653,In_2893,In_957);
nand U5654 (N_5654,In_2040,In_854);
and U5655 (N_5655,In_1627,In_1861);
nand U5656 (N_5656,In_1104,In_1500);
nor U5657 (N_5657,In_2772,In_1791);
nand U5658 (N_5658,In_2462,In_2439);
and U5659 (N_5659,In_731,In_233);
nand U5660 (N_5660,In_1090,In_1842);
nor U5661 (N_5661,In_1902,In_2084);
or U5662 (N_5662,In_1303,In_2657);
and U5663 (N_5663,In_1504,In_2731);
and U5664 (N_5664,In_851,In_2442);
nand U5665 (N_5665,In_2819,In_856);
xnor U5666 (N_5666,In_2132,In_633);
and U5667 (N_5667,In_700,In_2631);
nand U5668 (N_5668,In_2610,In_2206);
and U5669 (N_5669,In_879,In_653);
and U5670 (N_5670,In_1414,In_2655);
xor U5671 (N_5671,In_2348,In_306);
nor U5672 (N_5672,In_2517,In_1063);
nor U5673 (N_5673,In_1625,In_1279);
nor U5674 (N_5674,In_1980,In_209);
nand U5675 (N_5675,In_2872,In_262);
nor U5676 (N_5676,In_2463,In_1261);
and U5677 (N_5677,In_2406,In_209);
nor U5678 (N_5678,In_2933,In_2192);
or U5679 (N_5679,In_938,In_2186);
nor U5680 (N_5680,In_1136,In_631);
or U5681 (N_5681,In_2394,In_1392);
nand U5682 (N_5682,In_1751,In_2347);
and U5683 (N_5683,In_987,In_1765);
and U5684 (N_5684,In_1285,In_155);
nand U5685 (N_5685,In_2313,In_2078);
nor U5686 (N_5686,In_2898,In_2942);
xnor U5687 (N_5687,In_899,In_2002);
nor U5688 (N_5688,In_1528,In_1789);
and U5689 (N_5689,In_1458,In_391);
nand U5690 (N_5690,In_1001,In_2332);
xor U5691 (N_5691,In_484,In_2461);
xor U5692 (N_5692,In_764,In_1540);
nor U5693 (N_5693,In_52,In_2022);
nand U5694 (N_5694,In_1890,In_892);
nor U5695 (N_5695,In_394,In_1377);
nand U5696 (N_5696,In_2465,In_419);
and U5697 (N_5697,In_972,In_927);
and U5698 (N_5698,In_1273,In_708);
nand U5699 (N_5699,In_1918,In_2186);
nor U5700 (N_5700,In_2962,In_781);
and U5701 (N_5701,In_1863,In_32);
and U5702 (N_5702,In_1960,In_1390);
nand U5703 (N_5703,In_2953,In_2163);
and U5704 (N_5704,In_149,In_1253);
nand U5705 (N_5705,In_2244,In_1216);
or U5706 (N_5706,In_1687,In_2457);
xor U5707 (N_5707,In_69,In_134);
nor U5708 (N_5708,In_219,In_2922);
nand U5709 (N_5709,In_440,In_2409);
or U5710 (N_5710,In_552,In_947);
and U5711 (N_5711,In_201,In_1595);
nand U5712 (N_5712,In_2719,In_1958);
nor U5713 (N_5713,In_2132,In_996);
nand U5714 (N_5714,In_2551,In_948);
nor U5715 (N_5715,In_2886,In_2874);
xnor U5716 (N_5716,In_9,In_793);
nand U5717 (N_5717,In_793,In_149);
or U5718 (N_5718,In_1571,In_608);
xnor U5719 (N_5719,In_810,In_2808);
nand U5720 (N_5720,In_27,In_524);
nand U5721 (N_5721,In_2106,In_1192);
nand U5722 (N_5722,In_1531,In_1202);
or U5723 (N_5723,In_140,In_1137);
xor U5724 (N_5724,In_509,In_142);
nor U5725 (N_5725,In_2602,In_547);
and U5726 (N_5726,In_2186,In_2182);
nand U5727 (N_5727,In_1910,In_1392);
and U5728 (N_5728,In_696,In_2984);
xor U5729 (N_5729,In_2128,In_2580);
nor U5730 (N_5730,In_1554,In_903);
xnor U5731 (N_5731,In_786,In_1892);
xnor U5732 (N_5732,In_524,In_51);
xnor U5733 (N_5733,In_1450,In_2583);
and U5734 (N_5734,In_2754,In_2788);
xor U5735 (N_5735,In_2846,In_1699);
or U5736 (N_5736,In_419,In_498);
nand U5737 (N_5737,In_1348,In_2150);
and U5738 (N_5738,In_1613,In_1832);
and U5739 (N_5739,In_1952,In_2717);
xor U5740 (N_5740,In_314,In_1543);
or U5741 (N_5741,In_2068,In_177);
xor U5742 (N_5742,In_1882,In_100);
and U5743 (N_5743,In_2580,In_1081);
nand U5744 (N_5744,In_843,In_1036);
and U5745 (N_5745,In_1956,In_2726);
or U5746 (N_5746,In_1189,In_311);
and U5747 (N_5747,In_2951,In_1784);
xor U5748 (N_5748,In_2232,In_1886);
nor U5749 (N_5749,In_1419,In_2160);
or U5750 (N_5750,In_1110,In_641);
and U5751 (N_5751,In_598,In_2975);
nor U5752 (N_5752,In_2656,In_803);
xnor U5753 (N_5753,In_181,In_64);
nand U5754 (N_5754,In_2905,In_2518);
xnor U5755 (N_5755,In_8,In_1921);
nand U5756 (N_5756,In_2418,In_1916);
nand U5757 (N_5757,In_183,In_2281);
nor U5758 (N_5758,In_179,In_2536);
nor U5759 (N_5759,In_304,In_844);
and U5760 (N_5760,In_730,In_278);
nand U5761 (N_5761,In_1265,In_2041);
xnor U5762 (N_5762,In_570,In_750);
nor U5763 (N_5763,In_2054,In_2422);
nand U5764 (N_5764,In_2491,In_2405);
xor U5765 (N_5765,In_2293,In_1959);
or U5766 (N_5766,In_1860,In_891);
xnor U5767 (N_5767,In_1417,In_1583);
nor U5768 (N_5768,In_958,In_868);
nor U5769 (N_5769,In_829,In_2061);
nor U5770 (N_5770,In_1439,In_2827);
xnor U5771 (N_5771,In_1954,In_1562);
nand U5772 (N_5772,In_1864,In_2519);
or U5773 (N_5773,In_708,In_1496);
nand U5774 (N_5774,In_1012,In_2504);
nor U5775 (N_5775,In_2323,In_1245);
or U5776 (N_5776,In_310,In_1550);
and U5777 (N_5777,In_1469,In_1002);
and U5778 (N_5778,In_1687,In_418);
and U5779 (N_5779,In_961,In_1328);
or U5780 (N_5780,In_2759,In_2156);
or U5781 (N_5781,In_1653,In_729);
nor U5782 (N_5782,In_900,In_2472);
or U5783 (N_5783,In_2008,In_1469);
nor U5784 (N_5784,In_1733,In_1494);
and U5785 (N_5785,In_575,In_1422);
nand U5786 (N_5786,In_125,In_2924);
or U5787 (N_5787,In_823,In_1871);
or U5788 (N_5788,In_74,In_915);
nand U5789 (N_5789,In_487,In_2587);
or U5790 (N_5790,In_446,In_1108);
xnor U5791 (N_5791,In_1077,In_2353);
and U5792 (N_5792,In_1249,In_2275);
and U5793 (N_5793,In_1774,In_479);
or U5794 (N_5794,In_1067,In_1191);
and U5795 (N_5795,In_1219,In_1657);
xor U5796 (N_5796,In_2265,In_2183);
or U5797 (N_5797,In_156,In_669);
nand U5798 (N_5798,In_838,In_365);
or U5799 (N_5799,In_2288,In_2491);
or U5800 (N_5800,In_2038,In_790);
nand U5801 (N_5801,In_488,In_1790);
nand U5802 (N_5802,In_2361,In_2704);
xnor U5803 (N_5803,In_1374,In_2017);
nor U5804 (N_5804,In_131,In_2247);
nor U5805 (N_5805,In_1422,In_1369);
xor U5806 (N_5806,In_1636,In_2478);
and U5807 (N_5807,In_1574,In_923);
nor U5808 (N_5808,In_917,In_2182);
or U5809 (N_5809,In_507,In_765);
and U5810 (N_5810,In_2348,In_1301);
nor U5811 (N_5811,In_2010,In_746);
and U5812 (N_5812,In_2697,In_2413);
nand U5813 (N_5813,In_384,In_524);
or U5814 (N_5814,In_1575,In_2505);
and U5815 (N_5815,In_531,In_2654);
or U5816 (N_5816,In_1675,In_2872);
or U5817 (N_5817,In_339,In_249);
xnor U5818 (N_5818,In_1377,In_1796);
or U5819 (N_5819,In_1158,In_731);
or U5820 (N_5820,In_2346,In_2140);
and U5821 (N_5821,In_2957,In_2780);
xor U5822 (N_5822,In_1448,In_2826);
nor U5823 (N_5823,In_1562,In_1341);
or U5824 (N_5824,In_2347,In_2938);
or U5825 (N_5825,In_1541,In_1379);
or U5826 (N_5826,In_189,In_1965);
nand U5827 (N_5827,In_2561,In_882);
or U5828 (N_5828,In_1004,In_2691);
nor U5829 (N_5829,In_1219,In_2967);
nor U5830 (N_5830,In_2134,In_856);
or U5831 (N_5831,In_2501,In_921);
nor U5832 (N_5832,In_623,In_667);
nand U5833 (N_5833,In_2392,In_640);
or U5834 (N_5834,In_1498,In_2992);
and U5835 (N_5835,In_2503,In_303);
or U5836 (N_5836,In_165,In_503);
or U5837 (N_5837,In_2704,In_1565);
or U5838 (N_5838,In_560,In_994);
or U5839 (N_5839,In_96,In_407);
nand U5840 (N_5840,In_2,In_312);
nand U5841 (N_5841,In_1140,In_853);
nor U5842 (N_5842,In_2976,In_1563);
nor U5843 (N_5843,In_2446,In_1094);
and U5844 (N_5844,In_2422,In_183);
nor U5845 (N_5845,In_1240,In_2388);
and U5846 (N_5846,In_32,In_2282);
or U5847 (N_5847,In_2329,In_2317);
nand U5848 (N_5848,In_2881,In_2983);
xnor U5849 (N_5849,In_464,In_1903);
nand U5850 (N_5850,In_2977,In_911);
nor U5851 (N_5851,In_675,In_406);
and U5852 (N_5852,In_763,In_1182);
xor U5853 (N_5853,In_1771,In_2658);
or U5854 (N_5854,In_262,In_2431);
nor U5855 (N_5855,In_1112,In_1409);
xnor U5856 (N_5856,In_776,In_1737);
xnor U5857 (N_5857,In_1713,In_1817);
nand U5858 (N_5858,In_667,In_2024);
and U5859 (N_5859,In_2999,In_1617);
and U5860 (N_5860,In_1039,In_151);
and U5861 (N_5861,In_2199,In_965);
xnor U5862 (N_5862,In_733,In_576);
nor U5863 (N_5863,In_1040,In_1910);
nand U5864 (N_5864,In_1184,In_1111);
nor U5865 (N_5865,In_895,In_440);
nand U5866 (N_5866,In_2579,In_2399);
or U5867 (N_5867,In_2444,In_1476);
nand U5868 (N_5868,In_2668,In_1956);
xor U5869 (N_5869,In_953,In_2057);
nand U5870 (N_5870,In_569,In_1078);
nor U5871 (N_5871,In_2042,In_1694);
nand U5872 (N_5872,In_1931,In_2961);
xnor U5873 (N_5873,In_1679,In_1926);
xnor U5874 (N_5874,In_1480,In_2547);
nor U5875 (N_5875,In_1217,In_751);
nand U5876 (N_5876,In_754,In_2836);
nand U5877 (N_5877,In_2121,In_756);
or U5878 (N_5878,In_1900,In_1636);
nand U5879 (N_5879,In_2870,In_1208);
and U5880 (N_5880,In_963,In_2842);
nand U5881 (N_5881,In_1482,In_2971);
nor U5882 (N_5882,In_2354,In_1559);
nand U5883 (N_5883,In_2402,In_1270);
xnor U5884 (N_5884,In_976,In_2213);
nor U5885 (N_5885,In_1653,In_592);
or U5886 (N_5886,In_937,In_2657);
nor U5887 (N_5887,In_2883,In_2287);
xor U5888 (N_5888,In_1833,In_280);
xor U5889 (N_5889,In_997,In_1947);
nand U5890 (N_5890,In_2407,In_1274);
xor U5891 (N_5891,In_275,In_1779);
and U5892 (N_5892,In_863,In_1540);
nand U5893 (N_5893,In_685,In_1303);
and U5894 (N_5894,In_2304,In_2444);
xor U5895 (N_5895,In_797,In_1465);
xor U5896 (N_5896,In_1354,In_894);
or U5897 (N_5897,In_2125,In_643);
nand U5898 (N_5898,In_1207,In_1156);
or U5899 (N_5899,In_1218,In_2940);
xor U5900 (N_5900,In_1586,In_2084);
or U5901 (N_5901,In_133,In_1152);
xor U5902 (N_5902,In_2247,In_556);
nand U5903 (N_5903,In_798,In_183);
nor U5904 (N_5904,In_2154,In_1105);
or U5905 (N_5905,In_850,In_1768);
nor U5906 (N_5906,In_1118,In_1055);
xnor U5907 (N_5907,In_184,In_721);
or U5908 (N_5908,In_1716,In_1872);
and U5909 (N_5909,In_170,In_1288);
and U5910 (N_5910,In_2988,In_2163);
nor U5911 (N_5911,In_1523,In_2994);
nor U5912 (N_5912,In_261,In_284);
nand U5913 (N_5913,In_2538,In_784);
and U5914 (N_5914,In_2604,In_2072);
or U5915 (N_5915,In_1432,In_671);
and U5916 (N_5916,In_2088,In_604);
nor U5917 (N_5917,In_918,In_1443);
nor U5918 (N_5918,In_392,In_785);
and U5919 (N_5919,In_1028,In_2041);
and U5920 (N_5920,In_2315,In_1516);
nand U5921 (N_5921,In_367,In_1651);
xor U5922 (N_5922,In_2716,In_313);
nand U5923 (N_5923,In_2321,In_1756);
xor U5924 (N_5924,In_2566,In_480);
nor U5925 (N_5925,In_1400,In_1447);
nor U5926 (N_5926,In_2176,In_2663);
nand U5927 (N_5927,In_2120,In_1419);
xnor U5928 (N_5928,In_2792,In_1432);
nand U5929 (N_5929,In_1513,In_498);
nand U5930 (N_5930,In_2984,In_1334);
or U5931 (N_5931,In_812,In_957);
xnor U5932 (N_5932,In_2691,In_976);
and U5933 (N_5933,In_2828,In_197);
nand U5934 (N_5934,In_2525,In_2038);
nor U5935 (N_5935,In_2757,In_2131);
nand U5936 (N_5936,In_544,In_2377);
xnor U5937 (N_5937,In_1210,In_1769);
xnor U5938 (N_5938,In_1541,In_904);
nand U5939 (N_5939,In_2904,In_598);
nand U5940 (N_5940,In_2432,In_1483);
xnor U5941 (N_5941,In_470,In_180);
nor U5942 (N_5942,In_194,In_1022);
or U5943 (N_5943,In_353,In_2211);
nor U5944 (N_5944,In_1796,In_1013);
xor U5945 (N_5945,In_527,In_1513);
xnor U5946 (N_5946,In_1677,In_387);
xor U5947 (N_5947,In_1534,In_37);
and U5948 (N_5948,In_2832,In_2075);
nor U5949 (N_5949,In_898,In_572);
and U5950 (N_5950,In_188,In_2837);
xnor U5951 (N_5951,In_1124,In_1789);
and U5952 (N_5952,In_1259,In_1123);
or U5953 (N_5953,In_2678,In_2259);
or U5954 (N_5954,In_1432,In_2904);
and U5955 (N_5955,In_556,In_1997);
nor U5956 (N_5956,In_1377,In_1682);
nor U5957 (N_5957,In_1105,In_2957);
and U5958 (N_5958,In_236,In_1396);
nand U5959 (N_5959,In_547,In_2282);
nand U5960 (N_5960,In_2185,In_1388);
xor U5961 (N_5961,In_0,In_998);
or U5962 (N_5962,In_727,In_318);
xnor U5963 (N_5963,In_1985,In_1276);
xor U5964 (N_5964,In_2295,In_807);
nor U5965 (N_5965,In_1462,In_1371);
nand U5966 (N_5966,In_1266,In_2131);
nand U5967 (N_5967,In_646,In_1820);
nand U5968 (N_5968,In_668,In_510);
or U5969 (N_5969,In_1241,In_492);
xnor U5970 (N_5970,In_1855,In_641);
nand U5971 (N_5971,In_1562,In_2376);
xor U5972 (N_5972,In_1795,In_2459);
nor U5973 (N_5973,In_741,In_2733);
or U5974 (N_5974,In_944,In_2585);
nand U5975 (N_5975,In_1620,In_609);
and U5976 (N_5976,In_2031,In_830);
nor U5977 (N_5977,In_2107,In_2117);
nor U5978 (N_5978,In_2826,In_2208);
and U5979 (N_5979,In_2987,In_276);
and U5980 (N_5980,In_1823,In_2783);
or U5981 (N_5981,In_2117,In_64);
nor U5982 (N_5982,In_2633,In_1911);
xnor U5983 (N_5983,In_1878,In_2033);
xor U5984 (N_5984,In_1194,In_1156);
and U5985 (N_5985,In_2132,In_2309);
nor U5986 (N_5986,In_379,In_2178);
xnor U5987 (N_5987,In_2081,In_261);
or U5988 (N_5988,In_259,In_1565);
and U5989 (N_5989,In_2115,In_922);
and U5990 (N_5990,In_1785,In_2624);
xor U5991 (N_5991,In_585,In_1081);
and U5992 (N_5992,In_820,In_2819);
nand U5993 (N_5993,In_2806,In_2339);
and U5994 (N_5994,In_2537,In_228);
nand U5995 (N_5995,In_2116,In_605);
nand U5996 (N_5996,In_2716,In_1353);
xnor U5997 (N_5997,In_1064,In_69);
xor U5998 (N_5998,In_1788,In_1676);
and U5999 (N_5999,In_1361,In_930);
or U6000 (N_6000,N_3784,N_5477);
nor U6001 (N_6001,N_4998,N_3235);
and U6002 (N_6002,N_2494,N_5341);
or U6003 (N_6003,N_4127,N_3881);
xnor U6004 (N_6004,N_5597,N_5018);
or U6005 (N_6005,N_5628,N_3735);
and U6006 (N_6006,N_2049,N_2852);
or U6007 (N_6007,N_2511,N_2869);
xor U6008 (N_6008,N_5366,N_2155);
nor U6009 (N_6009,N_479,N_1842);
and U6010 (N_6010,N_4987,N_129);
nor U6011 (N_6011,N_4577,N_4593);
and U6012 (N_6012,N_554,N_672);
or U6013 (N_6013,N_5204,N_4483);
nand U6014 (N_6014,N_3211,N_4782);
nand U6015 (N_6015,N_4451,N_4909);
and U6016 (N_6016,N_2096,N_2676);
nor U6017 (N_6017,N_3236,N_1235);
nor U6018 (N_6018,N_1815,N_5070);
xnor U6019 (N_6019,N_2350,N_4213);
or U6020 (N_6020,N_1155,N_4729);
nor U6021 (N_6021,N_5337,N_1994);
xor U6022 (N_6022,N_5787,N_3829);
or U6023 (N_6023,N_3821,N_2132);
nand U6024 (N_6024,N_1531,N_1095);
or U6025 (N_6025,N_2481,N_1303);
xnor U6026 (N_6026,N_3799,N_1808);
nand U6027 (N_6027,N_1395,N_2864);
and U6028 (N_6028,N_900,N_3149);
and U6029 (N_6029,N_5472,N_1783);
or U6030 (N_6030,N_2865,N_5722);
nand U6031 (N_6031,N_70,N_3162);
or U6032 (N_6032,N_2754,N_1335);
xor U6033 (N_6033,N_1311,N_2739);
and U6034 (N_6034,N_3645,N_1968);
xor U6035 (N_6035,N_4529,N_3197);
or U6036 (N_6036,N_4034,N_3261);
and U6037 (N_6037,N_3414,N_1242);
nor U6038 (N_6038,N_2342,N_855);
nor U6039 (N_6039,N_4765,N_978);
nor U6040 (N_6040,N_1717,N_3516);
xnor U6041 (N_6041,N_861,N_754);
nand U6042 (N_6042,N_132,N_2745);
xnor U6043 (N_6043,N_2290,N_215);
nand U6044 (N_6044,N_1091,N_1868);
nand U6045 (N_6045,N_5620,N_1374);
nor U6046 (N_6046,N_5621,N_4573);
nor U6047 (N_6047,N_5563,N_190);
xnor U6048 (N_6048,N_2164,N_4221);
nor U6049 (N_6049,N_1066,N_113);
nor U6050 (N_6050,N_932,N_2982);
nor U6051 (N_6051,N_2561,N_4931);
xnor U6052 (N_6052,N_5413,N_366);
and U6053 (N_6053,N_3114,N_5290);
nand U6054 (N_6054,N_4315,N_57);
or U6055 (N_6055,N_2202,N_714);
and U6056 (N_6056,N_857,N_5524);
xnor U6057 (N_6057,N_95,N_5172);
and U6058 (N_6058,N_3520,N_2592);
nor U6059 (N_6059,N_5903,N_4245);
or U6060 (N_6060,N_3783,N_363);
xor U6061 (N_6061,N_2986,N_3122);
and U6062 (N_6062,N_5139,N_2156);
nand U6063 (N_6063,N_2875,N_3900);
xor U6064 (N_6064,N_3756,N_5004);
xnor U6065 (N_6065,N_4712,N_5704);
or U6066 (N_6066,N_1900,N_4328);
nor U6067 (N_6067,N_4912,N_3101);
nor U6068 (N_6068,N_5896,N_5325);
nor U6069 (N_6069,N_4187,N_3800);
and U6070 (N_6070,N_3708,N_1003);
nand U6071 (N_6071,N_2229,N_5520);
xor U6072 (N_6072,N_5774,N_1317);
nor U6073 (N_6073,N_955,N_3993);
nor U6074 (N_6074,N_1142,N_2034);
nand U6075 (N_6075,N_1969,N_2495);
and U6076 (N_6076,N_4851,N_984);
or U6077 (N_6077,N_1568,N_3712);
and U6078 (N_6078,N_2741,N_4053);
xor U6079 (N_6079,N_5226,N_1330);
and U6080 (N_6080,N_4805,N_3472);
or U6081 (N_6081,N_3852,N_5255);
and U6082 (N_6082,N_5791,N_1603);
or U6083 (N_6083,N_5693,N_2547);
and U6084 (N_6084,N_5258,N_2147);
and U6085 (N_6085,N_3500,N_5980);
or U6086 (N_6086,N_5819,N_304);
xor U6087 (N_6087,N_2503,N_5378);
xnor U6088 (N_6088,N_4362,N_1078);
nand U6089 (N_6089,N_5062,N_3487);
nand U6090 (N_6090,N_977,N_62);
nor U6091 (N_6091,N_5410,N_5024);
nand U6092 (N_6092,N_2037,N_4271);
and U6093 (N_6093,N_300,N_3766);
xnor U6094 (N_6094,N_5412,N_5992);
nand U6095 (N_6095,N_3097,N_1356);
nor U6096 (N_6096,N_5265,N_3091);
xnor U6097 (N_6097,N_2258,N_3192);
or U6098 (N_6098,N_5361,N_2432);
or U6099 (N_6099,N_1878,N_3662);
nand U6100 (N_6100,N_274,N_1033);
and U6101 (N_6101,N_3113,N_2305);
xnor U6102 (N_6102,N_2969,N_193);
nor U6103 (N_6103,N_4937,N_1965);
nand U6104 (N_6104,N_5556,N_5828);
xor U6105 (N_6105,N_3644,N_5531);
nand U6106 (N_6106,N_4896,N_4244);
nor U6107 (N_6107,N_3023,N_4429);
nand U6108 (N_6108,N_3711,N_4454);
xnor U6109 (N_6109,N_2346,N_982);
nand U6110 (N_6110,N_790,N_1856);
nand U6111 (N_6111,N_1296,N_249);
and U6112 (N_6112,N_3329,N_208);
nand U6113 (N_6113,N_1182,N_3253);
nand U6114 (N_6114,N_278,N_2450);
or U6115 (N_6115,N_3053,N_2944);
and U6116 (N_6116,N_2675,N_561);
xnor U6117 (N_6117,N_42,N_1136);
and U6118 (N_6118,N_1949,N_5568);
and U6119 (N_6119,N_605,N_5493);
or U6120 (N_6120,N_2338,N_882);
nand U6121 (N_6121,N_5987,N_2473);
nand U6122 (N_6122,N_77,N_1508);
and U6123 (N_6123,N_3966,N_4349);
or U6124 (N_6124,N_5632,N_2936);
and U6125 (N_6125,N_4789,N_4436);
xnor U6126 (N_6126,N_4218,N_1524);
or U6127 (N_6127,N_2681,N_1114);
or U6128 (N_6128,N_320,N_1711);
xnor U6129 (N_6129,N_3807,N_4168);
or U6130 (N_6130,N_4124,N_5071);
or U6131 (N_6131,N_1951,N_3088);
nor U6132 (N_6132,N_4389,N_4886);
and U6133 (N_6133,N_3209,N_2630);
nor U6134 (N_6134,N_5484,N_5550);
nand U6135 (N_6135,N_999,N_3095);
nor U6136 (N_6136,N_692,N_3439);
nor U6137 (N_6137,N_555,N_5129);
and U6138 (N_6138,N_2613,N_2172);
and U6139 (N_6139,N_1466,N_3579);
or U6140 (N_6140,N_2697,N_2218);
or U6141 (N_6141,N_2818,N_2386);
or U6142 (N_6142,N_2102,N_513);
nand U6143 (N_6143,N_671,N_1443);
and U6144 (N_6144,N_1082,N_3056);
xor U6145 (N_6145,N_1780,N_1805);
nand U6146 (N_6146,N_5033,N_795);
nand U6147 (N_6147,N_1191,N_611);
nor U6148 (N_6148,N_5869,N_1932);
nand U6149 (N_6149,N_2597,N_4859);
or U6150 (N_6150,N_2314,N_552);
nor U6151 (N_6151,N_2946,N_4522);
or U6152 (N_6152,N_1439,N_148);
nand U6153 (N_6153,N_5726,N_752);
xor U6154 (N_6154,N_593,N_5518);
nor U6155 (N_6155,N_4101,N_3482);
nand U6156 (N_6156,N_5430,N_5668);
or U6157 (N_6157,N_5114,N_4479);
or U6158 (N_6158,N_2966,N_3921);
or U6159 (N_6159,N_3320,N_5525);
nor U6160 (N_6160,N_2005,N_4040);
and U6161 (N_6161,N_4405,N_5800);
and U6162 (N_6162,N_4291,N_4832);
and U6163 (N_6163,N_4251,N_3188);
xor U6164 (N_6164,N_2988,N_68);
nand U6165 (N_6165,N_856,N_5465);
nand U6166 (N_6166,N_2576,N_5852);
nand U6167 (N_6167,N_1945,N_310);
xnor U6168 (N_6168,N_1791,N_1071);
and U6169 (N_6169,N_600,N_3626);
or U6170 (N_6170,N_1898,N_2786);
nor U6171 (N_6171,N_1505,N_2282);
or U6172 (N_6172,N_2500,N_1044);
and U6173 (N_6173,N_5134,N_4467);
nor U6174 (N_6174,N_3984,N_2371);
xnor U6175 (N_6175,N_241,N_5444);
nand U6176 (N_6176,N_1510,N_5535);
nand U6177 (N_6177,N_3586,N_47);
xor U6178 (N_6178,N_306,N_4706);
nor U6179 (N_6179,N_3350,N_41);
nand U6180 (N_6180,N_5393,N_2856);
nor U6181 (N_6181,N_4226,N_5399);
nand U6182 (N_6182,N_2385,N_3715);
or U6183 (N_6183,N_1040,N_154);
xor U6184 (N_6184,N_5857,N_1377);
xor U6185 (N_6185,N_136,N_3696);
nand U6186 (N_6186,N_5730,N_5578);
and U6187 (N_6187,N_4248,N_886);
xnor U6188 (N_6188,N_1297,N_230);
nand U6189 (N_6189,N_4686,N_3108);
and U6190 (N_6190,N_821,N_2478);
or U6191 (N_6191,N_5435,N_24);
xor U6192 (N_6192,N_840,N_3466);
or U6193 (N_6193,N_3292,N_2192);
nand U6194 (N_6194,N_3714,N_4818);
xor U6195 (N_6195,N_2884,N_5079);
xnor U6196 (N_6196,N_516,N_5553);
and U6197 (N_6197,N_4588,N_530);
xnor U6198 (N_6198,N_4310,N_2126);
nand U6199 (N_6199,N_811,N_1453);
xor U6200 (N_6200,N_1794,N_5935);
xor U6201 (N_6201,N_5183,N_4756);
or U6202 (N_6202,N_4376,N_5811);
nor U6203 (N_6203,N_2539,N_4863);
or U6204 (N_6204,N_5692,N_266);
or U6205 (N_6205,N_5585,N_5542);
or U6206 (N_6206,N_2079,N_1408);
nor U6207 (N_6207,N_4192,N_2110);
and U6208 (N_6208,N_2337,N_1336);
xor U6209 (N_6209,N_4512,N_2238);
and U6210 (N_6210,N_4509,N_5657);
nor U6211 (N_6211,N_724,N_3140);
nor U6212 (N_6212,N_2379,N_5873);
or U6213 (N_6213,N_5415,N_3264);
xnor U6214 (N_6214,N_2179,N_71);
or U6215 (N_6215,N_3266,N_4525);
nand U6216 (N_6216,N_4718,N_1626);
and U6217 (N_6217,N_3658,N_1425);
xor U6218 (N_6218,N_5087,N_616);
or U6219 (N_6219,N_146,N_4545);
and U6220 (N_6220,N_5534,N_850);
nor U6221 (N_6221,N_5608,N_1677);
xnor U6222 (N_6222,N_1052,N_5073);
nand U6223 (N_6223,N_5729,N_1762);
and U6224 (N_6224,N_3717,N_2970);
or U6225 (N_6225,N_3862,N_2502);
nand U6226 (N_6226,N_914,N_403);
nor U6227 (N_6227,N_5609,N_1778);
and U6228 (N_6228,N_2879,N_831);
nand U6229 (N_6229,N_662,N_4796);
or U6230 (N_6230,N_1576,N_4421);
xor U6231 (N_6231,N_5708,N_4627);
xor U6232 (N_6232,N_1790,N_1321);
or U6233 (N_6233,N_4704,N_3226);
xor U6234 (N_6234,N_1569,N_3032);
xnor U6235 (N_6235,N_5333,N_5326);
nand U6236 (N_6236,N_1300,N_4528);
nand U6237 (N_6237,N_5293,N_4901);
nand U6238 (N_6238,N_265,N_2727);
nand U6239 (N_6239,N_5453,N_825);
or U6240 (N_6240,N_2352,N_4883);
xnor U6241 (N_6241,N_2051,N_5470);
and U6242 (N_6242,N_387,N_1746);
or U6243 (N_6243,N_80,N_2104);
xor U6244 (N_6244,N_4270,N_694);
nor U6245 (N_6245,N_4866,N_1743);
or U6246 (N_6246,N_4254,N_3628);
and U6247 (N_6247,N_3259,N_4952);
nor U6248 (N_6248,N_3240,N_958);
or U6249 (N_6249,N_829,N_889);
or U6250 (N_6250,N_766,N_1387);
nor U6251 (N_6251,N_4878,N_3869);
nand U6252 (N_6252,N_3607,N_2999);
nor U6253 (N_6253,N_1039,N_5508);
or U6254 (N_6254,N_2203,N_4116);
nand U6255 (N_6255,N_2522,N_428);
nand U6256 (N_6256,N_5546,N_4196);
nor U6257 (N_6257,N_273,N_1516);
nor U6258 (N_6258,N_1064,N_5377);
xnor U6259 (N_6259,N_727,N_2178);
nor U6260 (N_6260,N_4430,N_580);
and U6261 (N_6261,N_2116,N_3443);
nor U6262 (N_6262,N_2713,N_4850);
xor U6263 (N_6263,N_16,N_2509);
or U6264 (N_6264,N_1134,N_5081);
nor U6265 (N_6265,N_2210,N_5058);
nand U6266 (N_6266,N_4957,N_698);
and U6267 (N_6267,N_3496,N_3647);
or U6268 (N_6268,N_19,N_1098);
xnor U6269 (N_6269,N_269,N_3392);
and U6270 (N_6270,N_5922,N_4766);
nand U6271 (N_6271,N_3217,N_4170);
and U6272 (N_6272,N_5458,N_4769);
xnor U6273 (N_6273,N_1083,N_5133);
and U6274 (N_6274,N_507,N_3962);
nand U6275 (N_6275,N_771,N_5923);
and U6276 (N_6276,N_2068,N_2762);
and U6277 (N_6277,N_383,N_4378);
nor U6278 (N_6278,N_2619,N_4334);
and U6279 (N_6279,N_3096,N_1964);
and U6280 (N_6280,N_4162,N_2973);
xnor U6281 (N_6281,N_3234,N_1348);
or U6282 (N_6282,N_4377,N_5502);
nor U6283 (N_6283,N_1515,N_3521);
nor U6284 (N_6284,N_121,N_910);
nor U6285 (N_6285,N_5771,N_4036);
xor U6286 (N_6286,N_342,N_891);
xor U6287 (N_6287,N_2382,N_5953);
or U6288 (N_6288,N_4930,N_3795);
xnor U6289 (N_6289,N_4616,N_4201);
nor U6290 (N_6290,N_5834,N_515);
nand U6291 (N_6291,N_2420,N_4771);
and U6292 (N_6292,N_2801,N_4535);
and U6293 (N_6293,N_5532,N_2044);
and U6294 (N_6294,N_4111,N_2082);
or U6295 (N_6295,N_5775,N_4665);
nand U6296 (N_6296,N_3702,N_1607);
xnor U6297 (N_6297,N_2223,N_1392);
nor U6298 (N_6298,N_4327,N_4680);
xor U6299 (N_6299,N_4469,N_520);
and U6300 (N_6300,N_3133,N_3815);
or U6301 (N_6301,N_1204,N_5084);
and U6302 (N_6302,N_2746,N_5674);
and U6303 (N_6303,N_2732,N_4643);
nand U6304 (N_6304,N_1167,N_1831);
nand U6305 (N_6305,N_4138,N_859);
nor U6306 (N_6306,N_3725,N_905);
nand U6307 (N_6307,N_3344,N_5711);
nand U6308 (N_6308,N_5208,N_5249);
and U6309 (N_6309,N_4239,N_4749);
xor U6310 (N_6310,N_2123,N_5191);
and U6311 (N_6311,N_3082,N_1470);
nor U6312 (N_6312,N_1539,N_789);
or U6313 (N_6313,N_4060,N_739);
nor U6314 (N_6314,N_1988,N_4956);
xor U6315 (N_6315,N_5901,N_2813);
nor U6316 (N_6316,N_1017,N_5276);
and U6317 (N_6317,N_736,N_1260);
nor U6318 (N_6318,N_1877,N_1995);
nor U6319 (N_6319,N_1776,N_3200);
nor U6320 (N_6320,N_2169,N_2531);
or U6321 (N_6321,N_1035,N_5120);
nor U6322 (N_6322,N_2186,N_729);
xor U6323 (N_6323,N_2039,N_3299);
nand U6324 (N_6324,N_3052,N_2206);
and U6325 (N_6325,N_673,N_5035);
and U6326 (N_6326,N_802,N_961);
and U6327 (N_6327,N_4698,N_259);
nand U6328 (N_6328,N_4417,N_4216);
and U6329 (N_6329,N_1504,N_2898);
xnor U6330 (N_6330,N_5408,N_395);
nand U6331 (N_6331,N_26,N_1821);
or U6332 (N_6332,N_484,N_5720);
xnor U6333 (N_6333,N_5779,N_930);
nand U6334 (N_6334,N_4795,N_1154);
nand U6335 (N_6335,N_2392,N_2872);
nor U6336 (N_6336,N_446,N_1146);
nor U6337 (N_6337,N_813,N_5314);
xor U6338 (N_6338,N_444,N_1616);
xnor U6339 (N_6339,N_5085,N_5786);
nand U6340 (N_6340,N_4985,N_2558);
nor U6341 (N_6341,N_581,N_443);
nand U6342 (N_6342,N_4275,N_74);
nor U6343 (N_6343,N_1554,N_5623);
xnor U6344 (N_6344,N_2439,N_3231);
nor U6345 (N_6345,N_2081,N_1563);
nor U6346 (N_6346,N_2569,N_296);
or U6347 (N_6347,N_1904,N_4614);
nor U6348 (N_6348,N_1653,N_1461);
xor U6349 (N_6349,N_1830,N_5911);
or U6350 (N_6350,N_5675,N_1529);
xor U6351 (N_6351,N_504,N_5880);
nand U6352 (N_6352,N_5101,N_2640);
xor U6353 (N_6353,N_2268,N_1481);
and U6354 (N_6354,N_1625,N_10);
nor U6355 (N_6355,N_2738,N_5492);
xnor U6356 (N_6356,N_38,N_492);
or U6357 (N_6357,N_4677,N_5591);
and U6358 (N_6358,N_1415,N_209);
xnor U6359 (N_6359,N_1641,N_3076);
nor U6360 (N_6360,N_4852,N_3761);
and U6361 (N_6361,N_3218,N_4158);
or U6362 (N_6362,N_1020,N_5936);
nand U6363 (N_6363,N_2878,N_5306);
or U6364 (N_6364,N_4716,N_627);
and U6365 (N_6365,N_5193,N_883);
and U6366 (N_6366,N_3641,N_5433);
xor U6367 (N_6367,N_5769,N_5978);
nand U6368 (N_6368,N_4048,N_3405);
nand U6369 (N_6369,N_2686,N_3823);
and U6370 (N_6370,N_1803,N_3423);
or U6371 (N_6371,N_2611,N_1250);
or U6372 (N_6372,N_2890,N_385);
and U6373 (N_6373,N_5115,N_5481);
xnor U6374 (N_6374,N_4077,N_5069);
nor U6375 (N_6375,N_4422,N_1249);
nand U6376 (N_6376,N_4633,N_494);
and U6377 (N_6377,N_1286,N_2167);
xor U6378 (N_6378,N_2855,N_2937);
or U6379 (N_6379,N_2508,N_5710);
xnor U6380 (N_6380,N_1946,N_2580);
and U6381 (N_6381,N_2029,N_615);
nand U6382 (N_6382,N_1474,N_5627);
nor U6383 (N_6383,N_757,N_5050);
nor U6384 (N_6384,N_1196,N_3001);
nand U6385 (N_6385,N_3832,N_1660);
nor U6386 (N_6386,N_473,N_3105);
nor U6387 (N_6387,N_2475,N_2491);
and U6388 (N_6388,N_503,N_5123);
and U6389 (N_6389,N_2776,N_2556);
or U6390 (N_6390,N_5218,N_5573);
nand U6391 (N_6391,N_1756,N_1661);
nand U6392 (N_6392,N_5949,N_1360);
nand U6393 (N_6393,N_5650,N_4856);
xnor U6394 (N_6394,N_4484,N_3239);
nand U6395 (N_6395,N_3413,N_5958);
and U6396 (N_6396,N_2634,N_3885);
and U6397 (N_6397,N_4758,N_4807);
or U6398 (N_6398,N_2482,N_1495);
or U6399 (N_6399,N_4470,N_364);
and U6400 (N_6400,N_3447,N_2365);
xor U6401 (N_6401,N_4656,N_2868);
or U6402 (N_6402,N_3590,N_2889);
nand U6403 (N_6403,N_3254,N_1521);
nor U6404 (N_6404,N_1061,N_3942);
xnor U6405 (N_6405,N_4755,N_2158);
nand U6406 (N_6406,N_4477,N_4563);
nand U6407 (N_6407,N_1446,N_5827);
xnor U6408 (N_6408,N_3036,N_5469);
or U6409 (N_6409,N_2730,N_5312);
xnor U6410 (N_6410,N_2673,N_3808);
and U6411 (N_6411,N_4829,N_5227);
and U6412 (N_6412,N_4876,N_164);
nand U6413 (N_6413,N_1939,N_5979);
nand U6414 (N_6414,N_4935,N_1367);
xor U6415 (N_6415,N_1719,N_2941);
xnor U6416 (N_6416,N_4503,N_4373);
xnor U6417 (N_6417,N_1857,N_1724);
or U6418 (N_6418,N_4432,N_4455);
nand U6419 (N_6419,N_2836,N_4202);
or U6420 (N_6420,N_1523,N_2978);
nor U6421 (N_6421,N_5931,N_699);
xor U6422 (N_6422,N_5856,N_5432);
nor U6423 (N_6423,N_2883,N_4604);
nand U6424 (N_6424,N_5658,N_2520);
nor U6425 (N_6425,N_5400,N_1272);
and U6426 (N_6426,N_3886,N_5392);
nor U6427 (N_6427,N_4471,N_402);
or U6428 (N_6428,N_3778,N_4409);
nor U6429 (N_6429,N_971,N_1430);
nand U6430 (N_6430,N_3168,N_5130);
xnor U6431 (N_6431,N_1934,N_1737);
or U6432 (N_6432,N_5054,N_1110);
and U6433 (N_6433,N_5862,N_550);
nand U6434 (N_6434,N_5239,N_1894);
nor U6435 (N_6435,N_248,N_1809);
xnor U6436 (N_6436,N_1157,N_4641);
or U6437 (N_6437,N_5135,N_3461);
or U6438 (N_6438,N_3260,N_420);
or U6439 (N_6439,N_3464,N_5749);
nor U6440 (N_6440,N_3436,N_3044);
or U6441 (N_6441,N_3833,N_4324);
nand U6442 (N_6442,N_5558,N_397);
and U6443 (N_6443,N_1604,N_634);
and U6444 (N_6444,N_5881,N_3939);
nand U6445 (N_6445,N_1145,N_3196);
or U6446 (N_6446,N_5803,N_2571);
and U6447 (N_6447,N_4980,N_4508);
xor U6448 (N_6448,N_170,N_493);
nand U6449 (N_6449,N_2026,N_3089);
nor U6450 (N_6450,N_4290,N_5042);
nand U6451 (N_6451,N_375,N_107);
nor U6452 (N_6452,N_4717,N_3399);
or U6453 (N_6453,N_5411,N_5288);
nor U6454 (N_6454,N_2084,N_3750);
nand U6455 (N_6455,N_2842,N_4887);
xor U6456 (N_6456,N_5930,N_92);
xor U6457 (N_6457,N_5629,N_5694);
xor U6458 (N_6458,N_4103,N_4705);
or U6459 (N_6459,N_3549,N_4933);
or U6460 (N_6460,N_5634,N_3119);
and U6461 (N_6461,N_5398,N_5991);
nand U6462 (N_6462,N_2415,N_1295);
or U6463 (N_6463,N_4493,N_225);
nand U6464 (N_6464,N_5626,N_5143);
or U6465 (N_6465,N_117,N_1271);
xnor U6466 (N_6466,N_628,N_1896);
and U6467 (N_6467,N_5519,N_58);
and U6468 (N_6468,N_389,N_4618);
nand U6469 (N_6469,N_2261,N_872);
xnor U6470 (N_6470,N_1646,N_1276);
and U6471 (N_6471,N_5918,N_4355);
nor U6472 (N_6472,N_3655,N_30);
and U6473 (N_6473,N_1006,N_445);
and U6474 (N_6474,N_5773,N_911);
xor U6475 (N_6475,N_4671,N_5487);
or U6476 (N_6476,N_1713,N_741);
xnor U6477 (N_6477,N_745,N_104);
nand U6478 (N_6478,N_5160,N_338);
nand U6479 (N_6479,N_4833,N_2269);
and U6480 (N_6480,N_195,N_4543);
xor U6481 (N_6481,N_2685,N_1895);
xor U6482 (N_6482,N_832,N_4287);
and U6483 (N_6483,N_3879,N_4434);
nor U6484 (N_6484,N_373,N_3749);
nor U6485 (N_6485,N_2677,N_332);
nand U6486 (N_6486,N_2705,N_3326);
nor U6487 (N_6487,N_3755,N_1268);
nor U6488 (N_6488,N_3765,N_5499);
and U6489 (N_6489,N_3619,N_788);
and U6490 (N_6490,N_5217,N_702);
nand U6491 (N_6491,N_5871,N_3182);
nand U6492 (N_6492,N_4017,N_4647);
nand U6493 (N_6493,N_1116,N_1642);
and U6494 (N_6494,N_743,N_1047);
and U6495 (N_6495,N_3724,N_160);
and U6496 (N_6496,N_450,N_5971);
and U6497 (N_6497,N_1143,N_5677);
xnor U6498 (N_6498,N_1889,N_3727);
nand U6499 (N_6499,N_1901,N_4157);
or U6500 (N_6500,N_483,N_2907);
and U6501 (N_6501,N_3614,N_5295);
or U6502 (N_6502,N_3334,N_5696);
or U6503 (N_6503,N_1839,N_1081);
nand U6504 (N_6504,N_528,N_262);
nand U6505 (N_6505,N_4465,N_3025);
nor U6506 (N_6506,N_2058,N_979);
or U6507 (N_6507,N_3222,N_4064);
nand U6508 (N_6508,N_826,N_4210);
and U6509 (N_6509,N_1594,N_5431);
nor U6510 (N_6510,N_44,N_5667);
nand U6511 (N_6511,N_5064,N_1262);
or U6512 (N_6512,N_798,N_340);
and U6513 (N_6513,N_330,N_5047);
xor U6514 (N_6514,N_2720,N_1881);
nor U6515 (N_6515,N_2809,N_792);
and U6516 (N_6516,N_3703,N_4694);
and U6517 (N_6517,N_2672,N_2751);
nand U6518 (N_6518,N_1156,N_78);
or U6519 (N_6519,N_4444,N_667);
and U6520 (N_6520,N_5555,N_5182);
nand U6521 (N_6521,N_4893,N_4517);
or U6522 (N_6522,N_5316,N_5080);
or U6523 (N_6523,N_404,N_2668);
xor U6524 (N_6524,N_1266,N_3587);
and U6525 (N_6525,N_2843,N_1591);
or U6526 (N_6526,N_5462,N_3567);
nor U6527 (N_6527,N_1623,N_119);
xor U6528 (N_6528,N_4300,N_2765);
and U6529 (N_6529,N_360,N_1873);
xnor U6530 (N_6530,N_11,N_5954);
and U6531 (N_6531,N_423,N_2281);
and U6532 (N_6532,N_3493,N_1967);
nand U6533 (N_6533,N_4842,N_2035);
xnor U6534 (N_6534,N_2614,N_1283);
and U6535 (N_6535,N_4760,N_499);
nand U6536 (N_6536,N_1292,N_5806);
nor U6537 (N_6537,N_4426,N_3408);
nor U6538 (N_6538,N_315,N_5438);
xnor U6539 (N_6539,N_2781,N_5660);
or U6540 (N_6540,N_1096,N_3297);
nand U6541 (N_6541,N_1552,N_3700);
or U6542 (N_6542,N_1577,N_1337);
nor U6543 (N_6543,N_3184,N_3035);
xnor U6544 (N_6544,N_1565,N_3632);
or U6545 (N_6545,N_3764,N_4079);
xor U6546 (N_6546,N_5343,N_3840);
and U6547 (N_6547,N_23,N_3215);
nor U6548 (N_6548,N_4284,N_784);
nor U6549 (N_6549,N_1958,N_3558);
nor U6550 (N_6550,N_5009,N_1555);
and U6551 (N_6551,N_3578,N_870);
nor U6552 (N_6552,N_2783,N_598);
nor U6553 (N_6553,N_2222,N_5428);
nor U6554 (N_6554,N_2541,N_1981);
and U6555 (N_6555,N_3440,N_2642);
or U6556 (N_6556,N_3068,N_3554);
or U6557 (N_6557,N_3572,N_2799);
nor U6558 (N_6558,N_3288,N_5792);
and U6559 (N_6559,N_3884,N_2804);
or U6560 (N_6560,N_256,N_3925);
and U6561 (N_6561,N_647,N_2911);
nand U6562 (N_6562,N_1076,N_5236);
xor U6563 (N_6563,N_5798,N_4780);
xor U6564 (N_6564,N_3528,N_3406);
nor U6565 (N_6565,N_4763,N_5474);
and U6566 (N_6566,N_2251,N_1582);
nor U6567 (N_6567,N_5601,N_3835);
nand U6568 (N_6568,N_2773,N_5164);
nor U6569 (N_6569,N_257,N_5820);
and U6570 (N_6570,N_1059,N_3713);
or U6571 (N_6571,N_4581,N_1175);
xor U6572 (N_6572,N_996,N_1090);
xor U6573 (N_6573,N_286,N_396);
nand U6574 (N_6574,N_1121,N_1043);
and U6575 (N_6575,N_2092,N_3825);
nor U6576 (N_6576,N_341,N_1199);
xor U6577 (N_6577,N_4553,N_2231);
xor U6578 (N_6578,N_1977,N_3760);
xnor U6579 (N_6579,N_369,N_4009);
xor U6580 (N_6580,N_3762,N_1910);
nand U6581 (N_6581,N_4181,N_1586);
and U6582 (N_6582,N_800,N_4076);
nor U6583 (N_6583,N_5441,N_5089);
nand U6584 (N_6584,N_102,N_1085);
nand U6585 (N_6585,N_5890,N_3826);
nand U6586 (N_6586,N_1548,N_4054);
and U6587 (N_6587,N_4757,N_178);
nand U6588 (N_6588,N_868,N_3454);
and U6589 (N_6589,N_2280,N_3946);
and U6590 (N_6590,N_2234,N_1170);
and U6591 (N_6591,N_252,N_1238);
nand U6592 (N_6592,N_1537,N_3067);
xor U6593 (N_6593,N_144,N_716);
nand U6594 (N_6594,N_3637,N_1701);
xor U6595 (N_6595,N_5809,N_1089);
and U6596 (N_6596,N_3505,N_1580);
and U6597 (N_6597,N_2111,N_5599);
or U6598 (N_6598,N_2,N_2758);
nor U6599 (N_6599,N_372,N_1437);
nand U6600 (N_6600,N_2639,N_2959);
or U6601 (N_6601,N_2285,N_2401);
and U6602 (N_6602,N_2426,N_3653);
nand U6603 (N_6603,N_5476,N_1131);
xor U6604 (N_6604,N_1479,N_2893);
or U6605 (N_6605,N_40,N_1789);
or U6606 (N_6606,N_2347,N_3092);
and U6607 (N_6607,N_5996,N_5743);
and U6608 (N_6608,N_3375,N_2187);
or U6609 (N_6609,N_542,N_4137);
nor U6610 (N_6610,N_5687,N_1538);
nand U6611 (N_6611,N_53,N_2953);
and U6612 (N_6612,N_4984,N_2935);
nand U6613 (N_6613,N_4365,N_1027);
or U6614 (N_6614,N_1458,N_1026);
xnor U6615 (N_6615,N_3978,N_2094);
nand U6616 (N_6616,N_5808,N_4055);
nor U6617 (N_6617,N_1115,N_66);
nand U6618 (N_6618,N_1612,N_5207);
and U6619 (N_6619,N_2598,N_506);
and U6620 (N_6620,N_228,N_3280);
or U6621 (N_6621,N_5745,N_1369);
nand U6622 (N_6622,N_2201,N_1370);
nand U6623 (N_6623,N_2933,N_3843);
nand U6624 (N_6624,N_240,N_860);
xnor U6625 (N_6625,N_4721,N_780);
nand U6626 (N_6626,N_1957,N_4203);
and U6627 (N_6627,N_4691,N_2564);
or U6628 (N_6628,N_5165,N_5395);
and U6629 (N_6629,N_2894,N_617);
or U6630 (N_6630,N_1477,N_764);
nor U6631 (N_6631,N_3074,N_5442);
nand U6632 (N_6632,N_5025,N_5715);
xor U6633 (N_6633,N_609,N_5521);
and U6634 (N_6634,N_4898,N_2715);
xnor U6635 (N_6635,N_5993,N_5283);
nor U6636 (N_6636,N_894,N_2160);
nand U6637 (N_6637,N_4904,N_1596);
nor U6638 (N_6638,N_1812,N_5455);
xnor U6639 (N_6639,N_1813,N_2529);
or U6640 (N_6640,N_4462,N_4448);
nor U6641 (N_6641,N_3983,N_223);
nand U6642 (N_6642,N_4252,N_1184);
nand U6643 (N_6643,N_4206,N_1650);
nand U6644 (N_6644,N_5374,N_5046);
nor U6645 (N_6645,N_2824,N_5406);
nand U6646 (N_6646,N_509,N_4450);
or U6647 (N_6647,N_5947,N_3109);
or U6648 (N_6648,N_939,N_1150);
nor U6649 (N_6649,N_814,N_2984);
and U6650 (N_6650,N_2245,N_3923);
nand U6651 (N_6651,N_2003,N_5309);
nand U6652 (N_6652,N_3296,N_2632);
xor U6653 (N_6653,N_4359,N_4172);
and U6654 (N_6654,N_1449,N_1973);
or U6655 (N_6655,N_2655,N_290);
nand U6656 (N_6656,N_5121,N_5338);
nor U6657 (N_6657,N_1129,N_4309);
or U6658 (N_6658,N_4446,N_4283);
or U6659 (N_6659,N_2185,N_522);
nor U6660 (N_6660,N_5043,N_2601);
nand U6661 (N_6661,N_3033,N_5059);
xor U6662 (N_6662,N_5912,N_865);
and U6663 (N_6663,N_756,N_2056);
nand U6664 (N_6664,N_1592,N_2696);
nor U6665 (N_6665,N_263,N_936);
and U6666 (N_6666,N_4399,N_1971);
and U6667 (N_6667,N_352,N_356);
nand U6668 (N_6668,N_2168,N_2004);
or U6669 (N_6669,N_4619,N_2402);
xor U6670 (N_6670,N_5419,N_5507);
xnor U6671 (N_6671,N_1427,N_2551);
and U6672 (N_6672,N_465,N_5848);
or U6673 (N_6673,N_539,N_1097);
nor U6674 (N_6674,N_2220,N_896);
and U6675 (N_6675,N_4474,N_1753);
nand U6676 (N_6676,N_4658,N_1551);
and U6677 (N_6677,N_2735,N_796);
nor U6678 (N_6678,N_1624,N_3455);
nor U6679 (N_6679,N_3695,N_4169);
xor U6680 (N_6680,N_438,N_69);
xnor U6681 (N_6681,N_496,N_904);
nand U6682 (N_6682,N_4862,N_2631);
and U6683 (N_6683,N_2925,N_4719);
nand U6684 (N_6684,N_3251,N_963);
nor U6685 (N_6685,N_327,N_5371);
or U6686 (N_6686,N_4595,N_5007);
xnor U6687 (N_6687,N_5032,N_2410);
nor U6688 (N_6688,N_5144,N_368);
or U6689 (N_6689,N_3523,N_3726);
xnor U6690 (N_6690,N_2289,N_5188);
nand U6691 (N_6691,N_3739,N_2526);
nor U6692 (N_6692,N_291,N_2940);
xor U6693 (N_6693,N_3013,N_5631);
and U6694 (N_6694,N_4848,N_4058);
nand U6695 (N_6695,N_1229,N_5274);
nand U6696 (N_6696,N_2774,N_5480);
and U6697 (N_6697,N_5661,N_1103);
xnor U6698 (N_6698,N_1740,N_4306);
or U6699 (N_6699,N_3498,N_1528);
xnor U6700 (N_6700,N_5616,N_1574);
or U6701 (N_6701,N_3045,N_4521);
or U6702 (N_6702,N_98,N_4117);
or U6703 (N_6703,N_5539,N_5788);
and U6704 (N_6704,N_4225,N_3643);
nand U6705 (N_6705,N_5695,N_421);
xnor U6706 (N_6706,N_5299,N_3685);
or U6707 (N_6707,N_4261,N_1084);
and U6708 (N_6708,N_621,N_1587);
nor U6709 (N_6709,N_2396,N_957);
or U6710 (N_6710,N_678,N_303);
nand U6711 (N_6711,N_3066,N_2484);
or U6712 (N_6712,N_3585,N_3284);
or U6713 (N_6713,N_2001,N_254);
nand U6714 (N_6714,N_4629,N_1828);
nor U6715 (N_6715,N_3343,N_1312);
xnor U6716 (N_6716,N_5607,N_2593);
xor U6717 (N_6717,N_4737,N_4999);
nand U6718 (N_6718,N_3174,N_3570);
or U6719 (N_6719,N_3214,N_3888);
nor U6720 (N_6720,N_2976,N_3009);
xor U6721 (N_6721,N_4331,N_2718);
nand U6722 (N_6722,N_2916,N_2019);
and U6723 (N_6723,N_3332,N_1333);
nor U6724 (N_6724,N_2333,N_5349);
nand U6725 (N_6725,N_4958,N_3330);
xor U6726 (N_6726,N_3988,N_3152);
xor U6727 (N_6727,N_4481,N_4964);
or U6728 (N_6728,N_5229,N_4867);
and U6729 (N_6729,N_2805,N_361);
nor U6730 (N_6730,N_1810,N_5180);
xnor U6731 (N_6731,N_3051,N_5617);
and U6732 (N_6732,N_34,N_3692);
nor U6733 (N_6733,N_2777,N_4514);
and U6734 (N_6734,N_4890,N_2154);
or U6735 (N_6735,N_1093,N_5673);
nand U6736 (N_6736,N_3897,N_4684);
nor U6737 (N_6737,N_4453,N_1021);
nor U6738 (N_6738,N_2263,N_5396);
nand U6739 (N_6739,N_4809,N_2629);
or U6740 (N_6740,N_4148,N_5353);
xnor U6741 (N_6741,N_4183,N_901);
and U6742 (N_6742,N_3610,N_115);
nor U6743 (N_6743,N_1844,N_1704);
nor U6744 (N_6744,N_3061,N_5835);
nor U6745 (N_6745,N_3043,N_314);
nand U6746 (N_6746,N_5206,N_664);
xor U6747 (N_6747,N_3223,N_3961);
and U6748 (N_6748,N_5202,N_72);
and U6749 (N_6749,N_3511,N_3265);
nand U6750 (N_6750,N_3752,N_4778);
and U6751 (N_6751,N_175,N_5286);
nor U6752 (N_6752,N_2072,N_3325);
or U6753 (N_6753,N_2862,N_2109);
and U6754 (N_6754,N_4480,N_5763);
or U6755 (N_6755,N_4959,N_5640);
nor U6756 (N_6756,N_5157,N_365);
nor U6757 (N_6757,N_1251,N_5641);
or U6758 (N_6758,N_2476,N_1566);
and U6759 (N_6759,N_4868,N_5404);
and U6760 (N_6760,N_5948,N_686);
nor U6761 (N_6761,N_5235,N_708);
nand U6762 (N_6762,N_2097,N_2046);
nand U6763 (N_6763,N_1221,N_3497);
and U6764 (N_6764,N_5647,N_5801);
xnor U6765 (N_6765,N_109,N_3740);
xor U6766 (N_6766,N_1243,N_5362);
nor U6767 (N_6767,N_2166,N_134);
or U6768 (N_6768,N_33,N_1560);
or U6769 (N_6769,N_5789,N_5874);
nor U6770 (N_6770,N_4672,N_4384);
nor U6771 (N_6771,N_4452,N_1557);
xnor U6772 (N_6772,N_467,N_1109);
nor U6773 (N_6773,N_1665,N_3502);
nor U6774 (N_6774,N_5966,N_2077);
or U6775 (N_6775,N_3494,N_1025);
and U6776 (N_6776,N_313,N_4791);
xnor U6777 (N_6777,N_871,N_1715);
nor U6778 (N_6778,N_4777,N_837);
or U6779 (N_6779,N_4634,N_2919);
and U6780 (N_6780,N_1469,N_65);
or U6781 (N_6781,N_3448,N_4768);
nand U6782 (N_6782,N_4348,N_759);
xnor U6783 (N_6783,N_4783,N_4810);
or U6784 (N_6784,N_3802,N_879);
xnor U6785 (N_6785,N_2286,N_3542);
nand U6786 (N_6786,N_1180,N_976);
or U6787 (N_6787,N_1190,N_1921);
xor U6788 (N_6788,N_67,N_4743);
nand U6789 (N_6789,N_211,N_1502);
and U6790 (N_6790,N_5590,N_1353);
and U6791 (N_6791,N_3471,N_2207);
xnor U6792 (N_6792,N_3566,N_3782);
nand U6793 (N_6793,N_3742,N_1731);
or U6794 (N_6794,N_2954,N_1181);
xnor U6795 (N_6795,N_2326,N_1597);
nand U6796 (N_6796,N_2825,N_1601);
xnor U6797 (N_6797,N_959,N_3054);
nor U6798 (N_6798,N_1640,N_177);
xnor U6799 (N_6799,N_1606,N_5479);
or U6800 (N_6800,N_3337,N_4590);
and U6801 (N_6801,N_1861,N_15);
xor U6802 (N_6802,N_5359,N_1375);
and U6803 (N_6803,N_1930,N_740);
or U6804 (N_6804,N_3075,N_5831);
nand U6805 (N_6805,N_1902,N_4066);
xnor U6806 (N_6806,N_2972,N_4307);
or U6807 (N_6807,N_4087,N_5466);
nand U6808 (N_6808,N_5733,N_3415);
nand U6809 (N_6809,N_5587,N_4460);
nand U6810 (N_6810,N_5434,N_691);
nand U6811 (N_6811,N_3926,N_4281);
nor U6812 (N_6812,N_765,N_3911);
nor U6813 (N_6813,N_116,N_2811);
nand U6814 (N_6814,N_4742,N_1164);
or U6815 (N_6815,N_1667,N_2979);
nand U6816 (N_6816,N_328,N_1986);
nand U6817 (N_6817,N_1745,N_5676);
or U6818 (N_6818,N_4049,N_5494);
or U6819 (N_6819,N_4397,N_5885);
nand U6820 (N_6820,N_5517,N_3580);
and U6821 (N_6821,N_1381,N_2575);
and U6822 (N_6822,N_5937,N_531);
xor U6823 (N_6823,N_4739,N_1622);
or U6824 (N_6824,N_4182,N_3704);
xnor U6825 (N_6825,N_3998,N_937);
and U6826 (N_6826,N_623,N_822);
xor U6827 (N_6827,N_5019,N_2565);
nand U6828 (N_6828,N_622,N_5889);
nand U6829 (N_6829,N_5976,N_5899);
nor U6830 (N_6830,N_2457,N_204);
nand U6831 (N_6831,N_2349,N_260);
xor U6832 (N_6832,N_1185,N_1310);
and U6833 (N_6833,N_5389,N_2204);
nand U6834 (N_6834,N_5988,N_1849);
xor U6835 (N_6835,N_2055,N_1907);
xnor U6836 (N_6836,N_5298,N_351);
nand U6837 (N_6837,N_3206,N_4788);
or U6838 (N_6838,N_4258,N_1693);
and U6839 (N_6839,N_3341,N_3577);
and U6840 (N_6840,N_3374,N_4630);
or U6841 (N_6841,N_3851,N_5076);
nand U6842 (N_6842,N_4354,N_5031);
and U6843 (N_6843,N_5092,N_5365);
nor U6844 (N_6844,N_2617,N_280);
and U6845 (N_6845,N_4993,N_448);
xor U6846 (N_6846,N_3575,N_5028);
xor U6847 (N_6847,N_5765,N_4846);
nand U6848 (N_6848,N_4382,N_4597);
or U6849 (N_6849,N_3386,N_558);
or U6850 (N_6850,N_3995,N_5596);
nand U6851 (N_6851,N_5266,N_5981);
nor U6852 (N_6852,N_3230,N_4969);
and U6853 (N_6853,N_234,N_4142);
or U6854 (N_6854,N_2359,N_3131);
xor U6855 (N_6855,N_3550,N_3506);
and U6856 (N_6856,N_498,N_2255);
nand U6857 (N_6857,N_277,N_2591);
nand U6858 (N_6858,N_2615,N_2066);
or U6859 (N_6859,N_1378,N_3258);
nor U6860 (N_6860,N_3377,N_5504);
nor U6861 (N_6861,N_1662,N_5997);
xnor U6862 (N_6862,N_2069,N_3323);
and U6863 (N_6863,N_5026,N_1355);
and U6864 (N_6864,N_3428,N_1050);
nor U6865 (N_6865,N_1678,N_4569);
xnor U6866 (N_6866,N_5685,N_3597);
and U6867 (N_6867,N_1852,N_723);
xor U6868 (N_6868,N_5222,N_781);
and U6869 (N_6869,N_4944,N_2098);
xor U6870 (N_6870,N_5074,N_2477);
and U6871 (N_6871,N_5648,N_2448);
or U6872 (N_6872,N_3943,N_1099);
nand U6873 (N_6873,N_2060,N_293);
and U6874 (N_6874,N_142,N_3904);
and U6875 (N_6875,N_4098,N_4090);
xnor U6876 (N_6876,N_5731,N_5664);
nand U6877 (N_6877,N_3902,N_3171);
xor U6878 (N_6878,N_1299,N_5575);
and U6879 (N_6879,N_97,N_3300);
nor U6880 (N_6880,N_418,N_1467);
xnor U6881 (N_6881,N_5083,N_88);
and U6882 (N_6882,N_2653,N_149);
or U6883 (N_6883,N_2949,N_4731);
nor U6884 (N_6884,N_1886,N_2691);
or U6885 (N_6885,N_3831,N_791);
nor U6886 (N_6886,N_5579,N_4330);
or U6887 (N_6887,N_5946,N_912);
nor U6888 (N_6888,N_461,N_3058);
or U6889 (N_6889,N_4916,N_1698);
or U6890 (N_6890,N_5381,N_5612);
and U6891 (N_6891,N_5358,N_4564);
xnor U6892 (N_6892,N_2183,N_3785);
or U6893 (N_6893,N_1435,N_940);
nand U6894 (N_6894,N_3768,N_5669);
nand U6895 (N_6895,N_5440,N_5782);
nor U6896 (N_6896,N_2608,N_4516);
and U6897 (N_6897,N_2790,N_1599);
nand U6898 (N_6898,N_1234,N_876);
nand U6899 (N_6899,N_794,N_2992);
or U6900 (N_6900,N_442,N_393);
nand U6901 (N_6901,N_5697,N_4971);
and U6902 (N_6902,N_2867,N_3369);
nor U6903 (N_6903,N_1779,N_2463);
or U6904 (N_6904,N_4016,N_603);
and U6905 (N_6905,N_1579,N_2716);
nand U6906 (N_6906,N_2582,N_3963);
xor U6907 (N_6907,N_2519,N_4345);
and U6908 (N_6908,N_4441,N_592);
nor U6909 (N_6909,N_3951,N_3268);
nand U6910 (N_6910,N_2095,N_3431);
or U6911 (N_6911,N_1009,N_4440);
xnor U6912 (N_6912,N_2904,N_3770);
nor U6913 (N_6913,N_3720,N_3220);
xnor U6914 (N_6914,N_2293,N_1074);
nor U6915 (N_6915,N_128,N_5457);
and U6916 (N_6916,N_3959,N_343);
or U6917 (N_6917,N_4979,N_5904);
xor U6918 (N_6918,N_1974,N_2224);
or U6919 (N_6919,N_1213,N_630);
or U6920 (N_6920,N_4531,N_4652);
nand U6921 (N_6921,N_519,N_5753);
nor U6922 (N_6922,N_3303,N_3394);
and U6923 (N_6923,N_880,N_4714);
xnor U6924 (N_6924,N_3640,N_5859);
and U6925 (N_6925,N_1388,N_4015);
nor U6926 (N_6926,N_399,N_2180);
nand U6927 (N_6927,N_1670,N_2654);
or U6928 (N_6928,N_2235,N_721);
and U6929 (N_6929,N_4961,N_3973);
nand U6930 (N_6930,N_3992,N_1132);
nor U6931 (N_6931,N_577,N_5810);
and U6932 (N_6932,N_4823,N_1996);
nand U6933 (N_6933,N_848,N_299);
and U6934 (N_6934,N_535,N_4108);
nand U6935 (N_6935,N_4143,N_1485);
nand U6936 (N_6936,N_1287,N_4028);
or U6937 (N_6937,N_635,N_4495);
or U6938 (N_6938,N_3936,N_4062);
xnor U6939 (N_6939,N_5574,N_2324);
nand U6940 (N_6940,N_770,N_5082);
or U6941 (N_6941,N_1241,N_2922);
nor U6942 (N_6942,N_1056,N_5020);
or U6943 (N_6943,N_2648,N_1102);
and U6944 (N_6944,N_3930,N_5443);
and U6945 (N_6945,N_4146,N_5639);
nor U6946 (N_6946,N_1547,N_4687);
xnor U6947 (N_6947,N_1126,N_4660);
and U6948 (N_6948,N_734,N_2709);
or U6949 (N_6949,N_537,N_4071);
xnor U6950 (N_6950,N_4208,N_3812);
or U6951 (N_6951,N_5928,N_2496);
nand U6952 (N_6952,N_5006,N_4713);
nor U6953 (N_6953,N_4892,N_4725);
or U6954 (N_6954,N_5959,N_5619);
xnor U6955 (N_6955,N_3098,N_1922);
nand U6956 (N_6956,N_3999,N_147);
nor U6957 (N_6957,N_312,N_1695);
nand U6958 (N_6958,N_4651,N_4601);
nor U6959 (N_6959,N_5097,N_2011);
nand U6960 (N_6960,N_508,N_924);
nand U6961 (N_6961,N_4967,N_576);
nor U6962 (N_6962,N_3315,N_4962);
nand U6963 (N_6963,N_84,N_1141);
and U6964 (N_6964,N_2253,N_512);
or U6965 (N_6965,N_815,N_3205);
nand U6966 (N_6966,N_4369,N_2574);
and U6967 (N_6967,N_3889,N_2497);
nand U6968 (N_6968,N_1581,N_1933);
or U6969 (N_6969,N_63,N_4125);
and U6970 (N_6970,N_2389,N_4329);
nor U6971 (N_6971,N_2567,N_4052);
xnor U6972 (N_6972,N_487,N_2041);
and U6973 (N_6973,N_3145,N_1380);
or U6974 (N_6974,N_5780,N_4113);
or U6975 (N_6975,N_1991,N_1784);
or U6976 (N_6976,N_2150,N_4176);
nor U6977 (N_6977,N_4804,N_1997);
nand U6978 (N_6978,N_4965,N_3365);
nor U6979 (N_6979,N_1811,N_1696);
nor U6980 (N_6980,N_1217,N_5983);
and U6981 (N_6981,N_2162,N_3031);
nand U6982 (N_6982,N_5250,N_5796);
nor U6983 (N_6983,N_4920,N_3603);
xor U6984 (N_6984,N_5907,N_4140);
nor U6985 (N_6985,N_3007,N_4404);
and U6986 (N_6986,N_2459,N_5955);
xor U6987 (N_6987,N_3387,N_3490);
and U6988 (N_6988,N_1985,N_1162);
and U6989 (N_6989,N_5702,N_2594);
xnor U6990 (N_6990,N_1668,N_998);
nor U6991 (N_6991,N_5606,N_3391);
nor U6992 (N_6992,N_5145,N_1774);
and U6993 (N_6993,N_5533,N_3421);
and U6994 (N_6994,N_2362,N_151);
xnor U6995 (N_6995,N_452,N_477);
xor U6996 (N_6996,N_231,N_5984);
nor U6997 (N_6997,N_2903,N_3005);
nor U6998 (N_6998,N_4692,N_1393);
xor U6999 (N_6999,N_4585,N_1386);
xor U7000 (N_7000,N_3691,N_2679);
and U7001 (N_7001,N_4072,N_2687);
xnor U7002 (N_7002,N_5275,N_4637);
nand U7003 (N_7003,N_4228,N_1211);
nand U7004 (N_7004,N_4010,N_2466);
or U7005 (N_7005,N_4500,N_282);
and U7006 (N_7006,N_1866,N_2638);
nor U7007 (N_7007,N_289,N_921);
and U7008 (N_7008,N_2669,N_5015);
and U7009 (N_7009,N_5757,N_4043);
nor U7010 (N_7010,N_5051,N_525);
nand U7011 (N_7011,N_2880,N_3613);
and U7012 (N_7012,N_5910,N_1797);
or U7013 (N_7013,N_3741,N_1823);
nand U7014 (N_7014,N_656,N_5388);
and U7015 (N_7015,N_4038,N_2405);
or U7016 (N_7016,N_3830,N_3539);
xnor U7017 (N_7017,N_3178,N_5867);
nand U7018 (N_7018,N_1018,N_3745);
nand U7019 (N_7019,N_5595,N_2125);
and U7020 (N_7020,N_5310,N_2375);
and U7021 (N_7021,N_2870,N_892);
nand U7022 (N_7022,N_4437,N_4519);
and U7023 (N_7023,N_207,N_1203);
xnor U7024 (N_7024,N_5,N_2501);
xor U7025 (N_7025,N_4215,N_1478);
nand U7026 (N_7026,N_237,N_4873);
nand U7027 (N_7027,N_527,N_5473);
or U7028 (N_7028,N_3847,N_3124);
or U7029 (N_7029,N_633,N_76);
nor U7030 (N_7030,N_378,N_4669);
nand U7031 (N_7031,N_1593,N_1383);
and U7032 (N_7032,N_712,N_5698);
xor U7033 (N_7033,N_318,N_2000);
nor U7034 (N_7034,N_2849,N_4745);
and U7035 (N_7035,N_227,N_463);
xnor U7036 (N_7036,N_4659,N_810);
xor U7037 (N_7037,N_1339,N_4114);
and U7038 (N_7038,N_4586,N_5103);
or U7039 (N_7039,N_1273,N_1426);
nand U7040 (N_7040,N_4592,N_4815);
or U7041 (N_7041,N_3107,N_2080);
or U7042 (N_7042,N_4625,N_2151);
nor U7043 (N_7043,N_1092,N_3285);
nor U7044 (N_7044,N_4428,N_546);
or U7045 (N_7045,N_2552,N_5228);
xnor U7046 (N_7046,N_2874,N_1879);
xnor U7047 (N_7047,N_4266,N_1371);
and U7048 (N_7048,N_2307,N_544);
and U7049 (N_7049,N_382,N_2036);
nand U7050 (N_7050,N_5939,N_1837);
xnor U7051 (N_7051,N_21,N_711);
or U7052 (N_7052,N_1694,N_1060);
and U7053 (N_7053,N_497,N_4612);
xnor U7054 (N_7054,N_2443,N_2996);
or U7055 (N_7055,N_5201,N_4679);
nor U7056 (N_7056,N_5152,N_390);
nand U7057 (N_7057,N_2232,N_3668);
nor U7058 (N_7058,N_5528,N_4344);
or U7059 (N_7059,N_1208,N_2683);
xnor U7060 (N_7060,N_2527,N_3630);
xnor U7061 (N_7061,N_407,N_4180);
xnor U7062 (N_7062,N_3081,N_4803);
and U7063 (N_7063,N_556,N_4490);
or U7064 (N_7064,N_2317,N_3345);
nor U7065 (N_7065,N_3112,N_3661);
or U7066 (N_7066,N_4534,N_5655);
and U7067 (N_7067,N_3757,N_2604);
nor U7068 (N_7068,N_4,N_1256);
xor U7069 (N_7069,N_4347,N_1739);
and U7070 (N_7070,N_5716,N_5864);
xnor U7071 (N_7071,N_3986,N_1223);
and U7072 (N_7072,N_3608,N_5347);
xor U7073 (N_7073,N_4368,N_5344);
or U7074 (N_7074,N_5700,N_944);
nor U7075 (N_7075,N_3479,N_1870);
xor U7076 (N_7076,N_4255,N_5557);
nand U7077 (N_7077,N_1708,N_2467);
nor U7078 (N_7078,N_2446,N_4081);
and U7079 (N_7079,N_5764,N_3364);
or U7080 (N_7080,N_2388,N_2010);
nor U7081 (N_7081,N_472,N_3533);
nor U7082 (N_7082,N_5016,N_4199);
or U7083 (N_7083,N_596,N_4822);
xor U7084 (N_7084,N_5916,N_1166);
xnor U7085 (N_7085,N_3426,N_4059);
nand U7086 (N_7086,N_5759,N_644);
or U7087 (N_7087,N_1672,N_4298);
and U7088 (N_7088,N_1492,N_3827);
and U7089 (N_7089,N_480,N_5385);
xnor U7090 (N_7090,N_4724,N_847);
xnor U7091 (N_7091,N_3038,N_4827);
xor U7092 (N_7092,N_2309,N_1259);
and U7093 (N_7093,N_5409,N_2743);
nand U7094 (N_7094,N_2678,N_5965);
nand U7095 (N_7095,N_5598,N_3687);
and U7096 (N_7096,N_2692,N_1329);
or U7097 (N_7097,N_3333,N_1655);
or U7098 (N_7098,N_2472,N_1309);
nor U7099 (N_7099,N_3813,N_2666);
nor U7100 (N_7100,N_1950,N_4942);
or U7101 (N_7101,N_2912,N_1073);
nor U7102 (N_7102,N_4574,N_5538);
xor U7103 (N_7103,N_2708,N_1277);
nor U7104 (N_7104,N_2014,N_1149);
or U7105 (N_7105,N_5061,N_5683);
nand U7106 (N_7106,N_5065,N_5691);
nor U7107 (N_7107,N_3524,N_5813);
or U7108 (N_7108,N_3507,N_1897);
nand U7109 (N_7109,N_4385,N_4250);
xnor U7110 (N_7110,N_573,N_4537);
xnor U7111 (N_7111,N_2540,N_1820);
and U7112 (N_7112,N_2882,N_5998);
xor U7113 (N_7113,N_3974,N_1382);
or U7114 (N_7114,N_4955,N_786);
or U7115 (N_7115,N_4265,N_1851);
and U7116 (N_7116,N_3796,N_1984);
nor U7117 (N_7117,N_2423,N_5919);
xor U7118 (N_7118,N_2938,N_4668);
xor U7119 (N_7119,N_441,N_1063);
and U7120 (N_7120,N_5582,N_4664);
or U7121 (N_7121,N_3404,N_2590);
nor U7122 (N_7122,N_3219,N_5030);
xnor U7123 (N_7123,N_2521,N_3589);
xor U7124 (N_7124,N_4046,N_5360);
nor U7125 (N_7125,N_3598,N_5108);
or U7126 (N_7126,N_5752,N_5171);
nand U7127 (N_7127,N_5614,N_588);
nor U7128 (N_7128,N_7,N_2216);
or U7129 (N_7129,N_3871,N_642);
and U7130 (N_7130,N_103,N_3287);
and U7131 (N_7131,N_28,N_3046);
nand U7132 (N_7132,N_4069,N_2826);
and U7133 (N_7133,N_2054,N_3675);
or U7134 (N_7134,N_4457,N_5367);
and U7135 (N_7135,N_3478,N_2328);
xnor U7136 (N_7136,N_5245,N_4864);
nand U7137 (N_7137,N_1088,N_2845);
nor U7138 (N_7138,N_4044,N_1880);
xor U7139 (N_7139,N_2071,N_5351);
nor U7140 (N_7140,N_4416,N_2212);
nor U7141 (N_7141,N_5785,N_2515);
and U7142 (N_7142,N_3102,N_2390);
and U7143 (N_7143,N_5467,N_2339);
xnor U7144 (N_7144,N_474,N_5559);
xor U7145 (N_7145,N_2714,N_3918);
and U7146 (N_7146,N_4151,N_2301);
and U7147 (N_7147,N_1177,N_3228);
and U7148 (N_7148,N_5403,N_4888);
and U7149 (N_7149,N_2771,N_1572);
or U7150 (N_7150,N_3674,N_1032);
and U7151 (N_7151,N_5118,N_5405);
nor U7152 (N_7152,N_2488,N_5510);
or U7153 (N_7153,N_4828,N_4475);
or U7154 (N_7154,N_422,N_3372);
nor U7155 (N_7155,N_3437,N_3743);
xor U7156 (N_7156,N_1553,N_1793);
or U7157 (N_7157,N_2533,N_3649);
and U7158 (N_7158,N_3470,N_1069);
nor U7159 (N_7159,N_2184,N_1752);
or U7160 (N_7160,N_5142,N_619);
and U7161 (N_7161,N_3967,N_3844);
and U7162 (N_7162,N_2798,N_3441);
xor U7163 (N_7163,N_5516,N_5190);
nand U7164 (N_7164,N_4816,N_4813);
or U7165 (N_7165,N_1825,N_348);
nor U7166 (N_7166,N_1445,N_2384);
nand U7167 (N_7167,N_4727,N_5615);
xor U7168 (N_7168,N_4141,N_2040);
nand U7169 (N_7169,N_354,N_2455);
and U7170 (N_7170,N_430,N_4311);
or U7171 (N_7171,N_4599,N_5203);
nor U7172 (N_7172,N_1159,N_3400);
xor U7173 (N_7173,N_250,N_4567);
or U7174 (N_7174,N_4188,N_5390);
or U7175 (N_7175,N_5986,N_1054);
and U7176 (N_7176,N_1559,N_1015);
or U7177 (N_7177,N_2474,N_5717);
nand U7178 (N_7178,N_48,N_3040);
nor U7179 (N_7179,N_1619,N_567);
or U7180 (N_7180,N_5583,N_3356);
xor U7181 (N_7181,N_4338,N_5376);
nand U7182 (N_7182,N_696,N_5439);
nand U7183 (N_7183,N_1424,N_1151);
and U7184 (N_7184,N_5278,N_1633);
xor U7185 (N_7185,N_1233,N_5886);
xnor U7186 (N_7186,N_2243,N_706);
xnor U7187 (N_7187,N_2528,N_3451);
xor U7188 (N_7188,N_4838,N_1514);
xnor U7189 (N_7189,N_242,N_1850);
nand U7190 (N_7190,N_3611,N_1257);
nand U7191 (N_7191,N_4891,N_5659);
and U7192 (N_7192,N_4106,N_3094);
and U7193 (N_7193,N_3368,N_4175);
nand U7194 (N_7194,N_1228,N_4297);
nor U7195 (N_7195,N_4821,N_3388);
or U7196 (N_7196,N_4973,N_4921);
xnor U7197 (N_7197,N_887,N_3773);
nor U7198 (N_7198,N_1230,N_5973);
nand U7199 (N_7199,N_4504,N_3279);
nand U7200 (N_7200,N_5174,N_1068);
and U7201 (N_7201,N_3877,N_4802);
nand U7202 (N_7202,N_4082,N_1338);
nor U7203 (N_7203,N_4025,N_5945);
nor U7204 (N_7204,N_5929,N_1890);
nor U7205 (N_7205,N_2009,N_3663);
nor U7206 (N_7206,N_2960,N_2744);
and U7207 (N_7207,N_3560,N_5475);
nor U7208 (N_7208,N_2876,N_5238);
xnor U7209 (N_7209,N_3639,N_1798);
nand U7210 (N_7210,N_5287,N_5684);
and U7211 (N_7211,N_2769,N_3681);
or U7212 (N_7212,N_2995,N_3697);
xnor U7213 (N_7213,N_707,N_1294);
nor U7214 (N_7214,N_213,N_1671);
nand U7215 (N_7215,N_5758,N_394);
xnor U7216 (N_7216,N_4532,N_5990);
xor U7217 (N_7217,N_335,N_5548);
xor U7218 (N_7218,N_4393,N_5426);
nor U7219 (N_7219,N_4853,N_3924);
nand U7220 (N_7220,N_553,N_991);
and U7221 (N_7221,N_5604,N_2211);
and U7222 (N_7222,N_1952,N_2504);
xor U7223 (N_7223,N_194,N_4747);
and U7224 (N_7224,N_2374,N_4858);
xnor U7225 (N_7225,N_4830,N_2628);
xor U7226 (N_7226,N_2859,N_3916);
or U7227 (N_7227,N_4379,N_5213);
or U7228 (N_7228,N_1999,N_174);
xnor U7229 (N_7229,N_1197,N_3186);
or U7230 (N_7230,N_3103,N_3039);
or U7231 (N_7231,N_737,N_2260);
xnor U7232 (N_7232,N_5327,N_2822);
or U7233 (N_7233,N_2821,N_4520);
nor U7234 (N_7234,N_4744,N_1320);
or U7235 (N_7235,N_5003,N_2544);
nand U7236 (N_7236,N_1647,N_4012);
and U7237 (N_7237,N_4676,N_3252);
nand U7238 (N_7238,N_2858,N_849);
xor U7239 (N_7239,N_1684,N_4366);
xor U7240 (N_7240,N_1832,N_3409);
nand U7241 (N_7241,N_4219,N_3508);
or U7242 (N_7242,N_491,N_3915);
nand U7243 (N_7243,N_774,N_4648);
or U7244 (N_7244,N_2015,N_2236);
and U7245 (N_7245,N_5526,N_4661);
nor U7246 (N_7246,N_3348,N_3449);
and U7247 (N_7247,N_5192,N_1016);
or U7248 (N_7248,N_5570,N_4974);
nor U7249 (N_7249,N_5321,N_5725);
nor U7250 (N_7250,N_2483,N_3380);
or U7251 (N_7251,N_413,N_3269);
nor U7252 (N_7252,N_4022,N_3390);
or U7253 (N_7253,N_5241,N_1128);
and U7254 (N_7254,N_4136,N_3242);
and U7255 (N_7255,N_747,N_1275);
nor U7256 (N_7256,N_4598,N_3803);
nand U7257 (N_7257,N_5454,N_1030);
xnor U7258 (N_7258,N_2427,N_1755);
and U7259 (N_7259,N_4363,N_5109);
nand U7260 (N_7260,N_2917,N_3232);
xor U7261 (N_7261,N_161,N_4968);
nand U7262 (N_7262,N_5603,N_4104);
nor U7263 (N_7263,N_1253,N_4539);
nand U7264 (N_7264,N_2099,N_972);
nand U7265 (N_7265,N_1106,N_2512);
and U7266 (N_7266,N_1070,N_3185);
and U7267 (N_7267,N_4296,N_2722);
xor U7268 (N_7268,N_5825,N_803);
xnor U7269 (N_7269,N_5721,N_4212);
nand U7270 (N_7270,N_4550,N_5893);
and U7271 (N_7271,N_4119,N_5969);
and U7272 (N_7272,N_3636,N_2403);
nor U7273 (N_7273,N_960,N_2647);
nor U7274 (N_7274,N_1125,N_4928);
and U7275 (N_7275,N_5368,N_5537);
xnor U7276 (N_7276,N_2114,N_4001);
or U7277 (N_7277,N_1298,N_2906);
xor U7278 (N_7278,N_2794,N_715);
or U7279 (N_7279,N_5242,N_4607);
nand U7280 (N_7280,N_2703,N_5436);
xnor U7281 (N_7281,N_4869,N_64);
or U7282 (N_7282,N_517,N_1615);
nand U7283 (N_7283,N_55,N_2543);
nor U7284 (N_7284,N_1942,N_137);
nand U7285 (N_7285,N_5995,N_2061);
nor U7286 (N_7286,N_1535,N_1899);
nand U7287 (N_7287,N_2753,N_3893);
nor U7288 (N_7288,N_2288,N_1845);
xnor U7289 (N_7289,N_5748,N_2217);
and U7290 (N_7290,N_43,N_435);
nor U7291 (N_7291,N_2341,N_5078);
nor U7292 (N_7292,N_2242,N_5262);
nand U7293 (N_7293,N_1709,N_5402);
xor U7294 (N_7294,N_658,N_2782);
and U7295 (N_7295,N_2589,N_1501);
and U7296 (N_7296,N_5505,N_4562);
nand U7297 (N_7297,N_3371,N_2411);
nor U7298 (N_7298,N_5416,N_5330);
and U7299 (N_7299,N_3144,N_4230);
xor U7300 (N_7300,N_1595,N_214);
nor U7301 (N_7301,N_281,N_988);
xnor U7302 (N_7302,N_639,N_3177);
and U7303 (N_7303,N_4917,N_143);
and U7304 (N_7304,N_3301,N_4774);
nand U7305 (N_7305,N_5319,N_1413);
and U7306 (N_7306,N_2670,N_1240);
and U7307 (N_7307,N_2143,N_4233);
nor U7308 (N_7308,N_5851,N_321);
and U7309 (N_7309,N_3853,N_91);
xnor U7310 (N_7310,N_1913,N_3517);
and U7311 (N_7311,N_5737,N_2400);
xnor U7312 (N_7312,N_3861,N_3787);
nor U7313 (N_7313,N_654,N_3204);
nand U7314 (N_7314,N_2196,N_3594);
xnor U7315 (N_7315,N_311,N_2174);
nand U7316 (N_7316,N_5933,N_1544);
or U7317 (N_7317,N_5847,N_2393);
nand U7318 (N_7318,N_14,N_3994);
and U7319 (N_7319,N_5551,N_384);
nand U7320 (N_7320,N_2828,N_5925);
nand U7321 (N_7321,N_4456,N_5105);
xor U7322 (N_7322,N_5117,N_1732);
xnor U7323 (N_7323,N_1838,N_3733);
and U7324 (N_7324,N_897,N_3263);
nand U7325 (N_7325,N_319,N_1629);
and U7326 (N_7326,N_1960,N_381);
nor U7327 (N_7327,N_1571,N_1954);
nor U7328 (N_7328,N_922,N_3438);
and U7329 (N_7329,N_3519,N_4626);
or U7330 (N_7330,N_4019,N_1346);
xnor U7331 (N_7331,N_4267,N_4710);
nor U7332 (N_7332,N_948,N_3042);
and U7333 (N_7333,N_2045,N_5185);
and U7334 (N_7334,N_5221,N_1041);
nor U7335 (N_7335,N_3248,N_2877);
nand U7336 (N_7336,N_1385,N_5364);
nand U7337 (N_7337,N_5017,N_1926);
nor U7338 (N_7338,N_2297,N_4530);
nor U7339 (N_7339,N_3679,N_4685);
nor U7340 (N_7340,N_5352,N_5277);
nor U7341 (N_7341,N_2658,N_3485);
nand U7342 (N_7342,N_4526,N_3887);
or U7343 (N_7343,N_538,N_3357);
nor U7344 (N_7344,N_2806,N_5379);
or U7345 (N_7345,N_4502,N_4449);
xnor U7346 (N_7346,N_995,N_3709);
nor U7347 (N_7347,N_1468,N_2820);
nand U7348 (N_7348,N_3346,N_5509);
and U7349 (N_7349,N_4321,N_3656);
nor U7350 (N_7350,N_36,N_1326);
and U7351 (N_7351,N_533,N_3845);
or U7352 (N_7352,N_4277,N_2355);
nand U7353 (N_7353,N_4094,N_4840);
or U7354 (N_7354,N_336,N_3971);
nor U7355 (N_7355,N_5260,N_3600);
nand U7356 (N_7356,N_5512,N_415);
nor U7357 (N_7357,N_4149,N_2327);
nand U7358 (N_7358,N_4923,N_3111);
nor U7359 (N_7359,N_5198,N_5414);
or U7360 (N_7360,N_1423,N_398);
nand U7361 (N_7361,N_2622,N_4280);
nor U7362 (N_7362,N_2620,N_1200);
nand U7363 (N_7363,N_2083,N_2997);
nand U7364 (N_7364,N_4308,N_4943);
or U7365 (N_7365,N_4364,N_4312);
nand U7366 (N_7366,N_4024,N_1632);
or U7367 (N_7367,N_4358,N_429);
and U7368 (N_7368,N_2188,N_4220);
nand U7369 (N_7369,N_4118,N_2726);
nand U7370 (N_7370,N_5237,N_1862);
nand U7371 (N_7371,N_3187,N_809);
nand U7372 (N_7372,N_1448,N_5488);
and U7373 (N_7373,N_5957,N_1511);
nand U7374 (N_7374,N_1585,N_2688);
xnor U7375 (N_7375,N_776,N_4997);
nor U7376 (N_7376,N_2618,N_1107);
xor U7377 (N_7377,N_2241,N_345);
or U7378 (N_7378,N_1703,N_3883);
nor U7379 (N_7379,N_3721,N_1786);
xnor U7380 (N_7380,N_5292,N_1111);
nand U7381 (N_7381,N_3459,N_1530);
nand U7382 (N_7382,N_4420,N_1609);
nand U7383 (N_7383,N_2030,N_5837);
nor U7384 (N_7384,N_3161,N_827);
nand U7385 (N_7385,N_5113,N_4476);
and U7386 (N_7386,N_3819,N_4990);
xor U7387 (N_7387,N_3193,N_414);
xnor U7388 (N_7388,N_2356,N_3559);
or U7389 (N_7389,N_3876,N_3716);
nor U7390 (N_7390,N_408,N_2760);
and U7391 (N_7391,N_3534,N_5581);
and U7392 (N_7392,N_1925,N_3281);
nor U7393 (N_7393,N_5307,N_726);
and U7394 (N_7394,N_4808,N_2834);
or U7395 (N_7395,N_3965,N_5545);
nand U7396 (N_7396,N_4459,N_575);
nand U7397 (N_7397,N_2537,N_2860);
or U7398 (N_7398,N_1072,N_285);
nor U7399 (N_7399,N_4947,N_4189);
nor U7400 (N_7400,N_5342,N_549);
nor U7401 (N_7401,N_4179,N_140);
and U7402 (N_7402,N_5680,N_1533);
and U7403 (N_7403,N_4642,N_3024);
nor U7404 (N_7404,N_3004,N_828);
nor U7405 (N_7405,N_3781,N_2490);
and U7406 (N_7406,N_5220,N_5938);
xnor U7407 (N_7407,N_3317,N_4690);
or U7408 (N_7408,N_3378,N_1007);
nor U7409 (N_7409,N_3304,N_2853);
xor U7410 (N_7410,N_5651,N_5637);
nand U7411 (N_7411,N_1341,N_986);
xnor U7412 (N_7412,N_4989,N_4773);
and U7413 (N_7413,N_2902,N_4105);
xor U7414 (N_7414,N_3213,N_4395);
nor U7415 (N_7415,N_4403,N_3746);
xor U7416 (N_7416,N_2283,N_1301);
or U7417 (N_7417,N_2149,N_3480);
and U7418 (N_7418,N_2429,N_37);
or U7419 (N_7419,N_1459,N_2530);
and U7420 (N_7420,N_1168,N_4491);
and U7421 (N_7421,N_3322,N_2832);
and U7422 (N_7422,N_5712,N_3949);
or U7423 (N_7423,N_5577,N_529);
or U7424 (N_7424,N_5100,N_1210);
or U7425 (N_7425,N_2702,N_1019);
xnor U7426 (N_7426,N_4135,N_2841);
or U7427 (N_7427,N_909,N_5750);
and U7428 (N_7428,N_873,N_649);
or U7429 (N_7429,N_5137,N_1305);
or U7430 (N_7430,N_2847,N_2173);
nand U7431 (N_7431,N_5741,N_2586);
nand U7432 (N_7432,N_1390,N_1627);
and U7433 (N_7433,N_2485,N_2886);
xnor U7434 (N_7434,N_5921,N_4013);
and U7435 (N_7435,N_5421,N_4764);
or U7436 (N_7436,N_3318,N_5515);
or U7437 (N_7437,N_4150,N_2165);
nor U7438 (N_7438,N_87,N_3160);
or U7439 (N_7439,N_3212,N_541);
nand U7440 (N_7440,N_5898,N_475);
or U7441 (N_7441,N_5572,N_5251);
nor U7442 (N_7442,N_3462,N_5149);
nor U7443 (N_7443,N_2690,N_4880);
nor U7444 (N_7444,N_1214,N_1909);
xor U7445 (N_7445,N_641,N_2073);
nand U7446 (N_7446,N_4061,N_1847);
and U7447 (N_7447,N_292,N_4940);
or U7448 (N_7448,N_2193,N_4427);
and U7449 (N_7449,N_3504,N_3137);
and U7450 (N_7450,N_5951,N_2329);
and U7451 (N_7451,N_3780,N_4035);
and U7452 (N_7452,N_45,N_2399);
xor U7453 (N_7453,N_5041,N_3139);
or U7454 (N_7454,N_801,N_2395);
nand U7455 (N_7455,N_432,N_4631);
and U7456 (N_7456,N_5845,N_2313);
xor U7457 (N_7457,N_106,N_2112);
or U7458 (N_7458,N_1785,N_2952);
nand U7459 (N_7459,N_3909,N_3648);
nor U7460 (N_7460,N_1500,N_4418);
or U7461 (N_7461,N_3130,N_5511);
nand U7462 (N_7462,N_4584,N_2434);
xnor U7463 (N_7463,N_502,N_717);
and U7464 (N_7464,N_997,N_1334);
xor U7465 (N_7465,N_172,N_1173);
nand U7466 (N_7466,N_1545,N_1319);
nand U7467 (N_7467,N_5807,N_3912);
or U7468 (N_7468,N_1561,N_1920);
or U7469 (N_7469,N_1038,N_3176);
or U7470 (N_7470,N_899,N_3401);
nand U7471 (N_7471,N_3393,N_4662);
xnor U7472 (N_7472,N_1583,N_3172);
nor U7473 (N_7473,N_5429,N_5452);
nand U7474 (N_7474,N_3730,N_2025);
nor U7475 (N_7475,N_3340,N_4542);
and U7476 (N_7476,N_3442,N_2900);
nand U7477 (N_7477,N_2252,N_4026);
xnor U7478 (N_7478,N_3956,N_4699);
and U7479 (N_7479,N_426,N_173);
nor U7480 (N_7480,N_3473,N_3605);
nand U7481 (N_7481,N_3801,N_5838);
nor U7482 (N_7482,N_60,N_2895);
or U7483 (N_7483,N_388,N_1037);
nand U7484 (N_7484,N_1176,N_5814);
and U7485 (N_7485,N_2050,N_3565);
nand U7486 (N_7486,N_5166,N_1712);
and U7487 (N_7487,N_4693,N_5565);
xor U7488 (N_7488,N_145,N_5908);
xnor U7489 (N_7489,N_3777,N_514);
nand U7490 (N_7490,N_877,N_5943);
and U7491 (N_7491,N_4222,N_2248);
and U7492 (N_7492,N_5483,N_4781);
xnor U7493 (N_7493,N_4678,N_4776);
and U7494 (N_7494,N_1764,N_4874);
nand U7495 (N_7495,N_3141,N_2090);
or U7496 (N_7496,N_2518,N_39);
and U7497 (N_7497,N_101,N_2171);
xnor U7498 (N_7498,N_2983,N_1389);
nand U7499 (N_7499,N_4670,N_2458);
xnor U7500 (N_7500,N_3000,N_951);
nand U7501 (N_7501,N_3452,N_5822);
or U7502 (N_7502,N_769,N_3728);
nand U7503 (N_7503,N_3699,N_3463);
xor U7504 (N_7504,N_5329,N_2381);
nand U7505 (N_7505,N_4126,N_5263);
or U7506 (N_7506,N_5354,N_5196);
nand U7507 (N_7507,N_2380,N_3536);
nand U7508 (N_7508,N_4793,N_4333);
and U7509 (N_7509,N_325,N_5091);
nand U7510 (N_7510,N_683,N_2134);
xor U7511 (N_7511,N_631,N_4031);
and U7512 (N_7512,N_2499,N_4356);
nand U7513 (N_7513,N_2200,N_1207);
xor U7514 (N_7514,N_406,N_2664);
or U7515 (N_7515,N_4303,N_1638);
nand U7516 (N_7516,N_587,N_5387);
xnor U7517 (N_7517,N_532,N_5642);
nor U7518 (N_7518,N_1410,N_2896);
nand U7519 (N_7519,N_5125,N_5163);
and U7520 (N_7520,N_981,N_5656);
nand U7521 (N_7521,N_5184,N_1264);
xnor U7522 (N_7522,N_1463,N_3291);
nand U7523 (N_7523,N_5247,N_5086);
or U7524 (N_7524,N_838,N_4184);
nand U7525 (N_7525,N_4095,N_1165);
nand U7526 (N_7526,N_5000,N_2833);
nand U7527 (N_7527,N_4443,N_2103);
nor U7528 (N_7528,N_5209,N_3633);
and U7529 (N_7529,N_1400,N_226);
nand U7530 (N_7530,N_3809,N_3532);
or U7531 (N_7531,N_1874,N_2948);
and U7532 (N_7532,N_1160,N_1428);
nand U7533 (N_7533,N_2546,N_4515);
nor U7534 (N_7534,N_155,N_1728);
xnor U7535 (N_7535,N_433,N_1884);
nor U7536 (N_7536,N_5690,N_5855);
or U7537 (N_7537,N_4894,N_255);
xnor U7538 (N_7538,N_3623,N_5324);
and U7539 (N_7539,N_983,N_1308);
or U7540 (N_7540,N_722,N_4775);
xnor U7541 (N_7541,N_5887,N_2557);
and U7542 (N_7542,N_3201,N_559);
nor U7543 (N_7543,N_2275,N_1848);
nand U7544 (N_7544,N_732,N_3175);
xnor U7545 (N_7545,N_471,N_108);
nor U7546 (N_7546,N_2737,N_56);
or U7547 (N_7547,N_3621,N_2623);
or U7548 (N_7548,N_4536,N_1681);
xor U7549 (N_7549,N_3358,N_3084);
xor U7550 (N_7550,N_1220,N_3244);
nor U7551 (N_7551,N_1227,N_3710);
xor U7552 (N_7552,N_5029,N_357);
nand U7553 (N_7553,N_1403,N_906);
nand U7554 (N_7554,N_4033,N_1100);
nor U7555 (N_7555,N_1938,N_1614);
xor U7556 (N_7556,N_1036,N_2908);
and U7557 (N_7557,N_3384,N_1436);
nor U7558 (N_7558,N_823,N_5882);
or U7559 (N_7559,N_3682,N_4732);
xnor U7560 (N_7560,N_2018,N_2048);
nand U7561 (N_7561,N_4709,N_114);
nor U7562 (N_7562,N_4513,N_2438);
or U7563 (N_7563,N_2464,N_5011);
and U7564 (N_7564,N_3435,N_2707);
or U7565 (N_7565,N_2298,N_4086);
xnor U7566 (N_7566,N_1244,N_862);
or U7567 (N_7567,N_2854,N_4700);
or U7568 (N_7568,N_4707,N_5894);
xnor U7569 (N_7569,N_13,N_807);
xnor U7570 (N_7570,N_2177,N_5397);
nor U7571 (N_7571,N_3086,N_4406);
xor U7572 (N_7572,N_4722,N_4461);
and U7573 (N_7573,N_4572,N_5495);
nor U7574 (N_7574,N_5926,N_3370);
and U7575 (N_7575,N_2779,N_83);
xnor U7576 (N_7576,N_1664,N_2991);
nor U7577 (N_7577,N_3642,N_2560);
xor U7578 (N_7578,N_3573,N_2662);
and U7579 (N_7579,N_4922,N_890);
xnor U7580 (N_7580,N_3302,N_2397);
nand U7581 (N_7581,N_3148,N_4854);
or U7582 (N_7582,N_5927,N_2057);
or U7583 (N_7583,N_4806,N_4205);
or U7584 (N_7584,N_4617,N_3336);
nand U7585 (N_7585,N_4190,N_2366);
xor U7586 (N_7586,N_1556,N_610);
xor U7587 (N_7587,N_1456,N_2489);
xnor U7588 (N_7588,N_3014,N_2121);
and U7589 (N_7589,N_5719,N_3670);
and U7590 (N_7590,N_4568,N_4950);
nor U7591 (N_7591,N_3306,N_3540);
and U7592 (N_7592,N_2981,N_5350);
or U7593 (N_7593,N_760,N_3127);
xor U7594 (N_7594,N_695,N_1691);
and U7595 (N_7595,N_5407,N_3734);
and U7596 (N_7596,N_1418,N_5861);
nand U7597 (N_7597,N_2300,N_27);
xor U7598 (N_7598,N_2465,N_3616);
nor U7599 (N_7599,N_4051,N_2660);
or U7600 (N_7600,N_5967,N_669);
xnor U7601 (N_7601,N_3474,N_2413);
xnor U7602 (N_7602,N_3385,N_4447);
xor U7603 (N_7603,N_1509,N_5093);
xor U7604 (N_7604,N_1421,N_4552);
xnor U7605 (N_7605,N_169,N_253);
nand U7606 (N_7606,N_1457,N_5449);
nand U7607 (N_7607,N_2299,N_1420);
xnor U7608 (N_7608,N_645,N_3615);
or U7609 (N_7609,N_3529,N_5665);
or U7610 (N_7610,N_3305,N_4571);
and U7611 (N_7611,N_460,N_4425);
xnor U7612 (N_7612,N_1158,N_2761);
xnor U7613 (N_7613,N_1183,N_1765);
nor U7614 (N_7614,N_2699,N_3146);
nor U7615 (N_7615,N_5942,N_915);
xor U7616 (N_7616,N_2602,N_4735);
xor U7617 (N_7617,N_1686,N_5075);
nand U7618 (N_7618,N_1248,N_5313);
xor U7619 (N_7619,N_1313,N_5622);
and U7620 (N_7620,N_391,N_844);
xnor U7621 (N_7621,N_400,N_3418);
nor U7622 (N_7622,N_1232,N_2357);
or U7623 (N_7623,N_184,N_4811);
and U7624 (N_7624,N_5232,N_929);
nand U7625 (N_7625,N_4242,N_2584);
xnor U7626 (N_7626,N_4320,N_4314);
nand U7627 (N_7627,N_1496,N_3906);
or U7628 (N_7628,N_2052,N_1506);
or U7629 (N_7629,N_2227,N_693);
and U7630 (N_7630,N_2360,N_3794);
xnor U7631 (N_7631,N_582,N_709);
xor U7632 (N_7632,N_3353,N_2140);
and U7633 (N_7633,N_5888,N_718);
nand U7634 (N_7634,N_1927,N_3444);
and U7635 (N_7635,N_5500,N_2671);
and U7636 (N_7636,N_5736,N_2124);
nand U7637 (N_7637,N_5770,N_3859);
and U7638 (N_7638,N_1611,N_2923);
nand U7639 (N_7639,N_323,N_3412);
and U7640 (N_7640,N_5756,N_3880);
and U7641 (N_7641,N_3381,N_2827);
xor U7642 (N_7642,N_2487,N_180);
xor U7643 (N_7643,N_1291,N_5977);
or U7644 (N_7644,N_4734,N_1192);
and U7645 (N_7645,N_3154,N_2831);
xnor U7646 (N_7646,N_18,N_4186);
xor U7647 (N_7647,N_2451,N_1075);
nand U7648 (N_7648,N_3117,N_2724);
nor U7649 (N_7649,N_1558,N_3899);
and U7650 (N_7650,N_4913,N_3115);
or U7651 (N_7651,N_3355,N_5892);
xnor U7652 (N_7652,N_5040,N_1304);
or U7653 (N_7653,N_3106,N_4408);
xor U7654 (N_7654,N_3158,N_1455);
nand U7655 (N_7655,N_2698,N_3138);
xnor U7656 (N_7656,N_4674,N_2800);
nor U7657 (N_7657,N_2958,N_3874);
and U7658 (N_7658,N_2042,N_3693);
xor U7659 (N_7659,N_5654,N_4497);
or U7660 (N_7660,N_3684,N_247);
and U7661 (N_7661,N_4855,N_968);
and U7662 (N_7662,N_2795,N_2943);
or U7663 (N_7663,N_1004,N_2344);
nand U7664 (N_7664,N_2913,N_1961);
or U7665 (N_7665,N_417,N_523);
xor U7666 (N_7666,N_1924,N_5230);
or U7667 (N_7667,N_3460,N_3481);
xnor U7668 (N_7668,N_5962,N_885);
and U7669 (N_7669,N_427,N_690);
or U7670 (N_7670,N_5068,N_3132);
and U7671 (N_7671,N_4772,N_5099);
nor U7672 (N_7672,N_431,N_3110);
and U7673 (N_7673,N_4269,N_4264);
nand U7674 (N_7674,N_4030,N_3165);
and U7675 (N_7675,N_2115,N_5794);
and U7676 (N_7676,N_1887,N_4505);
nand U7677 (N_7677,N_5795,N_689);
or U7678 (N_7678,N_458,N_4799);
nor U7679 (N_7679,N_3398,N_3060);
xnor U7680 (N_7680,N_4316,N_3837);
xnor U7681 (N_7681,N_1105,N_1193);
and U7682 (N_7682,N_2755,N_2372);
xor U7683 (N_7683,N_1733,N_2802);
or U7684 (N_7684,N_1846,N_4761);
or U7685 (N_7685,N_2942,N_2994);
and U7686 (N_7686,N_606,N_188);
nand U7687 (N_7687,N_3191,N_1935);
and U7688 (N_7688,N_386,N_2246);
xnor U7689 (N_7689,N_5382,N_2135);
nor U7690 (N_7690,N_1376,N_3224);
or U7691 (N_7691,N_3069,N_3680);
and U7692 (N_7692,N_4750,N_2230);
nor U7693 (N_7693,N_5320,N_920);
nor U7694 (N_7694,N_2931,N_81);
nor U7695 (N_7695,N_836,N_4288);
and U7696 (N_7696,N_5422,N_3672);
xnor U7697 (N_7697,N_3736,N_197);
nand U7698 (N_7698,N_4021,N_4381);
and U7699 (N_7699,N_0,N_4635);
and U7700 (N_7700,N_4383,N_1350);
xnor U7701 (N_7701,N_5053,N_864);
or U7702 (N_7702,N_3403,N_2422);
xnor U7703 (N_7703,N_5849,N_5832);
xor U7704 (N_7704,N_4153,N_2532);
xnor U7705 (N_7705,N_1358,N_4877);
nand U7706 (N_7706,N_966,N_3469);
xor U7707 (N_7707,N_564,N_2409);
nor U7708 (N_7708,N_3278,N_804);
or U7709 (N_7709,N_3806,N_1331);
or U7710 (N_7710,N_3790,N_5005);
and U7711 (N_7711,N_4860,N_5636);
nand U7712 (N_7712,N_787,N_3868);
nand U7713 (N_7713,N_1345,N_3908);
or U7714 (N_7714,N_2067,N_534);
nand U7715 (N_7715,N_4037,N_5187);
nand U7716 (N_7716,N_1707,N_4109);
or U7717 (N_7717,N_5489,N_5297);
or U7718 (N_7718,N_4753,N_73);
nand U7719 (N_7719,N_1127,N_2296);
nand U7720 (N_7720,N_2829,N_4986);
nand U7721 (N_7721,N_755,N_3002);
and U7722 (N_7722,N_2032,N_2453);
nand U7723 (N_7723,N_157,N_3872);
nand U7724 (N_7724,N_5766,N_2823);
and U7725 (N_7725,N_5635,N_3210);
nor U7726 (N_7726,N_405,N_135);
or U7727 (N_7727,N_3373,N_2734);
nor U7728 (N_7728,N_334,N_138);
xor U7729 (N_7729,N_2070,N_449);
nor U7730 (N_7730,N_5045,N_3034);
nor U7731 (N_7731,N_3818,N_5363);
xnor U7732 (N_7732,N_1679,N_2626);
nor U7733 (N_7733,N_3062,N_219);
and U7734 (N_7734,N_232,N_1488);
nand U7735 (N_7735,N_566,N_5751);
nor U7736 (N_7736,N_2244,N_5681);
or U7737 (N_7737,N_5176,N_1179);
nor U7738 (N_7738,N_5513,N_5724);
and U7739 (N_7739,N_1526,N_5688);
nand U7740 (N_7740,N_3987,N_5778);
and U7741 (N_7741,N_5605,N_1124);
and U7742 (N_7742,N_1351,N_511);
xor U7743 (N_7743,N_3838,N_4415);
xnor U7744 (N_7744,N_4050,N_4435);
xnor U7745 (N_7745,N_2062,N_4645);
xor U7746 (N_7746,N_224,N_416);
nor U7747 (N_7747,N_5072,N_3705);
nand U7748 (N_7748,N_2918,N_987);
xor U7749 (N_7749,N_797,N_5401);
or U7750 (N_7750,N_272,N_380);
or U7751 (N_7751,N_4549,N_1859);
nor U7752 (N_7752,N_5497,N_5131);
xnor U7753 (N_7753,N_4339,N_1630);
nand U7754 (N_7754,N_4576,N_3849);
nor U7755 (N_7755,N_1892,N_1792);
nand U7756 (N_7756,N_1536,N_1644);
nand U7757 (N_7757,N_100,N_526);
nand U7758 (N_7758,N_3601,N_2998);
or U7759 (N_7759,N_5884,N_1002);
and U7760 (N_7760,N_2256,N_3434);
and U7761 (N_7761,N_3022,N_4881);
xor U7762 (N_7762,N_2750,N_5014);
nand U7763 (N_7763,N_1685,N_1440);
or U7764 (N_7764,N_3747,N_3666);
and U7765 (N_7765,N_2053,N_2195);
or U7766 (N_7766,N_1450,N_5269);
xnor U7767 (N_7767,N_5878,N_2987);
or U7768 (N_7768,N_1274,N_4042);
nor U7769 (N_7769,N_3335,N_200);
nand U7770 (N_7770,N_3522,N_2637);
nand U7771 (N_7771,N_3944,N_2020);
xor U7772 (N_7772,N_2840,N_2142);
nor U7773 (N_7773,N_4632,N_3759);
and U7774 (N_7774,N_5566,N_4728);
and U7775 (N_7775,N_4492,N_3492);
xnor U7776 (N_7776,N_4977,N_2711);
nand U7777 (N_7777,N_2312,N_4020);
nand U7778 (N_7778,N_5012,N_5233);
nor U7779 (N_7779,N_79,N_5357);
nand U7780 (N_7780,N_500,N_4319);
or U7781 (N_7781,N_5584,N_462);
nor U7782 (N_7782,N_4992,N_5038);
and U7783 (N_7783,N_4256,N_4800);
nand U7784 (N_7784,N_3688,N_25);
nor U7785 (N_7785,N_2871,N_4145);
and U7786 (N_7786,N_4845,N_5754);
or U7787 (N_7787,N_5866,N_1891);
xnor U7788 (N_7788,N_1042,N_661);
or U7789 (N_7789,N_4653,N_1284);
xor U7790 (N_7790,N_3143,N_2323);
nor U7791 (N_7791,N_2866,N_5023);
or U7792 (N_7792,N_5370,N_2951);
nor U7793 (N_7793,N_2118,N_2757);
nand U7794 (N_7794,N_2616,N_1788);
or U7795 (N_7795,N_1328,N_4343);
or U7796 (N_7796,N_2605,N_579);
nor U7797 (N_7797,N_3651,N_5126);
nor U7798 (N_7798,N_2334,N_392);
nor U7799 (N_7799,N_701,N_1871);
and U7800 (N_7800,N_3272,N_4257);
xor U7801 (N_7801,N_181,N_5586);
nand U7802 (N_7802,N_3509,N_5816);
and U7803 (N_7803,N_3968,N_5858);
nor U7804 (N_7804,N_793,N_1600);
xnor U7805 (N_7805,N_2093,N_3701);
or U7806 (N_7806,N_5268,N_456);
nand U7807 (N_7807,N_1031,N_3314);
nor U7808 (N_7808,N_4102,N_5543);
or U7809 (N_7809,N_2358,N_1718);
xnor U7810 (N_7810,N_5950,N_4556);
or U7811 (N_7811,N_682,N_3841);
or U7812 (N_7812,N_5485,N_1835);
nand U7813 (N_7813,N_4322,N_875);
nor U7814 (N_7814,N_4960,N_2929);
and U7815 (N_7815,N_2768,N_5146);
and U7816 (N_7816,N_2767,N_938);
nor U7817 (N_7817,N_2152,N_2470);
xor U7818 (N_7818,N_1714,N_5940);
nor U7819 (N_7819,N_1513,N_5747);
nand U7820 (N_7820,N_5906,N_4918);
nor U7821 (N_7821,N_5663,N_5116);
nand U7822 (N_7822,N_2742,N_2796);
or U7823 (N_7823,N_5346,N_1065);
nand U7824 (N_7824,N_1867,N_1113);
or U7825 (N_7825,N_3290,N_2606);
nor U7826 (N_7826,N_3311,N_1929);
or U7827 (N_7827,N_2635,N_2031);
nor U7828 (N_7828,N_4879,N_5571);
xnor U7829 (N_7829,N_4247,N_4646);
and U7830 (N_7830,N_2803,N_1855);
and U7831 (N_7831,N_3958,N_1011);
xor U7832 (N_7832,N_2588,N_4784);
nand U7833 (N_7833,N_4837,N_3019);
xor U7834 (N_7834,N_5339,N_548);
nand U7835 (N_7835,N_5544,N_3563);
nand U7836 (N_7836,N_3941,N_3010);
nor U7837 (N_7837,N_805,N_4610);
and U7838 (N_7838,N_625,N_989);
and U7839 (N_7839,N_4498,N_437);
or U7840 (N_7840,N_4948,N_5420);
nand U7841 (N_7841,N_1541,N_1833);
nor U7842 (N_7842,N_1398,N_3555);
or U7843 (N_7843,N_4683,N_4754);
xnor U7844 (N_7844,N_3151,N_3179);
xor U7845 (N_7845,N_688,N_236);
nand U7846 (N_7846,N_5034,N_2549);
or U7847 (N_7847,N_3772,N_799);
and U7848 (N_7848,N_3791,N_3544);
nor U7849 (N_7849,N_331,N_3895);
xnor U7850 (N_7850,N_5448,N_4929);
and U7851 (N_7851,N_1034,N_1682);
xor U7852 (N_7852,N_1978,N_4752);
or U7853 (N_7853,N_1215,N_1618);
and U7854 (N_7854,N_1194,N_895);
or U7855 (N_7855,N_3631,N_4386);
and U7856 (N_7856,N_2599,N_4174);
xor U7857 (N_7857,N_4555,N_578);
nor U7858 (N_7858,N_2980,N_3588);
or U7859 (N_7859,N_5567,N_3255);
xnor U7860 (N_7860,N_1254,N_4394);
nor U7861 (N_7861,N_4073,N_3247);
or U7862 (N_7862,N_5728,N_1402);
nor U7863 (N_7863,N_4410,N_4946);
and U7864 (N_7864,N_4173,N_618);
or U7865 (N_7865,N_2197,N_3293);
xnor U7866 (N_7866,N_1324,N_3989);
or U7867 (N_7867,N_186,N_5781);
and U7868 (N_7868,N_5013,N_2932);
or U7869 (N_7869,N_3295,N_3203);
xor U7870 (N_7870,N_2950,N_4654);
nor U7871 (N_7871,N_1829,N_5471);
nand U7872 (N_7872,N_1404,N_2089);
nand U7873 (N_7873,N_1503,N_5985);
and U7874 (N_7874,N_5132,N_4560);
nand U7875 (N_7875,N_5162,N_2682);
nor U7876 (N_7876,N_4963,N_251);
xor U7877 (N_7877,N_834,N_2510);
nor U7878 (N_7878,N_1534,N_2209);
xor U7879 (N_7879,N_3850,N_5755);
xor U7880 (N_7880,N_3134,N_3914);
xnor U7881 (N_7881,N_3167,N_1379);
nor U7882 (N_7882,N_4236,N_4726);
xnor U7883 (N_7883,N_3731,N_3810);
nand U7884 (N_7884,N_5332,N_2596);
or U7885 (N_7885,N_3905,N_3797);
xnor U7886 (N_7886,N_5380,N_2006);
nand U7887 (N_7887,N_2665,N_1836);
or U7888 (N_7888,N_5279,N_3277);
or U7889 (N_7889,N_288,N_3227);
or U7890 (N_7890,N_4093,N_1484);
or U7891 (N_7891,N_750,N_735);
nor U7892 (N_7892,N_1610,N_3457);
and U7893 (N_7893,N_1391,N_4371);
xnor U7894 (N_7894,N_3309,N_3243);
nor U7895 (N_7895,N_4723,N_2810);
nor U7896 (N_7896,N_3595,N_2964);
or U7897 (N_7897,N_4332,N_931);
and U7898 (N_7898,N_907,N_3016);
or U7899 (N_7899,N_973,N_5369);
nor U7900 (N_7900,N_359,N_3489);
nor U7901 (N_7901,N_5225,N_2486);
or U7902 (N_7902,N_279,N_5569);
or U7903 (N_7903,N_4301,N_2265);
xnor U7904 (N_7904,N_5240,N_2844);
nor U7905 (N_7905,N_2421,N_1814);
nand U7906 (N_7906,N_2887,N_1493);
nand U7907 (N_7907,N_2610,N_5214);
nand U7908 (N_7908,N_5216,N_4357);
and U7909 (N_7909,N_2419,N_5815);
or U7910 (N_7910,N_5561,N_210);
xnor U7911 (N_7911,N_5486,N_2621);
nor U7912 (N_7912,N_586,N_4067);
and U7913 (N_7913,N_3569,N_4991);
and U7914 (N_7914,N_1840,N_2514);
or U7915 (N_7915,N_2107,N_4099);
and U7916 (N_7916,N_3225,N_4902);
nand U7917 (N_7917,N_1290,N_589);
and U7918 (N_7918,N_5423,N_1361);
or U7919 (N_7919,N_1589,N_3972);
nor U7920 (N_7920,N_1787,N_4689);
or U7921 (N_7921,N_5739,N_4246);
and U7922 (N_7922,N_613,N_1590);
nor U7923 (N_7923,N_1702,N_2797);
and U7924 (N_7924,N_4600,N_5027);
nand U7925 (N_7925,N_1912,N_1008);
nand U7926 (N_7926,N_3553,N_4903);
or U7927 (N_7927,N_2182,N_4730);
nor U7928 (N_7928,N_3622,N_5738);
nand U7929 (N_7929,N_970,N_4144);
xnor U7930 (N_7930,N_2440,N_346);
and U7931 (N_7931,N_3121,N_719);
nand U7932 (N_7932,N_4367,N_4820);
xnor U7933 (N_7933,N_3657,N_2493);
xnor U7934 (N_7934,N_454,N_1757);
nor U7935 (N_7935,N_4812,N_4259);
nor U7936 (N_7936,N_367,N_4390);
and U7937 (N_7937,N_2047,N_1014);
nor U7938 (N_7938,N_5008,N_1494);
or U7939 (N_7939,N_1258,N_4485);
nor U7940 (N_7940,N_884,N_3208);
or U7941 (N_7941,N_4506,N_2506);
nor U7942 (N_7942,N_1178,N_4882);
xor U7943 (N_7943,N_1237,N_2641);
xnor U7944 (N_7944,N_2190,N_2581);
nor U7945 (N_7945,N_663,N_2947);
xor U7946 (N_7946,N_1843,N_189);
and U7947 (N_7947,N_2225,N_2287);
or U7948 (N_7948,N_54,N_5723);
xnor U7949 (N_7949,N_2600,N_324);
nand U7950 (N_7950,N_4299,N_4231);
xor U7951 (N_7951,N_785,N_4636);
or U7952 (N_7952,N_1801,N_478);
xor U7953 (N_7953,N_4238,N_1983);
and U7954 (N_7954,N_3021,N_3901);
or U7955 (N_7955,N_2087,N_3237);
or U7956 (N_7956,N_3848,N_264);
nand U7957 (N_7957,N_5122,N_153);
or U7958 (N_7958,N_2270,N_5783);
nor U7959 (N_7959,N_3913,N_1948);
nor U7960 (N_7960,N_3283,N_3);
xnor U7961 (N_7961,N_2719,N_1721);
xnor U7962 (N_7962,N_4688,N_4708);
or U7963 (N_7963,N_2271,N_4982);
nand U7964 (N_7964,N_2442,N_866);
nand U7965 (N_7965,N_2740,N_4097);
xnor U7966 (N_7966,N_4293,N_2043);
nor U7967 (N_7967,N_595,N_4558);
or U7968 (N_7968,N_3354,N_3991);
xor U7969 (N_7969,N_3665,N_928);
nor U7970 (N_7970,N_61,N_1318);
nor U7971 (N_7971,N_4981,N_962);
nand U7972 (N_7972,N_1782,N_3811);
nor U7973 (N_7973,N_4720,N_3501);
nand U7974 (N_7974,N_5707,N_2644);
nor U7975 (N_7975,N_5760,N_5305);
or U7976 (N_7976,N_4494,N_1140);
and U7977 (N_7977,N_3596,N_5999);
and U7978 (N_7978,N_1773,N_1219);
xnor U7979 (N_7979,N_4787,N_4194);
nand U7980 (N_7980,N_5490,N_5762);
nand U7981 (N_7981,N_3495,N_1239);
nand U7982 (N_7982,N_2927,N_2555);
nand U7983 (N_7983,N_4224,N_2219);
or U7984 (N_7984,N_3503,N_2651);
nand U7985 (N_7985,N_2254,N_5159);
or U7986 (N_7986,N_1187,N_4548);
or U7987 (N_7987,N_1152,N_3142);
xnor U7988 (N_7988,N_376,N_5334);
or U7989 (N_7989,N_3635,N_952);
nand U7990 (N_7990,N_1216,N_851);
and U7991 (N_7991,N_4132,N_4240);
nand U7992 (N_7992,N_451,N_2302);
nand U7993 (N_7993,N_4085,N_3892);
nor U7994 (N_7994,N_2348,N_1472);
or U7995 (N_7995,N_3694,N_3055);
xnor U7996 (N_7996,N_4524,N_4160);
or U7997 (N_7997,N_3327,N_4268);
nor U7998 (N_7998,N_5768,N_2101);
xnor U7999 (N_7999,N_2990,N_2308);
nand U8000 (N_8000,N_3592,N_1700);
or U8001 (N_8001,N_4824,N_2534);
nor U8002 (N_8002,N_806,N_2144);
xnor U8003 (N_8003,N_4996,N_1771);
and U8004 (N_8004,N_1231,N_1754);
nand U8005 (N_8005,N_1340,N_4107);
and U8006 (N_8006,N_358,N_2835);
nand U8007 (N_8007,N_3433,N_5173);
and U8008 (N_8008,N_3150,N_1953);
xnor U8009 (N_8009,N_1914,N_235);
or U8010 (N_8010,N_5282,N_3273);
or U8011 (N_8011,N_495,N_591);
or U8012 (N_8012,N_2468,N_5478);
nand U8013 (N_8013,N_2278,N_4458);
xnor U8014 (N_8014,N_2643,N_3719);
and U8015 (N_8015,N_4463,N_2306);
xnor U8016 (N_8016,N_571,N_687);
xor U8017 (N_8017,N_3920,N_5273);
or U8018 (N_8018,N_3546,N_4675);
or U8019 (N_8019,N_5560,N_2793);
nor U8020 (N_8020,N_5705,N_2752);
nor U8021 (N_8021,N_3530,N_3241);
or U8022 (N_8022,N_2113,N_82);
and U8023 (N_8023,N_2861,N_657);
or U8024 (N_8024,N_125,N_5169);
or U8025 (N_8025,N_665,N_2452);
xnor U8026 (N_8026,N_4733,N_2704);
nand U8027 (N_8027,N_3049,N_2292);
or U8028 (N_8028,N_4861,N_4431);
xor U8029 (N_8029,N_1750,N_3456);
xnor U8030 (N_8030,N_670,N_1736);
nor U8031 (N_8031,N_2748,N_5056);
or U8032 (N_8032,N_5883,N_614);
nand U8033 (N_8033,N_926,N_4919);
and U8034 (N_8034,N_5941,N_4286);
nand U8035 (N_8035,N_2259,N_3822);
xnor U8036 (N_8036,N_839,N_5418);
or U8037 (N_8037,N_1763,N_543);
nor U8038 (N_8038,N_607,N_4227);
xnor U8039 (N_8039,N_4011,N_5141);
xor U8040 (N_8040,N_950,N_4580);
nor U8041 (N_8041,N_3551,N_3246);
and U8042 (N_8042,N_1542,N_5252);
xor U8043 (N_8043,N_3576,N_753);
and U8044 (N_8044,N_2627,N_4294);
and U8045 (N_8045,N_4335,N_1293);
and U8046 (N_8046,N_5732,N_1966);
nor U8047 (N_8047,N_457,N_5982);
and U8048 (N_8048,N_5523,N_4161);
nor U8049 (N_8049,N_1834,N_3427);
or U8050 (N_8050,N_3525,N_4039);
and U8051 (N_8051,N_1013,N_2471);
and U8052 (N_8052,N_4159,N_4325);
xnor U8053 (N_8053,N_470,N_4002);
or U8054 (N_8054,N_1148,N_1781);
xnor U8055 (N_8055,N_5821,N_643);
or U8056 (N_8056,N_3866,N_1992);
and U8057 (N_8057,N_1680,N_4972);
or U8058 (N_8058,N_3638,N_5915);
nand U8059 (N_8059,N_4501,N_626);
nor U8060 (N_8060,N_4402,N_5296);
nand U8061 (N_8061,N_2127,N_5383);
or U8062 (N_8062,N_1748,N_5839);
or U8063 (N_8063,N_1885,N_1770);
or U8064 (N_8064,N_2930,N_636);
nor U8065 (N_8065,N_1620,N_675);
and U8066 (N_8066,N_3207,N_2694);
xor U8067 (N_8067,N_5077,N_3233);
and U8068 (N_8068,N_1139,N_4387);
xnor U8069 (N_8069,N_191,N_4336);
nor U8070 (N_8070,N_4234,N_5461);
xnor U8071 (N_8071,N_1112,N_4663);
or U8072 (N_8072,N_1675,N_337);
xor U8073 (N_8073,N_1119,N_4640);
or U8074 (N_8074,N_5156,N_1687);
xor U8075 (N_8075,N_1635,N_1490);
and U8076 (N_8076,N_524,N_4032);
nor U8077 (N_8077,N_5830,N_705);
or U8078 (N_8078,N_1975,N_3789);
xor U8079 (N_8079,N_3041,N_1347);
and U8080 (N_8080,N_3351,N_167);
nand U8081 (N_8081,N_1343,N_5205);
nand U8082 (N_8082,N_1645,N_3775);
and U8083 (N_8083,N_3073,N_4899);
nand U8084 (N_8084,N_2086,N_4798);
xnor U8085 (N_8085,N_1289,N_874);
and U8086 (N_8086,N_4084,N_4147);
or U8087 (N_8087,N_4466,N_2736);
or U8088 (N_8088,N_934,N_1174);
nor U8089 (N_8089,N_2130,N_20);
or U8090 (N_8090,N_3008,N_5633);
xnor U8091 (N_8091,N_1261,N_31);
and U8092 (N_8092,N_2905,N_2205);
and U8093 (N_8093,N_5646,N_2021);
xnor U8094 (N_8094,N_5944,N_2807);
or U8095 (N_8095,N_4318,N_3707);
nor U8096 (N_8096,N_2262,N_2017);
or U8097 (N_8097,N_3676,N_5875);
nand U8098 (N_8098,N_2237,N_5036);
xor U8099 (N_8099,N_218,N_3940);
and U8100 (N_8100,N_4380,N_746);
and U8101 (N_8101,N_5491,N_5850);
nand U8102 (N_8102,N_5776,N_3624);
and U8103 (N_8103,N_162,N_3584);
nor U8104 (N_8104,N_4068,N_632);
and U8105 (N_8105,N_5212,N_5956);
xnor U8106 (N_8106,N_1841,N_1998);
or U8107 (N_8107,N_5863,N_5248);
or U8108 (N_8108,N_4711,N_4122);
nor U8109 (N_8109,N_2319,N_5897);
and U8110 (N_8110,N_1768,N_159);
or U8111 (N_8111,N_4615,N_476);
nand U8112 (N_8112,N_3667,N_4843);
and U8113 (N_8113,N_4715,N_1804);
nor U8114 (N_8114,N_990,N_46);
nor U8115 (N_8115,N_1744,N_2445);
and U8116 (N_8116,N_777,N_2462);
or U8117 (N_8117,N_4027,N_2523);
xor U8118 (N_8118,N_2993,N_3917);
or U8119 (N_8119,N_2780,N_5308);
or U8120 (N_8120,N_2725,N_854);
xnor U8121 (N_8121,N_1460,N_4794);
or U8122 (N_8122,N_6,N_4518);
nand U8123 (N_8123,N_1657,N_4115);
nor U8124 (N_8124,N_3173,N_1406);
nor U8125 (N_8125,N_5536,N_5281);
nand U8126 (N_8126,N_1826,N_2756);
xnor U8127 (N_8127,N_5611,N_2587);
or U8128 (N_8128,N_4232,N_1325);
nand U8129 (N_8129,N_1722,N_2417);
xor U8130 (N_8130,N_5645,N_212);
or U8131 (N_8131,N_733,N_2816);
or U8132 (N_8132,N_3047,N_1769);
nand U8133 (N_8133,N_5138,N_5315);
xor U8134 (N_8134,N_3064,N_4000);
or U8135 (N_8135,N_2189,N_51);
nand U8136 (N_8136,N_1617,N_1608);
xor U8137 (N_8137,N_5106,N_5211);
xor U8138 (N_8138,N_2554,N_4096);
nand U8139 (N_8139,N_3349,N_4970);
xnor U8140 (N_8140,N_5154,N_424);
nor U8141 (N_8141,N_469,N_646);
and U8142 (N_8142,N_5356,N_419);
xor U8143 (N_8143,N_2137,N_751);
or U8144 (N_8144,N_2838,N_4304);
nand U8145 (N_8145,N_1429,N_350);
and U8146 (N_8146,N_3411,N_3858);
nor U8147 (N_8147,N_1527,N_4488);
or U8148 (N_8148,N_833,N_5625);
nor U8149 (N_8149,N_2033,N_5323);
nand U8150 (N_8150,N_5052,N_5322);
or U8151 (N_8151,N_3397,N_5709);
and U8152 (N_8152,N_2583,N_5913);
or U8153 (N_8153,N_1822,N_4423);
and U8154 (N_8154,N_1438,N_3792);
and U8155 (N_8155,N_2145,N_1795);
or U8156 (N_8156,N_2199,N_3359);
or U8157 (N_8157,N_5110,N_3129);
or U8158 (N_8158,N_867,N_5630);
or U8159 (N_8159,N_4570,N_5215);
nand U8160 (N_8160,N_3249,N_1584);
and U8161 (N_8161,N_738,N_1001);
and U8162 (N_8162,N_2398,N_547);
nor U8163 (N_8163,N_1648,N_3313);
xor U8164 (N_8164,N_35,N_1738);
xor U8165 (N_8165,N_5194,N_3955);
nand U8166 (N_8166,N_3419,N_2345);
or U8167 (N_8167,N_4007,N_1943);
nor U8168 (N_8168,N_3754,N_590);
xor U8169 (N_8169,N_2808,N_3617);
nor U8170 (N_8170,N_4074,N_3003);
and U8171 (N_8171,N_5964,N_1222);
or U8172 (N_8172,N_2249,N_1189);
or U8173 (N_8173,N_3804,N_1045);
or U8174 (N_8174,N_1588,N_490);
nand U8175 (N_8175,N_4817,N_5136);
or U8176 (N_8176,N_326,N_5119);
nor U8177 (N_8177,N_1893,N_1281);
xnor U8178 (N_8178,N_629,N_2812);
or U8179 (N_8179,N_5021,N_5498);
and U8180 (N_8180,N_4779,N_4207);
and U8181 (N_8181,N_1117,N_3669);
and U8182 (N_8182,N_411,N_1323);
and U8183 (N_8183,N_3541,N_2294);
xnor U8184 (N_8184,N_2106,N_3945);
xnor U8185 (N_8185,N_985,N_563);
nand U8186 (N_8186,N_666,N_1307);
nor U8187 (N_8187,N_2492,N_2276);
or U8188 (N_8188,N_127,N_4433);
or U8189 (N_8189,N_5833,N_3997);
nand U8190 (N_8190,N_1730,N_5742);
or U8191 (N_8191,N_1917,N_574);
xor U8192 (N_8192,N_685,N_5386);
and U8193 (N_8193,N_2264,N_5734);
nand U8194 (N_8194,N_2649,N_1989);
nand U8195 (N_8195,N_2920,N_4849);
or U8196 (N_8196,N_1735,N_2971);
xor U8197 (N_8197,N_344,N_4559);
xor U8198 (N_8198,N_599,N_3910);
xor U8199 (N_8199,N_5618,N_3020);
nand U8200 (N_8200,N_1411,N_660);
nand U8201 (N_8201,N_5562,N_5158);
nand U8202 (N_8202,N_594,N_3779);
nor U8203 (N_8203,N_993,N_3420);
and U8204 (N_8204,N_5437,N_5701);
or U8205 (N_8205,N_2028,N_1860);
xnor U8206 (N_8206,N_3898,N_3245);
nand U8207 (N_8207,N_5170,N_2325);
and U8208 (N_8208,N_3048,N_3678);
nor U8209 (N_8209,N_3159,N_301);
nand U8210 (N_8210,N_2873,N_3467);
nor U8211 (N_8211,N_4353,N_4565);
nor U8212 (N_8212,N_684,N_1567);
and U8213 (N_8213,N_1475,N_1710);
xnor U8214 (N_8214,N_2456,N_720);
or U8215 (N_8215,N_4872,N_4317);
nand U8216 (N_8216,N_2957,N_5111);
xnor U8217 (N_8217,N_4374,N_585);
and U8218 (N_8218,N_1654,N_5872);
xor U8219 (N_8219,N_4400,N_4424);
xnor U8220 (N_8220,N_1225,N_2002);
nand U8221 (N_8221,N_203,N_1473);
nor U8222 (N_8222,N_3855,N_1802);
nand U8223 (N_8223,N_1246,N_5777);
nor U8224 (N_8224,N_1499,N_2027);
nor U8225 (N_8225,N_3929,N_5104);
or U8226 (N_8226,N_3932,N_2538);
or U8227 (N_8227,N_2789,N_2331);
nor U8228 (N_8228,N_3080,N_572);
nand U8229 (N_8229,N_158,N_3882);
or U8230 (N_8230,N_4004,N_2117);
xnor U8231 (N_8231,N_221,N_276);
or U8232 (N_8232,N_5854,N_1628);
nor U8233 (N_8233,N_5451,N_1067);
or U8234 (N_8234,N_1875,N_565);
and U8235 (N_8235,N_2701,N_5960);
and U8236 (N_8236,N_1761,N_355);
or U8237 (N_8237,N_2412,N_5090);
and U8238 (N_8238,N_1962,N_5714);
nor U8239 (N_8239,N_748,N_4083);
or U8240 (N_8240,N_217,N_3634);
or U8241 (N_8241,N_2139,N_3156);
and U8242 (N_8242,N_464,N_604);
nor U8243 (N_8243,N_5234,N_1205);
xnor U8244 (N_8244,N_2007,N_835);
nand U8245 (N_8245,N_2368,N_3422);
nor U8246 (N_8246,N_1028,N_3267);
nor U8247 (N_8247,N_2562,N_2267);
xor U8248 (N_8248,N_466,N_166);
nand U8249 (N_8249,N_3324,N_271);
nand U8250 (N_8250,N_2088,N_447);
nand U8251 (N_8251,N_2435,N_1195);
nand U8252 (N_8252,N_229,N_3547);
and U8253 (N_8253,N_5588,N_674);
xnor U8254 (N_8254,N_305,N_3072);
nor U8255 (N_8255,N_4388,N_3147);
nor U8256 (N_8256,N_5818,N_1858);
nor U8257 (N_8257,N_4411,N_2749);
nor U8258 (N_8258,N_267,N_5039);
or U8259 (N_8259,N_4253,N_1799);
or U8260 (N_8260,N_652,N_3402);
or U8261 (N_8261,N_4546,N_4123);
xnor U8262 (N_8262,N_1209,N_4608);
xnor U8263 (N_8263,N_1613,N_3977);
or U8264 (N_8264,N_4740,N_954);
and U8265 (N_8265,N_2897,N_2318);
and U8266 (N_8266,N_3312,N_4596);
or U8267 (N_8267,N_4047,N_2233);
nand U8268 (N_8268,N_1955,N_5589);
nor U8269 (N_8269,N_488,N_2848);
xor U8270 (N_8270,N_1564,N_1659);
nor U8271 (N_8271,N_1716,N_86);
nor U8272 (N_8272,N_1048,N_3798);
xnor U8273 (N_8273,N_3865,N_5445);
nand U8274 (N_8274,N_3363,N_5197);
and U8275 (N_8275,N_2914,N_3450);
or U8276 (N_8276,N_2850,N_4478);
nor U8277 (N_8277,N_3181,N_3842);
nor U8278 (N_8278,N_5140,N_2433);
nor U8279 (N_8279,N_3686,N_246);
or U8280 (N_8280,N_3383,N_5272);
nand U8281 (N_8281,N_239,N_3609);
nor U8282 (N_8282,N_2684,N_4346);
or U8283 (N_8283,N_946,N_4541);
or U8284 (N_8284,N_5846,N_964);
xnor U8285 (N_8285,N_2578,N_1649);
or U8286 (N_8286,N_4352,N_2373);
or U8287 (N_8287,N_1959,N_4295);
nand U8288 (N_8288,N_2391,N_1359);
and U8289 (N_8289,N_1422,N_1918);
or U8290 (N_8290,N_1357,N_5285);
or U8291 (N_8291,N_3593,N_2524);
nand U8292 (N_8292,N_4613,N_2266);
or U8293 (N_8293,N_4701,N_1726);
and U8294 (N_8294,N_2157,N_1705);
nand U8295 (N_8295,N_1876,N_2273);
or U8296 (N_8296,N_3153,N_3820);
xnor U8297 (N_8297,N_4263,N_3262);
xnor U8298 (N_8298,N_2404,N_245);
nand U8299 (N_8299,N_4006,N_5804);
xor U8300 (N_8300,N_4875,N_2008);
xor U8301 (N_8301,N_1888,N_994);
xnor U8302 (N_8302,N_1512,N_4041);
or U8303 (N_8303,N_1928,N_583);
nor U8304 (N_8304,N_2674,N_5231);
nor U8305 (N_8305,N_4413,N_2170);
xor U8306 (N_8306,N_2965,N_5682);
xor U8307 (N_8307,N_5703,N_2921);
and U8308 (N_8308,N_4193,N_2424);
nand U8309 (N_8309,N_5336,N_5970);
and U8310 (N_8310,N_653,N_5456);
or U8311 (N_8311,N_1656,N_5464);
nand U8312 (N_8312,N_3556,N_5063);
nand U8313 (N_8313,N_902,N_3574);
or U8314 (N_8314,N_2785,N_4370);
or U8315 (N_8315,N_5699,N_4372);
or U8316 (N_8316,N_5527,N_5067);
or U8317 (N_8317,N_4171,N_89);
and U8318 (N_8318,N_3028,N_5384);
or U8319 (N_8319,N_2934,N_2559);
nand U8320 (N_8320,N_2191,N_4313);
nor U8321 (N_8321,N_4065,N_5148);
xnor U8322 (N_8322,N_5328,N_1482);
and U8323 (N_8323,N_2985,N_2369);
nor U8324 (N_8324,N_4204,N_5463);
xnor U8325 (N_8325,N_3526,N_3870);
or U8326 (N_8326,N_1218,N_2764);
nand U8327 (N_8327,N_2316,N_201);
nor U8328 (N_8328,N_853,N_638);
and U8329 (N_8329,N_5686,N_2159);
or U8330 (N_8330,N_703,N_3136);
or U8331 (N_8331,N_5740,N_637);
xnor U8332 (N_8332,N_4439,N_1169);
or U8333 (N_8333,N_4908,N_3646);
or U8334 (N_8334,N_742,N_4130);
nor U8335 (N_8335,N_4934,N_4305);
and U8336 (N_8336,N_1206,N_2340);
xnor U8337 (N_8337,N_540,N_4582);
or U8338 (N_8338,N_4152,N_3606);
and U8339 (N_8339,N_935,N_1976);
nor U8340 (N_8340,N_4156,N_4561);
nand U8341 (N_8341,N_5095,N_4605);
or U8342 (N_8342,N_1236,N_3282);
nand U8343 (N_8343,N_1476,N_4323);
or U8344 (N_8344,N_1315,N_1683);
nor U8345 (N_8345,N_1451,N_3202);
xor U8346 (N_8346,N_1688,N_1906);
nor U8347 (N_8347,N_1306,N_505);
xor U8348 (N_8348,N_5375,N_3308);
and U8349 (N_8349,N_5812,N_3722);
and U8350 (N_8350,N_5254,N_4975);
nor U8351 (N_8351,N_5727,N_294);
nand U8352 (N_8352,N_1278,N_2772);
nor U8353 (N_8353,N_3486,N_5613);
nor U8354 (N_8354,N_2214,N_1434);
nor U8355 (N_8355,N_439,N_3856);
nor U8356 (N_8356,N_5210,N_568);
xor U8357 (N_8357,N_2819,N_1865);
xnor U8358 (N_8358,N_163,N_5345);
nor U8359 (N_8359,N_3331,N_4217);
nand U8360 (N_8360,N_953,N_3927);
nand U8361 (N_8361,N_4260,N_3545);
nand U8362 (N_8362,N_3180,N_2075);
nor U8363 (N_8363,N_1245,N_5424);
nor U8364 (N_8364,N_2955,N_3518);
nor U8365 (N_8365,N_3960,N_5678);
nor U8366 (N_8366,N_126,N_4100);
and U8367 (N_8367,N_339,N_1522);
nor U8368 (N_8368,N_4682,N_1280);
nor U8369 (N_8369,N_3030,N_819);
nor U8370 (N_8370,N_453,N_1447);
nand U8371 (N_8371,N_845,N_5394);
xnor U8372 (N_8372,N_3417,N_1172);
and U8373 (N_8373,N_3071,N_1639);
nand U8374 (N_8374,N_775,N_1573);
xor U8375 (N_8375,N_2881,N_4351);
nand U8376 (N_8376,N_3050,N_1373);
nor U8377 (N_8377,N_2924,N_4197);
or U8378 (N_8378,N_4927,N_123);
nand U8379 (N_8379,N_5128,N_3183);
nand U8380 (N_8380,N_2277,N_942);
xnor U8381 (N_8381,N_2731,N_2553);
or U8382 (N_8382,N_5624,N_3488);
nor U8383 (N_8383,N_5289,N_2194);
or U8384 (N_8384,N_3093,N_3257);
or U8385 (N_8385,N_2595,N_2577);
nand U8386 (N_8386,N_2013,N_5547);
xnor U8387 (N_8387,N_5425,N_5643);
xnor U8388 (N_8388,N_4900,N_1676);
or U8389 (N_8389,N_1441,N_4276);
xor U8390 (N_8390,N_1270,N_258);
nand U8391 (N_8391,N_1982,N_302);
nor U8392 (N_8392,N_1431,N_4591);
and U8393 (N_8393,N_2321,N_2215);
nand U8394 (N_8394,N_4412,N_3817);
nand U8395 (N_8395,N_2091,N_704);
xor U8396 (N_8396,N_1729,N_4191);
or U8397 (N_8397,N_5853,N_329);
nand U8398 (N_8398,N_5600,N_5891);
or U8399 (N_8399,N_2505,N_2387);
and U8400 (N_8400,N_2680,N_410);
nor U8401 (N_8401,N_244,N_4008);
xnor U8402 (N_8402,N_1854,N_597);
nand U8403 (N_8403,N_758,N_3083);
nand U8404 (N_8404,N_5793,N_4029);
and U8405 (N_8405,N_1444,N_1407);
or U8406 (N_8406,N_2770,N_4289);
and U8407 (N_8407,N_4445,N_362);
xnor U8408 (N_8408,N_2888,N_908);
and U8409 (N_8409,N_1399,N_1372);
nand U8410 (N_8410,N_4486,N_2525);
and U8411 (N_8411,N_3980,N_1990);
xnor U8412 (N_8412,N_1366,N_2846);
nor U8413 (N_8413,N_2928,N_878);
xor U8414 (N_8414,N_3271,N_3543);
or U8415 (N_8415,N_4624,N_3135);
and U8416 (N_8416,N_1405,N_4638);
nor U8417 (N_8417,N_268,N_3928);
nand U8418 (N_8418,N_974,N_3382);
xor U8419 (N_8419,N_3270,N_1651);
or U8420 (N_8420,N_2129,N_1122);
xor U8421 (N_8421,N_4939,N_4243);
nor U8422 (N_8422,N_425,N_205);
and U8423 (N_8423,N_2436,N_3465);
and U8424 (N_8424,N_5876,N_1491);
nor U8425 (N_8425,N_2548,N_4983);
and U8426 (N_8426,N_2247,N_2153);
and U8427 (N_8427,N_2291,N_5877);
or U8428 (N_8428,N_1578,N_5784);
nand U8429 (N_8429,N_5638,N_2367);
nor U8430 (N_8430,N_5649,N_2437);
and U8431 (N_8431,N_5355,N_4487);
and U8432 (N_8432,N_3947,N_3238);
or U8433 (N_8433,N_5530,N_4857);
and U8434 (N_8434,N_4499,N_3934);
nand U8435 (N_8435,N_602,N_3310);
nand U8436 (N_8436,N_5055,N_1171);
and U8437 (N_8437,N_1517,N_5662);
or U8438 (N_8438,N_5679,N_4790);
nand U8439 (N_8439,N_608,N_2120);
and U8440 (N_8440,N_4639,N_3767);
xor U8441 (N_8441,N_3274,N_2961);
nand U8442 (N_8442,N_261,N_3891);
xor U8443 (N_8443,N_5267,N_5098);
and U8444 (N_8444,N_2208,N_9);
or U8445 (N_8445,N_2146,N_1818);
and U8446 (N_8446,N_3198,N_2517);
and U8447 (N_8447,N_4907,N_1282);
nor U8448 (N_8448,N_2542,N_198);
nand U8449 (N_8449,N_75,N_5459);
xnor U8450 (N_8450,N_3969,N_3276);
and U8451 (N_8451,N_8,N_4865);
nor U8452 (N_8452,N_5552,N_4583);
or U8453 (N_8453,N_925,N_1751);
xnor U8454 (N_8454,N_3407,N_4057);
nor U8455 (N_8455,N_713,N_869);
nand U8456 (N_8456,N_1692,N_5843);
nor U8457 (N_8457,N_2550,N_482);
nand U8458 (N_8458,N_316,N_4936);
nand U8459 (N_8459,N_3294,N_4557);
nand U8460 (N_8460,N_3190,N_2612);
nand U8461 (N_8461,N_5602,N_1520);
or U8462 (N_8462,N_1690,N_3155);
and U8463 (N_8463,N_3814,N_2891);
nand U8464 (N_8464,N_852,N_5270);
or U8465 (N_8465,N_2418,N_1775);
xor U8466 (N_8466,N_3975,N_4978);
nand U8467 (N_8467,N_2926,N_1699);
nor U8468 (N_8468,N_4091,N_3922);
nor U8469 (N_8469,N_5243,N_2394);
and U8470 (N_8470,N_222,N_3319);
or U8471 (N_8471,N_5181,N_2710);
and U8472 (N_8472,N_4510,N_5049);
or U8473 (N_8473,N_4185,N_2059);
nand U8474 (N_8474,N_3689,N_2416);
and U8475 (N_8475,N_2310,N_4606);
nor U8476 (N_8476,N_842,N_1540);
xnor U8477 (N_8477,N_3564,N_2406);
xnor U8478 (N_8478,N_4120,N_1263);
nor U8479 (N_8479,N_5934,N_3583);
or U8480 (N_8480,N_5304,N_5147);
xor U8481 (N_8481,N_5302,N_3557);
nand U8482 (N_8482,N_1669,N_4702);
nor U8483 (N_8483,N_3424,N_1279);
and U8484 (N_8484,N_202,N_3953);
or U8485 (N_8485,N_2198,N_3763);
xnor U8486 (N_8486,N_3475,N_4134);
and U8487 (N_8487,N_3723,N_85);
xor U8488 (N_8488,N_2689,N_965);
or U8489 (N_8489,N_5189,N_1057);
nor U8490 (N_8490,N_4551,N_5870);
nand U8491 (N_8491,N_601,N_347);
nand U8492 (N_8492,N_1322,N_409);
nor U8493 (N_8493,N_2516,N_560);
xor U8494 (N_8494,N_648,N_4666);
and U8495 (N_8495,N_3788,N_767);
or U8496 (N_8496,N_4814,N_3059);
nor U8497 (N_8497,N_5653,N_3748);
nand U8498 (N_8498,N_4398,N_1863);
nand U8499 (N_8499,N_841,N_3673);
nor U8500 (N_8500,N_4177,N_2343);
and U8501 (N_8501,N_3538,N_2213);
nand U8502 (N_8502,N_1314,N_4279);
and U8503 (N_8503,N_1741,N_584);
nand U8504 (N_8504,N_5199,N_5902);
nor U8505 (N_8505,N_1368,N_4911);
nand U8506 (N_8506,N_5868,N_374);
xnor U8507 (N_8507,N_3286,N_4063);
xnor U8508 (N_8508,N_2330,N_4941);
nand U8509 (N_8509,N_1397,N_4797);
xor U8510 (N_8510,N_2038,N_1817);
nand U8511 (N_8511,N_2460,N_3189);
and U8512 (N_8512,N_3839,N_4741);
nor U8513 (N_8513,N_4538,N_570);
and U8514 (N_8514,N_486,N_4360);
or U8515 (N_8515,N_5670,N_4836);
nand U8516 (N_8516,N_5161,N_2717);
xor U8517 (N_8517,N_308,N_3118);
nor U8518 (N_8518,N_2723,N_5580);
or U8519 (N_8519,N_5879,N_3907);
nor U8520 (N_8520,N_1153,N_1354);
xnor U8521 (N_8521,N_3468,N_4375);
nand U8522 (N_8522,N_3484,N_1908);
nand U8523 (N_8523,N_4278,N_510);
xnor U8524 (N_8524,N_3816,N_768);
or U8525 (N_8525,N_2778,N_4133);
or U8526 (N_8526,N_2119,N_2759);
nor U8527 (N_8527,N_2336,N_1055);
xnor U8528 (N_8528,N_4088,N_945);
xnor U8529 (N_8529,N_2563,N_5594);
and U8530 (N_8530,N_3360,N_4801);
xnor U8531 (N_8531,N_50,N_196);
and U8532 (N_8532,N_3376,N_1419);
or U8533 (N_8533,N_5761,N_1285);
xor U8534 (N_8534,N_2122,N_4884);
xnor U8535 (N_8535,N_4237,N_3347);
nand U8536 (N_8536,N_5482,N_2311);
and U8537 (N_8537,N_4496,N_3671);
xnor U8538 (N_8538,N_3860,N_3548);
nand U8539 (N_8539,N_3510,N_1697);
and U8540 (N_8540,N_4511,N_3996);
nand U8541 (N_8541,N_5744,N_1442);
nor U8542 (N_8542,N_1489,N_4482);
and U8543 (N_8543,N_220,N_2320);
and U8544 (N_8544,N_2163,N_3864);
xor U8545 (N_8545,N_5037,N_93);
nor U8546 (N_8546,N_436,N_4650);
xnor U8547 (N_8547,N_2076,N_1364);
or U8548 (N_8548,N_773,N_5592);
xor U8549 (N_8549,N_2074,N_680);
nor U8550 (N_8550,N_4075,N_4018);
nand U8551 (N_8551,N_1643,N_1970);
nor U8552 (N_8552,N_5446,N_3769);
nand U8553 (N_8553,N_5107,N_1352);
xor U8554 (N_8554,N_3935,N_881);
and U8555 (N_8555,N_2454,N_820);
nand U8556 (N_8556,N_2975,N_3776);
xnor U8557 (N_8557,N_1979,N_3591);
and U8558 (N_8558,N_4110,N_5772);
nand U8559 (N_8559,N_295,N_1454);
or U8560 (N_8560,N_3950,N_903);
nand U8561 (N_8561,N_2659,N_3873);
or U8562 (N_8562,N_5975,N_1941);
and U8563 (N_8563,N_830,N_3221);
nand U8564 (N_8564,N_863,N_5022);
nand U8565 (N_8565,N_1923,N_5713);
xnor U8566 (N_8566,N_3744,N_2408);
and U8567 (N_8567,N_4438,N_1118);
nor U8568 (N_8568,N_2383,N_1734);
nor U8569 (N_8569,N_3476,N_401);
xnor U8570 (N_8570,N_1130,N_1749);
and U8571 (N_8571,N_5311,N_1634);
nand U8572 (N_8572,N_1,N_3834);
and U8573 (N_8573,N_3123,N_817);
nor U8574 (N_8574,N_1384,N_3805);
nor U8575 (N_8575,N_956,N_1086);
nand U8576 (N_8576,N_3933,N_2105);
or U8577 (N_8577,N_353,N_501);
xnor U8578 (N_8578,N_2570,N_4834);
xnor U8579 (N_8579,N_4578,N_4657);
or U8580 (N_8580,N_4273,N_5178);
and U8581 (N_8581,N_5153,N_1087);
nor U8582 (N_8582,N_168,N_3535);
xnor U8583 (N_8583,N_4139,N_1963);
nand U8584 (N_8584,N_4602,N_3006);
or U8585 (N_8585,N_3458,N_4554);
or U8586 (N_8586,N_5503,N_4523);
nor U8587 (N_8587,N_3116,N_2161);
or U8588 (N_8588,N_1673,N_1869);
or U8589 (N_8589,N_3328,N_2461);
xnor U8590 (N_8590,N_3867,N_1483);
nand U8591 (N_8591,N_1416,N_2721);
nand U8592 (N_8592,N_5790,N_1029);
and U8593 (N_8593,N_2817,N_5836);
or U8594 (N_8594,N_1663,N_1316);
and U8595 (N_8595,N_379,N_5317);
xnor U8596 (N_8596,N_5468,N_2414);
and U8597 (N_8597,N_4112,N_725);
and U8598 (N_8598,N_5280,N_4949);
or U8599 (N_8599,N_171,N_2228);
nand U8600 (N_8600,N_3729,N_2968);
or U8601 (N_8601,N_1806,N_3352);
or U8602 (N_8602,N_3514,N_2939);
or U8603 (N_8603,N_521,N_2573);
nand U8604 (N_8604,N_1487,N_2775);
or U8605 (N_8605,N_4951,N_2695);
xnor U8606 (N_8606,N_5373,N_2479);
and U8607 (N_8607,N_624,N_3771);
or U8608 (N_8608,N_5195,N_710);
nand U8609 (N_8609,N_1937,N_2830);
nand U8610 (N_8610,N_110,N_1049);
nand U8611 (N_8611,N_1288,N_270);
and U8612 (N_8612,N_5088,N_111);
nand U8613 (N_8613,N_3652,N_5303);
nand U8614 (N_8614,N_3446,N_1706);
nand U8615 (N_8615,N_3732,N_2609);
nand U8616 (N_8616,N_3527,N_5506);
nor U8617 (N_8617,N_681,N_2700);
nor U8618 (N_8618,N_2857,N_4924);
and U8619 (N_8619,N_943,N_3037);
and U8620 (N_8620,N_2507,N_2910);
and U8621 (N_8621,N_1224,N_4826);
xnor U8622 (N_8622,N_5549,N_17);
nor U8623 (N_8623,N_916,N_913);
or U8624 (N_8624,N_4128,N_3561);
xnor U8625 (N_8625,N_3100,N_2176);
or U8626 (N_8626,N_518,N_105);
xnor U8627 (N_8627,N_1543,N_5900);
nor U8628 (N_8628,N_1077,N_992);
xor U8629 (N_8629,N_1414,N_1349);
and U8630 (N_8630,N_307,N_2766);
nor U8631 (N_8631,N_3954,N_4249);
nor U8632 (N_8632,N_90,N_5823);
or U8633 (N_8633,N_569,N_843);
or U8634 (N_8634,N_4163,N_3250);
nand U8635 (N_8635,N_5501,N_2899);
nor U8636 (N_8636,N_3599,N_5044);
xor U8637 (N_8637,N_5124,N_1824);
nand U8638 (N_8638,N_4871,N_949);
nor U8639 (N_8639,N_2579,N_4533);
and U8640 (N_8640,N_3562,N_1362);
xor U8641 (N_8641,N_5905,N_4628);
and U8642 (N_8642,N_4350,N_1120);
and U8643 (N_8643,N_5271,N_179);
nand U8644 (N_8644,N_5920,N_2963);
or U8645 (N_8645,N_5010,N_122);
and U8646 (N_8646,N_3982,N_3537);
and U8647 (N_8647,N_2407,N_3099);
nand U8648 (N_8648,N_5175,N_1772);
xnor U8649 (N_8649,N_1816,N_1094);
and U8650 (N_8650,N_1519,N_4649);
and U8651 (N_8651,N_3361,N_3410);
nand U8652 (N_8652,N_2728,N_858);
and U8653 (N_8653,N_2787,N_3104);
nor U8654 (N_8654,N_3650,N_1518);
nand U8655 (N_8655,N_4621,N_5564);
nor U8656 (N_8656,N_283,N_1827);
and U8657 (N_8657,N_5963,N_4340);
xnor U8658 (N_8658,N_2148,N_4906);
xnor U8659 (N_8659,N_4945,N_1462);
xor U8660 (N_8660,N_5257,N_2885);
nor U8661 (N_8661,N_5514,N_3753);
or U8662 (N_8662,N_5244,N_96);
nor U8663 (N_8663,N_1903,N_744);
and U8664 (N_8664,N_923,N_2364);
nor U8665 (N_8665,N_1605,N_1202);
or U8666 (N_8666,N_1747,N_233);
and U8667 (N_8667,N_1101,N_3664);
xnor U8668 (N_8668,N_5917,N_4594);
nor U8669 (N_8669,N_5151,N_52);
nor U8670 (N_8670,N_2915,N_5096);
or U8671 (N_8671,N_49,N_2353);
and U8672 (N_8672,N_536,N_5048);
nor U8673 (N_8673,N_4841,N_3362);
nand U8674 (N_8674,N_2370,N_5300);
and U8675 (N_8675,N_620,N_640);
xor U8676 (N_8676,N_2428,N_120);
or U8677 (N_8677,N_5541,N_1807);
and U8678 (N_8678,N_918,N_1363);
xor U8679 (N_8679,N_5417,N_4166);
nor U8680 (N_8680,N_4736,N_4870);
nand U8681 (N_8681,N_3453,N_3970);
xnor U8682 (N_8682,N_1936,N_3957);
or U8683 (N_8683,N_3425,N_206);
nand U8684 (N_8684,N_3863,N_3552);
xnor U8685 (N_8685,N_4575,N_238);
nor U8686 (N_8686,N_1212,N_1767);
xnor U8687 (N_8687,N_1365,N_1944);
and U8688 (N_8688,N_3499,N_3077);
nand U8689 (N_8689,N_3321,N_2332);
xor U8690 (N_8690,N_4056,N_1666);
and U8691 (N_8691,N_5974,N_1226);
or U8692 (N_8692,N_2566,N_5167);
nor U8693 (N_8693,N_4609,N_3166);
nand U8694 (N_8694,N_309,N_2469);
and U8695 (N_8695,N_4396,N_2239);
and U8696 (N_8696,N_5865,N_4988);
xor U8697 (N_8697,N_4681,N_1046);
nor U8698 (N_8698,N_5972,N_2977);
nand U8699 (N_8699,N_4407,N_5264);
and U8700 (N_8700,N_3828,N_1631);
and U8701 (N_8701,N_3063,N_1201);
and U8702 (N_8702,N_5168,N_3629);
xor U8703 (N_8703,N_1760,N_3894);
or U8704 (N_8704,N_3275,N_730);
and U8705 (N_8705,N_4200,N_5671);
nand U8706 (N_8706,N_5450,N_3065);
or U8707 (N_8707,N_130,N_1080);
nor U8708 (N_8708,N_2133,N_2747);
nor U8709 (N_8709,N_3512,N_3786);
xor U8710 (N_8710,N_4953,N_5102);
or U8711 (N_8711,N_2763,N_2513);
nor U8712 (N_8712,N_2545,N_2815);
nand U8713 (N_8713,N_778,N_5799);
or U8714 (N_8714,N_5001,N_2221);
xor U8715 (N_8715,N_2274,N_4579);
nand U8716 (N_8716,N_5767,N_4489);
and U8717 (N_8717,N_3878,N_2377);
or U8718 (N_8718,N_1024,N_5002);
or U8719 (N_8719,N_1550,N_5961);
and U8720 (N_8720,N_5155,N_1198);
or U8721 (N_8721,N_919,N_3751);
nor U8722 (N_8722,N_3339,N_1570);
or U8723 (N_8723,N_4938,N_5223);
xnor U8724 (N_8724,N_5989,N_3366);
nor U8725 (N_8725,N_3229,N_1549);
xnor U8726 (N_8726,N_4472,N_4282);
nor U8727 (N_8727,N_3194,N_2480);
xor U8728 (N_8728,N_4154,N_3195);
and U8729 (N_8729,N_4262,N_5914);
nor U8730 (N_8730,N_3256,N_3571);
nand U8731 (N_8731,N_4235,N_5253);
nor U8732 (N_8732,N_3432,N_1940);
nand U8733 (N_8733,N_5112,N_3919);
xor U8734 (N_8734,N_1819,N_3979);
nand U8735 (N_8735,N_5840,N_2788);
nand U8736 (N_8736,N_1636,N_2065);
xor U8737 (N_8737,N_29,N_1012);
and U8738 (N_8738,N_2784,N_2136);
or U8739 (N_8739,N_2378,N_2603);
xor U8740 (N_8740,N_2572,N_2181);
nor U8741 (N_8741,N_1138,N_1956);
and U8742 (N_8742,N_3582,N_3824);
nand U8743 (N_8743,N_3027,N_3706);
or U8744 (N_8744,N_4468,N_1133);
xnor U8745 (N_8745,N_3367,N_4121);
nand U8746 (N_8746,N_1471,N_5735);
xor U8747 (N_8747,N_2363,N_2851);
xor U8748 (N_8748,N_3164,N_1915);
xor U8749 (N_8749,N_668,N_1796);
and U8750 (N_8750,N_5689,N_118);
or U8751 (N_8751,N_2064,N_4195);
or U8752 (N_8752,N_2661,N_1883);
nor U8753 (N_8753,N_1058,N_1727);
or U8754 (N_8754,N_3429,N_3307);
nor U8755 (N_8755,N_2607,N_4748);
nor U8756 (N_8756,N_4759,N_5968);
and U8757 (N_8757,N_2535,N_4014);
xor U8758 (N_8758,N_3903,N_4895);
xnor U8759 (N_8759,N_1269,N_1498);
xor U8760 (N_8760,N_4622,N_812);
xor U8761 (N_8761,N_2361,N_3938);
and U8762 (N_8762,N_4165,N_3846);
or U8763 (N_8763,N_5224,N_4839);
and U8764 (N_8764,N_4547,N_2693);
xor U8765 (N_8765,N_1872,N_5348);
xnor U8766 (N_8766,N_4914,N_761);
nor U8767 (N_8767,N_1432,N_4129);
xnor U8768 (N_8768,N_2295,N_779);
xor U8769 (N_8769,N_3875,N_1409);
and U8770 (N_8770,N_298,N_2240);
nand U8771 (N_8771,N_4341,N_2108);
nand U8772 (N_8772,N_3981,N_3690);
nand U8773 (N_8773,N_3087,N_4932);
or U8774 (N_8774,N_1546,N_5746);
or U8775 (N_8775,N_2837,N_1163);
nand U8776 (N_8776,N_5294,N_4164);
and U8777 (N_8777,N_3627,N_183);
nor U8778 (N_8778,N_1602,N_3126);
or U8779 (N_8779,N_3379,N_2322);
or U8780 (N_8780,N_1417,N_2284);
nand U8781 (N_8781,N_980,N_1000);
or U8782 (N_8782,N_3483,N_4155);
nor U8783 (N_8783,N_3216,N_2863);
nand U8784 (N_8784,N_545,N_888);
nor U8785 (N_8785,N_182,N_3604);
xnor U8786 (N_8786,N_4419,N_1598);
nand U8787 (N_8787,N_1344,N_2962);
or U8788 (N_8788,N_731,N_3120);
xnor U8789 (N_8789,N_2063,N_818);
xor U8790 (N_8790,N_2335,N_12);
nor U8791 (N_8791,N_377,N_933);
or U8792 (N_8792,N_5895,N_5150);
xor U8793 (N_8793,N_2012,N_4272);
nand U8794 (N_8794,N_165,N_5952);
xor U8795 (N_8795,N_782,N_1401);
or U8796 (N_8796,N_5829,N_412);
nor U8797 (N_8797,N_4751,N_3018);
nor U8798 (N_8798,N_1135,N_2447);
and U8799 (N_8799,N_5529,N_1947);
or U8800 (N_8800,N_3698,N_5301);
nand U8801 (N_8801,N_489,N_816);
nor U8802 (N_8802,N_1396,N_3342);
or U8803 (N_8803,N_3718,N_3931);
and U8804 (N_8804,N_141,N_4620);
or U8805 (N_8805,N_275,N_133);
and U8806 (N_8806,N_3612,N_1911);
xnor U8807 (N_8807,N_3017,N_3170);
and U8808 (N_8808,N_4540,N_4361);
or U8809 (N_8809,N_1108,N_3793);
xor U8810 (N_8810,N_2430,N_824);
nor U8811 (N_8811,N_4544,N_4209);
nor U8812 (N_8812,N_975,N_967);
and U8813 (N_8813,N_322,N_1931);
xnor U8814 (N_8814,N_2652,N_3125);
or U8815 (N_8815,N_4792,N_679);
xnor U8816 (N_8816,N_5994,N_3057);
or U8817 (N_8817,N_216,N_659);
nand U8818 (N_8818,N_3758,N_2967);
xnor U8819 (N_8819,N_762,N_4703);
and U8820 (N_8820,N_5460,N_152);
xor U8821 (N_8821,N_2814,N_22);
xnor U8822 (N_8822,N_5860,N_4302);
and U8823 (N_8823,N_1689,N_3952);
nand U8824 (N_8824,N_655,N_4767);
xnor U8825 (N_8825,N_808,N_349);
nand U8826 (N_8826,N_2645,N_3445);
or U8827 (N_8827,N_3985,N_4401);
xor U8828 (N_8828,N_1144,N_440);
xor U8829 (N_8829,N_1452,N_4285);
xnor U8830 (N_8830,N_5576,N_243);
or U8831 (N_8831,N_749,N_5066);
xnor U8832 (N_8832,N_124,N_150);
and U8833 (N_8833,N_2315,N_2100);
nor U8834 (N_8834,N_2425,N_4696);
xor U8835 (N_8835,N_2712,N_3654);
nand U8836 (N_8836,N_5666,N_677);
and U8837 (N_8837,N_3531,N_4527);
nor U8838 (N_8838,N_783,N_1464);
xor U8839 (N_8839,N_3029,N_4092);
nor U8840 (N_8840,N_2909,N_3890);
xnor U8841 (N_8841,N_3836,N_2376);
or U8842 (N_8842,N_3070,N_2279);
nand U8843 (N_8843,N_199,N_1051);
nand U8844 (N_8844,N_898,N_4785);
or U8845 (N_8845,N_3937,N_434);
or U8846 (N_8846,N_3677,N_4623);
and U8847 (N_8847,N_551,N_927);
nand U8848 (N_8848,N_5127,N_1480);
or U8849 (N_8849,N_481,N_1342);
or U8850 (N_8850,N_4885,N_2892);
and U8851 (N_8851,N_2667,N_5256);
and U8852 (N_8852,N_4003,N_4566);
xor U8853 (N_8853,N_2706,N_333);
nand U8854 (N_8854,N_139,N_4587);
nor U8855 (N_8855,N_4080,N_1919);
nand U8856 (N_8856,N_2650,N_32);
xnor U8857 (N_8857,N_3620,N_4274);
nand U8858 (N_8858,N_4131,N_2272);
nand U8859 (N_8859,N_4844,N_3085);
xnor U8860 (N_8860,N_3625,N_2022);
nor U8861 (N_8861,N_3289,N_5932);
nand U8862 (N_8862,N_2733,N_3396);
or U8863 (N_8863,N_1053,N_4342);
or U8864 (N_8864,N_1621,N_1010);
xnor U8865 (N_8865,N_4695,N_5706);
and U8866 (N_8866,N_485,N_5652);
xor U8867 (N_8867,N_5291,N_4507);
nor U8868 (N_8868,N_2354,N_1777);
or U8869 (N_8869,N_4178,N_2901);
xor U8870 (N_8870,N_4910,N_4746);
and U8871 (N_8871,N_5644,N_1433);
nor U8872 (N_8872,N_3430,N_4414);
or U8873 (N_8873,N_1507,N_192);
or U8874 (N_8874,N_4442,N_1532);
and U8875 (N_8875,N_2945,N_3078);
nand U8876 (N_8876,N_3659,N_3857);
nor U8877 (N_8877,N_4473,N_1882);
xnor U8878 (N_8878,N_1465,N_1147);
nand U8879 (N_8879,N_2141,N_5610);
or U8880 (N_8880,N_1104,N_4392);
and U8881 (N_8881,N_4915,N_5718);
nand U8882 (N_8882,N_2128,N_5246);
nand U8883 (N_8883,N_4223,N_4211);
xnor U8884 (N_8884,N_763,N_4905);
nand U8885 (N_8885,N_2431,N_370);
nor U8886 (N_8886,N_3618,N_1759);
or U8887 (N_8887,N_5340,N_557);
xor U8888 (N_8888,N_3683,N_5200);
nor U8889 (N_8889,N_3157,N_1394);
and U8890 (N_8890,N_1800,N_2633);
or U8891 (N_8891,N_2663,N_3128);
and U8892 (N_8892,N_5331,N_2304);
and U8893 (N_8893,N_5447,N_5496);
xnor U8894 (N_8894,N_846,N_5909);
nor U8895 (N_8895,N_3090,N_2257);
xor U8896 (N_8896,N_5259,N_2250);
or U8897 (N_8897,N_5179,N_4023);
or U8898 (N_8898,N_1980,N_2657);
nand U8899 (N_8899,N_4655,N_1674);
or U8900 (N_8900,N_2351,N_459);
xnor U8901 (N_8901,N_59,N_4667);
nand U8902 (N_8902,N_2791,N_5824);
xnor U8903 (N_8903,N_1916,N_1255);
nand U8904 (N_8904,N_112,N_4897);
xor U8905 (N_8905,N_1497,N_4925);
and U8906 (N_8906,N_3515,N_4045);
xnor U8907 (N_8907,N_1742,N_3990);
or U8908 (N_8908,N_700,N_3395);
and U8909 (N_8909,N_4825,N_2449);
nand U8910 (N_8910,N_3169,N_4995);
and U8911 (N_8911,N_3026,N_2656);
xnor U8912 (N_8912,N_2226,N_2303);
and U8913 (N_8913,N_1864,N_4770);
xnor U8914 (N_8914,N_3338,N_1562);
nor U8915 (N_8915,N_1766,N_676);
nor U8916 (N_8916,N_4089,N_3012);
xnor U8917 (N_8917,N_5924,N_3774);
xor U8918 (N_8918,N_2536,N_2568);
and U8919 (N_8919,N_2585,N_772);
and U8920 (N_8920,N_3079,N_5805);
xor U8921 (N_8921,N_3948,N_1853);
nor U8922 (N_8922,N_5261,N_468);
xor U8923 (N_8923,N_3416,N_2024);
nor U8924 (N_8924,N_2085,N_1332);
or U8925 (N_8925,N_3854,N_4966);
nor U8926 (N_8926,N_2989,N_187);
nand U8927 (N_8927,N_3513,N_893);
nor U8928 (N_8928,N_5540,N_3163);
or U8929 (N_8929,N_1267,N_651);
xor U8930 (N_8930,N_697,N_4926);
nand U8931 (N_8931,N_4994,N_2646);
xor U8932 (N_8932,N_5318,N_2498);
nor U8933 (N_8933,N_5094,N_3738);
xor U8934 (N_8934,N_1993,N_3660);
nand U8935 (N_8935,N_5593,N_94);
nor U8936 (N_8936,N_1079,N_2956);
or U8937 (N_8937,N_4835,N_3298);
xnor U8938 (N_8938,N_2624,N_4738);
xnor U8939 (N_8939,N_317,N_2625);
nand U8940 (N_8940,N_728,N_5219);
and U8941 (N_8941,N_2131,N_5427);
xnor U8942 (N_8942,N_4889,N_4229);
nor U8943 (N_8943,N_1575,N_1525);
or U8944 (N_8944,N_131,N_3964);
and U8945 (N_8945,N_4644,N_1161);
xnor U8946 (N_8946,N_5817,N_5391);
and U8947 (N_8947,N_4326,N_4198);
nand U8948 (N_8948,N_4337,N_5844);
nand U8949 (N_8949,N_5186,N_3568);
and U8950 (N_8950,N_4611,N_1123);
or U8951 (N_8951,N_1412,N_4673);
or U8952 (N_8952,N_2175,N_3477);
nand U8953 (N_8953,N_650,N_1637);
nor U8954 (N_8954,N_3737,N_1725);
xor U8955 (N_8955,N_5826,N_4167);
xor U8956 (N_8956,N_2016,N_4241);
xnor U8957 (N_8957,N_917,N_3976);
and U8958 (N_8958,N_4819,N_5797);
nor U8959 (N_8959,N_1247,N_5057);
xor U8960 (N_8960,N_1720,N_5335);
or U8961 (N_8961,N_1652,N_3581);
nor U8962 (N_8962,N_371,N_287);
xor U8963 (N_8963,N_4831,N_455);
xnor U8964 (N_8964,N_1486,N_2839);
nor U8965 (N_8965,N_562,N_1905);
xnor U8966 (N_8966,N_5554,N_4954);
xnor U8967 (N_8967,N_4976,N_2974);
nor U8968 (N_8968,N_176,N_5284);
nand U8969 (N_8969,N_1327,N_156);
and U8970 (N_8970,N_3602,N_5522);
nor U8971 (N_8971,N_2636,N_1005);
nand U8972 (N_8972,N_5672,N_2441);
xor U8973 (N_8973,N_2023,N_969);
nor U8974 (N_8974,N_2078,N_5060);
and U8975 (N_8975,N_941,N_99);
xor U8976 (N_8976,N_4391,N_4292);
or U8977 (N_8977,N_5177,N_3491);
and U8978 (N_8978,N_1972,N_3389);
xor U8979 (N_8979,N_4589,N_284);
xnor U8980 (N_8980,N_1023,N_1723);
nor U8981 (N_8981,N_1137,N_612);
and U8982 (N_8982,N_4762,N_1062);
nand U8983 (N_8983,N_4847,N_1758);
and U8984 (N_8984,N_2792,N_2444);
nand U8985 (N_8985,N_5372,N_1658);
and U8986 (N_8986,N_1188,N_4603);
xnor U8987 (N_8987,N_297,N_2729);
or U8988 (N_8988,N_5841,N_4005);
or U8989 (N_8989,N_5842,N_1265);
xor U8990 (N_8990,N_4070,N_3896);
or U8991 (N_8991,N_3199,N_1186);
and U8992 (N_8992,N_3015,N_947);
or U8993 (N_8993,N_4078,N_3316);
and U8994 (N_8994,N_185,N_3011);
xnor U8995 (N_8995,N_1987,N_2138);
or U8996 (N_8996,N_1252,N_4464);
and U8997 (N_8997,N_4697,N_4786);
nand U8998 (N_8998,N_5802,N_1022);
or U8999 (N_8999,N_4214,N_1302);
xor U9000 (N_9000,N_3881,N_2176);
or U9001 (N_9001,N_3091,N_5845);
nand U9002 (N_9002,N_3354,N_961);
nor U9003 (N_9003,N_1905,N_842);
nand U9004 (N_9004,N_2472,N_2535);
and U9005 (N_9005,N_2735,N_3715);
nor U9006 (N_9006,N_4952,N_1945);
or U9007 (N_9007,N_3239,N_1336);
nand U9008 (N_9008,N_2945,N_3395);
or U9009 (N_9009,N_2576,N_5611);
nand U9010 (N_9010,N_5585,N_3544);
or U9011 (N_9011,N_5606,N_3217);
or U9012 (N_9012,N_3662,N_1872);
and U9013 (N_9013,N_4792,N_3413);
nand U9014 (N_9014,N_2371,N_1848);
and U9015 (N_9015,N_1774,N_2058);
and U9016 (N_9016,N_1909,N_5022);
xor U9017 (N_9017,N_5711,N_2004);
and U9018 (N_9018,N_5685,N_1268);
xor U9019 (N_9019,N_2363,N_3264);
nand U9020 (N_9020,N_4930,N_2608);
and U9021 (N_9021,N_22,N_1952);
nand U9022 (N_9022,N_1520,N_5253);
or U9023 (N_9023,N_1448,N_4754);
nor U9024 (N_9024,N_5644,N_467);
nand U9025 (N_9025,N_4222,N_3979);
or U9026 (N_9026,N_1493,N_4789);
and U9027 (N_9027,N_5196,N_2450);
nand U9028 (N_9028,N_3103,N_4233);
xnor U9029 (N_9029,N_4682,N_3591);
and U9030 (N_9030,N_4246,N_3375);
or U9031 (N_9031,N_4158,N_1272);
or U9032 (N_9032,N_3083,N_1500);
nor U9033 (N_9033,N_1670,N_4631);
or U9034 (N_9034,N_3094,N_3609);
or U9035 (N_9035,N_475,N_773);
xor U9036 (N_9036,N_4224,N_1567);
or U9037 (N_9037,N_4048,N_648);
nor U9038 (N_9038,N_3822,N_5273);
xor U9039 (N_9039,N_1589,N_4806);
or U9040 (N_9040,N_5921,N_5307);
nand U9041 (N_9041,N_567,N_4622);
xnor U9042 (N_9042,N_5319,N_3935);
xor U9043 (N_9043,N_1387,N_212);
nand U9044 (N_9044,N_1536,N_3496);
nand U9045 (N_9045,N_4568,N_1324);
nor U9046 (N_9046,N_5409,N_4778);
nand U9047 (N_9047,N_3337,N_4923);
and U9048 (N_9048,N_3593,N_4999);
xor U9049 (N_9049,N_2789,N_4653);
xor U9050 (N_9050,N_910,N_5700);
or U9051 (N_9051,N_5516,N_644);
and U9052 (N_9052,N_1028,N_389);
xnor U9053 (N_9053,N_3194,N_882);
nor U9054 (N_9054,N_2665,N_4730);
nand U9055 (N_9055,N_2511,N_1727);
or U9056 (N_9056,N_742,N_856);
nor U9057 (N_9057,N_4978,N_4009);
xor U9058 (N_9058,N_2877,N_4578);
and U9059 (N_9059,N_3120,N_2152);
or U9060 (N_9060,N_2103,N_4101);
and U9061 (N_9061,N_5980,N_2499);
and U9062 (N_9062,N_1529,N_2568);
nand U9063 (N_9063,N_1691,N_4218);
nor U9064 (N_9064,N_608,N_1426);
or U9065 (N_9065,N_1628,N_3423);
xnor U9066 (N_9066,N_2524,N_2251);
or U9067 (N_9067,N_5951,N_3577);
or U9068 (N_9068,N_479,N_2421);
xor U9069 (N_9069,N_5804,N_2619);
and U9070 (N_9070,N_2188,N_602);
nand U9071 (N_9071,N_3657,N_5833);
or U9072 (N_9072,N_5109,N_4952);
xnor U9073 (N_9073,N_4541,N_5274);
nand U9074 (N_9074,N_1153,N_1515);
or U9075 (N_9075,N_730,N_628);
xor U9076 (N_9076,N_34,N_5574);
nor U9077 (N_9077,N_2469,N_332);
xor U9078 (N_9078,N_3771,N_716);
or U9079 (N_9079,N_824,N_874);
and U9080 (N_9080,N_2819,N_4851);
or U9081 (N_9081,N_422,N_2364);
nand U9082 (N_9082,N_3932,N_15);
and U9083 (N_9083,N_5741,N_3692);
nor U9084 (N_9084,N_2843,N_3176);
nand U9085 (N_9085,N_3138,N_1687);
or U9086 (N_9086,N_2847,N_1212);
xor U9087 (N_9087,N_1429,N_1330);
nand U9088 (N_9088,N_1183,N_4326);
nor U9089 (N_9089,N_5582,N_1995);
or U9090 (N_9090,N_4627,N_4784);
and U9091 (N_9091,N_3087,N_865);
and U9092 (N_9092,N_4808,N_4054);
xnor U9093 (N_9093,N_1896,N_1927);
and U9094 (N_9094,N_2209,N_3120);
nor U9095 (N_9095,N_100,N_2820);
and U9096 (N_9096,N_2772,N_2219);
or U9097 (N_9097,N_3749,N_4712);
nand U9098 (N_9098,N_4070,N_1855);
and U9099 (N_9099,N_1934,N_5585);
xor U9100 (N_9100,N_3588,N_632);
or U9101 (N_9101,N_5349,N_2072);
nand U9102 (N_9102,N_5320,N_4047);
or U9103 (N_9103,N_1358,N_5124);
or U9104 (N_9104,N_4861,N_3139);
xnor U9105 (N_9105,N_4013,N_1652);
nand U9106 (N_9106,N_2646,N_1018);
xnor U9107 (N_9107,N_4081,N_5420);
and U9108 (N_9108,N_4764,N_5494);
xor U9109 (N_9109,N_1685,N_5605);
nand U9110 (N_9110,N_418,N_979);
nand U9111 (N_9111,N_671,N_1045);
nor U9112 (N_9112,N_4028,N_3754);
nand U9113 (N_9113,N_619,N_5582);
or U9114 (N_9114,N_1335,N_3598);
and U9115 (N_9115,N_2771,N_3528);
nor U9116 (N_9116,N_268,N_4757);
or U9117 (N_9117,N_785,N_5975);
nor U9118 (N_9118,N_5098,N_5328);
nand U9119 (N_9119,N_3862,N_1206);
or U9120 (N_9120,N_916,N_5539);
xor U9121 (N_9121,N_285,N_1577);
and U9122 (N_9122,N_3163,N_3976);
xnor U9123 (N_9123,N_4785,N_2794);
and U9124 (N_9124,N_5815,N_2848);
nor U9125 (N_9125,N_1406,N_5162);
nor U9126 (N_9126,N_3547,N_1723);
nor U9127 (N_9127,N_3415,N_52);
xor U9128 (N_9128,N_4750,N_4646);
or U9129 (N_9129,N_2215,N_5516);
or U9130 (N_9130,N_3992,N_4910);
or U9131 (N_9131,N_287,N_2798);
nand U9132 (N_9132,N_5585,N_5865);
xnor U9133 (N_9133,N_1769,N_985);
nand U9134 (N_9134,N_1458,N_2126);
and U9135 (N_9135,N_907,N_238);
xnor U9136 (N_9136,N_5446,N_4021);
or U9137 (N_9137,N_3487,N_1498);
nor U9138 (N_9138,N_2182,N_1129);
nand U9139 (N_9139,N_2893,N_1019);
nor U9140 (N_9140,N_3401,N_5561);
nand U9141 (N_9141,N_539,N_2670);
nor U9142 (N_9142,N_3189,N_2758);
nand U9143 (N_9143,N_968,N_172);
xor U9144 (N_9144,N_2540,N_994);
xor U9145 (N_9145,N_2018,N_5017);
nor U9146 (N_9146,N_1012,N_5299);
nand U9147 (N_9147,N_2310,N_1864);
and U9148 (N_9148,N_1446,N_798);
and U9149 (N_9149,N_65,N_95);
or U9150 (N_9150,N_4999,N_4398);
and U9151 (N_9151,N_1138,N_3817);
or U9152 (N_9152,N_5793,N_102);
xor U9153 (N_9153,N_3917,N_3826);
or U9154 (N_9154,N_856,N_1322);
and U9155 (N_9155,N_1259,N_2431);
nor U9156 (N_9156,N_3966,N_2959);
nor U9157 (N_9157,N_2317,N_2722);
and U9158 (N_9158,N_2072,N_3524);
and U9159 (N_9159,N_1510,N_4442);
nor U9160 (N_9160,N_4465,N_2544);
nor U9161 (N_9161,N_4450,N_4325);
xnor U9162 (N_9162,N_4783,N_5267);
nand U9163 (N_9163,N_129,N_3616);
nand U9164 (N_9164,N_3836,N_4840);
and U9165 (N_9165,N_5411,N_3380);
and U9166 (N_9166,N_4388,N_5204);
nand U9167 (N_9167,N_2434,N_3895);
or U9168 (N_9168,N_3191,N_4348);
or U9169 (N_9169,N_2983,N_1761);
or U9170 (N_9170,N_4454,N_646);
nor U9171 (N_9171,N_3018,N_4334);
and U9172 (N_9172,N_4656,N_2338);
nand U9173 (N_9173,N_800,N_504);
and U9174 (N_9174,N_4759,N_5481);
xor U9175 (N_9175,N_4259,N_1251);
nand U9176 (N_9176,N_3111,N_5329);
or U9177 (N_9177,N_5846,N_3228);
nand U9178 (N_9178,N_5589,N_2774);
nand U9179 (N_9179,N_4728,N_4169);
nor U9180 (N_9180,N_5071,N_5749);
nand U9181 (N_9181,N_85,N_2217);
nor U9182 (N_9182,N_2825,N_3705);
nand U9183 (N_9183,N_2194,N_3385);
and U9184 (N_9184,N_2639,N_481);
nor U9185 (N_9185,N_3717,N_4404);
nand U9186 (N_9186,N_2417,N_2272);
nand U9187 (N_9187,N_1249,N_1215);
or U9188 (N_9188,N_1356,N_3036);
nand U9189 (N_9189,N_347,N_1797);
nand U9190 (N_9190,N_5054,N_42);
or U9191 (N_9191,N_4466,N_1585);
or U9192 (N_9192,N_4554,N_2184);
nand U9193 (N_9193,N_2239,N_408);
or U9194 (N_9194,N_4524,N_1092);
nor U9195 (N_9195,N_2250,N_604);
or U9196 (N_9196,N_1128,N_1751);
nor U9197 (N_9197,N_5941,N_5769);
and U9198 (N_9198,N_5357,N_2219);
nand U9199 (N_9199,N_2512,N_5753);
and U9200 (N_9200,N_2273,N_3186);
nand U9201 (N_9201,N_1458,N_3560);
xnor U9202 (N_9202,N_818,N_3809);
or U9203 (N_9203,N_3084,N_1590);
and U9204 (N_9204,N_2093,N_4617);
or U9205 (N_9205,N_3911,N_5428);
xor U9206 (N_9206,N_1639,N_4717);
nand U9207 (N_9207,N_5794,N_4769);
or U9208 (N_9208,N_3932,N_4764);
or U9209 (N_9209,N_2382,N_668);
xnor U9210 (N_9210,N_2909,N_2261);
nor U9211 (N_9211,N_5473,N_540);
and U9212 (N_9212,N_1465,N_4169);
xnor U9213 (N_9213,N_1849,N_2417);
nor U9214 (N_9214,N_5366,N_3833);
nor U9215 (N_9215,N_3089,N_2561);
nor U9216 (N_9216,N_5449,N_3473);
and U9217 (N_9217,N_2076,N_3000);
or U9218 (N_9218,N_2623,N_3055);
or U9219 (N_9219,N_368,N_762);
and U9220 (N_9220,N_5162,N_1657);
nand U9221 (N_9221,N_1165,N_1404);
nand U9222 (N_9222,N_530,N_522);
nand U9223 (N_9223,N_4101,N_2098);
and U9224 (N_9224,N_1,N_90);
nand U9225 (N_9225,N_673,N_1746);
and U9226 (N_9226,N_4439,N_2381);
nand U9227 (N_9227,N_5962,N_5204);
nand U9228 (N_9228,N_5313,N_2971);
nand U9229 (N_9229,N_1563,N_5550);
or U9230 (N_9230,N_4861,N_92);
nor U9231 (N_9231,N_5327,N_999);
and U9232 (N_9232,N_27,N_1795);
or U9233 (N_9233,N_1793,N_554);
or U9234 (N_9234,N_4909,N_3010);
or U9235 (N_9235,N_4846,N_5821);
or U9236 (N_9236,N_4229,N_2992);
nand U9237 (N_9237,N_4292,N_5140);
and U9238 (N_9238,N_5784,N_2663);
or U9239 (N_9239,N_792,N_2824);
and U9240 (N_9240,N_3436,N_5343);
and U9241 (N_9241,N_3764,N_3141);
or U9242 (N_9242,N_1058,N_5963);
nand U9243 (N_9243,N_2268,N_2883);
and U9244 (N_9244,N_124,N_290);
nor U9245 (N_9245,N_3671,N_578);
or U9246 (N_9246,N_2862,N_4724);
nor U9247 (N_9247,N_4229,N_3265);
nor U9248 (N_9248,N_5333,N_1501);
or U9249 (N_9249,N_1053,N_2257);
nand U9250 (N_9250,N_5504,N_2418);
nor U9251 (N_9251,N_4135,N_4051);
nand U9252 (N_9252,N_3325,N_5231);
xnor U9253 (N_9253,N_203,N_287);
nand U9254 (N_9254,N_2295,N_1314);
and U9255 (N_9255,N_4408,N_1811);
xor U9256 (N_9256,N_5025,N_2774);
nand U9257 (N_9257,N_1930,N_1164);
xnor U9258 (N_9258,N_2383,N_1890);
nor U9259 (N_9259,N_5771,N_2920);
and U9260 (N_9260,N_1355,N_841);
xnor U9261 (N_9261,N_4487,N_3974);
and U9262 (N_9262,N_1821,N_2266);
xor U9263 (N_9263,N_5682,N_1408);
or U9264 (N_9264,N_5764,N_4998);
nor U9265 (N_9265,N_3394,N_5867);
and U9266 (N_9266,N_3983,N_1473);
xnor U9267 (N_9267,N_2444,N_5638);
and U9268 (N_9268,N_2721,N_311);
and U9269 (N_9269,N_5411,N_976);
xor U9270 (N_9270,N_4751,N_3095);
and U9271 (N_9271,N_1041,N_3095);
nand U9272 (N_9272,N_4179,N_4635);
nand U9273 (N_9273,N_5246,N_4509);
nor U9274 (N_9274,N_3059,N_2380);
and U9275 (N_9275,N_756,N_802);
and U9276 (N_9276,N_906,N_5773);
nand U9277 (N_9277,N_5760,N_2890);
and U9278 (N_9278,N_4887,N_3718);
nor U9279 (N_9279,N_915,N_268);
and U9280 (N_9280,N_4159,N_4473);
or U9281 (N_9281,N_1813,N_2606);
or U9282 (N_9282,N_3935,N_5679);
nor U9283 (N_9283,N_1842,N_5192);
nor U9284 (N_9284,N_1536,N_1978);
and U9285 (N_9285,N_2737,N_1291);
or U9286 (N_9286,N_4314,N_5186);
or U9287 (N_9287,N_130,N_1972);
xor U9288 (N_9288,N_1482,N_4262);
nor U9289 (N_9289,N_3949,N_1086);
xnor U9290 (N_9290,N_773,N_4391);
nand U9291 (N_9291,N_4689,N_3171);
nand U9292 (N_9292,N_2796,N_2647);
nand U9293 (N_9293,N_1493,N_2233);
xnor U9294 (N_9294,N_1021,N_2292);
and U9295 (N_9295,N_5571,N_1266);
xnor U9296 (N_9296,N_3251,N_3386);
nand U9297 (N_9297,N_3158,N_292);
and U9298 (N_9298,N_5715,N_3278);
and U9299 (N_9299,N_234,N_2590);
xor U9300 (N_9300,N_2666,N_3325);
or U9301 (N_9301,N_570,N_2996);
nor U9302 (N_9302,N_3378,N_2714);
nor U9303 (N_9303,N_3731,N_5813);
and U9304 (N_9304,N_3175,N_443);
nor U9305 (N_9305,N_4017,N_4759);
nand U9306 (N_9306,N_3519,N_777);
or U9307 (N_9307,N_4737,N_1115);
nand U9308 (N_9308,N_3484,N_4287);
xnor U9309 (N_9309,N_1390,N_4494);
or U9310 (N_9310,N_2537,N_1732);
or U9311 (N_9311,N_4704,N_789);
or U9312 (N_9312,N_3083,N_351);
and U9313 (N_9313,N_5254,N_5579);
xor U9314 (N_9314,N_4529,N_626);
nand U9315 (N_9315,N_4886,N_292);
nand U9316 (N_9316,N_1138,N_1879);
nor U9317 (N_9317,N_5472,N_1145);
and U9318 (N_9318,N_3827,N_5919);
xor U9319 (N_9319,N_835,N_288);
or U9320 (N_9320,N_3878,N_1131);
nand U9321 (N_9321,N_3320,N_334);
nand U9322 (N_9322,N_5119,N_78);
and U9323 (N_9323,N_1619,N_790);
and U9324 (N_9324,N_2715,N_3203);
and U9325 (N_9325,N_5249,N_3263);
nor U9326 (N_9326,N_1620,N_2017);
nand U9327 (N_9327,N_3862,N_2481);
nor U9328 (N_9328,N_1887,N_3943);
or U9329 (N_9329,N_5703,N_2699);
and U9330 (N_9330,N_2970,N_5599);
or U9331 (N_9331,N_384,N_3621);
and U9332 (N_9332,N_5625,N_2565);
nand U9333 (N_9333,N_4266,N_1430);
xnor U9334 (N_9334,N_914,N_1461);
or U9335 (N_9335,N_2163,N_457);
nand U9336 (N_9336,N_733,N_4436);
nand U9337 (N_9337,N_1698,N_2012);
and U9338 (N_9338,N_2349,N_4034);
and U9339 (N_9339,N_3469,N_3412);
or U9340 (N_9340,N_5813,N_1750);
xor U9341 (N_9341,N_4252,N_2442);
or U9342 (N_9342,N_2682,N_2141);
or U9343 (N_9343,N_3857,N_2491);
nand U9344 (N_9344,N_2816,N_3492);
and U9345 (N_9345,N_974,N_1540);
or U9346 (N_9346,N_4216,N_3013);
nand U9347 (N_9347,N_793,N_2279);
and U9348 (N_9348,N_591,N_4836);
xor U9349 (N_9349,N_748,N_5420);
nand U9350 (N_9350,N_957,N_2878);
xor U9351 (N_9351,N_4614,N_888);
xor U9352 (N_9352,N_2444,N_103);
nor U9353 (N_9353,N_2981,N_3373);
nor U9354 (N_9354,N_5601,N_2922);
nor U9355 (N_9355,N_4269,N_3747);
nand U9356 (N_9356,N_519,N_5678);
or U9357 (N_9357,N_1597,N_1108);
xnor U9358 (N_9358,N_4728,N_3022);
nor U9359 (N_9359,N_4878,N_4138);
xnor U9360 (N_9360,N_2406,N_3378);
and U9361 (N_9361,N_4810,N_4319);
or U9362 (N_9362,N_1752,N_2767);
nand U9363 (N_9363,N_4551,N_1883);
xor U9364 (N_9364,N_5327,N_1991);
nor U9365 (N_9365,N_4253,N_1865);
and U9366 (N_9366,N_1437,N_5134);
nand U9367 (N_9367,N_1489,N_1087);
nand U9368 (N_9368,N_5767,N_756);
xnor U9369 (N_9369,N_749,N_1564);
and U9370 (N_9370,N_1631,N_1985);
nand U9371 (N_9371,N_5634,N_692);
nand U9372 (N_9372,N_2883,N_86);
or U9373 (N_9373,N_4265,N_4515);
nor U9374 (N_9374,N_3392,N_2338);
nor U9375 (N_9375,N_5831,N_1612);
xor U9376 (N_9376,N_3801,N_137);
nand U9377 (N_9377,N_4216,N_4199);
nor U9378 (N_9378,N_5100,N_2793);
nor U9379 (N_9379,N_3215,N_3708);
and U9380 (N_9380,N_2091,N_2740);
nor U9381 (N_9381,N_5111,N_752);
and U9382 (N_9382,N_4763,N_5637);
nand U9383 (N_9383,N_3556,N_654);
nand U9384 (N_9384,N_1245,N_881);
and U9385 (N_9385,N_5460,N_61);
nand U9386 (N_9386,N_3182,N_3670);
or U9387 (N_9387,N_2826,N_3262);
nor U9388 (N_9388,N_5978,N_5913);
xnor U9389 (N_9389,N_4669,N_2701);
or U9390 (N_9390,N_5342,N_4596);
xor U9391 (N_9391,N_4142,N_1145);
or U9392 (N_9392,N_5676,N_3969);
and U9393 (N_9393,N_5263,N_2847);
or U9394 (N_9394,N_1081,N_5034);
xnor U9395 (N_9395,N_3370,N_2857);
xor U9396 (N_9396,N_5502,N_1110);
nand U9397 (N_9397,N_3656,N_3119);
xor U9398 (N_9398,N_5880,N_4793);
or U9399 (N_9399,N_3431,N_1920);
xnor U9400 (N_9400,N_5370,N_248);
nor U9401 (N_9401,N_4358,N_1819);
and U9402 (N_9402,N_3016,N_4321);
nor U9403 (N_9403,N_140,N_2932);
xnor U9404 (N_9404,N_5840,N_120);
xnor U9405 (N_9405,N_2222,N_4087);
or U9406 (N_9406,N_3206,N_667);
or U9407 (N_9407,N_3687,N_571);
nor U9408 (N_9408,N_4048,N_2382);
and U9409 (N_9409,N_3253,N_4395);
xnor U9410 (N_9410,N_4113,N_2887);
nand U9411 (N_9411,N_1067,N_1970);
or U9412 (N_9412,N_3011,N_4831);
or U9413 (N_9413,N_29,N_2207);
xnor U9414 (N_9414,N_1633,N_3964);
nor U9415 (N_9415,N_4473,N_103);
or U9416 (N_9416,N_4768,N_4621);
nand U9417 (N_9417,N_2059,N_5384);
and U9418 (N_9418,N_3086,N_427);
nand U9419 (N_9419,N_4085,N_3099);
and U9420 (N_9420,N_2937,N_1514);
nor U9421 (N_9421,N_4368,N_989);
nand U9422 (N_9422,N_1075,N_3867);
xor U9423 (N_9423,N_3643,N_117);
nor U9424 (N_9424,N_1890,N_307);
or U9425 (N_9425,N_1377,N_119);
xnor U9426 (N_9426,N_5040,N_4189);
xor U9427 (N_9427,N_4727,N_1461);
nand U9428 (N_9428,N_2223,N_2763);
and U9429 (N_9429,N_2490,N_2065);
nor U9430 (N_9430,N_3596,N_1763);
nor U9431 (N_9431,N_2662,N_404);
nand U9432 (N_9432,N_5771,N_344);
xor U9433 (N_9433,N_657,N_2836);
xor U9434 (N_9434,N_1220,N_1671);
nor U9435 (N_9435,N_1092,N_5057);
and U9436 (N_9436,N_5391,N_3501);
nand U9437 (N_9437,N_4026,N_4663);
nor U9438 (N_9438,N_4127,N_5643);
or U9439 (N_9439,N_3312,N_2595);
nand U9440 (N_9440,N_1168,N_2042);
xor U9441 (N_9441,N_1842,N_3157);
xnor U9442 (N_9442,N_1996,N_2186);
nand U9443 (N_9443,N_2495,N_5157);
nand U9444 (N_9444,N_1161,N_5223);
nand U9445 (N_9445,N_3396,N_4507);
nand U9446 (N_9446,N_1057,N_1189);
xnor U9447 (N_9447,N_3857,N_952);
and U9448 (N_9448,N_1497,N_5877);
nor U9449 (N_9449,N_1297,N_625);
xor U9450 (N_9450,N_2541,N_4672);
xor U9451 (N_9451,N_2411,N_862);
nor U9452 (N_9452,N_4686,N_91);
nor U9453 (N_9453,N_959,N_383);
and U9454 (N_9454,N_5640,N_1171);
xnor U9455 (N_9455,N_1998,N_3974);
xnor U9456 (N_9456,N_4651,N_2145);
nand U9457 (N_9457,N_5244,N_693);
nor U9458 (N_9458,N_5410,N_4985);
and U9459 (N_9459,N_4897,N_258);
xor U9460 (N_9460,N_498,N_4712);
nand U9461 (N_9461,N_4931,N_5373);
and U9462 (N_9462,N_3223,N_1975);
or U9463 (N_9463,N_993,N_937);
nor U9464 (N_9464,N_5710,N_3500);
nand U9465 (N_9465,N_796,N_56);
or U9466 (N_9466,N_537,N_4711);
or U9467 (N_9467,N_4123,N_3303);
and U9468 (N_9468,N_278,N_4620);
nand U9469 (N_9469,N_4806,N_2527);
and U9470 (N_9470,N_1038,N_3900);
and U9471 (N_9471,N_5342,N_581);
or U9472 (N_9472,N_2562,N_3261);
xnor U9473 (N_9473,N_2711,N_289);
xor U9474 (N_9474,N_736,N_4109);
nand U9475 (N_9475,N_3040,N_2283);
and U9476 (N_9476,N_3598,N_3608);
nand U9477 (N_9477,N_1557,N_3498);
and U9478 (N_9478,N_5986,N_2899);
nand U9479 (N_9479,N_589,N_5013);
or U9480 (N_9480,N_2935,N_2609);
and U9481 (N_9481,N_1119,N_1257);
nand U9482 (N_9482,N_4332,N_5964);
and U9483 (N_9483,N_5909,N_4219);
nor U9484 (N_9484,N_971,N_5449);
xnor U9485 (N_9485,N_3583,N_4401);
and U9486 (N_9486,N_5951,N_5684);
xnor U9487 (N_9487,N_57,N_1826);
xnor U9488 (N_9488,N_1982,N_3560);
or U9489 (N_9489,N_4363,N_203);
xor U9490 (N_9490,N_1645,N_4123);
nand U9491 (N_9491,N_77,N_418);
or U9492 (N_9492,N_1280,N_3792);
nor U9493 (N_9493,N_4160,N_5033);
xnor U9494 (N_9494,N_3334,N_965);
nor U9495 (N_9495,N_5898,N_1335);
or U9496 (N_9496,N_1246,N_5211);
and U9497 (N_9497,N_877,N_5127);
or U9498 (N_9498,N_2117,N_5978);
nor U9499 (N_9499,N_1385,N_5305);
or U9500 (N_9500,N_4635,N_876);
and U9501 (N_9501,N_1037,N_385);
xnor U9502 (N_9502,N_136,N_2789);
and U9503 (N_9503,N_937,N_2192);
and U9504 (N_9504,N_3199,N_3729);
and U9505 (N_9505,N_5572,N_4342);
or U9506 (N_9506,N_5551,N_1677);
xor U9507 (N_9507,N_4239,N_5117);
nor U9508 (N_9508,N_60,N_506);
or U9509 (N_9509,N_4221,N_1142);
and U9510 (N_9510,N_2636,N_469);
nor U9511 (N_9511,N_838,N_4265);
xnor U9512 (N_9512,N_4312,N_5668);
nor U9513 (N_9513,N_2753,N_5597);
xor U9514 (N_9514,N_3751,N_3504);
and U9515 (N_9515,N_4674,N_2183);
and U9516 (N_9516,N_3505,N_3737);
and U9517 (N_9517,N_2804,N_5637);
nor U9518 (N_9518,N_5030,N_4202);
xnor U9519 (N_9519,N_572,N_4574);
xnor U9520 (N_9520,N_2669,N_5443);
nand U9521 (N_9521,N_4253,N_4602);
nor U9522 (N_9522,N_5077,N_278);
nand U9523 (N_9523,N_3636,N_4249);
xnor U9524 (N_9524,N_2233,N_5944);
or U9525 (N_9525,N_763,N_2102);
xor U9526 (N_9526,N_4831,N_2811);
or U9527 (N_9527,N_17,N_1504);
nand U9528 (N_9528,N_3334,N_839);
xor U9529 (N_9529,N_4137,N_2547);
nor U9530 (N_9530,N_3675,N_1094);
or U9531 (N_9531,N_1133,N_2305);
or U9532 (N_9532,N_1317,N_154);
nand U9533 (N_9533,N_4817,N_3815);
nor U9534 (N_9534,N_5203,N_3788);
and U9535 (N_9535,N_2060,N_3237);
or U9536 (N_9536,N_582,N_5897);
xnor U9537 (N_9537,N_1118,N_851);
and U9538 (N_9538,N_5629,N_4464);
or U9539 (N_9539,N_2528,N_3208);
nand U9540 (N_9540,N_2273,N_4402);
xor U9541 (N_9541,N_3036,N_2812);
nand U9542 (N_9542,N_4432,N_2178);
xor U9543 (N_9543,N_1588,N_1752);
nand U9544 (N_9544,N_2213,N_813);
xnor U9545 (N_9545,N_4165,N_1737);
nand U9546 (N_9546,N_1289,N_2885);
and U9547 (N_9547,N_5894,N_4716);
and U9548 (N_9548,N_5969,N_5458);
nor U9549 (N_9549,N_5832,N_1046);
nand U9550 (N_9550,N_133,N_1647);
and U9551 (N_9551,N_3859,N_1822);
nor U9552 (N_9552,N_5561,N_3257);
and U9553 (N_9553,N_4469,N_4954);
nand U9554 (N_9554,N_5242,N_2569);
nor U9555 (N_9555,N_123,N_1059);
nor U9556 (N_9556,N_1256,N_4698);
nor U9557 (N_9557,N_470,N_370);
nand U9558 (N_9558,N_1425,N_4811);
and U9559 (N_9559,N_4625,N_1636);
nand U9560 (N_9560,N_4672,N_3237);
and U9561 (N_9561,N_5752,N_3009);
xor U9562 (N_9562,N_2855,N_2963);
xnor U9563 (N_9563,N_5468,N_5544);
nand U9564 (N_9564,N_1790,N_5480);
or U9565 (N_9565,N_1987,N_3059);
nand U9566 (N_9566,N_4142,N_647);
nor U9567 (N_9567,N_2142,N_5754);
and U9568 (N_9568,N_474,N_4538);
nor U9569 (N_9569,N_1900,N_4321);
nand U9570 (N_9570,N_3555,N_3189);
nor U9571 (N_9571,N_3496,N_4266);
nor U9572 (N_9572,N_3362,N_5634);
xnor U9573 (N_9573,N_1266,N_5696);
nor U9574 (N_9574,N_3664,N_1091);
nor U9575 (N_9575,N_3572,N_3327);
nor U9576 (N_9576,N_1747,N_2664);
and U9577 (N_9577,N_1388,N_119);
xnor U9578 (N_9578,N_5315,N_236);
and U9579 (N_9579,N_867,N_4980);
or U9580 (N_9580,N_4037,N_5664);
nor U9581 (N_9581,N_434,N_4407);
nor U9582 (N_9582,N_912,N_1555);
and U9583 (N_9583,N_5199,N_2741);
nor U9584 (N_9584,N_4059,N_685);
xnor U9585 (N_9585,N_4558,N_4320);
nand U9586 (N_9586,N_5999,N_4962);
or U9587 (N_9587,N_2104,N_663);
nand U9588 (N_9588,N_5116,N_103);
or U9589 (N_9589,N_3485,N_1194);
xnor U9590 (N_9590,N_1862,N_5736);
and U9591 (N_9591,N_1464,N_2123);
nor U9592 (N_9592,N_1583,N_4366);
nor U9593 (N_9593,N_1144,N_1562);
or U9594 (N_9594,N_3234,N_3275);
nor U9595 (N_9595,N_2288,N_2760);
nor U9596 (N_9596,N_720,N_4741);
and U9597 (N_9597,N_3288,N_2836);
nor U9598 (N_9598,N_2697,N_49);
nor U9599 (N_9599,N_2398,N_374);
nand U9600 (N_9600,N_820,N_4538);
or U9601 (N_9601,N_5585,N_2867);
xnor U9602 (N_9602,N_3569,N_4588);
and U9603 (N_9603,N_1174,N_4455);
or U9604 (N_9604,N_264,N_2456);
nand U9605 (N_9605,N_2296,N_808);
nand U9606 (N_9606,N_1595,N_3916);
nor U9607 (N_9607,N_2487,N_1872);
nor U9608 (N_9608,N_2964,N_4170);
or U9609 (N_9609,N_2276,N_5479);
nor U9610 (N_9610,N_4461,N_2839);
and U9611 (N_9611,N_3614,N_3163);
and U9612 (N_9612,N_2744,N_857);
and U9613 (N_9613,N_4464,N_2111);
or U9614 (N_9614,N_5422,N_3940);
nand U9615 (N_9615,N_2977,N_5103);
nor U9616 (N_9616,N_5728,N_4541);
nor U9617 (N_9617,N_4276,N_3494);
nand U9618 (N_9618,N_5037,N_730);
nor U9619 (N_9619,N_3442,N_4150);
or U9620 (N_9620,N_1953,N_2136);
or U9621 (N_9621,N_1177,N_4219);
nand U9622 (N_9622,N_5857,N_1205);
and U9623 (N_9623,N_1543,N_2688);
or U9624 (N_9624,N_4813,N_1935);
xnor U9625 (N_9625,N_2895,N_5797);
or U9626 (N_9626,N_3196,N_5363);
xor U9627 (N_9627,N_188,N_1753);
or U9628 (N_9628,N_5781,N_2406);
nand U9629 (N_9629,N_1774,N_4030);
nor U9630 (N_9630,N_4525,N_5360);
xnor U9631 (N_9631,N_5454,N_813);
nand U9632 (N_9632,N_3045,N_1165);
and U9633 (N_9633,N_3451,N_2872);
nor U9634 (N_9634,N_2209,N_5200);
xor U9635 (N_9635,N_2429,N_5673);
nand U9636 (N_9636,N_1161,N_196);
nor U9637 (N_9637,N_4902,N_3288);
or U9638 (N_9638,N_3747,N_5523);
nor U9639 (N_9639,N_5822,N_5055);
xnor U9640 (N_9640,N_3780,N_4328);
nor U9641 (N_9641,N_4667,N_4489);
or U9642 (N_9642,N_915,N_5030);
or U9643 (N_9643,N_29,N_2838);
nand U9644 (N_9644,N_1062,N_3957);
nor U9645 (N_9645,N_2117,N_3583);
and U9646 (N_9646,N_5090,N_2398);
nand U9647 (N_9647,N_451,N_610);
and U9648 (N_9648,N_347,N_1210);
or U9649 (N_9649,N_5677,N_3931);
nor U9650 (N_9650,N_892,N_4963);
nand U9651 (N_9651,N_1646,N_2643);
and U9652 (N_9652,N_5309,N_4677);
nand U9653 (N_9653,N_2660,N_744);
nand U9654 (N_9654,N_2786,N_197);
xnor U9655 (N_9655,N_5670,N_1229);
nand U9656 (N_9656,N_1916,N_1174);
and U9657 (N_9657,N_1107,N_3697);
nand U9658 (N_9658,N_2535,N_1304);
or U9659 (N_9659,N_5867,N_51);
or U9660 (N_9660,N_3201,N_1939);
nor U9661 (N_9661,N_2847,N_5280);
and U9662 (N_9662,N_684,N_4042);
xnor U9663 (N_9663,N_4104,N_425);
nor U9664 (N_9664,N_5937,N_2302);
or U9665 (N_9665,N_1764,N_3577);
or U9666 (N_9666,N_915,N_3273);
and U9667 (N_9667,N_3824,N_194);
nor U9668 (N_9668,N_3632,N_2673);
or U9669 (N_9669,N_3987,N_1453);
nand U9670 (N_9670,N_4839,N_1720);
nand U9671 (N_9671,N_2466,N_5821);
xnor U9672 (N_9672,N_639,N_2685);
nand U9673 (N_9673,N_3989,N_19);
nand U9674 (N_9674,N_1264,N_2370);
nor U9675 (N_9675,N_4388,N_3016);
and U9676 (N_9676,N_1748,N_4748);
nor U9677 (N_9677,N_3231,N_4533);
and U9678 (N_9678,N_3454,N_5898);
or U9679 (N_9679,N_4915,N_2846);
nand U9680 (N_9680,N_2099,N_2915);
nand U9681 (N_9681,N_5960,N_5740);
nor U9682 (N_9682,N_5518,N_1149);
or U9683 (N_9683,N_2113,N_2838);
or U9684 (N_9684,N_963,N_2426);
nand U9685 (N_9685,N_245,N_2687);
nor U9686 (N_9686,N_2824,N_2352);
nand U9687 (N_9687,N_1413,N_1159);
nand U9688 (N_9688,N_1351,N_1788);
xor U9689 (N_9689,N_4459,N_5807);
or U9690 (N_9690,N_823,N_1201);
xor U9691 (N_9691,N_3895,N_3780);
or U9692 (N_9692,N_2255,N_1851);
nor U9693 (N_9693,N_2040,N_5889);
and U9694 (N_9694,N_3422,N_5016);
nor U9695 (N_9695,N_2668,N_3141);
xnor U9696 (N_9696,N_4739,N_2613);
or U9697 (N_9697,N_1397,N_4201);
xor U9698 (N_9698,N_5786,N_727);
or U9699 (N_9699,N_4653,N_5980);
or U9700 (N_9700,N_1498,N_5482);
nand U9701 (N_9701,N_1985,N_4121);
and U9702 (N_9702,N_2199,N_3117);
and U9703 (N_9703,N_3373,N_3688);
and U9704 (N_9704,N_3715,N_668);
nand U9705 (N_9705,N_5895,N_740);
and U9706 (N_9706,N_586,N_1846);
and U9707 (N_9707,N_3798,N_1641);
nor U9708 (N_9708,N_3989,N_4568);
nor U9709 (N_9709,N_3041,N_4648);
nor U9710 (N_9710,N_3136,N_4123);
and U9711 (N_9711,N_1545,N_2280);
nor U9712 (N_9712,N_577,N_701);
xnor U9713 (N_9713,N_3357,N_3282);
or U9714 (N_9714,N_764,N_5315);
or U9715 (N_9715,N_5680,N_495);
xnor U9716 (N_9716,N_1801,N_3589);
and U9717 (N_9717,N_3169,N_5997);
nand U9718 (N_9718,N_4464,N_171);
or U9719 (N_9719,N_4416,N_2693);
xor U9720 (N_9720,N_2318,N_1272);
nor U9721 (N_9721,N_2031,N_2487);
xnor U9722 (N_9722,N_1600,N_1755);
nand U9723 (N_9723,N_3352,N_2155);
nor U9724 (N_9724,N_5572,N_953);
nand U9725 (N_9725,N_4284,N_727);
nand U9726 (N_9726,N_2379,N_851);
or U9727 (N_9727,N_2925,N_5871);
and U9728 (N_9728,N_3362,N_3922);
xnor U9729 (N_9729,N_3876,N_5966);
nand U9730 (N_9730,N_1257,N_5954);
nand U9731 (N_9731,N_4532,N_426);
nand U9732 (N_9732,N_2581,N_4808);
and U9733 (N_9733,N_850,N_2835);
nor U9734 (N_9734,N_4448,N_1064);
and U9735 (N_9735,N_3761,N_4322);
and U9736 (N_9736,N_1400,N_5187);
nand U9737 (N_9737,N_3898,N_3056);
xor U9738 (N_9738,N_3559,N_3002);
or U9739 (N_9739,N_2687,N_3180);
and U9740 (N_9740,N_1934,N_4833);
or U9741 (N_9741,N_4352,N_5250);
xnor U9742 (N_9742,N_3649,N_1790);
nor U9743 (N_9743,N_3753,N_2202);
and U9744 (N_9744,N_4162,N_792);
nor U9745 (N_9745,N_1457,N_5659);
xnor U9746 (N_9746,N_3710,N_2011);
nor U9747 (N_9747,N_3059,N_4987);
nor U9748 (N_9748,N_5770,N_5116);
or U9749 (N_9749,N_5525,N_3371);
xor U9750 (N_9750,N_2563,N_5167);
and U9751 (N_9751,N_1004,N_2734);
nand U9752 (N_9752,N_1819,N_4592);
nand U9753 (N_9753,N_2328,N_773);
and U9754 (N_9754,N_282,N_1235);
nor U9755 (N_9755,N_5347,N_4884);
and U9756 (N_9756,N_5243,N_453);
nor U9757 (N_9757,N_4350,N_2614);
or U9758 (N_9758,N_701,N_3253);
and U9759 (N_9759,N_3460,N_2154);
xnor U9760 (N_9760,N_5879,N_345);
xnor U9761 (N_9761,N_2055,N_4137);
or U9762 (N_9762,N_416,N_5235);
nor U9763 (N_9763,N_4032,N_2372);
xor U9764 (N_9764,N_1260,N_2204);
nor U9765 (N_9765,N_2181,N_1032);
nand U9766 (N_9766,N_3618,N_4890);
nand U9767 (N_9767,N_5565,N_2658);
nand U9768 (N_9768,N_844,N_2852);
xor U9769 (N_9769,N_386,N_1229);
nand U9770 (N_9770,N_1505,N_5006);
xnor U9771 (N_9771,N_5605,N_943);
nor U9772 (N_9772,N_1255,N_2626);
nor U9773 (N_9773,N_4232,N_2790);
nand U9774 (N_9774,N_5794,N_80);
xor U9775 (N_9775,N_5704,N_1117);
or U9776 (N_9776,N_2279,N_2715);
and U9777 (N_9777,N_3454,N_2007);
nor U9778 (N_9778,N_3392,N_5797);
and U9779 (N_9779,N_2374,N_4469);
and U9780 (N_9780,N_895,N_997);
nor U9781 (N_9781,N_5960,N_5892);
and U9782 (N_9782,N_1805,N_5094);
and U9783 (N_9783,N_2787,N_3124);
nand U9784 (N_9784,N_2720,N_3758);
nor U9785 (N_9785,N_3411,N_2611);
and U9786 (N_9786,N_5409,N_4818);
nand U9787 (N_9787,N_5374,N_4235);
xnor U9788 (N_9788,N_407,N_1871);
nand U9789 (N_9789,N_4267,N_206);
or U9790 (N_9790,N_2206,N_3363);
nor U9791 (N_9791,N_4751,N_3624);
xnor U9792 (N_9792,N_5352,N_1390);
nor U9793 (N_9793,N_1392,N_1348);
or U9794 (N_9794,N_1954,N_26);
nor U9795 (N_9795,N_2648,N_3874);
and U9796 (N_9796,N_5043,N_3286);
nor U9797 (N_9797,N_20,N_4790);
xnor U9798 (N_9798,N_547,N_2271);
or U9799 (N_9799,N_3079,N_5481);
and U9800 (N_9800,N_3165,N_4728);
nor U9801 (N_9801,N_4035,N_3712);
and U9802 (N_9802,N_916,N_1904);
and U9803 (N_9803,N_3739,N_3553);
xnor U9804 (N_9804,N_3752,N_59);
or U9805 (N_9805,N_2852,N_1690);
and U9806 (N_9806,N_3321,N_3835);
or U9807 (N_9807,N_4659,N_2179);
nand U9808 (N_9808,N_3097,N_3865);
nor U9809 (N_9809,N_3484,N_1626);
and U9810 (N_9810,N_4266,N_5394);
or U9811 (N_9811,N_1927,N_516);
or U9812 (N_9812,N_3795,N_4246);
xnor U9813 (N_9813,N_2476,N_1001);
xor U9814 (N_9814,N_1496,N_5484);
nor U9815 (N_9815,N_1649,N_5913);
and U9816 (N_9816,N_905,N_5859);
nor U9817 (N_9817,N_4476,N_5059);
nand U9818 (N_9818,N_2755,N_4370);
xor U9819 (N_9819,N_3112,N_2739);
nor U9820 (N_9820,N_2809,N_4934);
or U9821 (N_9821,N_893,N_5753);
nor U9822 (N_9822,N_1419,N_4372);
nor U9823 (N_9823,N_21,N_4570);
nand U9824 (N_9824,N_1789,N_4236);
xnor U9825 (N_9825,N_521,N_2680);
and U9826 (N_9826,N_2855,N_4118);
xnor U9827 (N_9827,N_755,N_1808);
xor U9828 (N_9828,N_2589,N_4018);
or U9829 (N_9829,N_3586,N_2911);
and U9830 (N_9830,N_5882,N_4596);
xor U9831 (N_9831,N_4764,N_4725);
nor U9832 (N_9832,N_1357,N_4324);
nor U9833 (N_9833,N_49,N_2057);
nor U9834 (N_9834,N_878,N_5559);
or U9835 (N_9835,N_3362,N_3557);
xor U9836 (N_9836,N_3435,N_2528);
or U9837 (N_9837,N_891,N_473);
or U9838 (N_9838,N_363,N_3148);
or U9839 (N_9839,N_4855,N_690);
nand U9840 (N_9840,N_21,N_110);
nor U9841 (N_9841,N_1503,N_3966);
and U9842 (N_9842,N_2250,N_600);
or U9843 (N_9843,N_4706,N_4628);
nor U9844 (N_9844,N_1783,N_4144);
nand U9845 (N_9845,N_3144,N_4693);
or U9846 (N_9846,N_1118,N_1085);
and U9847 (N_9847,N_315,N_3868);
xor U9848 (N_9848,N_4741,N_2169);
and U9849 (N_9849,N_1355,N_5740);
xor U9850 (N_9850,N_2416,N_4048);
or U9851 (N_9851,N_3743,N_2113);
xnor U9852 (N_9852,N_4931,N_3587);
xnor U9853 (N_9853,N_3117,N_1369);
xor U9854 (N_9854,N_1137,N_4407);
nand U9855 (N_9855,N_5687,N_2417);
nor U9856 (N_9856,N_4495,N_2476);
and U9857 (N_9857,N_661,N_140);
xor U9858 (N_9858,N_5554,N_5232);
nand U9859 (N_9859,N_3825,N_439);
nor U9860 (N_9860,N_1506,N_101);
or U9861 (N_9861,N_2800,N_4285);
xnor U9862 (N_9862,N_3199,N_2825);
nor U9863 (N_9863,N_3756,N_3843);
nor U9864 (N_9864,N_257,N_961);
and U9865 (N_9865,N_1509,N_541);
nor U9866 (N_9866,N_4112,N_1927);
or U9867 (N_9867,N_1342,N_5438);
xor U9868 (N_9868,N_1691,N_1545);
nand U9869 (N_9869,N_5005,N_2968);
xnor U9870 (N_9870,N_3122,N_5176);
xor U9871 (N_9871,N_3107,N_3869);
nor U9872 (N_9872,N_4729,N_1104);
or U9873 (N_9873,N_4055,N_3619);
nand U9874 (N_9874,N_3399,N_1025);
and U9875 (N_9875,N_3878,N_2070);
or U9876 (N_9876,N_4924,N_3960);
or U9877 (N_9877,N_3569,N_4746);
and U9878 (N_9878,N_1469,N_4054);
nand U9879 (N_9879,N_3954,N_3535);
xor U9880 (N_9880,N_1727,N_5228);
xnor U9881 (N_9881,N_1891,N_4518);
nand U9882 (N_9882,N_3236,N_3272);
nor U9883 (N_9883,N_3251,N_4034);
xor U9884 (N_9884,N_608,N_1007);
or U9885 (N_9885,N_571,N_5099);
and U9886 (N_9886,N_2906,N_2180);
or U9887 (N_9887,N_2253,N_5123);
nor U9888 (N_9888,N_1336,N_2360);
nand U9889 (N_9889,N_2737,N_4849);
nor U9890 (N_9890,N_3196,N_1923);
nor U9891 (N_9891,N_4372,N_5716);
or U9892 (N_9892,N_2986,N_4992);
xor U9893 (N_9893,N_5616,N_3378);
or U9894 (N_9894,N_1337,N_3693);
nand U9895 (N_9895,N_5472,N_430);
nand U9896 (N_9896,N_286,N_4450);
xnor U9897 (N_9897,N_1859,N_3111);
xor U9898 (N_9898,N_5175,N_1129);
nand U9899 (N_9899,N_5404,N_4152);
xnor U9900 (N_9900,N_1556,N_4019);
nand U9901 (N_9901,N_5119,N_2010);
or U9902 (N_9902,N_1571,N_1274);
xor U9903 (N_9903,N_1825,N_5930);
nor U9904 (N_9904,N_5494,N_3209);
nand U9905 (N_9905,N_3724,N_2539);
or U9906 (N_9906,N_374,N_1376);
nand U9907 (N_9907,N_2390,N_2459);
nand U9908 (N_9908,N_3949,N_1746);
and U9909 (N_9909,N_2283,N_1018);
or U9910 (N_9910,N_1466,N_3928);
or U9911 (N_9911,N_3069,N_2890);
and U9912 (N_9912,N_3132,N_473);
and U9913 (N_9913,N_2858,N_3645);
xor U9914 (N_9914,N_1108,N_2282);
nor U9915 (N_9915,N_5170,N_3492);
and U9916 (N_9916,N_5166,N_933);
nand U9917 (N_9917,N_700,N_3281);
and U9918 (N_9918,N_464,N_3871);
xor U9919 (N_9919,N_5895,N_4264);
nand U9920 (N_9920,N_4413,N_2151);
nand U9921 (N_9921,N_3800,N_2430);
xor U9922 (N_9922,N_4732,N_3052);
xnor U9923 (N_9923,N_2831,N_2290);
and U9924 (N_9924,N_692,N_94);
or U9925 (N_9925,N_3585,N_2038);
or U9926 (N_9926,N_5019,N_4388);
or U9927 (N_9927,N_5838,N_4880);
nand U9928 (N_9928,N_442,N_1116);
nand U9929 (N_9929,N_4324,N_5205);
xor U9930 (N_9930,N_4846,N_759);
or U9931 (N_9931,N_4447,N_3808);
and U9932 (N_9932,N_1833,N_1642);
or U9933 (N_9933,N_1641,N_1827);
nor U9934 (N_9934,N_2813,N_2581);
and U9935 (N_9935,N_5805,N_3537);
nand U9936 (N_9936,N_5247,N_1177);
xnor U9937 (N_9937,N_1507,N_4236);
or U9938 (N_9938,N_4858,N_3256);
nand U9939 (N_9939,N_3489,N_2285);
or U9940 (N_9940,N_4953,N_137);
xnor U9941 (N_9941,N_5004,N_3014);
and U9942 (N_9942,N_4517,N_522);
and U9943 (N_9943,N_2549,N_1757);
or U9944 (N_9944,N_2869,N_4153);
or U9945 (N_9945,N_3176,N_2683);
xor U9946 (N_9946,N_382,N_4061);
nand U9947 (N_9947,N_782,N_5703);
nor U9948 (N_9948,N_4801,N_3797);
and U9949 (N_9949,N_4795,N_4881);
and U9950 (N_9950,N_3930,N_3149);
or U9951 (N_9951,N_2735,N_5621);
nand U9952 (N_9952,N_1856,N_5703);
xor U9953 (N_9953,N_2357,N_5206);
or U9954 (N_9954,N_3142,N_4910);
xnor U9955 (N_9955,N_452,N_1159);
xor U9956 (N_9956,N_283,N_5662);
nor U9957 (N_9957,N_2304,N_4175);
nor U9958 (N_9958,N_654,N_2553);
nand U9959 (N_9959,N_163,N_114);
xnor U9960 (N_9960,N_1156,N_3578);
or U9961 (N_9961,N_95,N_796);
xor U9962 (N_9962,N_1773,N_873);
nand U9963 (N_9963,N_4373,N_1473);
and U9964 (N_9964,N_2088,N_1238);
nand U9965 (N_9965,N_4003,N_2314);
nor U9966 (N_9966,N_4620,N_5068);
nand U9967 (N_9967,N_5343,N_5034);
nand U9968 (N_9968,N_479,N_340);
nand U9969 (N_9969,N_2920,N_4095);
nor U9970 (N_9970,N_3089,N_4967);
or U9971 (N_9971,N_768,N_2100);
nand U9972 (N_9972,N_5705,N_1222);
nand U9973 (N_9973,N_174,N_3132);
xor U9974 (N_9974,N_3088,N_4183);
nand U9975 (N_9975,N_2479,N_3233);
and U9976 (N_9976,N_2707,N_493);
xor U9977 (N_9977,N_3302,N_186);
xnor U9978 (N_9978,N_5994,N_3781);
nand U9979 (N_9979,N_3096,N_3414);
xor U9980 (N_9980,N_5295,N_1088);
xor U9981 (N_9981,N_2006,N_2734);
xnor U9982 (N_9982,N_2693,N_1316);
xnor U9983 (N_9983,N_3396,N_1079);
nor U9984 (N_9984,N_793,N_5784);
or U9985 (N_9985,N_509,N_4685);
xor U9986 (N_9986,N_3250,N_4124);
nor U9987 (N_9987,N_5447,N_975);
nor U9988 (N_9988,N_3966,N_168);
and U9989 (N_9989,N_5169,N_337);
or U9990 (N_9990,N_1932,N_1941);
or U9991 (N_9991,N_4989,N_1981);
and U9992 (N_9992,N_3424,N_1767);
nor U9993 (N_9993,N_4983,N_695);
and U9994 (N_9994,N_4238,N_3355);
xnor U9995 (N_9995,N_991,N_4956);
or U9996 (N_9996,N_1484,N_1073);
nand U9997 (N_9997,N_3596,N_3035);
and U9998 (N_9998,N_4688,N_1302);
nor U9999 (N_9999,N_3194,N_5716);
nor U10000 (N_10000,N_2168,N_3938);
nor U10001 (N_10001,N_5279,N_4369);
or U10002 (N_10002,N_5652,N_2330);
or U10003 (N_10003,N_873,N_1951);
nor U10004 (N_10004,N_1012,N_4847);
nand U10005 (N_10005,N_3293,N_1383);
xnor U10006 (N_10006,N_4692,N_2961);
nor U10007 (N_10007,N_960,N_1724);
and U10008 (N_10008,N_2162,N_3613);
nor U10009 (N_10009,N_4291,N_5741);
nor U10010 (N_10010,N_5490,N_5297);
xor U10011 (N_10011,N_316,N_1268);
nand U10012 (N_10012,N_5210,N_2508);
nor U10013 (N_10013,N_534,N_2037);
and U10014 (N_10014,N_4278,N_3201);
and U10015 (N_10015,N_3074,N_718);
nand U10016 (N_10016,N_4559,N_5318);
or U10017 (N_10017,N_2693,N_908);
nand U10018 (N_10018,N_958,N_1874);
and U10019 (N_10019,N_5952,N_5916);
nand U10020 (N_10020,N_73,N_5631);
nor U10021 (N_10021,N_269,N_2659);
and U10022 (N_10022,N_4065,N_176);
or U10023 (N_10023,N_3783,N_3310);
xnor U10024 (N_10024,N_4234,N_2324);
nor U10025 (N_10025,N_5727,N_3993);
or U10026 (N_10026,N_5939,N_40);
and U10027 (N_10027,N_5458,N_4826);
nand U10028 (N_10028,N_2208,N_2571);
nor U10029 (N_10029,N_3259,N_5671);
nor U10030 (N_10030,N_4956,N_4333);
xnor U10031 (N_10031,N_2529,N_5998);
nand U10032 (N_10032,N_4841,N_5502);
or U10033 (N_10033,N_5993,N_3011);
nor U10034 (N_10034,N_686,N_3049);
nand U10035 (N_10035,N_3828,N_5108);
nand U10036 (N_10036,N_1508,N_680);
nand U10037 (N_10037,N_1457,N_1461);
xor U10038 (N_10038,N_1656,N_4808);
nand U10039 (N_10039,N_5542,N_2060);
xor U10040 (N_10040,N_1388,N_2841);
nand U10041 (N_10041,N_2719,N_5708);
or U10042 (N_10042,N_2176,N_2969);
nand U10043 (N_10043,N_2598,N_1740);
nand U10044 (N_10044,N_5749,N_2202);
or U10045 (N_10045,N_3681,N_1360);
nor U10046 (N_10046,N_2873,N_2316);
and U10047 (N_10047,N_1711,N_2760);
xnor U10048 (N_10048,N_952,N_3022);
nand U10049 (N_10049,N_3076,N_4671);
nand U10050 (N_10050,N_5227,N_498);
xor U10051 (N_10051,N_1554,N_3538);
and U10052 (N_10052,N_169,N_1096);
or U10053 (N_10053,N_4975,N_1336);
nor U10054 (N_10054,N_4198,N_411);
nor U10055 (N_10055,N_2858,N_3280);
and U10056 (N_10056,N_2627,N_2415);
xor U10057 (N_10057,N_1377,N_5822);
nor U10058 (N_10058,N_2520,N_80);
and U10059 (N_10059,N_1853,N_4980);
nor U10060 (N_10060,N_5260,N_4463);
nand U10061 (N_10061,N_5220,N_99);
xor U10062 (N_10062,N_2583,N_229);
and U10063 (N_10063,N_834,N_1680);
nor U10064 (N_10064,N_3284,N_1641);
xor U10065 (N_10065,N_511,N_3602);
nand U10066 (N_10066,N_2990,N_1865);
nor U10067 (N_10067,N_5413,N_1869);
or U10068 (N_10068,N_5073,N_2022);
nand U10069 (N_10069,N_2318,N_1303);
xnor U10070 (N_10070,N_2381,N_3982);
xnor U10071 (N_10071,N_1987,N_4757);
xnor U10072 (N_10072,N_3162,N_1935);
nand U10073 (N_10073,N_113,N_4770);
and U10074 (N_10074,N_4596,N_4189);
and U10075 (N_10075,N_4818,N_879);
nor U10076 (N_10076,N_1231,N_4478);
and U10077 (N_10077,N_4322,N_3124);
nor U10078 (N_10078,N_3357,N_4551);
or U10079 (N_10079,N_1816,N_910);
or U10080 (N_10080,N_5574,N_4399);
xnor U10081 (N_10081,N_2910,N_3603);
xnor U10082 (N_10082,N_4226,N_4595);
nand U10083 (N_10083,N_5673,N_3157);
or U10084 (N_10084,N_109,N_43);
nand U10085 (N_10085,N_3998,N_2964);
or U10086 (N_10086,N_3268,N_3732);
or U10087 (N_10087,N_244,N_2593);
and U10088 (N_10088,N_1902,N_2918);
and U10089 (N_10089,N_2911,N_2167);
xnor U10090 (N_10090,N_3219,N_2777);
and U10091 (N_10091,N_4535,N_3257);
or U10092 (N_10092,N_5013,N_1222);
nand U10093 (N_10093,N_2874,N_2055);
and U10094 (N_10094,N_1887,N_699);
or U10095 (N_10095,N_5355,N_4671);
nor U10096 (N_10096,N_4695,N_3635);
nand U10097 (N_10097,N_4698,N_1709);
nand U10098 (N_10098,N_2733,N_3524);
or U10099 (N_10099,N_2366,N_3716);
and U10100 (N_10100,N_5719,N_1100);
and U10101 (N_10101,N_3460,N_4856);
nor U10102 (N_10102,N_113,N_4271);
and U10103 (N_10103,N_3125,N_998);
nor U10104 (N_10104,N_353,N_4055);
or U10105 (N_10105,N_60,N_3863);
or U10106 (N_10106,N_2386,N_4758);
nor U10107 (N_10107,N_4670,N_226);
nor U10108 (N_10108,N_1602,N_5349);
xnor U10109 (N_10109,N_3556,N_2722);
or U10110 (N_10110,N_597,N_1588);
or U10111 (N_10111,N_5439,N_3379);
and U10112 (N_10112,N_3618,N_382);
nor U10113 (N_10113,N_2371,N_4733);
and U10114 (N_10114,N_1474,N_2753);
nor U10115 (N_10115,N_5323,N_3904);
and U10116 (N_10116,N_4399,N_4132);
or U10117 (N_10117,N_2196,N_3462);
xnor U10118 (N_10118,N_4702,N_2585);
nor U10119 (N_10119,N_1174,N_4442);
nand U10120 (N_10120,N_2723,N_1260);
nor U10121 (N_10121,N_2760,N_3490);
or U10122 (N_10122,N_1464,N_253);
xnor U10123 (N_10123,N_3181,N_5949);
or U10124 (N_10124,N_4444,N_287);
nor U10125 (N_10125,N_5136,N_3337);
and U10126 (N_10126,N_3676,N_2898);
nand U10127 (N_10127,N_4079,N_4035);
nor U10128 (N_10128,N_1917,N_4848);
or U10129 (N_10129,N_5671,N_5029);
xor U10130 (N_10130,N_3527,N_752);
or U10131 (N_10131,N_5559,N_5745);
or U10132 (N_10132,N_4634,N_5584);
or U10133 (N_10133,N_3378,N_1909);
or U10134 (N_10134,N_2389,N_425);
xnor U10135 (N_10135,N_1948,N_4390);
nor U10136 (N_10136,N_4409,N_999);
or U10137 (N_10137,N_383,N_766);
nor U10138 (N_10138,N_3838,N_1965);
nand U10139 (N_10139,N_4593,N_1085);
nand U10140 (N_10140,N_4036,N_2592);
and U10141 (N_10141,N_3590,N_1057);
and U10142 (N_10142,N_385,N_2745);
nor U10143 (N_10143,N_4244,N_2214);
and U10144 (N_10144,N_1054,N_5463);
nor U10145 (N_10145,N_2702,N_3228);
xnor U10146 (N_10146,N_4775,N_1338);
or U10147 (N_10147,N_5375,N_878);
nor U10148 (N_10148,N_4926,N_5443);
nor U10149 (N_10149,N_4326,N_4775);
nor U10150 (N_10150,N_5680,N_3287);
or U10151 (N_10151,N_2734,N_3078);
nand U10152 (N_10152,N_334,N_3835);
or U10153 (N_10153,N_11,N_4904);
and U10154 (N_10154,N_5661,N_4533);
or U10155 (N_10155,N_1726,N_2588);
and U10156 (N_10156,N_1362,N_554);
nor U10157 (N_10157,N_327,N_996);
nor U10158 (N_10158,N_5110,N_4204);
nand U10159 (N_10159,N_5618,N_341);
nor U10160 (N_10160,N_1604,N_2018);
and U10161 (N_10161,N_432,N_5721);
nand U10162 (N_10162,N_20,N_2843);
nor U10163 (N_10163,N_5877,N_1648);
nor U10164 (N_10164,N_5335,N_2259);
nand U10165 (N_10165,N_4878,N_4163);
and U10166 (N_10166,N_4481,N_1416);
xnor U10167 (N_10167,N_3516,N_1094);
nor U10168 (N_10168,N_5964,N_1816);
nand U10169 (N_10169,N_3661,N_5039);
xor U10170 (N_10170,N_1137,N_702);
nand U10171 (N_10171,N_4707,N_5269);
or U10172 (N_10172,N_4568,N_4067);
or U10173 (N_10173,N_3577,N_3609);
nor U10174 (N_10174,N_3124,N_3644);
nand U10175 (N_10175,N_5550,N_1887);
and U10176 (N_10176,N_4757,N_4029);
nor U10177 (N_10177,N_1666,N_5565);
nand U10178 (N_10178,N_4995,N_4777);
and U10179 (N_10179,N_4407,N_1018);
xnor U10180 (N_10180,N_3929,N_3288);
or U10181 (N_10181,N_3132,N_2323);
and U10182 (N_10182,N_2169,N_1547);
and U10183 (N_10183,N_5735,N_1253);
xor U10184 (N_10184,N_5270,N_4159);
xnor U10185 (N_10185,N_3398,N_1018);
nor U10186 (N_10186,N_2088,N_219);
xor U10187 (N_10187,N_1191,N_3249);
nand U10188 (N_10188,N_5552,N_21);
nand U10189 (N_10189,N_5955,N_742);
or U10190 (N_10190,N_2933,N_4355);
nor U10191 (N_10191,N_2208,N_5656);
nor U10192 (N_10192,N_920,N_1292);
nand U10193 (N_10193,N_4362,N_4728);
xor U10194 (N_10194,N_1104,N_2266);
and U10195 (N_10195,N_4186,N_4397);
and U10196 (N_10196,N_3693,N_4975);
or U10197 (N_10197,N_4430,N_2561);
nor U10198 (N_10198,N_46,N_5921);
nor U10199 (N_10199,N_4335,N_1959);
nand U10200 (N_10200,N_1590,N_3948);
nand U10201 (N_10201,N_1002,N_4113);
nand U10202 (N_10202,N_2557,N_1392);
and U10203 (N_10203,N_183,N_4929);
nand U10204 (N_10204,N_1591,N_4581);
nand U10205 (N_10205,N_1325,N_1374);
or U10206 (N_10206,N_2542,N_3752);
xor U10207 (N_10207,N_1463,N_5202);
nor U10208 (N_10208,N_2357,N_3828);
and U10209 (N_10209,N_3343,N_1120);
nor U10210 (N_10210,N_1363,N_305);
or U10211 (N_10211,N_863,N_3679);
xnor U10212 (N_10212,N_2611,N_604);
xnor U10213 (N_10213,N_3405,N_1632);
and U10214 (N_10214,N_313,N_374);
nand U10215 (N_10215,N_1935,N_5849);
nand U10216 (N_10216,N_3422,N_5549);
nor U10217 (N_10217,N_5197,N_3446);
nand U10218 (N_10218,N_1884,N_3350);
xnor U10219 (N_10219,N_185,N_2835);
xnor U10220 (N_10220,N_5224,N_3338);
xnor U10221 (N_10221,N_4746,N_4859);
and U10222 (N_10222,N_1984,N_5749);
xnor U10223 (N_10223,N_3535,N_5272);
nor U10224 (N_10224,N_2600,N_3543);
nor U10225 (N_10225,N_3772,N_2459);
and U10226 (N_10226,N_412,N_4177);
and U10227 (N_10227,N_2391,N_2377);
and U10228 (N_10228,N_4971,N_2019);
nor U10229 (N_10229,N_5930,N_5226);
and U10230 (N_10230,N_3888,N_180);
or U10231 (N_10231,N_1444,N_2064);
xnor U10232 (N_10232,N_4675,N_233);
xnor U10233 (N_10233,N_5513,N_4677);
nand U10234 (N_10234,N_5926,N_5771);
xnor U10235 (N_10235,N_2641,N_2079);
and U10236 (N_10236,N_4099,N_2375);
or U10237 (N_10237,N_1364,N_2925);
nand U10238 (N_10238,N_3946,N_3629);
xnor U10239 (N_10239,N_1028,N_2518);
or U10240 (N_10240,N_906,N_2914);
and U10241 (N_10241,N_3188,N_476);
or U10242 (N_10242,N_5519,N_4089);
nor U10243 (N_10243,N_1635,N_1398);
nand U10244 (N_10244,N_5923,N_2489);
or U10245 (N_10245,N_1259,N_2898);
and U10246 (N_10246,N_888,N_3503);
nor U10247 (N_10247,N_4285,N_2497);
or U10248 (N_10248,N_3104,N_1757);
nor U10249 (N_10249,N_1026,N_5264);
or U10250 (N_10250,N_2961,N_4941);
xnor U10251 (N_10251,N_1530,N_2079);
nand U10252 (N_10252,N_317,N_1758);
and U10253 (N_10253,N_4439,N_2867);
and U10254 (N_10254,N_4502,N_5607);
nand U10255 (N_10255,N_1123,N_4120);
nor U10256 (N_10256,N_3921,N_5266);
and U10257 (N_10257,N_1581,N_3452);
nor U10258 (N_10258,N_2139,N_949);
and U10259 (N_10259,N_1930,N_4497);
or U10260 (N_10260,N_412,N_4717);
or U10261 (N_10261,N_1436,N_678);
xnor U10262 (N_10262,N_4600,N_2834);
or U10263 (N_10263,N_1803,N_3910);
and U10264 (N_10264,N_3056,N_5835);
nor U10265 (N_10265,N_4939,N_3180);
nor U10266 (N_10266,N_1384,N_2372);
nand U10267 (N_10267,N_2936,N_1683);
xor U10268 (N_10268,N_1123,N_1739);
nor U10269 (N_10269,N_3140,N_3780);
nor U10270 (N_10270,N_5009,N_2057);
or U10271 (N_10271,N_3252,N_4060);
nand U10272 (N_10272,N_4713,N_3966);
and U10273 (N_10273,N_3814,N_4081);
nand U10274 (N_10274,N_5470,N_4595);
and U10275 (N_10275,N_5549,N_5173);
xnor U10276 (N_10276,N_4132,N_3265);
nor U10277 (N_10277,N_5394,N_1045);
and U10278 (N_10278,N_4148,N_656);
and U10279 (N_10279,N_3524,N_3649);
nor U10280 (N_10280,N_1235,N_802);
nor U10281 (N_10281,N_4628,N_3708);
or U10282 (N_10282,N_894,N_3689);
and U10283 (N_10283,N_4949,N_4974);
nor U10284 (N_10284,N_3555,N_2355);
nor U10285 (N_10285,N_2522,N_1178);
and U10286 (N_10286,N_4608,N_3708);
or U10287 (N_10287,N_165,N_2569);
and U10288 (N_10288,N_4340,N_79);
and U10289 (N_10289,N_4401,N_5078);
nor U10290 (N_10290,N_1794,N_566);
nor U10291 (N_10291,N_2698,N_3874);
and U10292 (N_10292,N_4270,N_3423);
nor U10293 (N_10293,N_1034,N_1357);
nand U10294 (N_10294,N_2456,N_989);
xor U10295 (N_10295,N_5247,N_3910);
or U10296 (N_10296,N_1247,N_4239);
nand U10297 (N_10297,N_1067,N_4033);
nand U10298 (N_10298,N_753,N_1443);
xnor U10299 (N_10299,N_43,N_5897);
xnor U10300 (N_10300,N_2710,N_3363);
xnor U10301 (N_10301,N_403,N_4511);
nand U10302 (N_10302,N_436,N_1960);
nand U10303 (N_10303,N_2947,N_3976);
xnor U10304 (N_10304,N_5194,N_14);
nor U10305 (N_10305,N_3048,N_3449);
nor U10306 (N_10306,N_1798,N_153);
xor U10307 (N_10307,N_5852,N_406);
nand U10308 (N_10308,N_4986,N_4925);
and U10309 (N_10309,N_5308,N_1961);
nor U10310 (N_10310,N_1819,N_1649);
nand U10311 (N_10311,N_2022,N_2260);
nor U10312 (N_10312,N_1320,N_3854);
nor U10313 (N_10313,N_744,N_4823);
or U10314 (N_10314,N_963,N_1707);
xnor U10315 (N_10315,N_5613,N_4585);
and U10316 (N_10316,N_2594,N_1964);
or U10317 (N_10317,N_4651,N_5569);
nor U10318 (N_10318,N_4143,N_2029);
or U10319 (N_10319,N_2203,N_553);
or U10320 (N_10320,N_5144,N_4840);
nand U10321 (N_10321,N_4380,N_1771);
nand U10322 (N_10322,N_1486,N_1099);
nand U10323 (N_10323,N_1279,N_125);
nor U10324 (N_10324,N_5254,N_3724);
xnor U10325 (N_10325,N_3070,N_3079);
or U10326 (N_10326,N_5472,N_2624);
nand U10327 (N_10327,N_1871,N_1895);
nor U10328 (N_10328,N_3281,N_5957);
nand U10329 (N_10329,N_1435,N_3775);
nor U10330 (N_10330,N_5433,N_3224);
or U10331 (N_10331,N_3718,N_4196);
nand U10332 (N_10332,N_2124,N_4922);
or U10333 (N_10333,N_4296,N_3330);
and U10334 (N_10334,N_485,N_2357);
or U10335 (N_10335,N_5952,N_4348);
and U10336 (N_10336,N_4275,N_3745);
nor U10337 (N_10337,N_5814,N_4587);
or U10338 (N_10338,N_3630,N_1759);
nor U10339 (N_10339,N_5990,N_4718);
nor U10340 (N_10340,N_2006,N_3056);
and U10341 (N_10341,N_436,N_4868);
or U10342 (N_10342,N_1669,N_1788);
xnor U10343 (N_10343,N_2653,N_227);
nand U10344 (N_10344,N_676,N_2232);
and U10345 (N_10345,N_3454,N_4365);
and U10346 (N_10346,N_4580,N_5680);
nor U10347 (N_10347,N_1998,N_4274);
or U10348 (N_10348,N_3779,N_3414);
nand U10349 (N_10349,N_2459,N_4840);
nor U10350 (N_10350,N_4148,N_1719);
and U10351 (N_10351,N_3692,N_2099);
xnor U10352 (N_10352,N_423,N_5807);
nand U10353 (N_10353,N_5178,N_2216);
xnor U10354 (N_10354,N_5529,N_5280);
xnor U10355 (N_10355,N_2043,N_4233);
xor U10356 (N_10356,N_387,N_792);
nor U10357 (N_10357,N_3847,N_5286);
xnor U10358 (N_10358,N_2845,N_5545);
or U10359 (N_10359,N_1325,N_1168);
xnor U10360 (N_10360,N_3712,N_3778);
xor U10361 (N_10361,N_4397,N_2165);
xnor U10362 (N_10362,N_3973,N_3919);
or U10363 (N_10363,N_4634,N_1209);
nor U10364 (N_10364,N_4664,N_2585);
and U10365 (N_10365,N_2078,N_888);
or U10366 (N_10366,N_1017,N_2683);
nand U10367 (N_10367,N_1489,N_1142);
nor U10368 (N_10368,N_1309,N_5657);
and U10369 (N_10369,N_1821,N_256);
or U10370 (N_10370,N_3483,N_4869);
nor U10371 (N_10371,N_65,N_977);
xor U10372 (N_10372,N_5188,N_3292);
nand U10373 (N_10373,N_4845,N_594);
and U10374 (N_10374,N_3361,N_5329);
nor U10375 (N_10375,N_582,N_734);
xnor U10376 (N_10376,N_692,N_26);
xnor U10377 (N_10377,N_2438,N_1622);
nor U10378 (N_10378,N_5933,N_980);
nor U10379 (N_10379,N_5380,N_1274);
nor U10380 (N_10380,N_3967,N_5249);
xor U10381 (N_10381,N_3493,N_4338);
nand U10382 (N_10382,N_2203,N_5066);
or U10383 (N_10383,N_5419,N_755);
nor U10384 (N_10384,N_527,N_93);
nand U10385 (N_10385,N_4128,N_707);
xor U10386 (N_10386,N_5363,N_2525);
nand U10387 (N_10387,N_5594,N_832);
xor U10388 (N_10388,N_5511,N_5085);
nor U10389 (N_10389,N_3433,N_124);
or U10390 (N_10390,N_3971,N_5178);
xnor U10391 (N_10391,N_5062,N_5235);
nand U10392 (N_10392,N_2414,N_2470);
xor U10393 (N_10393,N_723,N_3317);
nand U10394 (N_10394,N_4088,N_1878);
xor U10395 (N_10395,N_3103,N_130);
xor U10396 (N_10396,N_5764,N_776);
nor U10397 (N_10397,N_4574,N_3196);
nand U10398 (N_10398,N_5816,N_863);
and U10399 (N_10399,N_2447,N_2548);
xnor U10400 (N_10400,N_3763,N_5152);
or U10401 (N_10401,N_4889,N_5658);
nand U10402 (N_10402,N_2038,N_3806);
and U10403 (N_10403,N_4333,N_1174);
nor U10404 (N_10404,N_1083,N_92);
and U10405 (N_10405,N_2591,N_618);
xnor U10406 (N_10406,N_976,N_1652);
nand U10407 (N_10407,N_4624,N_2134);
nor U10408 (N_10408,N_4426,N_4489);
nand U10409 (N_10409,N_3613,N_5185);
and U10410 (N_10410,N_5092,N_1871);
xor U10411 (N_10411,N_5789,N_137);
or U10412 (N_10412,N_2479,N_3941);
nand U10413 (N_10413,N_4073,N_3899);
nand U10414 (N_10414,N_1425,N_4014);
and U10415 (N_10415,N_1801,N_1302);
xnor U10416 (N_10416,N_2298,N_3547);
xor U10417 (N_10417,N_737,N_5174);
nor U10418 (N_10418,N_4128,N_4732);
nor U10419 (N_10419,N_259,N_2699);
and U10420 (N_10420,N_1590,N_3700);
nor U10421 (N_10421,N_5707,N_201);
xnor U10422 (N_10422,N_4798,N_437);
xnor U10423 (N_10423,N_1141,N_3124);
or U10424 (N_10424,N_3163,N_4654);
nor U10425 (N_10425,N_1599,N_2040);
or U10426 (N_10426,N_1417,N_1672);
nand U10427 (N_10427,N_616,N_1109);
and U10428 (N_10428,N_2977,N_284);
nand U10429 (N_10429,N_4038,N_3014);
xnor U10430 (N_10430,N_606,N_1368);
and U10431 (N_10431,N_177,N_4049);
nand U10432 (N_10432,N_4652,N_179);
nor U10433 (N_10433,N_3062,N_2412);
and U10434 (N_10434,N_4194,N_5479);
and U10435 (N_10435,N_5877,N_763);
xnor U10436 (N_10436,N_2611,N_4271);
nor U10437 (N_10437,N_131,N_3158);
xnor U10438 (N_10438,N_1040,N_807);
and U10439 (N_10439,N_358,N_1936);
nand U10440 (N_10440,N_370,N_5032);
nor U10441 (N_10441,N_5333,N_3183);
nor U10442 (N_10442,N_1516,N_4039);
or U10443 (N_10443,N_5858,N_1831);
and U10444 (N_10444,N_3264,N_543);
and U10445 (N_10445,N_4928,N_5696);
nor U10446 (N_10446,N_4378,N_1031);
xor U10447 (N_10447,N_5968,N_545);
nand U10448 (N_10448,N_1919,N_1706);
and U10449 (N_10449,N_2858,N_2487);
or U10450 (N_10450,N_2480,N_2585);
nand U10451 (N_10451,N_667,N_224);
nand U10452 (N_10452,N_5632,N_3029);
and U10453 (N_10453,N_5999,N_552);
nor U10454 (N_10454,N_3928,N_1046);
nor U10455 (N_10455,N_1960,N_1754);
and U10456 (N_10456,N_3955,N_1978);
or U10457 (N_10457,N_1242,N_393);
or U10458 (N_10458,N_502,N_5933);
or U10459 (N_10459,N_3539,N_894);
or U10460 (N_10460,N_4680,N_1597);
xnor U10461 (N_10461,N_3771,N_2352);
xor U10462 (N_10462,N_179,N_2572);
and U10463 (N_10463,N_4900,N_2776);
or U10464 (N_10464,N_3469,N_2650);
nand U10465 (N_10465,N_4249,N_4109);
nand U10466 (N_10466,N_4875,N_1631);
nand U10467 (N_10467,N_5584,N_5603);
nor U10468 (N_10468,N_4553,N_5107);
nor U10469 (N_10469,N_688,N_3021);
nand U10470 (N_10470,N_5885,N_5610);
and U10471 (N_10471,N_1385,N_1971);
and U10472 (N_10472,N_1736,N_2265);
and U10473 (N_10473,N_5199,N_4709);
nand U10474 (N_10474,N_1278,N_2211);
xnor U10475 (N_10475,N_3805,N_85);
xnor U10476 (N_10476,N_795,N_2831);
nor U10477 (N_10477,N_2196,N_5874);
and U10478 (N_10478,N_2649,N_3491);
nor U10479 (N_10479,N_810,N_5996);
nand U10480 (N_10480,N_4698,N_2601);
xor U10481 (N_10481,N_256,N_3747);
and U10482 (N_10482,N_5722,N_2162);
nor U10483 (N_10483,N_863,N_1165);
nand U10484 (N_10484,N_734,N_68);
nor U10485 (N_10485,N_254,N_3326);
or U10486 (N_10486,N_536,N_1173);
or U10487 (N_10487,N_3463,N_5540);
and U10488 (N_10488,N_4592,N_4539);
and U10489 (N_10489,N_1302,N_426);
xor U10490 (N_10490,N_1103,N_2728);
xnor U10491 (N_10491,N_1829,N_4460);
or U10492 (N_10492,N_743,N_2933);
and U10493 (N_10493,N_1148,N_3438);
or U10494 (N_10494,N_2664,N_3692);
xor U10495 (N_10495,N_1256,N_294);
nor U10496 (N_10496,N_2814,N_5424);
nand U10497 (N_10497,N_4853,N_1199);
and U10498 (N_10498,N_577,N_1654);
or U10499 (N_10499,N_1361,N_1349);
or U10500 (N_10500,N_5761,N_4987);
xnor U10501 (N_10501,N_882,N_5867);
and U10502 (N_10502,N_3715,N_4109);
nor U10503 (N_10503,N_195,N_3122);
or U10504 (N_10504,N_5971,N_1239);
or U10505 (N_10505,N_3725,N_2367);
and U10506 (N_10506,N_4689,N_5604);
or U10507 (N_10507,N_4158,N_1858);
nand U10508 (N_10508,N_4405,N_4811);
or U10509 (N_10509,N_555,N_535);
nand U10510 (N_10510,N_4530,N_904);
nor U10511 (N_10511,N_2970,N_3024);
or U10512 (N_10512,N_3734,N_3555);
nor U10513 (N_10513,N_202,N_3847);
nand U10514 (N_10514,N_4802,N_3017);
nand U10515 (N_10515,N_4966,N_2983);
and U10516 (N_10516,N_5803,N_1751);
nand U10517 (N_10517,N_3122,N_961);
nand U10518 (N_10518,N_882,N_519);
or U10519 (N_10519,N_2991,N_4073);
xor U10520 (N_10520,N_4915,N_5052);
nand U10521 (N_10521,N_3738,N_4366);
nand U10522 (N_10522,N_4406,N_1122);
xor U10523 (N_10523,N_2494,N_5875);
nand U10524 (N_10524,N_2631,N_1618);
and U10525 (N_10525,N_4510,N_1315);
and U10526 (N_10526,N_1075,N_3397);
xnor U10527 (N_10527,N_4462,N_1670);
and U10528 (N_10528,N_5757,N_4251);
and U10529 (N_10529,N_76,N_3246);
nor U10530 (N_10530,N_5197,N_1470);
xor U10531 (N_10531,N_4804,N_120);
nor U10532 (N_10532,N_3040,N_3435);
xor U10533 (N_10533,N_4125,N_4860);
nor U10534 (N_10534,N_909,N_4255);
xor U10535 (N_10535,N_166,N_2410);
and U10536 (N_10536,N_4166,N_5401);
nand U10537 (N_10537,N_3030,N_1680);
or U10538 (N_10538,N_5091,N_1864);
nand U10539 (N_10539,N_4466,N_2869);
nand U10540 (N_10540,N_1236,N_4815);
or U10541 (N_10541,N_477,N_3917);
nand U10542 (N_10542,N_2714,N_5776);
nand U10543 (N_10543,N_5602,N_2264);
nand U10544 (N_10544,N_4868,N_2763);
xor U10545 (N_10545,N_5321,N_4627);
xor U10546 (N_10546,N_2360,N_43);
nor U10547 (N_10547,N_1976,N_5793);
nor U10548 (N_10548,N_808,N_1871);
nor U10549 (N_10549,N_2475,N_4077);
xor U10550 (N_10550,N_205,N_2022);
nand U10551 (N_10551,N_5,N_3843);
nand U10552 (N_10552,N_5973,N_4750);
or U10553 (N_10553,N_3166,N_5662);
nor U10554 (N_10554,N_1851,N_665);
and U10555 (N_10555,N_522,N_1625);
xnor U10556 (N_10556,N_3432,N_4584);
nor U10557 (N_10557,N_3484,N_3080);
and U10558 (N_10558,N_3171,N_3020);
or U10559 (N_10559,N_4661,N_1420);
and U10560 (N_10560,N_4954,N_1030);
or U10561 (N_10561,N_3854,N_3423);
nand U10562 (N_10562,N_2940,N_650);
nor U10563 (N_10563,N_4861,N_2630);
nor U10564 (N_10564,N_3737,N_184);
xnor U10565 (N_10565,N_444,N_2227);
nor U10566 (N_10566,N_5211,N_2758);
and U10567 (N_10567,N_4969,N_1118);
xnor U10568 (N_10568,N_880,N_1059);
nor U10569 (N_10569,N_3897,N_3358);
nor U10570 (N_10570,N_5854,N_1318);
and U10571 (N_10571,N_5602,N_1577);
xnor U10572 (N_10572,N_3137,N_1221);
and U10573 (N_10573,N_422,N_4354);
nand U10574 (N_10574,N_956,N_1963);
nor U10575 (N_10575,N_229,N_2288);
nand U10576 (N_10576,N_1608,N_3249);
nor U10577 (N_10577,N_5505,N_760);
xor U10578 (N_10578,N_4204,N_4956);
nand U10579 (N_10579,N_3147,N_910);
xor U10580 (N_10580,N_5148,N_4677);
and U10581 (N_10581,N_4014,N_5899);
xor U10582 (N_10582,N_1732,N_5634);
xor U10583 (N_10583,N_5032,N_1261);
or U10584 (N_10584,N_1868,N_4627);
or U10585 (N_10585,N_4659,N_2614);
nor U10586 (N_10586,N_4928,N_5133);
or U10587 (N_10587,N_3674,N_3527);
xor U10588 (N_10588,N_2373,N_2376);
xnor U10589 (N_10589,N_1465,N_5077);
nor U10590 (N_10590,N_4311,N_4437);
or U10591 (N_10591,N_5665,N_5518);
or U10592 (N_10592,N_1911,N_3508);
xnor U10593 (N_10593,N_2010,N_5573);
xor U10594 (N_10594,N_5521,N_5631);
nor U10595 (N_10595,N_2414,N_2869);
and U10596 (N_10596,N_3638,N_729);
or U10597 (N_10597,N_3451,N_1373);
nor U10598 (N_10598,N_5120,N_2358);
and U10599 (N_10599,N_5740,N_5878);
and U10600 (N_10600,N_950,N_2538);
nand U10601 (N_10601,N_2050,N_3104);
nor U10602 (N_10602,N_5170,N_4461);
nand U10603 (N_10603,N_1756,N_1259);
or U10604 (N_10604,N_2279,N_394);
nor U10605 (N_10605,N_5912,N_222);
or U10606 (N_10606,N_856,N_276);
or U10607 (N_10607,N_4772,N_4811);
nand U10608 (N_10608,N_2010,N_1795);
nand U10609 (N_10609,N_4882,N_1360);
nor U10610 (N_10610,N_2201,N_848);
nand U10611 (N_10611,N_4174,N_405);
xor U10612 (N_10612,N_1066,N_773);
or U10613 (N_10613,N_5190,N_4474);
nor U10614 (N_10614,N_1448,N_411);
and U10615 (N_10615,N_4860,N_2232);
nand U10616 (N_10616,N_2439,N_4140);
nand U10617 (N_10617,N_1655,N_875);
xnor U10618 (N_10618,N_1765,N_123);
nand U10619 (N_10619,N_200,N_5751);
nand U10620 (N_10620,N_5,N_842);
and U10621 (N_10621,N_4705,N_4861);
or U10622 (N_10622,N_3955,N_1543);
or U10623 (N_10623,N_3588,N_5325);
xor U10624 (N_10624,N_1888,N_1132);
nand U10625 (N_10625,N_3681,N_2119);
and U10626 (N_10626,N_3908,N_2586);
and U10627 (N_10627,N_3521,N_5231);
or U10628 (N_10628,N_1946,N_5205);
and U10629 (N_10629,N_356,N_3804);
nand U10630 (N_10630,N_4035,N_1608);
xor U10631 (N_10631,N_5046,N_414);
xnor U10632 (N_10632,N_1217,N_5553);
xor U10633 (N_10633,N_3560,N_2110);
and U10634 (N_10634,N_5606,N_3785);
nor U10635 (N_10635,N_16,N_4576);
and U10636 (N_10636,N_2193,N_2315);
or U10637 (N_10637,N_153,N_2346);
and U10638 (N_10638,N_2188,N_819);
xnor U10639 (N_10639,N_5357,N_686);
or U10640 (N_10640,N_4839,N_2634);
nor U10641 (N_10641,N_2912,N_1882);
or U10642 (N_10642,N_4249,N_281);
nand U10643 (N_10643,N_1293,N_751);
nand U10644 (N_10644,N_1652,N_722);
and U10645 (N_10645,N_5371,N_5547);
nor U10646 (N_10646,N_1233,N_3046);
nand U10647 (N_10647,N_2592,N_5618);
or U10648 (N_10648,N_626,N_5073);
nor U10649 (N_10649,N_4457,N_3425);
nor U10650 (N_10650,N_1571,N_1803);
nor U10651 (N_10651,N_5209,N_1871);
and U10652 (N_10652,N_5554,N_1580);
nand U10653 (N_10653,N_4370,N_5434);
xnor U10654 (N_10654,N_133,N_1645);
xor U10655 (N_10655,N_4995,N_991);
and U10656 (N_10656,N_2322,N_5682);
nand U10657 (N_10657,N_2301,N_2256);
nor U10658 (N_10658,N_595,N_672);
nor U10659 (N_10659,N_2949,N_5173);
nand U10660 (N_10660,N_5317,N_1340);
or U10661 (N_10661,N_2409,N_1123);
xnor U10662 (N_10662,N_5111,N_3768);
nand U10663 (N_10663,N_1830,N_1226);
and U10664 (N_10664,N_1494,N_481);
nand U10665 (N_10665,N_5720,N_5198);
nor U10666 (N_10666,N_1029,N_849);
or U10667 (N_10667,N_5761,N_5178);
or U10668 (N_10668,N_199,N_3796);
nor U10669 (N_10669,N_5433,N_5477);
and U10670 (N_10670,N_5498,N_3224);
nand U10671 (N_10671,N_1111,N_5653);
and U10672 (N_10672,N_5460,N_1036);
or U10673 (N_10673,N_1928,N_1438);
or U10674 (N_10674,N_247,N_4258);
xor U10675 (N_10675,N_175,N_260);
or U10676 (N_10676,N_3270,N_1194);
xnor U10677 (N_10677,N_1012,N_3427);
nor U10678 (N_10678,N_159,N_2947);
or U10679 (N_10679,N_5861,N_3750);
nand U10680 (N_10680,N_2052,N_652);
and U10681 (N_10681,N_4152,N_4338);
and U10682 (N_10682,N_1340,N_3351);
nand U10683 (N_10683,N_3230,N_3524);
and U10684 (N_10684,N_705,N_2169);
xor U10685 (N_10685,N_4265,N_5819);
or U10686 (N_10686,N_719,N_5749);
or U10687 (N_10687,N_4662,N_4517);
xnor U10688 (N_10688,N_2462,N_3732);
xnor U10689 (N_10689,N_795,N_888);
xnor U10690 (N_10690,N_4307,N_5760);
or U10691 (N_10691,N_268,N_5950);
nand U10692 (N_10692,N_5715,N_1143);
nor U10693 (N_10693,N_1730,N_2976);
and U10694 (N_10694,N_5020,N_1341);
xnor U10695 (N_10695,N_5236,N_4044);
nand U10696 (N_10696,N_3410,N_5646);
xor U10697 (N_10697,N_273,N_4343);
xor U10698 (N_10698,N_1819,N_1180);
xor U10699 (N_10699,N_939,N_1897);
and U10700 (N_10700,N_3784,N_2434);
xor U10701 (N_10701,N_4711,N_3361);
or U10702 (N_10702,N_1202,N_3569);
and U10703 (N_10703,N_1805,N_5603);
and U10704 (N_10704,N_625,N_4894);
xor U10705 (N_10705,N_3475,N_2402);
xnor U10706 (N_10706,N_1669,N_3676);
nor U10707 (N_10707,N_3933,N_2197);
and U10708 (N_10708,N_3296,N_2317);
nand U10709 (N_10709,N_4748,N_288);
or U10710 (N_10710,N_235,N_1265);
xor U10711 (N_10711,N_208,N_1221);
xnor U10712 (N_10712,N_3753,N_3122);
and U10713 (N_10713,N_2717,N_5880);
or U10714 (N_10714,N_5746,N_3260);
xor U10715 (N_10715,N_3149,N_5765);
xor U10716 (N_10716,N_275,N_2639);
or U10717 (N_10717,N_4811,N_3559);
or U10718 (N_10718,N_5915,N_2239);
and U10719 (N_10719,N_4973,N_544);
xor U10720 (N_10720,N_1216,N_59);
xnor U10721 (N_10721,N_3016,N_4803);
xor U10722 (N_10722,N_2595,N_5535);
or U10723 (N_10723,N_3491,N_1776);
nand U10724 (N_10724,N_2957,N_1353);
nor U10725 (N_10725,N_822,N_1716);
and U10726 (N_10726,N_1052,N_1859);
nor U10727 (N_10727,N_3838,N_1478);
and U10728 (N_10728,N_3334,N_4563);
nor U10729 (N_10729,N_3613,N_730);
nand U10730 (N_10730,N_1742,N_4318);
or U10731 (N_10731,N_5054,N_1885);
xor U10732 (N_10732,N_2966,N_2414);
xnor U10733 (N_10733,N_97,N_3217);
nor U10734 (N_10734,N_570,N_3015);
or U10735 (N_10735,N_3714,N_4758);
nand U10736 (N_10736,N_4450,N_2952);
or U10737 (N_10737,N_4486,N_4872);
nand U10738 (N_10738,N_3331,N_1641);
xnor U10739 (N_10739,N_2152,N_4227);
xor U10740 (N_10740,N_2123,N_485);
nor U10741 (N_10741,N_3172,N_2516);
nand U10742 (N_10742,N_2868,N_5737);
or U10743 (N_10743,N_818,N_1286);
nand U10744 (N_10744,N_1688,N_5735);
and U10745 (N_10745,N_2061,N_950);
nand U10746 (N_10746,N_2874,N_2587);
xnor U10747 (N_10747,N_4646,N_514);
xor U10748 (N_10748,N_5470,N_5044);
nand U10749 (N_10749,N_3213,N_769);
nor U10750 (N_10750,N_997,N_2466);
nand U10751 (N_10751,N_269,N_884);
and U10752 (N_10752,N_4297,N_3379);
xnor U10753 (N_10753,N_345,N_5146);
nor U10754 (N_10754,N_1592,N_1555);
and U10755 (N_10755,N_5567,N_5444);
xor U10756 (N_10756,N_1786,N_5966);
xnor U10757 (N_10757,N_1396,N_3391);
nand U10758 (N_10758,N_761,N_3909);
or U10759 (N_10759,N_241,N_2027);
or U10760 (N_10760,N_1897,N_1465);
nor U10761 (N_10761,N_1088,N_5340);
xnor U10762 (N_10762,N_4787,N_2044);
nor U10763 (N_10763,N_2987,N_870);
xor U10764 (N_10764,N_3412,N_4652);
xnor U10765 (N_10765,N_385,N_4758);
and U10766 (N_10766,N_1017,N_1057);
xor U10767 (N_10767,N_1031,N_2712);
xor U10768 (N_10768,N_2787,N_2773);
nor U10769 (N_10769,N_5296,N_3613);
and U10770 (N_10770,N_449,N_3874);
and U10771 (N_10771,N_1537,N_3831);
nor U10772 (N_10772,N_2441,N_3462);
xnor U10773 (N_10773,N_1058,N_1938);
or U10774 (N_10774,N_970,N_2373);
nand U10775 (N_10775,N_4457,N_1530);
nor U10776 (N_10776,N_364,N_222);
xor U10777 (N_10777,N_2964,N_4189);
nand U10778 (N_10778,N_622,N_1664);
nor U10779 (N_10779,N_3533,N_1304);
nand U10780 (N_10780,N_5210,N_4196);
and U10781 (N_10781,N_1853,N_3373);
xor U10782 (N_10782,N_1057,N_1487);
nand U10783 (N_10783,N_3585,N_2483);
and U10784 (N_10784,N_4071,N_4548);
xnor U10785 (N_10785,N_4470,N_1236);
and U10786 (N_10786,N_4887,N_2698);
and U10787 (N_10787,N_2184,N_5376);
xnor U10788 (N_10788,N_3233,N_2453);
nor U10789 (N_10789,N_5505,N_2621);
nor U10790 (N_10790,N_5334,N_1329);
or U10791 (N_10791,N_3123,N_3184);
nor U10792 (N_10792,N_4274,N_126);
nand U10793 (N_10793,N_5678,N_864);
nor U10794 (N_10794,N_3922,N_4950);
nor U10795 (N_10795,N_1421,N_2070);
and U10796 (N_10796,N_5001,N_5353);
and U10797 (N_10797,N_2932,N_4983);
and U10798 (N_10798,N_1526,N_434);
xnor U10799 (N_10799,N_4576,N_2887);
or U10800 (N_10800,N_1722,N_5595);
nor U10801 (N_10801,N_211,N_4483);
xnor U10802 (N_10802,N_4883,N_708);
and U10803 (N_10803,N_4285,N_3035);
or U10804 (N_10804,N_4595,N_3898);
or U10805 (N_10805,N_4345,N_3800);
and U10806 (N_10806,N_3368,N_3035);
and U10807 (N_10807,N_5066,N_4713);
xor U10808 (N_10808,N_5157,N_3412);
and U10809 (N_10809,N_570,N_1788);
nand U10810 (N_10810,N_3285,N_2898);
nand U10811 (N_10811,N_4733,N_2101);
and U10812 (N_10812,N_2886,N_3388);
nand U10813 (N_10813,N_1405,N_1731);
nor U10814 (N_10814,N_3137,N_5209);
nand U10815 (N_10815,N_1968,N_154);
nor U10816 (N_10816,N_3853,N_766);
nand U10817 (N_10817,N_2898,N_544);
or U10818 (N_10818,N_5823,N_3217);
nor U10819 (N_10819,N_1560,N_5481);
xor U10820 (N_10820,N_1298,N_2511);
and U10821 (N_10821,N_3290,N_1176);
xor U10822 (N_10822,N_2996,N_2484);
nor U10823 (N_10823,N_1124,N_1557);
xnor U10824 (N_10824,N_921,N_4637);
and U10825 (N_10825,N_5504,N_316);
or U10826 (N_10826,N_2607,N_3672);
xnor U10827 (N_10827,N_1670,N_1534);
nor U10828 (N_10828,N_3670,N_4971);
nand U10829 (N_10829,N_4184,N_3624);
xor U10830 (N_10830,N_1864,N_3759);
or U10831 (N_10831,N_4306,N_4906);
nand U10832 (N_10832,N_1395,N_1291);
and U10833 (N_10833,N_690,N_5470);
nor U10834 (N_10834,N_1454,N_693);
nand U10835 (N_10835,N_2281,N_2564);
xnor U10836 (N_10836,N_283,N_656);
nor U10837 (N_10837,N_5051,N_987);
and U10838 (N_10838,N_4420,N_4224);
xor U10839 (N_10839,N_5592,N_2046);
or U10840 (N_10840,N_105,N_1390);
xor U10841 (N_10841,N_4739,N_72);
or U10842 (N_10842,N_1458,N_3070);
xnor U10843 (N_10843,N_4801,N_4455);
nor U10844 (N_10844,N_4315,N_4256);
nor U10845 (N_10845,N_5495,N_168);
xor U10846 (N_10846,N_1967,N_5987);
and U10847 (N_10847,N_5806,N_3683);
or U10848 (N_10848,N_3964,N_960);
xor U10849 (N_10849,N_3183,N_4395);
nand U10850 (N_10850,N_814,N_5117);
and U10851 (N_10851,N_2850,N_1214);
nand U10852 (N_10852,N_3206,N_1585);
and U10853 (N_10853,N_115,N_3878);
or U10854 (N_10854,N_108,N_4105);
xor U10855 (N_10855,N_2107,N_1915);
or U10856 (N_10856,N_2431,N_2201);
and U10857 (N_10857,N_3225,N_5976);
or U10858 (N_10858,N_4734,N_4357);
or U10859 (N_10859,N_5583,N_3879);
xnor U10860 (N_10860,N_3427,N_3977);
xnor U10861 (N_10861,N_4958,N_3347);
nor U10862 (N_10862,N_1261,N_5340);
xnor U10863 (N_10863,N_1738,N_5193);
nand U10864 (N_10864,N_5780,N_5421);
nor U10865 (N_10865,N_4280,N_1938);
xnor U10866 (N_10866,N_4661,N_3376);
nand U10867 (N_10867,N_531,N_1864);
and U10868 (N_10868,N_2606,N_1686);
and U10869 (N_10869,N_2471,N_2594);
or U10870 (N_10870,N_2143,N_2256);
nor U10871 (N_10871,N_2015,N_4396);
nor U10872 (N_10872,N_2492,N_3204);
nand U10873 (N_10873,N_3690,N_2270);
and U10874 (N_10874,N_355,N_5160);
nand U10875 (N_10875,N_1885,N_1528);
nand U10876 (N_10876,N_1026,N_4527);
or U10877 (N_10877,N_3707,N_4360);
nand U10878 (N_10878,N_3226,N_4321);
and U10879 (N_10879,N_5999,N_3440);
and U10880 (N_10880,N_5348,N_3776);
nand U10881 (N_10881,N_5068,N_5060);
nand U10882 (N_10882,N_3697,N_1896);
or U10883 (N_10883,N_4256,N_2187);
nor U10884 (N_10884,N_1652,N_464);
nor U10885 (N_10885,N_1617,N_4094);
xor U10886 (N_10886,N_3111,N_612);
xnor U10887 (N_10887,N_1199,N_2352);
and U10888 (N_10888,N_3149,N_3373);
xor U10889 (N_10889,N_3361,N_5359);
nand U10890 (N_10890,N_3535,N_3891);
or U10891 (N_10891,N_900,N_1142);
or U10892 (N_10892,N_5084,N_3641);
xnor U10893 (N_10893,N_2785,N_5056);
xnor U10894 (N_10894,N_619,N_1801);
xnor U10895 (N_10895,N_2885,N_4850);
xor U10896 (N_10896,N_666,N_3681);
and U10897 (N_10897,N_4371,N_939);
and U10898 (N_10898,N_3618,N_5674);
or U10899 (N_10899,N_1270,N_1136);
nand U10900 (N_10900,N_1722,N_4249);
or U10901 (N_10901,N_3189,N_2519);
xnor U10902 (N_10902,N_5759,N_3827);
nand U10903 (N_10903,N_5547,N_5083);
nand U10904 (N_10904,N_1520,N_3960);
nand U10905 (N_10905,N_4794,N_4155);
or U10906 (N_10906,N_2210,N_3691);
nor U10907 (N_10907,N_5078,N_5312);
or U10908 (N_10908,N_3805,N_2479);
and U10909 (N_10909,N_4410,N_5199);
xnor U10910 (N_10910,N_4897,N_5585);
or U10911 (N_10911,N_4787,N_1117);
xnor U10912 (N_10912,N_2511,N_3357);
and U10913 (N_10913,N_138,N_3693);
or U10914 (N_10914,N_1883,N_4755);
nor U10915 (N_10915,N_4527,N_1450);
nand U10916 (N_10916,N_1564,N_948);
and U10917 (N_10917,N_552,N_3917);
xnor U10918 (N_10918,N_4482,N_2473);
or U10919 (N_10919,N_5117,N_3428);
nand U10920 (N_10920,N_1551,N_1014);
or U10921 (N_10921,N_4848,N_613);
or U10922 (N_10922,N_1881,N_3102);
nor U10923 (N_10923,N_85,N_5328);
xnor U10924 (N_10924,N_2254,N_2040);
nand U10925 (N_10925,N_1978,N_795);
nor U10926 (N_10926,N_2883,N_4943);
and U10927 (N_10927,N_2802,N_1988);
nand U10928 (N_10928,N_4376,N_3953);
nor U10929 (N_10929,N_2492,N_3033);
or U10930 (N_10930,N_3040,N_5301);
and U10931 (N_10931,N_611,N_2899);
or U10932 (N_10932,N_3997,N_3417);
xnor U10933 (N_10933,N_5193,N_4841);
and U10934 (N_10934,N_1717,N_5962);
and U10935 (N_10935,N_1879,N_646);
and U10936 (N_10936,N_1890,N_637);
or U10937 (N_10937,N_1312,N_5376);
nand U10938 (N_10938,N_3065,N_5122);
nand U10939 (N_10939,N_4083,N_1133);
or U10940 (N_10940,N_2932,N_2002);
nand U10941 (N_10941,N_3402,N_1654);
or U10942 (N_10942,N_1275,N_3924);
nor U10943 (N_10943,N_1451,N_4353);
xor U10944 (N_10944,N_4895,N_165);
and U10945 (N_10945,N_264,N_4992);
or U10946 (N_10946,N_4467,N_2111);
or U10947 (N_10947,N_4686,N_730);
or U10948 (N_10948,N_4851,N_5900);
or U10949 (N_10949,N_5335,N_1289);
and U10950 (N_10950,N_4116,N_851);
or U10951 (N_10951,N_3393,N_1728);
nand U10952 (N_10952,N_1944,N_2880);
and U10953 (N_10953,N_4792,N_2911);
nor U10954 (N_10954,N_3832,N_1179);
nor U10955 (N_10955,N_2362,N_840);
and U10956 (N_10956,N_4403,N_5311);
xor U10957 (N_10957,N_3668,N_2600);
and U10958 (N_10958,N_5866,N_2947);
and U10959 (N_10959,N_4432,N_4357);
or U10960 (N_10960,N_250,N_294);
nor U10961 (N_10961,N_3388,N_1480);
xor U10962 (N_10962,N_298,N_937);
nand U10963 (N_10963,N_722,N_4511);
and U10964 (N_10964,N_4779,N_5044);
nand U10965 (N_10965,N_400,N_4062);
nand U10966 (N_10966,N_3728,N_695);
nor U10967 (N_10967,N_2972,N_3790);
or U10968 (N_10968,N_3333,N_2885);
nor U10969 (N_10969,N_4760,N_4066);
nor U10970 (N_10970,N_2744,N_2209);
and U10971 (N_10971,N_4925,N_472);
or U10972 (N_10972,N_88,N_3514);
nor U10973 (N_10973,N_241,N_651);
nand U10974 (N_10974,N_2121,N_2539);
or U10975 (N_10975,N_5046,N_3983);
nand U10976 (N_10976,N_112,N_4259);
nor U10977 (N_10977,N_3783,N_5651);
or U10978 (N_10978,N_2043,N_1193);
xor U10979 (N_10979,N_1648,N_5091);
or U10980 (N_10980,N_5073,N_2398);
or U10981 (N_10981,N_1195,N_325);
nor U10982 (N_10982,N_566,N_4401);
nor U10983 (N_10983,N_5608,N_3278);
xor U10984 (N_10984,N_5965,N_746);
nor U10985 (N_10985,N_4816,N_3749);
nand U10986 (N_10986,N_2892,N_5671);
and U10987 (N_10987,N_3726,N_2471);
or U10988 (N_10988,N_4347,N_1572);
nor U10989 (N_10989,N_5546,N_5107);
nand U10990 (N_10990,N_2894,N_4914);
nor U10991 (N_10991,N_3064,N_2461);
nand U10992 (N_10992,N_3980,N_2992);
or U10993 (N_10993,N_1583,N_5774);
nand U10994 (N_10994,N_5283,N_559);
and U10995 (N_10995,N_3480,N_5099);
nand U10996 (N_10996,N_3280,N_3835);
or U10997 (N_10997,N_2973,N_531);
or U10998 (N_10998,N_1745,N_5423);
xor U10999 (N_10999,N_3873,N_5954);
nand U11000 (N_11000,N_3314,N_2317);
nor U11001 (N_11001,N_41,N_5835);
or U11002 (N_11002,N_5541,N_3104);
or U11003 (N_11003,N_3907,N_1420);
xor U11004 (N_11004,N_2077,N_5240);
nand U11005 (N_11005,N_5016,N_4463);
nor U11006 (N_11006,N_56,N_5233);
nand U11007 (N_11007,N_4438,N_197);
nand U11008 (N_11008,N_5276,N_528);
nand U11009 (N_11009,N_385,N_1274);
nor U11010 (N_11010,N_4729,N_1838);
nor U11011 (N_11011,N_5344,N_501);
nor U11012 (N_11012,N_4036,N_3964);
or U11013 (N_11013,N_148,N_174);
nand U11014 (N_11014,N_3154,N_2448);
and U11015 (N_11015,N_4355,N_181);
or U11016 (N_11016,N_1818,N_5109);
nor U11017 (N_11017,N_5760,N_4137);
and U11018 (N_11018,N_2613,N_4499);
nor U11019 (N_11019,N_2586,N_3098);
nor U11020 (N_11020,N_711,N_5963);
nor U11021 (N_11021,N_1541,N_3819);
or U11022 (N_11022,N_815,N_456);
xnor U11023 (N_11023,N_1102,N_2917);
and U11024 (N_11024,N_1682,N_1541);
xor U11025 (N_11025,N_1340,N_5640);
or U11026 (N_11026,N_1670,N_1704);
nor U11027 (N_11027,N_2443,N_3298);
nand U11028 (N_11028,N_2028,N_839);
nand U11029 (N_11029,N_3835,N_5638);
or U11030 (N_11030,N_301,N_4484);
and U11031 (N_11031,N_2488,N_3469);
or U11032 (N_11032,N_2886,N_1969);
nor U11033 (N_11033,N_949,N_152);
xnor U11034 (N_11034,N_4859,N_81);
xnor U11035 (N_11035,N_718,N_3441);
nand U11036 (N_11036,N_3991,N_2677);
xor U11037 (N_11037,N_2535,N_581);
xnor U11038 (N_11038,N_862,N_1277);
nand U11039 (N_11039,N_2691,N_1941);
nand U11040 (N_11040,N_2899,N_4677);
nand U11041 (N_11041,N_5374,N_3420);
nor U11042 (N_11042,N_2714,N_1278);
nor U11043 (N_11043,N_3111,N_3365);
xor U11044 (N_11044,N_4582,N_2208);
xor U11045 (N_11045,N_4716,N_4772);
or U11046 (N_11046,N_4448,N_3540);
nand U11047 (N_11047,N_3700,N_1823);
and U11048 (N_11048,N_2253,N_833);
or U11049 (N_11049,N_5170,N_5367);
nand U11050 (N_11050,N_4216,N_4318);
nand U11051 (N_11051,N_1759,N_5556);
nand U11052 (N_11052,N_4242,N_4881);
and U11053 (N_11053,N_966,N_668);
xor U11054 (N_11054,N_1539,N_3860);
and U11055 (N_11055,N_5687,N_4576);
nand U11056 (N_11056,N_1536,N_81);
nand U11057 (N_11057,N_1793,N_534);
or U11058 (N_11058,N_222,N_3700);
nand U11059 (N_11059,N_2359,N_1814);
or U11060 (N_11060,N_5951,N_863);
nor U11061 (N_11061,N_1025,N_2749);
nand U11062 (N_11062,N_4,N_3463);
nand U11063 (N_11063,N_1873,N_4988);
nand U11064 (N_11064,N_3604,N_5563);
or U11065 (N_11065,N_4016,N_3244);
and U11066 (N_11066,N_5029,N_3695);
and U11067 (N_11067,N_4097,N_829);
and U11068 (N_11068,N_1347,N_4454);
nor U11069 (N_11069,N_4152,N_1822);
nand U11070 (N_11070,N_497,N_1325);
and U11071 (N_11071,N_1818,N_4273);
and U11072 (N_11072,N_3806,N_4088);
nand U11073 (N_11073,N_1378,N_1181);
nor U11074 (N_11074,N_4313,N_688);
and U11075 (N_11075,N_3056,N_3071);
xor U11076 (N_11076,N_5133,N_2919);
nand U11077 (N_11077,N_2261,N_4514);
nor U11078 (N_11078,N_899,N_5582);
nand U11079 (N_11079,N_1179,N_5372);
nor U11080 (N_11080,N_2148,N_3415);
or U11081 (N_11081,N_4642,N_1230);
nor U11082 (N_11082,N_5003,N_923);
and U11083 (N_11083,N_1121,N_3945);
xnor U11084 (N_11084,N_4180,N_1);
nor U11085 (N_11085,N_4588,N_4374);
xnor U11086 (N_11086,N_3710,N_776);
and U11087 (N_11087,N_1595,N_3924);
or U11088 (N_11088,N_4780,N_2389);
nor U11089 (N_11089,N_5617,N_5631);
nor U11090 (N_11090,N_4061,N_5939);
and U11091 (N_11091,N_4338,N_2693);
and U11092 (N_11092,N_5048,N_4572);
nand U11093 (N_11093,N_5213,N_3383);
nor U11094 (N_11094,N_681,N_5954);
xnor U11095 (N_11095,N_4724,N_4928);
nor U11096 (N_11096,N_4776,N_5291);
nand U11097 (N_11097,N_2329,N_5449);
nand U11098 (N_11098,N_5252,N_3258);
nor U11099 (N_11099,N_1921,N_4179);
nand U11100 (N_11100,N_2431,N_5985);
and U11101 (N_11101,N_3271,N_128);
or U11102 (N_11102,N_4106,N_2186);
or U11103 (N_11103,N_1483,N_1042);
and U11104 (N_11104,N_4127,N_2871);
nor U11105 (N_11105,N_570,N_1902);
and U11106 (N_11106,N_4480,N_5190);
or U11107 (N_11107,N_3062,N_3315);
and U11108 (N_11108,N_3285,N_2313);
and U11109 (N_11109,N_5262,N_1479);
xor U11110 (N_11110,N_714,N_1255);
nor U11111 (N_11111,N_1348,N_3971);
xnor U11112 (N_11112,N_3949,N_5984);
or U11113 (N_11113,N_3931,N_5741);
or U11114 (N_11114,N_2895,N_5938);
xnor U11115 (N_11115,N_1347,N_344);
or U11116 (N_11116,N_2414,N_862);
nand U11117 (N_11117,N_5596,N_5212);
xnor U11118 (N_11118,N_3844,N_5733);
or U11119 (N_11119,N_3445,N_663);
nor U11120 (N_11120,N_4690,N_4121);
nand U11121 (N_11121,N_5029,N_2959);
nand U11122 (N_11122,N_2176,N_4671);
and U11123 (N_11123,N_861,N_1821);
xnor U11124 (N_11124,N_3638,N_5809);
nand U11125 (N_11125,N_5843,N_5374);
xnor U11126 (N_11126,N_5976,N_739);
and U11127 (N_11127,N_825,N_4399);
and U11128 (N_11128,N_3178,N_3709);
or U11129 (N_11129,N_1793,N_4911);
and U11130 (N_11130,N_3569,N_2960);
and U11131 (N_11131,N_2998,N_2869);
or U11132 (N_11132,N_5174,N_347);
xnor U11133 (N_11133,N_3836,N_4712);
and U11134 (N_11134,N_5331,N_5415);
or U11135 (N_11135,N_1596,N_5380);
xor U11136 (N_11136,N_449,N_941);
or U11137 (N_11137,N_359,N_2785);
xor U11138 (N_11138,N_5232,N_2155);
and U11139 (N_11139,N_82,N_2135);
nor U11140 (N_11140,N_321,N_5743);
or U11141 (N_11141,N_984,N_844);
xor U11142 (N_11142,N_325,N_4962);
xor U11143 (N_11143,N_2284,N_4082);
xor U11144 (N_11144,N_329,N_1062);
and U11145 (N_11145,N_2791,N_2841);
or U11146 (N_11146,N_5963,N_2295);
or U11147 (N_11147,N_4613,N_5170);
xor U11148 (N_11148,N_852,N_3733);
and U11149 (N_11149,N_1823,N_2915);
and U11150 (N_11150,N_4053,N_4118);
and U11151 (N_11151,N_1558,N_5096);
nor U11152 (N_11152,N_1736,N_3388);
or U11153 (N_11153,N_465,N_3313);
xnor U11154 (N_11154,N_924,N_485);
nor U11155 (N_11155,N_3864,N_5776);
and U11156 (N_11156,N_3130,N_5080);
xor U11157 (N_11157,N_2380,N_906);
nor U11158 (N_11158,N_1773,N_3523);
and U11159 (N_11159,N_117,N_5108);
nor U11160 (N_11160,N_1075,N_4855);
or U11161 (N_11161,N_1817,N_2075);
nor U11162 (N_11162,N_34,N_5553);
and U11163 (N_11163,N_1686,N_1021);
xor U11164 (N_11164,N_2195,N_3506);
and U11165 (N_11165,N_340,N_5628);
or U11166 (N_11166,N_1029,N_2707);
xor U11167 (N_11167,N_1773,N_2376);
nand U11168 (N_11168,N_2424,N_30);
nor U11169 (N_11169,N_2608,N_4720);
nor U11170 (N_11170,N_2279,N_2158);
and U11171 (N_11171,N_1336,N_4944);
or U11172 (N_11172,N_85,N_5861);
nor U11173 (N_11173,N_5343,N_1905);
nor U11174 (N_11174,N_1757,N_230);
nor U11175 (N_11175,N_3289,N_493);
nor U11176 (N_11176,N_4406,N_4323);
xnor U11177 (N_11177,N_3340,N_4471);
nand U11178 (N_11178,N_3643,N_2243);
or U11179 (N_11179,N_3261,N_2711);
nand U11180 (N_11180,N_5543,N_1707);
nor U11181 (N_11181,N_2594,N_3093);
xor U11182 (N_11182,N_4013,N_3100);
nand U11183 (N_11183,N_5212,N_2524);
xor U11184 (N_11184,N_4755,N_5949);
xnor U11185 (N_11185,N_2001,N_4338);
xor U11186 (N_11186,N_2401,N_3613);
and U11187 (N_11187,N_5306,N_705);
and U11188 (N_11188,N_1876,N_3492);
and U11189 (N_11189,N_1766,N_3020);
and U11190 (N_11190,N_2432,N_2067);
nand U11191 (N_11191,N_4186,N_1700);
xor U11192 (N_11192,N_314,N_453);
xnor U11193 (N_11193,N_418,N_2396);
xor U11194 (N_11194,N_672,N_3330);
nor U11195 (N_11195,N_3495,N_2874);
nor U11196 (N_11196,N_3315,N_3378);
and U11197 (N_11197,N_2145,N_4747);
nand U11198 (N_11198,N_3206,N_4959);
nor U11199 (N_11199,N_4630,N_5341);
nor U11200 (N_11200,N_2492,N_2177);
nand U11201 (N_11201,N_404,N_2205);
or U11202 (N_11202,N_3175,N_2421);
and U11203 (N_11203,N_5610,N_3757);
or U11204 (N_11204,N_1045,N_2517);
nor U11205 (N_11205,N_4588,N_1835);
nand U11206 (N_11206,N_1757,N_415);
nor U11207 (N_11207,N_4804,N_3675);
and U11208 (N_11208,N_3173,N_3523);
xor U11209 (N_11209,N_2582,N_5718);
nand U11210 (N_11210,N_2069,N_235);
and U11211 (N_11211,N_3158,N_5192);
nand U11212 (N_11212,N_5495,N_5468);
nand U11213 (N_11213,N_4428,N_2695);
nand U11214 (N_11214,N_5772,N_1825);
xor U11215 (N_11215,N_5047,N_664);
xnor U11216 (N_11216,N_2081,N_2788);
and U11217 (N_11217,N_4117,N_2206);
and U11218 (N_11218,N_1206,N_428);
nor U11219 (N_11219,N_1736,N_678);
and U11220 (N_11220,N_5017,N_4344);
and U11221 (N_11221,N_2291,N_2091);
and U11222 (N_11222,N_5696,N_2522);
nand U11223 (N_11223,N_4229,N_5711);
or U11224 (N_11224,N_5862,N_5517);
and U11225 (N_11225,N_120,N_4932);
nand U11226 (N_11226,N_1713,N_2392);
or U11227 (N_11227,N_390,N_4563);
nand U11228 (N_11228,N_245,N_559);
and U11229 (N_11229,N_4026,N_2581);
and U11230 (N_11230,N_2279,N_2331);
or U11231 (N_11231,N_3240,N_1110);
and U11232 (N_11232,N_1619,N_5119);
nor U11233 (N_11233,N_2929,N_4035);
nand U11234 (N_11234,N_5919,N_2674);
nor U11235 (N_11235,N_2789,N_344);
nand U11236 (N_11236,N_715,N_52);
nor U11237 (N_11237,N_1985,N_1912);
xor U11238 (N_11238,N_1058,N_5756);
xnor U11239 (N_11239,N_454,N_2539);
nor U11240 (N_11240,N_4940,N_2554);
and U11241 (N_11241,N_2326,N_4282);
or U11242 (N_11242,N_2946,N_1249);
or U11243 (N_11243,N_4698,N_3573);
nor U11244 (N_11244,N_2515,N_13);
or U11245 (N_11245,N_3874,N_2015);
xnor U11246 (N_11246,N_1474,N_355);
nor U11247 (N_11247,N_1498,N_5650);
or U11248 (N_11248,N_4507,N_1367);
nand U11249 (N_11249,N_5774,N_1589);
or U11250 (N_11250,N_1204,N_3910);
xor U11251 (N_11251,N_1763,N_3278);
xor U11252 (N_11252,N_2506,N_3041);
or U11253 (N_11253,N_2073,N_3401);
nand U11254 (N_11254,N_296,N_3900);
and U11255 (N_11255,N_172,N_5113);
or U11256 (N_11256,N_300,N_3869);
xor U11257 (N_11257,N_5252,N_2935);
nand U11258 (N_11258,N_5361,N_1383);
nor U11259 (N_11259,N_5634,N_693);
or U11260 (N_11260,N_4704,N_5899);
nand U11261 (N_11261,N_1666,N_753);
xor U11262 (N_11262,N_2364,N_4815);
nor U11263 (N_11263,N_391,N_4021);
nor U11264 (N_11264,N_5384,N_634);
xnor U11265 (N_11265,N_1456,N_2727);
nor U11266 (N_11266,N_3925,N_5370);
nor U11267 (N_11267,N_5305,N_4051);
or U11268 (N_11268,N_5554,N_4270);
nand U11269 (N_11269,N_876,N_5675);
xnor U11270 (N_11270,N_957,N_1218);
nor U11271 (N_11271,N_1669,N_4117);
xnor U11272 (N_11272,N_3550,N_708);
and U11273 (N_11273,N_3769,N_1331);
nor U11274 (N_11274,N_992,N_2992);
nor U11275 (N_11275,N_3907,N_5168);
nand U11276 (N_11276,N_4430,N_4141);
or U11277 (N_11277,N_3782,N_1746);
nor U11278 (N_11278,N_2180,N_1943);
xnor U11279 (N_11279,N_1497,N_5623);
xor U11280 (N_11280,N_1860,N_4790);
or U11281 (N_11281,N_5540,N_3652);
or U11282 (N_11282,N_1939,N_778);
or U11283 (N_11283,N_1758,N_603);
or U11284 (N_11284,N_888,N_4055);
and U11285 (N_11285,N_5790,N_2277);
and U11286 (N_11286,N_2703,N_5968);
and U11287 (N_11287,N_3158,N_5253);
xnor U11288 (N_11288,N_3975,N_232);
nand U11289 (N_11289,N_5769,N_1282);
nand U11290 (N_11290,N_4477,N_4273);
nor U11291 (N_11291,N_5311,N_4792);
and U11292 (N_11292,N_688,N_1606);
or U11293 (N_11293,N_3015,N_5131);
nand U11294 (N_11294,N_4729,N_2233);
and U11295 (N_11295,N_5191,N_1687);
or U11296 (N_11296,N_4875,N_925);
nand U11297 (N_11297,N_4722,N_262);
nor U11298 (N_11298,N_974,N_3785);
xor U11299 (N_11299,N_4832,N_392);
nor U11300 (N_11300,N_605,N_5127);
and U11301 (N_11301,N_5391,N_3270);
or U11302 (N_11302,N_4980,N_325);
or U11303 (N_11303,N_4467,N_5822);
xor U11304 (N_11304,N_3892,N_488);
or U11305 (N_11305,N_3109,N_2103);
xor U11306 (N_11306,N_2502,N_2602);
or U11307 (N_11307,N_1209,N_430);
nand U11308 (N_11308,N_209,N_851);
and U11309 (N_11309,N_181,N_1475);
and U11310 (N_11310,N_5963,N_1384);
nand U11311 (N_11311,N_2060,N_982);
nand U11312 (N_11312,N_5429,N_3978);
xnor U11313 (N_11313,N_4170,N_4813);
xnor U11314 (N_11314,N_3128,N_4061);
xor U11315 (N_11315,N_3183,N_3065);
or U11316 (N_11316,N_3068,N_2020);
xor U11317 (N_11317,N_5433,N_4895);
and U11318 (N_11318,N_2235,N_4451);
and U11319 (N_11319,N_159,N_5501);
xnor U11320 (N_11320,N_288,N_5803);
nand U11321 (N_11321,N_3334,N_1905);
and U11322 (N_11322,N_2282,N_3303);
xor U11323 (N_11323,N_2245,N_756);
or U11324 (N_11324,N_440,N_5093);
nor U11325 (N_11325,N_3884,N_4324);
nor U11326 (N_11326,N_4178,N_586);
and U11327 (N_11327,N_2002,N_5893);
nand U11328 (N_11328,N_2473,N_2169);
nor U11329 (N_11329,N_5236,N_2351);
or U11330 (N_11330,N_213,N_5373);
and U11331 (N_11331,N_2188,N_5706);
xnor U11332 (N_11332,N_5153,N_978);
nor U11333 (N_11333,N_4993,N_3519);
nor U11334 (N_11334,N_2963,N_5724);
xnor U11335 (N_11335,N_1852,N_3345);
and U11336 (N_11336,N_5757,N_2742);
nand U11337 (N_11337,N_2713,N_1333);
nor U11338 (N_11338,N_3887,N_4895);
nor U11339 (N_11339,N_735,N_2190);
and U11340 (N_11340,N_850,N_5591);
nand U11341 (N_11341,N_1781,N_963);
xnor U11342 (N_11342,N_4515,N_2908);
xnor U11343 (N_11343,N_5177,N_2817);
and U11344 (N_11344,N_2063,N_5847);
nand U11345 (N_11345,N_975,N_3211);
nor U11346 (N_11346,N_1517,N_380);
or U11347 (N_11347,N_2195,N_4595);
xnor U11348 (N_11348,N_5376,N_3446);
or U11349 (N_11349,N_1887,N_3483);
nor U11350 (N_11350,N_2063,N_1919);
nand U11351 (N_11351,N_1657,N_2491);
nand U11352 (N_11352,N_3924,N_5667);
nand U11353 (N_11353,N_35,N_3692);
xor U11354 (N_11354,N_3860,N_5658);
and U11355 (N_11355,N_662,N_1742);
and U11356 (N_11356,N_5078,N_5943);
and U11357 (N_11357,N_1785,N_7);
nor U11358 (N_11358,N_3311,N_3751);
nand U11359 (N_11359,N_3928,N_948);
nand U11360 (N_11360,N_760,N_3790);
xor U11361 (N_11361,N_3053,N_5973);
and U11362 (N_11362,N_2578,N_694);
nand U11363 (N_11363,N_10,N_1941);
nand U11364 (N_11364,N_3871,N_4549);
nor U11365 (N_11365,N_3624,N_2359);
and U11366 (N_11366,N_1665,N_500);
xor U11367 (N_11367,N_947,N_4368);
or U11368 (N_11368,N_2465,N_4014);
xnor U11369 (N_11369,N_1218,N_2507);
xor U11370 (N_11370,N_3682,N_3626);
xor U11371 (N_11371,N_2722,N_5986);
xnor U11372 (N_11372,N_5119,N_3783);
or U11373 (N_11373,N_5340,N_2559);
nand U11374 (N_11374,N_4506,N_5901);
nand U11375 (N_11375,N_3962,N_3800);
xnor U11376 (N_11376,N_3165,N_379);
nor U11377 (N_11377,N_3194,N_1211);
nand U11378 (N_11378,N_4271,N_5432);
and U11379 (N_11379,N_1478,N_915);
xnor U11380 (N_11380,N_639,N_5325);
or U11381 (N_11381,N_1916,N_1151);
nor U11382 (N_11382,N_4234,N_5772);
nand U11383 (N_11383,N_4531,N_5156);
xor U11384 (N_11384,N_5273,N_4559);
xor U11385 (N_11385,N_106,N_272);
and U11386 (N_11386,N_4701,N_1619);
nand U11387 (N_11387,N_1513,N_4274);
nor U11388 (N_11388,N_4446,N_3826);
nand U11389 (N_11389,N_3355,N_2763);
nor U11390 (N_11390,N_3129,N_2408);
or U11391 (N_11391,N_5253,N_3769);
xnor U11392 (N_11392,N_704,N_2895);
xor U11393 (N_11393,N_5178,N_2673);
nor U11394 (N_11394,N_1561,N_2028);
nor U11395 (N_11395,N_1220,N_5979);
and U11396 (N_11396,N_5866,N_1712);
or U11397 (N_11397,N_5554,N_5932);
nor U11398 (N_11398,N_1346,N_1640);
and U11399 (N_11399,N_5287,N_2889);
or U11400 (N_11400,N_3074,N_4628);
xnor U11401 (N_11401,N_1188,N_4112);
or U11402 (N_11402,N_2282,N_4158);
and U11403 (N_11403,N_5600,N_1735);
xor U11404 (N_11404,N_139,N_1905);
nor U11405 (N_11405,N_5591,N_3518);
or U11406 (N_11406,N_473,N_1772);
xor U11407 (N_11407,N_98,N_5072);
xnor U11408 (N_11408,N_5369,N_320);
or U11409 (N_11409,N_4577,N_4983);
and U11410 (N_11410,N_1694,N_2621);
nand U11411 (N_11411,N_970,N_1199);
and U11412 (N_11412,N_3657,N_964);
and U11413 (N_11413,N_4274,N_5455);
xor U11414 (N_11414,N_1404,N_3302);
nand U11415 (N_11415,N_5429,N_4809);
or U11416 (N_11416,N_4904,N_2175);
xnor U11417 (N_11417,N_4909,N_5902);
xor U11418 (N_11418,N_3837,N_425);
nor U11419 (N_11419,N_587,N_3022);
nand U11420 (N_11420,N_3251,N_2259);
xor U11421 (N_11421,N_4868,N_3689);
nor U11422 (N_11422,N_2240,N_4408);
xor U11423 (N_11423,N_3314,N_5033);
nor U11424 (N_11424,N_5200,N_4046);
and U11425 (N_11425,N_3225,N_4432);
nand U11426 (N_11426,N_1675,N_5243);
nor U11427 (N_11427,N_5433,N_5681);
or U11428 (N_11428,N_1101,N_1134);
nor U11429 (N_11429,N_3138,N_2345);
and U11430 (N_11430,N_2153,N_5689);
nor U11431 (N_11431,N_2010,N_4790);
xnor U11432 (N_11432,N_5938,N_2714);
and U11433 (N_11433,N_4277,N_2842);
xor U11434 (N_11434,N_568,N_809);
and U11435 (N_11435,N_4478,N_5186);
nand U11436 (N_11436,N_1758,N_5386);
or U11437 (N_11437,N_3991,N_1654);
xor U11438 (N_11438,N_5804,N_5531);
and U11439 (N_11439,N_1357,N_3805);
nand U11440 (N_11440,N_961,N_5823);
nand U11441 (N_11441,N_1154,N_3329);
and U11442 (N_11442,N_4060,N_5033);
or U11443 (N_11443,N_1472,N_1515);
or U11444 (N_11444,N_3640,N_5125);
nand U11445 (N_11445,N_566,N_783);
nor U11446 (N_11446,N_3055,N_2434);
xnor U11447 (N_11447,N_4779,N_1784);
or U11448 (N_11448,N_3,N_5547);
nand U11449 (N_11449,N_5171,N_844);
or U11450 (N_11450,N_4425,N_5274);
xor U11451 (N_11451,N_5398,N_5782);
or U11452 (N_11452,N_1644,N_2232);
nand U11453 (N_11453,N_3071,N_21);
nor U11454 (N_11454,N_4265,N_1516);
xor U11455 (N_11455,N_2930,N_725);
and U11456 (N_11456,N_3529,N_3451);
xnor U11457 (N_11457,N_3851,N_1053);
xnor U11458 (N_11458,N_3937,N_4602);
nor U11459 (N_11459,N_4861,N_4996);
nor U11460 (N_11460,N_3859,N_3836);
nor U11461 (N_11461,N_3436,N_1497);
or U11462 (N_11462,N_5840,N_4851);
nor U11463 (N_11463,N_3551,N_2317);
nand U11464 (N_11464,N_5565,N_1325);
and U11465 (N_11465,N_4754,N_3425);
nor U11466 (N_11466,N_1802,N_553);
nand U11467 (N_11467,N_2806,N_5269);
nor U11468 (N_11468,N_4759,N_530);
nand U11469 (N_11469,N_3515,N_1869);
xor U11470 (N_11470,N_2957,N_2088);
nor U11471 (N_11471,N_4770,N_3225);
nand U11472 (N_11472,N_4486,N_13);
nand U11473 (N_11473,N_309,N_4122);
nor U11474 (N_11474,N_5301,N_147);
nand U11475 (N_11475,N_784,N_2970);
nor U11476 (N_11476,N_1965,N_3091);
nor U11477 (N_11477,N_4373,N_1910);
nand U11478 (N_11478,N_5598,N_3831);
xor U11479 (N_11479,N_2805,N_3493);
or U11480 (N_11480,N_3938,N_3365);
nor U11481 (N_11481,N_217,N_2283);
nor U11482 (N_11482,N_4690,N_448);
and U11483 (N_11483,N_2106,N_558);
nor U11484 (N_11484,N_1622,N_2597);
nor U11485 (N_11485,N_169,N_2669);
xor U11486 (N_11486,N_4406,N_1023);
or U11487 (N_11487,N_3080,N_2487);
xnor U11488 (N_11488,N_24,N_1518);
xnor U11489 (N_11489,N_4302,N_2605);
or U11490 (N_11490,N_3959,N_1393);
and U11491 (N_11491,N_3791,N_1540);
nor U11492 (N_11492,N_4778,N_1218);
nand U11493 (N_11493,N_5366,N_1452);
nor U11494 (N_11494,N_4979,N_3932);
nand U11495 (N_11495,N_1383,N_3263);
nand U11496 (N_11496,N_1502,N_5009);
xnor U11497 (N_11497,N_514,N_2633);
and U11498 (N_11498,N_5159,N_1280);
xnor U11499 (N_11499,N_2591,N_3809);
and U11500 (N_11500,N_28,N_2927);
and U11501 (N_11501,N_4978,N_5808);
nand U11502 (N_11502,N_1721,N_1246);
xor U11503 (N_11503,N_5327,N_5211);
or U11504 (N_11504,N_1615,N_5446);
xor U11505 (N_11505,N_3774,N_315);
xor U11506 (N_11506,N_5824,N_5961);
nand U11507 (N_11507,N_3117,N_3153);
or U11508 (N_11508,N_1544,N_4318);
or U11509 (N_11509,N_1705,N_2729);
nor U11510 (N_11510,N_4315,N_4548);
xnor U11511 (N_11511,N_178,N_1052);
xor U11512 (N_11512,N_1374,N_871);
and U11513 (N_11513,N_5304,N_1719);
nand U11514 (N_11514,N_3052,N_5551);
xnor U11515 (N_11515,N_2463,N_2502);
and U11516 (N_11516,N_705,N_1987);
nand U11517 (N_11517,N_2235,N_1845);
nand U11518 (N_11518,N_562,N_2311);
nand U11519 (N_11519,N_5499,N_2696);
nor U11520 (N_11520,N_2161,N_2030);
or U11521 (N_11521,N_5896,N_3846);
nand U11522 (N_11522,N_2241,N_2757);
nor U11523 (N_11523,N_5880,N_4329);
nand U11524 (N_11524,N_5287,N_1149);
nor U11525 (N_11525,N_5561,N_3171);
nand U11526 (N_11526,N_3497,N_2286);
and U11527 (N_11527,N_851,N_205);
nand U11528 (N_11528,N_3861,N_4011);
xnor U11529 (N_11529,N_819,N_1267);
and U11530 (N_11530,N_3012,N_4877);
and U11531 (N_11531,N_309,N_1981);
nor U11532 (N_11532,N_3234,N_3780);
and U11533 (N_11533,N_5647,N_5994);
and U11534 (N_11534,N_1602,N_4930);
nand U11535 (N_11535,N_602,N_1312);
and U11536 (N_11536,N_2081,N_834);
and U11537 (N_11537,N_4797,N_163);
nand U11538 (N_11538,N_1275,N_1166);
nand U11539 (N_11539,N_1776,N_3558);
nor U11540 (N_11540,N_5568,N_4065);
nor U11541 (N_11541,N_2638,N_1808);
nor U11542 (N_11542,N_5517,N_1245);
nand U11543 (N_11543,N_4921,N_5678);
and U11544 (N_11544,N_5234,N_619);
or U11545 (N_11545,N_2202,N_4102);
nor U11546 (N_11546,N_5113,N_1933);
xnor U11547 (N_11547,N_2449,N_4882);
or U11548 (N_11548,N_2199,N_2321);
nor U11549 (N_11549,N_5168,N_2701);
and U11550 (N_11550,N_4052,N_2482);
or U11551 (N_11551,N_4131,N_2834);
nor U11552 (N_11552,N_781,N_2495);
and U11553 (N_11553,N_5130,N_5111);
nor U11554 (N_11554,N_1882,N_213);
and U11555 (N_11555,N_5633,N_79);
xnor U11556 (N_11556,N_5808,N_2389);
and U11557 (N_11557,N_3710,N_2747);
xnor U11558 (N_11558,N_5571,N_1423);
nand U11559 (N_11559,N_3872,N_5800);
and U11560 (N_11560,N_4119,N_4205);
and U11561 (N_11561,N_999,N_1578);
nor U11562 (N_11562,N_3006,N_3037);
or U11563 (N_11563,N_1628,N_1436);
or U11564 (N_11564,N_4821,N_535);
and U11565 (N_11565,N_2255,N_3734);
nand U11566 (N_11566,N_5313,N_3886);
xnor U11567 (N_11567,N_1027,N_1802);
and U11568 (N_11568,N_5539,N_661);
xnor U11569 (N_11569,N_4037,N_4535);
xor U11570 (N_11570,N_2135,N_1556);
xor U11571 (N_11571,N_4356,N_4382);
nor U11572 (N_11572,N_3025,N_5647);
xor U11573 (N_11573,N_3620,N_2639);
xor U11574 (N_11574,N_1614,N_2621);
xnor U11575 (N_11575,N_117,N_565);
nand U11576 (N_11576,N_5303,N_2670);
xor U11577 (N_11577,N_1112,N_3282);
nand U11578 (N_11578,N_1042,N_2191);
nor U11579 (N_11579,N_3973,N_1507);
or U11580 (N_11580,N_4115,N_1637);
and U11581 (N_11581,N_5834,N_2458);
or U11582 (N_11582,N_5133,N_5137);
xor U11583 (N_11583,N_306,N_4307);
and U11584 (N_11584,N_5677,N_2573);
or U11585 (N_11585,N_2997,N_3794);
or U11586 (N_11586,N_5439,N_704);
xnor U11587 (N_11587,N_5211,N_2449);
and U11588 (N_11588,N_1997,N_702);
xnor U11589 (N_11589,N_3300,N_5998);
nand U11590 (N_11590,N_4928,N_342);
xnor U11591 (N_11591,N_739,N_5689);
nor U11592 (N_11592,N_5802,N_5141);
or U11593 (N_11593,N_3862,N_3232);
xnor U11594 (N_11594,N_3541,N_45);
xnor U11595 (N_11595,N_4567,N_1391);
and U11596 (N_11596,N_1993,N_3582);
or U11597 (N_11597,N_3059,N_4393);
nor U11598 (N_11598,N_5448,N_1737);
nand U11599 (N_11599,N_4610,N_5595);
nand U11600 (N_11600,N_2686,N_5508);
or U11601 (N_11601,N_5939,N_1516);
or U11602 (N_11602,N_4517,N_3800);
or U11603 (N_11603,N_2976,N_4612);
nor U11604 (N_11604,N_3531,N_5402);
nand U11605 (N_11605,N_4718,N_3248);
or U11606 (N_11606,N_2874,N_657);
xor U11607 (N_11607,N_315,N_5018);
xor U11608 (N_11608,N_447,N_1651);
or U11609 (N_11609,N_3224,N_5637);
xnor U11610 (N_11610,N_4585,N_5114);
nand U11611 (N_11611,N_3142,N_5094);
xor U11612 (N_11612,N_5720,N_637);
and U11613 (N_11613,N_4007,N_4734);
nor U11614 (N_11614,N_1447,N_2921);
xor U11615 (N_11615,N_1103,N_3211);
or U11616 (N_11616,N_4957,N_1600);
nor U11617 (N_11617,N_3743,N_1150);
nand U11618 (N_11618,N_3243,N_1770);
nand U11619 (N_11619,N_5843,N_3019);
or U11620 (N_11620,N_1048,N_236);
nor U11621 (N_11621,N_2791,N_851);
nand U11622 (N_11622,N_371,N_2898);
xnor U11623 (N_11623,N_3416,N_1919);
nand U11624 (N_11624,N_1317,N_233);
nor U11625 (N_11625,N_1,N_5756);
nand U11626 (N_11626,N_1795,N_1607);
nand U11627 (N_11627,N_1632,N_2963);
xnor U11628 (N_11628,N_3527,N_3995);
nand U11629 (N_11629,N_5378,N_1567);
and U11630 (N_11630,N_2697,N_231);
xnor U11631 (N_11631,N_540,N_645);
and U11632 (N_11632,N_5491,N_3334);
nand U11633 (N_11633,N_5750,N_5491);
nand U11634 (N_11634,N_4403,N_948);
nand U11635 (N_11635,N_1530,N_2839);
xnor U11636 (N_11636,N_1053,N_3912);
xnor U11637 (N_11637,N_3208,N_4884);
nor U11638 (N_11638,N_3890,N_1450);
or U11639 (N_11639,N_1108,N_3126);
nand U11640 (N_11640,N_3318,N_2851);
nand U11641 (N_11641,N_4047,N_4366);
and U11642 (N_11642,N_1296,N_5163);
or U11643 (N_11643,N_3342,N_1166);
or U11644 (N_11644,N_4024,N_5420);
nor U11645 (N_11645,N_4473,N_5841);
nor U11646 (N_11646,N_4493,N_388);
or U11647 (N_11647,N_5099,N_3227);
or U11648 (N_11648,N_3759,N_2150);
or U11649 (N_11649,N_4701,N_942);
xor U11650 (N_11650,N_1044,N_3995);
or U11651 (N_11651,N_3738,N_4950);
nand U11652 (N_11652,N_5838,N_4861);
and U11653 (N_11653,N_1557,N_4155);
and U11654 (N_11654,N_5587,N_160);
nand U11655 (N_11655,N_924,N_4738);
and U11656 (N_11656,N_1186,N_5461);
and U11657 (N_11657,N_3149,N_1146);
xnor U11658 (N_11658,N_2668,N_4178);
xnor U11659 (N_11659,N_1168,N_3859);
nand U11660 (N_11660,N_3748,N_5286);
nor U11661 (N_11661,N_3662,N_3374);
and U11662 (N_11662,N_2963,N_1877);
nand U11663 (N_11663,N_4880,N_1632);
and U11664 (N_11664,N_593,N_2000);
nand U11665 (N_11665,N_3829,N_1094);
nand U11666 (N_11666,N_4808,N_2962);
xnor U11667 (N_11667,N_5573,N_1200);
or U11668 (N_11668,N_48,N_1368);
or U11669 (N_11669,N_3746,N_5439);
nand U11670 (N_11670,N_3894,N_1891);
nor U11671 (N_11671,N_4724,N_1696);
xor U11672 (N_11672,N_3766,N_3459);
nand U11673 (N_11673,N_3492,N_1843);
or U11674 (N_11674,N_3785,N_3494);
nor U11675 (N_11675,N_5425,N_4994);
nand U11676 (N_11676,N_3025,N_5926);
and U11677 (N_11677,N_2045,N_2300);
xor U11678 (N_11678,N_313,N_3330);
or U11679 (N_11679,N_985,N_3915);
xor U11680 (N_11680,N_4615,N_1988);
or U11681 (N_11681,N_3897,N_1218);
or U11682 (N_11682,N_4927,N_1733);
nand U11683 (N_11683,N_3429,N_745);
xnor U11684 (N_11684,N_2928,N_2886);
or U11685 (N_11685,N_4736,N_4439);
nor U11686 (N_11686,N_2463,N_801);
xnor U11687 (N_11687,N_4027,N_5805);
nor U11688 (N_11688,N_5792,N_2678);
or U11689 (N_11689,N_3155,N_2072);
nand U11690 (N_11690,N_1219,N_4084);
nand U11691 (N_11691,N_4850,N_5840);
nor U11692 (N_11692,N_3196,N_4976);
nand U11693 (N_11693,N_1274,N_1049);
nor U11694 (N_11694,N_5816,N_5219);
and U11695 (N_11695,N_2698,N_4082);
xnor U11696 (N_11696,N_3922,N_4160);
and U11697 (N_11697,N_4742,N_202);
or U11698 (N_11698,N_3788,N_2058);
and U11699 (N_11699,N_5139,N_382);
xnor U11700 (N_11700,N_1873,N_2578);
nor U11701 (N_11701,N_1499,N_1013);
nand U11702 (N_11702,N_5194,N_368);
nor U11703 (N_11703,N_4448,N_5598);
nor U11704 (N_11704,N_4920,N_5726);
xor U11705 (N_11705,N_2507,N_2709);
xnor U11706 (N_11706,N_312,N_2652);
and U11707 (N_11707,N_2792,N_3304);
nor U11708 (N_11708,N_5470,N_2569);
xnor U11709 (N_11709,N_2068,N_419);
nand U11710 (N_11710,N_2164,N_546);
xnor U11711 (N_11711,N_3607,N_935);
nor U11712 (N_11712,N_474,N_4315);
or U11713 (N_11713,N_5044,N_625);
nor U11714 (N_11714,N_2237,N_305);
nor U11715 (N_11715,N_3804,N_461);
xnor U11716 (N_11716,N_5391,N_2268);
or U11717 (N_11717,N_5893,N_1201);
or U11718 (N_11718,N_2181,N_3889);
nand U11719 (N_11719,N_1851,N_4798);
nand U11720 (N_11720,N_1915,N_4783);
xor U11721 (N_11721,N_5560,N_343);
or U11722 (N_11722,N_1871,N_2177);
and U11723 (N_11723,N_78,N_3483);
or U11724 (N_11724,N_846,N_631);
and U11725 (N_11725,N_3901,N_2403);
nand U11726 (N_11726,N_2351,N_4770);
and U11727 (N_11727,N_5608,N_5203);
or U11728 (N_11728,N_5782,N_4544);
and U11729 (N_11729,N_4338,N_3191);
nand U11730 (N_11730,N_2007,N_1511);
nand U11731 (N_11731,N_2230,N_1093);
xor U11732 (N_11732,N_1591,N_2736);
or U11733 (N_11733,N_689,N_3264);
nor U11734 (N_11734,N_5482,N_1599);
nand U11735 (N_11735,N_5295,N_1446);
nor U11736 (N_11736,N_221,N_5689);
xnor U11737 (N_11737,N_4694,N_3414);
nor U11738 (N_11738,N_2820,N_428);
and U11739 (N_11739,N_137,N_3223);
or U11740 (N_11740,N_135,N_1444);
xor U11741 (N_11741,N_1354,N_4458);
or U11742 (N_11742,N_1342,N_4961);
nor U11743 (N_11743,N_56,N_2818);
nor U11744 (N_11744,N_2521,N_2532);
and U11745 (N_11745,N_4080,N_1281);
nand U11746 (N_11746,N_4521,N_2013);
and U11747 (N_11747,N_2331,N_1676);
nor U11748 (N_11748,N_2089,N_2502);
nand U11749 (N_11749,N_48,N_5113);
and U11750 (N_11750,N_5812,N_2501);
nor U11751 (N_11751,N_3203,N_680);
or U11752 (N_11752,N_2466,N_2268);
nor U11753 (N_11753,N_2039,N_4813);
and U11754 (N_11754,N_4696,N_937);
nor U11755 (N_11755,N_5076,N_5414);
and U11756 (N_11756,N_2482,N_1295);
and U11757 (N_11757,N_5561,N_5515);
or U11758 (N_11758,N_146,N_1970);
xor U11759 (N_11759,N_239,N_3325);
xnor U11760 (N_11760,N_3439,N_4537);
nand U11761 (N_11761,N_1763,N_115);
nor U11762 (N_11762,N_1151,N_5425);
xor U11763 (N_11763,N_5113,N_5575);
xor U11764 (N_11764,N_2158,N_2485);
nand U11765 (N_11765,N_1790,N_3745);
xnor U11766 (N_11766,N_20,N_5165);
and U11767 (N_11767,N_179,N_4627);
nor U11768 (N_11768,N_4545,N_130);
and U11769 (N_11769,N_688,N_407);
and U11770 (N_11770,N_5938,N_1050);
and U11771 (N_11771,N_3284,N_1925);
or U11772 (N_11772,N_2730,N_2502);
and U11773 (N_11773,N_3341,N_4253);
or U11774 (N_11774,N_355,N_4279);
or U11775 (N_11775,N_2572,N_1113);
xnor U11776 (N_11776,N_1015,N_20);
nand U11777 (N_11777,N_288,N_3050);
nand U11778 (N_11778,N_5008,N_4872);
nor U11779 (N_11779,N_3441,N_4403);
nand U11780 (N_11780,N_1672,N_4597);
nand U11781 (N_11781,N_1590,N_5226);
and U11782 (N_11782,N_2854,N_3152);
xor U11783 (N_11783,N_887,N_1548);
nand U11784 (N_11784,N_320,N_291);
nor U11785 (N_11785,N_3640,N_3948);
nor U11786 (N_11786,N_3979,N_1102);
nand U11787 (N_11787,N_3873,N_5265);
or U11788 (N_11788,N_3025,N_1172);
or U11789 (N_11789,N_3335,N_1385);
nand U11790 (N_11790,N_5377,N_3480);
xor U11791 (N_11791,N_1650,N_2853);
xor U11792 (N_11792,N_3879,N_4403);
and U11793 (N_11793,N_4460,N_4089);
nand U11794 (N_11794,N_1270,N_5642);
or U11795 (N_11795,N_1736,N_2603);
xnor U11796 (N_11796,N_1336,N_4752);
and U11797 (N_11797,N_4021,N_4638);
and U11798 (N_11798,N_1065,N_2217);
xnor U11799 (N_11799,N_234,N_5684);
nand U11800 (N_11800,N_559,N_4743);
and U11801 (N_11801,N_5432,N_1104);
xnor U11802 (N_11802,N_5087,N_181);
or U11803 (N_11803,N_4708,N_4832);
nor U11804 (N_11804,N_5446,N_438);
and U11805 (N_11805,N_4895,N_4493);
nand U11806 (N_11806,N_2135,N_399);
and U11807 (N_11807,N_2968,N_1286);
nand U11808 (N_11808,N_1012,N_5092);
xor U11809 (N_11809,N_4432,N_5525);
nor U11810 (N_11810,N_4471,N_4171);
and U11811 (N_11811,N_2909,N_5463);
nand U11812 (N_11812,N_737,N_5590);
or U11813 (N_11813,N_3350,N_5019);
nor U11814 (N_11814,N_4092,N_1122);
nand U11815 (N_11815,N_5644,N_2508);
xor U11816 (N_11816,N_987,N_3094);
and U11817 (N_11817,N_688,N_4339);
xor U11818 (N_11818,N_4024,N_3514);
nand U11819 (N_11819,N_2198,N_2870);
nand U11820 (N_11820,N_1481,N_5492);
nor U11821 (N_11821,N_2818,N_1125);
nor U11822 (N_11822,N_5704,N_2805);
or U11823 (N_11823,N_2633,N_2691);
and U11824 (N_11824,N_1724,N_1260);
or U11825 (N_11825,N_4178,N_5531);
and U11826 (N_11826,N_4766,N_651);
xor U11827 (N_11827,N_2797,N_4149);
nand U11828 (N_11828,N_4321,N_2247);
nor U11829 (N_11829,N_4805,N_3885);
xor U11830 (N_11830,N_715,N_4662);
nand U11831 (N_11831,N_5665,N_3053);
and U11832 (N_11832,N_2893,N_1215);
and U11833 (N_11833,N_2970,N_1259);
xor U11834 (N_11834,N_5165,N_4960);
nor U11835 (N_11835,N_3062,N_5714);
nand U11836 (N_11836,N_4470,N_4925);
xor U11837 (N_11837,N_3716,N_307);
nor U11838 (N_11838,N_2179,N_85);
nand U11839 (N_11839,N_399,N_4120);
and U11840 (N_11840,N_3286,N_5852);
xnor U11841 (N_11841,N_3387,N_5235);
nor U11842 (N_11842,N_1562,N_213);
nor U11843 (N_11843,N_5759,N_5757);
and U11844 (N_11844,N_1924,N_2649);
nand U11845 (N_11845,N_2565,N_1946);
nor U11846 (N_11846,N_3605,N_845);
and U11847 (N_11847,N_2754,N_2195);
and U11848 (N_11848,N_2675,N_3370);
xnor U11849 (N_11849,N_4910,N_3763);
nor U11850 (N_11850,N_5611,N_3372);
xor U11851 (N_11851,N_2090,N_2818);
and U11852 (N_11852,N_3020,N_1971);
xor U11853 (N_11853,N_589,N_764);
or U11854 (N_11854,N_2836,N_5422);
nand U11855 (N_11855,N_993,N_1463);
nand U11856 (N_11856,N_5986,N_1298);
nor U11857 (N_11857,N_4769,N_1445);
xnor U11858 (N_11858,N_2680,N_2371);
nand U11859 (N_11859,N_4456,N_312);
and U11860 (N_11860,N_4713,N_2322);
xnor U11861 (N_11861,N_2386,N_4375);
nor U11862 (N_11862,N_3271,N_3068);
xor U11863 (N_11863,N_1757,N_4704);
or U11864 (N_11864,N_1434,N_5629);
xor U11865 (N_11865,N_5647,N_3012);
and U11866 (N_11866,N_3641,N_453);
or U11867 (N_11867,N_5465,N_2256);
nor U11868 (N_11868,N_5411,N_1665);
nand U11869 (N_11869,N_346,N_3179);
xnor U11870 (N_11870,N_984,N_1977);
xnor U11871 (N_11871,N_2244,N_929);
xnor U11872 (N_11872,N_4073,N_1686);
nor U11873 (N_11873,N_989,N_1609);
nor U11874 (N_11874,N_87,N_3825);
xnor U11875 (N_11875,N_5109,N_2105);
and U11876 (N_11876,N_4453,N_3568);
nor U11877 (N_11877,N_1554,N_863);
xnor U11878 (N_11878,N_4183,N_3975);
xnor U11879 (N_11879,N_2332,N_4609);
or U11880 (N_11880,N_471,N_5871);
or U11881 (N_11881,N_3674,N_709);
and U11882 (N_11882,N_2815,N_3299);
or U11883 (N_11883,N_5550,N_622);
or U11884 (N_11884,N_435,N_3375);
or U11885 (N_11885,N_3083,N_1574);
nand U11886 (N_11886,N_756,N_609);
nor U11887 (N_11887,N_3369,N_2303);
xnor U11888 (N_11888,N_4908,N_1201);
nand U11889 (N_11889,N_11,N_5834);
and U11890 (N_11890,N_2115,N_3033);
xnor U11891 (N_11891,N_4656,N_784);
xor U11892 (N_11892,N_5029,N_213);
nand U11893 (N_11893,N_1115,N_5071);
or U11894 (N_11894,N_4364,N_5408);
xnor U11895 (N_11895,N_5779,N_4248);
or U11896 (N_11896,N_1159,N_3804);
nand U11897 (N_11897,N_1007,N_5265);
or U11898 (N_11898,N_1317,N_3663);
xor U11899 (N_11899,N_5977,N_1932);
xnor U11900 (N_11900,N_3861,N_1154);
nor U11901 (N_11901,N_5927,N_3252);
or U11902 (N_11902,N_1042,N_3854);
xor U11903 (N_11903,N_3467,N_4388);
or U11904 (N_11904,N_1747,N_5862);
xnor U11905 (N_11905,N_2607,N_4217);
and U11906 (N_11906,N_267,N_5438);
and U11907 (N_11907,N_5212,N_1163);
nand U11908 (N_11908,N_4508,N_4434);
xor U11909 (N_11909,N_842,N_2829);
nand U11910 (N_11910,N_3310,N_5169);
xor U11911 (N_11911,N_1932,N_5377);
and U11912 (N_11912,N_755,N_1563);
nor U11913 (N_11913,N_3466,N_1755);
nand U11914 (N_11914,N_1984,N_1894);
nor U11915 (N_11915,N_5490,N_714);
or U11916 (N_11916,N_1402,N_4861);
and U11917 (N_11917,N_750,N_4374);
or U11918 (N_11918,N_5974,N_2479);
nand U11919 (N_11919,N_1065,N_1821);
xor U11920 (N_11920,N_5056,N_1680);
xnor U11921 (N_11921,N_5596,N_3838);
and U11922 (N_11922,N_2183,N_3372);
or U11923 (N_11923,N_497,N_3345);
xor U11924 (N_11924,N_3258,N_2334);
nand U11925 (N_11925,N_128,N_4465);
nand U11926 (N_11926,N_3779,N_2750);
nand U11927 (N_11927,N_5577,N_3542);
nand U11928 (N_11928,N_967,N_3258);
nor U11929 (N_11929,N_1692,N_3471);
and U11930 (N_11930,N_201,N_3022);
nor U11931 (N_11931,N_514,N_20);
xnor U11932 (N_11932,N_1964,N_2876);
nor U11933 (N_11933,N_1752,N_2399);
nor U11934 (N_11934,N_2714,N_1173);
and U11935 (N_11935,N_925,N_5540);
xnor U11936 (N_11936,N_5811,N_2446);
or U11937 (N_11937,N_2469,N_3705);
xnor U11938 (N_11938,N_5237,N_2102);
and U11939 (N_11939,N_306,N_4488);
and U11940 (N_11940,N_3252,N_3432);
nand U11941 (N_11941,N_524,N_2542);
or U11942 (N_11942,N_3544,N_4060);
or U11943 (N_11943,N_2513,N_2748);
xor U11944 (N_11944,N_4909,N_2077);
nand U11945 (N_11945,N_1067,N_2943);
and U11946 (N_11946,N_4556,N_1866);
xnor U11947 (N_11947,N_2760,N_457);
nor U11948 (N_11948,N_193,N_540);
xnor U11949 (N_11949,N_1560,N_1891);
or U11950 (N_11950,N_5808,N_3866);
nand U11951 (N_11951,N_2287,N_3928);
and U11952 (N_11952,N_2599,N_5697);
nor U11953 (N_11953,N_4726,N_3087);
nor U11954 (N_11954,N_215,N_2382);
and U11955 (N_11955,N_127,N_4270);
and U11956 (N_11956,N_1043,N_2045);
or U11957 (N_11957,N_3196,N_4149);
nor U11958 (N_11958,N_3431,N_798);
xor U11959 (N_11959,N_118,N_3122);
or U11960 (N_11960,N_2522,N_5824);
and U11961 (N_11961,N_625,N_1483);
xnor U11962 (N_11962,N_4075,N_704);
or U11963 (N_11963,N_5302,N_5960);
nand U11964 (N_11964,N_1133,N_1609);
or U11965 (N_11965,N_4608,N_3068);
nor U11966 (N_11966,N_3872,N_4874);
nand U11967 (N_11967,N_4869,N_5409);
nor U11968 (N_11968,N_181,N_3152);
xor U11969 (N_11969,N_3195,N_5580);
and U11970 (N_11970,N_4725,N_345);
nand U11971 (N_11971,N_3074,N_3143);
or U11972 (N_11972,N_1890,N_4488);
nor U11973 (N_11973,N_3038,N_626);
xnor U11974 (N_11974,N_1985,N_2197);
nand U11975 (N_11975,N_5958,N_4015);
nor U11976 (N_11976,N_5205,N_5688);
nand U11977 (N_11977,N_5736,N_3856);
and U11978 (N_11978,N_3381,N_1986);
and U11979 (N_11979,N_284,N_2137);
or U11980 (N_11980,N_4315,N_3355);
and U11981 (N_11981,N_5531,N_5206);
xnor U11982 (N_11982,N_4679,N_4108);
or U11983 (N_11983,N_1092,N_5394);
nor U11984 (N_11984,N_5489,N_681);
nand U11985 (N_11985,N_1652,N_2020);
nand U11986 (N_11986,N_5139,N_2077);
and U11987 (N_11987,N_3926,N_1514);
nand U11988 (N_11988,N_5501,N_5339);
xnor U11989 (N_11989,N_2694,N_4497);
and U11990 (N_11990,N_2718,N_3149);
nand U11991 (N_11991,N_5394,N_4952);
xnor U11992 (N_11992,N_821,N_4794);
nand U11993 (N_11993,N_1406,N_1819);
nor U11994 (N_11994,N_3293,N_5505);
nor U11995 (N_11995,N_3502,N_111);
nor U11996 (N_11996,N_1100,N_2953);
nor U11997 (N_11997,N_4234,N_4570);
nand U11998 (N_11998,N_2540,N_4196);
and U11999 (N_11999,N_3020,N_2349);
nor U12000 (N_12000,N_9477,N_11516);
or U12001 (N_12001,N_7555,N_7013);
nor U12002 (N_12002,N_6207,N_9259);
nand U12003 (N_12003,N_6473,N_9541);
and U12004 (N_12004,N_11537,N_10895);
and U12005 (N_12005,N_7138,N_11740);
xor U12006 (N_12006,N_8673,N_9287);
or U12007 (N_12007,N_6464,N_8288);
xor U12008 (N_12008,N_7134,N_6851);
xnor U12009 (N_12009,N_9451,N_9819);
or U12010 (N_12010,N_9872,N_8156);
xor U12011 (N_12011,N_11329,N_6121);
xor U12012 (N_12012,N_9910,N_7588);
nand U12013 (N_12013,N_11906,N_7589);
or U12014 (N_12014,N_10432,N_6526);
nor U12015 (N_12015,N_11250,N_10325);
or U12016 (N_12016,N_10835,N_8666);
and U12017 (N_12017,N_9471,N_7225);
nand U12018 (N_12018,N_7707,N_10836);
nor U12019 (N_12019,N_7987,N_10048);
and U12020 (N_12020,N_9982,N_11052);
nor U12021 (N_12021,N_11571,N_6316);
and U12022 (N_12022,N_6096,N_11770);
nand U12023 (N_12023,N_11394,N_7105);
or U12024 (N_12024,N_8846,N_7903);
xnor U12025 (N_12025,N_9878,N_11878);
xnor U12026 (N_12026,N_6413,N_11092);
and U12027 (N_12027,N_7116,N_8902);
nor U12028 (N_12028,N_10877,N_8062);
and U12029 (N_12029,N_6354,N_11841);
or U12030 (N_12030,N_7294,N_8611);
nand U12031 (N_12031,N_6775,N_9296);
nand U12032 (N_12032,N_9509,N_10305);
nor U12033 (N_12033,N_7189,N_10685);
and U12034 (N_12034,N_11622,N_10857);
and U12035 (N_12035,N_9200,N_7535);
nand U12036 (N_12036,N_7177,N_10092);
or U12037 (N_12037,N_10374,N_8536);
nand U12038 (N_12038,N_11623,N_7875);
xnor U12039 (N_12039,N_11921,N_7212);
nand U12040 (N_12040,N_7241,N_11800);
xor U12041 (N_12041,N_8622,N_8686);
xnor U12042 (N_12042,N_9031,N_11214);
and U12043 (N_12043,N_9655,N_10255);
nor U12044 (N_12044,N_7191,N_6624);
and U12045 (N_12045,N_10172,N_6707);
or U12046 (N_12046,N_7208,N_7038);
xor U12047 (N_12047,N_11726,N_10645);
or U12048 (N_12048,N_7356,N_8096);
nor U12049 (N_12049,N_7991,N_9216);
xor U12050 (N_12050,N_10851,N_6152);
nand U12051 (N_12051,N_10587,N_7369);
nand U12052 (N_12052,N_11872,N_8829);
or U12053 (N_12053,N_9083,N_10021);
and U12054 (N_12054,N_11886,N_7259);
xor U12055 (N_12055,N_11003,N_7657);
and U12056 (N_12056,N_9968,N_6610);
xnor U12057 (N_12057,N_10639,N_11734);
nand U12058 (N_12058,N_6400,N_6367);
and U12059 (N_12059,N_7446,N_7056);
xor U12060 (N_12060,N_8135,N_9478);
xnor U12061 (N_12061,N_11318,N_8669);
and U12062 (N_12062,N_11897,N_9124);
xnor U12063 (N_12063,N_7395,N_7675);
nor U12064 (N_12064,N_10414,N_6757);
nor U12065 (N_12065,N_10691,N_6343);
and U12066 (N_12066,N_10964,N_9893);
or U12067 (N_12067,N_6195,N_7949);
nand U12068 (N_12068,N_9839,N_8940);
nand U12069 (N_12069,N_10119,N_9650);
nand U12070 (N_12070,N_7124,N_8596);
nor U12071 (N_12071,N_8993,N_11925);
xor U12072 (N_12072,N_11861,N_6669);
xnor U12073 (N_12073,N_8109,N_11371);
and U12074 (N_12074,N_9605,N_11065);
nor U12075 (N_12075,N_8687,N_6454);
xnor U12076 (N_12076,N_11446,N_11220);
or U12077 (N_12077,N_7080,N_10596);
and U12078 (N_12078,N_7227,N_7566);
nor U12079 (N_12079,N_8547,N_10553);
nand U12080 (N_12080,N_9534,N_10683);
xnor U12081 (N_12081,N_7711,N_11964);
nand U12082 (N_12082,N_8816,N_7130);
nor U12083 (N_12083,N_6412,N_11136);
nand U12084 (N_12084,N_10572,N_11422);
nor U12085 (N_12085,N_8986,N_6540);
or U12086 (N_12086,N_11833,N_7409);
nor U12087 (N_12087,N_10419,N_9028);
or U12088 (N_12088,N_10516,N_9074);
nor U12089 (N_12089,N_10404,N_6563);
and U12090 (N_12090,N_8269,N_7094);
xnor U12091 (N_12091,N_9535,N_6493);
and U12092 (N_12092,N_9504,N_9679);
nor U12093 (N_12093,N_9618,N_7978);
or U12094 (N_12094,N_7444,N_7417);
nand U12095 (N_12095,N_11236,N_9298);
and U12096 (N_12096,N_10850,N_8002);
nor U12097 (N_12097,N_10126,N_11188);
or U12098 (N_12098,N_6361,N_7643);
nand U12099 (N_12099,N_11752,N_10373);
nand U12100 (N_12100,N_11184,N_8644);
nand U12101 (N_12101,N_9578,N_7583);
or U12102 (N_12102,N_10881,N_8219);
or U12103 (N_12103,N_8994,N_8578);
and U12104 (N_12104,N_6293,N_9876);
or U12105 (N_12105,N_11807,N_9723);
or U12106 (N_12106,N_11570,N_10862);
or U12107 (N_12107,N_10847,N_10137);
nor U12108 (N_12108,N_10575,N_7497);
nand U12109 (N_12109,N_8082,N_9934);
and U12110 (N_12110,N_6709,N_6889);
or U12111 (N_12111,N_7916,N_6419);
xor U12112 (N_12112,N_6083,N_6007);
nand U12113 (N_12113,N_10193,N_6475);
nor U12114 (N_12114,N_9470,N_6070);
nand U12115 (N_12115,N_11439,N_7224);
or U12116 (N_12116,N_10214,N_11464);
xor U12117 (N_12117,N_10585,N_10403);
nor U12118 (N_12118,N_9719,N_6960);
nor U12119 (N_12119,N_11229,N_11776);
nor U12120 (N_12120,N_10701,N_8719);
nor U12121 (N_12121,N_6461,N_11292);
nor U12122 (N_12122,N_6603,N_6731);
or U12123 (N_12123,N_6375,N_10931);
and U12124 (N_12124,N_11745,N_9002);
xnor U12125 (N_12125,N_10460,N_8930);
xnor U12126 (N_12126,N_8475,N_11508);
nand U12127 (N_12127,N_6600,N_9737);
nand U12128 (N_12128,N_6448,N_11525);
nor U12129 (N_12129,N_9813,N_11685);
nand U12130 (N_12130,N_11661,N_7236);
xor U12131 (N_12131,N_7979,N_10535);
nand U12132 (N_12132,N_6398,N_7392);
nand U12133 (N_12133,N_6386,N_9962);
nor U12134 (N_12134,N_10574,N_9180);
nand U12135 (N_12135,N_10647,N_11451);
or U12136 (N_12136,N_10786,N_10943);
or U12137 (N_12137,N_11950,N_7967);
nand U12138 (N_12138,N_9887,N_9674);
xnor U12139 (N_12139,N_8005,N_10658);
and U12140 (N_12140,N_7065,N_11288);
nor U12141 (N_12141,N_11562,N_8814);
or U12142 (N_12142,N_8297,N_6873);
or U12143 (N_12143,N_6917,N_8922);
nor U12144 (N_12144,N_10693,N_11890);
and U12145 (N_12145,N_6767,N_11044);
and U12146 (N_12146,N_7343,N_10736);
or U12147 (N_12147,N_8663,N_10719);
or U12148 (N_12148,N_7524,N_6064);
or U12149 (N_12149,N_7419,N_9040);
or U12150 (N_12150,N_9621,N_11678);
xnor U12151 (N_12151,N_10762,N_6756);
xor U12152 (N_12152,N_10738,N_10858);
and U12153 (N_12153,N_8912,N_11199);
nand U12154 (N_12154,N_9167,N_10248);
nand U12155 (N_12155,N_9198,N_11594);
and U12156 (N_12156,N_11613,N_10774);
nand U12157 (N_12157,N_11021,N_9333);
nand U12158 (N_12158,N_8947,N_9967);
or U12159 (N_12159,N_8864,N_11204);
or U12160 (N_12160,N_6809,N_6685);
nor U12161 (N_12161,N_6269,N_7695);
xnor U12162 (N_12162,N_6481,N_7918);
and U12163 (N_12163,N_9165,N_11586);
xnor U12164 (N_12164,N_9126,N_10712);
xor U12165 (N_12165,N_11176,N_9145);
or U12166 (N_12166,N_6486,N_11390);
xor U12167 (N_12167,N_6380,N_6988);
nor U12168 (N_12168,N_11963,N_10488);
and U12169 (N_12169,N_9268,N_7968);
nor U12170 (N_12170,N_9408,N_11694);
nor U12171 (N_12171,N_6797,N_11163);
nor U12172 (N_12172,N_11829,N_9453);
and U12173 (N_12173,N_10152,N_7345);
and U12174 (N_12174,N_9808,N_9877);
nor U12175 (N_12175,N_10310,N_6492);
or U12176 (N_12176,N_8551,N_7686);
and U12177 (N_12177,N_11287,N_8268);
xor U12178 (N_12178,N_9340,N_6828);
xor U12179 (N_12179,N_9398,N_8018);
and U12180 (N_12180,N_10182,N_7393);
and U12181 (N_12181,N_8585,N_6717);
xnor U12182 (N_12182,N_7265,N_10165);
nand U12183 (N_12183,N_10930,N_11857);
or U12184 (N_12184,N_11108,N_9981);
nor U12185 (N_12185,N_7861,N_10016);
xor U12186 (N_12186,N_6758,N_11936);
nor U12187 (N_12187,N_10741,N_10948);
nor U12188 (N_12188,N_10003,N_10412);
nor U12189 (N_12189,N_8291,N_7107);
xor U12190 (N_12190,N_11299,N_6930);
and U12191 (N_12191,N_6935,N_9036);
nand U12192 (N_12192,N_7808,N_7192);
or U12193 (N_12193,N_7173,N_6311);
or U12194 (N_12194,N_8228,N_8813);
xor U12195 (N_12195,N_8679,N_8736);
xnor U12196 (N_12196,N_10849,N_6535);
or U12197 (N_12197,N_10203,N_8909);
and U12198 (N_12198,N_8099,N_8690);
nor U12199 (N_12199,N_6782,N_6665);
xor U12200 (N_12200,N_6019,N_6234);
nor U12201 (N_12201,N_11319,N_7893);
xor U12202 (N_12202,N_8318,N_9560);
or U12203 (N_12203,N_8981,N_11757);
nand U12204 (N_12204,N_8049,N_6940);
nand U12205 (N_12205,N_7155,N_7276);
and U12206 (N_12206,N_10700,N_6067);
nor U12207 (N_12207,N_10904,N_9190);
and U12208 (N_12208,N_9256,N_7304);
nand U12209 (N_12209,N_8404,N_11896);
or U12210 (N_12210,N_7036,N_10352);
xnor U12211 (N_12211,N_8988,N_8146);
nand U12212 (N_12212,N_10321,N_10630);
xnor U12213 (N_12213,N_11715,N_7472);
or U12214 (N_12214,N_9117,N_8371);
and U12215 (N_12215,N_7638,N_6625);
or U12216 (N_12216,N_10200,N_8285);
xnor U12217 (N_12217,N_11510,N_11768);
xor U12218 (N_12218,N_8901,N_7637);
nand U12219 (N_12219,N_7057,N_7059);
nand U12220 (N_12220,N_11893,N_7266);
nand U12221 (N_12221,N_6010,N_9899);
and U12222 (N_12222,N_11760,N_7884);
xor U12223 (N_12223,N_10327,N_8065);
nor U12224 (N_12224,N_7430,N_10989);
nor U12225 (N_12225,N_9115,N_6983);
nand U12226 (N_12226,N_7853,N_7015);
xor U12227 (N_12227,N_9798,N_8259);
nor U12228 (N_12228,N_11320,N_11102);
xor U12229 (N_12229,N_7088,N_11498);
nor U12230 (N_12230,N_6394,N_10199);
xnor U12231 (N_12231,N_10086,N_6221);
nand U12232 (N_12232,N_9607,N_11967);
nand U12233 (N_12233,N_6833,N_10994);
xor U12234 (N_12234,N_11290,N_10929);
or U12235 (N_12235,N_8327,N_6837);
or U12236 (N_12236,N_10898,N_6682);
and U12237 (N_12237,N_10186,N_8682);
nand U12238 (N_12238,N_8395,N_10684);
nor U12239 (N_12239,N_7466,N_8181);
and U12240 (N_12240,N_11459,N_10465);
nor U12241 (N_12241,N_11160,N_6456);
nand U12242 (N_12242,N_9995,N_8811);
or U12243 (N_12243,N_10246,N_11111);
xor U12244 (N_12244,N_9848,N_11333);
xnor U12245 (N_12245,N_9120,N_8387);
nor U12246 (N_12246,N_9303,N_11601);
nor U12247 (N_12247,N_8919,N_9410);
or U12248 (N_12248,N_11777,N_11995);
nand U12249 (N_12249,N_6870,N_9538);
xnor U12250 (N_12250,N_10106,N_11506);
nor U12251 (N_12251,N_10617,N_10865);
nand U12252 (N_12252,N_9923,N_8934);
or U12253 (N_12253,N_11644,N_11548);
or U12254 (N_12254,N_6643,N_9537);
or U12255 (N_12255,N_7198,N_9964);
or U12256 (N_12256,N_7242,N_6944);
or U12257 (N_12257,N_10552,N_8248);
and U12258 (N_12258,N_9546,N_8938);
or U12259 (N_12259,N_7097,N_9420);
nand U12260 (N_12260,N_7894,N_10218);
xnor U12261 (N_12261,N_6503,N_10845);
xnor U12262 (N_12262,N_9042,N_8881);
and U12263 (N_12263,N_10923,N_6093);
nor U12264 (N_12264,N_7231,N_9895);
nand U12265 (N_12265,N_6992,N_11465);
nand U12266 (N_12266,N_10974,N_7257);
or U12267 (N_12267,N_9464,N_11982);
nand U12268 (N_12268,N_11683,N_6118);
nand U12269 (N_12269,N_7499,N_7311);
nand U12270 (N_12270,N_10876,N_9599);
and U12271 (N_12271,N_6900,N_8473);
xor U12272 (N_12272,N_8931,N_10888);
nand U12273 (N_12273,N_9390,N_11335);
nand U12274 (N_12274,N_10996,N_8936);
nand U12275 (N_12275,N_10000,N_10411);
and U12276 (N_12276,N_10429,N_8385);
and U12277 (N_12277,N_10936,N_11793);
nand U12278 (N_12278,N_9414,N_10112);
and U12279 (N_12279,N_9095,N_10879);
or U12280 (N_12280,N_7014,N_8041);
nor U12281 (N_12281,N_11564,N_6662);
nor U12282 (N_12282,N_8625,N_8815);
and U12283 (N_12283,N_7671,N_8592);
or U12284 (N_12284,N_7612,N_7132);
nand U12285 (N_12285,N_8402,N_8384);
or U12286 (N_12286,N_10275,N_6778);
nor U12287 (N_12287,N_8311,N_7888);
and U12288 (N_12288,N_6657,N_11603);
nand U12289 (N_12289,N_6290,N_10754);
and U12290 (N_12290,N_9220,N_9006);
nand U12291 (N_12291,N_7620,N_6401);
nand U12292 (N_12292,N_8238,N_6292);
or U12293 (N_12293,N_9759,N_7399);
nor U12294 (N_12294,N_11472,N_11769);
nand U12295 (N_12295,N_7031,N_9343);
and U12296 (N_12296,N_9462,N_11182);
or U12297 (N_12297,N_11382,N_8672);
or U12298 (N_12298,N_8377,N_10269);
xor U12299 (N_12299,N_11519,N_9966);
xor U12300 (N_12300,N_8659,N_8312);
nor U12301 (N_12301,N_8483,N_9181);
and U12302 (N_12302,N_10566,N_7650);
nor U12303 (N_12303,N_6608,N_10391);
xnor U12304 (N_12304,N_8169,N_11069);
and U12305 (N_12305,N_8234,N_7052);
nor U12306 (N_12306,N_6794,N_7493);
and U12307 (N_12307,N_7522,N_9439);
and U12308 (N_12308,N_11692,N_6649);
xor U12309 (N_12309,N_7759,N_6100);
xor U12310 (N_12310,N_9937,N_10260);
nand U12311 (N_12311,N_7784,N_9519);
nand U12312 (N_12312,N_8159,N_11628);
nor U12313 (N_12313,N_7761,N_9107);
nor U12314 (N_12314,N_6071,N_8046);
xnor U12315 (N_12315,N_11235,N_7972);
or U12316 (N_12316,N_7724,N_9892);
nor U12317 (N_12317,N_10299,N_11255);
and U12318 (N_12318,N_6912,N_6076);
xor U12319 (N_12319,N_7858,N_11325);
nor U12320 (N_12320,N_10336,N_7791);
and U12321 (N_12321,N_7611,N_6230);
nor U12322 (N_12322,N_7725,N_7796);
and U12323 (N_12323,N_8556,N_6562);
nor U12324 (N_12324,N_8271,N_6634);
nor U12325 (N_12325,N_10052,N_6003);
or U12326 (N_12326,N_8990,N_8030);
nand U12327 (N_12327,N_8983,N_6278);
xor U12328 (N_12328,N_7228,N_9986);
xnor U12329 (N_12329,N_8283,N_9753);
or U12330 (N_12330,N_7182,N_10750);
xnor U12331 (N_12331,N_10846,N_9797);
nor U12332 (N_12332,N_7830,N_11442);
or U12333 (N_12333,N_9711,N_10920);
nor U12334 (N_12334,N_7997,N_11837);
nand U12335 (N_12335,N_10554,N_8910);
xor U12336 (N_12336,N_6953,N_10387);
nor U12337 (N_12337,N_11997,N_8961);
and U12338 (N_12338,N_10266,N_9377);
and U12339 (N_12339,N_11127,N_7253);
xor U12340 (N_12340,N_11616,N_11584);
nand U12341 (N_12341,N_6507,N_9603);
nor U12342 (N_12342,N_10853,N_10330);
and U12343 (N_12343,N_10211,N_7726);
nor U12344 (N_12344,N_10756,N_7391);
nor U12345 (N_12345,N_8917,N_7805);
nor U12346 (N_12346,N_8531,N_8114);
nand U12347 (N_12347,N_8150,N_9218);
nand U12348 (N_12348,N_6223,N_6420);
nor U12349 (N_12349,N_8341,N_10302);
nand U12350 (N_12350,N_10493,N_9830);
and U12351 (N_12351,N_7901,N_10887);
or U12352 (N_12352,N_6725,N_8498);
nor U12353 (N_12353,N_11655,N_6226);
and U12354 (N_12354,N_11973,N_7079);
nor U12355 (N_12355,N_9067,N_6165);
and U12356 (N_12356,N_6702,N_8292);
nor U12357 (N_12357,N_8681,N_10141);
or U12358 (N_12358,N_10605,N_7389);
nor U12359 (N_12359,N_9049,N_9499);
nor U12360 (N_12360,N_9514,N_10706);
or U12361 (N_12361,N_6573,N_6142);
nor U12362 (N_12362,N_7593,N_7290);
or U12363 (N_12363,N_10874,N_7093);
nand U12364 (N_12364,N_11419,N_6904);
nand U12365 (N_12365,N_8735,N_8427);
xor U12366 (N_12366,N_8208,N_10568);
or U12367 (N_12367,N_11326,N_11113);
xor U12368 (N_12368,N_9969,N_8440);
and U12369 (N_12369,N_9127,N_6170);
nor U12370 (N_12370,N_9474,N_7267);
or U12371 (N_12371,N_9327,N_9156);
and U12372 (N_12372,N_11923,N_10213);
or U12373 (N_12373,N_11783,N_8898);
and U12374 (N_12374,N_6597,N_8758);
nor U12375 (N_12375,N_9718,N_8260);
nand U12376 (N_12376,N_6344,N_10627);
and U12377 (N_12377,N_10817,N_6853);
or U12378 (N_12378,N_10332,N_9291);
nor U12379 (N_12379,N_11856,N_8474);
nor U12380 (N_12380,N_8807,N_9264);
nor U12381 (N_12381,N_10859,N_6356);
or U12382 (N_12382,N_7756,N_10356);
xor U12383 (N_12383,N_6591,N_6948);
and U12384 (N_12384,N_7779,N_7027);
or U12385 (N_12385,N_9014,N_6959);
and U12386 (N_12386,N_7434,N_10283);
nor U12387 (N_12387,N_11322,N_9212);
nor U12388 (N_12388,N_11134,N_6324);
nor U12389 (N_12389,N_10383,N_9996);
and U12390 (N_12390,N_8033,N_10818);
xnor U12391 (N_12391,N_7651,N_8247);
nor U12392 (N_12392,N_6670,N_6253);
xor U12393 (N_12393,N_8376,N_9004);
nor U12394 (N_12394,N_7214,N_6876);
or U12395 (N_12395,N_7547,N_11249);
and U12396 (N_12396,N_10220,N_6261);
xor U12397 (N_12397,N_9828,N_6060);
xnor U12398 (N_12398,N_7042,N_11951);
or U12399 (N_12399,N_9957,N_9825);
nor U12400 (N_12400,N_7973,N_8746);
and U12401 (N_12401,N_6556,N_10848);
nand U12402 (N_12402,N_7185,N_8835);
or U12403 (N_12403,N_6282,N_11316);
nor U12404 (N_12404,N_6140,N_10652);
xor U12405 (N_12405,N_11581,N_6890);
nor U12406 (N_12406,N_11985,N_7106);
xor U12407 (N_12407,N_10035,N_11971);
xnor U12408 (N_12408,N_11379,N_6294);
nand U12409 (N_12409,N_8230,N_6604);
nor U12410 (N_12410,N_10646,N_8246);
and U12411 (N_12411,N_7801,N_7303);
nand U12412 (N_12412,N_7141,N_9639);
and U12413 (N_12413,N_9236,N_10179);
nor U12414 (N_12414,N_7476,N_11294);
nand U12415 (N_12415,N_10714,N_11868);
xor U12416 (N_12416,N_6557,N_10292);
nor U12417 (N_12417,N_7904,N_10690);
and U12418 (N_12418,N_9143,N_9337);
and U12419 (N_12419,N_8623,N_11393);
xor U12420 (N_12420,N_10650,N_10623);
xnor U12421 (N_12421,N_10777,N_8013);
nand U12422 (N_12422,N_6506,N_11430);
nand U12423 (N_12423,N_9648,N_9297);
and U12424 (N_12424,N_11920,N_7832);
or U12425 (N_12425,N_6834,N_10416);
xor U12426 (N_12426,N_6204,N_10758);
or U12427 (N_12427,N_6219,N_6995);
and U12428 (N_12428,N_10398,N_8298);
xnor U12429 (N_12429,N_11077,N_7720);
nor U12430 (N_12430,N_6304,N_11877);
xor U12431 (N_12431,N_11209,N_10837);
or U12432 (N_12432,N_9109,N_7474);
or U12433 (N_12433,N_6126,N_9712);
nand U12434 (N_12434,N_10390,N_11858);
nand U12435 (N_12435,N_10270,N_8786);
xnor U12436 (N_12436,N_7026,N_11658);
and U12437 (N_12437,N_11552,N_8360);
or U12438 (N_12438,N_9505,N_7432);
xnor U12439 (N_12439,N_11349,N_9246);
nand U12440 (N_12440,N_8398,N_11270);
nor U12441 (N_12441,N_8462,N_10087);
or U12442 (N_12442,N_9290,N_7910);
and U12443 (N_12443,N_9713,N_8500);
xor U12444 (N_12444,N_9458,N_6047);
nor U12445 (N_12445,N_7677,N_10338);
or U12446 (N_12446,N_7148,N_9581);
nand U12447 (N_12447,N_9908,N_7041);
nand U12448 (N_12448,N_6262,N_7840);
nand U12449 (N_12449,N_6390,N_7635);
and U12450 (N_12450,N_7122,N_11344);
nand U12451 (N_12451,N_6399,N_10011);
xor U12452 (N_12452,N_6013,N_10868);
or U12453 (N_12453,N_11932,N_9855);
xor U12454 (N_12454,N_9761,N_8176);
or U12455 (N_12455,N_6521,N_11512);
and U12456 (N_12456,N_8027,N_6106);
nor U12457 (N_12457,N_7715,N_8039);
nor U12458 (N_12458,N_6256,N_7070);
nor U12459 (N_12459,N_9043,N_11358);
or U12460 (N_12460,N_9559,N_6842);
or U12461 (N_12461,N_11126,N_9666);
or U12462 (N_12462,N_10893,N_7486);
or U12463 (N_12463,N_7815,N_11990);
and U12464 (N_12464,N_10089,N_6467);
nand U12465 (N_12465,N_8774,N_7970);
xnor U12466 (N_12466,N_9622,N_8196);
nand U12467 (N_12467,N_9748,N_11007);
or U12468 (N_12468,N_9630,N_11306);
nand U12469 (N_12469,N_9722,N_9806);
or U12470 (N_12470,N_11130,N_11121);
or U12471 (N_12471,N_10396,N_8778);
and U12472 (N_12472,N_6903,N_6250);
nor U12473 (N_12473,N_11542,N_7324);
nand U12474 (N_12474,N_11875,N_7299);
xnor U12475 (N_12475,N_10927,N_11473);
nand U12476 (N_12476,N_6479,N_9931);
or U12477 (N_12477,N_7760,N_9846);
nand U12478 (N_12478,N_6281,N_8325);
and U12479 (N_12479,N_10147,N_10494);
nand U12480 (N_12480,N_11744,N_11313);
and U12481 (N_12481,N_8916,N_11070);
and U12482 (N_12482,N_8737,N_9206);
xor U12483 (N_12483,N_8060,N_9918);
xor U12484 (N_12484,N_6411,N_11028);
nand U12485 (N_12485,N_7537,N_9732);
and U12486 (N_12486,N_9428,N_10206);
nor U12487 (N_12487,N_10062,N_11492);
or U12488 (N_12488,N_9743,N_11736);
or U12489 (N_12489,N_8212,N_11696);
nor U12490 (N_12490,N_9954,N_10078);
and U12491 (N_12491,N_8953,N_10105);
or U12492 (N_12492,N_9378,N_9765);
xor U12493 (N_12493,N_11677,N_11904);
xor U12494 (N_12494,N_6954,N_11771);
or U12495 (N_12495,N_6303,N_8197);
nand U12496 (N_12496,N_7229,N_11873);
nand U12497 (N_12497,N_11507,N_9328);
xnor U12498 (N_12498,N_7271,N_8907);
nor U12499 (N_12499,N_7712,N_11234);
nand U12500 (N_12500,N_7912,N_9217);
nand U12501 (N_12501,N_6914,N_6309);
xor U12502 (N_12502,N_9730,N_10540);
and U12503 (N_12503,N_11577,N_6216);
xor U12504 (N_12504,N_9244,N_11033);
xor U12505 (N_12505,N_7965,N_10905);
nor U12506 (N_12506,N_10234,N_6814);
or U12507 (N_12507,N_9015,N_9692);
or U12508 (N_12508,N_10676,N_9641);
nor U12509 (N_12509,N_8110,N_11097);
xor U12510 (N_12510,N_11580,N_8870);
nand U12511 (N_12511,N_7451,N_7527);
nor U12512 (N_12512,N_9671,N_8233);
nor U12513 (N_12513,N_11023,N_10376);
nand U12514 (N_12514,N_8086,N_6081);
xor U12515 (N_12515,N_7777,N_9129);
xor U12516 (N_12516,N_8074,N_7119);
or U12517 (N_12517,N_10449,N_7067);
and U12518 (N_12518,N_9767,N_9058);
nand U12519 (N_12519,N_9500,N_7217);
and U12520 (N_12520,N_10482,N_7998);
and U12521 (N_12521,N_9977,N_7570);
xor U12522 (N_12522,N_7068,N_8945);
nand U12523 (N_12523,N_9081,N_6409);
nand U12524 (N_12524,N_6547,N_10175);
or U12525 (N_12525,N_10807,N_6231);
nand U12526 (N_12526,N_6698,N_11183);
or U12527 (N_12527,N_11952,N_11585);
nor U12528 (N_12528,N_9983,N_7511);
nand U12529 (N_12529,N_6307,N_11832);
nor U12530 (N_12530,N_8450,N_9257);
nand U12531 (N_12531,N_11271,N_11691);
nand U12532 (N_12532,N_8645,N_9365);
or U12533 (N_12533,N_8205,N_6160);
or U12534 (N_12534,N_10233,N_8194);
xnor U12535 (N_12535,N_11817,N_6233);
or U12536 (N_12536,N_8600,N_10190);
nor U12537 (N_12537,N_11802,N_9685);
or U12538 (N_12538,N_10573,N_6648);
and U12539 (N_12539,N_7774,N_8102);
or U12540 (N_12540,N_11641,N_11135);
nor U12541 (N_12541,N_9469,N_9262);
nor U12542 (N_12542,N_8245,N_11336);
xor U12543 (N_12543,N_7782,N_9935);
nor U12544 (N_12544,N_11152,N_9125);
nor U12545 (N_12545,N_10397,N_7307);
or U12546 (N_12546,N_6168,N_9959);
and U12547 (N_12547,N_6190,N_9086);
nand U12548 (N_12548,N_6136,N_8589);
xnor U12549 (N_12549,N_8229,N_10620);
xnor U12550 (N_12550,N_10100,N_6612);
or U12551 (N_12551,N_6021,N_10970);
nand U12552 (N_12552,N_7322,N_6452);
and U12553 (N_12553,N_11380,N_7713);
nor U12554 (N_12554,N_11883,N_10537);
or U12555 (N_12555,N_9638,N_10282);
xor U12556 (N_12556,N_7351,N_8432);
nor U12557 (N_12557,N_6519,N_11317);
and U12558 (N_12558,N_8137,N_8944);
or U12559 (N_12559,N_7350,N_7749);
and U12560 (N_12560,N_8670,N_6537);
or U12561 (N_12561,N_7170,N_7536);
nand U12562 (N_12562,N_9542,N_7728);
xor U12563 (N_12563,N_9802,N_7985);
or U12564 (N_12564,N_11758,N_6972);
nand U12565 (N_12565,N_11831,N_6158);
nor U12566 (N_12566,N_6962,N_7039);
xor U12567 (N_12567,N_11885,N_6549);
or U12568 (N_12568,N_6065,N_10558);
nor U12569 (N_12569,N_9920,N_11057);
nand U12570 (N_12570,N_9433,N_7323);
or U12571 (N_12571,N_8203,N_8061);
nand U12572 (N_12572,N_10399,N_8651);
nor U12573 (N_12573,N_7175,N_8691);
xor U12574 (N_12574,N_8982,N_8170);
xnor U12575 (N_12575,N_6055,N_9800);
nand U12576 (N_12576,N_10261,N_11177);
nand U12577 (N_12577,N_7773,N_9391);
or U12578 (N_12578,N_6595,N_9192);
nand U12579 (N_12579,N_7948,N_7238);
xnor U12580 (N_12580,N_7002,N_9976);
and U12581 (N_12581,N_7204,N_9583);
nand U12582 (N_12582,N_6120,N_6434);
nor U12583 (N_12583,N_8261,N_11854);
and U12584 (N_12584,N_10149,N_11977);
nor U12585 (N_12585,N_8968,N_8999);
or U12586 (N_12586,N_9669,N_9812);
nor U12587 (N_12587,N_6730,N_8287);
xor U12588 (N_12588,N_8676,N_7482);
or U12589 (N_12589,N_8890,N_8320);
nor U12590 (N_12590,N_11626,N_6862);
nand U12591 (N_12591,N_10599,N_10597);
or U12592 (N_12592,N_10979,N_10070);
nand U12593 (N_12593,N_6973,N_6002);
and U12594 (N_12594,N_9557,N_8615);
or U12595 (N_12595,N_6001,N_9011);
xor U12596 (N_12596,N_9501,N_6583);
nor U12597 (N_12597,N_7120,N_10663);
and U12598 (N_12598,N_11713,N_10405);
nor U12599 (N_12599,N_6006,N_10746);
nand U12600 (N_12600,N_7687,N_11772);
or U12601 (N_12601,N_10950,N_7574);
xnor U12602 (N_12602,N_9714,N_11728);
xor U12603 (N_12603,N_10355,N_7714);
nor U12604 (N_12604,N_9037,N_6129);
and U12605 (N_12605,N_10378,N_11870);
nor U12606 (N_12606,N_6738,N_6559);
or U12607 (N_12607,N_10790,N_6460);
xor U12608 (N_12608,N_11747,N_11815);
xor U12609 (N_12609,N_10513,N_9506);
or U12610 (N_12610,N_9310,N_7077);
nor U12611 (N_12611,N_9157,N_7442);
or U12612 (N_12612,N_10577,N_9245);
and U12613 (N_12613,N_8165,N_8482);
or U12614 (N_12614,N_11053,N_11124);
nand U12615 (N_12615,N_11231,N_8472);
and U12616 (N_12616,N_6276,N_11556);
nor U12617 (N_12617,N_8251,N_11086);
xor U12618 (N_12618,N_11216,N_11059);
and U12619 (N_12619,N_10184,N_7627);
and U12620 (N_12620,N_11224,N_10668);
nand U12621 (N_12621,N_7195,N_8124);
and U12622 (N_12622,N_6789,N_9792);
xor U12623 (N_12623,N_6716,N_11765);
and U12624 (N_12624,N_11927,N_9355);
nor U12625 (N_12625,N_8570,N_7174);
nand U12626 (N_12626,N_11527,N_10277);
xor U12627 (N_12627,N_11667,N_6671);
nand U12628 (N_12628,N_11279,N_6178);
or U12629 (N_12629,N_8448,N_10033);
xor U12630 (N_12630,N_11535,N_7478);
or U12631 (N_12631,N_10721,N_10911);
or U12632 (N_12632,N_11240,N_7448);
nand U12633 (N_12633,N_10518,N_8641);
nor U12634 (N_12634,N_7500,N_7117);
nor U12635 (N_12635,N_7990,N_11602);
nor U12636 (N_12636,N_7559,N_11470);
nor U12637 (N_12637,N_7960,N_11418);
and U12638 (N_12638,N_8549,N_9707);
or U12639 (N_12639,N_6297,N_9101);
and U12640 (N_12640,N_8451,N_9497);
nor U12641 (N_12641,N_9667,N_7873);
or U12642 (N_12642,N_8464,N_11157);
nand U12643 (N_12643,N_11269,N_8175);
and U12644 (N_12644,N_10058,N_9985);
nor U12645 (N_12645,N_9476,N_9643);
and U12646 (N_12646,N_11056,N_7986);
or U12647 (N_12647,N_10039,N_7440);
xnor U12648 (N_12648,N_6336,N_10783);
or U12649 (N_12649,N_6289,N_8365);
or U12650 (N_12650,N_11376,N_9949);
xor U12651 (N_12651,N_7413,N_7646);
or U12652 (N_12652,N_10542,N_11173);
or U12653 (N_12653,N_8355,N_8966);
nand U12654 (N_12654,N_10410,N_7269);
nor U12655 (N_12655,N_6306,N_8301);
or U12656 (N_12656,N_9885,N_8367);
nor U12657 (N_12657,N_9826,N_11450);
xor U12658 (N_12658,N_10532,N_8538);
or U12659 (N_12659,N_8106,N_8627);
and U12660 (N_12660,N_8134,N_7199);
xor U12661 (N_12661,N_8001,N_10054);
or U12662 (N_12662,N_10116,N_6139);
and U12663 (N_12663,N_6000,N_10588);
xor U12664 (N_12664,N_9247,N_6667);
nand U12665 (N_12665,N_11611,N_10469);
and U12666 (N_12666,N_9960,N_6104);
and U12667 (N_12667,N_11268,N_7789);
and U12668 (N_12668,N_8866,N_6552);
xnor U12669 (N_12669,N_10379,N_11666);
nand U12670 (N_12670,N_7301,N_7802);
xnor U12671 (N_12671,N_11258,N_11540);
xnor U12672 (N_12672,N_6132,N_10613);
nand U12673 (N_12673,N_8022,N_8342);
nor U12674 (N_12674,N_10464,N_6711);
nand U12675 (N_12675,N_6619,N_11693);
xnor U12676 (N_12676,N_8788,N_10603);
nor U12677 (N_12677,N_8857,N_11609);
nor U12678 (N_12678,N_10085,N_7463);
xor U12679 (N_12679,N_11314,N_9524);
or U12680 (N_12680,N_6299,N_8331);
or U12681 (N_12681,N_6748,N_10059);
xnor U12682 (N_12682,N_8925,N_10674);
or U12683 (N_12683,N_11403,N_10722);
nand U12684 (N_12684,N_7878,N_10771);
or U12685 (N_12685,N_10090,N_11780);
nor U12686 (N_12686,N_10924,N_8300);
and U12687 (N_12687,N_7709,N_8087);
xnor U12688 (N_12688,N_6177,N_10221);
and U12689 (N_12689,N_7412,N_6739);
or U12690 (N_12690,N_11438,N_8553);
nor U12691 (N_12691,N_9231,N_6878);
xnor U12692 (N_12692,N_8871,N_6395);
and U12693 (N_12693,N_11129,N_8173);
nor U12694 (N_12694,N_8545,N_6820);
xnor U12695 (N_12695,N_8698,N_10187);
nor U12696 (N_12696,N_6032,N_8955);
nand U12697 (N_12697,N_11708,N_8380);
xnor U12698 (N_12698,N_11513,N_9108);
nor U12699 (N_12699,N_8525,N_10239);
xnor U12700 (N_12700,N_6719,N_10041);
nand U12701 (N_12701,N_11159,N_6865);
xnor U12702 (N_12702,N_11848,N_6328);
nor U12703 (N_12703,N_6841,N_8379);
xor U12704 (N_12704,N_10828,N_8273);
and U12705 (N_12705,N_11918,N_6950);
xnor U12706 (N_12706,N_11819,N_6741);
nor U12707 (N_12707,N_10711,N_9048);
or U12708 (N_12708,N_10252,N_11420);
xnor U12709 (N_12709,N_7795,N_11795);
nor U12710 (N_12710,N_7221,N_8417);
nor U12711 (N_12711,N_7181,N_8696);
nand U12712 (N_12712,N_11175,N_6529);
nor U12713 (N_12713,N_9627,N_11634);
nor U12714 (N_12714,N_8858,N_11448);
nor U12715 (N_12715,N_9003,N_8865);
and U12716 (N_12716,N_8617,N_7398);
nand U12717 (N_12717,N_10524,N_10114);
or U12718 (N_12718,N_9770,N_11686);
nor U12719 (N_12719,N_9186,N_10463);
xnor U12720 (N_12720,N_6881,N_11291);
xor U12721 (N_12721,N_6239,N_10831);
xnor U12722 (N_12722,N_10545,N_10514);
xor U12723 (N_12723,N_6108,N_10692);
nor U12724 (N_12724,N_10761,N_10504);
and U12725 (N_12725,N_8878,N_8489);
xor U12726 (N_12726,N_7669,N_8503);
nand U12727 (N_12727,N_8050,N_6970);
or U12728 (N_12728,N_7698,N_8653);
nand U12729 (N_12729,N_8926,N_11254);
nor U12730 (N_12730,N_9656,N_9405);
and U12731 (N_12731,N_10393,N_11217);
and U12732 (N_12732,N_9703,N_6637);
xnor U12733 (N_12733,N_10670,N_10544);
nand U12734 (N_12734,N_8971,N_6705);
and U12735 (N_12735,N_6392,N_6938);
xnor U12736 (N_12736,N_6927,N_10177);
and U12737 (N_12737,N_10901,N_7844);
nand U12738 (N_12738,N_7306,N_7340);
xor U12739 (N_12739,N_7380,N_11732);
nand U12740 (N_12740,N_7156,N_9023);
or U12741 (N_12741,N_8765,N_9319);
and U12742 (N_12742,N_6613,N_11979);
nor U12743 (N_12743,N_11455,N_8168);
and U12744 (N_12744,N_8352,N_11816);
or U12745 (N_12745,N_7347,N_7277);
nor U12746 (N_12746,N_11986,N_8415);
nand U12747 (N_12747,N_7452,N_11698);
and U12748 (N_12748,N_10276,N_6863);
and U12749 (N_12749,N_8834,N_9883);
nand U12750 (N_12750,N_11042,N_9164);
and U12751 (N_12751,N_11647,N_9490);
and U12752 (N_12752,N_6607,N_6951);
and U12753 (N_12753,N_6568,N_6483);
nand U12754 (N_12754,N_9438,N_7666);
xor U12755 (N_12755,N_10369,N_6596);
xor U12756 (N_12756,N_8717,N_8037);
nand U12757 (N_12757,N_10362,N_10348);
nor U12758 (N_12758,N_7121,N_11265);
and U12759 (N_12759,N_9747,N_9061);
and U12760 (N_12760,N_9075,N_8609);
nand U12761 (N_12761,N_8817,N_9334);
nand U12762 (N_12762,N_9984,N_11850);
nor U12763 (N_12763,N_9035,N_11823);
nand U12764 (N_12764,N_6594,N_11475);
and U12765 (N_12765,N_7877,N_9057);
and U12766 (N_12766,N_6124,N_10238);
or U12767 (N_12767,N_6463,N_11411);
nand U12768 (N_12768,N_7771,N_6387);
or U12769 (N_12769,N_10688,N_8962);
nand U12770 (N_12770,N_6322,N_7431);
nand U12771 (N_12771,N_10640,N_9502);
and U12772 (N_12772,N_9768,N_7096);
or U12773 (N_12773,N_9555,N_11493);
or U12774 (N_12774,N_11730,N_11845);
nor U12775 (N_12775,N_7863,N_8707);
xor U12776 (N_12776,N_8985,N_10406);
nor U12777 (N_12777,N_9927,N_8728);
nor U12778 (N_12778,N_6764,N_6027);
nand U12779 (N_12779,N_8524,N_9616);
nand U12780 (N_12780,N_9370,N_8518);
and U12781 (N_12781,N_8335,N_9773);
nor U12782 (N_12782,N_6689,N_10014);
and U12783 (N_12783,N_6986,N_10450);
and U12784 (N_12784,N_7273,N_9591);
and U12785 (N_12785,N_10012,N_8567);
or U12786 (N_12786,N_10439,N_9997);
nand U12787 (N_12787,N_11227,N_7126);
nor U12788 (N_12788,N_6075,N_10547);
xor U12789 (N_12789,N_9059,N_10134);
nand U12790 (N_12790,N_7813,N_7678);
xnor U12791 (N_12791,N_8054,N_10675);
xor U12792 (N_12792,N_7694,N_10870);
nand U12793 (N_12793,N_6822,N_11839);
nand U12794 (N_12794,N_7428,N_8409);
xor U12795 (N_12795,N_9869,N_6345);
or U12796 (N_12796,N_10842,N_9171);
xor U12797 (N_12797,N_9461,N_7887);
or U12798 (N_12798,N_11466,N_10998);
nor U12799 (N_12799,N_8918,N_10272);
nor U12800 (N_12800,N_9901,N_6408);
xnor U12801 (N_12801,N_9403,N_10798);
and U12802 (N_12802,N_7161,N_9496);
nor U12803 (N_12803,N_6874,N_9139);
or U12804 (N_12804,N_11458,N_7314);
and U12805 (N_12805,N_6288,N_11505);
nand U12806 (N_12806,N_8833,N_11946);
or U12807 (N_12807,N_9289,N_8042);
xnor U12808 (N_12808,N_7563,N_9833);
xnor U12809 (N_12809,N_8339,N_11804);
nand U12810 (N_12810,N_7408,N_8403);
nor U12811 (N_12811,N_7137,N_7145);
and U12812 (N_12812,N_8113,N_7765);
and U12813 (N_12813,N_7923,N_10891);
xnor U12814 (N_12814,N_7072,N_7421);
nor U12815 (N_12815,N_10004,N_6964);
nand U12816 (N_12816,N_10766,N_7585);
nand U12817 (N_12817,N_6143,N_9521);
nand U12818 (N_12818,N_7104,N_8896);
and U12819 (N_12819,N_7144,N_11301);
and U12820 (N_12820,N_8739,N_7087);
nand U12821 (N_12821,N_7551,N_8548);
and U12822 (N_12822,N_7957,N_7827);
or U12823 (N_12823,N_9489,N_10196);
nand U12824 (N_12824,N_9781,N_9820);
xor U12825 (N_12825,N_9879,N_11663);
or U12826 (N_12826,N_9207,N_6300);
or U12827 (N_12827,N_6800,N_9113);
or U12828 (N_12828,N_9084,N_10448);
nand U12829 (N_12829,N_7099,N_6722);
or U12830 (N_12830,N_7060,N_10725);
and U12831 (N_12831,N_8439,N_7394);
xnor U12832 (N_12832,N_11161,N_9853);
or U12833 (N_12833,N_11228,N_9681);
or U12834 (N_12834,N_8797,N_11808);
nand U12835 (N_12835,N_11345,N_10967);
and U12836 (N_12836,N_8602,N_7898);
or U12837 (N_12837,N_11168,N_9975);
xnor U12838 (N_12838,N_6724,N_8867);
nand U12839 (N_12839,N_8307,N_11668);
or U12840 (N_12840,N_11244,N_9847);
and U12841 (N_12841,N_6085,N_10067);
nor U12842 (N_12842,N_10502,N_8202);
nand U12843 (N_12843,N_7866,N_9208);
xor U12844 (N_12844,N_8057,N_7680);
nor U12845 (N_12845,N_6798,N_6664);
and U12846 (N_12846,N_6517,N_8392);
and U12847 (N_12847,N_10146,N_11908);
or U12848 (N_12848,N_11572,N_8393);
nand U12849 (N_12849,N_7128,N_6385);
nand U12850 (N_12850,N_7165,N_8120);
or U12851 (N_12851,N_6199,N_8674);
nand U12852 (N_12852,N_11005,N_6751);
or U12853 (N_12853,N_6511,N_8872);
or U12854 (N_12854,N_10975,N_6425);
and U12855 (N_12855,N_6218,N_11378);
and U12856 (N_12856,N_8445,N_11637);
and U12857 (N_12857,N_9609,N_9052);
xor U12858 (N_12858,N_10838,N_11114);
nand U12859 (N_12859,N_8133,N_7426);
nand U12860 (N_12860,N_6117,N_8963);
and U12861 (N_12861,N_6796,N_6759);
and U12862 (N_12862,N_10938,N_7333);
and U12863 (N_12863,N_7461,N_11377);
nand U12864 (N_12864,N_10829,N_8015);
nor U12865 (N_12865,N_9435,N_6248);
nor U12866 (N_12866,N_8539,N_11916);
xnor U12867 (N_12867,N_6750,N_11405);
or U12868 (N_12868,N_11809,N_9827);
xnor U12869 (N_12869,N_8223,N_10631);
nor U12870 (N_12870,N_10614,N_10176);
and U12871 (N_12871,N_9402,N_7502);
and U12872 (N_12872,N_7820,N_9592);
nor U12873 (N_12873,N_8032,N_7554);
and U12874 (N_12874,N_6772,N_9457);
nand U12875 (N_12875,N_9237,N_7091);
nor U12876 (N_12876,N_11461,N_11528);
and U12877 (N_12877,N_8565,N_9320);
or U12878 (N_12878,N_10687,N_7999);
or U12879 (N_12879,N_11664,N_6807);
xor U12880 (N_12880,N_6319,N_6017);
nand U12881 (N_12881,N_6374,N_6478);
and U12882 (N_12882,N_7655,N_6543);
nor U12883 (N_12883,N_11332,N_11284);
xor U12884 (N_12884,N_11145,N_10578);
and U12885 (N_12885,N_9958,N_10322);
or U12886 (N_12886,N_7757,N_9645);
xor U12887 (N_12887,N_7994,N_8560);
nand U12888 (N_12888,N_10508,N_8052);
nand U12889 (N_12889,N_7629,N_10180);
nand U12890 (N_12890,N_9553,N_8642);
and U12891 (N_12891,N_6587,N_10576);
or U12892 (N_12892,N_6080,N_11699);
or U12893 (N_12893,N_11999,N_8949);
nor U12894 (N_12894,N_10363,N_6611);
and U12895 (N_12895,N_10731,N_10235);
or U12896 (N_12896,N_7250,N_11867);
xor U12897 (N_12897,N_10343,N_11887);
xor U12898 (N_12898,N_6894,N_10792);
nand U12899 (N_12899,N_9868,N_7751);
nor U12900 (N_12900,N_6620,N_8832);
xor U12901 (N_12901,N_7595,N_11487);
xor U12902 (N_12902,N_9933,N_10225);
and U12903 (N_12903,N_9570,N_6956);
nand U12904 (N_12904,N_7518,N_6255);
nor U12905 (N_12905,N_7816,N_11030);
and U12906 (N_12906,N_8843,N_10789);
nand U12907 (N_12907,N_9446,N_11589);
nand U12908 (N_12908,N_7180,N_11139);
xnor U12909 (N_12909,N_11247,N_6427);
and U12910 (N_12910,N_7248,N_8227);
or U12911 (N_12911,N_6241,N_11866);
and U12912 (N_12912,N_8006,N_10651);
or U12913 (N_12913,N_6088,N_8587);
xnor U12914 (N_12914,N_8743,N_10143);
or U12915 (N_12915,N_8956,N_6128);
nor U12916 (N_12916,N_11304,N_9051);
or U12917 (N_12917,N_6422,N_9729);
or U12918 (N_12918,N_11079,N_7920);
and U12919 (N_12919,N_11406,N_7754);
or U12920 (N_12920,N_6348,N_10556);
and U12921 (N_12921,N_7458,N_7849);
xnor U12922 (N_12922,N_6333,N_8064);
and U12923 (N_12923,N_7024,N_11039);
and U12924 (N_12924,N_8241,N_10295);
nand U12925 (N_12925,N_6171,N_8188);
or U12926 (N_12926,N_10166,N_7098);
xor U12927 (N_12927,N_10833,N_11640);
or U12928 (N_12928,N_10720,N_10458);
or U12929 (N_12929,N_8964,N_6677);
xor U12930 (N_12930,N_7368,N_6906);
xnor U12931 (N_12931,N_8487,N_7523);
or U12932 (N_12932,N_7100,N_9448);
nor U12933 (N_12933,N_7353,N_11485);
and U12934 (N_12934,N_11486,N_9415);
nand U12935 (N_12935,N_8097,N_6955);
xor U12936 (N_12936,N_6810,N_11751);
xor U12937 (N_12937,N_7073,N_10409);
and U12938 (N_12938,N_8756,N_10589);
nand U12939 (N_12939,N_10268,N_9936);
or U12940 (N_12940,N_9487,N_8928);
nand U12941 (N_12941,N_9636,N_10916);
and U12942 (N_12942,N_9794,N_6330);
or U12943 (N_12943,N_9338,N_7911);
and U12944 (N_12944,N_7790,N_11413);
and U12945 (N_12945,N_6308,N_6123);
nand U12946 (N_12946,N_6576,N_11286);
and U12947 (N_12947,N_10649,N_6079);
and U12948 (N_12948,N_8597,N_7285);
and U12949 (N_12949,N_9316,N_9278);
or U12950 (N_12950,N_6771,N_7924);
nand U12951 (N_12951,N_7044,N_11681);
xnor U12952 (N_12952,N_10802,N_8800);
nand U12953 (N_12953,N_8511,N_10727);
nor U12954 (N_12954,N_11500,N_10344);
or U12955 (N_12955,N_9897,N_7485);
nor U12956 (N_12956,N_8713,N_8211);
xor U12957 (N_12957,N_8048,N_9705);
or U12958 (N_12958,N_9528,N_6403);
xor U12959 (N_12959,N_8997,N_11558);
nor U12960 (N_12960,N_9329,N_10812);
or U12961 (N_12961,N_8334,N_9480);
or U12962 (N_12962,N_11720,N_8780);
and U12963 (N_12963,N_10364,N_9135);
nand U12964 (N_12964,N_6721,N_7900);
or U12965 (N_12965,N_8781,N_9595);
or U12966 (N_12966,N_9558,N_8761);
xor U12967 (N_12967,N_7179,N_6014);
nand U12968 (N_12968,N_8214,N_10952);
xor U12969 (N_12969,N_7115,N_10521);
xor U12970 (N_12970,N_9050,N_9486);
xnor U12971 (N_12971,N_9689,N_6078);
nor U12972 (N_12972,N_8730,N_6134);
xnor U12973 (N_12973,N_9384,N_8479);
nor U12974 (N_12974,N_11976,N_10197);
and U12975 (N_12975,N_9025,N_9793);
nand U12976 (N_12976,N_6675,N_8975);
xnor U12977 (N_12977,N_9317,N_6635);
and U12978 (N_12978,N_11034,N_11503);
or U12979 (N_12979,N_8405,N_6654);
nand U12980 (N_12980,N_7959,N_10099);
and U12981 (N_12981,N_8935,N_7374);
nor U12982 (N_12982,N_11488,N_9168);
or U12983 (N_12983,N_8527,N_10844);
xor U12984 (N_12984,N_8747,N_11724);
nand U12985 (N_12985,N_9864,N_6030);
or U12986 (N_12986,N_11962,N_11093);
nor U12987 (N_12987,N_7006,N_6490);
and U12988 (N_12988,N_10333,N_8466);
and U12989 (N_12989,N_7882,N_7101);
and U12990 (N_12990,N_10983,N_9226);
xnor U12991 (N_12991,N_10935,N_6815);
and U12992 (N_12992,N_6358,N_10629);
and U12993 (N_12993,N_9368,N_6570);
nor U12994 (N_12994,N_6921,N_11080);
and U12995 (N_12995,N_11196,N_6699);
xnor U12996 (N_12996,N_9019,N_8101);
or U12997 (N_12997,N_9105,N_7550);
or U12998 (N_12998,N_11449,N_10312);
nor U12999 (N_12999,N_10491,N_10884);
nand U13000 (N_13000,N_7316,N_11716);
or U13001 (N_13001,N_7037,N_6606);
nand U13002 (N_13002,N_10290,N_8382);
nor U13003 (N_13003,N_6879,N_7118);
xor U13004 (N_13004,N_9240,N_9018);
xor U13005 (N_13005,N_11178,N_7514);
xor U13006 (N_13006,N_8668,N_6446);
nor U13007 (N_13007,N_10990,N_8470);
or U13008 (N_13008,N_11888,N_11902);
nand U13009 (N_13009,N_7284,N_7176);
nand U13010 (N_13010,N_10477,N_11871);
or U13011 (N_13011,N_11123,N_7143);
nor U13012 (N_13012,N_8646,N_10509);
or U13013 (N_13013,N_7187,N_8853);
or U13014 (N_13014,N_11141,N_9223);
or U13015 (N_13015,N_10666,N_9693);
xor U13016 (N_13016,N_7422,N_7778);
nand U13017 (N_13017,N_7154,N_10335);
and U13018 (N_13018,N_10921,N_7708);
xnor U13019 (N_13019,N_10869,N_9924);
xnor U13020 (N_13020,N_6049,N_7656);
and U13021 (N_13021,N_7397,N_8084);
nor U13022 (N_13022,N_11820,N_7746);
and U13023 (N_13023,N_7549,N_8559);
and U13024 (N_13024,N_9114,N_10472);
nand U13025 (N_13025,N_9089,N_9013);
nor U13026 (N_13026,N_11399,N_11903);
xnor U13027 (N_13027,N_9715,N_7305);
and U13028 (N_13028,N_6450,N_7053);
nor U13029 (N_13029,N_11478,N_10013);
xor U13030 (N_13030,N_7467,N_7131);
or U13031 (N_13031,N_10341,N_11038);
xnor U13032 (N_13032,N_8541,N_10110);
or U13033 (N_13033,N_8633,N_6609);
or U13034 (N_13034,N_7519,N_6642);
xor U13035 (N_13035,N_11444,N_11431);
nor U13036 (N_13036,N_6901,N_9974);
nand U13037 (N_13037,N_11075,N_9556);
xnor U13038 (N_13038,N_9796,N_10005);
nand U13039 (N_13039,N_11087,N_7332);
and U13040 (N_13040,N_8766,N_6732);
nor U13041 (N_13041,N_6621,N_9345);
or U13042 (N_13042,N_6315,N_7571);
xor U13043 (N_13043,N_11501,N_11650);
xnor U13044 (N_13044,N_10962,N_10030);
nor U13045 (N_13045,N_10388,N_8299);
and U13046 (N_13046,N_8411,N_11071);
nand U13047 (N_13047,N_9540,N_8480);
xnor U13048 (N_13048,N_7665,N_7363);
nor U13049 (N_13049,N_9032,N_11032);
xor U13050 (N_13050,N_8793,N_8184);
or U13051 (N_13051,N_11598,N_8067);
or U13052 (N_13052,N_7625,N_11295);
nand U13053 (N_13053,N_7526,N_8528);
and U13054 (N_13054,N_9177,N_11094);
nor U13055 (N_13055,N_6545,N_8787);
nand U13056 (N_13056,N_9894,N_9840);
nor U13057 (N_13057,N_11432,N_11775);
nand U13058 (N_13058,N_8209,N_8147);
and U13059 (N_13059,N_10288,N_9421);
xnor U13060 (N_13060,N_7338,N_8555);
nor U13061 (N_13061,N_8848,N_9700);
or U13062 (N_13062,N_10959,N_9704);
nor U13063 (N_13063,N_11974,N_10636);
or U13064 (N_13064,N_9099,N_7553);
or U13065 (N_13065,N_6598,N_11081);
and U13066 (N_13066,N_11409,N_8347);
nor U13067 (N_13067,N_11388,N_10839);
or U13068 (N_13068,N_10072,N_10068);
nand U13069 (N_13069,N_10759,N_9673);
nor U13070 (N_13070,N_6971,N_9889);
nand U13071 (N_13071,N_10747,N_10232);
or U13072 (N_13072,N_10980,N_10139);
and U13073 (N_13073,N_8284,N_7996);
and U13074 (N_13074,N_7287,N_11009);
xor U13075 (N_13075,N_8213,N_11675);
or U13076 (N_13076,N_7129,N_10779);
nor U13077 (N_13077,N_8694,N_9330);
nand U13078 (N_13078,N_6895,N_6242);
nand U13079 (N_13079,N_9637,N_7220);
nor U13080 (N_13080,N_9565,N_9929);
xor U13081 (N_13081,N_11013,N_8894);
and U13082 (N_13082,N_9972,N_11412);
nor U13083 (N_13083,N_6114,N_7507);
or U13084 (N_13084,N_11062,N_11119);
nor U13085 (N_13085,N_7831,N_8695);
nand U13086 (N_13086,N_6558,N_9024);
nand U13087 (N_13087,N_8073,N_11891);
nor U13088 (N_13088,N_11357,N_11425);
nor U13089 (N_13089,N_10080,N_7578);
and U13090 (N_13090,N_11968,N_8680);
nand U13091 (N_13091,N_8324,N_8000);
nand U13092 (N_13092,N_7349,N_10867);
xnor U13093 (N_13093,N_10821,N_9407);
and U13094 (N_13094,N_9137,N_7494);
nand U13095 (N_13095,N_6936,N_6459);
or U13096 (N_13096,N_11818,N_7552);
and U13097 (N_13097,N_6206,N_6094);
nand U13098 (N_13098,N_7572,N_11278);
xnor U13099 (N_13099,N_7196,N_6565);
xor U13100 (N_13100,N_9766,N_11471);
nor U13101 (N_13101,N_11928,N_11187);
or U13102 (N_13102,N_6919,N_10340);
or U13103 (N_13103,N_10446,N_6966);
and U13104 (N_13104,N_7786,N_6147);
nand U13105 (N_13105,N_10699,N_11354);
or U13106 (N_13106,N_9367,N_7769);
nand U13107 (N_13107,N_6752,N_6808);
nor U13108 (N_13108,N_6779,N_8710);
nand U13109 (N_13109,N_6760,N_11614);
nand U13110 (N_13110,N_9531,N_11055);
nor U13111 (N_13111,N_10339,N_7166);
nand U13112 (N_13112,N_6381,N_9865);
nor U13113 (N_13113,N_7907,N_11575);
and U13114 (N_13114,N_11764,N_7945);
xor U13115 (N_13115,N_10044,N_6522);
and U13116 (N_13116,N_7047,N_6701);
nand U13117 (N_13117,N_7411,N_6482);
or U13118 (N_13118,N_11148,N_7516);
and U13119 (N_13119,N_9066,N_11395);
xnor U13120 (N_13120,N_11619,N_11060);
nor U13121 (N_13121,N_8509,N_10815);
and U13122 (N_13122,N_10130,N_6913);
and U13123 (N_13123,N_9243,N_9242);
xor U13124 (N_13124,N_11629,N_6349);
or U13125 (N_13125,N_10659,N_9261);
nor U13126 (N_13126,N_11421,N_8891);
and U13127 (N_13127,N_11323,N_8199);
nand U13128 (N_13128,N_10466,N_11978);
nand U13129 (N_13129,N_10810,N_9562);
nand U13130 (N_13130,N_11158,N_9239);
nor U13131 (N_13131,N_9366,N_11959);
or U13132 (N_13132,N_9241,N_8373);
xor U13133 (N_13133,N_8939,N_10245);
nand U13134 (N_13134,N_9341,N_7364);
and U13135 (N_13135,N_11789,N_11700);
nand U13136 (N_13136,N_8383,N_6923);
and U13137 (N_13137,N_7146,N_7260);
and U13138 (N_13138,N_9251,N_6727);
or U13139 (N_13139,N_8992,N_9940);
xnor U13140 (N_13140,N_11356,N_8085);
nand U13141 (N_13141,N_9741,N_6015);
xor U13142 (N_13142,N_9617,N_9613);
xnor U13143 (N_13143,N_10102,N_10281);
and U13144 (N_13144,N_6210,N_10634);
xnor U13145 (N_13145,N_11048,N_11339);
nand U13146 (N_13146,N_10548,N_6673);
xor U13147 (N_13147,N_9687,N_11635);
nor U13148 (N_13148,N_11372,N_7264);
nor U13149 (N_13149,N_11499,N_10056);
xnor U13150 (N_13150,N_7797,N_8523);
or U13151 (N_13151,N_7459,N_11415);
nand U13152 (N_13152,N_8127,N_9335);
and U13153 (N_13153,N_6314,N_6023);
and U13154 (N_13154,N_9861,N_6641);
nor U13155 (N_13155,N_6489,N_9484);
nand U13156 (N_13156,N_10717,N_8210);
and U13157 (N_13157,N_9870,N_8317);
and U13158 (N_13158,N_7693,N_6672);
nand U13159 (N_13159,N_9065,N_9263);
xor U13160 (N_13160,N_8400,N_7503);
nand U13161 (N_13161,N_7548,N_7295);
and U13162 (N_13162,N_11026,N_9293);
xnor U13163 (N_13163,N_6347,N_7584);
or U13164 (N_13164,N_9682,N_10161);
nand U13165 (N_13165,N_8927,N_10561);
or U13166 (N_13166,N_11960,N_10031);
nand U13167 (N_13167,N_10420,N_6283);
nor U13168 (N_13168,N_10457,N_10716);
and U13169 (N_13169,N_8724,N_9772);
xnor U13170 (N_13170,N_7471,N_9034);
nand U13171 (N_13171,N_7534,N_9837);
nor U13172 (N_13172,N_7058,N_7023);
or U13173 (N_13173,N_10499,N_6855);
or U13174 (N_13174,N_9739,N_8446);
nor U13175 (N_13175,N_6153,N_9342);
and U13176 (N_13176,N_9779,N_9680);
nor U13177 (N_13177,N_8322,N_6127);
nand U13178 (N_13178,N_11662,N_11520);
or U13179 (N_13179,N_8569,N_11373);
xor U13180 (N_13180,N_7691,N_7993);
xor U13181 (N_13181,N_11705,N_9817);
and U13182 (N_13182,N_11901,N_11922);
nor U13183 (N_13183,N_10185,N_10265);
nor U13184 (N_13184,N_11101,N_10740);
and U13185 (N_13185,N_6382,N_11012);
or U13186 (N_13186,N_8777,N_9307);
and U13187 (N_13187,N_11355,N_11281);
or U13188 (N_13188,N_11880,N_6151);
or U13189 (N_13189,N_9544,N_10019);
and U13190 (N_13190,N_11669,N_8537);
and U13191 (N_13191,N_8828,N_11116);
xnor U13192 (N_13192,N_8998,N_9973);
xnor U13193 (N_13193,N_11712,N_8070);
and U13194 (N_13194,N_10241,N_10314);
xor U13195 (N_13195,N_11263,N_6174);
xnor U13196 (N_13196,N_6058,N_6352);
or U13197 (N_13197,N_10698,N_9586);
or U13198 (N_13198,N_11140,N_6109);
xnor U13199 (N_13199,N_10237,N_8410);
nor U13200 (N_13200,N_7308,N_11194);
or U13201 (N_13201,N_11469,N_8847);
nor U13202 (N_13202,N_9873,N_11583);
nand U13203 (N_13203,N_9250,N_9087);
and U13204 (N_13204,N_6647,N_10075);
or U13205 (N_13205,N_11467,N_7021);
nand U13206 (N_13206,N_8024,N_11427);
xnor U13207 (N_13207,N_7019,N_6744);
nand U13208 (N_13208,N_8309,N_7234);
nand U13209 (N_13209,N_9552,N_6788);
and U13210 (N_13210,N_8155,N_11165);
xnor U13211 (N_13211,N_9574,N_10703);
xnor U13212 (N_13212,N_10624,N_10306);
nor U13213 (N_13213,N_6949,N_11759);
xor U13214 (N_13214,N_6351,N_8412);
and U13215 (N_13215,N_9577,N_9917);
nor U13216 (N_13216,N_11599,N_11068);
or U13217 (N_13217,N_9751,N_6627);
nor U13218 (N_13218,N_8844,N_11597);
nor U13219 (N_13219,N_10641,N_9020);
nand U13220 (N_13220,N_6690,N_6279);
xor U13221 (N_13221,N_6630,N_10329);
nand U13222 (N_13222,N_10071,N_6749);
nand U13223 (N_13223,N_11855,N_6569);
nand U13224 (N_13224,N_9103,N_9423);
xnor U13225 (N_13225,N_6743,N_9642);
nor U13226 (N_13226,N_11212,N_11353);
nand U13227 (N_13227,N_10782,N_7197);
or U13228 (N_13228,N_10438,N_7975);
nor U13229 (N_13229,N_9047,N_11749);
nor U13230 (N_13230,N_6551,N_7546);
or U13231 (N_13231,N_7480,N_6194);
xnor U13232 (N_13232,N_11494,N_10155);
xnor U13233 (N_13233,N_6994,N_8889);
nor U13234 (N_13234,N_8016,N_9441);
xnor U13235 (N_13235,N_6265,N_7414);
xor U13236 (N_13236,N_6766,N_7362);
nand U13237 (N_13237,N_7596,N_7543);
and U13238 (N_13238,N_10955,N_9651);
and U13239 (N_13239,N_9380,N_6296);
nor U13240 (N_13240,N_9756,N_10094);
nor U13241 (N_13241,N_11779,N_6934);
or U13242 (N_13242,N_7710,N_7931);
or U13243 (N_13243,N_10745,N_6504);
nor U13244 (N_13244,N_6209,N_11884);
xor U13245 (N_13245,N_8222,N_9442);
and U13246 (N_13246,N_11550,N_9867);
or U13247 (N_13247,N_6491,N_9738);
xnor U13248 (N_13248,N_6270,N_6712);
nand U13249 (N_13249,N_9634,N_11731);
nand U13250 (N_13250,N_9744,N_11362);
or U13251 (N_13251,N_9665,N_7766);
or U13252 (N_13252,N_9998,N_8879);
or U13253 (N_13253,N_9769,N_7360);
nor U13254 (N_13254,N_10949,N_10142);
xnor U13255 (N_13255,N_9073,N_9568);
nor U13256 (N_13256,N_9314,N_8812);
or U13257 (N_13257,N_8358,N_9857);
nor U13258 (N_13258,N_9916,N_8058);
xnor U13259 (N_13259,N_7510,N_7741);
nor U13260 (N_13260,N_9389,N_9063);
nand U13261 (N_13261,N_6287,N_11046);
or U13262 (N_13262,N_11865,N_11822);
nor U13263 (N_13263,N_8613,N_7929);
nand U13264 (N_13264,N_7964,N_6494);
xnor U13265 (N_13265,N_8425,N_7819);
and U13266 (N_13266,N_9473,N_9529);
nand U13267 (N_13267,N_10115,N_11457);
nor U13268 (N_13268,N_6280,N_10331);
or U13269 (N_13269,N_9771,N_10264);
or U13270 (N_13270,N_7218,N_7066);
xor U13271 (N_13271,N_10710,N_10267);
nand U13272 (N_13272,N_6034,N_7473);
and U13273 (N_13273,N_11695,N_11497);
and U13274 (N_13274,N_7186,N_8090);
and U13275 (N_13275,N_11517,N_8884);
xnor U13276 (N_13276,N_7780,N_7336);
xnor U13277 (N_13277,N_9045,N_8326);
or U13278 (N_13278,N_11709,N_8948);
xor U13279 (N_13279,N_9142,N_7206);
nand U13280 (N_13280,N_6740,N_7102);
nand U13281 (N_13281,N_8277,N_7539);
nor U13282 (N_13282,N_11682,N_6933);
xor U13283 (N_13283,N_11689,N_7852);
and U13284 (N_13284,N_6831,N_10586);
and U13285 (N_13285,N_8140,N_10501);
and U13286 (N_13286,N_10622,N_11957);
and U13287 (N_13287,N_11803,N_6208);
xor U13288 (N_13288,N_9677,N_9312);
and U13289 (N_13289,N_11436,N_7699);
nand U13290 (N_13290,N_8699,N_6404);
and U13291 (N_13291,N_6774,N_9510);
nand U13292 (N_13292,N_10969,N_11741);
or U13293 (N_13293,N_6993,N_9720);
nand U13294 (N_13294,N_7915,N_11761);
nor U13295 (N_13295,N_7660,N_10153);
nor U13296 (N_13296,N_7743,N_10653);
and U13297 (N_13297,N_8182,N_11632);
xnor U13298 (N_13298,N_7564,N_6861);
xnor U13299 (N_13299,N_8035,N_7895);
xnor U13300 (N_13300,N_6875,N_9882);
or U13301 (N_13301,N_8818,N_9516);
or U13302 (N_13302,N_6979,N_6539);
nand U13303 (N_13303,N_7889,N_10076);
xnor U13304 (N_13304,N_11463,N_11788);
nand U13305 (N_13305,N_9780,N_6039);
nand U13306 (N_13306,N_9418,N_11657);
nor U13307 (N_13307,N_9041,N_9001);
xor U13308 (N_13308,N_7963,N_11721);
or U13309 (N_13309,N_11753,N_8152);
xor U13310 (N_13310,N_7293,N_11621);
xnor U13311 (N_13311,N_8416,N_11280);
xor U13312 (N_13312,N_6237,N_10968);
or U13313 (N_13313,N_8419,N_6571);
and U13314 (N_13314,N_8595,N_11853);
and U13315 (N_13315,N_8929,N_9427);
and U13316 (N_13316,N_9280,N_9686);
nor U13317 (N_13317,N_6057,N_7331);
and U13318 (N_13318,N_6164,N_10247);
nor U13319 (N_13319,N_9763,N_11573);
or U13320 (N_13320,N_9483,N_9309);
and U13321 (N_13321,N_6447,N_11146);
nand U13322 (N_13322,N_8290,N_9956);
xor U13323 (N_13323,N_10101,N_11365);
and U13324 (N_13324,N_11790,N_8885);
nand U13325 (N_13325,N_9460,N_11147);
nor U13326 (N_13326,N_6342,N_7690);
nand U13327 (N_13327,N_9629,N_10037);
nor U13328 (N_13328,N_9232,N_9252);
nand U13329 (N_13329,N_11180,N_8845);
or U13330 (N_13330,N_7261,N_10816);
and U13331 (N_13331,N_7354,N_10734);
nor U13332 (N_13332,N_6214,N_7862);
and U13333 (N_13333,N_7167,N_6258);
nor U13334 (N_13334,N_7775,N_10841);
or U13335 (N_13335,N_9852,N_11117);
xnor U13336 (N_13336,N_8809,N_7649);
and U13337 (N_13337,N_9907,N_8430);
xnor U13338 (N_13338,N_8496,N_9746);
and U13339 (N_13339,N_11924,N_11400);
nand U13340 (N_13340,N_7909,N_7576);
nor U13341 (N_13341,N_10539,N_8946);
nand U13342 (N_13342,N_6777,N_9182);
nand U13343 (N_13343,N_10635,N_9925);
and U13344 (N_13344,N_10550,N_9202);
nor U13345 (N_13345,N_6437,N_10533);
and U13346 (N_13346,N_10805,N_9631);
nor U13347 (N_13347,N_6513,N_10389);
xnor U13348 (N_13348,N_7676,N_9871);
or U13349 (N_13349,N_9194,N_9589);
xnor U13350 (N_13350,N_7258,N_9582);
and U13351 (N_13351,N_8007,N_7977);
nand U13352 (N_13352,N_8206,N_6033);
nor U13353 (N_13353,N_7008,N_6327);
or U13354 (N_13354,N_7274,N_6368);
xnor U13355 (N_13355,N_9784,N_11526);
xnor U13356 (N_13356,N_9600,N_11025);
and U13357 (N_13357,N_7061,N_11321);
nor U13358 (N_13358,N_11812,N_9709);
nand U13359 (N_13359,N_9979,N_8447);
nand U13360 (N_13360,N_11723,N_11206);
xor U13361 (N_13361,N_6755,N_6786);
xnor U13362 (N_13362,N_6821,N_11267);
xor U13363 (N_13363,N_11690,N_7334);
and U13364 (N_13364,N_6696,N_7599);
nor U13365 (N_13365,N_8580,N_7685);
xnor U13366 (N_13366,N_6066,N_11654);
or U13367 (N_13367,N_6692,N_6090);
xor U13368 (N_13368,N_11814,N_10053);
or U13369 (N_13369,N_9610,N_7035);
or U13370 (N_13370,N_11024,N_6052);
xor U13371 (N_13371,N_9325,N_6213);
or U13372 (N_13372,N_9411,N_10655);
xnor U13373 (N_13373,N_6846,N_8166);
and U13374 (N_13374,N_8785,N_8336);
nor U13375 (N_13375,N_8584,N_8220);
or U13376 (N_13376,N_8652,N_11445);
nor U13377 (N_13377,N_8688,N_11143);
or U13378 (N_13378,N_6946,N_10426);
or U13379 (N_13379,N_10854,N_10262);
and U13380 (N_13380,N_8187,N_11047);
xnor U13381 (N_13381,N_10612,N_7366);
nand U13382 (N_13382,N_7961,N_8408);
nand U13383 (N_13383,N_9188,N_10040);
xor U13384 (N_13384,N_10487,N_10192);
or U13385 (N_13385,N_10820,N_9096);
and U13386 (N_13386,N_6768,N_11002);
xor U13387 (N_13387,N_7388,N_10498);
or U13388 (N_13388,N_9750,N_6388);
and U13389 (N_13389,N_7634,N_7034);
and U13390 (N_13390,N_8819,N_9227);
nor U13391 (N_13391,N_9455,N_6320);
nor U13392 (N_13392,N_9090,N_8201);
nand U13393 (N_13393,N_9598,N_6908);
or U13394 (N_13394,N_9539,N_8305);
nor U13395 (N_13395,N_8020,N_6926);
or U13396 (N_13396,N_9805,N_9005);
nand U13397 (N_13397,N_6005,N_11931);
or U13398 (N_13398,N_6335,N_6225);
xnor U13399 (N_13399,N_11230,N_11509);
nor U13400 (N_13400,N_7682,N_7237);
nand U13401 (N_13401,N_10896,N_7517);
or U13402 (N_13402,N_9789,N_7103);
and U13403 (N_13403,N_8139,N_6317);
xnor U13404 (N_13404,N_7367,N_11203);
xor U13405 (N_13405,N_7029,N_9253);
and U13406 (N_13406,N_9678,N_6193);
and U13407 (N_13407,N_9939,N_7089);
and U13408 (N_13408,N_7668,N_9382);
nor U13409 (N_13409,N_11495,N_10118);
nor U13410 (N_13410,N_7772,N_6582);
xnor U13411 (N_13411,N_9522,N_6793);
or U13412 (N_13412,N_8749,N_6527);
and U13413 (N_13413,N_11933,N_9440);
or U13414 (N_13414,N_10743,N_9030);
nor U13415 (N_13415,N_7806,N_6073);
and U13416 (N_13416,N_6852,N_6746);
and U13417 (N_13417,N_8321,N_8970);
nor U13418 (N_13418,N_8153,N_8029);
or U13419 (N_13419,N_8103,N_11559);
and U13420 (N_13420,N_8063,N_8003);
nand U13421 (N_13421,N_9136,N_10017);
nor U13422 (N_13422,N_6640,N_8089);
nor U13423 (N_13423,N_10401,N_9017);
xor U13424 (N_13424,N_6238,N_9823);
nand U13425 (N_13425,N_7533,N_9513);
and U13426 (N_13426,N_6985,N_7648);
xnor U13427 (N_13427,N_6843,N_7001);
xor U13428 (N_13428,N_7538,N_11426);
xnor U13429 (N_13429,N_9572,N_9691);
or U13430 (N_13430,N_8314,N_7379);
nor U13431 (N_13431,N_9804,N_10125);
or U13432 (N_13432,N_11591,N_9517);
xor U13433 (N_13433,N_9659,N_6989);
and U13434 (N_13434,N_6243,N_8115);
xor U13435 (N_13435,N_7908,N_8637);
and U13436 (N_13436,N_11360,N_9778);
xor U13437 (N_13437,N_9369,N_8031);
and U13438 (N_13438,N_7590,N_9994);
xnor U13439 (N_13439,N_7178,N_10083);
and U13440 (N_13440,N_9131,N_6189);
nor U13441 (N_13441,N_8235,N_7727);
or U13442 (N_13442,N_8805,N_9221);
or U13443 (N_13443,N_7579,N_7922);
and U13444 (N_13444,N_9597,N_11398);
or U13445 (N_13445,N_7937,N_10009);
xnor U13446 (N_13446,N_7561,N_8160);
xnor U13447 (N_13447,N_8861,N_7781);
and U13448 (N_13448,N_11625,N_9176);
xnor U13449 (N_13449,N_7647,N_6860);
and U13450 (N_13450,N_10228,N_7902);
nor U13451 (N_13451,N_9100,N_8722);
nor U13452 (N_13452,N_6567,N_6835);
and U13453 (N_13453,N_10981,N_6273);
xor U13454 (N_13454,N_9323,N_9313);
nor U13455 (N_13455,N_6377,N_6542);
nor U13456 (N_13456,N_8692,N_10863);
nor U13457 (N_13457,N_11551,N_8399);
or U13458 (N_13458,N_9394,N_6376);
nor U13459 (N_13459,N_8504,N_7385);
or U13460 (N_13460,N_10023,N_6910);
xnor U13461 (N_13461,N_6059,N_11900);
or U13462 (N_13462,N_10797,N_8903);
nand U13463 (N_13463,N_9417,N_9371);
nand U13464 (N_13464,N_10584,N_10093);
or U13465 (N_13465,N_11243,N_8370);
or U13466 (N_13466,N_10480,N_6975);
xor U13467 (N_13467,N_6415,N_10156);
nand U13468 (N_13468,N_8980,N_9459);
nor U13469 (N_13469,N_8017,N_6277);
nand U13470 (N_13470,N_11801,N_11874);
or U13471 (N_13471,N_9214,N_11221);
xor U13472 (N_13472,N_6590,N_9456);
nand U13473 (N_13473,N_9121,N_6589);
or U13474 (N_13474,N_10462,N_8621);
nor U13475 (N_13475,N_7586,N_10907);
xor U13476 (N_13476,N_11729,N_10785);
nor U13477 (N_13477,N_9068,N_8348);
or U13478 (N_13478,N_10191,N_7003);
or U13479 (N_13479,N_8859,N_9698);
or U13480 (N_13480,N_11636,N_7597);
nand U13481 (N_13481,N_7592,N_6115);
xor U13482 (N_13482,N_8769,N_10875);
or U13483 (N_13483,N_9854,N_9431);
and U13484 (N_13484,N_7048,N_11001);
or U13485 (N_13485,N_9364,N_7423);
nand U13486 (N_13486,N_11082,N_6091);
nand U13487 (N_13487,N_7955,N_9726);
and U13488 (N_13488,N_6130,N_7542);
or U13489 (N_13489,N_8593,N_10111);
xnor U13490 (N_13490,N_7335,N_10320);
and U13491 (N_13491,N_8558,N_6697);
nor U13492 (N_13492,N_11211,N_10705);
nand U13493 (N_13493,N_10689,N_9658);
nor U13494 (N_13494,N_8520,N_9315);
nand U13495 (N_13495,N_7007,N_10250);
nor U13496 (N_13496,N_10291,N_8353);
nand U13497 (N_13497,N_11679,N_6332);
nor U13498 (N_13498,N_11441,N_6029);
xor U13499 (N_13499,N_10707,N_10351);
nand U13500 (N_13500,N_11090,N_10447);
and U13501 (N_13501,N_6629,N_11648);
nand U13502 (N_13502,N_8726,N_8254);
or U13503 (N_13503,N_9653,N_10319);
nor U13504 (N_13504,N_10563,N_7598);
xor U13505 (N_13505,N_7633,N_6157);
nand U13506 (N_13506,N_7905,N_7487);
and U13507 (N_13507,N_10606,N_8424);
nor U13508 (N_13508,N_11085,N_8083);
xor U13509 (N_13509,N_6155,N_8782);
nor U13510 (N_13510,N_8095,N_6252);
and U13511 (N_13511,N_8759,N_8512);
and U13512 (N_13512,N_7557,N_7081);
and U13513 (N_13513,N_9856,N_9888);
xnor U13514 (N_13514,N_6260,N_10107);
nor U13515 (N_13515,N_6310,N_9915);
or U13516 (N_13516,N_7529,N_11560);
xnor U13517 (N_13517,N_6468,N_9098);
xor U13518 (N_13518,N_8128,N_7479);
or U13519 (N_13519,N_9611,N_9363);
nand U13520 (N_13520,N_8107,N_6291);
nand U13521 (N_13521,N_6222,N_8530);
xor U13522 (N_13522,N_10730,N_9550);
xnor U13523 (N_13523,N_7092,N_6502);
and U13524 (N_13524,N_10022,N_10910);
xnor U13525 (N_13525,N_9990,N_10256);
xor U13526 (N_13526,N_11155,N_8821);
and U13527 (N_13527,N_7653,N_10025);
or U13528 (N_13528,N_10788,N_6776);
and U13529 (N_13529,N_9425,N_7930);
nand U13530 (N_13530,N_8563,N_10227);
xor U13531 (N_13531,N_7127,N_6054);
xnor U13532 (N_13532,N_8575,N_7325);
xnor U13533 (N_13533,N_7498,N_6244);
or U13534 (N_13534,N_9322,N_10834);
nand U13535 (N_13535,N_8397,N_10890);
nand U13536 (N_13536,N_9782,N_11334);
nor U13537 (N_13537,N_11242,N_9204);
and U13538 (N_13538,N_11198,N_7470);
or U13539 (N_13539,N_6631,N_11785);
or U13540 (N_13540,N_8092,N_9452);
or U13541 (N_13541,N_11201,N_7254);
nor U13542 (N_13542,N_7630,N_10430);
nand U13543 (N_13543,N_9044,N_6469);
or U13544 (N_13544,N_11711,N_9601);
or U13545 (N_13545,N_9302,N_10323);
nor U13546 (N_13546,N_8264,N_8731);
xnor U13547 (N_13547,N_10976,N_8908);
xnor U13548 (N_13548,N_6016,N_10050);
nor U13549 (N_13549,N_7078,N_11171);
and U13550 (N_13550,N_8441,N_8218);
or U13551 (N_13551,N_6633,N_10407);
nand U13552 (N_13552,N_9160,N_10590);
and U13553 (N_13553,N_9169,N_10307);
nand U13554 (N_13554,N_9155,N_7125);
or U13555 (N_13555,N_10481,N_10778);
and U13556 (N_13556,N_8647,N_7275);
xor U13557 (N_13557,N_6192,N_7591);
xor U13558 (N_13558,N_7983,N_10593);
xnor U13559 (N_13559,N_8693,N_9195);
and U13560 (N_13560,N_10947,N_8661);
nand U13561 (N_13561,N_8546,N_7410);
nor U13562 (N_13562,N_6184,N_10528);
or U13563 (N_13563,N_7243,N_10171);
xnor U13564 (N_13564,N_10029,N_10208);
and U13565 (N_13565,N_10217,N_6247);
nor U13566 (N_13566,N_8366,N_9624);
nand U13567 (N_13567,N_7848,N_6383);
and U13568 (N_13568,N_7469,N_9694);
nand U13569 (N_13569,N_6173,N_8849);
and U13570 (N_13570,N_7876,N_10495);
nor U13571 (N_13571,N_8125,N_11714);
nand U13572 (N_13572,N_11592,N_6618);
or U13573 (N_13573,N_11697,N_11142);
xor U13574 (N_13574,N_10795,N_10889);
and U13575 (N_13575,N_7233,N_6466);
nand U13576 (N_13576,N_10296,N_10694);
xor U13577 (N_13577,N_9567,N_8158);
and U13578 (N_13578,N_7565,N_8631);
nor U13579 (N_13579,N_6826,N_11049);
xnor U13580 (N_13580,N_6424,N_6146);
nand U13581 (N_13581,N_6043,N_7606);
xnor U13582 (N_13582,N_8507,N_7845);
xor U13583 (N_13583,N_11246,N_7153);
and U13584 (N_13584,N_6659,N_11934);
or U13585 (N_13585,N_11782,N_8581);
and U13586 (N_13586,N_6232,N_11484);
or U13587 (N_13587,N_8841,N_9662);
nand U13588 (N_13588,N_10010,N_10163);
nand U13589 (N_13589,N_11569,N_10908);
or U13590 (N_13590,N_10223,N_10571);
xor U13591 (N_13591,N_10347,N_10309);
nand U13592 (N_13592,N_11237,N_9374);
xor U13593 (N_13593,N_10814,N_7622);
nand U13594 (N_13594,N_9569,N_8748);
or U13595 (N_13595,N_10473,N_11219);
nor U13596 (N_13596,N_6370,N_9351);
nand U13597 (N_13597,N_8572,N_9526);
and U13598 (N_13598,N_9141,N_8969);
nor U13599 (N_13599,N_8117,N_8490);
or U13600 (N_13600,N_10823,N_10918);
xnor U13601 (N_13601,N_8795,N_6031);
nand U13602 (N_13602,N_8009,N_10204);
xnor U13603 (N_13603,N_6942,N_11213);
nor U13604 (N_13604,N_11860,N_10380);
nand U13605 (N_13605,N_6856,N_7262);
nor U13606 (N_13606,N_10148,N_9445);
or U13607 (N_13607,N_11813,N_7203);
xnor U13608 (N_13608,N_6718,N_10278);
xnor U13609 (N_13609,N_6026,N_9657);
or U13610 (N_13610,N_10034,N_8648);
or U13611 (N_13611,N_9097,N_11474);
and U13612 (N_13612,N_8418,N_8258);
nor U13613 (N_13613,N_8720,N_6700);
nor U13614 (N_13614,N_10564,N_11483);
and U13615 (N_13615,N_9326,N_9874);
nand U13616 (N_13616,N_6734,N_7855);
nor U13617 (N_13617,N_10144,N_11061);
or U13618 (N_13618,N_11653,N_10201);
nand U13619 (N_13619,N_6436,N_7319);
or U13620 (N_13620,N_10178,N_6584);
or U13621 (N_13621,N_7742,N_11011);
nand U13622 (N_13622,N_7012,N_8289);
and U13623 (N_13623,N_6156,N_11433);
xor U13624 (N_13624,N_10971,N_7992);
nand U13625 (N_13625,N_10215,N_6325);
nand U13626 (N_13626,N_8877,N_9463);
and U13627 (N_13627,N_10098,N_7016);
nor U13628 (N_13628,N_10066,N_9963);
or U13629 (N_13629,N_8655,N_6679);
nand U13630 (N_13630,N_9305,N_7475);
nand U13631 (N_13631,N_8104,N_6829);
and U13632 (N_13632,N_6175,N_10800);
nor U13633 (N_13633,N_10337,N_8790);
nand U13634 (N_13634,N_10506,N_7488);
nor U13635 (N_13635,N_10437,N_6350);
nand U13636 (N_13636,N_10942,N_8378);
xor U13637 (N_13637,N_11546,N_11369);
nor U13638 (N_13638,N_7286,N_7640);
and U13639 (N_13639,N_11910,N_8723);
nor U13640 (N_13640,N_8915,N_10546);
nor U13641 (N_13641,N_11195,N_11239);
nand U13642 (N_13642,N_8612,N_8011);
and U13643 (N_13643,N_8984,N_10679);
or U13644 (N_13644,N_8590,N_7158);
nor U13645 (N_13645,N_6449,N_11563);
or U13646 (N_13646,N_8250,N_11000);
nand U13647 (N_13647,N_9077,N_8192);
or U13648 (N_13648,N_7946,N_10972);
nand U13649 (N_13649,N_11955,N_11274);
nand U13650 (N_13650,N_10830,N_8974);
or U13651 (N_13651,N_8977,N_10077);
xnor U13652 (N_13652,N_8573,N_8605);
and U13653 (N_13653,N_7667,N_6220);
xnor U13654 (N_13654,N_11502,N_6869);
or U13655 (N_13655,N_7223,N_8343);
xor U13656 (N_13656,N_10860,N_6116);
nor U13657 (N_13657,N_6074,N_11131);
nor U13658 (N_13658,N_10657,N_10195);
nand U13659 (N_13659,N_8091,N_8142);
and U13660 (N_13660,N_11208,N_8059);
and U13661 (N_13661,N_6691,N_8098);
and U13662 (N_13662,N_8004,N_7521);
and U13663 (N_13663,N_11630,N_8803);
or U13664 (N_13664,N_8564,N_7159);
and U13665 (N_13665,N_10806,N_6229);
or U13666 (N_13666,N_8491,N_8495);
nor U13667 (N_13667,N_10285,N_9475);
nor U13668 (N_13668,N_10940,N_11181);
xnor U13669 (N_13669,N_10840,N_7183);
or U13670 (N_13670,N_8941,N_7989);
xnor U13671 (N_13671,N_11375,N_6714);
nor U13672 (N_13672,N_9955,N_11646);
xnor U13673 (N_13673,N_6602,N_8226);
nor U13674 (N_13674,N_8138,N_6044);
nand U13675 (N_13675,N_11443,N_7758);
or U13676 (N_13676,N_8461,N_7289);
nor U13677 (N_13677,N_10308,N_10230);
or U13678 (N_13678,N_8460,N_9000);
nand U13679 (N_13679,N_7684,N_11945);
nor U13680 (N_13680,N_8913,N_8079);
nand U13681 (N_13681,N_8683,N_6892);
nor U13682 (N_13682,N_9999,N_11370);
nor U13683 (N_13683,N_6515,N_8665);
and U13684 (N_13684,N_9162,N_8463);
or U13685 (N_13685,N_10915,N_11215);
or U13686 (N_13686,N_10421,N_11167);
or U13687 (N_13687,N_7794,N_11988);
and U13688 (N_13688,N_7933,N_7841);
nor U13689 (N_13689,N_6806,N_11557);
or U13690 (N_13690,N_10852,N_7309);
xnor U13691 (N_13691,N_10662,N_9530);
and U13692 (N_13692,N_10365,N_10517);
or U13693 (N_13693,N_7798,N_8429);
nand U13694 (N_13694,N_11088,N_9548);
or U13695 (N_13695,N_9948,N_11245);
nand U13696 (N_13696,N_9373,N_9491);
nand U13697 (N_13697,N_7792,N_6686);
nor U13698 (N_13698,N_11343,N_10096);
xor U13699 (N_13699,N_11651,N_6144);
nand U13700 (N_13700,N_11179,N_10318);
nor U13701 (N_13701,N_7729,N_8882);
nand U13702 (N_13702,N_7839,N_10444);
xnor U13703 (N_13703,N_9944,N_6524);
nor U13704 (N_13704,N_8077,N_7679);
xnor U13705 (N_13705,N_11293,N_11456);
nor U13706 (N_13706,N_9727,N_6601);
xor U13707 (N_13707,N_7050,N_11233);
xnor U13708 (N_13708,N_6441,N_8143);
or U13709 (N_13709,N_7291,N_7244);
or U13710 (N_13710,N_11437,N_11827);
xor U13711 (N_13711,N_10560,N_6011);
nand U13712 (N_13712,N_8880,N_8468);
xnor U13713 (N_13713,N_10880,N_6616);
nand U13714 (N_13714,N_7950,N_7617);
nor U13715 (N_13715,N_7370,N_7407);
nand U13716 (N_13716,N_11773,N_8469);
nand U13717 (N_13717,N_9422,N_8958);
nor U13718 (N_13718,N_7142,N_10212);
or U13719 (N_13719,N_8216,N_11337);
nor U13720 (N_13720,N_8820,N_7613);
nand U13721 (N_13721,N_10360,N_8628);
and U13722 (N_13722,N_10739,N_9880);
or U13723 (N_13723,N_11567,N_8991);
nor U13724 (N_13724,N_10953,N_10253);
nand U13725 (N_13725,N_11791,N_10280);
xor U13726 (N_13726,N_6830,N_6931);
nand U13727 (N_13727,N_10079,N_6257);
xnor U13728 (N_13728,N_6470,N_6538);
nand U13729 (N_13729,N_9615,N_11826);
nand U13730 (N_13730,N_11702,N_10682);
or U13731 (N_13731,N_11040,N_6346);
nor U13732 (N_13732,N_9432,N_7865);
or U13733 (N_13733,N_6295,N_11496);
nand U13734 (N_13734,N_8021,N_8231);
and U13735 (N_13735,N_11652,N_10123);
nor U13736 (N_13736,N_8854,N_6172);
or U13737 (N_13737,N_7108,N_9062);
and U13738 (N_13738,N_11162,N_10136);
xnor U13739 (N_13739,N_9387,N_9801);
and U13740 (N_13740,N_10897,N_10372);
or U13741 (N_13741,N_11633,N_10963);
nor U13742 (N_13742,N_11144,N_11707);
or U13743 (N_13743,N_11410,N_9992);
xnor U13744 (N_13744,N_11554,N_6150);
nand U13745 (N_13745,N_11095,N_7084);
or U13746 (N_13746,N_9549,N_8636);
and U13747 (N_13747,N_11223,N_10026);
nand U13748 (N_13748,N_8751,N_11238);
and U13749 (N_13749,N_8905,N_8779);
nor U13750 (N_13750,N_6337,N_11615);
nor U13751 (N_13751,N_11260,N_11435);
nor U13752 (N_13752,N_9201,N_7560);
nor U13753 (N_13753,N_6575,N_6430);
nand U13754 (N_13754,N_6465,N_9708);
nand U13755 (N_13755,N_6655,N_7958);
nor U13756 (N_13756,N_8244,N_8851);
and U13757 (N_13757,N_7313,N_8529);
or U13758 (N_13758,N_9619,N_8526);
nand U13759 (N_13759,N_10475,N_8036);
nand U13760 (N_13760,N_6266,N_8332);
xor U13761 (N_13761,N_11645,N_8119);
nor U13762 (N_13762,N_7515,N_10695);
nand U13763 (N_13763,N_10036,N_8863);
nand U13764 (N_13764,N_7803,N_7745);
nor U13765 (N_13765,N_6384,N_8315);
xor U13766 (N_13766,N_9078,N_6363);
or U13767 (N_13767,N_11582,N_8516);
nor U13768 (N_13768,N_8561,N_6188);
nor U13769 (N_13769,N_10557,N_8794);
nor U13770 (N_13770,N_6212,N_8275);
nand U13771 (N_13771,N_6302,N_7508);
xor U13772 (N_13772,N_8540,N_10775);
nor U13773 (N_13773,N_6205,N_11037);
xnor U13774 (N_13774,N_8764,N_9716);
and U13775 (N_13775,N_10809,N_7418);
or U13776 (N_13776,N_7826,N_6268);
or U13777 (N_13777,N_11704,N_9173);
nand U13778 (N_13778,N_7312,N_7200);
and U13779 (N_13779,N_7846,N_9383);
and U13780 (N_13780,N_10543,N_10794);
nand U13781 (N_13781,N_7618,N_8550);
xnor U13782 (N_13782,N_8279,N_11164);
and U13783 (N_13783,N_8716,N_8638);
xor U13784 (N_13784,N_8144,N_9392);
and U13785 (N_13785,N_11972,N_6501);
xor U13786 (N_13786,N_11544,N_7085);
nand U13787 (N_13787,N_6984,N_10583);
nor U13788 (N_13788,N_7420,N_10673);
and U13789 (N_13789,N_9467,N_7936);
nand U13790 (N_13790,N_8808,N_11482);
nor U13791 (N_13791,N_9911,N_8437);
nor U13792 (N_13792,N_8767,N_10787);
xor U13793 (N_13793,N_9580,N_11083);
and U13794 (N_13794,N_8294,N_10503);
xnor U13795 (N_13795,N_11307,N_11824);
nand U13796 (N_13796,N_9010,N_9566);
or U13797 (N_13797,N_6179,N_10873);
nand U13798 (N_13798,N_10669,N_8267);
and U13799 (N_13799,N_8306,N_8576);
nor U13800 (N_13800,N_10140,N_6186);
or U13801 (N_13801,N_10082,N_6341);
or U13802 (N_13802,N_7913,N_11929);
or U13803 (N_13803,N_9082,N_11232);
nand U13804 (N_13804,N_7939,N_6961);
or U13805 (N_13805,N_10394,N_8363);
or U13806 (N_13806,N_6877,N_10055);
nand U13807 (N_13807,N_6580,N_11408);
or U13808 (N_13808,N_10018,N_8582);
xor U13809 (N_13809,N_6018,N_11656);
xor U13810 (N_13810,N_8310,N_10311);
nor U13811 (N_13811,N_7424,N_7860);
and U13812 (N_13812,N_9203,N_11847);
nor U13813 (N_13813,N_6783,N_10486);
nor U13814 (N_13814,N_8660,N_9258);
nor U13815 (N_13815,N_10108,N_7568);
xnor U13816 (N_13816,N_6397,N_6107);
xnor U13817 (N_13817,N_11273,N_9623);
and U13818 (N_13818,N_7513,N_11610);
or U13819 (N_13819,N_9026,N_6652);
or U13820 (N_13820,N_10496,N_7149);
and U13821 (N_13821,N_7009,N_9902);
nor U13822 (N_13822,N_6360,N_7603);
xor U13823 (N_13823,N_11941,N_11911);
nor U13824 (N_13824,N_10592,N_7706);
or U13825 (N_13825,N_9286,N_10937);
and U13826 (N_13826,N_11156,N_9702);
or U13827 (N_13827,N_10511,N_11676);
nand U13828 (N_13828,N_9515,N_8614);
nand U13829 (N_13829,N_8643,N_7074);
or U13830 (N_13830,N_9284,N_7330);
nand U13831 (N_13831,N_9814,N_11303);
xor U13832 (N_13832,N_6089,N_6191);
nand U13833 (N_13833,N_8263,N_11659);
xor U13834 (N_13834,N_10530,N_6035);
xnor U13835 (N_13835,N_7454,N_8179);
or U13836 (N_13836,N_9930,N_8571);
nand U13837 (N_13837,N_7226,N_11840);
or U13838 (N_13838,N_6240,N_8727);
and U13839 (N_13839,N_6518,N_11984);
xor U13840 (N_13840,N_9140,N_8640);
and U13841 (N_13841,N_6451,N_11359);
or U13842 (N_13842,N_10060,N_11189);
and U13843 (N_13843,N_9283,N_7390);
nand U13844 (N_13844,N_7747,N_9604);
nor U13845 (N_13845,N_8874,N_9072);
nand U13846 (N_13846,N_9495,N_7872);
nand U13847 (N_13847,N_6945,N_8217);
nand U13848 (N_13848,N_8750,N_9279);
xor U13849 (N_13849,N_7835,N_6141);
or U13850 (N_13850,N_7213,N_7468);
and U13851 (N_13851,N_8426,N_6046);
nor U13852 (N_13852,N_8510,N_8634);
nor U13853 (N_13853,N_6359,N_9518);
or U13854 (N_13854,N_6457,N_11578);
and U13855 (N_13855,N_9740,N_6991);
and U13856 (N_13856,N_10452,N_7940);
xor U13857 (N_13857,N_9070,N_11518);
xnor U13858 (N_13858,N_6925,N_8839);
and U13859 (N_13859,N_7310,N_7296);
and U13860 (N_13860,N_6977,N_6098);
or U13861 (N_13861,N_10334,N_9683);
nor U13862 (N_13862,N_9270,N_6967);
nand U13863 (N_13863,N_9468,N_8685);
and U13864 (N_13864,N_7051,N_7222);
nor U13865 (N_13865,N_9166,N_10279);
or U13866 (N_13866,N_10667,N_10926);
or U13867 (N_13867,N_8454,N_11912);
and U13868 (N_13868,N_11434,N_6102);
nand U13869 (N_13869,N_11429,N_7387);
or U13870 (N_13870,N_9942,N_10680);
nor U13871 (N_13871,N_7785,N_9646);
xor U13872 (N_13872,N_11937,N_6887);
and U13873 (N_13873,N_10951,N_6024);
nor U13874 (N_13874,N_11350,N_8515);
xnor U13875 (N_13875,N_10258,N_6227);
or U13876 (N_13876,N_6723,N_9787);
and U13877 (N_13877,N_6228,N_6267);
nor U13878 (N_13878,N_11363,N_7184);
or U13879 (N_13879,N_7384,N_6844);
nor U13880 (N_13880,N_11058,N_9755);
xor U13881 (N_13881,N_7941,N_7433);
xnor U13882 (N_13882,N_8240,N_9991);
xnor U13883 (N_13883,N_6803,N_10886);
and U13884 (N_13884,N_8118,N_10415);
xnor U13885 (N_13885,N_10555,N_7268);
or U13886 (N_13886,N_11756,N_6523);
nand U13887 (N_13887,N_8093,N_9525);
nor U13888 (N_13888,N_6791,N_8215);
or U13889 (N_13889,N_9154,N_8438);
or U13890 (N_13890,N_8236,N_11746);
nand U13891 (N_13891,N_7406,N_6729);
nor U13892 (N_13892,N_11099,N_11154);
and U13893 (N_13893,N_10370,N_10966);
or U13894 (N_13894,N_11843,N_6836);
and U13895 (N_13895,N_10987,N_8608);
or U13896 (N_13896,N_6845,N_6847);
and U13897 (N_13897,N_10902,N_9357);
and U13898 (N_13898,N_7194,N_8501);
nand U13899 (N_13899,N_10091,N_7854);
and U13900 (N_13900,N_9116,N_10718);
xor U13901 (N_13901,N_6742,N_11489);
nand U13902 (N_13902,N_7327,N_10298);
xnor U13903 (N_13903,N_10485,N_10796);
xnor U13904 (N_13904,N_8154,N_10289);
and U13905 (N_13905,N_8357,N_8869);
nand U13906 (N_13906,N_9056,N_9336);
nor U13907 (N_13907,N_10382,N_9786);
nor U13908 (N_13908,N_10581,N_6710);
xor U13909 (N_13909,N_6561,N_10073);
nor U13910 (N_13910,N_10991,N_11396);
or U13911 (N_13911,N_9353,N_6259);
nor U13912 (N_13912,N_7450,N_10436);
and U13913 (N_13913,N_6653,N_7010);
or U13914 (N_13914,N_7811,N_9233);
nor U13915 (N_13915,N_11315,N_6981);
nor U13916 (N_13916,N_10027,N_6378);
nor U13917 (N_13917,N_8506,N_9388);
and U13918 (N_13918,N_7615,N_8921);
nand U13919 (N_13919,N_10826,N_10229);
nand U13920 (N_13920,N_6431,N_7697);
or U13921 (N_13921,N_6520,N_11285);
nand U13922 (N_13922,N_8616,N_9444);
xnor U13923 (N_13923,N_11750,N_8406);
or U13924 (N_13924,N_8075,N_6036);
or U13925 (N_13925,N_8105,N_9576);
and U13926 (N_13926,N_10476,N_11738);
or U13927 (N_13927,N_6823,N_10569);
or U13928 (N_13928,N_8278,N_7581);
nor U13929 (N_13929,N_9386,N_10315);
and U13930 (N_13930,N_6628,N_6495);
xnor U13931 (N_13931,N_8072,N_7626);
xnor U13932 (N_13932,N_8796,N_7022);
or U13933 (N_13933,N_9395,N_9875);
nand U13934 (N_13934,N_9695,N_7892);
and U13935 (N_13935,N_7821,N_10057);
and U13936 (N_13936,N_8255,N_8313);
xnor U13937 (N_13937,N_11892,N_10371);
and U13938 (N_13938,N_10349,N_9055);
nand U13939 (N_13939,N_8784,N_7886);
nor U13940 (N_13940,N_11261,N_8588);
xnor U13941 (N_13941,N_8773,N_11066);
xor U13942 (N_13942,N_9818,N_7490);
or U13943 (N_13943,N_11774,N_8191);
nand U13944 (N_13944,N_9593,N_10497);
nor U13945 (N_13945,N_7748,N_10244);
nor U13946 (N_13946,N_7899,N_10713);
nand U13947 (N_13947,N_8697,N_11949);
or U13948 (N_13948,N_11966,N_9579);
nor U13949 (N_13949,N_9606,N_7216);
and U13950 (N_13950,N_11428,N_9903);
or U13951 (N_13951,N_10386,N_10801);
or U13952 (N_13952,N_6416,N_9843);
or U13953 (N_13953,N_7602,N_8257);
xnor U13954 (N_13954,N_11132,N_9921);
or U13955 (N_13955,N_11342,N_10294);
and U13956 (N_13956,N_6365,N_8733);
nand U13957 (N_13957,N_7594,N_10121);
and U13958 (N_13958,N_10158,N_9106);
xnor U13959 (N_13959,N_9721,N_11796);
nand U13960 (N_13960,N_7857,N_7927);
nor U13961 (N_13961,N_10455,N_6138);
nor U13962 (N_13962,N_9170,N_6069);
and U13963 (N_13963,N_8452,N_10500);
and U13964 (N_13964,N_7352,N_8876);
and U13965 (N_13965,N_9354,N_9274);
xnor U13966 (N_13966,N_8783,N_9647);
nand U13967 (N_13967,N_6765,N_7375);
or U13968 (N_13968,N_6864,N_6340);
nand U13969 (N_13969,N_9397,N_7717);
and U13970 (N_13970,N_11423,N_9158);
xnor U13971 (N_13971,N_9199,N_7355);
and U13972 (N_13972,N_11701,N_11680);
or U13973 (N_13973,N_6651,N_7600);
nand U13974 (N_13974,N_11909,N_7947);
or U13975 (N_13975,N_6025,N_11014);
nor U13976 (N_13976,N_10317,N_10625);
or U13977 (N_13977,N_8776,N_11671);
and U13978 (N_13978,N_11617,N_9728);
and U13979 (N_13979,N_8875,N_10257);
xnor U13980 (N_13980,N_9255,N_9104);
or U13981 (N_13981,N_11639,N_10431);
and U13982 (N_13982,N_7346,N_11618);
and U13983 (N_13983,N_10129,N_9507);
nor U13984 (N_13984,N_6687,N_7209);
xnor U13985 (N_13985,N_8675,N_7988);
or U13986 (N_13986,N_8714,N_6533);
nor U13987 (N_13987,N_10696,N_9788);
or U13988 (N_13988,N_9803,N_6087);
nor U13989 (N_13989,N_8088,N_10642);
nand U13990 (N_13990,N_9697,N_11523);
nand U13991 (N_13991,N_7139,N_7049);
nand U13992 (N_13992,N_8026,N_6666);
nor U13993 (N_13993,N_9914,N_8486);
xor U13994 (N_13994,N_8762,N_8282);
xnor U13995 (N_13995,N_10803,N_10856);
or U13996 (N_13996,N_9890,N_11538);
xnor U13997 (N_13997,N_11078,N_6331);
and U13998 (N_13998,N_11259,N_10932);
xor U13999 (N_13999,N_8836,N_9133);
nor U14000 (N_14000,N_7317,N_7436);
nand U14001 (N_14001,N_9437,N_10958);
nand U14002 (N_14002,N_11606,N_6458);
and U14003 (N_14003,N_10174,N_9620);
and U14004 (N_14004,N_9119,N_10715);
xor U14005 (N_14005,N_8770,N_10219);
nand U14006 (N_14006,N_7926,N_10159);
nor U14007 (N_14007,N_9575,N_6588);
and U14008 (N_14008,N_9652,N_10735);
nand U14009 (N_14009,N_11309,N_7512);
nor U14010 (N_14010,N_11386,N_6145);
or U14011 (N_14011,N_7028,N_8328);
nand U14012 (N_14012,N_11787,N_10878);
nand U14013 (N_14013,N_10113,N_11407);
xor U14014 (N_14014,N_11991,N_10671);
and U14015 (N_14015,N_11106,N_7255);
nor U14016 (N_14016,N_6574,N_11115);
and U14017 (N_14017,N_9260,N_8069);
nor U14018 (N_14018,N_7658,N_11590);
and U14019 (N_14019,N_7837,N_10313);
nand U14020 (N_14020,N_7770,N_10912);
nand U14021 (N_14021,N_8249,N_9016);
xor U14022 (N_14022,N_11706,N_7378);
xnor U14023 (N_14023,N_7569,N_6824);
or U14024 (N_14024,N_6541,N_8401);
xnor U14025 (N_14025,N_11687,N_11940);
nand U14026 (N_14026,N_10427,N_11283);
nor U14027 (N_14027,N_7917,N_11784);
xor U14028 (N_14028,N_6082,N_6684);
nand U14029 (N_14029,N_11638,N_11811);
xor U14030 (N_14030,N_10637,N_7373);
xnor U14031 (N_14031,N_11838,N_10209);
nor U14032 (N_14032,N_11521,N_9360);
and U14033 (N_14033,N_10832,N_11566);
nor U14034 (N_14034,N_11402,N_10392);
nor U14035 (N_14035,N_6488,N_6131);
nor U14036 (N_14036,N_10063,N_9584);
or U14037 (N_14037,N_9608,N_6882);
or U14038 (N_14038,N_7344,N_7163);
or U14039 (N_14039,N_8599,N_6968);
nor U14040 (N_14040,N_9271,N_11008);
nand U14041 (N_14041,N_10939,N_6680);
and U14042 (N_14042,N_7361,N_8768);
xor U14043 (N_14043,N_7880,N_10768);
and U14044 (N_14044,N_8771,N_7017);
and U14045 (N_14045,N_6784,N_9941);
and U14046 (N_14046,N_10591,N_8045);
or U14047 (N_14047,N_7341,N_11018);
nand U14048 (N_14048,N_6888,N_8111);
nand U14049 (N_14049,N_11341,N_10366);
xor U14050 (N_14050,N_9412,N_11328);
and U14051 (N_14051,N_10527,N_9735);
nor U14052 (N_14052,N_9811,N_6735);
and U14053 (N_14053,N_6577,N_8924);
xnor U14054 (N_14054,N_11347,N_11330);
xor U14055 (N_14055,N_8423,N_10784);
xnor U14056 (N_14056,N_8649,N_9163);
nor U14057 (N_14057,N_8014,N_7239);
and U14058 (N_14058,N_7136,N_6048);
xnor U14059 (N_14059,N_10618,N_10001);
or U14060 (N_14060,N_11490,N_8591);
and U14061 (N_14061,N_10024,N_8650);
nand U14062 (N_14062,N_6050,N_9900);
and U14063 (N_14063,N_10357,N_9276);
nand U14064 (N_14064,N_6339,N_6040);
nor U14065 (N_14065,N_7788,N_6009);
or U14066 (N_14066,N_6554,N_7885);
nand U14067 (N_14067,N_9450,N_8081);
and U14068 (N_14068,N_10549,N_7095);
xnor U14069 (N_14069,N_8744,N_9866);
xor U14070 (N_14070,N_7734,N_10061);
and U14071 (N_14071,N_8040,N_7004);
nor U14072 (N_14072,N_8354,N_10944);
or U14073 (N_14073,N_11312,N_11200);
and U14074 (N_14074,N_6859,N_11739);
and U14075 (N_14075,N_9485,N_7735);
nor U14076 (N_14076,N_11529,N_10109);
and U14077 (N_14077,N_8789,N_6720);
and U14078 (N_14078,N_9736,N_11404);
or U14079 (N_14079,N_8193,N_9831);
and U14080 (N_14080,N_11600,N_11553);
nor U14081 (N_14081,N_11297,N_6566);
xnor U14082 (N_14082,N_11296,N_10611);
and U14083 (N_14083,N_10626,N_8112);
nor U14084 (N_14084,N_9094,N_10484);
and U14085 (N_14085,N_7982,N_9838);
and U14086 (N_14086,N_8471,N_10442);
xor U14087 (N_14087,N_6868,N_9299);
nor U14088 (N_14088,N_9640,N_8066);
nor U14089 (N_14089,N_7541,N_10189);
xnor U14090 (N_14090,N_7890,N_8667);
or U14091 (N_14091,N_9676,N_7673);
nor U14092 (N_14092,N_9573,N_8684);
nand U14093 (N_14093,N_11849,N_11277);
nor U14094 (N_14094,N_9447,N_10793);
and U14095 (N_14095,N_11031,N_9132);
nor U14096 (N_14096,N_9551,N_8449);
nor U14097 (N_14097,N_10293,N_6534);
and U14098 (N_14098,N_7188,N_7492);
nor U14099 (N_14099,N_8701,N_10084);
and U14100 (N_14100,N_8662,N_11767);
nor U14101 (N_14101,N_8162,N_7491);
nand U14102 (N_14102,N_9234,N_10150);
nor U14103 (N_14103,N_10541,N_7082);
or U14104 (N_14104,N_7737,N_6042);
xnor U14105 (N_14105,N_8657,N_11895);
xnor U14106 (N_14106,N_9144,N_9564);
and U14107 (N_14107,N_8344,N_6251);
nor U14108 (N_14108,N_6932,N_8987);
xnor U14109 (N_14109,N_6585,N_9632);
nor U14110 (N_14110,N_10776,N_8721);
or U14111 (N_14111,N_7914,N_10251);
nand U14112 (N_14112,N_8303,N_10164);
xor U14113 (N_14113,N_11252,N_11917);
nand U14114 (N_14114,N_7850,N_6898);
and U14115 (N_14115,N_9563,N_8568);
xnor U14116 (N_14116,N_11958,N_6092);
xnor U14117 (N_14117,N_11915,N_6396);
nand U14118 (N_14118,N_9401,N_8012);
nor U14119 (N_14119,N_11980,N_6525);
nand U14120 (N_14120,N_8729,N_7064);
nand U14121 (N_14121,N_11631,N_8080);
nor U14122 (N_14122,N_6484,N_9733);
or U14123 (N_14123,N_8654,N_7953);
and U14124 (N_14124,N_10441,N_8801);
and U14125 (N_14125,N_7843,N_9860);
xnor U14126 (N_14126,N_10565,N_10609);
nor U14127 (N_14127,N_11898,N_8574);
nor U14128 (N_14128,N_9663,N_7147);
nor U14129 (N_14129,N_11364,N_9189);
xor U14130 (N_14130,N_10236,N_9331);
or U14131 (N_14131,N_11781,N_7020);
nand U14132 (N_14132,N_10615,N_10954);
or U14133 (N_14133,N_7232,N_6364);
nor U14134 (N_14134,N_7869,N_6905);
xnor U14135 (N_14135,N_7807,N_9690);
or U14136 (N_14136,N_10686,N_6510);
xor U14137 (N_14137,N_7245,N_11192);
xnor U14138 (N_14138,N_10453,N_8481);
nor U14139 (N_14139,N_7447,N_7763);
or U14140 (N_14140,N_11778,N_7619);
xor U14141 (N_14141,N_10598,N_10207);
nor U14142 (N_14142,N_9265,N_6063);
nand U14143 (N_14143,N_9406,N_9429);
or U14144 (N_14144,N_9807,N_7587);
nor U14145 (N_14145,N_8056,N_8340);
nand U14146 (N_14146,N_8775,N_9905);
nor U14147 (N_14147,N_7558,N_6298);
or U14148 (N_14148,N_6825,N_9091);
and U14149 (N_14149,N_10765,N_11981);
nand U14150 (N_14150,N_11190,N_11447);
nor U14151 (N_14151,N_10181,N_8860);
nor U14152 (N_14152,N_9881,N_7689);
nor U14153 (N_14153,N_11806,N_8364);
nor U14154 (N_14154,N_8705,N_7283);
nand U14155 (N_14155,N_7783,N_7716);
xor U14156 (N_14156,N_10534,N_6795);
nand U14157 (N_14157,N_7896,N_11643);
and U14158 (N_14158,N_6531,N_9668);
nor U14159 (N_14159,N_7032,N_8186);
nor U14160 (N_14160,N_7642,N_10709);
or U14161 (N_14161,N_8799,N_7733);
nor U14162 (N_14162,N_9022,N_7376);
xnor U14163 (N_14163,N_10941,N_8151);
or U14164 (N_14164,N_11549,N_10906);
and U14165 (N_14165,N_11191,N_11118);
nor U14166 (N_14166,N_10358,N_9896);
nor U14167 (N_14167,N_7944,N_9134);
nor U14168 (N_14168,N_11733,N_11835);
or U14169 (N_14169,N_6366,N_10864);
and U14170 (N_14170,N_8421,N_9356);
or U14171 (N_14171,N_10467,N_9481);
and U14172 (N_14172,N_11185,N_6312);
and U14173 (N_14173,N_9731,N_11074);
nor U14174 (N_14174,N_11300,N_10145);
nor U14175 (N_14175,N_8838,N_8734);
nand U14176 (N_14176,N_8225,N_9294);
nor U14177 (N_14177,N_6440,N_6880);
xnor U14178 (N_14178,N_11568,N_8350);
nand U14179 (N_14179,N_8996,N_7641);
or U14180 (N_14180,N_7624,N_8183);
and U14181 (N_14181,N_10770,N_10728);
nand U14182 (N_14182,N_6472,N_11953);
nor U14183 (N_14183,N_8476,N_11019);
and U14184 (N_14184,N_7462,N_10510);
nor U14185 (N_14185,N_8702,N_7662);
nand U14186 (N_14186,N_9884,N_11029);
nand U14187 (N_14187,N_8034,N_10226);
xor U14188 (N_14188,N_7925,N_6432);
nor U14189 (N_14189,N_8129,N_9492);
nor U14190 (N_14190,N_9344,N_9358);
and U14191 (N_14191,N_8163,N_6326);
nand U14192 (N_14192,N_9080,N_11076);
xnor U14193 (N_14193,N_9810,N_7400);
nand U14194 (N_14194,N_8738,N_6886);
and U14195 (N_14195,N_10582,N_11105);
nand U14196 (N_14196,N_10672,N_9213);
nand U14197 (N_14197,N_9069,N_9215);
and U14198 (N_14198,N_10367,N_11882);
or U14199 (N_14199,N_7851,N_7723);
and U14200 (N_14200,N_6586,N_6185);
nand U14201 (N_14201,N_9434,N_10843);
nand U14202 (N_14202,N_11073,N_9842);
and U14203 (N_14203,N_10751,N_11627);
and U14204 (N_14204,N_10047,N_11476);
nand U14205 (N_14205,N_11852,N_8019);
nor U14206 (N_14206,N_6286,N_8620);
and U14207 (N_14207,N_6885,N_6037);
nor U14208 (N_14208,N_7681,N_6180);
nor U14209 (N_14209,N_8131,N_7823);
nand U14210 (N_14210,N_7075,N_8434);
nand U14211 (N_14211,N_10579,N_7966);
nand U14212 (N_14212,N_11565,N_11041);
xor U14213 (N_14213,N_6663,N_7623);
nor U14214 (N_14214,N_9938,N_10202);
and U14215 (N_14215,N_10827,N_10737);
nor U14216 (N_14216,N_10103,N_9799);
or U14217 (N_14217,N_7465,N_11112);
nand U14218 (N_14218,N_11596,N_6622);
nand U14219 (N_14219,N_7738,N_9409);
nor U14220 (N_14220,N_9318,N_11374);
and U14221 (N_14221,N_11067,N_8276);
and U14222 (N_14222,N_11256,N_10008);
nand U14223 (N_14223,N_8265,N_9614);
and U14224 (N_14224,N_7055,N_9654);
or U14225 (N_14225,N_6284,N_6176);
xnor U14226 (N_14226,N_9943,N_10160);
nand U14227 (N_14227,N_8754,N_11103);
and U14228 (N_14228,N_11385,N_8892);
or U14229 (N_14229,N_8978,N_7506);
xor U14230 (N_14230,N_6235,N_11798);
nor U14231 (N_14231,N_9093,N_7405);
nor U14232 (N_14232,N_8583,N_6485);
xor U14233 (N_14233,N_8044,N_9102);
or U14234 (N_14234,N_9649,N_8965);
or U14235 (N_14235,N_10507,N_7372);
or U14236 (N_14236,N_10811,N_7545);
nor U14237 (N_14237,N_9150,N_9230);
and U14238 (N_14238,N_7525,N_10993);
or U14239 (N_14239,N_9970,N_9184);
xnor U14240 (N_14240,N_7110,N_9699);
nor U14241 (N_14241,N_11930,N_11545);
nand U14242 (N_14242,N_10644,N_6313);
xor U14243 (N_14243,N_11016,N_10088);
nand U14244 (N_14244,N_10654,N_10982);
or U14245 (N_14245,N_7870,N_10600);
or U14246 (N_14246,N_8772,N_8732);
nor U14247 (N_14247,N_6169,N_8433);
nor U14248 (N_14248,N_10395,N_11907);
xor U14249 (N_14249,N_11943,N_10273);
or U14250 (N_14250,N_8519,N_6909);
nand U14251 (N_14251,N_6496,N_8619);
nand U14252 (N_14252,N_8368,N_7083);
nor U14253 (N_14253,N_8888,N_6077);
and U14254 (N_14254,N_9027,N_6812);
xor U14255 (N_14255,N_6555,N_7984);
or U14256 (N_14256,N_6159,N_8436);
xor U14257 (N_14257,N_10985,N_11794);
nand U14258 (N_14258,N_10128,N_6928);
or U14259 (N_14259,N_8047,N_8562);
and U14260 (N_14260,N_7951,N_9815);
nand U14261 (N_14261,N_6801,N_7150);
nand U14262 (N_14262,N_8792,N_10621);
and U14263 (N_14263,N_8492,N_6893);
nor U14264 (N_14264,N_6133,N_7443);
nand U14265 (N_14265,N_8508,N_10377);
and U14266 (N_14266,N_11842,N_6474);
nand U14267 (N_14267,N_9545,N_6476);
xnor U14268 (N_14268,N_11241,N_6181);
nor U14269 (N_14269,N_8522,N_6646);
xnor U14270 (N_14270,N_8232,N_9757);
or U14271 (N_14271,N_10872,N_8979);
or U14272 (N_14272,N_6550,N_10702);
nor U14273 (N_14273,N_7404,N_7954);
and U14274 (N_14274,N_10855,N_9372);
and U14275 (N_14275,N_8025,N_7732);
nand U14276 (N_14276,N_8374,N_9859);
nor U14277 (N_14277,N_7580,N_8207);
or U14278 (N_14278,N_6417,N_11604);
or U14279 (N_14279,N_7043,N_8933);
or U14280 (N_14280,N_9498,N_10799);
or U14281 (N_14281,N_10697,N_11742);
xor U14282 (N_14282,N_9306,N_6614);
xor U14283 (N_14283,N_10665,N_7767);
nor U14284 (N_14284,N_11006,N_6528);
nor U14285 (N_14285,N_10210,N_7956);
xor U14286 (N_14286,N_11207,N_6211);
nand U14287 (N_14287,N_6626,N_11754);
and U14288 (N_14288,N_6632,N_9587);
and U14289 (N_14289,N_7090,N_11324);
or U14290 (N_14290,N_9523,N_9266);
or U14291 (N_14291,N_8937,N_7252);
xor U14292 (N_14292,N_8850,N_10324);
xnor U14293 (N_14293,N_8873,N_10773);
nor U14294 (N_14294,N_10752,N_7453);
nor U14295 (N_14295,N_7952,N_11797);
xnor U14296 (N_14296,N_7135,N_7381);
xor U14297 (N_14297,N_7484,N_10032);
xnor U14298 (N_14298,N_6644,N_6099);
xnor U14299 (N_14299,N_7705,N_7445);
nor U14300 (N_14300,N_9926,N_6445);
or U14301 (N_14301,N_8497,N_7140);
or U14302 (N_14302,N_11588,N_7207);
and U14303 (N_14303,N_6084,N_10602);
or U14304 (N_14304,N_6362,N_9950);
or U14305 (N_14305,N_9951,N_8414);
xnor U14306 (N_14306,N_10984,N_10899);
nor U14307 (N_14307,N_6471,N_11107);
nor U14308 (N_14308,N_9945,N_6428);
or U14309 (N_14309,N_9706,N_6660);
nand U14310 (N_14310,N_9269,N_6615);
or U14311 (N_14311,N_8823,N_9922);
nor U14312 (N_14312,N_11547,N_10973);
and U14313 (N_14313,N_8626,N_7817);
or U14314 (N_14314,N_11416,N_9153);
and U14315 (N_14315,N_9352,N_7505);
and U14316 (N_14316,N_8171,N_8272);
nor U14317 (N_14317,N_9385,N_8639);
and U14318 (N_14318,N_10297,N_8455);
nand U14319 (N_14319,N_6110,N_6838);
nor U14320 (N_14320,N_6435,N_7152);
nor U14321 (N_14321,N_6318,N_7046);
xnor U14322 (N_14322,N_9790,N_9110);
and U14323 (N_14323,N_8323,N_6693);
or U14324 (N_14324,N_11305,N_7636);
or U14325 (N_14325,N_6737,N_9791);
nor U14326 (N_14326,N_8499,N_9076);
or U14327 (N_14327,N_9928,N_10538);
or U14328 (N_14328,N_7928,N_11091);
or U14329 (N_14329,N_6987,N_9701);
nor U14330 (N_14330,N_8967,N_7639);
nor U14331 (N_14331,N_10381,N_6990);
nor U14332 (N_14332,N_10755,N_9508);
or U14333 (N_14333,N_8453,N_10243);
or U14334 (N_14334,N_7609,N_8488);
and U14335 (N_14335,N_9304,N_6135);
xor U14336 (N_14336,N_7577,N_8351);
or U14337 (N_14337,N_6334,N_7114);
nand U14338 (N_14338,N_9536,N_10742);
nor U14339 (N_14339,N_7318,N_8995);
or U14340 (N_14340,N_8333,N_7063);
nor U14341 (N_14341,N_10435,N_7556);
and U14342 (N_14342,N_8130,N_8157);
or U14343 (N_14343,N_8513,N_8678);
or U14344 (N_14344,N_8076,N_6546);
and U14345 (N_14345,N_9626,N_11036);
and U14346 (N_14346,N_6799,N_8038);
or U14347 (N_14347,N_10304,N_7528);
nand U14348 (N_14348,N_6198,N_7297);
nand U14349 (N_14349,N_9588,N_8904);
nor U14350 (N_14350,N_6884,N_6068);
xnor U14351 (N_14351,N_8493,N_10934);
nor U14352 (N_14352,N_8372,N_8635);
and U14353 (N_14353,N_6999,N_6858);
nor U14354 (N_14354,N_7123,N_10961);
and U14355 (N_14355,N_7976,N_8319);
nand U14356 (N_14356,N_6937,N_6274);
or U14357 (N_14357,N_8825,N_10894);
and U14358 (N_14358,N_7481,N_10729);
and U14359 (N_14359,N_11017,N_11218);
or U14360 (N_14360,N_10804,N_6072);
nor U14361 (N_14361,N_11275,N_8543);
and U14362 (N_14362,N_10678,N_10900);
and U14363 (N_14363,N_7112,N_7251);
and U14364 (N_14364,N_11440,N_8094);
xnor U14365 (N_14365,N_11532,N_6246);
or U14366 (N_14366,N_9021,N_7496);
and U14367 (N_14367,N_9400,N_10677);
nor U14368 (N_14368,N_8190,N_9147);
nor U14369 (N_14369,N_6505,N_7190);
and U14370 (N_14370,N_7532,N_6902);
xor U14371 (N_14371,N_6438,N_6922);
nor U14372 (N_14372,N_11717,N_10946);
or U14373 (N_14373,N_6564,N_6866);
nand U14374 (N_14374,N_11120,N_8381);
and U14375 (N_14375,N_7157,N_8356);
nand U14376 (N_14376,N_8959,N_11805);
xnor U14377 (N_14377,N_9054,N_11642);
and U14378 (N_14378,N_7616,N_9149);
or U14379 (N_14379,N_9844,N_6916);
or U14380 (N_14380,N_8428,N_10616);
nand U14381 (N_14381,N_8008,N_6426);
nor U14382 (N_14382,N_7664,N_10433);
nor U14383 (N_14383,N_7871,N_8856);
and U14384 (N_14384,N_11969,N_8178);
nor U14385 (N_14385,N_6645,N_9612);
nand U14386 (N_14386,N_9512,N_9858);
and U14387 (N_14387,N_10445,N_6112);
xnor U14388 (N_14388,N_7567,N_9443);
or U14389 (N_14389,N_7076,N_11248);
nand U14390 (N_14390,N_11688,N_9038);
nor U14391 (N_14391,N_11170,N_6442);
xor U14392 (N_14392,N_10002,N_11996);
nand U14393 (N_14393,N_11401,N_9590);
xnor U14394 (N_14394,N_7663,N_7342);
nand U14395 (N_14395,N_8606,N_11100);
and U14396 (N_14396,N_9346,N_11710);
nor U14397 (N_14397,N_10167,N_10117);
and U14398 (N_14398,N_9785,N_6579);
xor U14399 (N_14399,N_11514,N_10661);
or U14400 (N_14400,N_9849,N_8338);
or U14401 (N_14401,N_7288,N_8544);
xor U14402 (N_14402,N_7935,N_6623);
and U14403 (N_14403,N_7040,N_8164);
or U14404 (N_14404,N_7464,N_6477);
xor U14405 (N_14405,N_7799,N_6285);
or U14406 (N_14406,N_11862,N_7654);
nand U14407 (N_14407,N_6254,N_6263);
or U14408 (N_14408,N_6038,N_7509);
xnor U14409 (N_14409,N_8329,N_7425);
or U14410 (N_14410,N_9919,N_11210);
or U14411 (N_14411,N_7441,N_11387);
nor U14412 (N_14412,N_8100,N_9684);
and U14413 (N_14413,N_7718,N_11593);
nand U14414 (N_14414,N_6726,N_9185);
nand U14415 (N_14415,N_9273,N_8256);
nand U14416 (N_14416,N_7133,N_10170);
or U14417 (N_14417,N_9197,N_6530);
xnor U14418 (N_14418,N_9547,N_7520);
nor U14419 (N_14419,N_10326,N_8763);
nand U14420 (N_14420,N_8198,N_11308);
nand U14421 (N_14421,N_9965,N_6762);
or U14422 (N_14422,N_7302,N_6802);
xor U14423 (N_14423,N_10992,N_6780);
nor U14424 (N_14424,N_6423,N_8677);
nand U14425 (N_14425,N_7847,N_8802);
nand U14426 (N_14426,N_9836,N_6958);
xnor U14427 (N_14427,N_6978,N_11947);
nor U14428 (N_14428,N_11272,N_8239);
nand U14429 (N_14429,N_8632,N_7864);
nand U14430 (N_14430,N_10633,N_7460);
and U14431 (N_14431,N_7495,N_10681);
nand U14432 (N_14432,N_7278,N_6638);
xor U14433 (N_14433,N_7731,N_6605);
or U14434 (N_14434,N_11110,N_9493);
and U14435 (N_14435,N_6678,N_8293);
and U14436 (N_14436,N_9696,N_10925);
nand U14437 (N_14437,N_9482,N_11104);
or U14438 (N_14438,N_7824,N_9347);
xnor U14439 (N_14439,N_10051,N_8920);
and U14440 (N_14440,N_6051,N_7202);
xnor U14441 (N_14441,N_10825,N_6462);
and U14442 (N_14442,N_10354,N_11462);
and U14443 (N_14443,N_11830,N_7247);
nand U14444 (N_14444,N_6769,N_8923);
nand U14445 (N_14445,N_11098,N_8055);
nand U14446 (N_14446,N_7740,N_11786);
nand U14447 (N_14447,N_10368,N_9904);
and U14448 (N_14448,N_8532,N_10271);
xnor U14449 (N_14449,N_11480,N_6763);
xor U14450 (N_14450,N_10249,N_10866);
and U14451 (N_14451,N_6113,N_11392);
or U14452 (N_14452,N_7932,N_10660);
or U14453 (N_14453,N_8386,N_11186);
nor U14454 (N_14454,N_11993,N_10643);
and U14455 (N_14455,N_9111,N_11205);
or U14456 (N_14456,N_10744,N_9717);
or U14457 (N_14457,N_11914,N_6840);
nand U14458 (N_14458,N_6264,N_8494);
or U14459 (N_14459,N_6137,N_7644);
nor U14460 (N_14460,N_10628,N_8459);
xor U14461 (N_14461,N_7359,N_8051);
or U14462 (N_14462,N_7201,N_8123);
nor U14463 (N_14463,N_7456,N_8752);
and U14464 (N_14464,N_6028,N_8610);
xnor U14465 (N_14465,N_11810,N_7631);
xor U14466 (N_14466,N_7793,N_9762);
or U14467 (N_14467,N_9399,N_11673);
and U14468 (N_14468,N_6998,N_10095);
or U14469 (N_14469,N_9776,N_11737);
or U14470 (N_14470,N_10483,N_10913);
or U14471 (N_14471,N_7575,N_9361);
nand U14472 (N_14472,N_6202,N_6544);
or U14473 (N_14473,N_7000,N_11022);
xor U14474 (N_14474,N_8413,N_10914);
and U14475 (N_14475,N_11539,N_8185);
and U14476 (N_14476,N_8174,N_7270);
nor U14477 (N_14477,N_6455,N_10780);
xor U14478 (N_14478,N_8346,N_6406);
xor U14479 (N_14479,N_10440,N_7018);
nand U14480 (N_14480,N_6443,N_7281);
and U14481 (N_14481,N_11351,N_8671);
or U14482 (N_14482,N_10977,N_9159);
or U14483 (N_14483,N_7415,N_9596);
nand U14484 (N_14484,N_8942,N_8023);
nor U14485 (N_14485,N_11004,N_8422);
xor U14486 (N_14486,N_10704,N_6683);
xnor U14487 (N_14487,N_6924,N_8071);
nor U14488 (N_14488,N_8709,N_8420);
xor U14489 (N_14489,N_11961,N_6980);
xnor U14490 (N_14490,N_9295,N_6105);
nand U14491 (N_14491,N_11346,N_9008);
or U14492 (N_14492,N_10478,N_8149);
nor U14493 (N_14493,N_6203,N_9122);
and U14494 (N_14494,N_11096,N_9532);
nand U14495 (N_14495,N_11311,N_7168);
nand U14496 (N_14496,N_8822,N_9824);
or U14497 (N_14497,N_7776,N_9633);
nand U14498 (N_14498,N_8952,N_6819);
and U14499 (N_14499,N_8458,N_11864);
nor U14500 (N_14500,N_8742,N_11894);
nand U14501 (N_14501,N_10928,N_10097);
nor U14502 (N_14502,N_8972,N_6045);
or U14503 (N_14503,N_10708,N_8976);
or U14504 (N_14504,N_9850,N_9161);
xor U14505 (N_14505,N_7897,N_11948);
nand U14506 (N_14506,N_7162,N_11050);
and U14507 (N_14507,N_10183,N_10303);
nand U14508 (N_14508,N_11389,N_10903);
nand U14509 (N_14509,N_6323,N_11579);
nor U14510 (N_14510,N_11722,N_6636);
or U14511 (N_14511,N_6061,N_6355);
nand U14512 (N_14512,N_10519,N_10254);
xor U14513 (N_14513,N_6617,N_7670);
and U14514 (N_14514,N_6154,N_8465);
or U14515 (N_14515,N_10194,N_6379);
nand U14516 (N_14516,N_11454,N_9821);
xor U14517 (N_14517,N_8837,N_10135);
and U14518 (N_14518,N_11128,N_9436);
and U14519 (N_14519,N_10763,N_9349);
or U14520 (N_14520,N_10726,N_7814);
nand U14521 (N_14521,N_8132,N_7339);
and U14522 (N_14522,N_6650,N_8388);
nand U14523 (N_14523,N_7429,N_10454);
nor U14524 (N_14524,N_11524,N_8274);
nand U14525 (N_14525,N_8478,N_7337);
nand U14526 (N_14526,N_10808,N_9909);
and U14527 (N_14527,N_8145,N_7822);
nor U14528 (N_14528,N_9362,N_7169);
and U14529 (N_14529,N_6008,N_10065);
and U14530 (N_14530,N_11561,N_8224);
or U14531 (N_14531,N_10423,N_6850);
nor U14532 (N_14532,N_8629,N_7438);
nor U14533 (N_14533,N_9724,N_10772);
nor U14534 (N_14534,N_10169,N_9795);
and U14535 (N_14535,N_7263,N_6514);
or U14536 (N_14536,N_10723,N_11020);
xnor U14537 (N_14537,N_10468,N_6498);
or U14538 (N_14538,N_10945,N_11015);
xnor U14539 (N_14539,N_9670,N_11169);
or U14540 (N_14540,N_10231,N_6754);
or U14541 (N_14541,N_9426,N_6393);
or U14542 (N_14542,N_9118,N_10120);
nor U14543 (N_14543,N_6041,N_8435);
nand U14544 (N_14544,N_8895,N_7205);
and U14545 (N_14545,N_11340,N_10664);
or U14546 (N_14546,N_10922,N_9783);
xnor U14547 (N_14547,N_10284,N_8689);
nor U14548 (N_14548,N_11735,N_11799);
nand U14549 (N_14549,N_7531,N_11302);
or U14550 (N_14550,N_6182,N_7033);
nand U14551 (N_14551,N_8704,N_6745);
xnor U14552 (N_14552,N_10162,N_8718);
nand U14553 (N_14553,N_6444,N_8932);
nor U14554 (N_14554,N_6062,N_8607);
nor U14555 (N_14555,N_11453,N_6305);
or U14556 (N_14556,N_11327,N_11534);
nand U14557 (N_14557,N_6167,N_6453);
and U14558 (N_14558,N_8010,N_9664);
or U14559 (N_14559,N_9554,N_6947);
nor U14560 (N_14560,N_11660,N_10594);
nor U14561 (N_14561,N_11905,N_6704);
or U14562 (N_14562,N_11954,N_7396);
nor U14563 (N_14563,N_6389,N_6372);
and U14564 (N_14564,N_9219,N_9913);
and U14565 (N_14565,N_7582,N_9148);
and U14566 (N_14566,N_9822,N_7688);
or U14567 (N_14567,N_6867,N_8116);
nor U14568 (N_14568,N_11743,N_9339);
and U14569 (N_14569,N_8316,N_11310);
and U14570 (N_14570,N_9430,N_7573);
or U14571 (N_14571,N_10791,N_7435);
nand U14572 (N_14572,N_8407,N_6439);
or U14573 (N_14573,N_6532,N_6369);
or U14574 (N_14574,N_10286,N_10824);
nor U14575 (N_14575,N_6941,N_9060);
nor U14576 (N_14576,N_10986,N_9777);
nand U14577 (N_14577,N_7833,N_7403);
or U14578 (N_14578,N_10222,N_10046);
and U14579 (N_14579,N_7943,N_11253);
nor U14580 (N_14580,N_10764,N_10353);
nand U14581 (N_14581,N_10648,N_10490);
nand U14582 (N_14582,N_8280,N_7842);
nand U14583 (N_14583,N_9472,N_11607);
nor U14584 (N_14584,N_11844,N_7357);
nand U14585 (N_14585,N_6957,N_9494);
or U14586 (N_14586,N_11670,N_9688);
xnor U14587 (N_14587,N_9248,N_10133);
nor U14588 (N_14588,N_11276,N_7427);
xnor U14589 (N_14589,N_8396,N_7661);
xnor U14590 (N_14590,N_11859,N_9424);
nor U14591 (N_14591,N_6161,N_10562);
nor U14592 (N_14592,N_11289,N_6733);
and U14593 (N_14593,N_9465,N_6805);
or U14594 (N_14594,N_7980,N_11125);
or U14595 (N_14595,N_11137,N_8914);
and U14596 (N_14596,N_11792,N_8126);
and U14597 (N_14597,N_11264,N_7804);
or U14598 (N_14598,N_10732,N_11942);
nor U14599 (N_14599,N_11876,N_11063);
nor U14600 (N_14600,N_10274,N_8827);
nand U14601 (N_14601,N_8359,N_6217);
nor U14602 (N_14602,N_6915,N_6813);
or U14603 (N_14603,N_7919,N_9561);
nand U14604 (N_14604,N_11391,N_7750);
xnor U14605 (N_14605,N_11331,N_6770);
and U14606 (N_14606,N_7457,N_8745);
and U14607 (N_14607,N_9989,N_6536);
nand U14608 (N_14608,N_8757,N_10505);
nand U14609 (N_14609,N_7836,N_6402);
or U14610 (N_14610,N_6095,N_11821);
and U14611 (N_14611,N_10400,N_7838);
nor U14612 (N_14612,N_8852,N_9196);
nor U14613 (N_14613,N_8658,N_11202);
nor U14614 (N_14614,N_8810,N_11282);
nor U14615 (N_14615,N_7883,N_8172);
nand U14616 (N_14616,N_6656,N_6480);
or U14617 (N_14617,N_8443,N_11970);
and U14618 (N_14618,N_7604,N_6433);
xor U14619 (N_14619,N_6703,N_9178);
nand U14620 (N_14620,N_11718,N_11504);
or U14621 (N_14621,N_10413,N_7005);
xnor U14622 (N_14622,N_11035,N_6896);
nor U14623 (N_14623,N_8389,N_7062);
and U14624 (N_14624,N_9007,N_8603);
and U14625 (N_14625,N_6321,N_6275);
and U14626 (N_14626,N_6548,N_9635);
nand U14627 (N_14627,N_6053,N_10595);
nand U14628 (N_14628,N_8824,N_9235);
xor U14629 (N_14629,N_7562,N_7700);
and U14630 (N_14630,N_6391,N_10757);
or U14631 (N_14631,N_8253,N_9841);
nand U14632 (N_14632,N_10428,N_8830);
or U14633 (N_14633,N_11574,N_6560);
or U14634 (N_14634,N_7652,N_7971);
nor U14635 (N_14635,N_11944,N_11975);
and U14636 (N_14636,N_10069,N_9174);
xor U14637 (N_14637,N_8740,N_8521);
and U14638 (N_14638,N_10124,N_6421);
or U14639 (N_14639,N_9321,N_6224);
nor U14640 (N_14640,N_9285,N_8189);
nor U14641 (N_14641,N_8361,N_9672);
nand U14642 (N_14642,N_10999,N_7934);
or U14643 (N_14643,N_6817,N_6163);
or U14644 (N_14644,N_6952,N_6849);
and U14645 (N_14645,N_6187,N_11133);
nand U14646 (N_14646,N_6236,N_11755);
or U14647 (N_14647,N_10064,N_8161);
xor U14648 (N_14648,N_9281,N_7605);
nand U14649 (N_14649,N_6245,N_6183);
nand U14650 (N_14650,N_8502,N_8295);
xnor U14651 (N_14651,N_10417,N_7172);
nor U14652 (N_14652,N_11674,N_8594);
xnor U14653 (N_14653,N_6101,N_9152);
nand U14654 (N_14654,N_9760,N_10043);
nand U14655 (N_14655,N_11397,N_6982);
nand U14656 (N_14656,N_7632,N_10402);
xnor U14657 (N_14657,N_11054,N_6688);
nand U14658 (N_14658,N_6508,N_6249);
and U14659 (N_14659,N_9079,N_7030);
and U14660 (N_14660,N_9288,N_7719);
nor U14661 (N_14661,N_6872,N_10422);
and U14662 (N_14662,N_11298,N_9862);
or U14663 (N_14663,N_11424,N_8604);
or U14664 (N_14664,N_6907,N_8542);
nand U14665 (N_14665,N_10443,N_10933);
nor U14666 (N_14666,N_10384,N_6020);
nor U14667 (N_14667,N_9661,N_9834);
nor U14668 (N_14668,N_8656,N_10733);
nand U14669 (N_14669,N_10769,N_6499);
xor U14670 (N_14670,N_7672,N_11939);
or U14671 (N_14671,N_9396,N_9381);
nor U14672 (N_14672,N_11965,N_7151);
nor U14673 (N_14673,N_6301,N_11846);
nor U14674 (N_14674,N_11522,N_6271);
nand U14675 (N_14675,N_6405,N_6761);
nand U14676 (N_14676,N_7401,N_8122);
nand U14677 (N_14677,N_7868,N_10316);
and U14678 (N_14678,N_8349,N_10619);
or U14679 (N_14679,N_10461,N_10608);
or U14680 (N_14680,N_9675,N_8043);
and U14681 (N_14681,N_6708,N_9816);
xor U14682 (N_14682,N_8855,N_7071);
xor U14683 (N_14683,N_11367,N_8911);
and U14684 (N_14684,N_7752,N_6899);
nand U14685 (N_14685,N_8514,N_11064);
nand U14686 (N_14686,N_6197,N_11515);
and U14687 (N_14687,N_6418,N_8485);
nand U14688 (N_14688,N_6713,N_8457);
or U14689 (N_14689,N_11998,N_9952);
nand U14690 (N_14690,N_7981,N_10580);
nand U14691 (N_14691,N_8304,N_10551);
nand U14692 (N_14692,N_10205,N_11151);
nor U14693 (N_14693,N_6410,N_9625);
xor U14694 (N_14694,N_11045,N_9311);
and U14695 (N_14695,N_8957,N_10375);
nand U14696 (N_14696,N_7659,N_10601);
nand U14697 (N_14697,N_8394,N_9947);
and U14698 (N_14698,N_8725,N_9479);
nand U14699 (N_14699,N_7240,N_9845);
xnor U14700 (N_14700,N_10451,N_8221);
xor U14701 (N_14701,N_7025,N_9301);
nor U14702 (N_14702,N_8477,N_7938);
nand U14703 (N_14703,N_11672,N_8390);
nor U14704 (N_14704,N_8442,N_11725);
xor U14705 (N_14705,N_10520,N_9404);
nand U14706 (N_14706,N_8804,N_11828);
nand U14707 (N_14707,N_11889,N_10131);
or U14708 (N_14708,N_11084,N_11762);
and U14709 (N_14709,N_6918,N_11166);
or U14710 (N_14710,N_8554,N_7402);
or U14711 (N_14711,N_8601,N_9993);
xnor U14712 (N_14712,N_9987,N_7601);
nor U14713 (N_14713,N_10885,N_7279);
or U14714 (N_14714,N_8906,N_9225);
nor U14715 (N_14715,N_9829,N_7881);
nand U14716 (N_14716,N_6500,N_6848);
or U14717 (N_14717,N_10871,N_6272);
nand U14718 (N_14718,N_11983,N_8708);
nand U14719 (N_14719,N_6592,N_11587);
nand U14720 (N_14720,N_10760,N_9466);
or U14721 (N_14721,N_10753,N_8943);
nor U14722 (N_14722,N_11193,N_10385);
and U14723 (N_14723,N_11531,N_10570);
xor U14724 (N_14724,N_7683,N_7416);
nand U14725 (N_14725,N_7812,N_10216);
and U14726 (N_14726,N_11913,N_10489);
nand U14727 (N_14727,N_9660,N_9906);
or U14728 (N_14728,N_7365,N_7272);
or U14729 (N_14729,N_11624,N_10045);
xnor U14730 (N_14730,N_10474,N_8177);
or U14731 (N_14731,N_9224,N_9229);
and U14732 (N_14732,N_11414,N_9033);
xnor U14733 (N_14733,N_7011,N_6839);
or U14734 (N_14734,N_10526,N_8204);
and U14735 (N_14735,N_10287,N_6694);
nand U14736 (N_14736,N_9533,N_6373);
or U14737 (N_14737,N_11935,N_10567);
or U14738 (N_14738,N_10749,N_8715);
nor U14739 (N_14739,N_10122,N_9946);
nor U14740 (N_14740,N_8200,N_6509);
or U14741 (N_14741,N_9130,N_6086);
or U14742 (N_14742,N_10529,N_6200);
nor U14743 (N_14743,N_10813,N_7382);
and U14744 (N_14744,N_8121,N_11477);
or U14745 (N_14745,N_6854,N_10242);
nor U14746 (N_14746,N_9416,N_8741);
nand U14747 (N_14747,N_6572,N_9932);
xnor U14748 (N_14748,N_10301,N_9053);
or U14749 (N_14749,N_11266,N_8136);
and U14750 (N_14750,N_10960,N_6639);
or U14751 (N_14751,N_7962,N_8630);
nor U14752 (N_14752,N_9128,N_6329);
and U14753 (N_14753,N_8141,N_7867);
and U14754 (N_14754,N_11222,N_11027);
nand U14755 (N_14755,N_9725,N_9752);
nand U14756 (N_14756,N_8053,N_6414);
or U14757 (N_14757,N_10224,N_6939);
and U14758 (N_14758,N_8755,N_10995);
or U14759 (N_14759,N_10610,N_7320);
nor U14760 (N_14760,N_8444,N_7483);
nor U14761 (N_14761,N_7874,N_9809);
xor U14762 (N_14762,N_7809,N_11836);
or U14763 (N_14763,N_6974,N_9209);
and U14764 (N_14764,N_8989,N_7504);
xor U14765 (N_14765,N_6429,N_6119);
xor U14766 (N_14766,N_7768,N_8753);
xor U14767 (N_14767,N_6920,N_7329);
nand U14768 (N_14768,N_11956,N_10861);
xor U14769 (N_14769,N_10028,N_10456);
or U14770 (N_14770,N_6201,N_11727);
nand U14771 (N_14771,N_6787,N_7628);
nor U14772 (N_14772,N_7230,N_8868);
and U14773 (N_14773,N_11543,N_6487);
xor U14774 (N_14774,N_6661,N_11612);
and U14775 (N_14775,N_7995,N_9238);
nand U14776 (N_14776,N_10822,N_9210);
and U14777 (N_14777,N_7942,N_7974);
nand U14778 (N_14778,N_9745,N_6012);
or U14779 (N_14779,N_9193,N_10263);
xnor U14780 (N_14780,N_10157,N_11460);
xor U14781 (N_14781,N_10471,N_7730);
or U14782 (N_14782,N_6818,N_8180);
nor U14783 (N_14783,N_10138,N_8900);
nor U14784 (N_14784,N_9332,N_7449);
nand U14785 (N_14785,N_10492,N_10892);
nand U14786 (N_14786,N_9092,N_10038);
and U14787 (N_14787,N_9503,N_10781);
or U14788 (N_14788,N_7610,N_9179);
nor U14789 (N_14789,N_8886,N_11541);
and U14790 (N_14790,N_7755,N_10198);
or U14791 (N_14791,N_8954,N_7054);
and U14792 (N_14792,N_9775,N_11172);
nand U14793 (N_14793,N_10132,N_9585);
nand U14794 (N_14794,N_6658,N_9971);
xnor U14795 (N_14795,N_11491,N_7829);
xnor U14796 (N_14796,N_8068,N_6122);
nand U14797 (N_14797,N_6871,N_10240);
or U14798 (N_14798,N_10006,N_10459);
nand U14799 (N_14799,N_10988,N_9348);
and U14800 (N_14800,N_11348,N_11763);
and U14801 (N_14801,N_10909,N_6965);
or U14802 (N_14802,N_10015,N_11153);
nor U14803 (N_14803,N_6963,N_9350);
xnor U14804 (N_14804,N_8798,N_11051);
and U14805 (N_14805,N_7358,N_10819);
nand U14806 (N_14806,N_9520,N_7315);
nor U14807 (N_14807,N_8369,N_9891);
nor U14808 (N_14808,N_6785,N_9183);
xnor U14809 (N_14809,N_11530,N_6581);
xor U14810 (N_14810,N_7219,N_6097);
and U14811 (N_14811,N_7211,N_8308);
xnor U14812 (N_14812,N_10956,N_6728);
nand U14813 (N_14813,N_7210,N_11089);
or U14814 (N_14814,N_8456,N_7856);
nand U14815 (N_14815,N_8893,N_8252);
nor U14816 (N_14816,N_9085,N_10425);
and U14817 (N_14817,N_6706,N_10049);
and U14818 (N_14818,N_6497,N_11149);
and U14819 (N_14819,N_11899,N_8831);
xor U14820 (N_14820,N_7818,N_8840);
or U14821 (N_14821,N_11072,N_6857);
or U14822 (N_14822,N_7800,N_11620);
or U14823 (N_14823,N_7321,N_7292);
and U14824 (N_14824,N_10020,N_6149);
and U14825 (N_14825,N_6353,N_6676);
xor U14826 (N_14826,N_9953,N_10883);
or U14827 (N_14827,N_9009,N_8566);
nand U14828 (N_14828,N_9071,N_11417);
nand U14829 (N_14829,N_10418,N_9594);
nor U14830 (N_14830,N_6022,N_8535);
nand U14831 (N_14831,N_10512,N_6371);
nand U14832 (N_14832,N_8598,N_8862);
nor U14833 (N_14833,N_6599,N_11010);
nand U14834 (N_14834,N_11352,N_8552);
nand U14835 (N_14835,N_9146,N_10479);
nor U14836 (N_14836,N_8243,N_10346);
or U14837 (N_14837,N_8345,N_9511);
nor U14838 (N_14838,N_10965,N_10536);
or U14839 (N_14839,N_8266,N_6773);
xor U14840 (N_14840,N_6125,N_7921);
xnor U14841 (N_14841,N_10522,N_6407);
nor U14842 (N_14842,N_9980,N_9012);
and U14843 (N_14843,N_10424,N_11863);
and U14844 (N_14844,N_7193,N_9758);
nand U14845 (N_14845,N_6715,N_11225);
or U14846 (N_14846,N_6897,N_10559);
nand U14847 (N_14847,N_11226,N_9988);
nor U14848 (N_14848,N_6004,N_6891);
nor U14849 (N_14849,N_11381,N_7544);
xor U14850 (N_14850,N_11684,N_6593);
xor U14851 (N_14851,N_11703,N_7721);
xor U14852 (N_14852,N_7246,N_9211);
nand U14853 (N_14853,N_7704,N_11361);
nand U14854 (N_14854,N_10345,N_6338);
nand U14855 (N_14855,N_10656,N_9275);
nand U14856 (N_14856,N_10919,N_8791);
nand U14857 (N_14857,N_11109,N_8337);
and U14858 (N_14858,N_11926,N_7891);
and U14859 (N_14859,N_8760,N_8703);
xor U14860 (N_14860,N_6695,N_8467);
and U14861 (N_14861,N_8951,N_8078);
or U14862 (N_14862,N_7540,N_11536);
or U14863 (N_14863,N_8700,N_6056);
or U14864 (N_14864,N_10342,N_7530);
and U14865 (N_14865,N_7256,N_8577);
nand U14866 (N_14866,N_7828,N_7621);
xnor U14867 (N_14867,N_7489,N_10127);
and U14868 (N_14868,N_7377,N_10074);
or U14869 (N_14869,N_8842,N_10978);
nand U14870 (N_14870,N_7109,N_9419);
nand U14871 (N_14871,N_9628,N_6681);
or U14872 (N_14872,N_8195,N_11368);
nor U14873 (N_14873,N_7298,N_9454);
or U14874 (N_14874,N_7439,N_11479);
and U14875 (N_14875,N_7164,N_7674);
and U14876 (N_14876,N_8330,N_9254);
nand U14877 (N_14877,N_7736,N_11262);
and U14878 (N_14878,N_8296,N_9886);
nor U14879 (N_14879,N_7235,N_9272);
nor U14880 (N_14880,N_11834,N_6103);
and U14881 (N_14881,N_11174,N_11992);
nor U14882 (N_14882,N_11987,N_6512);
nor U14883 (N_14883,N_8281,N_11608);
nand U14884 (N_14884,N_11766,N_11719);
nor U14885 (N_14885,N_9742,N_6832);
and U14886 (N_14886,N_10359,N_9449);
and U14887 (N_14887,N_7371,N_7326);
or U14888 (N_14888,N_9277,N_9832);
and U14889 (N_14889,N_8484,N_6516);
and U14890 (N_14890,N_10434,N_10632);
xnor U14891 (N_14891,N_7969,N_11555);
or U14892 (N_14892,N_8960,N_9413);
xor U14893 (N_14893,N_7834,N_10361);
nor U14894 (N_14894,N_9379,N_10767);
xnor U14895 (N_14895,N_10638,N_9282);
and U14896 (N_14896,N_6943,N_8624);
xor U14897 (N_14897,N_7455,N_11481);
and U14898 (N_14898,N_8391,N_11881);
nor U14899 (N_14899,N_10408,N_7348);
or U14900 (N_14900,N_6736,N_9187);
or U14901 (N_14901,N_8533,N_11665);
nor U14902 (N_14902,N_10748,N_8897);
or U14903 (N_14903,N_11251,N_6111);
nor U14904 (N_14904,N_7702,N_7645);
or U14905 (N_14905,N_9754,N_8286);
xnor U14906 (N_14906,N_11994,N_8237);
or U14907 (N_14907,N_10007,N_11825);
nor U14908 (N_14908,N_8712,N_9175);
and U14909 (N_14909,N_9308,N_7300);
nor U14910 (N_14910,N_7477,N_8534);
nand U14911 (N_14911,N_10154,N_11576);
or U14912 (N_14912,N_10259,N_7386);
xor U14913 (N_14913,N_11338,N_10104);
or U14914 (N_14914,N_10188,N_9749);
nand U14915 (N_14915,N_6827,N_8167);
or U14916 (N_14916,N_8586,N_7692);
or U14917 (N_14917,N_8883,N_11605);
nand U14918 (N_14918,N_9228,N_10525);
or U14919 (N_14919,N_6196,N_11150);
nand U14920 (N_14920,N_6747,N_11938);
xor U14921 (N_14921,N_8505,N_9151);
xnor U14922 (N_14922,N_8375,N_8826);
nand U14923 (N_14923,N_8028,N_9029);
or U14924 (N_14924,N_9734,N_7744);
or U14925 (N_14925,N_7879,N_9710);
nor U14926 (N_14926,N_9912,N_10882);
and U14927 (N_14927,N_11919,N_9488);
nand U14928 (N_14928,N_11366,N_6969);
nor U14929 (N_14929,N_11384,N_10168);
xnor U14930 (N_14930,N_9644,N_11879);
xor U14931 (N_14931,N_7249,N_6674);
xor U14932 (N_14932,N_6578,N_11511);
nand U14933 (N_14933,N_7825,N_9064);
nor U14934 (N_14934,N_9249,N_9376);
or U14935 (N_14935,N_8517,N_6215);
nor U14936 (N_14936,N_6929,N_8711);
nor U14937 (N_14937,N_10604,N_10328);
nand U14938 (N_14938,N_11383,N_9527);
or U14939 (N_14939,N_7703,N_10470);
and U14940 (N_14940,N_6553,N_10515);
or U14941 (N_14941,N_7215,N_6816);
or U14942 (N_14942,N_9863,N_10173);
nand U14943 (N_14943,N_9292,N_7086);
and U14944 (N_14944,N_10350,N_10607);
nor U14945 (N_14945,N_11043,N_9172);
nand U14946 (N_14946,N_7859,N_8262);
nand U14947 (N_14947,N_7437,N_8806);
or U14948 (N_14948,N_9112,N_7160);
nor U14949 (N_14949,N_9222,N_7762);
nor U14950 (N_14950,N_6357,N_6997);
and U14951 (N_14951,N_9046,N_7810);
and U14952 (N_14952,N_9764,N_8950);
or U14953 (N_14953,N_7614,N_7787);
nand U14954 (N_14954,N_7607,N_11748);
nor U14955 (N_14955,N_7739,N_10917);
and U14956 (N_14956,N_9898,N_7753);
or U14957 (N_14957,N_11257,N_11869);
xnor U14958 (N_14958,N_6976,N_6790);
nand U14959 (N_14959,N_8618,N_10042);
xnor U14960 (N_14960,N_9543,N_9961);
xnor U14961 (N_14961,N_10724,N_8148);
xnor U14962 (N_14962,N_8242,N_8108);
nand U14963 (N_14963,N_6804,N_9267);
and U14964 (N_14964,N_11197,N_7383);
xnor U14965 (N_14965,N_10997,N_11595);
and U14966 (N_14966,N_8557,N_8362);
and U14967 (N_14967,N_11851,N_6166);
nand U14968 (N_14968,N_11649,N_9300);
xnor U14969 (N_14969,N_11989,N_9205);
xor U14970 (N_14970,N_11122,N_10300);
and U14971 (N_14971,N_8887,N_7045);
nor U14972 (N_14972,N_6883,N_6148);
and U14973 (N_14973,N_8270,N_8579);
nor U14974 (N_14974,N_7608,N_7171);
nor U14975 (N_14975,N_6668,N_9324);
xnor U14976 (N_14976,N_7701,N_9375);
or U14977 (N_14977,N_8302,N_6792);
and U14978 (N_14978,N_8973,N_7501);
nor U14979 (N_14979,N_7328,N_6781);
xnor U14980 (N_14980,N_6996,N_6811);
and U14981 (N_14981,N_7282,N_10531);
or U14982 (N_14982,N_8664,N_9088);
nand U14983 (N_14983,N_9835,N_7113);
nand U14984 (N_14984,N_6162,N_9123);
or U14985 (N_14985,N_10957,N_8706);
nor U14986 (N_14986,N_7722,N_7906);
nor U14987 (N_14987,N_10081,N_9359);
and U14988 (N_14988,N_10523,N_9039);
nand U14989 (N_14989,N_11452,N_6753);
and U14990 (N_14990,N_9774,N_9851);
nand U14991 (N_14991,N_7069,N_9191);
nand U14992 (N_14992,N_6911,N_11138);
and U14993 (N_14993,N_11533,N_7280);
or U14994 (N_14994,N_11468,N_7111);
nand U14995 (N_14995,N_9978,N_9138);
xor U14996 (N_14996,N_8431,N_7764);
nor U14997 (N_14997,N_7696,N_9602);
nor U14998 (N_14998,N_9393,N_10151);
nor U14999 (N_14999,N_8899,N_9571);
or U15000 (N_15000,N_11176,N_10522);
xnor U15001 (N_15001,N_11336,N_6831);
nor U15002 (N_15002,N_8241,N_11068);
and U15003 (N_15003,N_6045,N_11102);
and U15004 (N_15004,N_10125,N_7954);
nor U15005 (N_15005,N_9704,N_8713);
and U15006 (N_15006,N_8542,N_8681);
or U15007 (N_15007,N_6650,N_6050);
nand U15008 (N_15008,N_9745,N_9213);
nor U15009 (N_15009,N_8578,N_11459);
and U15010 (N_15010,N_10680,N_11443);
xor U15011 (N_15011,N_7364,N_6258);
nand U15012 (N_15012,N_10809,N_6761);
and U15013 (N_15013,N_10171,N_9275);
nand U15014 (N_15014,N_7231,N_7702);
nor U15015 (N_15015,N_6899,N_10335);
xor U15016 (N_15016,N_6871,N_6542);
and U15017 (N_15017,N_7706,N_11323);
or U15018 (N_15018,N_11950,N_6171);
nor U15019 (N_15019,N_10791,N_8150);
or U15020 (N_15020,N_10352,N_6775);
nor U15021 (N_15021,N_11344,N_7699);
nand U15022 (N_15022,N_8351,N_6719);
nand U15023 (N_15023,N_8738,N_9913);
and U15024 (N_15024,N_6979,N_9725);
xor U15025 (N_15025,N_7192,N_9724);
and U15026 (N_15026,N_6195,N_6644);
xnor U15027 (N_15027,N_6733,N_8886);
nor U15028 (N_15028,N_10487,N_7909);
nand U15029 (N_15029,N_8246,N_8761);
nand U15030 (N_15030,N_7224,N_8367);
or U15031 (N_15031,N_8012,N_10506);
xnor U15032 (N_15032,N_10289,N_11995);
xnor U15033 (N_15033,N_7214,N_10504);
or U15034 (N_15034,N_9014,N_8227);
nor U15035 (N_15035,N_7142,N_7742);
nand U15036 (N_15036,N_8376,N_9677);
nor U15037 (N_15037,N_7779,N_10381);
xor U15038 (N_15038,N_6565,N_6627);
or U15039 (N_15039,N_7116,N_9958);
and U15040 (N_15040,N_9390,N_9228);
nand U15041 (N_15041,N_9541,N_7679);
xor U15042 (N_15042,N_8280,N_8032);
nand U15043 (N_15043,N_10269,N_9544);
xor U15044 (N_15044,N_7243,N_7591);
or U15045 (N_15045,N_6776,N_7215);
xor U15046 (N_15046,N_7520,N_11044);
and U15047 (N_15047,N_6861,N_10995);
xnor U15048 (N_15048,N_6308,N_11175);
nor U15049 (N_15049,N_10241,N_7725);
nor U15050 (N_15050,N_8829,N_10792);
xnor U15051 (N_15051,N_7801,N_6358);
nor U15052 (N_15052,N_7441,N_7579);
xnor U15053 (N_15053,N_9167,N_6214);
or U15054 (N_15054,N_9545,N_11283);
or U15055 (N_15055,N_11731,N_6184);
and U15056 (N_15056,N_7670,N_8975);
nor U15057 (N_15057,N_11694,N_7566);
and U15058 (N_15058,N_10111,N_10597);
nor U15059 (N_15059,N_11757,N_11300);
or U15060 (N_15060,N_11031,N_7184);
xnor U15061 (N_15061,N_9237,N_6921);
and U15062 (N_15062,N_10130,N_8255);
nand U15063 (N_15063,N_6797,N_10191);
xor U15064 (N_15064,N_8347,N_6249);
or U15065 (N_15065,N_9327,N_9068);
xor U15066 (N_15066,N_6999,N_11315);
xor U15067 (N_15067,N_9891,N_6651);
xor U15068 (N_15068,N_11185,N_8746);
and U15069 (N_15069,N_9102,N_6870);
xnor U15070 (N_15070,N_9040,N_10583);
and U15071 (N_15071,N_6531,N_6439);
nor U15072 (N_15072,N_11569,N_7416);
or U15073 (N_15073,N_11548,N_11219);
nand U15074 (N_15074,N_6376,N_8694);
xor U15075 (N_15075,N_7135,N_9245);
nand U15076 (N_15076,N_9182,N_6156);
or U15077 (N_15077,N_9392,N_8539);
xnor U15078 (N_15078,N_11597,N_10801);
nor U15079 (N_15079,N_11448,N_10132);
nor U15080 (N_15080,N_10438,N_9638);
and U15081 (N_15081,N_10365,N_7002);
nand U15082 (N_15082,N_7225,N_9190);
nor U15083 (N_15083,N_8064,N_10879);
xnor U15084 (N_15084,N_7457,N_9200);
and U15085 (N_15085,N_8905,N_9388);
xnor U15086 (N_15086,N_7752,N_9065);
xnor U15087 (N_15087,N_6402,N_11110);
nand U15088 (N_15088,N_7401,N_8092);
nor U15089 (N_15089,N_8817,N_11561);
and U15090 (N_15090,N_10109,N_11887);
nor U15091 (N_15091,N_6906,N_7395);
nor U15092 (N_15092,N_8107,N_8392);
nand U15093 (N_15093,N_9696,N_6997);
and U15094 (N_15094,N_9733,N_6271);
or U15095 (N_15095,N_10038,N_6986);
nor U15096 (N_15096,N_7748,N_11064);
xor U15097 (N_15097,N_8767,N_6045);
xor U15098 (N_15098,N_6676,N_9860);
nand U15099 (N_15099,N_8828,N_10069);
nor U15100 (N_15100,N_8352,N_11997);
and U15101 (N_15101,N_10429,N_11393);
and U15102 (N_15102,N_9821,N_11078);
nor U15103 (N_15103,N_10347,N_7029);
xor U15104 (N_15104,N_11237,N_9610);
nand U15105 (N_15105,N_11197,N_11310);
or U15106 (N_15106,N_9416,N_10083);
nor U15107 (N_15107,N_9120,N_7099);
nor U15108 (N_15108,N_6657,N_8697);
and U15109 (N_15109,N_10183,N_7577);
or U15110 (N_15110,N_9761,N_6996);
xor U15111 (N_15111,N_10841,N_10986);
and U15112 (N_15112,N_8747,N_10886);
and U15113 (N_15113,N_7668,N_9462);
nor U15114 (N_15114,N_9316,N_9584);
or U15115 (N_15115,N_11475,N_9848);
and U15116 (N_15116,N_7294,N_9206);
nor U15117 (N_15117,N_7766,N_9608);
and U15118 (N_15118,N_9634,N_10170);
or U15119 (N_15119,N_9153,N_11337);
nand U15120 (N_15120,N_10758,N_11781);
nor U15121 (N_15121,N_8622,N_9185);
and U15122 (N_15122,N_11337,N_7045);
nand U15123 (N_15123,N_9826,N_11482);
and U15124 (N_15124,N_8198,N_9181);
and U15125 (N_15125,N_9276,N_7191);
and U15126 (N_15126,N_10948,N_6667);
nand U15127 (N_15127,N_11773,N_8746);
nand U15128 (N_15128,N_10893,N_7144);
nand U15129 (N_15129,N_9971,N_7921);
or U15130 (N_15130,N_10942,N_10160);
nor U15131 (N_15131,N_11708,N_9322);
xor U15132 (N_15132,N_10398,N_7279);
nand U15133 (N_15133,N_10235,N_6406);
nor U15134 (N_15134,N_6058,N_9952);
xnor U15135 (N_15135,N_11831,N_6134);
nand U15136 (N_15136,N_9366,N_6176);
and U15137 (N_15137,N_8327,N_7892);
xor U15138 (N_15138,N_11693,N_8673);
xor U15139 (N_15139,N_7935,N_11468);
nand U15140 (N_15140,N_6955,N_6685);
nor U15141 (N_15141,N_6813,N_7901);
nor U15142 (N_15142,N_7920,N_11946);
nor U15143 (N_15143,N_7975,N_7923);
or U15144 (N_15144,N_7371,N_6694);
nor U15145 (N_15145,N_11346,N_10416);
and U15146 (N_15146,N_10321,N_6108);
or U15147 (N_15147,N_7418,N_7338);
xor U15148 (N_15148,N_9140,N_6824);
or U15149 (N_15149,N_6263,N_8332);
xnor U15150 (N_15150,N_8437,N_8039);
nor U15151 (N_15151,N_9714,N_6597);
xnor U15152 (N_15152,N_7431,N_11222);
xnor U15153 (N_15153,N_7481,N_10798);
or U15154 (N_15154,N_6634,N_9326);
xnor U15155 (N_15155,N_10545,N_10139);
nor U15156 (N_15156,N_6837,N_7254);
and U15157 (N_15157,N_7328,N_7694);
xnor U15158 (N_15158,N_7614,N_6339);
or U15159 (N_15159,N_8387,N_10254);
nand U15160 (N_15160,N_7306,N_10031);
or U15161 (N_15161,N_6727,N_9054);
nor U15162 (N_15162,N_11533,N_9559);
or U15163 (N_15163,N_7708,N_6987);
or U15164 (N_15164,N_7469,N_9054);
or U15165 (N_15165,N_7675,N_6487);
nor U15166 (N_15166,N_6129,N_6970);
or U15167 (N_15167,N_8166,N_10543);
or U15168 (N_15168,N_11328,N_7019);
xor U15169 (N_15169,N_9938,N_10367);
nand U15170 (N_15170,N_6593,N_9685);
xnor U15171 (N_15171,N_11291,N_6415);
nand U15172 (N_15172,N_7936,N_11947);
xor U15173 (N_15173,N_11106,N_10523);
xnor U15174 (N_15174,N_6998,N_6037);
nor U15175 (N_15175,N_9043,N_6217);
nor U15176 (N_15176,N_9447,N_7822);
and U15177 (N_15177,N_6180,N_6612);
nand U15178 (N_15178,N_7292,N_8554);
nand U15179 (N_15179,N_10853,N_11868);
nand U15180 (N_15180,N_10951,N_6697);
nor U15181 (N_15181,N_7093,N_7789);
xor U15182 (N_15182,N_7738,N_10919);
xnor U15183 (N_15183,N_9710,N_6540);
and U15184 (N_15184,N_10732,N_11347);
or U15185 (N_15185,N_11204,N_8697);
or U15186 (N_15186,N_8024,N_6450);
xnor U15187 (N_15187,N_9146,N_10896);
nand U15188 (N_15188,N_9767,N_11284);
nor U15189 (N_15189,N_6773,N_6087);
nand U15190 (N_15190,N_7862,N_11994);
or U15191 (N_15191,N_7186,N_7481);
or U15192 (N_15192,N_6009,N_9496);
xor U15193 (N_15193,N_8312,N_9455);
nand U15194 (N_15194,N_7895,N_8703);
xnor U15195 (N_15195,N_10529,N_10923);
nand U15196 (N_15196,N_10361,N_9218);
nor U15197 (N_15197,N_9760,N_11434);
or U15198 (N_15198,N_11083,N_7730);
xnor U15199 (N_15199,N_10350,N_11844);
or U15200 (N_15200,N_9493,N_6883);
nor U15201 (N_15201,N_8879,N_9711);
nand U15202 (N_15202,N_7448,N_9649);
or U15203 (N_15203,N_11813,N_10372);
and U15204 (N_15204,N_10027,N_9058);
nand U15205 (N_15205,N_9494,N_10194);
nor U15206 (N_15206,N_9845,N_9256);
or U15207 (N_15207,N_7376,N_8744);
and U15208 (N_15208,N_8677,N_6634);
xor U15209 (N_15209,N_11659,N_7289);
xor U15210 (N_15210,N_10161,N_6916);
and U15211 (N_15211,N_8988,N_7190);
or U15212 (N_15212,N_11934,N_10837);
xor U15213 (N_15213,N_10826,N_8784);
xor U15214 (N_15214,N_10336,N_10282);
nor U15215 (N_15215,N_6613,N_8529);
and U15216 (N_15216,N_6135,N_9578);
xnor U15217 (N_15217,N_11268,N_9575);
xnor U15218 (N_15218,N_6962,N_11801);
nand U15219 (N_15219,N_8891,N_6272);
xnor U15220 (N_15220,N_8452,N_9024);
nand U15221 (N_15221,N_8853,N_10651);
nor U15222 (N_15222,N_7237,N_7805);
and U15223 (N_15223,N_10180,N_11606);
xor U15224 (N_15224,N_9038,N_11088);
nand U15225 (N_15225,N_6825,N_7145);
and U15226 (N_15226,N_8144,N_9272);
nor U15227 (N_15227,N_10208,N_11328);
and U15228 (N_15228,N_6625,N_8937);
nor U15229 (N_15229,N_10953,N_11968);
or U15230 (N_15230,N_8269,N_7044);
xor U15231 (N_15231,N_9284,N_7723);
or U15232 (N_15232,N_7875,N_9625);
xor U15233 (N_15233,N_10599,N_11150);
xnor U15234 (N_15234,N_11280,N_8329);
xnor U15235 (N_15235,N_11869,N_8588);
xnor U15236 (N_15236,N_11352,N_10088);
nand U15237 (N_15237,N_9066,N_9438);
and U15238 (N_15238,N_9102,N_9011);
or U15239 (N_15239,N_10715,N_9100);
and U15240 (N_15240,N_10116,N_10633);
nand U15241 (N_15241,N_10225,N_11234);
nand U15242 (N_15242,N_7377,N_9738);
and U15243 (N_15243,N_6470,N_11114);
nor U15244 (N_15244,N_8112,N_6919);
or U15245 (N_15245,N_9489,N_10306);
or U15246 (N_15246,N_8752,N_11060);
and U15247 (N_15247,N_11569,N_9150);
nor U15248 (N_15248,N_10802,N_10166);
xnor U15249 (N_15249,N_8251,N_11567);
or U15250 (N_15250,N_6795,N_7071);
and U15251 (N_15251,N_11901,N_7234);
and U15252 (N_15252,N_6827,N_8784);
xor U15253 (N_15253,N_7911,N_9473);
nor U15254 (N_15254,N_6049,N_8494);
nor U15255 (N_15255,N_10249,N_10803);
nand U15256 (N_15256,N_11699,N_6334);
nand U15257 (N_15257,N_6476,N_10285);
nor U15258 (N_15258,N_9279,N_8256);
and U15259 (N_15259,N_10907,N_6747);
and U15260 (N_15260,N_8638,N_11975);
or U15261 (N_15261,N_10920,N_6954);
or U15262 (N_15262,N_9151,N_9207);
nand U15263 (N_15263,N_7257,N_7614);
and U15264 (N_15264,N_10242,N_7702);
nand U15265 (N_15265,N_7967,N_10055);
nor U15266 (N_15266,N_10574,N_11360);
nor U15267 (N_15267,N_6564,N_11945);
nand U15268 (N_15268,N_8698,N_8623);
nand U15269 (N_15269,N_11592,N_10235);
and U15270 (N_15270,N_8046,N_9002);
nor U15271 (N_15271,N_9533,N_7302);
and U15272 (N_15272,N_9237,N_10018);
xnor U15273 (N_15273,N_10568,N_6967);
and U15274 (N_15274,N_7816,N_10063);
nor U15275 (N_15275,N_9392,N_8993);
or U15276 (N_15276,N_6572,N_10692);
or U15277 (N_15277,N_6369,N_8399);
nand U15278 (N_15278,N_6527,N_11081);
and U15279 (N_15279,N_7074,N_7055);
and U15280 (N_15280,N_11162,N_6888);
or U15281 (N_15281,N_8850,N_10855);
nand U15282 (N_15282,N_8370,N_7285);
and U15283 (N_15283,N_7639,N_7979);
and U15284 (N_15284,N_7091,N_10369);
nor U15285 (N_15285,N_7718,N_8847);
xnor U15286 (N_15286,N_10252,N_11127);
or U15287 (N_15287,N_7134,N_7924);
xor U15288 (N_15288,N_11952,N_10013);
xor U15289 (N_15289,N_8527,N_7505);
nand U15290 (N_15290,N_8915,N_9008);
or U15291 (N_15291,N_9356,N_8474);
xnor U15292 (N_15292,N_8814,N_11471);
or U15293 (N_15293,N_11736,N_8657);
nand U15294 (N_15294,N_8217,N_7318);
nor U15295 (N_15295,N_11714,N_8671);
nor U15296 (N_15296,N_10435,N_8308);
nor U15297 (N_15297,N_10043,N_10451);
nor U15298 (N_15298,N_6104,N_7034);
xnor U15299 (N_15299,N_10353,N_7652);
nand U15300 (N_15300,N_7335,N_7547);
and U15301 (N_15301,N_10220,N_8320);
and U15302 (N_15302,N_9874,N_11821);
nand U15303 (N_15303,N_8065,N_9926);
or U15304 (N_15304,N_9525,N_6751);
nand U15305 (N_15305,N_11424,N_10227);
nor U15306 (N_15306,N_11054,N_8484);
xor U15307 (N_15307,N_8426,N_10548);
xnor U15308 (N_15308,N_11168,N_8224);
and U15309 (N_15309,N_7085,N_11700);
xor U15310 (N_15310,N_7669,N_8526);
and U15311 (N_15311,N_11386,N_7514);
xor U15312 (N_15312,N_7675,N_7579);
or U15313 (N_15313,N_10712,N_8149);
xnor U15314 (N_15314,N_7766,N_7942);
xor U15315 (N_15315,N_10792,N_9972);
or U15316 (N_15316,N_7416,N_6244);
or U15317 (N_15317,N_8247,N_6133);
or U15318 (N_15318,N_6765,N_8602);
nand U15319 (N_15319,N_6314,N_11733);
and U15320 (N_15320,N_8427,N_6950);
nor U15321 (N_15321,N_11246,N_7976);
or U15322 (N_15322,N_9122,N_11412);
or U15323 (N_15323,N_6374,N_6182);
nor U15324 (N_15324,N_8911,N_7387);
xor U15325 (N_15325,N_8487,N_7876);
nor U15326 (N_15326,N_10508,N_11185);
and U15327 (N_15327,N_8584,N_9879);
xnor U15328 (N_15328,N_8729,N_7791);
and U15329 (N_15329,N_6382,N_10761);
xor U15330 (N_15330,N_10247,N_11296);
nand U15331 (N_15331,N_7701,N_7892);
and U15332 (N_15332,N_9707,N_6455);
or U15333 (N_15333,N_10144,N_9179);
and U15334 (N_15334,N_8958,N_7154);
and U15335 (N_15335,N_9651,N_7324);
and U15336 (N_15336,N_11520,N_9599);
nor U15337 (N_15337,N_10881,N_10565);
and U15338 (N_15338,N_6091,N_11712);
and U15339 (N_15339,N_11154,N_11980);
nand U15340 (N_15340,N_7339,N_10087);
nand U15341 (N_15341,N_7387,N_10362);
xor U15342 (N_15342,N_9058,N_10028);
and U15343 (N_15343,N_7796,N_7324);
nor U15344 (N_15344,N_7444,N_6978);
nor U15345 (N_15345,N_11619,N_8887);
nand U15346 (N_15346,N_7942,N_11342);
nor U15347 (N_15347,N_11566,N_8645);
xnor U15348 (N_15348,N_6505,N_6287);
nor U15349 (N_15349,N_6931,N_10470);
or U15350 (N_15350,N_8678,N_11007);
or U15351 (N_15351,N_6445,N_10022);
xor U15352 (N_15352,N_10287,N_10824);
and U15353 (N_15353,N_8654,N_9432);
nor U15354 (N_15354,N_10282,N_11325);
nand U15355 (N_15355,N_8777,N_7167);
and U15356 (N_15356,N_6787,N_8556);
xor U15357 (N_15357,N_8582,N_9840);
or U15358 (N_15358,N_11003,N_7442);
nand U15359 (N_15359,N_7705,N_7006);
xor U15360 (N_15360,N_9620,N_6978);
or U15361 (N_15361,N_7077,N_9903);
or U15362 (N_15362,N_10928,N_6575);
xor U15363 (N_15363,N_8511,N_6097);
or U15364 (N_15364,N_10892,N_7394);
nand U15365 (N_15365,N_10305,N_7686);
and U15366 (N_15366,N_10503,N_11401);
or U15367 (N_15367,N_6240,N_7793);
nand U15368 (N_15368,N_6114,N_11195);
nand U15369 (N_15369,N_6486,N_8249);
nand U15370 (N_15370,N_8755,N_6935);
nand U15371 (N_15371,N_11483,N_6668);
and U15372 (N_15372,N_9019,N_8251);
xor U15373 (N_15373,N_10679,N_11733);
and U15374 (N_15374,N_11608,N_10067);
nand U15375 (N_15375,N_8183,N_6315);
or U15376 (N_15376,N_9929,N_7978);
nor U15377 (N_15377,N_11716,N_6782);
xnor U15378 (N_15378,N_7055,N_7343);
and U15379 (N_15379,N_6220,N_7324);
or U15380 (N_15380,N_8979,N_7157);
and U15381 (N_15381,N_11834,N_11670);
or U15382 (N_15382,N_7662,N_7886);
nor U15383 (N_15383,N_6112,N_8207);
xnor U15384 (N_15384,N_10434,N_7539);
or U15385 (N_15385,N_10582,N_6008);
nor U15386 (N_15386,N_7637,N_10053);
nand U15387 (N_15387,N_10820,N_9272);
nand U15388 (N_15388,N_10313,N_9482);
or U15389 (N_15389,N_9264,N_6802);
or U15390 (N_15390,N_7304,N_9960);
and U15391 (N_15391,N_10287,N_10427);
xnor U15392 (N_15392,N_9328,N_9990);
nor U15393 (N_15393,N_8346,N_11161);
nand U15394 (N_15394,N_8594,N_8274);
and U15395 (N_15395,N_7698,N_9382);
and U15396 (N_15396,N_6842,N_9226);
nand U15397 (N_15397,N_7290,N_8417);
nand U15398 (N_15398,N_7568,N_8015);
xor U15399 (N_15399,N_8013,N_9796);
or U15400 (N_15400,N_10797,N_8458);
xor U15401 (N_15401,N_10748,N_11400);
nand U15402 (N_15402,N_10212,N_10665);
and U15403 (N_15403,N_6524,N_9668);
and U15404 (N_15404,N_10696,N_11274);
nor U15405 (N_15405,N_10511,N_11243);
nor U15406 (N_15406,N_10367,N_11049);
nor U15407 (N_15407,N_7356,N_8969);
or U15408 (N_15408,N_8926,N_8906);
and U15409 (N_15409,N_7581,N_9178);
nor U15410 (N_15410,N_10079,N_9173);
nand U15411 (N_15411,N_11914,N_10774);
or U15412 (N_15412,N_6548,N_8748);
and U15413 (N_15413,N_11056,N_10511);
or U15414 (N_15414,N_7913,N_11846);
xor U15415 (N_15415,N_9028,N_11004);
or U15416 (N_15416,N_10474,N_7747);
nor U15417 (N_15417,N_9648,N_7074);
nor U15418 (N_15418,N_6102,N_9800);
or U15419 (N_15419,N_7118,N_6218);
and U15420 (N_15420,N_10170,N_11563);
nor U15421 (N_15421,N_8678,N_10626);
and U15422 (N_15422,N_8102,N_7524);
nand U15423 (N_15423,N_10123,N_11692);
nand U15424 (N_15424,N_10485,N_11960);
xor U15425 (N_15425,N_11854,N_9356);
and U15426 (N_15426,N_10593,N_9993);
xnor U15427 (N_15427,N_9258,N_8887);
nand U15428 (N_15428,N_10271,N_9167);
and U15429 (N_15429,N_11060,N_10810);
nand U15430 (N_15430,N_8379,N_10168);
nand U15431 (N_15431,N_9216,N_10692);
xnor U15432 (N_15432,N_11763,N_7949);
xor U15433 (N_15433,N_11350,N_8186);
nand U15434 (N_15434,N_6416,N_8219);
or U15435 (N_15435,N_8673,N_7129);
nand U15436 (N_15436,N_7937,N_6921);
or U15437 (N_15437,N_8236,N_8617);
nand U15438 (N_15438,N_10086,N_6675);
nand U15439 (N_15439,N_8081,N_11796);
xnor U15440 (N_15440,N_7488,N_11681);
or U15441 (N_15441,N_8019,N_11607);
xor U15442 (N_15442,N_7907,N_7480);
or U15443 (N_15443,N_9418,N_8615);
xor U15444 (N_15444,N_11839,N_11381);
nor U15445 (N_15445,N_10627,N_7428);
nand U15446 (N_15446,N_10364,N_11575);
xnor U15447 (N_15447,N_6097,N_11164);
or U15448 (N_15448,N_8910,N_11053);
xnor U15449 (N_15449,N_9869,N_8025);
nor U15450 (N_15450,N_11406,N_9735);
and U15451 (N_15451,N_10822,N_9090);
xor U15452 (N_15452,N_6104,N_11906);
xnor U15453 (N_15453,N_10416,N_11989);
xnor U15454 (N_15454,N_6615,N_9731);
xnor U15455 (N_15455,N_11024,N_11591);
xor U15456 (N_15456,N_8758,N_9701);
nand U15457 (N_15457,N_6574,N_10527);
or U15458 (N_15458,N_8891,N_6003);
and U15459 (N_15459,N_6563,N_10667);
nand U15460 (N_15460,N_6190,N_9540);
nand U15461 (N_15461,N_6321,N_10400);
xnor U15462 (N_15462,N_10171,N_7894);
or U15463 (N_15463,N_8424,N_10403);
nand U15464 (N_15464,N_11804,N_10261);
and U15465 (N_15465,N_7357,N_7108);
or U15466 (N_15466,N_8588,N_7154);
and U15467 (N_15467,N_9502,N_6215);
nor U15468 (N_15468,N_8955,N_10866);
or U15469 (N_15469,N_9339,N_11505);
and U15470 (N_15470,N_10019,N_6923);
nand U15471 (N_15471,N_8948,N_7470);
xnor U15472 (N_15472,N_9956,N_9503);
and U15473 (N_15473,N_10551,N_9293);
and U15474 (N_15474,N_8460,N_6023);
nor U15475 (N_15475,N_10636,N_10531);
nor U15476 (N_15476,N_6124,N_7300);
nand U15477 (N_15477,N_9705,N_7586);
or U15478 (N_15478,N_10843,N_6721);
nor U15479 (N_15479,N_7883,N_11561);
nand U15480 (N_15480,N_8327,N_9569);
nor U15481 (N_15481,N_10426,N_9289);
and U15482 (N_15482,N_10514,N_6369);
or U15483 (N_15483,N_8073,N_11632);
nor U15484 (N_15484,N_7479,N_6752);
and U15485 (N_15485,N_11617,N_6391);
and U15486 (N_15486,N_10539,N_10369);
xor U15487 (N_15487,N_7805,N_8744);
nand U15488 (N_15488,N_9793,N_8941);
xnor U15489 (N_15489,N_10710,N_11252);
xnor U15490 (N_15490,N_11523,N_10469);
xor U15491 (N_15491,N_10184,N_7554);
xor U15492 (N_15492,N_8988,N_11621);
or U15493 (N_15493,N_11680,N_7428);
nor U15494 (N_15494,N_9230,N_10835);
or U15495 (N_15495,N_11675,N_10089);
xor U15496 (N_15496,N_10071,N_7702);
or U15497 (N_15497,N_11778,N_8771);
nor U15498 (N_15498,N_10755,N_6552);
and U15499 (N_15499,N_7020,N_6763);
and U15500 (N_15500,N_6773,N_8339);
nor U15501 (N_15501,N_7806,N_9500);
xnor U15502 (N_15502,N_7878,N_6141);
nand U15503 (N_15503,N_10785,N_7356);
nor U15504 (N_15504,N_6615,N_7514);
nor U15505 (N_15505,N_7208,N_9226);
or U15506 (N_15506,N_10774,N_7967);
and U15507 (N_15507,N_7937,N_11918);
nor U15508 (N_15508,N_6519,N_11098);
nor U15509 (N_15509,N_11356,N_9016);
or U15510 (N_15510,N_8767,N_11327);
or U15511 (N_15511,N_6347,N_7999);
or U15512 (N_15512,N_10675,N_6186);
nand U15513 (N_15513,N_9727,N_6463);
nand U15514 (N_15514,N_11735,N_8605);
or U15515 (N_15515,N_8639,N_6061);
nor U15516 (N_15516,N_8651,N_8746);
xnor U15517 (N_15517,N_7318,N_11681);
and U15518 (N_15518,N_11126,N_7865);
nand U15519 (N_15519,N_8323,N_7516);
nor U15520 (N_15520,N_9569,N_8405);
or U15521 (N_15521,N_10788,N_9735);
nor U15522 (N_15522,N_8474,N_6207);
nor U15523 (N_15523,N_10525,N_9687);
nor U15524 (N_15524,N_6748,N_10286);
nand U15525 (N_15525,N_11599,N_7200);
nand U15526 (N_15526,N_8154,N_7604);
or U15527 (N_15527,N_8100,N_7748);
or U15528 (N_15528,N_6950,N_6052);
or U15529 (N_15529,N_6454,N_6240);
and U15530 (N_15530,N_9071,N_11609);
or U15531 (N_15531,N_6594,N_7174);
or U15532 (N_15532,N_11588,N_11450);
and U15533 (N_15533,N_8673,N_9698);
or U15534 (N_15534,N_10613,N_11773);
and U15535 (N_15535,N_9426,N_7548);
xnor U15536 (N_15536,N_9739,N_8240);
and U15537 (N_15537,N_6597,N_10525);
nand U15538 (N_15538,N_11294,N_8615);
or U15539 (N_15539,N_10117,N_7976);
or U15540 (N_15540,N_9605,N_6291);
and U15541 (N_15541,N_11329,N_11056);
nand U15542 (N_15542,N_9344,N_6030);
nand U15543 (N_15543,N_9710,N_6906);
or U15544 (N_15544,N_8254,N_7961);
nand U15545 (N_15545,N_9463,N_8605);
or U15546 (N_15546,N_7404,N_8266);
xor U15547 (N_15547,N_7523,N_6367);
or U15548 (N_15548,N_8267,N_9420);
nor U15549 (N_15549,N_11491,N_11826);
nand U15550 (N_15550,N_10656,N_11363);
and U15551 (N_15551,N_10335,N_6447);
nor U15552 (N_15552,N_10864,N_6174);
or U15553 (N_15553,N_8328,N_7001);
nor U15554 (N_15554,N_6182,N_8957);
nor U15555 (N_15555,N_10976,N_11457);
nor U15556 (N_15556,N_10337,N_8913);
nor U15557 (N_15557,N_11776,N_8978);
xor U15558 (N_15558,N_11703,N_7473);
xor U15559 (N_15559,N_10848,N_11421);
or U15560 (N_15560,N_9970,N_8639);
xnor U15561 (N_15561,N_9317,N_10341);
and U15562 (N_15562,N_7007,N_7231);
or U15563 (N_15563,N_7200,N_10373);
nor U15564 (N_15564,N_8203,N_11932);
xnor U15565 (N_15565,N_11444,N_10152);
and U15566 (N_15566,N_10168,N_9986);
or U15567 (N_15567,N_6613,N_8235);
and U15568 (N_15568,N_6513,N_6356);
and U15569 (N_15569,N_6604,N_9694);
xor U15570 (N_15570,N_9757,N_8833);
nand U15571 (N_15571,N_8191,N_10322);
nor U15572 (N_15572,N_9752,N_6208);
or U15573 (N_15573,N_8215,N_9194);
or U15574 (N_15574,N_8485,N_9742);
xor U15575 (N_15575,N_10710,N_8615);
or U15576 (N_15576,N_7646,N_9071);
xnor U15577 (N_15577,N_10301,N_6957);
nand U15578 (N_15578,N_11400,N_11091);
and U15579 (N_15579,N_11603,N_11662);
or U15580 (N_15580,N_10426,N_11218);
nand U15581 (N_15581,N_11761,N_6750);
and U15582 (N_15582,N_11089,N_11341);
and U15583 (N_15583,N_11213,N_11225);
nand U15584 (N_15584,N_9884,N_6248);
and U15585 (N_15585,N_6595,N_8291);
xnor U15586 (N_15586,N_8484,N_8508);
nor U15587 (N_15587,N_11120,N_6518);
xnor U15588 (N_15588,N_11019,N_11441);
nand U15589 (N_15589,N_7777,N_11215);
or U15590 (N_15590,N_7002,N_7017);
xor U15591 (N_15591,N_6639,N_10197);
and U15592 (N_15592,N_8608,N_9932);
or U15593 (N_15593,N_7485,N_9630);
and U15594 (N_15594,N_9023,N_9906);
nor U15595 (N_15595,N_7249,N_7826);
xnor U15596 (N_15596,N_11876,N_10399);
nor U15597 (N_15597,N_8882,N_7246);
nand U15598 (N_15598,N_11205,N_7561);
and U15599 (N_15599,N_6115,N_6940);
nor U15600 (N_15600,N_6036,N_7103);
nand U15601 (N_15601,N_6001,N_10553);
and U15602 (N_15602,N_10258,N_6141);
and U15603 (N_15603,N_7277,N_11270);
or U15604 (N_15604,N_11969,N_6905);
xor U15605 (N_15605,N_8837,N_9143);
nand U15606 (N_15606,N_10293,N_10152);
nand U15607 (N_15607,N_8006,N_10646);
and U15608 (N_15608,N_8531,N_8686);
nor U15609 (N_15609,N_6975,N_8330);
nand U15610 (N_15610,N_11396,N_10915);
or U15611 (N_15611,N_7951,N_7905);
nor U15612 (N_15612,N_10422,N_7652);
or U15613 (N_15613,N_7494,N_7236);
nand U15614 (N_15614,N_8128,N_10222);
xnor U15615 (N_15615,N_11847,N_9554);
nand U15616 (N_15616,N_6051,N_7580);
nor U15617 (N_15617,N_6142,N_7452);
or U15618 (N_15618,N_9061,N_11731);
or U15619 (N_15619,N_8119,N_11314);
nand U15620 (N_15620,N_8008,N_8741);
or U15621 (N_15621,N_10396,N_8259);
nor U15622 (N_15622,N_11743,N_8514);
and U15623 (N_15623,N_8948,N_11026);
nand U15624 (N_15624,N_9651,N_7938);
nand U15625 (N_15625,N_10231,N_7330);
or U15626 (N_15626,N_6848,N_11244);
or U15627 (N_15627,N_7451,N_6266);
or U15628 (N_15628,N_9905,N_8766);
or U15629 (N_15629,N_6708,N_8527);
xor U15630 (N_15630,N_6944,N_10438);
or U15631 (N_15631,N_7906,N_10445);
xnor U15632 (N_15632,N_8410,N_7105);
nor U15633 (N_15633,N_8715,N_7683);
nor U15634 (N_15634,N_7860,N_10706);
nor U15635 (N_15635,N_6568,N_7136);
nand U15636 (N_15636,N_9439,N_11725);
xnor U15637 (N_15637,N_9848,N_6353);
or U15638 (N_15638,N_10340,N_11600);
or U15639 (N_15639,N_9280,N_10807);
and U15640 (N_15640,N_6606,N_6268);
and U15641 (N_15641,N_6693,N_6153);
or U15642 (N_15642,N_6180,N_10626);
or U15643 (N_15643,N_11652,N_8978);
nand U15644 (N_15644,N_11259,N_6869);
and U15645 (N_15645,N_6967,N_7294);
nand U15646 (N_15646,N_8268,N_11867);
and U15647 (N_15647,N_8028,N_7972);
nand U15648 (N_15648,N_6116,N_8877);
nor U15649 (N_15649,N_6777,N_8618);
nor U15650 (N_15650,N_10088,N_10962);
nand U15651 (N_15651,N_6367,N_6621);
xnor U15652 (N_15652,N_7613,N_7329);
and U15653 (N_15653,N_11035,N_7889);
and U15654 (N_15654,N_6164,N_6130);
and U15655 (N_15655,N_7124,N_7828);
nor U15656 (N_15656,N_8443,N_8241);
nand U15657 (N_15657,N_9624,N_9810);
or U15658 (N_15658,N_10936,N_6827);
or U15659 (N_15659,N_9177,N_9834);
nor U15660 (N_15660,N_9532,N_9011);
xor U15661 (N_15661,N_7560,N_7846);
or U15662 (N_15662,N_10547,N_9042);
nor U15663 (N_15663,N_7888,N_9907);
and U15664 (N_15664,N_7348,N_8194);
xnor U15665 (N_15665,N_7477,N_7679);
xor U15666 (N_15666,N_11236,N_10228);
and U15667 (N_15667,N_6005,N_9241);
nand U15668 (N_15668,N_9938,N_8545);
or U15669 (N_15669,N_9438,N_9804);
nand U15670 (N_15670,N_10161,N_7741);
nand U15671 (N_15671,N_7365,N_8452);
or U15672 (N_15672,N_6840,N_10515);
nand U15673 (N_15673,N_7271,N_9334);
and U15674 (N_15674,N_6302,N_7438);
xnor U15675 (N_15675,N_11277,N_6617);
nor U15676 (N_15676,N_10017,N_6557);
or U15677 (N_15677,N_10978,N_6361);
nand U15678 (N_15678,N_8432,N_10999);
nand U15679 (N_15679,N_9028,N_6317);
xor U15680 (N_15680,N_8621,N_9259);
nand U15681 (N_15681,N_10471,N_10005);
nor U15682 (N_15682,N_8324,N_10466);
and U15683 (N_15683,N_9328,N_10528);
or U15684 (N_15684,N_11256,N_11188);
nor U15685 (N_15685,N_10248,N_10875);
xnor U15686 (N_15686,N_11043,N_9080);
xnor U15687 (N_15687,N_11818,N_7923);
xnor U15688 (N_15688,N_8541,N_11469);
nand U15689 (N_15689,N_6881,N_11624);
and U15690 (N_15690,N_11828,N_9455);
nor U15691 (N_15691,N_6019,N_10601);
xnor U15692 (N_15692,N_8538,N_8755);
xor U15693 (N_15693,N_7908,N_7205);
or U15694 (N_15694,N_9025,N_10750);
xor U15695 (N_15695,N_6995,N_7449);
xnor U15696 (N_15696,N_10680,N_6026);
or U15697 (N_15697,N_10294,N_7233);
xor U15698 (N_15698,N_10513,N_10099);
nand U15699 (N_15699,N_7582,N_11774);
nor U15700 (N_15700,N_9555,N_7957);
or U15701 (N_15701,N_11558,N_10498);
or U15702 (N_15702,N_11844,N_6385);
nor U15703 (N_15703,N_9791,N_8421);
or U15704 (N_15704,N_9748,N_7292);
xor U15705 (N_15705,N_7831,N_7930);
and U15706 (N_15706,N_10385,N_11130);
nor U15707 (N_15707,N_6208,N_8919);
or U15708 (N_15708,N_8515,N_6839);
nand U15709 (N_15709,N_10654,N_10570);
or U15710 (N_15710,N_9321,N_6345);
nand U15711 (N_15711,N_9822,N_8031);
xor U15712 (N_15712,N_9054,N_10062);
nor U15713 (N_15713,N_7060,N_11981);
xor U15714 (N_15714,N_10710,N_11505);
or U15715 (N_15715,N_6292,N_6183);
or U15716 (N_15716,N_6893,N_6056);
and U15717 (N_15717,N_6065,N_11111);
nor U15718 (N_15718,N_11058,N_9656);
nor U15719 (N_15719,N_7744,N_9298);
or U15720 (N_15720,N_11039,N_10394);
nand U15721 (N_15721,N_7630,N_9853);
nand U15722 (N_15722,N_9886,N_10269);
xor U15723 (N_15723,N_9112,N_8713);
or U15724 (N_15724,N_10293,N_6189);
and U15725 (N_15725,N_11615,N_10097);
or U15726 (N_15726,N_11252,N_7767);
or U15727 (N_15727,N_7278,N_11219);
or U15728 (N_15728,N_6635,N_11864);
or U15729 (N_15729,N_6783,N_8014);
or U15730 (N_15730,N_10424,N_9545);
and U15731 (N_15731,N_7384,N_7799);
or U15732 (N_15732,N_8482,N_10155);
and U15733 (N_15733,N_7893,N_8669);
nor U15734 (N_15734,N_7790,N_6222);
nor U15735 (N_15735,N_7063,N_10962);
xor U15736 (N_15736,N_9531,N_6935);
nor U15737 (N_15737,N_11493,N_10252);
or U15738 (N_15738,N_7349,N_10000);
or U15739 (N_15739,N_7611,N_8557);
or U15740 (N_15740,N_9766,N_8781);
xor U15741 (N_15741,N_11149,N_7992);
and U15742 (N_15742,N_7507,N_8480);
xor U15743 (N_15743,N_6492,N_11149);
xor U15744 (N_15744,N_7661,N_7629);
or U15745 (N_15745,N_6877,N_10885);
nor U15746 (N_15746,N_8816,N_9381);
or U15747 (N_15747,N_8823,N_10017);
nand U15748 (N_15748,N_11344,N_10315);
xnor U15749 (N_15749,N_6749,N_11772);
or U15750 (N_15750,N_11701,N_7349);
xor U15751 (N_15751,N_10869,N_7962);
nand U15752 (N_15752,N_6677,N_7443);
nand U15753 (N_15753,N_9639,N_8812);
or U15754 (N_15754,N_11808,N_8424);
nor U15755 (N_15755,N_11860,N_11535);
nand U15756 (N_15756,N_10652,N_10583);
nor U15757 (N_15757,N_6305,N_11948);
and U15758 (N_15758,N_9035,N_8537);
nor U15759 (N_15759,N_7401,N_7282);
xnor U15760 (N_15760,N_6606,N_7232);
nand U15761 (N_15761,N_6611,N_8214);
nor U15762 (N_15762,N_8206,N_7323);
nor U15763 (N_15763,N_9641,N_7014);
nor U15764 (N_15764,N_11028,N_7903);
xor U15765 (N_15765,N_10815,N_9213);
xnor U15766 (N_15766,N_11557,N_10906);
nor U15767 (N_15767,N_11455,N_6530);
or U15768 (N_15768,N_9551,N_7926);
nand U15769 (N_15769,N_10161,N_11324);
xnor U15770 (N_15770,N_10401,N_7274);
nor U15771 (N_15771,N_11662,N_8732);
and U15772 (N_15772,N_10861,N_6737);
and U15773 (N_15773,N_6375,N_8205);
nand U15774 (N_15774,N_11326,N_8913);
nand U15775 (N_15775,N_8418,N_6151);
nor U15776 (N_15776,N_6118,N_8989);
nand U15777 (N_15777,N_10847,N_8414);
nand U15778 (N_15778,N_11698,N_10197);
or U15779 (N_15779,N_6917,N_8032);
nor U15780 (N_15780,N_10736,N_9031);
xor U15781 (N_15781,N_11262,N_11510);
or U15782 (N_15782,N_9893,N_8394);
and U15783 (N_15783,N_11789,N_10858);
or U15784 (N_15784,N_6338,N_9008);
and U15785 (N_15785,N_11343,N_8364);
and U15786 (N_15786,N_8187,N_8226);
and U15787 (N_15787,N_7217,N_7385);
or U15788 (N_15788,N_9801,N_7201);
nor U15789 (N_15789,N_11789,N_10921);
or U15790 (N_15790,N_11961,N_8187);
and U15791 (N_15791,N_11445,N_9307);
nand U15792 (N_15792,N_11151,N_10098);
or U15793 (N_15793,N_9795,N_8234);
nor U15794 (N_15794,N_8552,N_8305);
nor U15795 (N_15795,N_8370,N_10670);
nand U15796 (N_15796,N_9638,N_11073);
nor U15797 (N_15797,N_8739,N_10092);
nand U15798 (N_15798,N_10831,N_8333);
xnor U15799 (N_15799,N_6246,N_8444);
xor U15800 (N_15800,N_6108,N_6726);
or U15801 (N_15801,N_10746,N_11330);
nand U15802 (N_15802,N_9834,N_7355);
or U15803 (N_15803,N_8414,N_6768);
or U15804 (N_15804,N_10009,N_11126);
or U15805 (N_15805,N_10748,N_7588);
nor U15806 (N_15806,N_9290,N_6157);
xnor U15807 (N_15807,N_9390,N_10125);
nor U15808 (N_15808,N_10970,N_6450);
or U15809 (N_15809,N_9119,N_6155);
nor U15810 (N_15810,N_9140,N_8154);
or U15811 (N_15811,N_7021,N_11905);
nor U15812 (N_15812,N_9086,N_11243);
nand U15813 (N_15813,N_10749,N_8319);
nand U15814 (N_15814,N_10789,N_6449);
xnor U15815 (N_15815,N_8311,N_10369);
nor U15816 (N_15816,N_10377,N_7997);
nor U15817 (N_15817,N_9477,N_7095);
and U15818 (N_15818,N_10393,N_6816);
nand U15819 (N_15819,N_11240,N_9993);
and U15820 (N_15820,N_10631,N_11078);
and U15821 (N_15821,N_9682,N_8116);
or U15822 (N_15822,N_10370,N_10328);
nand U15823 (N_15823,N_10789,N_7881);
nand U15824 (N_15824,N_7225,N_8627);
or U15825 (N_15825,N_8817,N_7317);
nand U15826 (N_15826,N_9223,N_11060);
and U15827 (N_15827,N_9594,N_10368);
and U15828 (N_15828,N_6557,N_6726);
xnor U15829 (N_15829,N_8869,N_6261);
nand U15830 (N_15830,N_8380,N_6842);
xnor U15831 (N_15831,N_6975,N_9704);
nand U15832 (N_15832,N_10155,N_6275);
xnor U15833 (N_15833,N_9495,N_10175);
nor U15834 (N_15834,N_8685,N_9282);
xnor U15835 (N_15835,N_9655,N_11549);
and U15836 (N_15836,N_10116,N_9851);
xnor U15837 (N_15837,N_6046,N_7490);
nor U15838 (N_15838,N_7067,N_6156);
nor U15839 (N_15839,N_10039,N_11724);
nor U15840 (N_15840,N_8194,N_8448);
or U15841 (N_15841,N_11878,N_6835);
nor U15842 (N_15842,N_10848,N_10238);
nand U15843 (N_15843,N_7518,N_7774);
and U15844 (N_15844,N_6772,N_8277);
xnor U15845 (N_15845,N_8139,N_9287);
xnor U15846 (N_15846,N_10264,N_8604);
xor U15847 (N_15847,N_10225,N_11971);
nand U15848 (N_15848,N_9825,N_8576);
xor U15849 (N_15849,N_9976,N_6845);
nor U15850 (N_15850,N_8692,N_6575);
and U15851 (N_15851,N_11105,N_6978);
or U15852 (N_15852,N_6546,N_8252);
or U15853 (N_15853,N_11385,N_8047);
or U15854 (N_15854,N_8270,N_6623);
or U15855 (N_15855,N_6671,N_8025);
nand U15856 (N_15856,N_8156,N_11472);
or U15857 (N_15857,N_9550,N_9045);
nor U15858 (N_15858,N_6798,N_10223);
and U15859 (N_15859,N_9654,N_7332);
and U15860 (N_15860,N_11448,N_6718);
and U15861 (N_15861,N_10181,N_10820);
nor U15862 (N_15862,N_9564,N_9456);
or U15863 (N_15863,N_7826,N_11370);
and U15864 (N_15864,N_8716,N_9707);
and U15865 (N_15865,N_10110,N_7406);
xnor U15866 (N_15866,N_8293,N_11994);
and U15867 (N_15867,N_6259,N_10984);
xnor U15868 (N_15868,N_6479,N_8517);
or U15869 (N_15869,N_10642,N_7789);
xnor U15870 (N_15870,N_6563,N_6379);
and U15871 (N_15871,N_9654,N_8688);
nor U15872 (N_15872,N_11981,N_7136);
or U15873 (N_15873,N_10326,N_6644);
nand U15874 (N_15874,N_10644,N_11825);
xor U15875 (N_15875,N_10105,N_11325);
and U15876 (N_15876,N_10971,N_9747);
or U15877 (N_15877,N_6817,N_9285);
xor U15878 (N_15878,N_6640,N_9000);
xor U15879 (N_15879,N_11660,N_8728);
nor U15880 (N_15880,N_10957,N_7829);
nor U15881 (N_15881,N_7341,N_8641);
or U15882 (N_15882,N_6442,N_8832);
nor U15883 (N_15883,N_9833,N_8693);
xnor U15884 (N_15884,N_8552,N_8985);
and U15885 (N_15885,N_7360,N_9213);
xor U15886 (N_15886,N_6567,N_11755);
xnor U15887 (N_15887,N_9508,N_11525);
xor U15888 (N_15888,N_7917,N_9857);
nor U15889 (N_15889,N_10556,N_9574);
nor U15890 (N_15890,N_6248,N_10737);
or U15891 (N_15891,N_8226,N_9663);
and U15892 (N_15892,N_10823,N_10430);
and U15893 (N_15893,N_6344,N_8332);
or U15894 (N_15894,N_8996,N_6316);
and U15895 (N_15895,N_8594,N_7024);
nand U15896 (N_15896,N_6838,N_11831);
nand U15897 (N_15897,N_7426,N_11091);
nor U15898 (N_15898,N_11861,N_8041);
or U15899 (N_15899,N_6530,N_11737);
nor U15900 (N_15900,N_11352,N_11645);
nor U15901 (N_15901,N_8116,N_6204);
xor U15902 (N_15902,N_11806,N_8856);
xor U15903 (N_15903,N_7523,N_6680);
nor U15904 (N_15904,N_8641,N_6556);
or U15905 (N_15905,N_8750,N_10133);
xnor U15906 (N_15906,N_7794,N_10904);
or U15907 (N_15907,N_9300,N_9812);
xor U15908 (N_15908,N_9740,N_9572);
xor U15909 (N_15909,N_11776,N_6985);
or U15910 (N_15910,N_6143,N_7198);
nor U15911 (N_15911,N_9349,N_8869);
or U15912 (N_15912,N_6904,N_11221);
nand U15913 (N_15913,N_11293,N_9235);
xor U15914 (N_15914,N_10819,N_7818);
nor U15915 (N_15915,N_11468,N_10544);
nor U15916 (N_15916,N_11662,N_10442);
or U15917 (N_15917,N_10171,N_10824);
nand U15918 (N_15918,N_11186,N_6900);
and U15919 (N_15919,N_8179,N_11655);
nand U15920 (N_15920,N_6667,N_7441);
or U15921 (N_15921,N_7025,N_11595);
or U15922 (N_15922,N_6265,N_8238);
and U15923 (N_15923,N_11810,N_8601);
nand U15924 (N_15924,N_8212,N_10897);
nand U15925 (N_15925,N_7188,N_11408);
and U15926 (N_15926,N_11549,N_11531);
or U15927 (N_15927,N_7418,N_8899);
nand U15928 (N_15928,N_10520,N_11728);
and U15929 (N_15929,N_11540,N_11834);
xnor U15930 (N_15930,N_8754,N_9293);
xor U15931 (N_15931,N_11476,N_10754);
nand U15932 (N_15932,N_8861,N_7604);
and U15933 (N_15933,N_9963,N_6483);
xnor U15934 (N_15934,N_7659,N_6223);
or U15935 (N_15935,N_11238,N_11344);
and U15936 (N_15936,N_10867,N_7026);
and U15937 (N_15937,N_7495,N_8293);
or U15938 (N_15938,N_8174,N_7290);
xnor U15939 (N_15939,N_9376,N_10562);
and U15940 (N_15940,N_11293,N_7797);
and U15941 (N_15941,N_11557,N_6523);
nand U15942 (N_15942,N_6609,N_9493);
xnor U15943 (N_15943,N_8199,N_6013);
nor U15944 (N_15944,N_8094,N_11505);
nor U15945 (N_15945,N_9656,N_9207);
nand U15946 (N_15946,N_11995,N_9182);
nor U15947 (N_15947,N_6098,N_8982);
nor U15948 (N_15948,N_8778,N_6615);
xor U15949 (N_15949,N_7909,N_9213);
nor U15950 (N_15950,N_9516,N_9751);
or U15951 (N_15951,N_8332,N_11955);
xor U15952 (N_15952,N_7577,N_8033);
or U15953 (N_15953,N_6190,N_7011);
nand U15954 (N_15954,N_11818,N_6836);
nand U15955 (N_15955,N_6595,N_11990);
nor U15956 (N_15956,N_6551,N_6822);
and U15957 (N_15957,N_9191,N_7931);
nor U15958 (N_15958,N_10236,N_8464);
nand U15959 (N_15959,N_7687,N_10697);
nand U15960 (N_15960,N_9383,N_6807);
or U15961 (N_15961,N_10364,N_10060);
and U15962 (N_15962,N_6209,N_7382);
nand U15963 (N_15963,N_8916,N_7837);
and U15964 (N_15964,N_10645,N_11285);
and U15965 (N_15965,N_10452,N_8591);
and U15966 (N_15966,N_7192,N_6470);
and U15967 (N_15967,N_8227,N_11420);
or U15968 (N_15968,N_8964,N_6441);
nor U15969 (N_15969,N_8602,N_7736);
or U15970 (N_15970,N_10832,N_10336);
and U15971 (N_15971,N_7360,N_6302);
nand U15972 (N_15972,N_10294,N_11830);
nor U15973 (N_15973,N_9870,N_8654);
nor U15974 (N_15974,N_8651,N_6029);
or U15975 (N_15975,N_9322,N_7732);
nor U15976 (N_15976,N_6898,N_11346);
nand U15977 (N_15977,N_11784,N_9263);
xnor U15978 (N_15978,N_11441,N_11503);
or U15979 (N_15979,N_6142,N_7219);
nand U15980 (N_15980,N_7515,N_10225);
and U15981 (N_15981,N_11203,N_7701);
or U15982 (N_15982,N_6854,N_11045);
or U15983 (N_15983,N_10968,N_11123);
and U15984 (N_15984,N_7763,N_9546);
nand U15985 (N_15985,N_8094,N_6213);
nor U15986 (N_15986,N_7169,N_8913);
or U15987 (N_15987,N_7883,N_6622);
and U15988 (N_15988,N_8750,N_7973);
nand U15989 (N_15989,N_8272,N_11874);
or U15990 (N_15990,N_7866,N_10216);
nand U15991 (N_15991,N_6226,N_10858);
or U15992 (N_15992,N_8312,N_6460);
and U15993 (N_15993,N_11737,N_8176);
xor U15994 (N_15994,N_10277,N_8026);
xor U15995 (N_15995,N_9200,N_9111);
or U15996 (N_15996,N_8251,N_10289);
and U15997 (N_15997,N_6420,N_8198);
or U15998 (N_15998,N_11522,N_11126);
or U15999 (N_15999,N_11150,N_6863);
and U16000 (N_16000,N_7078,N_11409);
or U16001 (N_16001,N_11097,N_7788);
and U16002 (N_16002,N_9255,N_9079);
nand U16003 (N_16003,N_7101,N_10093);
and U16004 (N_16004,N_8560,N_7741);
xnor U16005 (N_16005,N_10089,N_7625);
and U16006 (N_16006,N_6938,N_8596);
nor U16007 (N_16007,N_9706,N_9129);
nor U16008 (N_16008,N_6000,N_8440);
nand U16009 (N_16009,N_11101,N_11601);
nand U16010 (N_16010,N_6876,N_7114);
and U16011 (N_16011,N_7687,N_10308);
nand U16012 (N_16012,N_7122,N_9046);
nand U16013 (N_16013,N_9656,N_11822);
xnor U16014 (N_16014,N_8419,N_10300);
nand U16015 (N_16015,N_10840,N_8883);
nor U16016 (N_16016,N_8363,N_7636);
or U16017 (N_16017,N_8534,N_9185);
xor U16018 (N_16018,N_8901,N_11644);
xnor U16019 (N_16019,N_10118,N_11856);
nor U16020 (N_16020,N_6191,N_8443);
nand U16021 (N_16021,N_9483,N_7709);
and U16022 (N_16022,N_11784,N_11094);
xor U16023 (N_16023,N_7259,N_11984);
and U16024 (N_16024,N_7326,N_10266);
or U16025 (N_16025,N_9052,N_10997);
xnor U16026 (N_16026,N_6038,N_8395);
nor U16027 (N_16027,N_10362,N_7242);
or U16028 (N_16028,N_9847,N_7270);
nor U16029 (N_16029,N_10553,N_7212);
nor U16030 (N_16030,N_9828,N_8105);
xnor U16031 (N_16031,N_6679,N_11833);
xnor U16032 (N_16032,N_6184,N_9568);
nand U16033 (N_16033,N_9805,N_10982);
nand U16034 (N_16034,N_7816,N_10005);
nand U16035 (N_16035,N_10639,N_8135);
or U16036 (N_16036,N_8434,N_11834);
nand U16037 (N_16037,N_6088,N_11612);
nand U16038 (N_16038,N_11616,N_9774);
nor U16039 (N_16039,N_8864,N_7037);
nand U16040 (N_16040,N_10843,N_7248);
xnor U16041 (N_16041,N_6576,N_10431);
nor U16042 (N_16042,N_7570,N_6402);
nand U16043 (N_16043,N_6190,N_8177);
xor U16044 (N_16044,N_11984,N_11560);
and U16045 (N_16045,N_8244,N_7134);
or U16046 (N_16046,N_9065,N_7497);
nor U16047 (N_16047,N_10009,N_7882);
xor U16048 (N_16048,N_7535,N_6427);
and U16049 (N_16049,N_6400,N_11144);
nor U16050 (N_16050,N_6762,N_8221);
xnor U16051 (N_16051,N_6545,N_9471);
nand U16052 (N_16052,N_11539,N_11446);
xor U16053 (N_16053,N_6735,N_9093);
xor U16054 (N_16054,N_6747,N_7265);
and U16055 (N_16055,N_6270,N_8487);
xnor U16056 (N_16056,N_6231,N_11239);
nand U16057 (N_16057,N_8528,N_8061);
xor U16058 (N_16058,N_11191,N_7627);
xor U16059 (N_16059,N_7167,N_6695);
or U16060 (N_16060,N_6113,N_9474);
xor U16061 (N_16061,N_9986,N_6671);
nor U16062 (N_16062,N_10500,N_10923);
nor U16063 (N_16063,N_6079,N_11917);
nand U16064 (N_16064,N_9111,N_9045);
nand U16065 (N_16065,N_11443,N_7387);
nor U16066 (N_16066,N_10764,N_6511);
or U16067 (N_16067,N_7969,N_6309);
or U16068 (N_16068,N_7253,N_6674);
nor U16069 (N_16069,N_11144,N_8256);
nand U16070 (N_16070,N_10759,N_9198);
and U16071 (N_16071,N_6130,N_6074);
and U16072 (N_16072,N_10650,N_11689);
and U16073 (N_16073,N_9997,N_8738);
xnor U16074 (N_16074,N_9029,N_7045);
nor U16075 (N_16075,N_6583,N_11715);
and U16076 (N_16076,N_8425,N_11989);
or U16077 (N_16077,N_11839,N_10429);
nor U16078 (N_16078,N_9811,N_9116);
xor U16079 (N_16079,N_10954,N_10631);
or U16080 (N_16080,N_8752,N_11468);
and U16081 (N_16081,N_11301,N_9402);
nand U16082 (N_16082,N_6143,N_8835);
xnor U16083 (N_16083,N_8089,N_8020);
and U16084 (N_16084,N_8857,N_8554);
nand U16085 (N_16085,N_7886,N_9436);
nor U16086 (N_16086,N_9138,N_9552);
xor U16087 (N_16087,N_7718,N_7154);
and U16088 (N_16088,N_7161,N_7877);
or U16089 (N_16089,N_9669,N_9386);
or U16090 (N_16090,N_6511,N_9092);
and U16091 (N_16091,N_6995,N_10958);
nor U16092 (N_16092,N_8442,N_8681);
xor U16093 (N_16093,N_8901,N_10627);
and U16094 (N_16094,N_9197,N_8226);
and U16095 (N_16095,N_11318,N_10362);
or U16096 (N_16096,N_11234,N_6815);
xnor U16097 (N_16097,N_6441,N_6221);
xor U16098 (N_16098,N_9680,N_6815);
or U16099 (N_16099,N_8162,N_8664);
nor U16100 (N_16100,N_6083,N_8920);
nand U16101 (N_16101,N_8650,N_10724);
nor U16102 (N_16102,N_6562,N_10192);
xnor U16103 (N_16103,N_10385,N_7331);
or U16104 (N_16104,N_6188,N_9196);
and U16105 (N_16105,N_8012,N_11500);
nand U16106 (N_16106,N_10625,N_7704);
nor U16107 (N_16107,N_10504,N_10547);
and U16108 (N_16108,N_9913,N_9761);
and U16109 (N_16109,N_8641,N_8228);
nand U16110 (N_16110,N_6369,N_6114);
or U16111 (N_16111,N_6297,N_6713);
nand U16112 (N_16112,N_11285,N_10754);
nor U16113 (N_16113,N_9948,N_9618);
nor U16114 (N_16114,N_8182,N_7959);
nand U16115 (N_16115,N_6639,N_9780);
xor U16116 (N_16116,N_11259,N_10604);
xnor U16117 (N_16117,N_6342,N_9743);
nor U16118 (N_16118,N_11325,N_7167);
nand U16119 (N_16119,N_10958,N_7933);
nand U16120 (N_16120,N_9160,N_6002);
nor U16121 (N_16121,N_8742,N_8951);
xnor U16122 (N_16122,N_6730,N_7676);
nand U16123 (N_16123,N_6052,N_10586);
nor U16124 (N_16124,N_7656,N_9691);
or U16125 (N_16125,N_8221,N_9163);
nor U16126 (N_16126,N_10977,N_6786);
nor U16127 (N_16127,N_6071,N_9428);
and U16128 (N_16128,N_10916,N_11727);
nand U16129 (N_16129,N_7653,N_8382);
and U16130 (N_16130,N_6648,N_11130);
xor U16131 (N_16131,N_10528,N_7360);
or U16132 (N_16132,N_8622,N_10057);
and U16133 (N_16133,N_8751,N_11167);
or U16134 (N_16134,N_8851,N_9817);
and U16135 (N_16135,N_9251,N_10334);
nor U16136 (N_16136,N_9691,N_7993);
xnor U16137 (N_16137,N_7537,N_10850);
nor U16138 (N_16138,N_9413,N_8487);
and U16139 (N_16139,N_9477,N_9605);
or U16140 (N_16140,N_10691,N_11565);
nand U16141 (N_16141,N_6699,N_11967);
nor U16142 (N_16142,N_9312,N_7102);
nand U16143 (N_16143,N_8263,N_11392);
and U16144 (N_16144,N_10585,N_8274);
or U16145 (N_16145,N_8684,N_9817);
nor U16146 (N_16146,N_10226,N_11142);
nor U16147 (N_16147,N_8553,N_8078);
xnor U16148 (N_16148,N_9289,N_6430);
nand U16149 (N_16149,N_9636,N_9675);
nand U16150 (N_16150,N_11386,N_8212);
nor U16151 (N_16151,N_9022,N_6578);
nor U16152 (N_16152,N_11039,N_9450);
nand U16153 (N_16153,N_6371,N_9604);
xor U16154 (N_16154,N_10570,N_9539);
and U16155 (N_16155,N_7347,N_9251);
and U16156 (N_16156,N_10642,N_7958);
xnor U16157 (N_16157,N_11331,N_8316);
or U16158 (N_16158,N_9496,N_10874);
nor U16159 (N_16159,N_10652,N_10719);
and U16160 (N_16160,N_9073,N_11461);
nor U16161 (N_16161,N_11243,N_11425);
xor U16162 (N_16162,N_8951,N_6220);
nand U16163 (N_16163,N_9105,N_7131);
nor U16164 (N_16164,N_10317,N_6031);
and U16165 (N_16165,N_7527,N_6444);
and U16166 (N_16166,N_10440,N_6464);
nand U16167 (N_16167,N_7477,N_7680);
nand U16168 (N_16168,N_9645,N_7259);
or U16169 (N_16169,N_8719,N_9299);
xor U16170 (N_16170,N_9929,N_8094);
xnor U16171 (N_16171,N_7464,N_7135);
nor U16172 (N_16172,N_10629,N_8223);
and U16173 (N_16173,N_11015,N_9819);
nand U16174 (N_16174,N_11608,N_9853);
nand U16175 (N_16175,N_11084,N_10108);
nand U16176 (N_16176,N_8561,N_10941);
xor U16177 (N_16177,N_8915,N_8671);
nor U16178 (N_16178,N_11200,N_11163);
and U16179 (N_16179,N_11892,N_6212);
xnor U16180 (N_16180,N_6207,N_9836);
or U16181 (N_16181,N_7148,N_11215);
or U16182 (N_16182,N_6020,N_11272);
and U16183 (N_16183,N_7520,N_6031);
nand U16184 (N_16184,N_8153,N_7682);
xnor U16185 (N_16185,N_10943,N_8677);
or U16186 (N_16186,N_10385,N_7343);
nand U16187 (N_16187,N_10251,N_9865);
nand U16188 (N_16188,N_11761,N_8801);
or U16189 (N_16189,N_11151,N_6465);
xor U16190 (N_16190,N_7849,N_10862);
or U16191 (N_16191,N_6571,N_6748);
and U16192 (N_16192,N_11514,N_11622);
nor U16193 (N_16193,N_10743,N_9187);
or U16194 (N_16194,N_10741,N_11315);
xnor U16195 (N_16195,N_9399,N_10646);
xor U16196 (N_16196,N_8639,N_10164);
nand U16197 (N_16197,N_8868,N_7383);
nor U16198 (N_16198,N_6232,N_11802);
nand U16199 (N_16199,N_7711,N_6393);
nor U16200 (N_16200,N_8855,N_7317);
and U16201 (N_16201,N_8430,N_8774);
or U16202 (N_16202,N_7993,N_10487);
nand U16203 (N_16203,N_10600,N_9643);
nor U16204 (N_16204,N_6286,N_8078);
nand U16205 (N_16205,N_7574,N_9895);
and U16206 (N_16206,N_7506,N_7896);
and U16207 (N_16207,N_10080,N_6015);
and U16208 (N_16208,N_10643,N_7505);
nand U16209 (N_16209,N_7185,N_10057);
nand U16210 (N_16210,N_7762,N_7872);
xnor U16211 (N_16211,N_10056,N_9940);
nor U16212 (N_16212,N_7787,N_6566);
nand U16213 (N_16213,N_9273,N_7084);
xor U16214 (N_16214,N_10592,N_11514);
and U16215 (N_16215,N_7579,N_11884);
and U16216 (N_16216,N_10048,N_8136);
and U16217 (N_16217,N_7393,N_11718);
xnor U16218 (N_16218,N_7576,N_7501);
nor U16219 (N_16219,N_8162,N_7575);
nor U16220 (N_16220,N_8216,N_8821);
nor U16221 (N_16221,N_7220,N_7415);
and U16222 (N_16222,N_6625,N_7116);
and U16223 (N_16223,N_8662,N_8443);
and U16224 (N_16224,N_7051,N_11532);
nand U16225 (N_16225,N_8924,N_11454);
nand U16226 (N_16226,N_10391,N_8579);
or U16227 (N_16227,N_9716,N_10835);
or U16228 (N_16228,N_10899,N_8957);
or U16229 (N_16229,N_8285,N_6533);
and U16230 (N_16230,N_11586,N_11706);
and U16231 (N_16231,N_7300,N_11610);
or U16232 (N_16232,N_10586,N_8679);
xor U16233 (N_16233,N_10329,N_8419);
nor U16234 (N_16234,N_8679,N_6370);
or U16235 (N_16235,N_9273,N_9744);
and U16236 (N_16236,N_8268,N_10893);
or U16237 (N_16237,N_6566,N_8090);
nor U16238 (N_16238,N_7664,N_6458);
or U16239 (N_16239,N_8361,N_10025);
xor U16240 (N_16240,N_6311,N_10186);
nand U16241 (N_16241,N_8066,N_7952);
and U16242 (N_16242,N_11833,N_11505);
and U16243 (N_16243,N_10152,N_8838);
nor U16244 (N_16244,N_6022,N_6310);
and U16245 (N_16245,N_7034,N_8147);
nand U16246 (N_16246,N_8453,N_10475);
nand U16247 (N_16247,N_7848,N_11883);
and U16248 (N_16248,N_6933,N_8031);
or U16249 (N_16249,N_9977,N_8497);
or U16250 (N_16250,N_7141,N_8468);
and U16251 (N_16251,N_7080,N_6972);
or U16252 (N_16252,N_7706,N_6163);
and U16253 (N_16253,N_7148,N_9789);
and U16254 (N_16254,N_11365,N_9929);
and U16255 (N_16255,N_6119,N_9746);
xnor U16256 (N_16256,N_10515,N_8317);
nand U16257 (N_16257,N_10076,N_9458);
or U16258 (N_16258,N_9992,N_7140);
nand U16259 (N_16259,N_10020,N_11478);
and U16260 (N_16260,N_11644,N_7396);
nand U16261 (N_16261,N_11581,N_6565);
nor U16262 (N_16262,N_8911,N_8232);
or U16263 (N_16263,N_7180,N_10075);
nor U16264 (N_16264,N_8119,N_11918);
or U16265 (N_16265,N_11274,N_9027);
nand U16266 (N_16266,N_10768,N_11560);
nor U16267 (N_16267,N_7036,N_9589);
nor U16268 (N_16268,N_9200,N_6587);
or U16269 (N_16269,N_8924,N_10721);
nor U16270 (N_16270,N_9484,N_10223);
nand U16271 (N_16271,N_10764,N_8368);
and U16272 (N_16272,N_11027,N_11147);
or U16273 (N_16273,N_6943,N_10299);
and U16274 (N_16274,N_8736,N_8325);
or U16275 (N_16275,N_7542,N_8835);
nor U16276 (N_16276,N_8311,N_11030);
nor U16277 (N_16277,N_11703,N_6180);
and U16278 (N_16278,N_8616,N_10442);
xor U16279 (N_16279,N_11268,N_11953);
nand U16280 (N_16280,N_11716,N_10952);
nor U16281 (N_16281,N_7622,N_9583);
or U16282 (N_16282,N_10842,N_11797);
and U16283 (N_16283,N_7903,N_7273);
nor U16284 (N_16284,N_7210,N_11490);
or U16285 (N_16285,N_11872,N_10330);
xor U16286 (N_16286,N_10193,N_6958);
nand U16287 (N_16287,N_8665,N_10057);
and U16288 (N_16288,N_8484,N_7734);
xnor U16289 (N_16289,N_7029,N_7731);
xnor U16290 (N_16290,N_7727,N_9048);
nand U16291 (N_16291,N_10423,N_10564);
or U16292 (N_16292,N_9443,N_8711);
nor U16293 (N_16293,N_10433,N_10217);
or U16294 (N_16294,N_8448,N_11448);
nor U16295 (N_16295,N_9255,N_9281);
nand U16296 (N_16296,N_6262,N_7734);
and U16297 (N_16297,N_8500,N_9489);
nand U16298 (N_16298,N_8020,N_9758);
xor U16299 (N_16299,N_9619,N_7794);
nand U16300 (N_16300,N_6890,N_7578);
xnor U16301 (N_16301,N_9181,N_6304);
nand U16302 (N_16302,N_9488,N_6862);
and U16303 (N_16303,N_10520,N_7170);
xor U16304 (N_16304,N_11434,N_10295);
nand U16305 (N_16305,N_7690,N_6112);
nor U16306 (N_16306,N_8221,N_8663);
xor U16307 (N_16307,N_10531,N_11664);
or U16308 (N_16308,N_9139,N_7670);
or U16309 (N_16309,N_6441,N_6466);
nor U16310 (N_16310,N_6297,N_7944);
xnor U16311 (N_16311,N_10664,N_6246);
and U16312 (N_16312,N_8158,N_11591);
nor U16313 (N_16313,N_6357,N_9897);
or U16314 (N_16314,N_9754,N_10500);
nor U16315 (N_16315,N_6132,N_8374);
nand U16316 (N_16316,N_11745,N_8821);
nor U16317 (N_16317,N_11560,N_10787);
xor U16318 (N_16318,N_7831,N_7341);
and U16319 (N_16319,N_6729,N_7172);
or U16320 (N_16320,N_9543,N_6440);
or U16321 (N_16321,N_10061,N_11580);
nand U16322 (N_16322,N_11237,N_11058);
or U16323 (N_16323,N_11878,N_9793);
nand U16324 (N_16324,N_6742,N_11273);
or U16325 (N_16325,N_6193,N_10353);
or U16326 (N_16326,N_7108,N_9958);
and U16327 (N_16327,N_10830,N_9672);
xnor U16328 (N_16328,N_9973,N_11812);
and U16329 (N_16329,N_9623,N_9458);
nand U16330 (N_16330,N_8902,N_8791);
and U16331 (N_16331,N_11181,N_7481);
xnor U16332 (N_16332,N_6449,N_11489);
or U16333 (N_16333,N_9820,N_8216);
or U16334 (N_16334,N_8891,N_10893);
or U16335 (N_16335,N_8742,N_6158);
nor U16336 (N_16336,N_7057,N_11354);
nor U16337 (N_16337,N_9794,N_10397);
and U16338 (N_16338,N_7121,N_9990);
or U16339 (N_16339,N_7694,N_8703);
or U16340 (N_16340,N_7701,N_11358);
nand U16341 (N_16341,N_9627,N_11418);
or U16342 (N_16342,N_7443,N_10054);
nand U16343 (N_16343,N_11317,N_8725);
and U16344 (N_16344,N_7717,N_7107);
xor U16345 (N_16345,N_8779,N_11673);
nand U16346 (N_16346,N_6971,N_10550);
nor U16347 (N_16347,N_10282,N_10131);
and U16348 (N_16348,N_8798,N_7651);
and U16349 (N_16349,N_6927,N_11059);
xnor U16350 (N_16350,N_9220,N_11001);
or U16351 (N_16351,N_7884,N_8746);
xor U16352 (N_16352,N_7412,N_8030);
and U16353 (N_16353,N_11243,N_7729);
and U16354 (N_16354,N_6674,N_10153);
and U16355 (N_16355,N_6544,N_11941);
nand U16356 (N_16356,N_10995,N_7949);
nand U16357 (N_16357,N_7681,N_8803);
xnor U16358 (N_16358,N_7956,N_11594);
and U16359 (N_16359,N_11113,N_8286);
or U16360 (N_16360,N_7438,N_11900);
nor U16361 (N_16361,N_11648,N_7626);
or U16362 (N_16362,N_9136,N_6668);
or U16363 (N_16363,N_6275,N_10359);
nor U16364 (N_16364,N_10094,N_6329);
xor U16365 (N_16365,N_11505,N_9659);
nor U16366 (N_16366,N_8004,N_10547);
nor U16367 (N_16367,N_11698,N_8814);
nor U16368 (N_16368,N_9990,N_7895);
xnor U16369 (N_16369,N_10928,N_8547);
nand U16370 (N_16370,N_10663,N_10089);
xnor U16371 (N_16371,N_7817,N_8440);
and U16372 (N_16372,N_7899,N_9318);
nor U16373 (N_16373,N_10649,N_11461);
nor U16374 (N_16374,N_6076,N_9738);
nor U16375 (N_16375,N_10979,N_9915);
nand U16376 (N_16376,N_10641,N_9705);
nor U16377 (N_16377,N_9528,N_10880);
or U16378 (N_16378,N_6724,N_8672);
xor U16379 (N_16379,N_9693,N_10171);
and U16380 (N_16380,N_7542,N_7505);
or U16381 (N_16381,N_8340,N_6577);
xor U16382 (N_16382,N_11019,N_8808);
xnor U16383 (N_16383,N_11012,N_6708);
xor U16384 (N_16384,N_9375,N_10481);
and U16385 (N_16385,N_8304,N_11041);
nand U16386 (N_16386,N_8310,N_8235);
xnor U16387 (N_16387,N_7123,N_6334);
and U16388 (N_16388,N_6995,N_9236);
nand U16389 (N_16389,N_6093,N_9571);
nor U16390 (N_16390,N_10963,N_10005);
or U16391 (N_16391,N_7758,N_8181);
and U16392 (N_16392,N_11493,N_10158);
nor U16393 (N_16393,N_6976,N_11757);
nand U16394 (N_16394,N_8534,N_11717);
or U16395 (N_16395,N_9710,N_8862);
and U16396 (N_16396,N_7507,N_10354);
nand U16397 (N_16397,N_8659,N_7296);
or U16398 (N_16398,N_8077,N_7013);
xnor U16399 (N_16399,N_6865,N_10613);
nand U16400 (N_16400,N_7129,N_9429);
and U16401 (N_16401,N_6159,N_9681);
nor U16402 (N_16402,N_7043,N_6543);
and U16403 (N_16403,N_6277,N_8680);
and U16404 (N_16404,N_11624,N_8215);
nand U16405 (N_16405,N_7311,N_11344);
nand U16406 (N_16406,N_7006,N_6449);
nor U16407 (N_16407,N_8722,N_9688);
and U16408 (N_16408,N_11783,N_7542);
and U16409 (N_16409,N_9269,N_7291);
or U16410 (N_16410,N_9614,N_7942);
or U16411 (N_16411,N_7930,N_11559);
xnor U16412 (N_16412,N_9380,N_9866);
nand U16413 (N_16413,N_8854,N_6617);
and U16414 (N_16414,N_11746,N_8256);
or U16415 (N_16415,N_10211,N_10401);
nand U16416 (N_16416,N_10814,N_7476);
nor U16417 (N_16417,N_8659,N_10338);
xnor U16418 (N_16418,N_9080,N_11370);
nor U16419 (N_16419,N_11443,N_9315);
nor U16420 (N_16420,N_7575,N_7469);
nor U16421 (N_16421,N_9951,N_6122);
nand U16422 (N_16422,N_7233,N_6202);
or U16423 (N_16423,N_11940,N_6550);
xnor U16424 (N_16424,N_11648,N_11505);
nor U16425 (N_16425,N_7785,N_7960);
nand U16426 (N_16426,N_8171,N_8600);
or U16427 (N_16427,N_8845,N_11267);
nand U16428 (N_16428,N_11383,N_8704);
and U16429 (N_16429,N_8975,N_11140);
and U16430 (N_16430,N_6921,N_8399);
nor U16431 (N_16431,N_11368,N_6651);
xnor U16432 (N_16432,N_9687,N_9387);
xor U16433 (N_16433,N_9718,N_7958);
xor U16434 (N_16434,N_7553,N_8862);
xnor U16435 (N_16435,N_7937,N_10151);
nand U16436 (N_16436,N_8613,N_6643);
nor U16437 (N_16437,N_7268,N_7133);
or U16438 (N_16438,N_9727,N_6270);
nand U16439 (N_16439,N_7152,N_10813);
nor U16440 (N_16440,N_6487,N_7387);
xnor U16441 (N_16441,N_11154,N_8665);
xor U16442 (N_16442,N_7601,N_10542);
nand U16443 (N_16443,N_8727,N_6650);
nor U16444 (N_16444,N_11034,N_8302);
xnor U16445 (N_16445,N_7414,N_11980);
and U16446 (N_16446,N_10551,N_8415);
or U16447 (N_16447,N_6867,N_8485);
nor U16448 (N_16448,N_8268,N_10765);
nand U16449 (N_16449,N_9257,N_11545);
nand U16450 (N_16450,N_11111,N_10868);
xnor U16451 (N_16451,N_6687,N_8207);
nor U16452 (N_16452,N_10436,N_6229);
and U16453 (N_16453,N_10452,N_8618);
nand U16454 (N_16454,N_6435,N_10542);
nor U16455 (N_16455,N_10573,N_11051);
nand U16456 (N_16456,N_10784,N_8079);
xnor U16457 (N_16457,N_9122,N_9431);
nand U16458 (N_16458,N_6614,N_6174);
nand U16459 (N_16459,N_8292,N_8890);
nand U16460 (N_16460,N_8578,N_11714);
or U16461 (N_16461,N_9716,N_8378);
and U16462 (N_16462,N_10344,N_11832);
nor U16463 (N_16463,N_6682,N_6776);
nor U16464 (N_16464,N_6791,N_11896);
or U16465 (N_16465,N_8681,N_8061);
or U16466 (N_16466,N_8457,N_8918);
or U16467 (N_16467,N_6278,N_9849);
nor U16468 (N_16468,N_8043,N_10524);
or U16469 (N_16469,N_9883,N_10089);
or U16470 (N_16470,N_9832,N_10634);
and U16471 (N_16471,N_10050,N_11407);
or U16472 (N_16472,N_6052,N_7055);
nand U16473 (N_16473,N_6449,N_7574);
xnor U16474 (N_16474,N_11912,N_7796);
xnor U16475 (N_16475,N_7299,N_10358);
and U16476 (N_16476,N_11002,N_8670);
nor U16477 (N_16477,N_11454,N_6651);
or U16478 (N_16478,N_10281,N_11333);
nand U16479 (N_16479,N_8297,N_6294);
nor U16480 (N_16480,N_8021,N_10941);
nor U16481 (N_16481,N_10948,N_10287);
or U16482 (N_16482,N_9637,N_9446);
xnor U16483 (N_16483,N_7284,N_6308);
xnor U16484 (N_16484,N_8732,N_11436);
xnor U16485 (N_16485,N_6928,N_11148);
nor U16486 (N_16486,N_9930,N_10442);
xor U16487 (N_16487,N_11463,N_7415);
nand U16488 (N_16488,N_9905,N_10305);
nor U16489 (N_16489,N_9654,N_11393);
and U16490 (N_16490,N_10320,N_11614);
nor U16491 (N_16491,N_8331,N_8587);
or U16492 (N_16492,N_7141,N_9357);
xor U16493 (N_16493,N_6184,N_7582);
xor U16494 (N_16494,N_7107,N_8263);
nand U16495 (N_16495,N_7654,N_11027);
nand U16496 (N_16496,N_8912,N_6176);
or U16497 (N_16497,N_6924,N_9187);
and U16498 (N_16498,N_11821,N_9519);
nand U16499 (N_16499,N_8488,N_6234);
nand U16500 (N_16500,N_7405,N_10584);
nor U16501 (N_16501,N_11805,N_7004);
and U16502 (N_16502,N_8711,N_11709);
nand U16503 (N_16503,N_10261,N_6881);
nand U16504 (N_16504,N_10670,N_8110);
xor U16505 (N_16505,N_6385,N_10073);
xnor U16506 (N_16506,N_8793,N_6837);
or U16507 (N_16507,N_7665,N_9746);
xnor U16508 (N_16508,N_7916,N_11396);
nand U16509 (N_16509,N_8909,N_10218);
nor U16510 (N_16510,N_8040,N_7508);
xnor U16511 (N_16511,N_8309,N_10780);
nor U16512 (N_16512,N_9600,N_10621);
nor U16513 (N_16513,N_10685,N_6229);
and U16514 (N_16514,N_10362,N_8250);
xnor U16515 (N_16515,N_8839,N_9549);
xor U16516 (N_16516,N_7794,N_8090);
nor U16517 (N_16517,N_11884,N_7571);
or U16518 (N_16518,N_8336,N_11642);
nor U16519 (N_16519,N_8162,N_9937);
xor U16520 (N_16520,N_9803,N_8930);
or U16521 (N_16521,N_8310,N_11194);
or U16522 (N_16522,N_8412,N_7225);
xor U16523 (N_16523,N_9475,N_8434);
nor U16524 (N_16524,N_8218,N_11485);
and U16525 (N_16525,N_6629,N_6716);
xor U16526 (N_16526,N_8197,N_7286);
xor U16527 (N_16527,N_6866,N_10325);
and U16528 (N_16528,N_10225,N_7089);
or U16529 (N_16529,N_9321,N_7230);
or U16530 (N_16530,N_7575,N_7167);
nor U16531 (N_16531,N_7887,N_9605);
or U16532 (N_16532,N_9370,N_10778);
nor U16533 (N_16533,N_11791,N_7711);
or U16534 (N_16534,N_7409,N_6984);
nor U16535 (N_16535,N_9389,N_10968);
nor U16536 (N_16536,N_6779,N_9610);
and U16537 (N_16537,N_8799,N_6492);
or U16538 (N_16538,N_9803,N_11395);
nor U16539 (N_16539,N_10435,N_11188);
nor U16540 (N_16540,N_6031,N_6643);
nand U16541 (N_16541,N_10522,N_7760);
xnor U16542 (N_16542,N_10523,N_9261);
nor U16543 (N_16543,N_7591,N_10172);
nor U16544 (N_16544,N_7421,N_9239);
and U16545 (N_16545,N_11306,N_6432);
nor U16546 (N_16546,N_8723,N_11805);
nor U16547 (N_16547,N_8466,N_11933);
nor U16548 (N_16548,N_11496,N_9629);
nand U16549 (N_16549,N_7703,N_11050);
nor U16550 (N_16550,N_7179,N_6306);
and U16551 (N_16551,N_7124,N_10531);
xor U16552 (N_16552,N_8246,N_11580);
nand U16553 (N_16553,N_7813,N_9648);
nor U16554 (N_16554,N_11773,N_7781);
nor U16555 (N_16555,N_11719,N_8113);
xnor U16556 (N_16556,N_8510,N_10976);
nand U16557 (N_16557,N_8412,N_9265);
nand U16558 (N_16558,N_11471,N_8569);
xor U16559 (N_16559,N_8539,N_9731);
and U16560 (N_16560,N_6043,N_8566);
nor U16561 (N_16561,N_8108,N_8986);
nor U16562 (N_16562,N_7075,N_11018);
nor U16563 (N_16563,N_11286,N_8315);
or U16564 (N_16564,N_9222,N_6921);
xnor U16565 (N_16565,N_11171,N_9162);
nor U16566 (N_16566,N_11349,N_10626);
nor U16567 (N_16567,N_9719,N_8063);
xnor U16568 (N_16568,N_7870,N_8317);
nor U16569 (N_16569,N_8829,N_9652);
nand U16570 (N_16570,N_11776,N_9584);
or U16571 (N_16571,N_8531,N_7997);
and U16572 (N_16572,N_8650,N_8899);
nor U16573 (N_16573,N_9315,N_7150);
xor U16574 (N_16574,N_6767,N_6848);
xor U16575 (N_16575,N_7109,N_10288);
nor U16576 (N_16576,N_8378,N_7234);
xnor U16577 (N_16577,N_7078,N_9422);
nor U16578 (N_16578,N_9337,N_6067);
and U16579 (N_16579,N_10703,N_11460);
xnor U16580 (N_16580,N_6357,N_11028);
nand U16581 (N_16581,N_6642,N_7973);
xor U16582 (N_16582,N_11611,N_11667);
xnor U16583 (N_16583,N_10078,N_11632);
xor U16584 (N_16584,N_6677,N_8751);
xnor U16585 (N_16585,N_9354,N_11609);
nand U16586 (N_16586,N_8928,N_8913);
nand U16587 (N_16587,N_10992,N_11547);
or U16588 (N_16588,N_7066,N_7662);
nand U16589 (N_16589,N_6998,N_8213);
xnor U16590 (N_16590,N_7875,N_8558);
nor U16591 (N_16591,N_7349,N_10693);
nand U16592 (N_16592,N_9038,N_8435);
nand U16593 (N_16593,N_6268,N_9520);
nand U16594 (N_16594,N_10685,N_9495);
nand U16595 (N_16595,N_11347,N_8110);
nor U16596 (N_16596,N_11911,N_11632);
or U16597 (N_16597,N_9168,N_7676);
or U16598 (N_16598,N_11873,N_11766);
nor U16599 (N_16599,N_9853,N_6717);
or U16600 (N_16600,N_8180,N_9840);
nor U16601 (N_16601,N_9389,N_8597);
nand U16602 (N_16602,N_10585,N_8076);
and U16603 (N_16603,N_10278,N_9708);
nor U16604 (N_16604,N_11858,N_9433);
xor U16605 (N_16605,N_7527,N_10379);
nand U16606 (N_16606,N_10783,N_6203);
and U16607 (N_16607,N_6147,N_9552);
and U16608 (N_16608,N_11583,N_6891);
or U16609 (N_16609,N_11506,N_11301);
and U16610 (N_16610,N_11124,N_8662);
nand U16611 (N_16611,N_10250,N_11944);
nor U16612 (N_16612,N_8652,N_11481);
nor U16613 (N_16613,N_8205,N_9926);
nand U16614 (N_16614,N_10924,N_6592);
xor U16615 (N_16615,N_10755,N_11413);
and U16616 (N_16616,N_6335,N_8523);
or U16617 (N_16617,N_9166,N_6353);
nand U16618 (N_16618,N_9986,N_9356);
nor U16619 (N_16619,N_11291,N_11964);
nand U16620 (N_16620,N_11459,N_10694);
or U16621 (N_16621,N_7196,N_8478);
nand U16622 (N_16622,N_11210,N_6664);
nand U16623 (N_16623,N_9786,N_6159);
nand U16624 (N_16624,N_6342,N_6351);
or U16625 (N_16625,N_7997,N_7459);
nor U16626 (N_16626,N_9394,N_7509);
and U16627 (N_16627,N_10455,N_7235);
nand U16628 (N_16628,N_8712,N_7971);
xor U16629 (N_16629,N_7531,N_7603);
nand U16630 (N_16630,N_8799,N_7432);
nor U16631 (N_16631,N_6214,N_11467);
nor U16632 (N_16632,N_9277,N_11375);
nand U16633 (N_16633,N_6785,N_8577);
nand U16634 (N_16634,N_9903,N_7118);
and U16635 (N_16635,N_8998,N_9569);
and U16636 (N_16636,N_11831,N_8043);
xnor U16637 (N_16637,N_7410,N_7836);
xor U16638 (N_16638,N_11646,N_9845);
or U16639 (N_16639,N_11026,N_11613);
and U16640 (N_16640,N_11164,N_11705);
or U16641 (N_16641,N_11355,N_7763);
nor U16642 (N_16642,N_8026,N_6162);
nand U16643 (N_16643,N_10655,N_11192);
xnor U16644 (N_16644,N_6935,N_8907);
or U16645 (N_16645,N_6560,N_11383);
and U16646 (N_16646,N_11461,N_10701);
nor U16647 (N_16647,N_8936,N_6017);
xnor U16648 (N_16648,N_8128,N_8071);
xnor U16649 (N_16649,N_11849,N_11441);
xor U16650 (N_16650,N_7268,N_6820);
or U16651 (N_16651,N_7770,N_6554);
or U16652 (N_16652,N_11840,N_6932);
and U16653 (N_16653,N_9641,N_9468);
nor U16654 (N_16654,N_11517,N_9536);
and U16655 (N_16655,N_7774,N_8815);
and U16656 (N_16656,N_9182,N_6727);
nor U16657 (N_16657,N_11159,N_8621);
and U16658 (N_16658,N_7958,N_7108);
or U16659 (N_16659,N_7355,N_9011);
or U16660 (N_16660,N_10150,N_7905);
nand U16661 (N_16661,N_8942,N_8614);
and U16662 (N_16662,N_9291,N_10697);
xor U16663 (N_16663,N_11625,N_7279);
or U16664 (N_16664,N_11914,N_11612);
nor U16665 (N_16665,N_11708,N_8084);
and U16666 (N_16666,N_11816,N_7367);
and U16667 (N_16667,N_7245,N_9113);
xor U16668 (N_16668,N_6927,N_6333);
xor U16669 (N_16669,N_7813,N_7085);
or U16670 (N_16670,N_9921,N_10093);
and U16671 (N_16671,N_8478,N_7377);
nand U16672 (N_16672,N_8248,N_9426);
or U16673 (N_16673,N_11228,N_6329);
nor U16674 (N_16674,N_9569,N_6422);
or U16675 (N_16675,N_11678,N_8477);
or U16676 (N_16676,N_10962,N_11533);
and U16677 (N_16677,N_8039,N_10934);
xnor U16678 (N_16678,N_9735,N_11979);
or U16679 (N_16679,N_9152,N_11447);
or U16680 (N_16680,N_10765,N_10184);
and U16681 (N_16681,N_8869,N_11038);
nand U16682 (N_16682,N_6856,N_9448);
nand U16683 (N_16683,N_8261,N_7555);
xnor U16684 (N_16684,N_7030,N_6736);
xnor U16685 (N_16685,N_11649,N_6910);
xor U16686 (N_16686,N_8475,N_10216);
xnor U16687 (N_16687,N_6185,N_6241);
and U16688 (N_16688,N_7126,N_10827);
nand U16689 (N_16689,N_10491,N_9048);
or U16690 (N_16690,N_8431,N_11794);
nand U16691 (N_16691,N_7093,N_7330);
nor U16692 (N_16692,N_10962,N_7940);
and U16693 (N_16693,N_6082,N_6644);
xor U16694 (N_16694,N_10816,N_10761);
or U16695 (N_16695,N_7645,N_6270);
nand U16696 (N_16696,N_10943,N_11716);
xor U16697 (N_16697,N_11087,N_7089);
nor U16698 (N_16698,N_11297,N_9644);
and U16699 (N_16699,N_10774,N_6834);
or U16700 (N_16700,N_9540,N_11601);
nand U16701 (N_16701,N_6735,N_6964);
nor U16702 (N_16702,N_7802,N_7919);
and U16703 (N_16703,N_10561,N_8502);
xnor U16704 (N_16704,N_8501,N_7144);
and U16705 (N_16705,N_11780,N_8676);
xnor U16706 (N_16706,N_7693,N_8167);
nor U16707 (N_16707,N_7724,N_6295);
nand U16708 (N_16708,N_7457,N_8252);
or U16709 (N_16709,N_7039,N_9710);
nor U16710 (N_16710,N_7293,N_10002);
or U16711 (N_16711,N_9348,N_7967);
or U16712 (N_16712,N_6242,N_6335);
nor U16713 (N_16713,N_6776,N_11515);
nor U16714 (N_16714,N_6313,N_10150);
or U16715 (N_16715,N_10949,N_6633);
and U16716 (N_16716,N_6983,N_9354);
and U16717 (N_16717,N_6837,N_10537);
nand U16718 (N_16718,N_10591,N_7855);
or U16719 (N_16719,N_10929,N_11944);
xor U16720 (N_16720,N_8084,N_8071);
or U16721 (N_16721,N_10937,N_10189);
nor U16722 (N_16722,N_7777,N_6542);
xnor U16723 (N_16723,N_11911,N_6653);
nor U16724 (N_16724,N_11681,N_6018);
nand U16725 (N_16725,N_6179,N_8390);
nor U16726 (N_16726,N_8561,N_8269);
and U16727 (N_16727,N_11985,N_10833);
nor U16728 (N_16728,N_8710,N_10662);
xor U16729 (N_16729,N_8819,N_8256);
and U16730 (N_16730,N_8324,N_6152);
xnor U16731 (N_16731,N_8423,N_8943);
and U16732 (N_16732,N_8664,N_6754);
nor U16733 (N_16733,N_9644,N_8326);
xnor U16734 (N_16734,N_7588,N_9391);
nor U16735 (N_16735,N_10089,N_10595);
nor U16736 (N_16736,N_8383,N_8637);
nand U16737 (N_16737,N_11982,N_6824);
nand U16738 (N_16738,N_6332,N_7707);
or U16739 (N_16739,N_11999,N_10737);
nor U16740 (N_16740,N_7994,N_6572);
or U16741 (N_16741,N_6546,N_7065);
or U16742 (N_16742,N_6114,N_11477);
nand U16743 (N_16743,N_8135,N_11776);
xnor U16744 (N_16744,N_9570,N_6952);
xor U16745 (N_16745,N_6583,N_11497);
xnor U16746 (N_16746,N_6647,N_8474);
xor U16747 (N_16747,N_6032,N_9900);
nor U16748 (N_16748,N_8580,N_8188);
xor U16749 (N_16749,N_10882,N_11449);
xnor U16750 (N_16750,N_10175,N_7794);
or U16751 (N_16751,N_11146,N_8158);
and U16752 (N_16752,N_9538,N_8425);
or U16753 (N_16753,N_6225,N_8261);
xor U16754 (N_16754,N_11983,N_9076);
or U16755 (N_16755,N_6967,N_6621);
or U16756 (N_16756,N_8065,N_9549);
nor U16757 (N_16757,N_6295,N_7880);
or U16758 (N_16758,N_7230,N_6541);
and U16759 (N_16759,N_9217,N_7080);
xor U16760 (N_16760,N_10635,N_6391);
or U16761 (N_16761,N_6005,N_6891);
and U16762 (N_16762,N_6427,N_10943);
nand U16763 (N_16763,N_8834,N_9385);
and U16764 (N_16764,N_7443,N_7940);
and U16765 (N_16765,N_11197,N_7814);
xor U16766 (N_16766,N_8059,N_10704);
nand U16767 (N_16767,N_10550,N_6941);
nor U16768 (N_16768,N_6076,N_6058);
nor U16769 (N_16769,N_6852,N_7978);
or U16770 (N_16770,N_9305,N_9584);
and U16771 (N_16771,N_9499,N_8989);
nand U16772 (N_16772,N_7536,N_7260);
xor U16773 (N_16773,N_9856,N_8592);
and U16774 (N_16774,N_6193,N_6884);
nand U16775 (N_16775,N_6061,N_6202);
xor U16776 (N_16776,N_8251,N_9770);
nor U16777 (N_16777,N_6846,N_11717);
nand U16778 (N_16778,N_9190,N_6821);
xor U16779 (N_16779,N_10858,N_7979);
nand U16780 (N_16780,N_7338,N_8936);
xnor U16781 (N_16781,N_7538,N_9767);
or U16782 (N_16782,N_10559,N_7545);
nor U16783 (N_16783,N_8377,N_8112);
xor U16784 (N_16784,N_10408,N_7414);
or U16785 (N_16785,N_7258,N_8220);
nor U16786 (N_16786,N_9840,N_8924);
nor U16787 (N_16787,N_10929,N_9543);
xnor U16788 (N_16788,N_9320,N_10049);
or U16789 (N_16789,N_10733,N_7895);
xor U16790 (N_16790,N_8770,N_8885);
xnor U16791 (N_16791,N_10027,N_6837);
and U16792 (N_16792,N_8238,N_7305);
xor U16793 (N_16793,N_9693,N_7455);
nor U16794 (N_16794,N_10503,N_6730);
nand U16795 (N_16795,N_8629,N_7468);
and U16796 (N_16796,N_10566,N_7004);
or U16797 (N_16797,N_9895,N_10264);
and U16798 (N_16798,N_8846,N_9086);
or U16799 (N_16799,N_7284,N_7244);
nand U16800 (N_16800,N_10270,N_9350);
or U16801 (N_16801,N_8412,N_8798);
nor U16802 (N_16802,N_7999,N_11928);
and U16803 (N_16803,N_11847,N_6989);
and U16804 (N_16804,N_8197,N_9284);
nand U16805 (N_16805,N_11324,N_7152);
nor U16806 (N_16806,N_6293,N_8673);
nand U16807 (N_16807,N_8898,N_9244);
xnor U16808 (N_16808,N_10634,N_7326);
or U16809 (N_16809,N_7419,N_7046);
xor U16810 (N_16810,N_8887,N_6319);
and U16811 (N_16811,N_6623,N_6852);
and U16812 (N_16812,N_8410,N_7693);
or U16813 (N_16813,N_11515,N_8914);
and U16814 (N_16814,N_7322,N_9601);
nor U16815 (N_16815,N_11353,N_11619);
and U16816 (N_16816,N_10706,N_8611);
nand U16817 (N_16817,N_10901,N_7861);
and U16818 (N_16818,N_9987,N_8150);
nand U16819 (N_16819,N_8661,N_7918);
or U16820 (N_16820,N_7151,N_6279);
and U16821 (N_16821,N_11227,N_10869);
nand U16822 (N_16822,N_10872,N_6343);
nand U16823 (N_16823,N_6762,N_11450);
xor U16824 (N_16824,N_6659,N_7865);
and U16825 (N_16825,N_11416,N_8912);
or U16826 (N_16826,N_8226,N_10625);
nor U16827 (N_16827,N_8589,N_10044);
xor U16828 (N_16828,N_9811,N_8009);
nor U16829 (N_16829,N_10822,N_11230);
xor U16830 (N_16830,N_10794,N_6822);
xor U16831 (N_16831,N_7957,N_10052);
and U16832 (N_16832,N_11888,N_10203);
or U16833 (N_16833,N_8425,N_8993);
nand U16834 (N_16834,N_11364,N_7981);
nor U16835 (N_16835,N_7354,N_7765);
and U16836 (N_16836,N_8836,N_11285);
nand U16837 (N_16837,N_11689,N_10804);
or U16838 (N_16838,N_7450,N_11813);
xor U16839 (N_16839,N_9021,N_7765);
or U16840 (N_16840,N_6658,N_11846);
or U16841 (N_16841,N_10714,N_6664);
xor U16842 (N_16842,N_7403,N_6655);
and U16843 (N_16843,N_6917,N_8057);
nor U16844 (N_16844,N_7010,N_7980);
or U16845 (N_16845,N_6318,N_11826);
xor U16846 (N_16846,N_11844,N_11246);
nand U16847 (N_16847,N_11391,N_10717);
and U16848 (N_16848,N_7912,N_9007);
xor U16849 (N_16849,N_8655,N_10343);
or U16850 (N_16850,N_6016,N_7834);
nand U16851 (N_16851,N_10437,N_11511);
and U16852 (N_16852,N_6204,N_10414);
and U16853 (N_16853,N_6239,N_9011);
xnor U16854 (N_16854,N_10989,N_11596);
xnor U16855 (N_16855,N_11821,N_6387);
nor U16856 (N_16856,N_9442,N_8121);
or U16857 (N_16857,N_10794,N_6194);
nand U16858 (N_16858,N_7314,N_9164);
and U16859 (N_16859,N_8081,N_9943);
and U16860 (N_16860,N_9891,N_10759);
xnor U16861 (N_16861,N_6076,N_7483);
or U16862 (N_16862,N_8459,N_10116);
nand U16863 (N_16863,N_11877,N_8364);
and U16864 (N_16864,N_8012,N_8292);
and U16865 (N_16865,N_7349,N_6204);
nand U16866 (N_16866,N_10182,N_9520);
or U16867 (N_16867,N_9085,N_8344);
nand U16868 (N_16868,N_8406,N_9484);
and U16869 (N_16869,N_8921,N_10983);
or U16870 (N_16870,N_6477,N_9285);
nor U16871 (N_16871,N_9826,N_9427);
nand U16872 (N_16872,N_11373,N_7113);
xnor U16873 (N_16873,N_11011,N_8328);
nand U16874 (N_16874,N_9764,N_11881);
xnor U16875 (N_16875,N_6793,N_10084);
nand U16876 (N_16876,N_9961,N_9497);
xnor U16877 (N_16877,N_10604,N_6619);
and U16878 (N_16878,N_6696,N_9113);
nor U16879 (N_16879,N_7616,N_11940);
nor U16880 (N_16880,N_11759,N_8301);
and U16881 (N_16881,N_11349,N_11866);
nor U16882 (N_16882,N_6855,N_6085);
nor U16883 (N_16883,N_9647,N_11937);
nor U16884 (N_16884,N_7063,N_9991);
or U16885 (N_16885,N_8070,N_6993);
and U16886 (N_16886,N_9801,N_7296);
or U16887 (N_16887,N_8037,N_6181);
nand U16888 (N_16888,N_9710,N_7395);
or U16889 (N_16889,N_9828,N_6873);
and U16890 (N_16890,N_8162,N_9019);
nor U16891 (N_16891,N_7066,N_6613);
nor U16892 (N_16892,N_7154,N_6279);
and U16893 (N_16893,N_6566,N_8907);
or U16894 (N_16894,N_9118,N_11913);
nor U16895 (N_16895,N_6079,N_11585);
and U16896 (N_16896,N_10925,N_6805);
or U16897 (N_16897,N_10375,N_9633);
nand U16898 (N_16898,N_6235,N_6895);
or U16899 (N_16899,N_6523,N_11585);
nand U16900 (N_16900,N_9822,N_6397);
nor U16901 (N_16901,N_8800,N_9241);
nand U16902 (N_16902,N_11716,N_9517);
or U16903 (N_16903,N_9887,N_11362);
and U16904 (N_16904,N_6378,N_8167);
xnor U16905 (N_16905,N_8578,N_7078);
or U16906 (N_16906,N_8822,N_10025);
and U16907 (N_16907,N_6042,N_9432);
xnor U16908 (N_16908,N_6370,N_7872);
and U16909 (N_16909,N_7751,N_11166);
xnor U16910 (N_16910,N_8100,N_8435);
nor U16911 (N_16911,N_8664,N_11879);
and U16912 (N_16912,N_10473,N_7679);
or U16913 (N_16913,N_10045,N_10180);
nand U16914 (N_16914,N_8841,N_7926);
nand U16915 (N_16915,N_8225,N_11925);
nor U16916 (N_16916,N_7075,N_8147);
and U16917 (N_16917,N_7238,N_9517);
nand U16918 (N_16918,N_8255,N_10485);
and U16919 (N_16919,N_10341,N_10346);
and U16920 (N_16920,N_6030,N_11534);
or U16921 (N_16921,N_10502,N_6035);
nor U16922 (N_16922,N_11932,N_11955);
or U16923 (N_16923,N_11259,N_6811);
xnor U16924 (N_16924,N_7649,N_11332);
or U16925 (N_16925,N_9510,N_6970);
or U16926 (N_16926,N_11630,N_7373);
and U16927 (N_16927,N_10973,N_11894);
or U16928 (N_16928,N_10337,N_10074);
and U16929 (N_16929,N_8144,N_9775);
xor U16930 (N_16930,N_9960,N_6069);
or U16931 (N_16931,N_6717,N_6533);
or U16932 (N_16932,N_11085,N_6687);
and U16933 (N_16933,N_7461,N_10102);
nand U16934 (N_16934,N_10775,N_7157);
or U16935 (N_16935,N_11714,N_8617);
nand U16936 (N_16936,N_7534,N_9281);
and U16937 (N_16937,N_7703,N_11499);
nor U16938 (N_16938,N_10379,N_9452);
nor U16939 (N_16939,N_7914,N_8085);
and U16940 (N_16940,N_11313,N_8030);
xnor U16941 (N_16941,N_6302,N_6770);
and U16942 (N_16942,N_8595,N_8395);
nand U16943 (N_16943,N_9222,N_11789);
nand U16944 (N_16944,N_9879,N_7918);
and U16945 (N_16945,N_9123,N_11140);
and U16946 (N_16946,N_6312,N_11992);
xor U16947 (N_16947,N_8775,N_11368);
and U16948 (N_16948,N_10776,N_10827);
and U16949 (N_16949,N_6029,N_10119);
or U16950 (N_16950,N_8723,N_7288);
or U16951 (N_16951,N_10119,N_6927);
xnor U16952 (N_16952,N_9327,N_10909);
and U16953 (N_16953,N_10553,N_11317);
nand U16954 (N_16954,N_10604,N_8401);
nor U16955 (N_16955,N_8621,N_8755);
nor U16956 (N_16956,N_9051,N_7999);
nor U16957 (N_16957,N_9915,N_8479);
xor U16958 (N_16958,N_10508,N_6284);
or U16959 (N_16959,N_6983,N_11341);
xnor U16960 (N_16960,N_8492,N_10141);
nand U16961 (N_16961,N_7057,N_7221);
or U16962 (N_16962,N_10960,N_9470);
or U16963 (N_16963,N_10624,N_6135);
and U16964 (N_16964,N_8330,N_8486);
xnor U16965 (N_16965,N_9011,N_7917);
nor U16966 (N_16966,N_6143,N_6167);
nor U16967 (N_16967,N_8451,N_6329);
nand U16968 (N_16968,N_7752,N_10974);
or U16969 (N_16969,N_6858,N_11344);
nor U16970 (N_16970,N_10092,N_8285);
nand U16971 (N_16971,N_9019,N_6604);
and U16972 (N_16972,N_11716,N_11807);
xor U16973 (N_16973,N_7670,N_9426);
nor U16974 (N_16974,N_9023,N_9875);
or U16975 (N_16975,N_11687,N_8982);
xor U16976 (N_16976,N_11169,N_10620);
and U16977 (N_16977,N_10968,N_8890);
nor U16978 (N_16978,N_8880,N_8372);
xnor U16979 (N_16979,N_7367,N_10512);
xor U16980 (N_16980,N_6721,N_9797);
xor U16981 (N_16981,N_6223,N_10138);
nor U16982 (N_16982,N_6692,N_10644);
or U16983 (N_16983,N_11811,N_9655);
nor U16984 (N_16984,N_7511,N_9073);
or U16985 (N_16985,N_10024,N_6597);
and U16986 (N_16986,N_8656,N_8397);
and U16987 (N_16987,N_10810,N_9489);
nor U16988 (N_16988,N_8924,N_8570);
or U16989 (N_16989,N_11328,N_10351);
or U16990 (N_16990,N_6623,N_8279);
or U16991 (N_16991,N_11024,N_7707);
and U16992 (N_16992,N_9250,N_8399);
nor U16993 (N_16993,N_8627,N_8254);
or U16994 (N_16994,N_7519,N_6829);
or U16995 (N_16995,N_10513,N_8437);
and U16996 (N_16996,N_6138,N_8895);
nor U16997 (N_16997,N_8380,N_8666);
and U16998 (N_16998,N_7946,N_6359);
nor U16999 (N_16999,N_11552,N_11323);
xor U17000 (N_17000,N_7296,N_8421);
and U17001 (N_17001,N_10248,N_6485);
nand U17002 (N_17002,N_8820,N_9105);
nand U17003 (N_17003,N_6405,N_11785);
or U17004 (N_17004,N_6801,N_6960);
nand U17005 (N_17005,N_8301,N_8854);
and U17006 (N_17006,N_11632,N_8475);
nor U17007 (N_17007,N_9723,N_9129);
and U17008 (N_17008,N_6945,N_11034);
or U17009 (N_17009,N_10348,N_8169);
or U17010 (N_17010,N_8284,N_9035);
or U17011 (N_17011,N_11463,N_8564);
xnor U17012 (N_17012,N_11637,N_6527);
and U17013 (N_17013,N_9386,N_6438);
and U17014 (N_17014,N_7717,N_7200);
xor U17015 (N_17015,N_11798,N_6320);
and U17016 (N_17016,N_7417,N_6958);
or U17017 (N_17017,N_7527,N_7638);
and U17018 (N_17018,N_8306,N_7829);
nand U17019 (N_17019,N_10685,N_11982);
nand U17020 (N_17020,N_6414,N_11128);
and U17021 (N_17021,N_11788,N_8041);
nand U17022 (N_17022,N_11414,N_6139);
or U17023 (N_17023,N_7077,N_10218);
nand U17024 (N_17024,N_7721,N_7533);
xnor U17025 (N_17025,N_7474,N_10630);
nand U17026 (N_17026,N_11203,N_7762);
nor U17027 (N_17027,N_10694,N_6429);
xnor U17028 (N_17028,N_7180,N_8024);
nor U17029 (N_17029,N_9260,N_8037);
nor U17030 (N_17030,N_7689,N_10055);
or U17031 (N_17031,N_6617,N_8078);
and U17032 (N_17032,N_6944,N_8060);
nand U17033 (N_17033,N_9208,N_7202);
nand U17034 (N_17034,N_10536,N_10272);
nand U17035 (N_17035,N_6072,N_8254);
nand U17036 (N_17036,N_11039,N_7934);
or U17037 (N_17037,N_7583,N_7401);
or U17038 (N_17038,N_8413,N_7406);
and U17039 (N_17039,N_9119,N_6615);
xnor U17040 (N_17040,N_11178,N_7190);
and U17041 (N_17041,N_6318,N_7802);
or U17042 (N_17042,N_6673,N_11996);
and U17043 (N_17043,N_11781,N_8537);
nand U17044 (N_17044,N_10544,N_11527);
or U17045 (N_17045,N_10089,N_9129);
nand U17046 (N_17046,N_9198,N_11173);
nand U17047 (N_17047,N_9473,N_10411);
nor U17048 (N_17048,N_11227,N_8708);
nor U17049 (N_17049,N_6754,N_9787);
or U17050 (N_17050,N_9292,N_8700);
and U17051 (N_17051,N_6703,N_9643);
and U17052 (N_17052,N_7562,N_6810);
nand U17053 (N_17053,N_9093,N_6606);
nor U17054 (N_17054,N_6290,N_11266);
or U17055 (N_17055,N_6212,N_10464);
nor U17056 (N_17056,N_6332,N_10039);
nor U17057 (N_17057,N_8136,N_6915);
and U17058 (N_17058,N_7239,N_7835);
and U17059 (N_17059,N_6986,N_6400);
xnor U17060 (N_17060,N_11457,N_8388);
xnor U17061 (N_17061,N_10581,N_6622);
and U17062 (N_17062,N_9812,N_7100);
and U17063 (N_17063,N_6408,N_11387);
xnor U17064 (N_17064,N_11246,N_7897);
nand U17065 (N_17065,N_9945,N_11868);
nand U17066 (N_17066,N_10549,N_10078);
nor U17067 (N_17067,N_7865,N_10851);
and U17068 (N_17068,N_7203,N_6632);
nor U17069 (N_17069,N_7222,N_10473);
nor U17070 (N_17070,N_6132,N_6910);
and U17071 (N_17071,N_7027,N_11434);
xor U17072 (N_17072,N_7995,N_6505);
and U17073 (N_17073,N_8980,N_8894);
and U17074 (N_17074,N_6523,N_10525);
nor U17075 (N_17075,N_11810,N_11387);
or U17076 (N_17076,N_11418,N_11106);
nand U17077 (N_17077,N_6278,N_7803);
nor U17078 (N_17078,N_8786,N_11703);
xor U17079 (N_17079,N_10263,N_11675);
nor U17080 (N_17080,N_6350,N_8038);
nor U17081 (N_17081,N_7912,N_10413);
nand U17082 (N_17082,N_8511,N_6831);
or U17083 (N_17083,N_8254,N_7649);
xor U17084 (N_17084,N_9054,N_8751);
or U17085 (N_17085,N_7626,N_10679);
and U17086 (N_17086,N_7209,N_9027);
nor U17087 (N_17087,N_11126,N_11547);
and U17088 (N_17088,N_6129,N_8356);
or U17089 (N_17089,N_6023,N_10597);
and U17090 (N_17090,N_6385,N_8781);
nor U17091 (N_17091,N_6992,N_11661);
and U17092 (N_17092,N_7396,N_11922);
xnor U17093 (N_17093,N_9816,N_6637);
nor U17094 (N_17094,N_8529,N_10650);
nand U17095 (N_17095,N_11109,N_11355);
nor U17096 (N_17096,N_8449,N_8427);
or U17097 (N_17097,N_11713,N_10859);
xor U17098 (N_17098,N_11014,N_6690);
xor U17099 (N_17099,N_11300,N_11709);
or U17100 (N_17100,N_9030,N_7850);
or U17101 (N_17101,N_8221,N_9292);
nor U17102 (N_17102,N_6956,N_6190);
and U17103 (N_17103,N_7074,N_10323);
nand U17104 (N_17104,N_7393,N_10366);
nand U17105 (N_17105,N_6465,N_9957);
xnor U17106 (N_17106,N_10730,N_11383);
or U17107 (N_17107,N_11467,N_8145);
xor U17108 (N_17108,N_9580,N_10329);
or U17109 (N_17109,N_7101,N_6480);
nor U17110 (N_17110,N_10900,N_7965);
nor U17111 (N_17111,N_10087,N_8652);
or U17112 (N_17112,N_8727,N_6030);
and U17113 (N_17113,N_7581,N_8830);
or U17114 (N_17114,N_9647,N_7996);
nand U17115 (N_17115,N_8046,N_6206);
nor U17116 (N_17116,N_11385,N_9394);
nand U17117 (N_17117,N_8948,N_11874);
nand U17118 (N_17118,N_9180,N_11172);
nor U17119 (N_17119,N_10660,N_10488);
nor U17120 (N_17120,N_6581,N_9097);
nor U17121 (N_17121,N_6766,N_11712);
xnor U17122 (N_17122,N_6399,N_10734);
xnor U17123 (N_17123,N_9239,N_9478);
or U17124 (N_17124,N_9822,N_9654);
and U17125 (N_17125,N_8679,N_10863);
xor U17126 (N_17126,N_6106,N_11568);
xnor U17127 (N_17127,N_9304,N_7889);
nor U17128 (N_17128,N_9018,N_6035);
nand U17129 (N_17129,N_10159,N_9671);
nand U17130 (N_17130,N_9845,N_9621);
xor U17131 (N_17131,N_8423,N_11869);
nor U17132 (N_17132,N_6057,N_11946);
nor U17133 (N_17133,N_7966,N_9385);
nand U17134 (N_17134,N_10920,N_7006);
or U17135 (N_17135,N_7972,N_6120);
xor U17136 (N_17136,N_10067,N_9175);
nand U17137 (N_17137,N_6067,N_9071);
nor U17138 (N_17138,N_9501,N_8051);
xnor U17139 (N_17139,N_6547,N_10012);
nand U17140 (N_17140,N_6756,N_11997);
nand U17141 (N_17141,N_8232,N_11012);
nor U17142 (N_17142,N_6983,N_7367);
nand U17143 (N_17143,N_10537,N_8154);
or U17144 (N_17144,N_11460,N_6214);
or U17145 (N_17145,N_11194,N_9617);
or U17146 (N_17146,N_7063,N_8024);
nor U17147 (N_17147,N_6941,N_10466);
nand U17148 (N_17148,N_10425,N_7237);
or U17149 (N_17149,N_8823,N_10549);
nor U17150 (N_17150,N_10322,N_10730);
nor U17151 (N_17151,N_8912,N_6299);
or U17152 (N_17152,N_9150,N_11415);
nand U17153 (N_17153,N_8349,N_9603);
or U17154 (N_17154,N_9274,N_11839);
or U17155 (N_17155,N_7044,N_10574);
or U17156 (N_17156,N_10732,N_11424);
nor U17157 (N_17157,N_8545,N_11735);
xor U17158 (N_17158,N_8234,N_11077);
and U17159 (N_17159,N_10347,N_11707);
xor U17160 (N_17160,N_8273,N_8466);
nand U17161 (N_17161,N_11735,N_7738);
and U17162 (N_17162,N_7479,N_8378);
or U17163 (N_17163,N_6245,N_7713);
nand U17164 (N_17164,N_7124,N_8685);
or U17165 (N_17165,N_9740,N_9594);
xor U17166 (N_17166,N_10232,N_9077);
nand U17167 (N_17167,N_11857,N_11331);
xnor U17168 (N_17168,N_10409,N_8086);
or U17169 (N_17169,N_9263,N_10241);
nand U17170 (N_17170,N_9242,N_9081);
nor U17171 (N_17171,N_9019,N_10657);
or U17172 (N_17172,N_6356,N_6690);
or U17173 (N_17173,N_6856,N_8656);
or U17174 (N_17174,N_7648,N_7292);
or U17175 (N_17175,N_8670,N_6771);
or U17176 (N_17176,N_8933,N_11584);
or U17177 (N_17177,N_6985,N_11386);
nand U17178 (N_17178,N_6747,N_9032);
nor U17179 (N_17179,N_10076,N_11684);
nor U17180 (N_17180,N_11962,N_7331);
and U17181 (N_17181,N_11954,N_7817);
nor U17182 (N_17182,N_11958,N_7557);
nand U17183 (N_17183,N_10012,N_8183);
or U17184 (N_17184,N_10190,N_6387);
or U17185 (N_17185,N_7260,N_8975);
and U17186 (N_17186,N_11218,N_11336);
and U17187 (N_17187,N_7625,N_8064);
xnor U17188 (N_17188,N_7660,N_8263);
and U17189 (N_17189,N_8579,N_6105);
and U17190 (N_17190,N_7747,N_7326);
nor U17191 (N_17191,N_7627,N_10793);
and U17192 (N_17192,N_8670,N_11059);
or U17193 (N_17193,N_9822,N_10235);
or U17194 (N_17194,N_7584,N_9645);
and U17195 (N_17195,N_9666,N_11231);
or U17196 (N_17196,N_10798,N_10099);
xor U17197 (N_17197,N_6872,N_10633);
or U17198 (N_17198,N_7209,N_9097);
xor U17199 (N_17199,N_7662,N_10735);
xnor U17200 (N_17200,N_9154,N_8160);
xor U17201 (N_17201,N_11560,N_7054);
xnor U17202 (N_17202,N_7494,N_7248);
or U17203 (N_17203,N_10656,N_7230);
or U17204 (N_17204,N_7051,N_9079);
and U17205 (N_17205,N_7097,N_6012);
xor U17206 (N_17206,N_9372,N_8590);
nor U17207 (N_17207,N_9396,N_7603);
xnor U17208 (N_17208,N_11531,N_9725);
and U17209 (N_17209,N_6407,N_6964);
nor U17210 (N_17210,N_8244,N_10131);
and U17211 (N_17211,N_9991,N_6891);
and U17212 (N_17212,N_10086,N_10206);
nor U17213 (N_17213,N_7876,N_7440);
xnor U17214 (N_17214,N_10553,N_7131);
or U17215 (N_17215,N_10454,N_11457);
nand U17216 (N_17216,N_11253,N_8005);
nor U17217 (N_17217,N_9668,N_9930);
nor U17218 (N_17218,N_7477,N_9355);
nor U17219 (N_17219,N_9517,N_7485);
nor U17220 (N_17220,N_6028,N_6184);
xnor U17221 (N_17221,N_8438,N_6403);
xnor U17222 (N_17222,N_10735,N_8592);
xnor U17223 (N_17223,N_10532,N_6972);
nand U17224 (N_17224,N_11907,N_7602);
nand U17225 (N_17225,N_10879,N_7238);
nand U17226 (N_17226,N_11899,N_11994);
nor U17227 (N_17227,N_7472,N_10853);
xnor U17228 (N_17228,N_8991,N_10096);
nand U17229 (N_17229,N_9312,N_9937);
and U17230 (N_17230,N_8341,N_7522);
nor U17231 (N_17231,N_8373,N_11263);
nor U17232 (N_17232,N_11977,N_9541);
xnor U17233 (N_17233,N_6526,N_8706);
and U17234 (N_17234,N_11686,N_7437);
or U17235 (N_17235,N_9103,N_8504);
or U17236 (N_17236,N_11623,N_7305);
xnor U17237 (N_17237,N_6169,N_7317);
nand U17238 (N_17238,N_10724,N_8893);
nand U17239 (N_17239,N_8495,N_10978);
nand U17240 (N_17240,N_8290,N_7175);
or U17241 (N_17241,N_7326,N_8590);
xnor U17242 (N_17242,N_9286,N_11491);
nor U17243 (N_17243,N_7005,N_9595);
xnor U17244 (N_17244,N_8436,N_8107);
nand U17245 (N_17245,N_7364,N_7551);
or U17246 (N_17246,N_8912,N_7072);
nor U17247 (N_17247,N_11195,N_6172);
nor U17248 (N_17248,N_11409,N_11449);
or U17249 (N_17249,N_11813,N_6192);
nor U17250 (N_17250,N_9598,N_11964);
and U17251 (N_17251,N_6513,N_6915);
or U17252 (N_17252,N_10451,N_11089);
or U17253 (N_17253,N_6397,N_8308);
xor U17254 (N_17254,N_9233,N_10410);
or U17255 (N_17255,N_9927,N_8339);
xnor U17256 (N_17256,N_10091,N_6866);
or U17257 (N_17257,N_7119,N_11265);
xnor U17258 (N_17258,N_11270,N_11003);
and U17259 (N_17259,N_7203,N_8507);
xor U17260 (N_17260,N_11766,N_11922);
xnor U17261 (N_17261,N_6635,N_11524);
and U17262 (N_17262,N_6509,N_8909);
xor U17263 (N_17263,N_9809,N_6860);
nand U17264 (N_17264,N_9696,N_6334);
and U17265 (N_17265,N_6850,N_7473);
xnor U17266 (N_17266,N_8211,N_8664);
xnor U17267 (N_17267,N_7851,N_7774);
or U17268 (N_17268,N_9285,N_9835);
nor U17269 (N_17269,N_8497,N_10937);
and U17270 (N_17270,N_11754,N_10915);
nor U17271 (N_17271,N_9675,N_6577);
nor U17272 (N_17272,N_6141,N_10932);
nand U17273 (N_17273,N_9502,N_7572);
xnor U17274 (N_17274,N_7118,N_8031);
nand U17275 (N_17275,N_6443,N_10253);
xnor U17276 (N_17276,N_6732,N_8463);
nand U17277 (N_17277,N_11414,N_8855);
nand U17278 (N_17278,N_8593,N_7581);
nor U17279 (N_17279,N_8356,N_7084);
or U17280 (N_17280,N_10972,N_6732);
or U17281 (N_17281,N_6658,N_10370);
or U17282 (N_17282,N_10712,N_10083);
or U17283 (N_17283,N_11936,N_6415);
xor U17284 (N_17284,N_10580,N_9049);
or U17285 (N_17285,N_8907,N_6262);
and U17286 (N_17286,N_9901,N_10555);
nand U17287 (N_17287,N_7727,N_6647);
nor U17288 (N_17288,N_7718,N_11745);
or U17289 (N_17289,N_11023,N_10265);
or U17290 (N_17290,N_11760,N_8297);
and U17291 (N_17291,N_10031,N_10549);
and U17292 (N_17292,N_7378,N_9912);
nand U17293 (N_17293,N_10992,N_8627);
nand U17294 (N_17294,N_11251,N_9050);
nor U17295 (N_17295,N_9790,N_9527);
or U17296 (N_17296,N_11104,N_6877);
and U17297 (N_17297,N_8718,N_8523);
or U17298 (N_17298,N_10485,N_11228);
nand U17299 (N_17299,N_11053,N_11536);
and U17300 (N_17300,N_9011,N_11832);
nor U17301 (N_17301,N_6852,N_11816);
or U17302 (N_17302,N_7244,N_6494);
or U17303 (N_17303,N_11365,N_11317);
and U17304 (N_17304,N_7395,N_11606);
xor U17305 (N_17305,N_11123,N_10053);
or U17306 (N_17306,N_6469,N_6712);
xor U17307 (N_17307,N_7443,N_6108);
nor U17308 (N_17308,N_8739,N_8251);
nand U17309 (N_17309,N_7602,N_7710);
or U17310 (N_17310,N_7513,N_11869);
nand U17311 (N_17311,N_9054,N_10015);
nand U17312 (N_17312,N_6128,N_6310);
xor U17313 (N_17313,N_8325,N_10667);
or U17314 (N_17314,N_8764,N_9380);
xnor U17315 (N_17315,N_7135,N_11359);
nand U17316 (N_17316,N_11032,N_10935);
and U17317 (N_17317,N_7473,N_10348);
nor U17318 (N_17318,N_7391,N_10224);
nor U17319 (N_17319,N_7278,N_8720);
xor U17320 (N_17320,N_9104,N_7034);
nor U17321 (N_17321,N_9806,N_9609);
or U17322 (N_17322,N_7405,N_11361);
xnor U17323 (N_17323,N_7890,N_9929);
or U17324 (N_17324,N_7257,N_10302);
xor U17325 (N_17325,N_10916,N_9797);
and U17326 (N_17326,N_6493,N_6698);
and U17327 (N_17327,N_10325,N_11691);
and U17328 (N_17328,N_6438,N_8703);
or U17329 (N_17329,N_6551,N_6736);
or U17330 (N_17330,N_7825,N_6353);
xor U17331 (N_17331,N_8604,N_11552);
nor U17332 (N_17332,N_9672,N_8602);
and U17333 (N_17333,N_6596,N_6374);
xor U17334 (N_17334,N_11639,N_9219);
nand U17335 (N_17335,N_9510,N_6372);
xor U17336 (N_17336,N_9807,N_9810);
xor U17337 (N_17337,N_7154,N_11397);
nor U17338 (N_17338,N_8170,N_10812);
and U17339 (N_17339,N_11342,N_9172);
nand U17340 (N_17340,N_7421,N_6928);
nor U17341 (N_17341,N_8013,N_6630);
and U17342 (N_17342,N_10680,N_11289);
or U17343 (N_17343,N_10415,N_8447);
or U17344 (N_17344,N_7497,N_6168);
nor U17345 (N_17345,N_10564,N_7126);
nor U17346 (N_17346,N_9250,N_11761);
xnor U17347 (N_17347,N_7506,N_10345);
nor U17348 (N_17348,N_8999,N_6584);
nand U17349 (N_17349,N_7611,N_10215);
xnor U17350 (N_17350,N_9529,N_8921);
nor U17351 (N_17351,N_11966,N_11146);
xnor U17352 (N_17352,N_9680,N_9484);
xor U17353 (N_17353,N_9179,N_11629);
nand U17354 (N_17354,N_11811,N_9090);
nor U17355 (N_17355,N_9620,N_8039);
or U17356 (N_17356,N_9047,N_9481);
or U17357 (N_17357,N_6825,N_9025);
or U17358 (N_17358,N_7136,N_8722);
nor U17359 (N_17359,N_6522,N_8295);
nand U17360 (N_17360,N_7027,N_10256);
nand U17361 (N_17361,N_10175,N_6777);
nor U17362 (N_17362,N_8264,N_9884);
nor U17363 (N_17363,N_7541,N_6757);
or U17364 (N_17364,N_6709,N_6877);
and U17365 (N_17365,N_8851,N_6528);
nor U17366 (N_17366,N_6883,N_10560);
nor U17367 (N_17367,N_7101,N_6513);
and U17368 (N_17368,N_8234,N_11666);
or U17369 (N_17369,N_7335,N_11110);
xnor U17370 (N_17370,N_10170,N_9951);
and U17371 (N_17371,N_11987,N_8272);
and U17372 (N_17372,N_6085,N_9618);
and U17373 (N_17373,N_7638,N_9092);
nand U17374 (N_17374,N_8229,N_8951);
or U17375 (N_17375,N_10324,N_8404);
or U17376 (N_17376,N_9067,N_10505);
xor U17377 (N_17377,N_6303,N_11985);
nor U17378 (N_17378,N_8793,N_9184);
or U17379 (N_17379,N_8896,N_7052);
and U17380 (N_17380,N_7473,N_10577);
xnor U17381 (N_17381,N_7104,N_8277);
nor U17382 (N_17382,N_8131,N_8281);
or U17383 (N_17383,N_10249,N_8254);
nor U17384 (N_17384,N_6272,N_10889);
or U17385 (N_17385,N_6634,N_10163);
or U17386 (N_17386,N_7104,N_7722);
xor U17387 (N_17387,N_7012,N_11953);
nand U17388 (N_17388,N_7883,N_7233);
and U17389 (N_17389,N_9078,N_8857);
or U17390 (N_17390,N_11927,N_10299);
and U17391 (N_17391,N_7070,N_7743);
xor U17392 (N_17392,N_7073,N_11713);
nand U17393 (N_17393,N_7597,N_8075);
or U17394 (N_17394,N_11115,N_11638);
nand U17395 (N_17395,N_6236,N_9362);
nand U17396 (N_17396,N_7010,N_7537);
and U17397 (N_17397,N_11375,N_9595);
and U17398 (N_17398,N_8662,N_8314);
nand U17399 (N_17399,N_9494,N_7221);
nor U17400 (N_17400,N_6749,N_10576);
xor U17401 (N_17401,N_10130,N_7131);
and U17402 (N_17402,N_8623,N_10346);
or U17403 (N_17403,N_9343,N_10796);
nand U17404 (N_17404,N_8005,N_8280);
or U17405 (N_17405,N_10728,N_6853);
or U17406 (N_17406,N_9812,N_8635);
or U17407 (N_17407,N_6342,N_7249);
or U17408 (N_17408,N_10176,N_10679);
or U17409 (N_17409,N_9844,N_8055);
nor U17410 (N_17410,N_6328,N_9300);
or U17411 (N_17411,N_7954,N_10205);
xnor U17412 (N_17412,N_7072,N_11592);
or U17413 (N_17413,N_11306,N_11541);
or U17414 (N_17414,N_8108,N_10492);
xor U17415 (N_17415,N_10137,N_9859);
or U17416 (N_17416,N_9623,N_11848);
or U17417 (N_17417,N_7508,N_11270);
and U17418 (N_17418,N_10639,N_9727);
nor U17419 (N_17419,N_11875,N_11302);
nand U17420 (N_17420,N_10152,N_6194);
nor U17421 (N_17421,N_9586,N_9832);
and U17422 (N_17422,N_7127,N_6099);
nand U17423 (N_17423,N_8938,N_11689);
xnor U17424 (N_17424,N_6219,N_7602);
and U17425 (N_17425,N_8584,N_11839);
nor U17426 (N_17426,N_10846,N_10678);
or U17427 (N_17427,N_11818,N_7875);
and U17428 (N_17428,N_11904,N_10676);
nor U17429 (N_17429,N_9023,N_8733);
and U17430 (N_17430,N_9194,N_8630);
or U17431 (N_17431,N_7204,N_11215);
nor U17432 (N_17432,N_10186,N_7480);
and U17433 (N_17433,N_10173,N_6190);
nor U17434 (N_17434,N_7508,N_6240);
and U17435 (N_17435,N_11733,N_9589);
and U17436 (N_17436,N_11891,N_10008);
and U17437 (N_17437,N_6940,N_9891);
or U17438 (N_17438,N_7302,N_11087);
nand U17439 (N_17439,N_9829,N_6433);
xor U17440 (N_17440,N_10747,N_7912);
nor U17441 (N_17441,N_7616,N_10904);
or U17442 (N_17442,N_6075,N_6493);
or U17443 (N_17443,N_11155,N_10822);
nand U17444 (N_17444,N_8586,N_10154);
xnor U17445 (N_17445,N_11542,N_11055);
xnor U17446 (N_17446,N_10865,N_6384);
nor U17447 (N_17447,N_6954,N_10437);
nor U17448 (N_17448,N_10350,N_9247);
xor U17449 (N_17449,N_11503,N_6503);
nand U17450 (N_17450,N_7823,N_11442);
xnor U17451 (N_17451,N_9043,N_6166);
xor U17452 (N_17452,N_9979,N_11325);
or U17453 (N_17453,N_7447,N_8666);
xor U17454 (N_17454,N_9355,N_8040);
nand U17455 (N_17455,N_6654,N_8741);
and U17456 (N_17456,N_8922,N_6200);
xnor U17457 (N_17457,N_8458,N_6344);
or U17458 (N_17458,N_11713,N_6392);
nand U17459 (N_17459,N_8203,N_7133);
or U17460 (N_17460,N_7916,N_10645);
xor U17461 (N_17461,N_8174,N_7781);
and U17462 (N_17462,N_10240,N_10942);
and U17463 (N_17463,N_11947,N_9348);
nor U17464 (N_17464,N_9670,N_8537);
nor U17465 (N_17465,N_10618,N_7451);
nor U17466 (N_17466,N_9802,N_6258);
nand U17467 (N_17467,N_10253,N_7135);
and U17468 (N_17468,N_7113,N_9134);
or U17469 (N_17469,N_11756,N_8603);
xnor U17470 (N_17470,N_10927,N_11698);
and U17471 (N_17471,N_10341,N_9768);
nor U17472 (N_17472,N_6503,N_9264);
nor U17473 (N_17473,N_10846,N_10628);
xor U17474 (N_17474,N_7138,N_7659);
or U17475 (N_17475,N_8955,N_6873);
or U17476 (N_17476,N_8330,N_6591);
nand U17477 (N_17477,N_8425,N_6751);
xor U17478 (N_17478,N_7473,N_7338);
xnor U17479 (N_17479,N_10235,N_8813);
nand U17480 (N_17480,N_9467,N_10698);
and U17481 (N_17481,N_6482,N_7617);
or U17482 (N_17482,N_10998,N_6436);
nor U17483 (N_17483,N_11340,N_10153);
or U17484 (N_17484,N_9112,N_9436);
nor U17485 (N_17485,N_6265,N_6917);
nor U17486 (N_17486,N_6236,N_8564);
nor U17487 (N_17487,N_11781,N_8119);
and U17488 (N_17488,N_6394,N_10457);
and U17489 (N_17489,N_11084,N_6034);
or U17490 (N_17490,N_11455,N_11915);
nor U17491 (N_17491,N_11511,N_6203);
nand U17492 (N_17492,N_7546,N_6432);
nor U17493 (N_17493,N_6789,N_8469);
xnor U17494 (N_17494,N_11758,N_9891);
nor U17495 (N_17495,N_7976,N_10225);
or U17496 (N_17496,N_6621,N_7632);
xnor U17497 (N_17497,N_9249,N_6892);
xor U17498 (N_17498,N_6856,N_11259);
xor U17499 (N_17499,N_7021,N_7430);
and U17500 (N_17500,N_10967,N_11210);
xnor U17501 (N_17501,N_11083,N_8074);
and U17502 (N_17502,N_6942,N_9569);
xnor U17503 (N_17503,N_6090,N_8190);
nand U17504 (N_17504,N_11790,N_8399);
nor U17505 (N_17505,N_7375,N_9482);
and U17506 (N_17506,N_11885,N_6297);
xnor U17507 (N_17507,N_6376,N_7034);
xor U17508 (N_17508,N_7375,N_9174);
nor U17509 (N_17509,N_7774,N_6359);
xnor U17510 (N_17510,N_9002,N_7990);
or U17511 (N_17511,N_11428,N_6447);
xnor U17512 (N_17512,N_6231,N_9289);
xnor U17513 (N_17513,N_10189,N_9612);
nor U17514 (N_17514,N_6402,N_6592);
nand U17515 (N_17515,N_9916,N_8855);
or U17516 (N_17516,N_8415,N_8852);
xnor U17517 (N_17517,N_11447,N_11761);
or U17518 (N_17518,N_10510,N_11186);
nor U17519 (N_17519,N_11332,N_9099);
and U17520 (N_17520,N_9355,N_11329);
and U17521 (N_17521,N_7199,N_8706);
xor U17522 (N_17522,N_10486,N_6965);
and U17523 (N_17523,N_10404,N_6644);
nor U17524 (N_17524,N_10136,N_9783);
and U17525 (N_17525,N_11923,N_10205);
and U17526 (N_17526,N_10138,N_9571);
or U17527 (N_17527,N_6689,N_10451);
nor U17528 (N_17528,N_8611,N_8820);
xor U17529 (N_17529,N_8844,N_10593);
nor U17530 (N_17530,N_10495,N_6188);
and U17531 (N_17531,N_10674,N_9930);
xnor U17532 (N_17532,N_7180,N_7072);
xor U17533 (N_17533,N_6165,N_8864);
and U17534 (N_17534,N_7344,N_7877);
xor U17535 (N_17535,N_7734,N_11048);
or U17536 (N_17536,N_8978,N_8516);
xor U17537 (N_17537,N_11551,N_10517);
and U17538 (N_17538,N_6144,N_7053);
nor U17539 (N_17539,N_8616,N_6992);
and U17540 (N_17540,N_11022,N_9250);
nor U17541 (N_17541,N_9694,N_7934);
or U17542 (N_17542,N_11039,N_7850);
and U17543 (N_17543,N_6071,N_10791);
nor U17544 (N_17544,N_11058,N_11225);
xor U17545 (N_17545,N_8090,N_10110);
or U17546 (N_17546,N_9662,N_7683);
and U17547 (N_17547,N_10641,N_9269);
or U17548 (N_17548,N_11833,N_10125);
xor U17549 (N_17549,N_6260,N_9293);
xor U17550 (N_17550,N_7995,N_9956);
or U17551 (N_17551,N_8853,N_9229);
or U17552 (N_17552,N_6186,N_10657);
nor U17553 (N_17553,N_7336,N_11917);
or U17554 (N_17554,N_8308,N_9803);
nand U17555 (N_17555,N_8651,N_9531);
and U17556 (N_17556,N_11619,N_7468);
nor U17557 (N_17557,N_11889,N_6115);
or U17558 (N_17558,N_7407,N_11087);
or U17559 (N_17559,N_10129,N_10996);
nand U17560 (N_17560,N_10445,N_9754);
nand U17561 (N_17561,N_6493,N_7473);
nand U17562 (N_17562,N_7636,N_11430);
xnor U17563 (N_17563,N_9838,N_9670);
or U17564 (N_17564,N_10293,N_6752);
nor U17565 (N_17565,N_11799,N_9535);
nand U17566 (N_17566,N_7118,N_9792);
xor U17567 (N_17567,N_8653,N_7124);
nand U17568 (N_17568,N_7711,N_9218);
and U17569 (N_17569,N_6225,N_7253);
nor U17570 (N_17570,N_6066,N_10567);
xnor U17571 (N_17571,N_6183,N_6665);
and U17572 (N_17572,N_11465,N_8122);
nand U17573 (N_17573,N_6071,N_9371);
nor U17574 (N_17574,N_11042,N_7072);
nor U17575 (N_17575,N_7910,N_9345);
xor U17576 (N_17576,N_9691,N_8801);
and U17577 (N_17577,N_9071,N_10425);
nand U17578 (N_17578,N_8826,N_10326);
and U17579 (N_17579,N_8696,N_10469);
nor U17580 (N_17580,N_11727,N_11524);
xnor U17581 (N_17581,N_6541,N_10796);
and U17582 (N_17582,N_8354,N_7209);
and U17583 (N_17583,N_11586,N_8518);
xnor U17584 (N_17584,N_11152,N_11586);
xnor U17585 (N_17585,N_11629,N_7960);
or U17586 (N_17586,N_7826,N_9438);
or U17587 (N_17587,N_6079,N_7840);
or U17588 (N_17588,N_8850,N_6308);
nand U17589 (N_17589,N_8302,N_9910);
nand U17590 (N_17590,N_8103,N_7323);
or U17591 (N_17591,N_9194,N_6204);
nor U17592 (N_17592,N_6959,N_7186);
nor U17593 (N_17593,N_6962,N_7447);
nand U17594 (N_17594,N_9754,N_8175);
nor U17595 (N_17595,N_6602,N_7298);
nand U17596 (N_17596,N_6277,N_8415);
nand U17597 (N_17597,N_6438,N_8912);
nor U17598 (N_17598,N_10546,N_10066);
nand U17599 (N_17599,N_9493,N_11603);
nor U17600 (N_17600,N_6545,N_7100);
nor U17601 (N_17601,N_6533,N_6844);
nand U17602 (N_17602,N_10546,N_9878);
nor U17603 (N_17603,N_7817,N_8984);
xor U17604 (N_17604,N_11400,N_10828);
nor U17605 (N_17605,N_6487,N_10332);
nand U17606 (N_17606,N_9086,N_11995);
and U17607 (N_17607,N_6496,N_8854);
or U17608 (N_17608,N_9494,N_11249);
and U17609 (N_17609,N_11584,N_11235);
and U17610 (N_17610,N_10792,N_11056);
xnor U17611 (N_17611,N_6108,N_8342);
nor U17612 (N_17612,N_11626,N_9412);
nor U17613 (N_17613,N_11923,N_10765);
and U17614 (N_17614,N_9013,N_6567);
nand U17615 (N_17615,N_10788,N_8493);
xnor U17616 (N_17616,N_9097,N_11040);
nor U17617 (N_17617,N_6325,N_7327);
and U17618 (N_17618,N_10978,N_7938);
xor U17619 (N_17619,N_10655,N_7489);
xor U17620 (N_17620,N_11053,N_10711);
and U17621 (N_17621,N_8599,N_8347);
xor U17622 (N_17622,N_10518,N_8840);
nor U17623 (N_17623,N_8135,N_11273);
and U17624 (N_17624,N_6273,N_9999);
and U17625 (N_17625,N_10613,N_7640);
nor U17626 (N_17626,N_11969,N_9264);
xor U17627 (N_17627,N_7100,N_8560);
and U17628 (N_17628,N_11372,N_6210);
xnor U17629 (N_17629,N_9316,N_6990);
or U17630 (N_17630,N_8138,N_11908);
nand U17631 (N_17631,N_6045,N_9001);
and U17632 (N_17632,N_6225,N_6258);
nor U17633 (N_17633,N_9752,N_10908);
nand U17634 (N_17634,N_8212,N_8942);
and U17635 (N_17635,N_7277,N_7748);
and U17636 (N_17636,N_6900,N_10564);
or U17637 (N_17637,N_6604,N_8319);
or U17638 (N_17638,N_6685,N_7454);
xnor U17639 (N_17639,N_9125,N_8534);
and U17640 (N_17640,N_9097,N_11768);
xnor U17641 (N_17641,N_6217,N_8660);
xor U17642 (N_17642,N_11219,N_8220);
xnor U17643 (N_17643,N_9855,N_7932);
and U17644 (N_17644,N_7825,N_11463);
or U17645 (N_17645,N_10229,N_9003);
and U17646 (N_17646,N_6589,N_9245);
or U17647 (N_17647,N_9943,N_7961);
or U17648 (N_17648,N_11820,N_6390);
or U17649 (N_17649,N_9029,N_6335);
nor U17650 (N_17650,N_10294,N_11199);
or U17651 (N_17651,N_8947,N_7078);
nand U17652 (N_17652,N_8648,N_8926);
nor U17653 (N_17653,N_11934,N_6449);
xnor U17654 (N_17654,N_10903,N_8843);
xnor U17655 (N_17655,N_11089,N_7561);
nand U17656 (N_17656,N_11904,N_11885);
and U17657 (N_17657,N_9964,N_8369);
nor U17658 (N_17658,N_9490,N_11612);
nand U17659 (N_17659,N_11075,N_7883);
xor U17660 (N_17660,N_11428,N_8920);
xnor U17661 (N_17661,N_10415,N_6991);
and U17662 (N_17662,N_9585,N_11627);
nor U17663 (N_17663,N_6595,N_11766);
or U17664 (N_17664,N_6157,N_6239);
nand U17665 (N_17665,N_11106,N_9295);
xnor U17666 (N_17666,N_10560,N_11755);
nand U17667 (N_17667,N_8114,N_9579);
and U17668 (N_17668,N_7295,N_11756);
and U17669 (N_17669,N_7821,N_7830);
or U17670 (N_17670,N_7874,N_7391);
and U17671 (N_17671,N_8798,N_7134);
nand U17672 (N_17672,N_9285,N_7719);
nand U17673 (N_17673,N_8592,N_7721);
xnor U17674 (N_17674,N_6224,N_11492);
nor U17675 (N_17675,N_9462,N_10168);
nand U17676 (N_17676,N_7821,N_6642);
or U17677 (N_17677,N_11472,N_6952);
or U17678 (N_17678,N_8337,N_6297);
or U17679 (N_17679,N_10849,N_9740);
or U17680 (N_17680,N_10168,N_9437);
nand U17681 (N_17681,N_8751,N_10109);
or U17682 (N_17682,N_11720,N_7383);
or U17683 (N_17683,N_9688,N_10991);
or U17684 (N_17684,N_6971,N_10828);
or U17685 (N_17685,N_7858,N_8784);
and U17686 (N_17686,N_7102,N_8113);
xnor U17687 (N_17687,N_6711,N_10649);
nor U17688 (N_17688,N_6254,N_7940);
nand U17689 (N_17689,N_7796,N_6720);
or U17690 (N_17690,N_6384,N_10511);
or U17691 (N_17691,N_10249,N_8351);
xnor U17692 (N_17692,N_6510,N_11024);
nor U17693 (N_17693,N_6637,N_6461);
or U17694 (N_17694,N_11741,N_7694);
and U17695 (N_17695,N_11687,N_6200);
and U17696 (N_17696,N_6757,N_10009);
or U17697 (N_17697,N_7208,N_10501);
nand U17698 (N_17698,N_11807,N_8233);
xnor U17699 (N_17699,N_6559,N_7315);
and U17700 (N_17700,N_7332,N_9358);
xnor U17701 (N_17701,N_8373,N_10776);
and U17702 (N_17702,N_7293,N_9661);
nand U17703 (N_17703,N_7235,N_11333);
and U17704 (N_17704,N_6377,N_8727);
and U17705 (N_17705,N_10048,N_11798);
xnor U17706 (N_17706,N_10396,N_6717);
nand U17707 (N_17707,N_8543,N_6448);
nor U17708 (N_17708,N_8448,N_7866);
xnor U17709 (N_17709,N_7334,N_7842);
nand U17710 (N_17710,N_6200,N_6074);
nand U17711 (N_17711,N_6085,N_8875);
xor U17712 (N_17712,N_6548,N_11456);
or U17713 (N_17713,N_9046,N_6373);
nor U17714 (N_17714,N_9427,N_11925);
nor U17715 (N_17715,N_7075,N_7309);
nand U17716 (N_17716,N_9330,N_8566);
or U17717 (N_17717,N_6526,N_10159);
nand U17718 (N_17718,N_8423,N_10650);
and U17719 (N_17719,N_6642,N_10684);
and U17720 (N_17720,N_6277,N_9031);
or U17721 (N_17721,N_7193,N_9563);
nor U17722 (N_17722,N_11752,N_10589);
or U17723 (N_17723,N_7297,N_10516);
xnor U17724 (N_17724,N_10736,N_11192);
or U17725 (N_17725,N_6636,N_7860);
and U17726 (N_17726,N_6753,N_9613);
nor U17727 (N_17727,N_9288,N_7400);
nand U17728 (N_17728,N_10586,N_10364);
or U17729 (N_17729,N_11286,N_10384);
and U17730 (N_17730,N_11197,N_8882);
and U17731 (N_17731,N_11652,N_8948);
xnor U17732 (N_17732,N_7508,N_8110);
nor U17733 (N_17733,N_8632,N_9829);
and U17734 (N_17734,N_8485,N_7655);
or U17735 (N_17735,N_7548,N_11460);
nor U17736 (N_17736,N_10827,N_11571);
or U17737 (N_17737,N_9200,N_11682);
or U17738 (N_17738,N_8879,N_8553);
nand U17739 (N_17739,N_6525,N_11360);
or U17740 (N_17740,N_11929,N_10602);
nand U17741 (N_17741,N_10024,N_11605);
xnor U17742 (N_17742,N_6937,N_10385);
xnor U17743 (N_17743,N_6229,N_10904);
nor U17744 (N_17744,N_6607,N_9119);
and U17745 (N_17745,N_9503,N_6760);
and U17746 (N_17746,N_10976,N_6306);
and U17747 (N_17747,N_10536,N_7949);
nand U17748 (N_17748,N_8538,N_11110);
nand U17749 (N_17749,N_7340,N_6477);
xnor U17750 (N_17750,N_11674,N_8551);
nor U17751 (N_17751,N_11962,N_10129);
nand U17752 (N_17752,N_11808,N_10255);
xnor U17753 (N_17753,N_11038,N_10092);
nor U17754 (N_17754,N_11857,N_6595);
and U17755 (N_17755,N_8320,N_11325);
and U17756 (N_17756,N_11236,N_8980);
and U17757 (N_17757,N_7020,N_11400);
xor U17758 (N_17758,N_7638,N_8807);
and U17759 (N_17759,N_11561,N_6114);
xnor U17760 (N_17760,N_7435,N_7636);
and U17761 (N_17761,N_9715,N_6370);
or U17762 (N_17762,N_8874,N_10566);
nor U17763 (N_17763,N_10600,N_10635);
xnor U17764 (N_17764,N_8215,N_7010);
xnor U17765 (N_17765,N_7710,N_7029);
or U17766 (N_17766,N_9996,N_9519);
nand U17767 (N_17767,N_11189,N_8713);
or U17768 (N_17768,N_10775,N_10957);
nand U17769 (N_17769,N_9190,N_10299);
xor U17770 (N_17770,N_9791,N_9568);
nor U17771 (N_17771,N_10871,N_6369);
nor U17772 (N_17772,N_8684,N_10826);
and U17773 (N_17773,N_6395,N_9750);
or U17774 (N_17774,N_7748,N_6395);
xnor U17775 (N_17775,N_6308,N_9020);
nor U17776 (N_17776,N_8970,N_11395);
nand U17777 (N_17777,N_7110,N_10689);
or U17778 (N_17778,N_9833,N_10904);
nor U17779 (N_17779,N_8671,N_10460);
or U17780 (N_17780,N_7545,N_9155);
nand U17781 (N_17781,N_6745,N_6555);
xor U17782 (N_17782,N_11129,N_10965);
xor U17783 (N_17783,N_7891,N_10431);
or U17784 (N_17784,N_11956,N_9399);
or U17785 (N_17785,N_10530,N_6958);
nand U17786 (N_17786,N_7016,N_7176);
nor U17787 (N_17787,N_9901,N_7022);
and U17788 (N_17788,N_9067,N_8678);
or U17789 (N_17789,N_7703,N_11680);
xor U17790 (N_17790,N_7848,N_6334);
nor U17791 (N_17791,N_8607,N_8227);
xnor U17792 (N_17792,N_10283,N_6752);
and U17793 (N_17793,N_8489,N_8700);
or U17794 (N_17794,N_10361,N_9429);
xor U17795 (N_17795,N_11842,N_10895);
and U17796 (N_17796,N_8006,N_9723);
nand U17797 (N_17797,N_10414,N_8749);
xor U17798 (N_17798,N_7413,N_11276);
or U17799 (N_17799,N_6067,N_6026);
or U17800 (N_17800,N_11117,N_9619);
nand U17801 (N_17801,N_9492,N_10994);
nor U17802 (N_17802,N_11809,N_6071);
xor U17803 (N_17803,N_7016,N_9315);
or U17804 (N_17804,N_9048,N_9681);
nor U17805 (N_17805,N_6350,N_7979);
nand U17806 (N_17806,N_11467,N_7925);
xnor U17807 (N_17807,N_11623,N_7659);
and U17808 (N_17808,N_11214,N_11495);
and U17809 (N_17809,N_9451,N_8329);
xnor U17810 (N_17810,N_11892,N_7254);
nand U17811 (N_17811,N_7205,N_6957);
nand U17812 (N_17812,N_6547,N_9016);
or U17813 (N_17813,N_8201,N_8695);
and U17814 (N_17814,N_6789,N_7589);
nor U17815 (N_17815,N_11373,N_11859);
nand U17816 (N_17816,N_9757,N_9475);
nor U17817 (N_17817,N_7285,N_10051);
nand U17818 (N_17818,N_9142,N_9795);
xor U17819 (N_17819,N_11840,N_9409);
xnor U17820 (N_17820,N_11149,N_9587);
and U17821 (N_17821,N_9007,N_8031);
and U17822 (N_17822,N_11572,N_6974);
and U17823 (N_17823,N_10956,N_6240);
nand U17824 (N_17824,N_7188,N_10643);
or U17825 (N_17825,N_6703,N_7890);
nor U17826 (N_17826,N_9601,N_11291);
nand U17827 (N_17827,N_6440,N_9143);
xnor U17828 (N_17828,N_6727,N_7416);
or U17829 (N_17829,N_11071,N_8013);
nand U17830 (N_17830,N_11148,N_7121);
nand U17831 (N_17831,N_10965,N_7113);
nand U17832 (N_17832,N_6235,N_7957);
xnor U17833 (N_17833,N_8655,N_6485);
xnor U17834 (N_17834,N_7916,N_6141);
and U17835 (N_17835,N_9829,N_7144);
or U17836 (N_17836,N_7878,N_6891);
or U17837 (N_17837,N_10685,N_7965);
xor U17838 (N_17838,N_9536,N_10737);
or U17839 (N_17839,N_10104,N_7988);
nor U17840 (N_17840,N_6285,N_10608);
or U17841 (N_17841,N_6037,N_10355);
nand U17842 (N_17842,N_7803,N_11493);
nand U17843 (N_17843,N_8427,N_8832);
or U17844 (N_17844,N_10926,N_6664);
nand U17845 (N_17845,N_6794,N_8459);
xor U17846 (N_17846,N_9703,N_8594);
and U17847 (N_17847,N_10408,N_11175);
or U17848 (N_17848,N_8528,N_8256);
xnor U17849 (N_17849,N_11820,N_11138);
nor U17850 (N_17850,N_10560,N_11523);
nand U17851 (N_17851,N_6701,N_10635);
xor U17852 (N_17852,N_11448,N_6484);
xnor U17853 (N_17853,N_10915,N_11493);
nor U17854 (N_17854,N_6711,N_6301);
nor U17855 (N_17855,N_7639,N_7758);
xor U17856 (N_17856,N_8078,N_8263);
xor U17857 (N_17857,N_6697,N_6787);
xor U17858 (N_17858,N_8636,N_6314);
and U17859 (N_17859,N_10839,N_10580);
nor U17860 (N_17860,N_7271,N_8600);
or U17861 (N_17861,N_7544,N_11277);
nor U17862 (N_17862,N_7865,N_9280);
and U17863 (N_17863,N_9837,N_7489);
and U17864 (N_17864,N_11539,N_9501);
and U17865 (N_17865,N_6424,N_8720);
or U17866 (N_17866,N_8326,N_6317);
nor U17867 (N_17867,N_7620,N_6460);
xnor U17868 (N_17868,N_7931,N_7028);
nor U17869 (N_17869,N_9480,N_6690);
and U17870 (N_17870,N_11069,N_8122);
xnor U17871 (N_17871,N_11314,N_6334);
nor U17872 (N_17872,N_11195,N_10194);
nor U17873 (N_17873,N_7980,N_8010);
xnor U17874 (N_17874,N_11701,N_11872);
and U17875 (N_17875,N_8519,N_9768);
nor U17876 (N_17876,N_7219,N_8452);
xnor U17877 (N_17877,N_11646,N_7536);
xnor U17878 (N_17878,N_10860,N_10924);
xor U17879 (N_17879,N_8780,N_8755);
nand U17880 (N_17880,N_9663,N_6559);
and U17881 (N_17881,N_7883,N_11468);
and U17882 (N_17882,N_9414,N_8956);
nor U17883 (N_17883,N_9467,N_9558);
xnor U17884 (N_17884,N_6180,N_7024);
xnor U17885 (N_17885,N_11159,N_11878);
or U17886 (N_17886,N_9791,N_7351);
nor U17887 (N_17887,N_10583,N_6161);
or U17888 (N_17888,N_9721,N_11089);
or U17889 (N_17889,N_9684,N_7318);
nor U17890 (N_17890,N_6009,N_7925);
and U17891 (N_17891,N_11056,N_11791);
nand U17892 (N_17892,N_10042,N_6689);
and U17893 (N_17893,N_6708,N_8105);
nand U17894 (N_17894,N_7836,N_7801);
or U17895 (N_17895,N_10189,N_6625);
or U17896 (N_17896,N_8303,N_7945);
nand U17897 (N_17897,N_10040,N_10738);
or U17898 (N_17898,N_10503,N_9827);
xnor U17899 (N_17899,N_9508,N_9470);
and U17900 (N_17900,N_9931,N_6588);
or U17901 (N_17901,N_9051,N_11594);
and U17902 (N_17902,N_9473,N_11664);
nor U17903 (N_17903,N_11679,N_11868);
xnor U17904 (N_17904,N_7561,N_7688);
nand U17905 (N_17905,N_8545,N_10919);
and U17906 (N_17906,N_10139,N_11229);
xnor U17907 (N_17907,N_10798,N_10164);
nor U17908 (N_17908,N_6655,N_8198);
nand U17909 (N_17909,N_7513,N_6385);
or U17910 (N_17910,N_6969,N_10983);
or U17911 (N_17911,N_6089,N_8978);
nand U17912 (N_17912,N_10145,N_10929);
nand U17913 (N_17913,N_8350,N_10082);
and U17914 (N_17914,N_9268,N_11376);
and U17915 (N_17915,N_6404,N_7975);
xor U17916 (N_17916,N_10576,N_11381);
xnor U17917 (N_17917,N_8514,N_8522);
nor U17918 (N_17918,N_7348,N_9212);
nor U17919 (N_17919,N_8579,N_6674);
nor U17920 (N_17920,N_8693,N_8429);
or U17921 (N_17921,N_6933,N_10658);
xnor U17922 (N_17922,N_6517,N_6432);
nand U17923 (N_17923,N_8145,N_8232);
nand U17924 (N_17924,N_9965,N_8683);
or U17925 (N_17925,N_8853,N_7451);
xnor U17926 (N_17926,N_10191,N_10589);
and U17927 (N_17927,N_9969,N_11507);
nand U17928 (N_17928,N_7452,N_8736);
xnor U17929 (N_17929,N_8065,N_7291);
nand U17930 (N_17930,N_6391,N_6054);
and U17931 (N_17931,N_9352,N_9662);
xnor U17932 (N_17932,N_6342,N_11835);
and U17933 (N_17933,N_9268,N_6330);
or U17934 (N_17934,N_8347,N_10812);
nor U17935 (N_17935,N_10793,N_7147);
or U17936 (N_17936,N_8370,N_7504);
and U17937 (N_17937,N_7436,N_6984);
xnor U17938 (N_17938,N_10633,N_8251);
and U17939 (N_17939,N_6706,N_8330);
xor U17940 (N_17940,N_8469,N_11498);
or U17941 (N_17941,N_10066,N_8059);
nor U17942 (N_17942,N_6339,N_6395);
nand U17943 (N_17943,N_9353,N_9137);
or U17944 (N_17944,N_9921,N_9257);
nand U17945 (N_17945,N_10966,N_10348);
nand U17946 (N_17946,N_7892,N_6764);
nand U17947 (N_17947,N_11632,N_11566);
nand U17948 (N_17948,N_9405,N_8689);
nand U17949 (N_17949,N_8099,N_10939);
and U17950 (N_17950,N_10176,N_7526);
xnor U17951 (N_17951,N_11507,N_7025);
and U17952 (N_17952,N_6167,N_9524);
and U17953 (N_17953,N_7623,N_6472);
or U17954 (N_17954,N_7865,N_7217);
or U17955 (N_17955,N_11573,N_8418);
or U17956 (N_17956,N_7976,N_6626);
nor U17957 (N_17957,N_8199,N_9389);
nor U17958 (N_17958,N_9638,N_6090);
xor U17959 (N_17959,N_10682,N_6776);
and U17960 (N_17960,N_8429,N_7303);
nor U17961 (N_17961,N_9555,N_11477);
nand U17962 (N_17962,N_7372,N_9604);
and U17963 (N_17963,N_6186,N_11349);
nor U17964 (N_17964,N_10797,N_11299);
nand U17965 (N_17965,N_7048,N_9833);
and U17966 (N_17966,N_6562,N_11366);
nand U17967 (N_17967,N_8168,N_7010);
and U17968 (N_17968,N_8977,N_11869);
and U17969 (N_17969,N_9402,N_6414);
nor U17970 (N_17970,N_9273,N_9293);
nand U17971 (N_17971,N_11552,N_10057);
nor U17972 (N_17972,N_6254,N_8157);
or U17973 (N_17973,N_7123,N_7776);
nor U17974 (N_17974,N_9459,N_10202);
and U17975 (N_17975,N_8040,N_10015);
or U17976 (N_17976,N_9903,N_7313);
xnor U17977 (N_17977,N_10449,N_8777);
or U17978 (N_17978,N_11755,N_10808);
nand U17979 (N_17979,N_11725,N_11863);
or U17980 (N_17980,N_9532,N_7086);
and U17981 (N_17981,N_9980,N_10661);
nand U17982 (N_17982,N_11521,N_11289);
or U17983 (N_17983,N_7820,N_11563);
nand U17984 (N_17984,N_9655,N_7321);
nor U17985 (N_17985,N_10480,N_7445);
and U17986 (N_17986,N_9896,N_7894);
nor U17987 (N_17987,N_7248,N_9035);
or U17988 (N_17988,N_11341,N_9668);
nand U17989 (N_17989,N_6329,N_11074);
or U17990 (N_17990,N_9907,N_7072);
nor U17991 (N_17991,N_6508,N_11670);
nand U17992 (N_17992,N_9145,N_9500);
nand U17993 (N_17993,N_6158,N_6698);
nor U17994 (N_17994,N_6498,N_9183);
and U17995 (N_17995,N_7936,N_7256);
or U17996 (N_17996,N_8626,N_7761);
and U17997 (N_17997,N_9655,N_8257);
xnor U17998 (N_17998,N_11108,N_6872);
and U17999 (N_17999,N_7899,N_9527);
xnor U18000 (N_18000,N_15947,N_16714);
nand U18001 (N_18001,N_14913,N_17775);
xnor U18002 (N_18002,N_15522,N_17553);
nand U18003 (N_18003,N_12373,N_13622);
xor U18004 (N_18004,N_12673,N_16035);
nand U18005 (N_18005,N_14798,N_14336);
nand U18006 (N_18006,N_16437,N_14437);
nand U18007 (N_18007,N_17792,N_16897);
nor U18008 (N_18008,N_14388,N_15722);
or U18009 (N_18009,N_15463,N_15971);
or U18010 (N_18010,N_17758,N_16625);
and U18011 (N_18011,N_17748,N_16224);
nand U18012 (N_18012,N_13018,N_15901);
nand U18013 (N_18013,N_17299,N_16737);
and U18014 (N_18014,N_13507,N_12076);
or U18015 (N_18015,N_14276,N_12528);
nor U18016 (N_18016,N_15919,N_13669);
or U18017 (N_18017,N_15850,N_17128);
nor U18018 (N_18018,N_17439,N_12607);
xnor U18019 (N_18019,N_16918,N_16116);
xor U18020 (N_18020,N_15593,N_15026);
or U18021 (N_18021,N_14701,N_12288);
xor U18022 (N_18022,N_15363,N_13445);
and U18023 (N_18023,N_14571,N_14522);
nand U18024 (N_18024,N_12220,N_16923);
nor U18025 (N_18025,N_16922,N_14268);
or U18026 (N_18026,N_15196,N_12201);
nor U18027 (N_18027,N_17222,N_17002);
nor U18028 (N_18028,N_16377,N_12928);
nor U18029 (N_18029,N_12548,N_14319);
nand U18030 (N_18030,N_13460,N_16599);
nand U18031 (N_18031,N_12275,N_13878);
nand U18032 (N_18032,N_13231,N_17443);
or U18033 (N_18033,N_12139,N_15879);
nor U18034 (N_18034,N_15200,N_16171);
or U18035 (N_18035,N_12137,N_16121);
nand U18036 (N_18036,N_15863,N_12209);
nand U18037 (N_18037,N_17802,N_14552);
and U18038 (N_18038,N_15348,N_17018);
nand U18039 (N_18039,N_14289,N_13391);
xnor U18040 (N_18040,N_15712,N_15686);
nand U18041 (N_18041,N_13162,N_13952);
and U18042 (N_18042,N_14012,N_14057);
or U18043 (N_18043,N_13191,N_17692);
and U18044 (N_18044,N_13384,N_14929);
xor U18045 (N_18045,N_17753,N_13850);
xnor U18046 (N_18046,N_13113,N_16088);
or U18047 (N_18047,N_17209,N_16279);
nor U18048 (N_18048,N_17764,N_14860);
nor U18049 (N_18049,N_15965,N_17142);
or U18050 (N_18050,N_16663,N_17939);
nand U18051 (N_18051,N_17776,N_13814);
xnor U18052 (N_18052,N_15680,N_12223);
or U18053 (N_18053,N_13419,N_12508);
nand U18054 (N_18054,N_15380,N_13332);
or U18055 (N_18055,N_16677,N_17712);
or U18056 (N_18056,N_14524,N_13809);
xor U18057 (N_18057,N_14055,N_17216);
xor U18058 (N_18058,N_13681,N_12540);
and U18059 (N_18059,N_15643,N_12334);
or U18060 (N_18060,N_16765,N_13706);
xnor U18061 (N_18061,N_14361,N_17480);
nand U18062 (N_18062,N_14517,N_16881);
nor U18063 (N_18063,N_17635,N_13940);
nor U18064 (N_18064,N_15549,N_13103);
and U18065 (N_18065,N_14627,N_12907);
xor U18066 (N_18066,N_13239,N_17253);
xnor U18067 (N_18067,N_12065,N_15498);
nand U18068 (N_18068,N_14611,N_15271);
nand U18069 (N_18069,N_16685,N_14778);
or U18070 (N_18070,N_15295,N_12460);
nand U18071 (N_18071,N_13229,N_14290);
nor U18072 (N_18072,N_16410,N_14312);
nor U18073 (N_18073,N_12513,N_15562);
nor U18074 (N_18074,N_14294,N_15246);
and U18075 (N_18075,N_15467,N_16866);
nor U18076 (N_18076,N_16096,N_17741);
or U18077 (N_18077,N_14354,N_12775);
nor U18078 (N_18078,N_15563,N_12984);
and U18079 (N_18079,N_15984,N_16278);
nand U18080 (N_18080,N_13274,N_16013);
nand U18081 (N_18081,N_12785,N_14813);
nand U18082 (N_18082,N_13275,N_12180);
nor U18083 (N_18083,N_17115,N_13314);
and U18084 (N_18084,N_17583,N_16488);
and U18085 (N_18085,N_14563,N_13825);
nand U18086 (N_18086,N_16733,N_16791);
or U18087 (N_18087,N_17965,N_12215);
nor U18088 (N_18088,N_17352,N_17261);
or U18089 (N_18089,N_12880,N_16125);
and U18090 (N_18090,N_16011,N_13715);
and U18091 (N_18091,N_13582,N_17586);
nand U18092 (N_18092,N_17033,N_13840);
nor U18093 (N_18093,N_14063,N_12127);
or U18094 (N_18094,N_16548,N_15437);
and U18095 (N_18095,N_12178,N_17199);
nor U18096 (N_18096,N_13614,N_14352);
nor U18097 (N_18097,N_15660,N_12897);
and U18098 (N_18098,N_16296,N_17448);
or U18099 (N_18099,N_14954,N_15761);
xnor U18100 (N_18100,N_13546,N_14265);
xor U18101 (N_18101,N_16168,N_13693);
nor U18102 (N_18102,N_16858,N_17742);
nor U18103 (N_18103,N_15827,N_16212);
nor U18104 (N_18104,N_12336,N_12779);
and U18105 (N_18105,N_14349,N_17403);
and U18106 (N_18106,N_14904,N_12463);
and U18107 (N_18107,N_17623,N_12794);
and U18108 (N_18108,N_12703,N_12555);
nand U18109 (N_18109,N_13765,N_12530);
nand U18110 (N_18110,N_15410,N_13659);
xor U18111 (N_18111,N_15320,N_16645);
nand U18112 (N_18112,N_17987,N_16855);
or U18113 (N_18113,N_15935,N_12154);
nand U18114 (N_18114,N_14187,N_12877);
nor U18115 (N_18115,N_16758,N_14178);
nor U18116 (N_18116,N_15442,N_13476);
xor U18117 (N_18117,N_12527,N_13657);
and U18118 (N_18118,N_15951,N_13615);
nor U18119 (N_18119,N_12677,N_13766);
and U18120 (N_18120,N_17752,N_15378);
xor U18121 (N_18121,N_12533,N_12744);
nor U18122 (N_18122,N_13217,N_13966);
nor U18123 (N_18123,N_15881,N_15094);
nor U18124 (N_18124,N_15351,N_14831);
xnor U18125 (N_18125,N_15021,N_12312);
nand U18126 (N_18126,N_13104,N_17750);
and U18127 (N_18127,N_12253,N_16823);
xnor U18128 (N_18128,N_14123,N_15603);
xor U18129 (N_18129,N_13673,N_14987);
and U18130 (N_18130,N_17052,N_12683);
nor U18131 (N_18131,N_13632,N_15400);
and U18132 (N_18132,N_16953,N_12939);
nand U18133 (N_18133,N_16556,N_17551);
and U18134 (N_18134,N_14084,N_17360);
nand U18135 (N_18135,N_13491,N_17933);
nor U18136 (N_18136,N_15068,N_15849);
nor U18137 (N_18137,N_14826,N_17871);
nand U18138 (N_18138,N_13490,N_17864);
xor U18139 (N_18139,N_14003,N_12791);
nor U18140 (N_18140,N_17993,N_12261);
or U18141 (N_18141,N_15610,N_16103);
or U18142 (N_18142,N_13980,N_16945);
or U18143 (N_18143,N_16266,N_13779);
nor U18144 (N_18144,N_14089,N_17349);
xnor U18145 (N_18145,N_14341,N_17361);
nor U18146 (N_18146,N_17807,N_13876);
nor U18147 (N_18147,N_13260,N_14328);
nor U18148 (N_18148,N_13728,N_12222);
xnor U18149 (N_18149,N_12048,N_13487);
and U18150 (N_18150,N_12204,N_16308);
or U18151 (N_18151,N_15720,N_17540);
nand U18152 (N_18152,N_12698,N_12413);
nand U18153 (N_18153,N_13945,N_13888);
xnor U18154 (N_18154,N_14953,N_12562);
nand U18155 (N_18155,N_16948,N_14539);
nand U18156 (N_18156,N_17044,N_16433);
xor U18157 (N_18157,N_12476,N_15174);
and U18158 (N_18158,N_17098,N_12458);
nand U18159 (N_18159,N_13080,N_13283);
or U18160 (N_18160,N_12612,N_14148);
nor U18161 (N_18161,N_17683,N_17240);
and U18162 (N_18162,N_13355,N_13551);
nor U18163 (N_18163,N_17985,N_16751);
nand U18164 (N_18164,N_13819,N_13864);
nor U18165 (N_18165,N_14261,N_12608);
nand U18166 (N_18166,N_15359,N_16317);
and U18167 (N_18167,N_13707,N_16339);
nand U18168 (N_18168,N_13999,N_14194);
nand U18169 (N_18169,N_17339,N_12024);
or U18170 (N_18170,N_12447,N_16098);
or U18171 (N_18171,N_14947,N_14587);
and U18172 (N_18172,N_16331,N_16336);
nand U18173 (N_18173,N_15873,N_15303);
xnor U18174 (N_18174,N_16844,N_14252);
xnor U18175 (N_18175,N_14879,N_15353);
and U18176 (N_18176,N_16459,N_17020);
nor U18177 (N_18177,N_14795,N_12181);
nor U18178 (N_18178,N_16190,N_14966);
or U18179 (N_18179,N_15817,N_15786);
and U18180 (N_18180,N_15818,N_16184);
or U18181 (N_18181,N_17949,N_13421);
or U18182 (N_18182,N_13379,N_12625);
and U18183 (N_18183,N_13039,N_16977);
nand U18184 (N_18184,N_15001,N_14781);
nand U18185 (N_18185,N_12022,N_16407);
and U18186 (N_18186,N_12848,N_14203);
nor U18187 (N_18187,N_16661,N_16817);
and U18188 (N_18188,N_14130,N_13292);
or U18189 (N_18189,N_14287,N_15236);
xor U18190 (N_18190,N_15531,N_15515);
or U18191 (N_18191,N_17212,N_14416);
xor U18192 (N_18192,N_17878,N_13059);
nor U18193 (N_18193,N_16469,N_12218);
and U18194 (N_18194,N_13932,N_17724);
xor U18195 (N_18195,N_15733,N_14930);
nand U18196 (N_18196,N_14565,N_17693);
xor U18197 (N_18197,N_15650,N_16099);
nand U18198 (N_18198,N_12506,N_12242);
and U18199 (N_18199,N_13442,N_17231);
nand U18200 (N_18200,N_12667,N_16983);
and U18201 (N_18201,N_17035,N_17326);
nand U18202 (N_18202,N_15355,N_16623);
nor U18203 (N_18203,N_16853,N_16762);
xnor U18204 (N_18204,N_14286,N_16890);
and U18205 (N_18205,N_12961,N_17524);
nor U18206 (N_18206,N_13015,N_17182);
or U18207 (N_18207,N_14711,N_13957);
nand U18208 (N_18208,N_14050,N_15691);
nor U18209 (N_18209,N_16448,N_15737);
xor U18210 (N_18210,N_14880,N_13913);
xnor U18211 (N_18211,N_14511,N_12751);
or U18212 (N_18212,N_17913,N_13408);
or U18213 (N_18213,N_16540,N_14193);
nand U18214 (N_18214,N_12094,N_16759);
xor U18215 (N_18215,N_17766,N_14535);
xnor U18216 (N_18216,N_16474,N_12063);
and U18217 (N_18217,N_13061,N_15006);
or U18218 (N_18218,N_17073,N_17196);
nor U18219 (N_18219,N_14878,N_16535);
xnor U18220 (N_18220,N_13738,N_12002);
xnor U18221 (N_18221,N_15699,N_12882);
or U18222 (N_18222,N_16005,N_12115);
nand U18223 (N_18223,N_13081,N_12274);
or U18224 (N_18224,N_17607,N_12498);
nand U18225 (N_18225,N_12773,N_13433);
xnor U18226 (N_18226,N_15809,N_16213);
and U18227 (N_18227,N_12500,N_13197);
nor U18228 (N_18228,N_13782,N_14374);
nand U18229 (N_18229,N_12681,N_16624);
xnor U18230 (N_18230,N_17050,N_12472);
or U18231 (N_18231,N_14083,N_12487);
nor U18232 (N_18232,N_15461,N_16829);
and U18233 (N_18233,N_15941,N_12596);
xor U18234 (N_18234,N_12095,N_14121);
and U18235 (N_18235,N_16343,N_15128);
nor U18236 (N_18236,N_12372,N_12466);
or U18237 (N_18237,N_17247,N_12292);
or U18238 (N_18238,N_12719,N_17272);
xor U18239 (N_18239,N_14212,N_17120);
nand U18240 (N_18240,N_17608,N_17264);
nand U18241 (N_18241,N_13121,N_14686);
and U18242 (N_18242,N_12584,N_17566);
and U18243 (N_18243,N_13639,N_15061);
nor U18244 (N_18244,N_16041,N_16076);
and U18245 (N_18245,N_13203,N_14292);
xnor U18246 (N_18246,N_14997,N_15771);
nand U18247 (N_18247,N_13316,N_17704);
nor U18248 (N_18248,N_13106,N_13858);
and U18249 (N_18249,N_16723,N_16659);
or U18250 (N_18250,N_15018,N_13063);
and U18251 (N_18251,N_13526,N_14972);
nand U18252 (N_18252,N_14496,N_15264);
nand U18253 (N_18253,N_12806,N_16430);
nor U18254 (N_18254,N_16263,N_15474);
nand U18255 (N_18255,N_16238,N_17463);
nor U18256 (N_18256,N_12817,N_14177);
and U18257 (N_18257,N_16697,N_17945);
nand U18258 (N_18258,N_17706,N_15429);
xor U18259 (N_18259,N_15548,N_15744);
or U18260 (N_18260,N_12769,N_14072);
and U18261 (N_18261,N_12400,N_16452);
and U18262 (N_18262,N_13611,N_16175);
xor U18263 (N_18263,N_12924,N_12718);
nand U18264 (N_18264,N_16141,N_17307);
and U18265 (N_18265,N_16773,N_12066);
nand U18266 (N_18266,N_15729,N_12490);
nor U18267 (N_18267,N_16027,N_17007);
nand U18268 (N_18268,N_16143,N_14030);
or U18269 (N_18269,N_17080,N_15109);
and U18270 (N_18270,N_12863,N_13584);
and U18271 (N_18271,N_15826,N_17702);
and U18272 (N_18272,N_17657,N_14493);
nor U18273 (N_18273,N_12245,N_16669);
and U18274 (N_18274,N_15917,N_17058);
xor U18275 (N_18275,N_15226,N_14410);
or U18276 (N_18276,N_16439,N_15981);
or U18277 (N_18277,N_17428,N_17885);
or U18278 (N_18278,N_14054,N_13296);
or U18279 (N_18279,N_15685,N_12384);
nor U18280 (N_18280,N_15677,N_14936);
nor U18281 (N_18281,N_13906,N_14305);
and U18282 (N_18282,N_16649,N_16609);
nor U18283 (N_18283,N_15465,N_15605);
nor U18284 (N_18284,N_12529,N_14747);
and U18285 (N_18285,N_17631,N_14236);
or U18286 (N_18286,N_16257,N_16491);
nor U18287 (N_18287,N_13247,N_15112);
or U18288 (N_18288,N_13192,N_17300);
nand U18289 (N_18289,N_16929,N_14401);
xnor U18290 (N_18290,N_12231,N_15915);
and U18291 (N_18291,N_16460,N_15052);
and U18292 (N_18292,N_14132,N_13482);
xnor U18293 (N_18293,N_17109,N_13310);
nor U18294 (N_18294,N_14803,N_13363);
or U18295 (N_18295,N_13323,N_17350);
xnor U18296 (N_18296,N_15375,N_17685);
or U18297 (N_18297,N_17681,N_13534);
xnor U18298 (N_18298,N_15622,N_12659);
or U18299 (N_18299,N_14209,N_13590);
xor U18300 (N_18300,N_12816,N_14351);
or U18301 (N_18301,N_17102,N_15512);
nor U18302 (N_18302,N_12097,N_14149);
and U18303 (N_18303,N_16424,N_16490);
nor U18304 (N_18304,N_13093,N_14028);
nor U18305 (N_18305,N_13443,N_12309);
or U18306 (N_18306,N_15801,N_16050);
nor U18307 (N_18307,N_13591,N_14777);
xnor U18308 (N_18308,N_12333,N_12355);
nor U18309 (N_18309,N_16062,N_14845);
or U18310 (N_18310,N_17411,N_15399);
and U18311 (N_18311,N_16290,N_14489);
and U18312 (N_18312,N_14939,N_12235);
nor U18313 (N_18313,N_17267,N_15511);
nor U18314 (N_18314,N_13056,N_12303);
nor U18315 (N_18315,N_14949,N_13117);
or U18316 (N_18316,N_15417,N_14830);
nor U18317 (N_18317,N_16235,N_12229);
nand U18318 (N_18318,N_16384,N_12868);
and U18319 (N_18319,N_14670,N_15851);
and U18320 (N_18320,N_13802,N_15087);
or U18321 (N_18321,N_14582,N_16668);
or U18322 (N_18322,N_17368,N_13633);
nor U18323 (N_18323,N_13578,N_16306);
xnor U18324 (N_18324,N_14449,N_16501);
and U18325 (N_18325,N_14179,N_12564);
and U18326 (N_18326,N_13086,N_17356);
xnor U18327 (N_18327,N_15185,N_16323);
or U18328 (N_18328,N_17250,N_17729);
and U18329 (N_18329,N_13020,N_15521);
or U18330 (N_18330,N_12774,N_16223);
and U18331 (N_18331,N_15913,N_16557);
nor U18332 (N_18332,N_16509,N_17423);
or U18333 (N_18333,N_13222,N_13986);
and U18334 (N_18334,N_17152,N_15518);
nor U18335 (N_18335,N_14785,N_16916);
and U18336 (N_18336,N_16788,N_12890);
or U18337 (N_18337,N_15985,N_15110);
nor U18338 (N_18338,N_15779,N_16389);
nor U18339 (N_18339,N_16613,N_15898);
nand U18340 (N_18340,N_14636,N_15445);
nand U18341 (N_18341,N_16149,N_16978);
and U18342 (N_18342,N_17866,N_16741);
xor U18343 (N_18343,N_12313,N_14256);
and U18344 (N_18344,N_16691,N_12249);
nor U18345 (N_18345,N_13612,N_17535);
or U18346 (N_18346,N_15231,N_17208);
xnor U18347 (N_18347,N_15938,N_12386);
or U18348 (N_18348,N_14591,N_13270);
nand U18349 (N_18349,N_13955,N_12704);
nand U18350 (N_18350,N_14060,N_14792);
or U18351 (N_18351,N_17552,N_13418);
or U18352 (N_18352,N_16170,N_12379);
nand U18353 (N_18353,N_13392,N_14473);
or U18354 (N_18354,N_16217,N_13756);
nor U18355 (N_18355,N_13874,N_13087);
and U18356 (N_18356,N_13827,N_13930);
xnor U18357 (N_18357,N_13359,N_16255);
and U18358 (N_18358,N_16322,N_14327);
nand U18359 (N_18359,N_13923,N_16552);
xnor U18360 (N_18360,N_15103,N_13522);
or U18361 (N_18361,N_16568,N_17343);
xor U18362 (N_18362,N_12834,N_13778);
xor U18363 (N_18363,N_15386,N_14288);
xnor U18364 (N_18364,N_13905,N_12573);
and U18365 (N_18365,N_17316,N_16467);
and U18366 (N_18366,N_13299,N_17176);
nor U18367 (N_18367,N_17771,N_16462);
xnor U18368 (N_18368,N_13640,N_12501);
and U18369 (N_18369,N_17141,N_14850);
xnor U18370 (N_18370,N_15148,N_17429);
and U18371 (N_18371,N_12759,N_15332);
nand U18372 (N_18372,N_14669,N_17075);
xnor U18373 (N_18373,N_15130,N_12503);
nor U18374 (N_18374,N_17589,N_13025);
or U18375 (N_18375,N_15239,N_16689);
xor U18376 (N_18376,N_16973,N_14748);
nand U18377 (N_18377,N_13894,N_15811);
nand U18378 (N_18378,N_15299,N_15910);
xnor U18379 (N_18379,N_12109,N_12944);
and U18380 (N_18380,N_14460,N_12662);
xor U18381 (N_18381,N_13513,N_17698);
or U18382 (N_18382,N_16642,N_13023);
and U18383 (N_18383,N_17996,N_14921);
nor U18384 (N_18384,N_12597,N_15944);
and U18385 (N_18385,N_17558,N_16966);
and U18386 (N_18386,N_16284,N_13860);
nand U18387 (N_18387,N_17404,N_12053);
nor U18388 (N_18388,N_17042,N_14697);
nand U18389 (N_18389,N_17907,N_17230);
or U18390 (N_18390,N_17498,N_13708);
or U18391 (N_18391,N_16361,N_17943);
nor U18392 (N_18392,N_13245,N_17687);
and U18393 (N_18393,N_15591,N_15015);
or U18394 (N_18394,N_15413,N_12566);
or U18395 (N_18395,N_13798,N_13474);
xnor U18396 (N_18396,N_15431,N_15928);
nand U18397 (N_18397,N_16493,N_15409);
nor U18398 (N_18398,N_15020,N_14903);
nand U18399 (N_18399,N_15080,N_15621);
and U18400 (N_18400,N_13548,N_12323);
nor U18401 (N_18401,N_12427,N_15450);
or U18402 (N_18402,N_15436,N_17600);
and U18403 (N_18403,N_12046,N_14544);
nor U18404 (N_18404,N_13336,N_12823);
nor U18405 (N_18405,N_12391,N_15244);
xor U18406 (N_18406,N_16340,N_16589);
or U18407 (N_18407,N_17386,N_13190);
nand U18408 (N_18408,N_16730,N_14757);
or U18409 (N_18409,N_13069,N_13184);
nor U18410 (N_18410,N_16161,N_14569);
xor U18411 (N_18411,N_12800,N_17351);
nor U18412 (N_18412,N_17082,N_14906);
or U18413 (N_18413,N_17405,N_12227);
nor U18414 (N_18414,N_16662,N_14694);
and U18415 (N_18415,N_12987,N_16517);
nand U18416 (N_18416,N_15261,N_14521);
and U18417 (N_18417,N_12434,N_12068);
nand U18418 (N_18418,N_14868,N_15608);
nand U18419 (N_18419,N_17280,N_16478);
nor U18420 (N_18420,N_17767,N_17735);
nand U18421 (N_18421,N_15478,N_13154);
nor U18422 (N_18422,N_12314,N_12788);
xnor U18423 (N_18423,N_12795,N_16242);
xor U18424 (N_18424,N_12202,N_16716);
nor U18425 (N_18425,N_16100,N_14750);
xnor U18426 (N_18426,N_12230,N_15497);
nand U18427 (N_18427,N_15854,N_15575);
or U18428 (N_18428,N_17140,N_15337);
nand U18429 (N_18429,N_16109,N_16803);
and U18430 (N_18430,N_17015,N_16288);
nor U18431 (N_18431,N_12731,N_16138);
nand U18432 (N_18432,N_16409,N_13434);
or U18433 (N_18433,N_12102,N_12299);
or U18434 (N_18434,N_17482,N_14106);
and U18435 (N_18435,N_13322,N_13959);
or U18436 (N_18436,N_16394,N_16270);
or U18437 (N_18437,N_13238,N_15255);
nor U18438 (N_18438,N_14926,N_15657);
or U18439 (N_18439,N_13908,N_12971);
or U18440 (N_18440,N_12916,N_13468);
xnor U18441 (N_18441,N_13109,N_16083);
or U18442 (N_18442,N_17110,N_16933);
nor U18443 (N_18443,N_14267,N_15457);
nor U18444 (N_18444,N_17399,N_17220);
or U18445 (N_18445,N_16180,N_16291);
xnor U18446 (N_18446,N_15049,N_14973);
and U18447 (N_18447,N_12544,N_16570);
nor U18448 (N_18448,N_15262,N_16167);
and U18449 (N_18449,N_15560,N_13409);
or U18450 (N_18450,N_14441,N_13563);
nor U18451 (N_18451,N_14963,N_15750);
xnor U18452 (N_18452,N_15510,N_15287);
xnor U18453 (N_18453,N_13100,N_15194);
and U18454 (N_18454,N_16513,N_12128);
nor U18455 (N_18455,N_12219,N_12898);
xor U18456 (N_18456,N_16499,N_14301);
or U18457 (N_18457,N_14841,N_17249);
nand U18458 (N_18458,N_12468,N_13593);
or U18459 (N_18459,N_15085,N_17714);
nor U18460 (N_18460,N_17389,N_16174);
xnor U18461 (N_18461,N_12349,N_15684);
nand U18462 (N_18462,N_14505,N_13941);
nor U18463 (N_18463,N_17779,N_12614);
or U18464 (N_18464,N_17625,N_16672);
xor U18465 (N_18465,N_14481,N_16806);
nor U18466 (N_18466,N_13007,N_16782);
nor U18467 (N_18467,N_16392,N_16172);
xor U18468 (N_18468,N_14783,N_16422);
and U18469 (N_18469,N_13510,N_12895);
or U18470 (N_18470,N_12524,N_15808);
and U18471 (N_18471,N_14993,N_15064);
and U18472 (N_18472,N_13603,N_16840);
nor U18473 (N_18473,N_12159,N_12353);
xnor U18474 (N_18474,N_17045,N_17195);
nor U18475 (N_18475,N_16396,N_17946);
nand U18476 (N_18476,N_15289,N_15707);
or U18477 (N_18477,N_12870,N_13459);
or U18478 (N_18478,N_13805,N_12482);
nor U18479 (N_18479,N_12492,N_15379);
nor U18480 (N_18480,N_16991,N_17257);
nand U18481 (N_18481,N_13464,N_15115);
xnor U18482 (N_18482,N_17202,N_15252);
nand U18483 (N_18483,N_15290,N_13366);
nor U18484 (N_18484,N_17129,N_16781);
nor U18485 (N_18485,N_16952,N_14630);
xor U18486 (N_18486,N_14938,N_16163);
or U18487 (N_18487,N_12894,N_12151);
and U18488 (N_18488,N_17972,N_17438);
xnor U18489 (N_18489,N_17135,N_16411);
nor U18490 (N_18490,N_14674,N_15710);
xor U18491 (N_18491,N_17223,N_17150);
nand U18492 (N_18492,N_15743,N_13796);
nand U18493 (N_18493,N_16004,N_17301);
and U18494 (N_18494,N_16947,N_12058);
or U18495 (N_18495,N_17296,N_12602);
xnor U18496 (N_18496,N_17994,N_12734);
or U18497 (N_18497,N_15775,N_16502);
nand U18498 (N_18498,N_16877,N_17757);
xor U18499 (N_18499,N_16944,N_14719);
or U18500 (N_18500,N_12887,N_17157);
or U18501 (N_18501,N_14210,N_17582);
and U18502 (N_18502,N_16770,N_16763);
nor U18503 (N_18503,N_12193,N_14604);
nor U18504 (N_18504,N_15909,N_14242);
or U18505 (N_18505,N_17557,N_16956);
nor U18506 (N_18506,N_12325,N_13842);
and U18507 (N_18507,N_17393,N_12093);
nand U18508 (N_18508,N_17923,N_16931);
nor U18509 (N_18509,N_17827,N_16379);
nand U18510 (N_18510,N_16114,N_17062);
xor U18511 (N_18511,N_17621,N_17294);
nor U18512 (N_18512,N_16198,N_16547);
or U18513 (N_18513,N_13564,N_13988);
and U18514 (N_18514,N_16720,N_16383);
xnor U18515 (N_18515,N_12889,N_15234);
nand U18516 (N_18516,N_13733,N_16153);
xor U18517 (N_18517,N_16381,N_13174);
xor U18518 (N_18518,N_12329,N_12514);
or U18519 (N_18519,N_17710,N_12161);
nor U18520 (N_18520,N_16312,N_14542);
nor U18521 (N_18521,N_17911,N_13315);
and U18522 (N_18522,N_15772,N_13241);
or U18523 (N_18523,N_13989,N_13248);
nor U18524 (N_18524,N_14971,N_15084);
and U18525 (N_18525,N_13009,N_12854);
nand U18526 (N_18526,N_12622,N_12687);
or U18527 (N_18527,N_17134,N_17915);
xor U18528 (N_18528,N_13370,N_13764);
nand U18529 (N_18529,N_14262,N_15412);
xnor U18530 (N_18530,N_17021,N_15609);
xor U18531 (N_18531,N_16295,N_12164);
nand U18532 (N_18532,N_17534,N_12583);
xor U18533 (N_18533,N_17794,N_15166);
nor U18534 (N_18534,N_17440,N_13968);
and U18535 (N_18535,N_16302,N_12551);
xnor U18536 (N_18536,N_13138,N_14408);
nor U18537 (N_18537,N_16102,N_16398);
nor U18538 (N_18538,N_17156,N_15611);
or U18539 (N_18539,N_15335,N_14730);
nand U18540 (N_18540,N_16528,N_14486);
nand U18541 (N_18541,N_17454,N_14566);
nor U18542 (N_18542,N_13592,N_17270);
and U18543 (N_18543,N_15994,N_16193);
nand U18544 (N_18544,N_16033,N_14466);
nor U18545 (N_18545,N_14735,N_16992);
nand U18546 (N_18546,N_13900,N_15118);
xnor U18547 (N_18547,N_16755,N_17036);
or U18548 (N_18548,N_14293,N_16955);
nor U18549 (N_18549,N_16608,N_17457);
or U18550 (N_18550,N_16387,N_12361);
or U18551 (N_18551,N_15306,N_14000);
and U18552 (N_18552,N_16285,N_17358);
nand U18553 (N_18553,N_13996,N_13698);
xnor U18554 (N_18554,N_12525,N_17975);
and U18555 (N_18555,N_17990,N_14923);
xor U18556 (N_18556,N_16214,N_16523);
nor U18557 (N_18557,N_12112,N_17584);
and U18558 (N_18558,N_17611,N_14677);
or U18559 (N_18559,N_17610,N_16903);
or U18560 (N_18560,N_12824,N_12835);
nand U18561 (N_18561,N_12799,N_17675);
xor U18562 (N_18562,N_15574,N_15922);
nor U18563 (N_18563,N_12156,N_16969);
nand U18564 (N_18564,N_14738,N_14198);
and U18565 (N_18565,N_14482,N_17497);
nand U18566 (N_18566,N_16971,N_15098);
nand U18567 (N_18567,N_16412,N_12884);
or U18568 (N_18568,N_17896,N_12695);
nor U18569 (N_18569,N_15868,N_16177);
nor U18570 (N_18570,N_16246,N_16464);
xor U18571 (N_18571,N_12936,N_17780);
xnor U18572 (N_18572,N_16577,N_12541);
nand U18573 (N_18573,N_14403,N_12712);
nand U18574 (N_18574,N_14185,N_14806);
and U18575 (N_18575,N_16333,N_15945);
nand U18576 (N_18576,N_17854,N_15652);
nor U18577 (N_18577,N_13172,N_17633);
nor U18578 (N_18578,N_12184,N_15003);
nor U18579 (N_18579,N_13630,N_12031);
or U18580 (N_18580,N_12485,N_14760);
xor U18581 (N_18581,N_15486,N_14284);
xor U18582 (N_18582,N_14197,N_15315);
and U18583 (N_18583,N_14532,N_12014);
nor U18584 (N_18584,N_12951,N_14439);
xor U18585 (N_18585,N_15173,N_16309);
or U18586 (N_18586,N_17163,N_17648);
or U18587 (N_18587,N_17521,N_12431);
xor U18588 (N_18588,N_12320,N_17263);
xor U18589 (N_18589,N_17942,N_15216);
xnor U18590 (N_18590,N_16602,N_16869);
and U18591 (N_18591,N_17555,N_12973);
xor U18592 (N_18592,N_16395,N_13397);
nor U18593 (N_18593,N_12956,N_17254);
xnor U18594 (N_18594,N_15207,N_14714);
and U18595 (N_18595,N_14272,N_14126);
nand U18596 (N_18596,N_12910,N_14251);
nor U18597 (N_18597,N_14779,N_12813);
nand U18598 (N_18598,N_17432,N_15878);
xnor U18599 (N_18599,N_14821,N_14547);
nor U18600 (N_18600,N_15120,N_13290);
xnor U18601 (N_18601,N_14551,N_12586);
nor U18602 (N_18602,N_13532,N_14513);
and U18603 (N_18603,N_17153,N_15745);
nand U18604 (N_18604,N_16385,N_16251);
nand U18605 (N_18605,N_13494,N_15493);
or U18606 (N_18606,N_14311,N_13886);
nand U18607 (N_18607,N_15663,N_14548);
and U18608 (N_18608,N_14530,N_15282);
and U18609 (N_18609,N_12212,N_14069);
and U18610 (N_18610,N_17215,N_17256);
nor U18611 (N_18611,N_12020,N_16843);
nor U18612 (N_18612,N_17906,N_12642);
or U18613 (N_18613,N_15833,N_14353);
xnor U18614 (N_18614,N_17636,N_17620);
nand U18615 (N_18615,N_17470,N_12904);
nand U18616 (N_18616,N_14946,N_14010);
nand U18617 (N_18617,N_17210,N_13875);
and U18618 (N_18618,N_16209,N_16048);
and U18619 (N_18619,N_12730,N_17720);
or U18620 (N_18620,N_17359,N_12302);
xnor U18621 (N_18621,N_16614,N_12803);
nand U18622 (N_18622,N_14269,N_13567);
nand U18623 (N_18623,N_17916,N_12761);
nand U18624 (N_18624,N_15304,N_13685);
xor U18625 (N_18625,N_16105,N_12366);
nand U18626 (N_18626,N_17982,N_14641);
or U18627 (N_18627,N_17362,N_14141);
nor U18628 (N_18628,N_14870,N_13743);
nand U18629 (N_18629,N_16710,N_12663);
and U18630 (N_18630,N_17969,N_16095);
xor U18631 (N_18631,N_13912,N_13401);
nand U18632 (N_18632,N_15394,N_12407);
and U18633 (N_18633,N_13128,N_14044);
nand U18634 (N_18634,N_15158,N_13909);
xnor U18635 (N_18635,N_15912,N_15292);
or U18636 (N_18636,N_17198,N_14295);
nand U18637 (N_18637,N_16899,N_17839);
or U18638 (N_18638,N_13097,N_17616);
nand U18639 (N_18639,N_13992,N_16274);
nor U18640 (N_18640,N_15250,N_15724);
xor U18641 (N_18641,N_16181,N_14567);
and U18642 (N_18642,N_14699,N_13646);
and U18643 (N_18643,N_16130,N_16546);
xor U18644 (N_18644,N_17663,N_15129);
and U18645 (N_18645,N_16696,N_14739);
or U18646 (N_18646,N_15342,N_17894);
xnor U18647 (N_18647,N_14306,N_16236);
nor U18648 (N_18648,N_14412,N_16965);
nand U18649 (N_18649,N_14969,N_13373);
xor U18650 (N_18650,N_16793,N_15638);
xnor U18651 (N_18651,N_13461,N_13972);
nand U18652 (N_18652,N_15727,N_14724);
nor U18653 (N_18653,N_12989,N_14490);
and U18654 (N_18654,N_15648,N_16244);
and U18655 (N_18655,N_15093,N_17921);
or U18656 (N_18656,N_14593,N_14864);
and U18657 (N_18657,N_17594,N_15132);
or U18658 (N_18658,N_12411,N_13565);
xor U18659 (N_18659,N_16397,N_13927);
and U18660 (N_18660,N_12228,N_16824);
nor U18661 (N_18661,N_14553,N_16702);
and U18662 (N_18662,N_12509,N_16935);
nand U18663 (N_18663,N_17290,N_17746);
nor U18664 (N_18664,N_15957,N_14142);
or U18665 (N_18665,N_15658,N_15149);
nor U18666 (N_18666,N_12917,N_17988);
or U18667 (N_18667,N_12424,N_14775);
xor U18668 (N_18668,N_12798,N_12082);
nor U18669 (N_18669,N_15979,N_15501);
xor U18670 (N_18670,N_17697,N_12187);
nand U18671 (N_18671,N_16690,N_14955);
and U18672 (N_18672,N_17197,N_14502);
and U18673 (N_18673,N_14161,N_12243);
and U18674 (N_18674,N_15179,N_12364);
nand U18675 (N_18675,N_13161,N_17989);
nor U18676 (N_18676,N_16938,N_16834);
and U18677 (N_18677,N_12037,N_14737);
or U18678 (N_18678,N_14990,N_14304);
and U18679 (N_18679,N_12842,N_12021);
and U18680 (N_18680,N_17904,N_14464);
xor U18681 (N_18681,N_17219,N_16656);
xnor U18682 (N_18682,N_16538,N_14090);
xor U18683 (N_18683,N_14423,N_14220);
and U18684 (N_18684,N_16486,N_12419);
nor U18685 (N_18685,N_16003,N_12489);
nand U18686 (N_18686,N_15248,N_15836);
or U18687 (N_18687,N_16777,N_15017);
nor U18688 (N_18688,N_14560,N_17145);
xnor U18689 (N_18689,N_17785,N_14685);
nor U18690 (N_18690,N_15565,N_13732);
or U18691 (N_18691,N_14847,N_15494);
nor U18692 (N_18692,N_16772,N_12909);
nand U18693 (N_18693,N_15402,N_14586);
nand U18694 (N_18694,N_16150,N_13943);
and U18695 (N_18695,N_17853,N_16921);
and U18696 (N_18696,N_16058,N_17941);
and U18697 (N_18697,N_15573,N_15632);
xnor U18698 (N_18698,N_13166,N_15784);
and U18699 (N_18699,N_16543,N_13346);
or U18700 (N_18700,N_12699,N_16776);
or U18701 (N_18701,N_14838,N_12701);
nand U18702 (N_18702,N_16137,N_12862);
nor U18703 (N_18703,N_15056,N_12422);
nand U18704 (N_18704,N_16734,N_13910);
xor U18705 (N_18705,N_15237,N_14964);
nand U18706 (N_18706,N_12829,N_17111);
or U18707 (N_18707,N_16942,N_12872);
or U18708 (N_18708,N_16597,N_14254);
xnor U18709 (N_18709,N_14406,N_14648);
or U18710 (N_18710,N_14202,N_17136);
nor U18711 (N_18711,N_13012,N_13202);
and U18712 (N_18712,N_15396,N_15008);
and U18713 (N_18713,N_17245,N_12963);
nor U18714 (N_18714,N_15147,N_15076);
nor U18715 (N_18715,N_17475,N_13918);
xor U18716 (N_18716,N_15803,N_12985);
or U18717 (N_18717,N_16164,N_15446);
or U18718 (N_18718,N_15321,N_13588);
xnor U18719 (N_18719,N_17431,N_14852);
nand U18720 (N_18720,N_16814,N_17321);
nand U18721 (N_18721,N_15254,N_13122);
or U18722 (N_18722,N_16673,N_16633);
nand U18723 (N_18723,N_15805,N_15366);
and U18724 (N_18724,N_13124,N_14886);
nand U18725 (N_18725,N_13947,N_17314);
or U18726 (N_18726,N_12554,N_15027);
or U18727 (N_18727,N_16639,N_12246);
or U18728 (N_18728,N_15186,N_13183);
nand U18729 (N_18729,N_13899,N_12426);
nor U18730 (N_18730,N_17071,N_16294);
nor U18731 (N_18731,N_13566,N_16431);
or U18732 (N_18732,N_14988,N_13695);
and U18733 (N_18733,N_13374,N_12101);
nor U18734 (N_18734,N_17127,N_14888);
xnor U18735 (N_18735,N_12997,N_14073);
nor U18736 (N_18736,N_12077,N_17597);
and U18737 (N_18737,N_15916,N_17227);
or U18738 (N_18738,N_13784,N_17486);
and U18739 (N_18739,N_13406,N_12359);
nand U18740 (N_18740,N_13571,N_14417);
and U18741 (N_18741,N_12420,N_15580);
and U18742 (N_18742,N_13424,N_16726);
and U18743 (N_18743,N_12397,N_15983);
xnor U18744 (N_18744,N_17673,N_15296);
xor U18745 (N_18745,N_14840,N_16374);
xor U18746 (N_18746,N_17688,N_12289);
xnor U18747 (N_18747,N_15641,N_16094);
or U18748 (N_18748,N_16442,N_16009);
nor U18749 (N_18749,N_16056,N_16026);
nor U18750 (N_18750,N_12526,N_13164);
and U18751 (N_18751,N_12396,N_12342);
xnor U18752 (N_18752,N_17345,N_12856);
xor U18753 (N_18753,N_15338,N_16314);
xor U18754 (N_18754,N_12310,N_15253);
or U18755 (N_18755,N_17571,N_15520);
nand U18756 (N_18756,N_12940,N_12637);
or U18757 (N_18757,N_17234,N_15219);
or U18758 (N_18758,N_17041,N_16957);
xor U18759 (N_18759,N_12934,N_13889);
or U18760 (N_18760,N_14599,N_15153);
xnor U18761 (N_18761,N_16283,N_15847);
and U18762 (N_18762,N_13033,N_12720);
nor U18763 (N_18763,N_13094,N_14959);
nor U18764 (N_18764,N_16950,N_16974);
nand U18765 (N_18765,N_17458,N_12282);
or U18766 (N_18766,N_16055,N_14260);
nor U18767 (N_18767,N_15390,N_17315);
and U18768 (N_18768,N_12648,N_17329);
or U18769 (N_18769,N_17269,N_15517);
and U18770 (N_18770,N_12441,N_17369);
nand U18771 (N_18771,N_16928,N_12927);
or U18772 (N_18772,N_17074,N_17282);
nand U18773 (N_18773,N_16551,N_15206);
nand U18774 (N_18774,N_17672,N_14426);
nand U18775 (N_18775,N_15678,N_15749);
or U18776 (N_18776,N_14893,N_16352);
nand U18777 (N_18777,N_17338,N_16482);
nor U18778 (N_18778,N_14657,N_15777);
nand U18779 (N_18779,N_14751,N_13001);
and U18780 (N_18780,N_17512,N_12653);
nand U18781 (N_18781,N_13727,N_12495);
nor U18782 (N_18782,N_12454,N_12958);
and U18783 (N_18783,N_14029,N_17394);
xor U18784 (N_18784,N_14128,N_12938);
or U18785 (N_18785,N_12291,N_15169);
or U18786 (N_18786,N_12825,N_16148);
nand U18787 (N_18787,N_12696,N_14362);
nand U18788 (N_18788,N_13060,N_15381);
xnor U18789 (N_18789,N_14575,N_15165);
xnor U18790 (N_18790,N_13783,N_14635);
or U18791 (N_18791,N_13204,N_16453);
and U18792 (N_18792,N_13425,N_12881);
or U18793 (N_18793,N_16740,N_16315);
nand U18794 (N_18794,N_14541,N_12543);
xor U18795 (N_18795,N_15986,N_17516);
or U18796 (N_18796,N_12390,N_12605);
nand U18797 (N_18797,N_13873,N_12741);
and U18798 (N_18798,N_17713,N_12007);
nand U18799 (N_18799,N_13378,N_15739);
xnor U18800 (N_18800,N_13090,N_12593);
xnor U18801 (N_18801,N_13046,N_14650);
or U18802 (N_18802,N_15241,N_17063);
and U18803 (N_18803,N_12901,N_15586);
or U18804 (N_18804,N_12237,N_14382);
xnor U18805 (N_18805,N_12467,N_14308);
and U18806 (N_18806,N_13277,N_12012);
and U18807 (N_18807,N_12891,N_14595);
and U18808 (N_18808,N_17100,N_12822);
nor U18809 (N_18809,N_12011,N_15042);
or U18810 (N_18810,N_16126,N_15674);
or U18811 (N_18811,N_13365,N_12756);
and U18812 (N_18812,N_14037,N_14950);
nor U18813 (N_18813,N_15585,N_16927);
and U18814 (N_18814,N_13142,N_17656);
and U18815 (N_18815,N_15667,N_17095);
and U18816 (N_18816,N_17605,N_17305);
or U18817 (N_18817,N_15444,N_17851);
and U18818 (N_18818,N_13210,N_14316);
nand U18819 (N_18819,N_16879,N_12669);
nor U18820 (N_18820,N_13252,N_16483);
or U18821 (N_18821,N_12120,N_14867);
and U18822 (N_18822,N_17833,N_16985);
and U18823 (N_18823,N_13531,N_17279);
and U18824 (N_18824,N_14664,N_12786);
and U18825 (N_18825,N_13726,N_13752);
and U18826 (N_18826,N_12168,N_15301);
or U18827 (N_18827,N_12493,N_13348);
xnor U18828 (N_18828,N_14790,N_12001);
nor U18829 (N_18829,N_16960,N_16586);
xnor U18830 (N_18830,N_17798,N_15875);
nor U18831 (N_18831,N_12255,N_12976);
nor U18832 (N_18832,N_16364,N_16408);
and U18833 (N_18833,N_17991,N_15277);
nor U18834 (N_18834,N_15681,N_14624);
or U18835 (N_18835,N_17808,N_16332);
nand U18836 (N_18836,N_17384,N_12176);
nand U18837 (N_18837,N_15079,N_16818);
nor U18838 (N_18838,N_15063,N_17879);
xnor U18839 (N_18839,N_13790,N_15561);
or U18840 (N_18840,N_14300,N_17717);
nand U18841 (N_18841,N_15140,N_14725);
nor U18842 (N_18842,N_14673,N_16585);
or U18843 (N_18843,N_16416,N_13372);
xor U18844 (N_18844,N_13880,N_14399);
nand U18845 (N_18845,N_17320,N_16958);
or U18846 (N_18846,N_17848,N_15418);
nand U18847 (N_18847,N_14764,N_16699);
and U18848 (N_18848,N_15432,N_13168);
or U18849 (N_18849,N_14652,N_14703);
or U18850 (N_18850,N_15626,N_13709);
nor U18851 (N_18851,N_17529,N_12966);
or U18852 (N_18852,N_13218,N_13073);
xnor U18853 (N_18853,N_13689,N_12356);
or U18854 (N_18854,N_14991,N_14160);
nand U18855 (N_18855,N_16107,N_17467);
nand U18856 (N_18856,N_15035,N_13472);
nor U18857 (N_18857,N_13262,N_13846);
nand U18858 (N_18858,N_15168,N_16456);
nor U18859 (N_18859,N_16618,N_13446);
nand U18860 (N_18860,N_15108,N_15464);
and U18861 (N_18861,N_13440,N_13200);
nand U18862 (N_18862,N_14155,N_15317);
nand U18863 (N_18863,N_14483,N_12285);
nor U18864 (N_18864,N_12145,N_16269);
xnor U18865 (N_18865,N_17016,N_13799);
or U18866 (N_18866,N_17947,N_15884);
nor U18867 (N_18867,N_14434,N_16316);
nor U18868 (N_18868,N_17929,N_16717);
nand U18869 (N_18869,N_13572,N_13047);
xnor U18870 (N_18870,N_13473,N_14282);
xnor U18871 (N_18871,N_17980,N_12070);
and U18872 (N_18872,N_17184,N_16949);
or U18873 (N_18873,N_12979,N_13368);
and U18874 (N_18874,N_14665,N_12381);
xor U18875 (N_18875,N_14851,N_14019);
nand U18876 (N_18876,N_16220,N_13021);
nor U18877 (N_18877,N_12098,N_13969);
or U18878 (N_18878,N_14900,N_17427);
and U18879 (N_18879,N_16605,N_13786);
nor U18880 (N_18880,N_13024,N_17437);
nand U18881 (N_18881,N_13177,N_14755);
nand U18882 (N_18882,N_15247,N_16436);
nor U18883 (N_18883,N_16970,N_15888);
and U18884 (N_18884,N_16320,N_13246);
nor U18885 (N_18885,N_16419,N_12992);
and U18886 (N_18886,N_16792,N_12330);
and U18887 (N_18887,N_13907,N_15005);
and U18888 (N_18888,N_13862,N_17615);
xnor U18889 (N_18889,N_14400,N_12284);
xnor U18890 (N_18890,N_14614,N_12380);
nand U18891 (N_18891,N_15133,N_13496);
nor U18892 (N_18892,N_12523,N_17834);
and U18893 (N_18893,N_14892,N_14446);
nor U18894 (N_18894,N_15959,N_12155);
nand U18895 (N_18895,N_13130,N_17828);
xor U18896 (N_18896,N_17466,N_13761);
nor U18897 (N_18897,N_12475,N_17069);
and U18898 (N_18898,N_15212,N_16541);
xor U18899 (N_18899,N_17265,N_13641);
and U18900 (N_18900,N_17421,N_17084);
nor U18901 (N_18901,N_17211,N_12190);
or U18902 (N_18902,N_15902,N_12086);
and U18903 (N_18903,N_15187,N_12167);
or U18904 (N_18904,N_13029,N_13215);
or U18905 (N_18905,N_14223,N_14172);
and U18906 (N_18906,N_15834,N_12170);
xnor U18907 (N_18907,N_12793,N_16812);
and U18908 (N_18908,N_14574,N_15624);
or U18909 (N_18909,N_15671,N_16604);
nor U18910 (N_18910,N_14046,N_12404);
xor U18911 (N_18911,N_14390,N_17868);
or U18912 (N_18912,N_16444,N_12609);
or U18913 (N_18913,N_15275,N_15356);
xor U18914 (N_18914,N_15022,N_14017);
or U18915 (N_18915,N_15007,N_14863);
nor U18916 (N_18916,N_12921,N_16124);
xnor U18917 (N_18917,N_12616,N_13255);
or U18918 (N_18918,N_15082,N_12217);
and U18919 (N_18919,N_17564,N_15374);
and U18920 (N_18920,N_14070,N_17244);
nand U18921 (N_18921,N_16549,N_13076);
xor U18922 (N_18922,N_17577,N_14059);
nand U18923 (N_18923,N_15111,N_12196);
nand U18924 (N_18924,N_14576,N_15210);
or U18925 (N_18925,N_13718,N_14984);
or U18926 (N_18926,N_17328,N_13077);
xor U18927 (N_18927,N_16140,N_14945);
nand U18928 (N_18928,N_16199,N_12192);
xor U18929 (N_18929,N_17377,N_13179);
nand U18930 (N_18930,N_13537,N_12418);
nand U18931 (N_18931,N_16767,N_16226);
or U18932 (N_18932,N_17508,N_12207);
nand U18933 (N_18933,N_15537,N_17066);
xnor U18934 (N_18934,N_13092,N_16261);
nand U18935 (N_18935,N_16908,N_14205);
and U18936 (N_18936,N_14384,N_12416);
or U18937 (N_18937,N_13893,N_16529);
and U18938 (N_18938,N_16473,N_13751);
nand U18939 (N_18939,N_17910,N_15637);
xnor U18940 (N_18940,N_15831,N_14397);
nand U18941 (N_18941,N_13579,N_14396);
nor U18942 (N_18942,N_15800,N_14186);
nand U18943 (N_18943,N_13787,N_14333);
nand U18944 (N_18944,N_16982,N_12852);
and U18945 (N_18945,N_15904,N_13683);
xor U18946 (N_18946,N_15867,N_12580);
or U18947 (N_18947,N_17954,N_13116);
and U18948 (N_18948,N_12581,N_16463);
nand U18949 (N_18949,N_16808,N_13774);
or U18950 (N_18950,N_14510,N_17644);
or U18951 (N_18951,N_15571,N_15783);
or U18952 (N_18952,N_16701,N_17831);
or U18953 (N_18953,N_15397,N_16481);
xnor U18954 (N_18954,N_12869,N_15955);
nand U18955 (N_18955,N_15411,N_17085);
nand U18956 (N_18956,N_16423,N_16964);
xnor U18957 (N_18957,N_16122,N_15440);
nand U18958 (N_18958,N_16514,N_17680);
and U18959 (N_18959,N_12347,N_13436);
and U18960 (N_18960,N_12724,N_16293);
nand U18961 (N_18961,N_15074,N_12857);
or U18962 (N_18962,N_16046,N_13163);
nand U18963 (N_18963,N_12385,N_17769);
or U18964 (N_18964,N_14745,N_14135);
xnor U18965 (N_18965,N_17418,N_14905);
and U18966 (N_18966,N_15865,N_17835);
xnor U18967 (N_18967,N_12321,N_14199);
xnor U18968 (N_18968,N_12080,N_14910);
nand U18969 (N_18969,N_17637,N_15635);
nor U18970 (N_18970,N_14452,N_12480);
xnor U18971 (N_18971,N_16563,N_17009);
and U18972 (N_18972,N_15438,N_16961);
nor U18973 (N_18973,N_15048,N_14957);
nor U18974 (N_18974,N_12113,N_15599);
or U18975 (N_18975,N_14519,N_15280);
nand U18976 (N_18976,N_15391,N_17162);
and U18977 (N_18977,N_14395,N_15403);
or U18978 (N_18978,N_15004,N_14066);
and U18979 (N_18979,N_14092,N_15482);
xor U18980 (N_18980,N_17408,N_17048);
nor U18981 (N_18981,N_12764,N_14492);
and U18982 (N_18982,N_15589,N_13700);
and U18983 (N_18983,N_14702,N_15242);
or U18984 (N_18984,N_16531,N_16429);
nand U18985 (N_18985,N_13674,N_13158);
and U18986 (N_18986,N_17013,N_17576);
nor U18987 (N_18987,N_13665,N_12401);
xor U18988 (N_18988,N_15601,N_17346);
xor U18989 (N_18989,N_14967,N_16441);
or U18990 (N_18990,N_14935,N_17373);
nor U18991 (N_18991,N_17053,N_14436);
or U18992 (N_18992,N_14942,N_15788);
xnor U18993 (N_18993,N_12646,N_12023);
nor U18994 (N_18994,N_13386,N_12632);
or U18995 (N_18995,N_15793,N_16704);
nor U18996 (N_18996,N_17003,N_12032);
and U18997 (N_18997,N_15887,N_17715);
nor U18998 (N_18998,N_13797,N_15554);
and U18999 (N_18999,N_17395,N_13542);
or U19000 (N_19000,N_17914,N_16644);
xnor U19001 (N_19001,N_14527,N_17190);
xnor U19002 (N_19002,N_15892,N_17619);
or U19003 (N_19003,N_17286,N_14996);
nand U19004 (N_19004,N_12537,N_12727);
or U19005 (N_19005,N_16247,N_12248);
nor U19006 (N_19006,N_15630,N_16738);
and U19007 (N_19007,N_17613,N_15408);
and U19008 (N_19008,N_15675,N_13118);
nand U19009 (N_19009,N_13062,N_16967);
and U19010 (N_19010,N_15692,N_13173);
and U19011 (N_19011,N_17490,N_13303);
nand U19012 (N_19012,N_13550,N_14889);
or U19013 (N_19013,N_14898,N_14820);
or U19014 (N_19014,N_15347,N_16560);
xor U19015 (N_19015,N_16655,N_16920);
nand U19016 (N_19016,N_12096,N_15874);
and U19017 (N_19017,N_15044,N_12433);
or U19018 (N_19018,N_15721,N_15746);
nor U19019 (N_19019,N_15459,N_12682);
nand U19020 (N_19020,N_12571,N_12913);
xor U19021 (N_19021,N_17049,N_12457);
or U19022 (N_19022,N_14243,N_13423);
xor U19023 (N_19023,N_15891,N_12322);
and U19024 (N_19024,N_15011,N_16647);
and U19025 (N_19025,N_14717,N_16358);
nor U19026 (N_19026,N_16936,N_15855);
nor U19027 (N_19027,N_16752,N_16678);
nand U19028 (N_19028,N_13617,N_12517);
xnor U19029 (N_19029,N_14683,N_13731);
or U19030 (N_19030,N_16632,N_16194);
and U19031 (N_19031,N_17526,N_12262);
or U19032 (N_19032,N_15544,N_14549);
or U19033 (N_19033,N_14283,N_16864);
xor U19034 (N_19034,N_14834,N_12999);
xor U19035 (N_19035,N_13581,N_17365);
nor U19036 (N_19036,N_17538,N_15101);
nand U19037 (N_19037,N_13068,N_12516);
and U19038 (N_19038,N_12933,N_14409);
nand U19039 (N_19039,N_14035,N_14237);
nand U19040 (N_19040,N_16883,N_12315);
or U19041 (N_19041,N_14248,N_12326);
xor U19042 (N_19042,N_12518,N_17107);
and U19043 (N_19043,N_17355,N_12740);
xnor U19044 (N_19044,N_14378,N_14918);
or U19045 (N_19045,N_12613,N_17677);
or U19046 (N_19046,N_14330,N_12598);
xor U19047 (N_19047,N_12136,N_12423);
and U19048 (N_19048,N_15203,N_17795);
xnor U19049 (N_19049,N_14015,N_12542);
and U19050 (N_19050,N_14658,N_12238);
nand U19051 (N_19051,N_14407,N_17984);
and U19052 (N_19052,N_14600,N_13613);
and U19053 (N_19053,N_15089,N_12784);
nor U19054 (N_19054,N_13964,N_13165);
nand U19055 (N_19055,N_16695,N_17420);
or U19056 (N_19056,N_17590,N_14480);
nand U19057 (N_19057,N_16544,N_16582);
or U19058 (N_19058,N_13493,N_15730);
nand U19059 (N_19059,N_17492,N_15701);
nor U19060 (N_19060,N_17297,N_17089);
or U19061 (N_19061,N_14226,N_15524);
xor U19062 (N_19062,N_14528,N_16789);
xnor U19063 (N_19063,N_12393,N_12804);
and U19064 (N_19064,N_17167,N_16222);
nor U19065 (N_19065,N_12726,N_14082);
nor U19066 (N_19066,N_16606,N_15405);
xnor U19067 (N_19067,N_14691,N_16091);
nand U19068 (N_19068,N_12071,N_13356);
and U19069 (N_19069,N_17001,N_14922);
nor U19070 (N_19070,N_12738,N_13450);
or U19071 (N_19071,N_12132,N_16245);
and U19072 (N_19072,N_15223,N_15769);
and U19073 (N_19073,N_15462,N_13692);
and U19074 (N_19074,N_16939,N_14093);
nor U19075 (N_19075,N_12923,N_12206);
and U19076 (N_19076,N_17060,N_16440);
and U19077 (N_19077,N_13148,N_13811);
xor U19078 (N_19078,N_14120,N_16882);
nand U19079 (N_19079,N_13803,N_16826);
and U19080 (N_19080,N_15666,N_16664);
and U19081 (N_19081,N_15013,N_15617);
nand U19082 (N_19082,N_17347,N_13358);
nor U19083 (N_19083,N_13325,N_17090);
xor U19084 (N_19084,N_12874,N_14211);
nor U19085 (N_19085,N_12672,N_13620);
or U19086 (N_19086,N_17691,N_16532);
or U19087 (N_19087,N_13831,N_17745);
and U19088 (N_19088,N_17472,N_17883);
xnor U19089 (N_19089,N_15852,N_15131);
and U19090 (N_19090,N_14455,N_12486);
and U19091 (N_19091,N_17311,N_15882);
and U19092 (N_19092,N_13557,N_13719);
nand U19093 (N_19093,N_16739,N_15612);
xor U19094 (N_19094,N_17707,N_17892);
or U19095 (N_19095,N_13232,N_14744);
nor U19096 (N_19096,N_14934,N_17609);
nand U19097 (N_19097,N_15188,N_16197);
and U19098 (N_19098,N_14545,N_17283);
nand U19099 (N_19099,N_14529,N_14456);
and U19100 (N_19100,N_17669,N_13832);
nand U19101 (N_19101,N_15016,N_15000);
or U19102 (N_19102,N_12389,N_14104);
or U19103 (N_19103,N_17563,N_12876);
nor U19104 (N_19104,N_12346,N_13569);
xor U19105 (N_19105,N_14887,N_13729);
nor U19106 (N_19106,N_15150,N_16510);
nor U19107 (N_19107,N_12815,N_13697);
xnor U19108 (N_19108,N_13701,N_17039);
and U19109 (N_19109,N_16749,N_15753);
or U19110 (N_19110,N_16631,N_14651);
or U19111 (N_19111,N_12557,N_16029);
nor U19112 (N_19112,N_12362,N_13544);
and U19113 (N_19113,N_17462,N_12969);
and U19114 (N_19114,N_14700,N_13753);
nand U19115 (N_19115,N_15759,N_17930);
nor U19116 (N_19116,N_12611,N_15545);
nor U19117 (N_19117,N_17180,N_12265);
and U19118 (N_19118,N_16764,N_14359);
or U19119 (N_19119,N_13413,N_16630);
xnor U19120 (N_19120,N_17446,N_15258);
and U19121 (N_19121,N_13555,N_12676);
nand U19122 (N_19122,N_17416,N_12811);
nand U19123 (N_19123,N_17514,N_16426);
or U19124 (N_19124,N_16112,N_14698);
nor U19125 (N_19125,N_16249,N_13539);
nor U19126 (N_19126,N_16999,N_12172);
or U19127 (N_19127,N_14047,N_16674);
nor U19128 (N_19128,N_16887,N_14763);
xnor U19129 (N_19129,N_14693,N_14676);
or U19130 (N_19130,N_12535,N_16008);
and U19131 (N_19131,N_14656,N_12174);
nor U19132 (N_19132,N_14471,N_13680);
or U19133 (N_19133,N_16128,N_12947);
or U19134 (N_19134,N_17151,N_15535);
nor U19135 (N_19135,N_12331,N_15092);
and U19136 (N_19136,N_15302,N_13082);
xor U19137 (N_19137,N_16391,N_15291);
or U19138 (N_19138,N_14603,N_13872);
xor U19139 (N_19139,N_13775,N_16837);
and U19140 (N_19140,N_17260,N_13269);
and U19141 (N_19141,N_14095,N_12808);
nand U19142 (N_19142,N_13871,N_16268);
and U19143 (N_19143,N_12271,N_17246);
nand U19144 (N_19144,N_13049,N_15477);
and U19145 (N_19145,N_16895,N_16787);
nor U19146 (N_19146,N_12988,N_13696);
and U19147 (N_19147,N_16709,N_16558);
xor U19148 (N_19148,N_17375,N_12269);
nand U19149 (N_19149,N_15728,N_14259);
xnor U19150 (N_19150,N_12778,N_12208);
nand U19151 (N_19151,N_15861,N_15058);
and U19152 (N_19152,N_14021,N_16583);
nor U19153 (N_19153,N_16802,N_13182);
or U19154 (N_19154,N_15385,N_17028);
and U19155 (N_19155,N_16182,N_16372);
or U19156 (N_19156,N_17449,N_13089);
xor U19157 (N_19157,N_12247,N_16943);
and U19158 (N_19158,N_14961,N_15895);
xor U19159 (N_19159,N_15698,N_17172);
or U19160 (N_19160,N_17580,N_17544);
or U19161 (N_19161,N_13107,N_14558);
nand U19162 (N_19162,N_12470,N_15146);
nor U19163 (N_19163,N_17905,N_13794);
nand U19164 (N_19164,N_16963,N_13631);
nand U19165 (N_19165,N_13517,N_13540);
or U19166 (N_19166,N_15903,N_13882);
nand U19167 (N_19167,N_13404,N_15222);
xor U19168 (N_19168,N_15328,N_16060);
nor U19169 (N_19169,N_13454,N_14628);
nor U19170 (N_19170,N_14981,N_17522);
nand U19171 (N_19171,N_16042,N_15259);
nand U19172 (N_19172,N_14214,N_16951);
nor U19173 (N_19173,N_16064,N_14338);
and U19174 (N_19174,N_15550,N_15523);
or U19175 (N_19175,N_14690,N_16337);
or U19176 (N_19176,N_15755,N_14387);
and U19177 (N_19177,N_16231,N_14531);
nor U19178 (N_19178,N_15828,N_13273);
xnor U19179 (N_19179,N_17101,N_16925);
xor U19180 (N_19180,N_16346,N_15672);
or U19181 (N_19181,N_13817,N_12383);
nor U19182 (N_19182,N_12107,N_16434);
nor U19183 (N_19183,N_12354,N_17598);
or U19184 (N_19184,N_14468,N_17887);
xnor U19185 (N_19185,N_13212,N_12165);
nor U19186 (N_19186,N_12297,N_12905);
nor U19187 (N_19187,N_13268,N_13830);
nand U19188 (N_19188,N_14761,N_15476);
xnor U19189 (N_19189,N_13293,N_17441);
nor U19190 (N_19190,N_12721,N_12279);
xnor U19191 (N_19191,N_17596,N_17725);
and U19192 (N_19192,N_13236,N_15989);
and U19193 (N_19193,N_14561,N_15257);
and U19194 (N_19194,N_12946,N_13650);
nor U19195 (N_19195,N_16896,N_13594);
or U19196 (N_19196,N_12974,N_17957);
or U19197 (N_19197,N_14925,N_14680);
nor U19198 (N_19198,N_17877,N_17632);
or U19199 (N_19199,N_17962,N_17444);
or U19200 (N_19200,N_17148,N_16359);
and U19201 (N_19201,N_14122,N_17574);
nor U19202 (N_19202,N_13883,N_15341);
nor U19203 (N_19203,N_16401,N_16891);
nor U19204 (N_19204,N_14978,N_16233);
nand U19205 (N_19205,N_14753,N_17203);
and U19206 (N_19206,N_16457,N_12069);
or U19207 (N_19207,N_12343,N_16348);
and U19208 (N_19208,N_17335,N_12512);
or U19209 (N_19209,N_12345,N_16037);
and U19210 (N_19210,N_17888,N_15948);
xnor U19211 (N_19211,N_15613,N_12995);
or U19212 (N_19212,N_13267,N_15095);
and U19213 (N_19213,N_17217,N_13266);
and U19214 (N_19214,N_13216,N_13335);
or U19215 (N_19215,N_16158,N_13520);
and U19216 (N_19216,N_17671,N_12327);
nand U19217 (N_19217,N_15040,N_16360);
and U19218 (N_19218,N_12036,N_14629);
or U19219 (N_19219,N_15859,N_16975);
nor U19220 (N_19220,N_14096,N_13249);
and U19221 (N_19221,N_12055,N_14133);
xnor U19222 (N_19222,N_14688,N_14067);
xnor U19223 (N_19223,N_15596,N_16708);
and U19224 (N_19224,N_14042,N_15377);
and U19225 (N_19225,N_13415,N_16147);
and U19226 (N_19226,N_16210,N_12150);
xnor U19227 (N_19227,N_17057,N_17870);
or U19228 (N_19228,N_17958,N_13960);
nand U19229 (N_19229,N_12337,N_14865);
or U19230 (N_19230,N_17836,N_12638);
and U19231 (N_19231,N_15344,N_13682);
nor U19232 (N_19232,N_15285,N_15180);
and U19233 (N_19233,N_17005,N_16572);
nor U19234 (N_19234,N_12008,N_14728);
or U19235 (N_19235,N_14543,N_14371);
and U19236 (N_19236,N_12711,N_15914);
nor U19237 (N_19237,N_12339,N_13856);
or U19238 (N_19238,N_16086,N_14299);
nand U19239 (N_19239,N_14297,N_13261);
or U19240 (N_19240,N_13828,N_15714);
nor U19241 (N_19241,N_16146,N_17912);
or U19242 (N_19242,N_15558,N_15604);
or U19243 (N_19243,N_15468,N_16275);
or U19244 (N_19244,N_16484,N_13136);
nor U19245 (N_19245,N_12251,N_12748);
xnor U19246 (N_19246,N_14138,N_14127);
or U19247 (N_19247,N_12534,N_14590);
xor U19248 (N_19248,N_14204,N_13892);
or U19249 (N_19249,N_16913,N_16382);
nor U19250 (N_19250,N_12814,N_14164);
and U19251 (N_19251,N_15159,N_14345);
nand U19252 (N_19252,N_15530,N_15555);
or U19253 (N_19253,N_17867,N_15741);
nor U19254 (N_19254,N_13922,N_13859);
or U19255 (N_19255,N_16506,N_16849);
or U19256 (N_19256,N_17731,N_12594);
xor U19257 (N_19257,N_12892,N_16021);
or U19258 (N_19258,N_14240,N_12965);
xor U19259 (N_19259,N_15546,N_12750);
xor U19260 (N_19260,N_12955,N_13619);
nor U19261 (N_19261,N_14491,N_12214);
nor U19262 (N_19262,N_14585,N_13634);
nand U19263 (N_19263,N_17639,N_12757);
and U19264 (N_19264,N_14876,N_12146);
xnor U19265 (N_19265,N_13845,N_17863);
nand U19266 (N_19266,N_17106,N_14100);
xnor U19267 (N_19267,N_14504,N_15577);
xor U19268 (N_19268,N_14375,N_16889);
and U19269 (N_19269,N_14477,N_13065);
xor U19270 (N_19270,N_14307,N_16110);
xor U19271 (N_19271,N_14537,N_12437);
nand U19272 (N_19272,N_14512,N_16981);
xor U19273 (N_19273,N_12188,N_15668);
nand U19274 (N_19274,N_17595,N_13375);
or U19275 (N_19275,N_15958,N_15974);
or U19276 (N_19276,N_16712,N_14581);
nand U19277 (N_19277,N_13791,N_16216);
nor U19278 (N_19278,N_15346,N_13108);
nand U19279 (N_19279,N_15414,N_15309);
xor U19280 (N_19280,N_17372,N_13157);
or U19281 (N_19281,N_17813,N_16304);
or U19282 (N_19282,N_17881,N_14602);
nand U19283 (N_19283,N_13147,N_15123);
and U19284 (N_19284,N_17504,N_12626);
nor U19285 (N_19285,N_14331,N_13754);
or U19286 (N_19286,N_14145,N_16134);
and U19287 (N_19287,N_15702,N_15333);
or U19288 (N_19288,N_15533,N_17903);
or U19289 (N_19289,N_13150,N_14425);
or U19290 (N_19290,N_16089,N_17520);
nand U19291 (N_19291,N_15392,N_13605);
and U19292 (N_19292,N_12827,N_17030);
xor U19293 (N_19293,N_15213,N_15742);
xor U19294 (N_19294,N_13598,N_12375);
nand U19295 (N_19295,N_15127,N_16610);
nand U19296 (N_19296,N_15631,N_17133);
xor U19297 (N_19297,N_16313,N_13946);
xnor U19298 (N_19298,N_12332,N_15595);
and U19299 (N_19299,N_17065,N_16203);
nand U19300 (N_19300,N_17192,N_16766);
and U19301 (N_19301,N_13195,N_15435);
xor U19302 (N_19302,N_17705,N_15731);
and U19303 (N_19303,N_17814,N_15053);
or U19304 (N_19304,N_16652,N_15706);
nand U19305 (N_19305,N_13508,N_13175);
xor U19306 (N_19306,N_14180,N_15527);
xor U19307 (N_19307,N_16524,N_13257);
nand U19308 (N_19308,N_14111,N_13483);
xor U19309 (N_19309,N_14131,N_17966);
or U19310 (N_19310,N_16653,N_13070);
nor U19311 (N_19311,N_13272,N_14931);
and U19312 (N_19312,N_15960,N_16807);
and U19313 (N_19313,N_14011,N_16911);
and U19314 (N_19314,N_12840,N_16400);
and U19315 (N_19315,N_13755,N_12919);
nand U19316 (N_19316,N_17502,N_12558);
nand U19317 (N_19317,N_17846,N_16455);
and U19318 (N_19318,N_16519,N_12621);
xor U19319 (N_19319,N_14713,N_13135);
xor U19320 (N_19320,N_12693,N_13035);
or U19321 (N_19321,N_16569,N_15893);
nor U19322 (N_19322,N_15426,N_15579);
nand U19323 (N_19323,N_17528,N_15991);
xor U19324 (N_19324,N_16237,N_16525);
or U19325 (N_19325,N_13602,N_12059);
xor U19326 (N_19326,N_13914,N_12293);
nor U19327 (N_19327,N_17390,N_13626);
xnor U19328 (N_19328,N_15505,N_15393);
or U19329 (N_19329,N_16683,N_13428);
xor U19330 (N_19330,N_14983,N_17549);
nor U19331 (N_19331,N_17354,N_14773);
nand U19332 (N_19332,N_14671,N_16836);
and U19333 (N_19333,N_16505,N_15872);
or U19334 (N_19334,N_12832,N_12216);
nor U19335 (N_19335,N_14550,N_12932);
and U19336 (N_19336,N_15956,N_17530);
and U19337 (N_19337,N_17511,N_17660);
xnor U19338 (N_19338,N_16131,N_17161);
xor U19339 (N_19339,N_13816,N_15756);
nor U19340 (N_19340,N_12705,N_17953);
xor U19341 (N_19341,N_13227,N_12448);
or U19342 (N_19342,N_15031,N_12263);
or U19343 (N_19343,N_12152,N_12056);
nand U19344 (N_19344,N_15718,N_15961);
and U19345 (N_19345,N_13587,N_17599);
or U19346 (N_19346,N_13884,N_16402);
or U19347 (N_19347,N_17963,N_17191);
and U19348 (N_19348,N_16259,N_17010);
and U19349 (N_19349,N_12858,N_13263);
xnor U19350 (N_19350,N_17684,N_16873);
nand U19351 (N_19351,N_14958,N_13702);
and U19352 (N_19352,N_14625,N_16155);
xor U19353 (N_19353,N_17334,N_12896);
nand U19354 (N_19354,N_13145,N_14811);
nor U19355 (N_19355,N_14277,N_14722);
or U19356 (N_19356,N_16813,N_16870);
xor U19357 (N_19357,N_12123,N_16273);
xnor U19358 (N_19358,N_14780,N_12617);
or U19359 (N_19359,N_17696,N_16123);
and U19360 (N_19360,N_14444,N_16335);
and U19361 (N_19361,N_14791,N_12357);
xor U19362 (N_19362,N_14171,N_14320);
or U19363 (N_19363,N_17575,N_13387);
nand U19364 (N_19364,N_16856,N_12599);
nor U19365 (N_19365,N_13030,N_16721);
nor U19366 (N_19366,N_17761,N_15471);
nor U19367 (N_19367,N_15033,N_13486);
and U19368 (N_19368,N_13541,N_17076);
or U19369 (N_19369,N_17366,N_17661);
xor U19370 (N_19370,N_12173,N_15162);
or U19371 (N_19371,N_16321,N_13958);
or U19372 (N_19372,N_14506,N_15557);
xor U19373 (N_19373,N_13780,N_14771);
xor U19374 (N_19374,N_14474,N_17032);
nor U19375 (N_19375,N_12491,N_17064);
and U19376 (N_19376,N_15908,N_14169);
and U19377 (N_19377,N_15235,N_16845);
nand U19378 (N_19378,N_17079,N_13950);
xnor U19379 (N_19379,N_16495,N_13389);
and U19380 (N_19380,N_13645,N_13396);
nor U19381 (N_19381,N_17235,N_12213);
and U19382 (N_19382,N_12604,N_15238);
nor U19383 (N_19383,N_15688,N_17517);
nor U19384 (N_19384,N_14807,N_17379);
or U19385 (N_19385,N_17927,N_15387);
and U19386 (N_19386,N_12763,N_16771);
and U19387 (N_19387,N_15823,N_15656);
and U19388 (N_19388,N_15369,N_12918);
nand U19389 (N_19389,N_12078,N_15936);
xnor U19390 (N_19390,N_16595,N_12519);
nand U19391 (N_19391,N_13815,N_17154);
xor U19392 (N_19392,N_14518,N_13672);
or U19393 (N_19393,N_15104,N_13600);
nand U19394 (N_19394,N_14756,N_15773);
nor U19395 (N_19395,N_13075,N_17481);
nor U19396 (N_19396,N_17489,N_16376);
and U19397 (N_19397,N_17690,N_16479);
xnor U19398 (N_19398,N_13360,N_16040);
xnor U19399 (N_19399,N_15659,N_16476);
and U19400 (N_19400,N_14218,N_16496);
nand U19401 (N_19401,N_17459,N_15067);
nand U19402 (N_19402,N_13298,N_13220);
and U19403 (N_19403,N_15899,N_13079);
xor U19404 (N_19404,N_14008,N_14157);
or U19405 (N_19405,N_13484,N_15466);
nor U19406 (N_19406,N_12767,N_15682);
and U19407 (N_19407,N_14469,N_16201);
xnor U19408 (N_19408,N_16369,N_14857);
or U19409 (N_19409,N_14638,N_16657);
or U19410 (N_19410,N_15890,N_17040);
xor U19411 (N_19411,N_14380,N_17274);
xor U19412 (N_19412,N_12451,N_15830);
nand U19413 (N_19413,N_17348,N_14678);
xnor U19414 (N_19414,N_13549,N_13253);
and U19415 (N_19415,N_15204,N_15225);
nor U19416 (N_19416,N_14485,N_15764);
nor U19417 (N_19417,N_12129,N_17170);
and U19418 (N_19418,N_12954,N_16357);
xnor U19419 (N_19419,N_16228,N_13944);
and U19420 (N_19420,N_13481,N_17803);
xor U19421 (N_19421,N_15804,N_16196);
nor U19422 (N_19422,N_12360,N_16867);
or U19423 (N_19423,N_16032,N_14742);
or U19424 (N_19424,N_15060,N_13901);
nand U19425 (N_19425,N_12241,N_14181);
and U19426 (N_19426,N_17160,N_12471);
and U19427 (N_19427,N_13661,N_16262);
xnor U19428 (N_19428,N_14151,N_16930);
xor U19429 (N_19429,N_12781,N_16298);
nor U19430 (N_19430,N_17944,N_17143);
or U19431 (N_19431,N_17509,N_15500);
xnor U19432 (N_19432,N_14429,N_13225);
xor U19433 (N_19433,N_15789,N_17797);
and U19434 (N_19434,N_12504,N_12860);
and U19435 (N_19435,N_16301,N_14110);
nor U19436 (N_19436,N_12931,N_15543);
and U19437 (N_19437,N_12841,N_13088);
and U19438 (N_19438,N_17436,N_13995);
nor U19439 (N_19439,N_15458,N_14031);
xor U19440 (N_19440,N_16277,N_13576);
and U19441 (N_19441,N_17796,N_12133);
or U19442 (N_19442,N_12257,N_14617);
and U19443 (N_19443,N_13621,N_13489);
or U19444 (N_19444,N_13896,N_15323);
xor U19445 (N_19445,N_17059,N_14989);
nor U19446 (N_19446,N_16666,N_16884);
and U19447 (N_19447,N_14623,N_12839);
nor U19448 (N_19448,N_14882,N_16902);
nor U19449 (N_19449,N_13758,N_17017);
and U19450 (N_19450,N_17336,N_13045);
or U19451 (N_19451,N_17374,N_15508);
and U19452 (N_19452,N_12144,N_12603);
nand U19453 (N_19453,N_17055,N_17023);
nor U19454 (N_19454,N_12620,N_13949);
or U19455 (N_19455,N_12439,N_15507);
nand U19456 (N_19456,N_12060,N_15620);
nor U19457 (N_19457,N_16417,N_17308);
xor U19458 (N_19458,N_13915,N_14501);
nand U19459 (N_19459,N_17433,N_16628);
or U19460 (N_19460,N_14642,N_12267);
nand U19461 (N_19461,N_17087,N_15695);
nor U19462 (N_19462,N_17452,N_12092);
xor U19463 (N_19463,N_15929,N_12801);
nand U19464 (N_19464,N_13504,N_12341);
or U19465 (N_19465,N_12873,N_12560);
and U19466 (N_19466,N_14919,N_13895);
nand U19467 (N_19467,N_17805,N_13469);
or U19468 (N_19468,N_17970,N_16159);
nand U19469 (N_19469,N_12952,N_13979);
nor U19470 (N_19470,N_12792,N_12957);
nor U19471 (N_19471,N_17402,N_13848);
nand U19472 (N_19472,N_17588,N_15735);
or U19473 (N_19473,N_15794,N_13981);
or U19474 (N_19474,N_16754,N_13777);
nor U19475 (N_19475,N_13016,N_15640);
nand U19476 (N_19476,N_16629,N_12408);
or U19477 (N_19477,N_13304,N_12106);
xnor U19478 (N_19478,N_14816,N_17430);
and U19479 (N_19479,N_13064,N_16264);
or U19480 (N_19480,N_13824,N_14933);
nor U19481 (N_19481,N_12270,N_12244);
nand U19482 (N_19482,N_17132,N_14622);
nand U19483 (N_19483,N_17168,N_12358);
nor U19484 (N_19484,N_17787,N_15866);
nand U19485 (N_19485,N_17138,N_12680);
nand U19486 (N_19486,N_16368,N_13388);
xor U19487 (N_19487,N_12733,N_14419);
nand U19488 (N_19488,N_15325,N_15288);
nor U19489 (N_19489,N_14666,N_12264);
nor U19490 (N_19490,N_14064,N_17306);
nor U19491 (N_19491,N_17011,N_16485);
nor U19492 (N_19492,N_13478,N_12033);
nand U19493 (N_19493,N_17723,N_14255);
nor U19494 (N_19494,N_17451,N_17638);
or U19495 (N_19495,N_17233,N_15281);
or U19496 (N_19496,N_16289,N_17852);
and U19497 (N_19497,N_12430,N_17537);
nand U19498 (N_19498,N_17744,N_15711);
and U19499 (N_19499,N_12837,N_16937);
xnor U19500 (N_19500,N_12624,N_17789);
and U19501 (N_19501,N_14608,N_16072);
and U19502 (N_19502,N_13437,N_14976);
or U19503 (N_19503,N_17676,N_13199);
nand U19504 (N_19504,N_15703,N_13818);
nor U19505 (N_19505,N_15357,N_12260);
and U19506 (N_19506,N_17592,N_13666);
and U19507 (N_19507,N_15526,N_13091);
xnor U19508 (N_19508,N_15428,N_17118);
nand U19509 (N_19509,N_16373,N_17218);
xnor U19510 (N_19510,N_12079,N_12015);
nor U19511 (N_19511,N_14770,N_16497);
xnor U19512 (N_19512,N_16135,N_15747);
nand U19513 (N_19513,N_16804,N_15361);
xor U19514 (N_19514,N_17367,N_17276);
nand U19515 (N_19515,N_14244,N_14579);
xnor U19516 (N_19516,N_12796,N_13867);
and U19517 (N_19517,N_15192,N_17298);
and U19518 (N_19518,N_13022,N_14296);
xnor U19519 (N_19519,N_17166,N_17483);
nand U19520 (N_19520,N_14451,N_14153);
nand U19521 (N_19521,N_16349,N_12805);
and U19522 (N_19522,N_12717,N_14102);
xor U19523 (N_19523,N_17547,N_17816);
or U19524 (N_19524,N_17603,N_16186);
xor U19525 (N_19525,N_15655,N_13330);
nand U19526 (N_19526,N_13031,N_15582);
or U19527 (N_19527,N_13887,N_16851);
xnor U19528 (N_19528,N_16968,N_16085);
xnor U19529 (N_19529,N_15653,N_14309);
and U19530 (N_19530,N_16438,N_17763);
and U19531 (N_19531,N_16119,N_13951);
nor U19532 (N_19532,N_17546,N_15813);
or U19533 (N_19533,N_12949,N_13320);
nand U19534 (N_19534,N_13309,N_16047);
xnor U19535 (N_19535,N_14508,N_16815);
nor U19536 (N_19536,N_14116,N_12643);
nor U19537 (N_19537,N_16946,N_13967);
and U19538 (N_19538,N_14995,N_12670);
or U19539 (N_19539,N_14965,N_13431);
xor U19540 (N_19540,N_12232,N_15336);
or U19541 (N_19541,N_14523,N_14594);
or U19542 (N_19542,N_17722,N_12735);
nor U19543 (N_19543,N_13186,N_12134);
or U19544 (N_19544,N_12743,N_13455);
xor U19545 (N_19545,N_13781,N_13917);
or U19546 (N_19546,N_12634,N_16471);
nand U19547 (N_19547,N_16868,N_16565);
or U19548 (N_19548,N_17873,N_16061);
xnor U19549 (N_19549,N_16637,N_17843);
nand U19550 (N_19550,N_17099,N_12410);
nand U19551 (N_19551,N_12465,N_16559);
xnor U19552 (N_19552,N_17572,N_13300);
nand U19553 (N_19553,N_17046,N_17181);
and U19554 (N_19554,N_15540,N_17385);
or U19555 (N_19555,N_14802,N_13477);
and U19556 (N_19556,N_17973,N_13499);
nand U19557 (N_19557,N_17655,N_14712);
or U19558 (N_19558,N_17476,N_12950);
or U19559 (N_19559,N_15969,N_14024);
xor U19560 (N_19560,N_14839,N_13101);
and U19561 (N_19561,N_16375,N_16390);
and U19562 (N_19562,N_12484,N_12004);
and U19563 (N_19563,N_12736,N_16660);
nand U19564 (N_19564,N_13694,N_14443);
nand U19565 (N_19565,N_12141,N_15615);
or U19566 (N_19566,N_13638,N_12737);
nor U19567 (N_19567,N_15419,N_12038);
xnor U19568 (N_19568,N_13324,N_12446);
nor U19569 (N_19569,N_12610,N_12126);
xor U19570 (N_19570,N_15091,N_15176);
and U19571 (N_19571,N_12240,N_14540);
and U19572 (N_19572,N_12499,N_15937);
or U19573 (N_19573,N_16345,N_16744);
nor U19574 (N_19574,N_17364,N_16414);
nor U19575 (N_19575,N_13869,N_15962);
or U19576 (N_19576,N_16819,N_13776);
or U19577 (N_19577,N_15646,N_16611);
nand U19578 (N_19578,N_14940,N_14219);
xor U19579 (N_19579,N_13675,N_15066);
xor U19580 (N_19580,N_12714,N_13306);
nand U19581 (N_19581,N_17874,N_17872);
or U19582 (N_19582,N_14183,N_17205);
nand U19583 (N_19583,N_14462,N_12124);
nand U19584 (N_19584,N_16706,N_17077);
or U19585 (N_19585,N_17976,N_16550);
or U19586 (N_19586,N_12588,N_14899);
nor U19587 (N_19587,N_16554,N_17070);
or U19588 (N_19588,N_16727,N_13110);
and U19589 (N_19589,N_13185,N_16561);
nand U19590 (N_19590,N_14818,N_12866);
nor U19591 (N_19591,N_13823,N_13337);
or U19592 (N_19592,N_12962,N_16786);
nor U19593 (N_19593,N_13328,N_12912);
nand U19594 (N_19594,N_14347,N_17646);
nor U19595 (N_19595,N_15717,N_13497);
xnor U19596 (N_19596,N_15665,N_16521);
nor U19597 (N_19597,N_15590,N_16670);
nor U19598 (N_19598,N_16297,N_13456);
nand U19599 (N_19599,N_17519,N_13085);
nor U19600 (N_19600,N_15704,N_14743);
xor U19601 (N_19601,N_16176,N_13452);
xor U19602 (N_19602,N_15184,N_12415);
or U19603 (N_19603,N_12807,N_14114);
nand U19604 (N_19604,N_17897,N_17027);
nor U19605 (N_19605,N_14824,N_12865);
nor U19606 (N_19606,N_17736,N_15952);
nor U19607 (N_19607,N_13558,N_16195);
and U19608 (N_19608,N_15199,N_17716);
nand U19609 (N_19609,N_12684,N_15382);
nand U19610 (N_19610,N_15559,N_17678);
or U19611 (N_19611,N_15125,N_16192);
or U19612 (N_19612,N_12394,N_16225);
or U19613 (N_19613,N_16588,N_15869);
or U19614 (N_19614,N_12618,N_12298);
and U19615 (N_19615,N_15644,N_13849);
nor U19616 (N_19616,N_12772,N_17749);
nand U19617 (N_19617,N_17679,N_12859);
and U19618 (N_19618,N_15322,N_13562);
nor U19619 (N_19619,N_12713,N_15251);
nand U19620 (N_19620,N_14411,N_16607);
or U19621 (N_19621,N_14634,N_13058);
and U19622 (N_19622,N_16067,N_12344);
nor U19623 (N_19623,N_16054,N_16700);
and U19624 (N_19624,N_13321,N_14079);
nand U19625 (N_19625,N_16252,N_13953);
or U19626 (N_19626,N_14231,N_14041);
and U19627 (N_19627,N_13500,N_14786);
or U19628 (N_19628,N_13004,N_15228);
or U19629 (N_19629,N_15723,N_12993);
and U19630 (N_19630,N_17668,N_17445);
nor U19631 (N_19631,N_12510,N_15243);
nor U19632 (N_19632,N_17241,N_17961);
nor U19633 (N_19633,N_15371,N_14213);
and U19634 (N_19634,N_14206,N_17614);
or U19635 (N_19635,N_16477,N_12085);
nor U19636 (N_19636,N_16353,N_12194);
and U19637 (N_19637,N_12812,N_13837);
or U19638 (N_19638,N_16393,N_13350);
xor U19639 (N_19639,N_17383,N_17900);
nand U19640 (N_19640,N_14440,N_17004);
nor U19641 (N_19641,N_15883,N_15019);
nand U19642 (N_19642,N_14568,N_15584);
nand U19643 (N_19643,N_15263,N_13835);
and U19644 (N_19644,N_15812,N_16620);
and U19645 (N_19645,N_16185,N_16822);
nor U19646 (N_19646,N_14188,N_15999);
and U19647 (N_19647,N_15583,N_14610);
xor U19648 (N_19648,N_14143,N_17380);
and U19649 (N_19649,N_13586,N_17645);
nand U19650 (N_19650,N_14430,N_14494);
or U19651 (N_19651,N_13044,N_12568);
and U19652 (N_19652,N_16017,N_13448);
nand U19653 (N_19653,N_15738,N_14166);
or U19654 (N_19654,N_14516,N_14619);
and U19655 (N_19655,N_15871,N_15245);
xnor U19656 (N_19656,N_15078,N_16795);
or U19657 (N_19657,N_13920,N_17686);
xor U19658 (N_19658,N_13120,N_15757);
and U19659 (N_19659,N_15633,N_14442);
nand U19660 (N_19660,N_15933,N_16748);
xor U19661 (N_19661,N_14741,N_16654);
and U19662 (N_19662,N_14762,N_14812);
xnor U19663 (N_19663,N_16798,N_16173);
or U19664 (N_19664,N_14433,N_16693);
and U19665 (N_19665,N_16418,N_17932);
and U19666 (N_19666,N_14774,N_14736);
and U19667 (N_19667,N_12203,N_17773);
or U19668 (N_19668,N_13196,N_15273);
nand U19669 (N_19669,N_17471,N_17188);
or U19670 (N_19670,N_13987,N_12166);
and U19671 (N_19671,N_12010,N_12316);
and U19672 (N_19672,N_16616,N_15142);
nand U19673 (N_19673,N_12057,N_12100);
and U19674 (N_19674,N_15725,N_13098);
xnor U19675 (N_19675,N_17258,N_16200);
xor U19676 (N_19676,N_12175,N_17122);
nor U19677 (N_19677,N_14278,N_16984);
nand U19678 (N_19678,N_12780,N_15155);
nand U19679 (N_19679,N_13535,N_13123);
nor U19680 (N_19680,N_17207,N_17901);
nor U19681 (N_19681,N_16520,N_16651);
xnor U19682 (N_19682,N_13416,N_15195);
xor U19683 (N_19683,N_16626,N_16253);
nor U19684 (N_19684,N_14982,N_14343);
nor U19685 (N_19685,N_12318,N_14970);
or U19686 (N_19686,N_13916,N_16747);
or U19687 (N_19687,N_12239,N_13385);
or U19688 (N_19688,N_14189,N_17125);
and U19689 (N_19689,N_12042,N_15099);
nand U19690 (N_19690,N_12378,N_17525);
and U19691 (N_19691,N_15230,N_17146);
xnor U19692 (N_19692,N_13740,N_17532);
nand U19693 (N_19693,N_15057,N_14928);
and U19694 (N_19694,N_12707,N_15853);
xor U19695 (N_19695,N_17999,N_17956);
xor U19696 (N_19696,N_14873,N_15072);
nand U19697 (N_19697,N_15885,N_12280);
or U19698 (N_19698,N_12821,N_17068);
xor U19699 (N_19699,N_15010,N_15310);
xor U19700 (N_19700,N_16979,N_17755);
or U19701 (N_19701,N_17022,N_17760);
or U19702 (N_19702,N_17008,N_14394);
or U19703 (N_19703,N_16299,N_14707);
nor U19704 (N_19704,N_12459,N_16894);
or U19705 (N_19705,N_16636,N_14476);
nand U19706 (N_19706,N_15807,N_13042);
or U19707 (N_19707,N_16875,N_12983);
nand U19708 (N_19708,N_16152,N_13521);
nand U19709 (N_19709,N_15977,N_15926);
nor U19710 (N_19710,N_17259,N_13939);
or U19711 (N_19711,N_12119,N_17237);
nor U19712 (N_19712,N_15422,N_13704);
nor U19713 (N_19713,N_12674,N_14943);
nand U19714 (N_19714,N_13750,N_16545);
or U19715 (N_19715,N_16404,N_13984);
xor U19716 (N_19716,N_13903,N_12233);
xnor U19717 (N_19717,N_12043,N_12140);
nor U19718 (N_19718,N_12296,N_12511);
nand U19719 (N_19719,N_15693,N_17114);
nor U19720 (N_19720,N_13839,N_16305);
xor U19721 (N_19721,N_14944,N_13160);
nand U19722 (N_19722,N_13868,N_17284);
nand U19723 (N_19723,N_13902,N_14583);
nor U19724 (N_19724,N_16071,N_14174);
nand U19725 (N_19725,N_17126,N_15810);
nand U19726 (N_19726,N_16909,N_17689);
or U19727 (N_19727,N_14661,N_12157);
nor U19728 (N_19728,N_14270,N_14077);
or U19729 (N_19729,N_16527,N_17266);
nor U19730 (N_19730,N_12405,N_17568);
xor U19731 (N_19731,N_15790,N_17622);
and U19732 (N_19732,N_13426,N_13891);
and U19733 (N_19733,N_13994,N_14606);
nand U19734 (N_19734,N_12453,N_14952);
xor U19735 (N_19735,N_17313,N_17501);
or U19736 (N_19736,N_16797,N_12589);
nand U19737 (N_19737,N_14075,N_15982);
and U19738 (N_19738,N_14009,N_13962);
and U19739 (N_19739,N_15298,N_15025);
or U19740 (N_19740,N_13655,N_15050);
or U19741 (N_19741,N_12960,N_15842);
nor U19742 (N_19742,N_15448,N_15182);
xnor U19743 (N_19743,N_17858,N_14862);
nand U19744 (N_19744,N_12797,N_14655);
nand U19745 (N_19745,N_16399,N_17762);
nand U19746 (N_19746,N_16188,N_17104);
or U19747 (N_19747,N_13857,N_12148);
xnor U19748 (N_19748,N_15365,N_16318);
nand U19749 (N_19749,N_17323,N_13400);
or U19750 (N_19750,N_12595,N_14708);
and U19751 (N_19751,N_14117,N_14099);
and U19752 (N_19752,N_16428,N_17602);
nand U19753 (N_19753,N_16075,N_17559);
nand U19754 (N_19754,N_12268,N_12049);
or U19755 (N_19755,N_13281,N_12205);
nor U19756 (N_19756,N_13067,N_15876);
xor U19757 (N_19757,N_15949,N_15968);
nor U19758 (N_19758,N_14340,N_17487);
and U19759 (N_19759,N_16745,N_12689);
and U19760 (N_19760,N_16451,N_13133);
nand U19761 (N_19761,N_16234,N_16063);
nand U19762 (N_19762,N_16002,N_13034);
xnor U19763 (N_19763,N_16578,N_15978);
nor U19764 (N_19764,N_12789,N_15139);
nor U19765 (N_19765,N_14994,N_14115);
xnor U19766 (N_19766,N_17273,N_15029);
and U19767 (N_19767,N_12304,N_13008);
and U19768 (N_19768,N_17865,N_16640);
and U19769 (N_19769,N_12650,N_16919);
or U19770 (N_19770,N_17918,N_15838);
or U19771 (N_19771,N_17859,N_14828);
nor U19772 (N_19772,N_13449,N_17928);
or U19773 (N_19773,N_13187,N_13344);
or U19774 (N_19774,N_12081,N_14509);
or U19775 (N_19775,N_13380,N_16998);
or U19776 (N_19776,N_12853,N_16686);
nand U19777 (N_19777,N_17662,N_13568);
and U19778 (N_19778,N_12435,N_15996);
or U19779 (N_19779,N_15077,N_16406);
nor U19780 (N_19780,N_15102,N_12044);
xor U19781 (N_19781,N_13770,N_13533);
xnor U19782 (N_19782,N_16207,N_12317);
xnor U19783 (N_19783,N_15946,N_16366);
and U19784 (N_19784,N_15791,N_17806);
nor U19785 (N_19785,N_16784,N_15373);
xnor U19786 (N_19786,N_13134,N_14159);
nand U19787 (N_19787,N_12902,N_14647);
nand U19788 (N_19788,N_13926,N_15940);
nor U19789 (N_19789,N_17342,N_15970);
and U19790 (N_19790,N_15492,N_14626);
nor U19791 (N_19791,N_12576,N_14271);
and U19792 (N_19792,N_17627,N_17665);
xor U19793 (N_19793,N_15368,N_13724);
xnor U19794 (N_19794,N_17817,N_14573);
nand U19795 (N_19795,N_15569,N_15197);
or U19796 (N_19796,N_14103,N_15566);
nor U19797 (N_19797,N_14058,N_17732);
nor U19798 (N_19798,N_12831,N_13254);
or U19799 (N_19799,N_12005,N_14048);
nor U19800 (N_19800,N_15662,N_15270);
nor U19801 (N_19801,N_15424,N_12655);
and U19802 (N_19802,N_13877,N_12392);
or U19803 (N_19803,N_14689,N_15160);
and U19804 (N_19804,N_16579,N_17793);
nand U19805 (N_19805,N_17177,N_12067);
or U19806 (N_19806,N_13367,N_17754);
nor U19807 (N_19807,N_17837,N_13432);
nand U19808 (N_19808,N_17453,N_13441);
or U19809 (N_19809,N_17997,N_14281);
nand U19810 (N_19810,N_15284,N_13005);
xnor U19811 (N_19811,N_13560,N_15964);
or U19812 (N_19812,N_15279,N_16030);
xnor U19813 (N_19813,N_16475,N_17674);
xor U19814 (N_19814,N_12406,N_14291);
xnor U19815 (N_19815,N_13317,N_17513);
nand U19816 (N_19816,N_17641,N_15770);
or U19817 (N_19817,N_13713,N_16707);
nand U19818 (N_19818,N_13954,N_13881);
xor U19819 (N_19819,N_14835,N_13235);
nand U19820 (N_19820,N_14020,N_14810);
nand U19821 (N_19821,N_15995,N_17397);
and U19822 (N_19822,N_12335,N_13153);
or U19823 (N_19823,N_13364,N_12644);
nor U19824 (N_19824,N_17043,N_14716);
nor U19825 (N_19825,N_12328,N_14420);
nand U19826 (N_19826,N_12709,N_15987);
or U19827 (N_19827,N_16841,N_13055);
and U19828 (N_19828,N_14357,N_17477);
or U19829 (N_19829,N_13982,N_12830);
xor U19830 (N_19830,N_13345,N_14369);
xor U19831 (N_19831,N_13861,N_15137);
xor U19832 (N_19832,N_17890,N_15367);
or U19833 (N_19833,N_12040,N_17550);
or U19834 (N_19834,N_12290,N_17737);
and U19835 (N_19835,N_17847,N_15754);
and U19836 (N_19836,N_16025,N_12843);
nand U19837 (N_19837,N_12199,N_15038);
nand U19838 (N_19838,N_13739,N_15286);
nor U19839 (N_19839,N_17822,N_17801);
or U19840 (N_19840,N_13211,N_13800);
nor U19841 (N_19841,N_12009,N_14827);
and U19842 (N_19842,N_15439,N_17371);
or U19843 (N_19843,N_16816,N_15806);
xnor U19844 (N_19844,N_14646,N_14960);
nor U19845 (N_19845,N_16667,N_13515);
or U19846 (N_19846,N_16311,N_16421);
nand U19847 (N_19847,N_17578,N_17456);
nor U19848 (N_19848,N_15534,N_15183);
xor U19849 (N_19849,N_12664,N_16915);
or U19850 (N_19850,N_15748,N_16854);
nor U19851 (N_19851,N_12922,N_16074);
and U19852 (N_19852,N_12083,N_13002);
and U19853 (N_19853,N_17624,N_13286);
nor U19854 (N_19854,N_13596,N_14026);
or U19855 (N_19855,N_15352,N_16239);
nand U19856 (N_19856,N_15045,N_17014);
or U19857 (N_19857,N_12121,N_12376);
or U19858 (N_19858,N_17649,N_16443);
nor U19859 (N_19859,N_12967,N_17951);
nand U19860 (N_19860,N_13822,N_13503);
xor U19861 (N_19861,N_15551,N_14800);
nand U19862 (N_19862,N_14577,N_14470);
xnor U19863 (N_19863,N_16801,N_12688);
or U19864 (N_19864,N_17960,N_13458);
nand U19865 (N_19865,N_15815,N_13735);
xnor U19866 (N_19866,N_17239,N_14596);
or U19867 (N_19867,N_12911,N_14588);
or U19868 (N_19868,N_14190,N_12710);
or U19869 (N_19869,N_14038,N_17860);
nor U19870 (N_19870,N_17112,N_16850);
or U19871 (N_19871,N_13977,N_12893);
nor U19872 (N_19872,N_15116,N_15318);
nand U19873 (N_19873,N_14875,N_13838);
and U19874 (N_19874,N_17981,N_12412);
xor U19875 (N_19875,N_15719,N_14454);
nand U19876 (N_19876,N_14373,N_17097);
and U19877 (N_19877,N_13279,N_14076);
and U19878 (N_19878,N_15822,N_14450);
nand U19879 (N_19879,N_12547,N_16794);
and U19880 (N_19880,N_14445,N_15588);
and U19881 (N_19881,N_14578,N_15740);
nand U19882 (N_19882,N_16350,N_16907);
nor U19883 (N_19883,N_12234,N_13214);
nor U19884 (N_19884,N_14916,N_17820);
xor U19885 (N_19885,N_12432,N_16324);
and U19886 (N_19886,N_12783,N_15539);
nor U19887 (N_19887,N_12522,N_14418);
xor U19888 (N_19888,N_12073,N_15312);
and U19889 (N_19889,N_16926,N_14894);
nand U19890 (N_19890,N_12899,N_15453);
and U19891 (N_19891,N_16835,N_16646);
nor U19892 (N_19892,N_14597,N_15269);
xnor U19893 (N_19893,N_14247,N_12943);
nor U19894 (N_19894,N_12135,N_15694);
and U19895 (N_19895,N_14249,N_12307);
nand U19896 (N_19896,N_13812,N_12606);
nand U19897 (N_19897,N_13935,N_12538);
nor U19898 (N_19898,N_16272,N_14653);
xnor U19899 (N_19899,N_15117,N_17165);
xor U19900 (N_19900,N_17658,N_13763);
xor U19901 (N_19901,N_16828,N_17950);
nand U19902 (N_19902,N_16449,N_14660);
nand U19903 (N_19903,N_15330,N_15014);
or U19904 (N_19904,N_13651,N_12122);
and U19905 (N_19905,N_17201,N_12776);
and U19906 (N_19906,N_16241,N_15157);
xor U19907 (N_19907,N_14534,N_13313);
nand U19908 (N_19908,N_15039,N_12425);
or U19909 (N_19909,N_15106,N_17844);
xnor U19910 (N_19910,N_17072,N_17291);
or U19911 (N_19911,N_16761,N_14554);
nor U19912 (N_19912,N_14986,N_14263);
nor U19913 (N_19913,N_16265,N_12968);
or U19914 (N_19914,N_17096,N_15858);
or U19915 (N_19915,N_15489,N_16785);
xnor U19916 (N_19916,N_16722,N_15525);
nor U19917 (N_19917,N_15143,N_13451);
nand U19918 (N_19918,N_13129,N_15896);
nor U19919 (N_19919,N_13467,N_15581);
xnor U19920 (N_19920,N_15293,N_12851);
nor U19921 (N_19921,N_14230,N_16757);
nand U19922 (N_19922,N_12749,N_12259);
or U19923 (N_19923,N_13361,N_14787);
or U19924 (N_19924,N_13965,N_16731);
and U19925 (N_19925,N_16059,N_12450);
and U19926 (N_19926,N_14006,N_17400);
xnor U19927 (N_19927,N_15683,N_13288);
nand U19928 (N_19928,N_14413,N_13264);
xnor U19929 (N_19929,N_12013,N_16330);
or U19930 (N_19930,N_15383,N_13347);
xnor U19931 (N_19931,N_13010,N_16023);
or U19932 (N_19932,N_17784,N_13580);
nor U19933 (N_19933,N_14108,N_12930);
and U19934 (N_19934,N_17232,N_13111);
or U19935 (N_19935,N_15734,N_14367);
nand U19936 (N_19936,N_16065,N_15340);
or U19937 (N_19937,N_16113,N_16564);
nand U19938 (N_19938,N_13911,N_17768);
and U19939 (N_19939,N_13627,N_12765);
nor U19940 (N_19940,N_12828,N_17786);
nor U19941 (N_19941,N_17238,N_13624);
nand U19942 (N_19942,N_16990,N_14342);
nand U19943 (N_19943,N_14909,N_13730);
nor U19944 (N_19944,N_13457,N_15124);
xor U19945 (N_19945,N_17159,N_14389);
or U19946 (N_19946,N_14229,N_12641);
nand U19947 (N_19947,N_12507,N_16687);
xor U19948 (N_19948,N_14368,N_16612);
nor U19949 (N_19949,N_16049,N_13879);
xor U19950 (N_19950,N_13144,N_15894);
and U19951 (N_19951,N_16178,N_12665);
xor U19952 (N_19952,N_12920,N_13405);
xor U19953 (N_19953,N_13180,N_16593);
nor U19954 (N_19954,N_12768,N_17228);
nand U19955 (N_19955,N_15265,N_17856);
and U19956 (N_19956,N_12697,N_15416);
nand U19957 (N_19957,N_15362,N_13649);
nor U19958 (N_19958,N_16831,N_14883);
or U19959 (N_19959,N_15154,N_13340);
nand U19960 (N_19960,N_17479,N_12131);
xor U19961 (N_19961,N_17968,N_16713);
nor U19962 (N_19962,N_16838,N_17756);
xor U19963 (N_19963,N_13577,N_12945);
nor U19964 (N_19964,N_16468,N_16445);
xor U19965 (N_19965,N_13747,N_13115);
and U19966 (N_19966,N_17938,N_13381);
xnor U19967 (N_19967,N_14266,N_13151);
nand U19968 (N_19968,N_13556,N_15736);
nor U19969 (N_19969,N_17093,N_13767);
nand U19970 (N_19970,N_17790,N_15845);
nand U19971 (N_19971,N_13181,N_12273);
nand U19972 (N_19972,N_12903,N_15541);
nand U19973 (N_19973,N_17088,N_14086);
xnor U19974 (N_19974,N_12179,N_13663);
xnor U19975 (N_19975,N_17425,N_12746);
nand U19976 (N_19976,N_14280,N_16480);
or U19977 (N_19977,N_16077,N_12197);
and U19978 (N_19978,N_16910,N_14891);
nand U19979 (N_19979,N_16045,N_16681);
xnor U19980 (N_19980,N_13705,N_14139);
nor U19981 (N_19981,N_15532,N_15781);
xnor U19982 (N_19982,N_14556,N_17288);
xor U19983 (N_19983,N_14759,N_12169);
nand U19984 (N_19984,N_16760,N_17139);
and U19985 (N_19985,N_16014,N_14274);
or U19986 (N_19986,N_13865,N_13498);
and U19987 (N_19987,N_15993,N_13319);
or U19988 (N_19988,N_16053,N_14463);
xnor U19989 (N_19989,N_16940,N_12369);
and U19990 (N_19990,N_13444,N_13492);
nand U19991 (N_19991,N_17119,N_13234);
nor U19992 (N_19992,N_14370,N_12790);
nand U19993 (N_19993,N_16643,N_16187);
or U19994 (N_19994,N_14119,N_15360);
nand U19995 (N_19995,N_12278,N_14438);
nor U19996 (N_19996,N_12941,N_16934);
nor U19997 (N_19997,N_15768,N_12520);
nor U19998 (N_19998,N_13305,N_12142);
xnor U19999 (N_19999,N_14074,N_12570);
nor U20000 (N_20000,N_17830,N_14310);
or U20001 (N_20001,N_17051,N_16641);
xor U20002 (N_20002,N_14726,N_16833);
and U20003 (N_20003,N_13357,N_13146);
nand U20004 (N_20004,N_16892,N_16989);
nor U20005 (N_20005,N_12351,N_13506);
or U20006 (N_20006,N_14915,N_15889);
nor U20007 (N_20007,N_15086,N_12153);
nand U20008 (N_20008,N_17523,N_14146);
xor U20009 (N_20009,N_16472,N_15715);
nand U20010 (N_20010,N_17791,N_12382);
xor U20011 (N_20011,N_12926,N_15973);
and U20012 (N_20012,N_14156,N_16118);
nor U20013 (N_20013,N_15297,N_14644);
nor U20014 (N_20014,N_16000,N_12577);
nand U20015 (N_20015,N_14695,N_15358);
nand U20016 (N_20016,N_15395,N_14313);
nand U20017 (N_20017,N_12867,N_13543);
and U20018 (N_20018,N_13529,N_13420);
nor U20019 (N_20019,N_12103,N_17935);
xnor U20020 (N_20020,N_15857,N_17468);
nand U20021 (N_20021,N_15504,N_16070);
or U20022 (N_20022,N_13536,N_17507);
or U20023 (N_20023,N_17992,N_16997);
and U20024 (N_20024,N_14215,N_17123);
and U20025 (N_20025,N_15923,N_14752);
xor U20026 (N_20026,N_16256,N_14195);
nand U20027 (N_20027,N_17895,N_15193);
or U20028 (N_20028,N_15870,N_14200);
xor U20029 (N_20029,N_13390,N_13820);
nand U20030 (N_20030,N_13017,N_13208);
nand U20031 (N_20031,N_12295,N_12582);
and U20032 (N_20032,N_17083,N_12445);
and U20033 (N_20033,N_12276,N_16221);
xor U20034 (N_20034,N_17174,N_14767);
nor U20035 (N_20035,N_14846,N_17499);
nand U20036 (N_20036,N_15491,N_13125);
and U20037 (N_20037,N_16750,N_15848);
or U20038 (N_20038,N_16775,N_15370);
nor U20039 (N_20039,N_14908,N_14856);
or U20040 (N_20040,N_12054,N_16386);
and U20041 (N_20041,N_14032,N_12787);
xnor U20042 (N_20042,N_14257,N_12671);
or U20043 (N_20043,N_14224,N_17920);
xnor U20044 (N_20044,N_17382,N_14105);
xor U20045 (N_20045,N_17922,N_12627);
xnor U20046 (N_20046,N_17699,N_13119);
xor U20047 (N_20047,N_15553,N_17478);
and U20048 (N_20048,N_14772,N_15997);
or U20049 (N_20049,N_13789,N_17461);
and U20050 (N_20050,N_13352,N_13343);
xor U20051 (N_20051,N_16871,N_13561);
nand U20052 (N_20052,N_17357,N_15528);
nand U20053 (N_20053,N_14023,N_14897);
or U20054 (N_20054,N_15930,N_15597);
and U20055 (N_20055,N_13327,N_16347);
xor U20056 (N_20056,N_17424,N_14227);
xor U20057 (N_20057,N_14570,N_16117);
xor U20058 (N_20058,N_16435,N_15339);
and U20059 (N_20059,N_14823,N_17484);
nand U20060 (N_20060,N_13637,N_13985);
and U20061 (N_20061,N_14640,N_14170);
nor U20062 (N_20062,N_13289,N_14013);
and U20063 (N_20063,N_13126,N_14920);
or U20064 (N_20064,N_16344,N_16487);
or U20065 (N_20065,N_15877,N_13991);
nand U20066 (N_20066,N_16590,N_15576);
nand U20067 (N_20067,N_13512,N_13919);
or U20068 (N_20068,N_13998,N_13853);
nand U20069 (N_20069,N_14515,N_13760);
nor U20070 (N_20070,N_14848,N_16334);
or U20071 (N_20071,N_14720,N_15976);
nand U20072 (N_20072,N_17855,N_13643);
nand U20073 (N_20073,N_16044,N_17255);
xnor U20074 (N_20074,N_14208,N_14018);
nor U20075 (N_20075,N_13207,N_15181);
nand U20076 (N_20076,N_12118,N_12452);
or U20077 (N_20077,N_13140,N_16142);
nor U20078 (N_20078,N_13417,N_16286);
and U20079 (N_20079,N_14951,N_12409);
nand U20080 (N_20080,N_15670,N_17047);
nand U20081 (N_20081,N_14618,N_12708);
xnor U20082 (N_20082,N_14315,N_15051);
nand U20083 (N_20083,N_16534,N_12050);
or U20084 (N_20084,N_13656,N_13480);
and U20085 (N_20085,N_15483,N_15519);
nand U20086 (N_20086,N_14001,N_12497);
xnor U20087 (N_20087,N_12464,N_16676);
xnor U20088 (N_20088,N_17401,N_15427);
or U20089 (N_20089,N_14022,N_13721);
or U20090 (N_20090,N_13511,N_17337);
xor U20091 (N_20091,N_17287,N_16028);
nand U20092 (N_20092,N_17948,N_15433);
xor U20093 (N_20093,N_15907,N_17422);
xor U20094 (N_20094,N_17882,N_16530);
xor U20095 (N_20095,N_15953,N_12722);
and U20096 (N_20096,N_12250,N_16988);
and U20097 (N_20097,N_14379,N_13687);
or U20098 (N_20098,N_12935,N_12074);
nand U20099 (N_20099,N_14754,N_14232);
xnor U20100 (N_20100,N_16367,N_16976);
nor U20101 (N_20101,N_15046,N_12766);
or U20102 (N_20102,N_12158,N_12027);
nand U20103 (N_20103,N_16090,N_14386);
or U20104 (N_20104,N_14094,N_12003);
and U20105 (N_20105,N_13976,N_12702);
xnor U20106 (N_20106,N_16018,N_14765);
and U20107 (N_20107,N_16465,N_13635);
and U20108 (N_20108,N_13897,N_16327);
or U20109 (N_20109,N_16591,N_17548);
nand U20110 (N_20110,N_17617,N_15998);
xnor U20111 (N_20111,N_12619,N_17536);
or U20112 (N_20112,N_13102,N_13833);
xnor U20113 (N_20113,N_17312,N_15988);
or U20114 (N_20114,N_17643,N_14298);
or U20115 (N_20115,N_16522,N_16111);
nor U20116 (N_20116,N_15028,N_13411);
nand U20117 (N_20117,N_13810,N_12906);
nand U20118 (N_20118,N_13013,N_14435);
or U20119 (N_20119,N_17494,N_15032);
nand U20120 (N_20120,N_17719,N_12652);
nor U20121 (N_20121,N_16057,N_15844);
or U20122 (N_20122,N_15134,N_17169);
nand U20123 (N_20123,N_12742,N_13078);
or U20124 (N_20124,N_17144,N_14087);
nand U20125 (N_20125,N_12061,N_13228);
xor U20126 (N_20126,N_12417,N_13412);
xor U20127 (N_20127,N_16573,N_14620);
nor U20128 (N_20128,N_17319,N_14165);
xor U20129 (N_20129,N_13198,N_13664);
nand U20130 (N_20130,N_12546,N_14805);
nor U20131 (N_20131,N_16136,N_16703);
and U20132 (N_20132,N_14536,N_17419);
and U20133 (N_20133,N_14804,N_15126);
and U20134 (N_20134,N_14346,N_14794);
xor U20135 (N_20135,N_15943,N_16736);
and U20136 (N_20136,N_15636,N_17061);
nand U20137 (N_20137,N_16068,N_16151);
nand U20138 (N_20138,N_17310,N_15434);
nor U20139 (N_20139,N_17173,N_16862);
nor U20140 (N_20140,N_15634,N_13066);
and U20141 (N_20141,N_12630,N_14849);
or U20142 (N_20142,N_16507,N_17937);
or U20143 (N_20143,N_12088,N_14822);
and U20144 (N_20144,N_15598,N_16260);
nand U20145 (N_20145,N_15202,N_14681);
and U20146 (N_20146,N_13904,N_16580);
xnor U20147 (N_20147,N_15697,N_17067);
nand U20148 (N_20148,N_14766,N_15443);
and U20149 (N_20149,N_12762,N_15990);
nand U20150 (N_20150,N_14484,N_15488);
xnor U20151 (N_20151,N_12838,N_15664);
and U20152 (N_20152,N_16627,N_15469);
and U20153 (N_20153,N_15233,N_12861);
or U20154 (N_20154,N_17601,N_15542);
xnor U20155 (N_20155,N_14372,N_14192);
and U20156 (N_20156,N_14962,N_16281);
nand U20157 (N_20157,N_13933,N_14081);
nor U20158 (N_20158,N_13836,N_17271);
or U20159 (N_20159,N_13213,N_15421);
nor U20160 (N_20160,N_13382,N_14776);
and U20161 (N_20161,N_17187,N_17091);
nand U20162 (N_20162,N_12654,N_17670);
xor U20163 (N_20163,N_17738,N_13052);
xor U20164 (N_20164,N_17506,N_15201);
nand U20165 (N_20165,N_14154,N_14137);
and U20166 (N_20166,N_17727,N_16675);
or U20167 (N_20167,N_12442,N_14684);
or U20168 (N_20168,N_14890,N_13690);
nor U20169 (N_20169,N_13223,N_13616);
nor U20170 (N_20170,N_17224,N_16325);
xnor U20171 (N_20171,N_17387,N_17251);
nand U20172 (N_20172,N_12515,N_13749);
xnor U20173 (N_20173,N_14809,N_12099);
nor U20174 (N_20174,N_14733,N_13574);
nor U20175 (N_20175,N_14448,N_14107);
nor U20176 (N_20176,N_17275,N_17971);
nor U20177 (N_20177,N_13043,N_14718);
and U20178 (N_20178,N_16566,N_15083);
and U20179 (N_20179,N_17842,N_14253);
xnor U20180 (N_20180,N_16179,N_14679);
xnor U20181 (N_20181,N_16993,N_13152);
nor U20182 (N_20182,N_12875,N_15447);
xnor U20183 (N_20183,N_14842,N_14632);
xnor U20184 (N_20184,N_15765,N_16328);
and U20185 (N_20185,N_15841,N_15942);
xnor U20186 (N_20186,N_15592,N_14796);
xnor U20187 (N_20187,N_15456,N_13294);
nor U20188 (N_20188,N_13625,N_14789);
or U20189 (N_20189,N_14924,N_17396);
xor U20190 (N_20190,N_12075,N_14366);
xor U20191 (N_20191,N_17131,N_17772);
or U20192 (N_20192,N_14927,N_15177);
or U20193 (N_20193,N_14182,N_13975);
and U20194 (N_20194,N_17363,N_14323);
and U20195 (N_20195,N_16512,N_13677);
or U20196 (N_20196,N_17659,N_15616);
nor U20197 (N_20197,N_13334,N_17979);
and U20198 (N_20198,N_16860,N_14475);
xnor U20199 (N_20199,N_16351,N_15071);
or U20200 (N_20200,N_13658,N_13230);
nor U20201 (N_20201,N_17378,N_17515);
and U20202 (N_20202,N_14175,N_13027);
or U20203 (N_20203,N_17019,N_12579);
nand U20204 (N_20204,N_13516,N_15645);
or U20205 (N_20205,N_16425,N_13114);
xnor U20206 (N_20206,N_12306,N_12084);
nand U20207 (N_20207,N_14844,N_17591);
xor U20208 (N_20208,N_16684,N_15156);
and U20209 (N_20209,N_14453,N_14637);
and U20210 (N_20210,N_16267,N_13354);
nand U20211 (N_20211,N_13938,N_16106);
and U20212 (N_20212,N_15430,N_17924);
nor U20213 (N_20213,N_13898,N_13746);
nor U20214 (N_20214,N_12844,N_16016);
nand U20215 (N_20215,N_15043,N_17293);
or U20216 (N_20216,N_13326,N_17094);
nand U20217 (N_20217,N_15506,N_16711);
nand U20218 (N_20218,N_12977,N_14065);
nand U20219 (N_20219,N_17783,N_12028);
nor U20220 (N_20220,N_15314,N_14525);
nand U20221 (N_20221,N_14514,N_13250);
or U20222 (N_20222,N_16508,N_14235);
nand U20223 (N_20223,N_15100,N_12039);
xor U20224 (N_20224,N_12138,N_13050);
nand U20225 (N_20225,N_13244,N_15708);
nor U20226 (N_20226,N_17700,N_12171);
or U20227 (N_20227,N_14884,N_12440);
or U20228 (N_20228,N_13575,N_12438);
nand U20229 (N_20229,N_15260,N_12657);
nor U20230 (N_20230,N_14705,N_13475);
nor U20231 (N_20231,N_16596,N_13338);
or U20232 (N_20232,N_12000,N_14358);
or U20233 (N_20233,N_14980,N_15307);
nor U20234 (N_20234,N_15267,N_14769);
or U20235 (N_20235,N_16638,N_13301);
or U20236 (N_20236,N_13854,N_12110);
or U20237 (N_20237,N_12116,N_17908);
nand U20238 (N_20238,N_17606,N_15776);
xor U20239 (N_20239,N_16728,N_16729);
xor U20240 (N_20240,N_14129,N_13668);
nand U20241 (N_20241,N_17303,N_15272);
and U20242 (N_20242,N_16144,N_17826);
xor U20243 (N_20243,N_16120,N_14829);
xnor U20244 (N_20244,N_15449,N_16986);
or U20245 (N_20245,N_16872,N_12716);
and U20246 (N_20246,N_13026,N_15311);
or U20247 (N_20247,N_17739,N_16518);
nor U20248 (N_20248,N_17666,N_13524);
and U20249 (N_20249,N_12888,N_16743);
nor U20250 (N_20250,N_16715,N_17543);
nand U20251 (N_20251,N_16084,N_15651);
and U20252 (N_20252,N_16007,N_17370);
and U20253 (N_20253,N_14052,N_12421);
xor U20254 (N_20254,N_12363,N_14098);
nor U20255 (N_20255,N_14217,N_16066);
xor U20256 (N_20256,N_17086,N_13329);
xnor U20257 (N_20257,N_16619,N_14721);
xnor U20258 (N_20258,N_16980,N_13807);
and U20259 (N_20259,N_12365,N_15587);
or U20260 (N_20260,N_15762,N_14793);
nand U20261 (N_20261,N_16243,N_14869);
nand U20262 (N_20262,N_13942,N_15980);
and U20263 (N_20263,N_12553,N_13041);
and U20264 (N_20264,N_14854,N_13847);
nand U20265 (N_20265,N_13722,N_17983);
or U20266 (N_20266,N_15452,N_14709);
nand U20267 (N_20267,N_12572,N_13233);
and U20268 (N_20268,N_12686,N_16038);
and U20269 (N_20269,N_15451,N_14039);
nor U20270 (N_20270,N_13169,N_14176);
nor U20271 (N_20271,N_13973,N_17117);
nand U20272 (N_20272,N_17959,N_16051);
nand U20273 (N_20273,N_17751,N_12981);
or U20274 (N_20274,N_17850,N_13773);
or U20275 (N_20275,N_12600,N_13855);
nor U20276 (N_20276,N_16954,N_17899);
or U20277 (N_20277,N_16500,N_14091);
nand U20278 (N_20278,N_14101,N_17248);
or U20279 (N_20279,N_13604,N_14317);
and U20280 (N_20280,N_14914,N_16603);
xnor U20281 (N_20281,N_17327,N_13188);
or U20282 (N_20282,N_17893,N_16183);
xnor U20283 (N_20283,N_15364,N_12277);
or U20284 (N_20284,N_13583,N_17919);
or U20285 (N_20285,N_17527,N_16139);
nor U20286 (N_20286,N_15415,N_12455);
nor U20287 (N_20287,N_12635,N_16466);
nand U20288 (N_20288,N_13671,N_12615);
and U20289 (N_20289,N_13610,N_14710);
xnor U20290 (N_20290,N_12725,N_14832);
xnor U20291 (N_20291,N_17711,N_13678);
nand U20292 (N_20292,N_14356,N_13801);
and U20293 (N_20293,N_13589,N_17450);
nor U20294 (N_20294,N_13194,N_16594);
nor U20295 (N_20295,N_17455,N_15816);
nor U20296 (N_20296,N_16846,N_17510);
xnor U20297 (N_20297,N_13176,N_12539);
or U20298 (N_20298,N_14461,N_17413);
nand U20299 (N_20299,N_13312,N_14704);
or U20300 (N_20300,N_12449,N_16248);
or U20301 (N_20301,N_15152,N_15198);
nand U20302 (N_20302,N_17488,N_12660);
xnor U20303 (N_20303,N_13806,N_12254);
nand U20304 (N_20304,N_15785,N_13159);
and U20305 (N_20305,N_17612,N_15343);
xnor U20306 (N_20306,N_13788,N_12996);
nor U20307 (N_20307,N_17341,N_14168);
xor U20308 (N_20308,N_15249,N_15570);
nor U20309 (N_20309,N_12645,N_16069);
or U20310 (N_20310,N_14855,N_16905);
nor U20311 (N_20311,N_16719,N_15138);
xor U20312 (N_20312,N_16303,N_15934);
xnor U20313 (N_20313,N_14225,N_15327);
xnor U20314 (N_20314,N_13237,N_13921);
or U20315 (N_20315,N_14414,N_15713);
or U20316 (N_20316,N_16825,N_12087);
or U20317 (N_20317,N_17376,N_16034);
nor U20318 (N_20318,N_12236,N_14377);
xor U20319 (N_20319,N_16080,N_15860);
xnor U20320 (N_20320,N_14167,N_15037);
nor U20321 (N_20321,N_14612,N_16162);
nand U20322 (N_20322,N_15839,N_13741);
or U20323 (N_20323,N_13795,N_17652);
xor U20324 (N_20324,N_16679,N_12640);
nor U20325 (N_20325,N_17179,N_12496);
nor U20326 (N_20326,N_17809,N_15485);
and U20327 (N_20327,N_14616,N_12628);
nand U20328 (N_20328,N_14715,N_15054);
nand U20329 (N_20329,N_14228,N_15495);
or U20330 (N_20330,N_17823,N_12051);
xnor U20331 (N_20331,N_16012,N_15088);
nand U20332 (N_20332,N_12370,N_16859);
xor U20333 (N_20333,N_15460,N_17496);
nor U20334 (N_20334,N_13772,N_16820);
or U20335 (N_20335,N_14881,N_13331);
nor U20336 (N_20336,N_15767,N_16893);
xor U20337 (N_20337,N_17978,N_16093);
xor U20338 (N_20338,N_16901,N_14016);
or U20339 (N_20339,N_17116,N_15690);
nand U20340 (N_20340,N_16450,N_15161);
or U20341 (N_20341,N_17518,N_14999);
nand U20342 (N_20342,N_12802,N_14885);
and U20343 (N_20343,N_17121,N_15649);
nand U20344 (N_20344,N_17485,N_12585);
xnor U20345 (N_20345,N_16852,N_13302);
nor U20346 (N_20346,N_13141,N_16019);
nor U20347 (N_20347,N_15055,N_14746);
nand U20348 (N_20348,N_15954,N_14729);
and U20349 (N_20349,N_14649,N_13019);
and U20350 (N_20350,N_17604,N_17243);
and U20351 (N_20351,N_17618,N_17214);
nand U20352 (N_20352,N_16780,N_12091);
nand U20353 (N_20353,N_12025,N_16250);
nor U20354 (N_20354,N_17955,N_12592);
xor U20355 (N_20355,N_12143,N_12550);
and U20356 (N_20356,N_14339,N_17936);
nor U20357 (N_20357,N_17902,N_15820);
or U20358 (N_20358,N_13495,N_17194);
and U20359 (N_20359,N_15552,N_15002);
xnor U20360 (N_20360,N_15905,N_16515);
or U20361 (N_20361,N_16615,N_16536);
xnor U20362 (N_20362,N_17025,N_12111);
xnor U20363 (N_20363,N_12972,N_12281);
and U20364 (N_20364,N_12846,N_13053);
nor U20365 (N_20365,N_14258,N_12836);
xor U20366 (N_20366,N_12016,N_13970);
nor U20367 (N_20367,N_17292,N_17229);
nor U20368 (N_20368,N_12114,N_16010);
nand U20369 (N_20369,N_12964,N_17765);
nor U20370 (N_20370,N_17629,N_13291);
nor U20371 (N_20371,N_15023,N_14723);
xnor U20372 (N_20372,N_16878,N_14901);
xor U20373 (N_20373,N_17545,N_16378);
or U20374 (N_20374,N_15354,N_13890);
or U20375 (N_20375,N_15294,N_12729);
xnor U20376 (N_20376,N_13852,N_15846);
and U20377 (N_20377,N_16805,N_12266);
and U20378 (N_20378,N_12034,N_13167);
nor U20379 (N_20379,N_14497,N_13349);
xor U20380 (N_20380,N_15529,N_15843);
nor U20381 (N_20381,N_14668,N_15614);
nand U20382 (N_20382,N_13821,N_15499);
xor U20383 (N_20383,N_16403,N_13759);
and U20384 (N_20384,N_12429,N_12978);
or U20385 (N_20385,N_16413,N_16494);
xor U20386 (N_20386,N_13226,N_16682);
xnor U20387 (N_20387,N_17469,N_12398);
and U20388 (N_20388,N_13608,N_15795);
and U20389 (N_20389,N_13573,N_12474);
xor U20390 (N_20390,N_16129,N_12473);
nor U20391 (N_20391,N_17804,N_12948);
nand U20392 (N_20392,N_16371,N_14782);
nand U20393 (N_20393,N_13528,N_13074);
nand U20394 (N_20394,N_17318,N_15389);
xnor U20395 (N_20395,N_13488,N_17682);
xnor U20396 (N_20396,N_12026,N_15921);
or U20397 (N_20397,N_15215,N_15334);
or U20398 (N_20398,N_16232,N_17344);
xnor U20399 (N_20399,N_12574,N_17869);
nand U20400 (N_20400,N_15227,N_17728);
nand U20401 (N_20401,N_12679,N_17880);
nor U20402 (N_20402,N_12444,N_12521);
and U20403 (N_20403,N_15480,N_15455);
or U20404 (N_20404,N_12189,N_13547);
and U20405 (N_20405,N_12636,N_12739);
nor U20406 (N_20406,N_13928,N_14968);
nand U20407 (N_20407,N_15274,N_16865);
nor U20408 (N_20408,N_16388,N_12982);
or U20409 (N_20409,N_15799,N_17812);
nand U20410 (N_20410,N_16574,N_12045);
and U20411 (N_20411,N_16427,N_13841);
nand U20412 (N_20412,N_17000,N_15036);
and U20413 (N_20413,N_16504,N_12998);
nand U20414 (N_20414,N_13048,N_16575);
and U20415 (N_20415,N_15350,N_15832);
and U20416 (N_20416,N_13278,N_17730);
or U20417 (N_20417,N_13054,N_13439);
nand U20418 (N_20418,N_15324,N_14580);
xor U20419 (N_20419,N_15062,N_13395);
or U20420 (N_20420,N_14383,N_12030);
nand U20421 (N_20421,N_17409,N_15220);
xor U20422 (N_20422,N_15030,N_16205);
or U20423 (N_20423,N_12706,N_14727);
xor U20424 (N_20424,N_16380,N_17242);
nand U20425 (N_20425,N_13170,N_12908);
xor U20426 (N_20426,N_17569,N_13219);
and U20427 (N_20427,N_13258,N_17974);
or U20428 (N_20428,N_17474,N_16810);
and U20429 (N_20429,N_17164,N_13623);
nand U20430 (N_20430,N_17539,N_16132);
or U20431 (N_20431,N_12403,N_15619);
nand U20432 (N_20432,N_15208,N_16888);
and U20433 (N_20433,N_13983,N_17026);
nand U20434 (N_20434,N_14866,N_13095);
or U20435 (N_20435,N_16809,N_16204);
nand U20436 (N_20436,N_17777,N_13642);
and U20437 (N_20437,N_12478,N_14808);
or U20438 (N_20438,N_17200,N_17105);
or U20439 (N_20439,N_13654,N_12272);
xnor U20440 (N_20440,N_14902,N_15047);
and U20441 (N_20441,N_17407,N_14250);
and U20442 (N_20442,N_13149,N_12443);
nand U20443 (N_20443,N_12340,N_12436);
nor U20444 (N_20444,N_14801,N_15513);
xor U20445 (N_20445,N_12578,N_17998);
nand U20446 (N_20446,N_16553,N_16329);
and U20447 (N_20447,N_16079,N_16904);
or U20448 (N_20448,N_13725,N_13618);
nand U20449 (N_20449,N_12728,N_13447);
xnor U20450 (N_20450,N_13734,N_13362);
nor U20451 (N_20451,N_12258,N_17653);
and U20452 (N_20452,N_14150,N_15472);
and U20453 (N_20453,N_14912,N_13978);
and U20454 (N_20454,N_12183,N_13399);
and U20455 (N_20455,N_12256,N_13925);
xor U20456 (N_20456,N_17268,N_17189);
xnor U20457 (N_20457,N_12631,N_15425);
nor U20458 (N_20458,N_13414,N_12198);
nand U20459 (N_20459,N_12308,N_16600);
xnor U20460 (N_20460,N_15514,N_12820);
nand U20461 (N_20461,N_12536,N_16115);
xnor U20462 (N_20462,N_13737,N_17815);
nand U20463 (N_20463,N_15536,N_16917);
xor U20464 (N_20464,N_14264,N_13353);
and U20465 (N_20465,N_14871,N_12130);
and U20466 (N_20466,N_15782,N_15420);
nand U20467 (N_20467,N_13997,N_16356);
nand U20468 (N_20468,N_12833,N_14005);
or U20469 (N_20469,N_15642,N_13040);
and U20470 (N_20470,N_13924,N_12374);
and U20471 (N_20471,N_13224,N_14061);
or U20472 (N_20472,N_14080,N_12601);
nor U20473 (N_20473,N_16240,N_16617);
nor U20474 (N_20474,N_14402,N_12723);
or U20475 (N_20475,N_17721,N_15096);
and U20476 (N_20476,N_13221,N_15687);
nand U20477 (N_20477,N_14682,N_17006);
nand U20478 (N_20478,N_14062,N_13771);
xor U20479 (N_20479,N_12324,N_16994);
nand U20480 (N_20480,N_17964,N_13465);
xor U20481 (N_20481,N_16832,N_14498);
nand U20482 (N_20482,N_16790,N_17734);
nand U20483 (N_20483,N_14302,N_16839);
and U20484 (N_20484,N_16924,N_17442);
and U20485 (N_20485,N_12770,N_15256);
and U20486 (N_20486,N_15401,N_14607);
xnor U20487 (N_20487,N_12047,N_14662);
and U20488 (N_20488,N_15218,N_14740);
xor U20489 (N_20489,N_15931,N_14538);
nand U20490 (N_20490,N_17909,N_17849);
or U20491 (N_20491,N_14731,N_13559);
and U20492 (N_20492,N_17654,N_14088);
and U20493 (N_20493,N_12561,N_15629);
or U20494 (N_20494,N_12210,N_13502);
nand U20495 (N_20495,N_13711,N_17810);
or U20496 (N_20496,N_12319,N_16811);
nand U20497 (N_20497,N_15407,N_16015);
nor U20498 (N_20498,N_14932,N_17825);
xnor U20499 (N_20499,N_13295,N_14672);
or U20500 (N_20500,N_12019,N_16735);
xor U20501 (N_20501,N_13851,N_13826);
nor U20502 (N_20502,N_14859,N_12286);
or U20503 (N_20503,N_16271,N_15705);
and U20504 (N_20504,N_17302,N_15276);
nor U20505 (N_20505,N_12388,N_17995);
and U20506 (N_20506,N_15602,N_17398);
or U20507 (N_20507,N_17289,N_15268);
nor U20508 (N_20508,N_17818,N_17821);
or U20509 (N_20509,N_15097,N_17579);
nor U20510 (N_20510,N_16634,N_17137);
or U20511 (N_20511,N_12488,N_16635);
nand U20512 (N_20512,N_14392,N_16778);
and U20513 (N_20513,N_16078,N_13193);
or U20514 (N_20514,N_17278,N_16097);
nand U20515 (N_20515,N_14459,N_17740);
nand U20516 (N_20516,N_13096,N_13383);
nand U20517 (N_20517,N_13171,N_15752);
or U20518 (N_20518,N_13112,N_16447);
nand U20519 (N_20519,N_17640,N_16022);
xor U20520 (N_20520,N_16774,N_17593);
nor U20521 (N_20521,N_14034,N_16533);
nor U20522 (N_20522,N_17505,N_13870);
nand U20523 (N_20523,N_13785,N_13297);
xnor U20524 (N_20524,N_13333,N_13552);
and U20525 (N_20525,N_17774,N_14355);
and U20526 (N_20526,N_16215,N_13178);
nand U20527 (N_20527,N_17186,N_12252);
xor U20528 (N_20528,N_13393,N_12879);
and U20529 (N_20529,N_17435,N_15918);
nand U20530 (N_20530,N_14002,N_12864);
and U20531 (N_20531,N_15221,N_14948);
or U20532 (N_20532,N_16880,N_17917);
or U20533 (N_20533,N_17391,N_14285);
nor U20534 (N_20534,N_12311,N_12745);
xnor U20535 (N_20535,N_17819,N_17556);
nor U20536 (N_20536,N_15669,N_14234);
xor U20537 (N_20537,N_13553,N_17447);
xnor U20538 (N_20538,N_15618,N_15164);
xor U20539 (N_20539,N_15041,N_14472);
nor U20540 (N_20540,N_14025,N_17417);
and U20541 (N_20541,N_17845,N_17473);
xnor U20542 (N_20542,N_16886,N_17800);
xnor U20543 (N_20543,N_16742,N_16365);
nor U20544 (N_20544,N_14085,N_14113);
xnor U20545 (N_20545,N_17570,N_13376);
and U20546 (N_20546,N_13963,N_17884);
xnor U20547 (N_20547,N_14979,N_15709);
or U20548 (N_20548,N_13792,N_15760);
and U20549 (N_20549,N_16698,N_13519);
nand U20550 (N_20550,N_13438,N_14004);
nor U20551 (N_20551,N_13652,N_16258);
or U20552 (N_20552,N_13311,N_17664);
nor U20553 (N_20553,N_17309,N_12177);
nand U20554 (N_20554,N_17862,N_16555);
or U20555 (N_20555,N_16694,N_13099);
xor U20556 (N_20556,N_14977,N_16995);
or U20557 (N_20557,N_13131,N_12587);
and U20558 (N_20558,N_17967,N_17381);
or U20559 (N_20559,N_17493,N_15490);
nand U20560 (N_20560,N_15966,N_17587);
or U20561 (N_20561,N_14533,N_17824);
and U20562 (N_20562,N_14350,N_14385);
nand U20563 (N_20563,N_13736,N_14458);
xor U20564 (N_20564,N_14853,N_12200);
or U20565 (N_20565,N_14557,N_13479);
and U20566 (N_20566,N_17295,N_14427);
and U20567 (N_20567,N_16542,N_13403);
nand U20568 (N_20568,N_17651,N_16338);
or U20569 (N_20569,N_13662,N_15175);
or U20570 (N_20570,N_13599,N_14334);
and U20571 (N_20571,N_16779,N_15716);
nor U20572 (N_20572,N_13028,N_13699);
nand U20573 (N_20573,N_14819,N_13453);
nand U20574 (N_20574,N_15487,N_16300);
nand U20575 (N_20575,N_14507,N_16354);
and U20576 (N_20576,N_15932,N_12678);
xor U20577 (N_20577,N_13530,N_15475);
or U20578 (N_20578,N_12549,N_13670);
and U20579 (N_20579,N_12754,N_12367);
nor U20580 (N_20580,N_14329,N_15009);
nand U20581 (N_20581,N_13948,N_15484);
or U20582 (N_20582,N_16821,N_14797);
and U20583 (N_20583,N_17206,N_12886);
xnor U20584 (N_20584,N_12035,N_14768);
or U20585 (N_20585,N_17333,N_15214);
xnor U20586 (N_20586,N_17838,N_13377);
and U20587 (N_20587,N_13629,N_12661);
and U20588 (N_20588,N_17236,N_16108);
or U20589 (N_20589,N_12871,N_12377);
xor U20590 (N_20590,N_15372,N_13609);
and U20591 (N_20591,N_12029,N_13679);
nor U20592 (N_20592,N_16020,N_14479);
xor U20593 (N_20593,N_14173,N_13256);
and U20594 (N_20594,N_13505,N_14428);
and U20595 (N_20595,N_14222,N_16341);
nand U20596 (N_20596,N_17585,N_16581);
nor U20597 (N_20597,N_13710,N_17426);
nor U20598 (N_20598,N_12064,N_14221);
xor U20599 (N_20599,N_12428,N_12668);
or U20600 (N_20600,N_12651,N_13072);
or U20601 (N_20601,N_13644,N_14589);
nor U20602 (N_20602,N_17977,N_15696);
xnor U20603 (N_20603,N_17886,N_12986);
and U20604 (N_20604,N_13466,N_16280);
nor U20605 (N_20605,N_12782,N_14246);
xnor U20606 (N_20606,N_13538,N_14097);
and U20607 (N_20607,N_13648,N_16876);
and U20608 (N_20608,N_16282,N_17092);
or U20609 (N_20609,N_16081,N_13523);
nand U20610 (N_20610,N_12191,N_17832);
and U20611 (N_20611,N_16906,N_17554);
nand U20612 (N_20612,N_12666,N_13527);
or U20613 (N_20613,N_17799,N_17034);
nand U20614 (N_20614,N_16206,N_12117);
xor U20615 (N_20615,N_16959,N_12575);
or U20616 (N_20616,N_16584,N_17573);
and U20617 (N_20617,N_14478,N_16848);
and U20618 (N_20618,N_16601,N_15689);
or U20619 (N_20619,N_13829,N_16043);
or U20620 (N_20620,N_12915,N_15780);
nand U20621 (N_20621,N_17647,N_15726);
nand U20622 (N_20622,N_14376,N_12185);
xor U20623 (N_20623,N_14162,N_12108);
nand U20624 (N_20624,N_13518,N_17171);
xor U20625 (N_20625,N_15388,N_14216);
nor U20626 (N_20626,N_15190,N_16470);
and U20627 (N_20627,N_17330,N_13606);
nand U20628 (N_20628,N_14815,N_15406);
or U20629 (N_20629,N_12590,N_17565);
or U20630 (N_20630,N_17986,N_12647);
or U20631 (N_20631,N_15073,N_13554);
and U20632 (N_20632,N_16526,N_16370);
xnor U20633 (N_20633,N_15673,N_14877);
nor U20634 (N_20634,N_16598,N_14663);
nand U20635 (N_20635,N_17747,N_13243);
nor U20636 (N_20636,N_15113,N_14158);
nand U20637 (N_20637,N_16587,N_17718);
or U20638 (N_20638,N_14381,N_16492);
xnor U20639 (N_20639,N_16307,N_17024);
or U20640 (N_20640,N_12545,N_15567);
nand U20641 (N_20641,N_14621,N_13937);
nand U20642 (N_20642,N_13808,N_12591);
xnor U20643 (N_20643,N_17322,N_16874);
and U20644 (N_20644,N_15012,N_14907);
xor U20645 (N_20645,N_16796,N_13036);
nand U20646 (N_20646,N_16208,N_17392);
or U20647 (N_20647,N_14201,N_16688);
and U20648 (N_20648,N_12826,N_14562);
and U20649 (N_20649,N_14687,N_12878);
and U20650 (N_20650,N_17464,N_13762);
xor U20651 (N_20651,N_14322,N_14056);
and U20652 (N_20652,N_12182,N_12461);
or U20653 (N_20653,N_14078,N_17185);
or U20654 (N_20654,N_14837,N_12225);
nor U20655 (N_20655,N_15034,N_12350);
nand U20656 (N_20656,N_17891,N_16511);
nor U20657 (N_20657,N_14643,N_15349);
nand U20658 (N_20658,N_17108,N_12819);
or U20659 (N_20659,N_12494,N_13000);
nand U20660 (N_20660,N_13240,N_17841);
xor U20661 (N_20661,N_13341,N_14584);
nor U20662 (N_20662,N_13038,N_16415);
nand U20663 (N_20663,N_15840,N_14324);
or U20664 (N_20664,N_15607,N_12850);
and U20665 (N_20665,N_13032,N_13407);
or U20666 (N_20666,N_14431,N_12629);
nor U20667 (N_20667,N_12694,N_16827);
nand U20668 (N_20668,N_17889,N_16622);
xnor U20669 (N_20669,N_14415,N_17406);
xnor U20670 (N_20670,N_13282,N_14007);
and U20671 (N_20671,N_14546,N_14335);
nor U20672 (N_20672,N_12462,N_15114);
nor U20673 (N_20673,N_17561,N_13206);
nand U20674 (N_20674,N_12818,N_16211);
nand U20675 (N_20675,N_13660,N_13308);
xnor U20676 (N_20676,N_13956,N_13285);
nand U20677 (N_20677,N_13993,N_15837);
nand U20678 (N_20678,N_12149,N_15814);
nand U20679 (N_20679,N_14692,N_12771);
or U20680 (N_20680,N_14861,N_14817);
nor U20681 (N_20681,N_13804,N_14788);
nor U20682 (N_20682,N_14937,N_17331);
xor U20683 (N_20683,N_12532,N_13597);
and U20684 (N_20684,N_14985,N_15319);
nor U20685 (N_20685,N_13342,N_13714);
nor U20686 (N_20686,N_15090,N_16073);
nand U20687 (N_20687,N_12300,N_14564);
and U20688 (N_20688,N_14152,N_15217);
xnor U20689 (N_20689,N_12089,N_13271);
xor U20690 (N_20690,N_12752,N_12477);
nor U20691 (N_20691,N_12692,N_17056);
nor U20692 (N_20692,N_15081,N_14457);
nor U20693 (N_20693,N_15763,N_16705);
or U20694 (N_20694,N_17038,N_13501);
nand U20695 (N_20695,N_14233,N_14033);
xnor U20696 (N_20696,N_14053,N_14467);
nand U20697 (N_20697,N_16156,N_16087);
nand U20698 (N_20698,N_16567,N_17876);
and U20699 (N_20699,N_13394,N_16830);
nand U20700 (N_20700,N_14799,N_17332);
xor U20701 (N_20701,N_13757,N_14068);
nor U20702 (N_20702,N_17650,N_12552);
nand U20703 (N_20703,N_13318,N_14405);
nand U20704 (N_20704,N_15798,N_12226);
and U20705 (N_20705,N_14147,N_16648);
and U20706 (N_20706,N_14421,N_12991);
or U20707 (N_20707,N_14911,N_15191);
and U20708 (N_20708,N_16405,N_13971);
or U20709 (N_20709,N_14325,N_12195);
nand U20710 (N_20710,N_14609,N_17193);
nand U20711 (N_20711,N_13422,N_15481);
nor U20712 (N_20712,N_15240,N_15578);
xor U20713 (N_20713,N_15503,N_17281);
nor U20714 (N_20714,N_16799,N_14071);
xor U20715 (N_20715,N_17709,N_15911);
and U20716 (N_20716,N_13628,N_15496);
or U20717 (N_20717,N_14040,N_17925);
nand U20718 (N_20718,N_12847,N_13929);
and U20719 (N_20719,N_17626,N_17324);
or U20720 (N_20720,N_12747,N_16319);
xnor U20721 (N_20721,N_15316,N_16006);
nor U20722 (N_20722,N_12700,N_12352);
xor U20723 (N_20723,N_12649,N_14836);
and U20724 (N_20724,N_16461,N_17581);
nand U20725 (N_20725,N_14495,N_13137);
nor U20726 (N_20726,N_16127,N_17934);
and U20727 (N_20727,N_13866,N_16783);
nand U20728 (N_20728,N_17829,N_15135);
and U20729 (N_20729,N_14391,N_17531);
or U20730 (N_20730,N_15205,N_15384);
and U20731 (N_20731,N_17226,N_16432);
or U20732 (N_20732,N_14814,N_16165);
nor U20733 (N_20733,N_17081,N_14140);
or U20734 (N_20734,N_12758,N_13132);
and U20735 (N_20735,N_14348,N_13990);
nor U20736 (N_20736,N_15473,N_15950);
xnor U20737 (N_20737,N_15283,N_14645);
nand U20738 (N_20738,N_12565,N_12990);
or U20739 (N_20739,N_14825,N_16800);
and U20740 (N_20740,N_17415,N_15345);
nor U20741 (N_20741,N_13139,N_15676);
or U20742 (N_20742,N_15679,N_14555);
or U20743 (N_20743,N_12639,N_16724);
xor U20744 (N_20744,N_14858,N_12970);
nand U20745 (N_20745,N_15070,N_16987);
nand U20746 (N_20746,N_15479,N_14633);
and U20747 (N_20747,N_15556,N_14134);
and U20748 (N_20748,N_15792,N_13742);
nand U20749 (N_20749,N_13601,N_15069);
nand U20750 (N_20750,N_16227,N_13768);
nor U20751 (N_20751,N_14049,N_17541);
xnor U20752 (N_20752,N_13684,N_12883);
and U20753 (N_20753,N_15163,N_12305);
and U20754 (N_20754,N_15897,N_17434);
and U20755 (N_20755,N_17353,N_13676);
nand U20756 (N_20756,N_12953,N_16972);
and U20757 (N_20757,N_16861,N_16576);
or U20758 (N_20758,N_12371,N_14941);
xor U20759 (N_20759,N_13371,N_16941);
nand U20760 (N_20760,N_12900,N_14654);
xnor U20761 (N_20761,N_15305,N_15824);
or U20762 (N_20762,N_17743,N_15171);
or U20763 (N_20763,N_17031,N_16363);
or U20764 (N_20764,N_13430,N_15172);
or U20765 (N_20765,N_14344,N_16914);
nor U20766 (N_20766,N_15024,N_13716);
nor U20767 (N_20767,N_14639,N_17898);
nor U20768 (N_20768,N_16539,N_15963);
nor U20769 (N_20769,N_15700,N_14998);
xnor U20770 (N_20770,N_14605,N_15639);
and U20771 (N_20771,N_13006,N_15121);
or U20772 (N_20772,N_14125,N_17628);
xor U20773 (N_20773,N_17029,N_14874);
nor U20774 (N_20774,N_14843,N_16912);
nor U20775 (N_20775,N_15547,N_15331);
nor U20776 (N_20776,N_13339,N_13514);
and U20777 (N_20777,N_15189,N_17252);
nor U20778 (N_20778,N_13667,N_14659);
xnor U20779 (N_20779,N_13607,N_16218);
xor U20780 (N_20780,N_12006,N_16189);
nor U20781 (N_20781,N_13934,N_17630);
nor U20782 (N_20782,N_15313,N_14526);
and U20783 (N_20783,N_15796,N_14027);
nand U20784 (N_20784,N_14422,N_15906);
nand U20785 (N_20785,N_17926,N_17155);
nor U20786 (N_20786,N_17861,N_12559);
or U20787 (N_20787,N_12656,N_15141);
and U20788 (N_20788,N_16885,N_16857);
or U20789 (N_20789,N_17781,N_13570);
nand U20790 (N_20790,N_12301,N_15229);
and U20791 (N_20791,N_16342,N_15778);
nor U20792 (N_20792,N_14332,N_13844);
or U20793 (N_20793,N_16756,N_15900);
nand U20794 (N_20794,N_14432,N_16996);
nor U20795 (N_20795,N_12914,N_12395);
xnor U20796 (N_20796,N_16024,N_13276);
or U20797 (N_20797,N_15308,N_14956);
xor U20798 (N_20798,N_15864,N_15145);
nor U20799 (N_20799,N_16133,N_13284);
nor U20800 (N_20800,N_16160,N_15992);
and U20801 (N_20801,N_14559,N_15211);
nand U20802 (N_20802,N_14447,N_17759);
nand U20803 (N_20803,N_15232,N_17567);
and U20804 (N_20804,N_13463,N_14895);
and U20805 (N_20805,N_15594,N_14241);
or U20806 (N_20806,N_12469,N_14245);
or U20807 (N_20807,N_15075,N_17782);
nor U20808 (N_20808,N_14279,N_13885);
xor U20809 (N_20809,N_15136,N_15821);
and U20810 (N_20810,N_13720,N_13427);
nor U20811 (N_20811,N_16276,N_16898);
xnor U20812 (N_20812,N_12855,N_14014);
or U20813 (N_20813,N_16420,N_13769);
nor U20814 (N_20814,N_12072,N_16169);
or U20815 (N_20815,N_15967,N_17500);
or U20816 (N_20816,N_16665,N_17178);
nand U20817 (N_20817,N_16082,N_15774);
xnor U20818 (N_20818,N_14872,N_14974);
xnor U20819 (N_20819,N_15600,N_16104);
xor U20820 (N_20820,N_14273,N_13265);
xor U20821 (N_20821,N_14572,N_16863);
or U20822 (N_20822,N_13471,N_16768);
xor U20823 (N_20823,N_13251,N_16746);
nand U20824 (N_20824,N_17495,N_14184);
and U20825 (N_20825,N_13686,N_17634);
and U20826 (N_20826,N_13242,N_14036);
nor U20827 (N_20827,N_13748,N_17285);
xnor U20828 (N_20828,N_17388,N_14833);
nor U20829 (N_20829,N_17952,N_12162);
and U20830 (N_20830,N_16145,N_12368);
nand U20831 (N_20831,N_12090,N_12690);
nor U20832 (N_20832,N_17667,N_12211);
or U20833 (N_20833,N_15326,N_15119);
nand U20834 (N_20834,N_15835,N_13014);
xnor U20835 (N_20835,N_13410,N_13307);
xnor U20836 (N_20836,N_12163,N_15628);
and U20837 (N_20837,N_12569,N_17414);
nor U20838 (N_20838,N_12224,N_12732);
and U20839 (N_20839,N_12691,N_17770);
nand U20840 (N_20840,N_14615,N_12925);
xor U20841 (N_20841,N_16446,N_17733);
and U20842 (N_20842,N_12937,N_17491);
nand U20843 (N_20843,N_17204,N_14118);
nand U20844 (N_20844,N_17317,N_12849);
or U20845 (N_20845,N_13155,N_14136);
nor U20846 (N_20846,N_13723,N_13429);
nor U20847 (N_20847,N_12481,N_17708);
xnor U20848 (N_20848,N_16718,N_13402);
xnor U20849 (N_20849,N_12658,N_16092);
nor U20850 (N_20850,N_15266,N_13084);
and U20851 (N_20851,N_13974,N_17465);
nand U20852 (N_20852,N_15167,N_16671);
xor U20853 (N_20853,N_13462,N_13057);
xor U20854 (N_20854,N_14191,N_16031);
nand U20855 (N_20855,N_15927,N_12777);
nor U20856 (N_20856,N_16355,N_12505);
nor U20857 (N_20857,N_15516,N_13813);
or U20858 (N_20858,N_12186,N_14499);
and U20859 (N_20859,N_13259,N_12348);
and U20860 (N_20860,N_12160,N_15880);
or U20861 (N_20861,N_16292,N_15065);
nor U20862 (N_20862,N_14051,N_17642);
xor U20863 (N_20863,N_17560,N_14318);
xnor U20864 (N_20864,N_15151,N_14314);
or U20865 (N_20865,N_16592,N_12753);
nor U20866 (N_20866,N_14321,N_15398);
nor U20867 (N_20867,N_16454,N_17694);
xnor U20868 (N_20868,N_16842,N_12929);
xor U20869 (N_20869,N_15886,N_15972);
nor U20870 (N_20870,N_16039,N_17124);
nand U20871 (N_20871,N_15509,N_16537);
nand U20872 (N_20872,N_14749,N_14601);
xor U20873 (N_20873,N_12456,N_12685);
nand U20874 (N_20874,N_16847,N_16489);
or U20875 (N_20875,N_13793,N_12287);
and U20876 (N_20876,N_17012,N_14045);
xor U20877 (N_20877,N_12885,N_15564);
and U20878 (N_20878,N_15329,N_15627);
nand U20879 (N_20879,N_17183,N_15300);
or U20880 (N_20880,N_13647,N_15209);
nand U20881 (N_20881,N_17325,N_12414);
and U20882 (N_20882,N_15502,N_14207);
and U20883 (N_20883,N_12294,N_14631);
and U20884 (N_20884,N_17778,N_16154);
nor U20885 (N_20885,N_14992,N_16362);
nor U20886 (N_20886,N_13105,N_13509);
nand U20887 (N_20887,N_12715,N_14404);
and U20888 (N_20888,N_16157,N_17277);
or U20889 (N_20889,N_12221,N_12502);
nor U20890 (N_20890,N_16101,N_12402);
nor U20891 (N_20891,N_16052,N_14238);
nand U20892 (N_20892,N_12062,N_13083);
or U20893 (N_20893,N_16458,N_16310);
or U20894 (N_20894,N_16658,N_12942);
nand U20895 (N_20895,N_16191,N_15825);
and U20896 (N_20896,N_15423,N_14613);
nor U20897 (N_20897,N_14326,N_16498);
nor U20898 (N_20898,N_13545,N_17726);
and U20899 (N_20899,N_13843,N_13143);
nor U20900 (N_20900,N_17542,N_13485);
xor U20901 (N_20901,N_13351,N_15661);
nand U20902 (N_20902,N_14598,N_14706);
and U20903 (N_20903,N_17562,N_15924);
nor U20904 (N_20904,N_15122,N_15766);
xor U20905 (N_20905,N_15797,N_15647);
or U20906 (N_20906,N_16219,N_12809);
nand U20907 (N_20907,N_12563,N_14337);
and U20908 (N_20908,N_17078,N_14363);
and U20909 (N_20909,N_16900,N_17213);
and U20910 (N_20910,N_12104,N_14734);
xnor U20911 (N_20911,N_14487,N_15939);
and U20912 (N_20912,N_13003,N_14112);
and U20913 (N_20913,N_17225,N_15623);
xnor U20914 (N_20914,N_12623,N_16326);
xnor U20915 (N_20915,N_15441,N_14365);
xor U20916 (N_20916,N_12980,N_12556);
nand U20917 (N_20917,N_17304,N_12387);
and U20918 (N_20918,N_17221,N_13863);
or U20919 (N_20919,N_14784,N_14696);
or U20920 (N_20920,N_13470,N_15059);
nor U20921 (N_20921,N_15787,N_17037);
nor U20922 (N_20922,N_14758,N_13745);
and U20923 (N_20923,N_12760,N_15105);
nor U20924 (N_20924,N_15107,N_15819);
or U20925 (N_20925,N_13051,N_15751);
or U20926 (N_20926,N_13595,N_13717);
nor U20927 (N_20927,N_12633,N_17054);
xor U20928 (N_20928,N_13712,N_12567);
and U20929 (N_20929,N_13744,N_15732);
and U20930 (N_20930,N_16503,N_16732);
nand U20931 (N_20931,N_12041,N_14917);
xor U20932 (N_20932,N_13209,N_17875);
nor U20933 (N_20933,N_17857,N_16650);
nor U20934 (N_20934,N_17130,N_15224);
nand U20935 (N_20935,N_13834,N_12283);
and U20936 (N_20936,N_13585,N_16692);
or U20937 (N_20937,N_16287,N_12018);
nor U20938 (N_20938,N_17103,N_13205);
or U20939 (N_20939,N_17940,N_15376);
xnor U20940 (N_20940,N_14398,N_14364);
nand U20941 (N_20941,N_16254,N_14592);
nand U20942 (N_20942,N_17412,N_17701);
nand U20943 (N_20943,N_16230,N_14109);
and U20944 (N_20944,N_17695,N_13398);
or U20945 (N_20945,N_13071,N_17158);
or U20946 (N_20946,N_14520,N_14360);
or U20947 (N_20947,N_13688,N_15862);
xnor U20948 (N_20948,N_15454,N_12105);
or U20949 (N_20949,N_17175,N_13037);
xor U20950 (N_20950,N_14239,N_17340);
or U20951 (N_20951,N_16229,N_13703);
xor U20952 (N_20952,N_16036,N_14275);
xor U20953 (N_20953,N_16725,N_13156);
and U20954 (N_20954,N_17113,N_14732);
xnor U20955 (N_20955,N_12479,N_16571);
nand U20956 (N_20956,N_15802,N_13127);
nor U20957 (N_20957,N_15856,N_15625);
nand U20958 (N_20958,N_14675,N_13931);
or U20959 (N_20959,N_14163,N_12017);
nand U20960 (N_20960,N_13287,N_14043);
nand U20961 (N_20961,N_12531,N_12399);
nand U20962 (N_20962,N_17788,N_12975);
xnor U20963 (N_20963,N_14975,N_16769);
xnor U20964 (N_20964,N_16516,N_16932);
or U20965 (N_20965,N_12675,N_15758);
nor U20966 (N_20966,N_12994,N_17811);
or U20967 (N_20967,N_14488,N_17840);
xor U20968 (N_20968,N_12338,N_17503);
and U20969 (N_20969,N_14500,N_14144);
nand U20970 (N_20970,N_15404,N_15654);
nand U20971 (N_20971,N_12959,N_12483);
or U20972 (N_20972,N_12052,N_15170);
nand U20973 (N_20973,N_15829,N_13435);
or U20974 (N_20974,N_14124,N_13936);
and U20975 (N_20975,N_17262,N_17931);
or U20976 (N_20976,N_12125,N_15538);
or U20977 (N_20977,N_14465,N_17703);
or U20978 (N_20978,N_13011,N_17147);
xor U20979 (N_20979,N_14196,N_14896);
nand U20980 (N_20980,N_13691,N_13636);
nand U20981 (N_20981,N_15568,N_16621);
and U20982 (N_20982,N_15572,N_14303);
nand U20983 (N_20983,N_12755,N_13653);
nor U20984 (N_20984,N_15144,N_12845);
and U20985 (N_20985,N_12147,N_16753);
and U20986 (N_20986,N_16962,N_15975);
and U20987 (N_20987,N_12810,N_16001);
nor U20988 (N_20988,N_13525,N_13961);
or U20989 (N_20989,N_13201,N_16202);
nor U20990 (N_20990,N_14393,N_17533);
xnor U20991 (N_20991,N_13280,N_16166);
and U20992 (N_20992,N_14424,N_15470);
nand U20993 (N_20993,N_17460,N_15920);
or U20994 (N_20994,N_16680,N_15606);
and U20995 (N_20995,N_13369,N_14667);
and U20996 (N_20996,N_17149,N_17410);
or U20997 (N_20997,N_16562,N_14503);
nor U20998 (N_20998,N_15178,N_15925);
nor U20999 (N_20999,N_15278,N_13189);
xnor U21000 (N_21000,N_14049,N_15746);
and U21001 (N_21001,N_13860,N_16976);
nor U21002 (N_21002,N_13109,N_17566);
or U21003 (N_21003,N_15991,N_14298);
nor U21004 (N_21004,N_17244,N_13781);
or U21005 (N_21005,N_12272,N_14277);
or U21006 (N_21006,N_16551,N_13965);
xor U21007 (N_21007,N_12613,N_16766);
and U21008 (N_21008,N_13373,N_15499);
nor U21009 (N_21009,N_17137,N_13200);
or U21010 (N_21010,N_12778,N_17670);
nand U21011 (N_21011,N_12632,N_14453);
or U21012 (N_21012,N_14783,N_15967);
or U21013 (N_21013,N_12308,N_15303);
and U21014 (N_21014,N_15546,N_15683);
or U21015 (N_21015,N_15260,N_16256);
or U21016 (N_21016,N_17780,N_17506);
nand U21017 (N_21017,N_13390,N_16675);
or U21018 (N_21018,N_12510,N_16358);
and U21019 (N_21019,N_17279,N_16310);
or U21020 (N_21020,N_16029,N_13021);
and U21021 (N_21021,N_16836,N_17262);
nor U21022 (N_21022,N_15229,N_12863);
nand U21023 (N_21023,N_15643,N_12261);
or U21024 (N_21024,N_14868,N_12457);
nand U21025 (N_21025,N_17608,N_14742);
nand U21026 (N_21026,N_17203,N_12245);
xor U21027 (N_21027,N_13470,N_17466);
nor U21028 (N_21028,N_17628,N_15615);
nand U21029 (N_21029,N_14545,N_15872);
nor U21030 (N_21030,N_14497,N_13707);
xor U21031 (N_21031,N_14708,N_12990);
nor U21032 (N_21032,N_13342,N_12253);
and U21033 (N_21033,N_13136,N_17190);
nor U21034 (N_21034,N_14212,N_16728);
nand U21035 (N_21035,N_12387,N_14906);
nor U21036 (N_21036,N_17961,N_12971);
and U21037 (N_21037,N_12112,N_14027);
xnor U21038 (N_21038,N_16809,N_16671);
nor U21039 (N_21039,N_14549,N_13745);
nor U21040 (N_21040,N_16055,N_16513);
and U21041 (N_21041,N_17506,N_16751);
xnor U21042 (N_21042,N_17834,N_12825);
and U21043 (N_21043,N_15828,N_17619);
nand U21044 (N_21044,N_15306,N_15088);
xnor U21045 (N_21045,N_17733,N_15196);
or U21046 (N_21046,N_13177,N_16765);
and U21047 (N_21047,N_16506,N_13444);
xnor U21048 (N_21048,N_12172,N_13440);
and U21049 (N_21049,N_15865,N_15929);
nor U21050 (N_21050,N_12627,N_16508);
and U21051 (N_21051,N_15014,N_14407);
and U21052 (N_21052,N_12341,N_15406);
and U21053 (N_21053,N_13695,N_12068);
or U21054 (N_21054,N_13387,N_13806);
nand U21055 (N_21055,N_17329,N_17754);
or U21056 (N_21056,N_14222,N_17441);
and U21057 (N_21057,N_15631,N_13836);
nand U21058 (N_21058,N_12773,N_17097);
and U21059 (N_21059,N_12906,N_14577);
nor U21060 (N_21060,N_16631,N_13573);
and U21061 (N_21061,N_16882,N_13486);
or U21062 (N_21062,N_16995,N_12575);
xnor U21063 (N_21063,N_13876,N_16264);
xnor U21064 (N_21064,N_17522,N_16159);
and U21065 (N_21065,N_16512,N_12732);
and U21066 (N_21066,N_15195,N_15556);
and U21067 (N_21067,N_15458,N_16756);
or U21068 (N_21068,N_17893,N_14538);
xor U21069 (N_21069,N_16514,N_16795);
or U21070 (N_21070,N_12901,N_16094);
or U21071 (N_21071,N_17279,N_15893);
nand U21072 (N_21072,N_12901,N_14077);
and U21073 (N_21073,N_15469,N_17131);
or U21074 (N_21074,N_16963,N_14762);
nand U21075 (N_21075,N_13974,N_16750);
and U21076 (N_21076,N_14079,N_14276);
nor U21077 (N_21077,N_14922,N_15704);
xor U21078 (N_21078,N_15426,N_12095);
nand U21079 (N_21079,N_14284,N_12780);
xor U21080 (N_21080,N_16515,N_16700);
nor U21081 (N_21081,N_12873,N_15448);
and U21082 (N_21082,N_13255,N_14246);
nor U21083 (N_21083,N_15601,N_13222);
xor U21084 (N_21084,N_12235,N_17438);
xnor U21085 (N_21085,N_13340,N_14585);
xnor U21086 (N_21086,N_12990,N_14591);
nor U21087 (N_21087,N_15114,N_16468);
xor U21088 (N_21088,N_13473,N_14723);
or U21089 (N_21089,N_12154,N_16797);
nor U21090 (N_21090,N_16508,N_12271);
or U21091 (N_21091,N_17850,N_14380);
or U21092 (N_21092,N_16692,N_12447);
nand U21093 (N_21093,N_12411,N_17681);
xnor U21094 (N_21094,N_12319,N_13339);
nor U21095 (N_21095,N_13526,N_14220);
or U21096 (N_21096,N_12303,N_15324);
and U21097 (N_21097,N_13336,N_17182);
nor U21098 (N_21098,N_13375,N_16705);
nor U21099 (N_21099,N_14005,N_13150);
nor U21100 (N_21100,N_17923,N_12217);
and U21101 (N_21101,N_17289,N_13789);
nand U21102 (N_21102,N_13020,N_13840);
or U21103 (N_21103,N_13871,N_16606);
xor U21104 (N_21104,N_17028,N_14246);
and U21105 (N_21105,N_15128,N_15767);
nand U21106 (N_21106,N_15463,N_16409);
or U21107 (N_21107,N_14064,N_12719);
nor U21108 (N_21108,N_13780,N_14205);
or U21109 (N_21109,N_17703,N_12806);
xnor U21110 (N_21110,N_16724,N_12205);
or U21111 (N_21111,N_14999,N_13209);
nor U21112 (N_21112,N_12436,N_15215);
nand U21113 (N_21113,N_15472,N_12357);
nand U21114 (N_21114,N_15977,N_14471);
nand U21115 (N_21115,N_15500,N_15226);
xor U21116 (N_21116,N_17706,N_14554);
or U21117 (N_21117,N_16283,N_12973);
nor U21118 (N_21118,N_15659,N_13564);
or U21119 (N_21119,N_16612,N_16483);
or U21120 (N_21120,N_15230,N_14596);
and U21121 (N_21121,N_16329,N_14889);
nand U21122 (N_21122,N_12909,N_12592);
and U21123 (N_21123,N_17298,N_13565);
xor U21124 (N_21124,N_16542,N_14941);
or U21125 (N_21125,N_15343,N_12487);
and U21126 (N_21126,N_17837,N_17367);
nand U21127 (N_21127,N_17122,N_12260);
nand U21128 (N_21128,N_16487,N_13394);
and U21129 (N_21129,N_17533,N_15660);
xnor U21130 (N_21130,N_13853,N_16178);
or U21131 (N_21131,N_15452,N_16856);
nor U21132 (N_21132,N_15227,N_13804);
nor U21133 (N_21133,N_16245,N_16189);
xnor U21134 (N_21134,N_14841,N_16104);
nand U21135 (N_21135,N_14878,N_14452);
xor U21136 (N_21136,N_14273,N_13809);
xor U21137 (N_21137,N_16674,N_12274);
xor U21138 (N_21138,N_15004,N_14962);
or U21139 (N_21139,N_13899,N_16573);
nor U21140 (N_21140,N_16395,N_15289);
nor U21141 (N_21141,N_13602,N_14244);
or U21142 (N_21142,N_13025,N_12813);
and U21143 (N_21143,N_16900,N_17349);
or U21144 (N_21144,N_13805,N_12891);
nor U21145 (N_21145,N_16872,N_16496);
nor U21146 (N_21146,N_17506,N_12907);
nor U21147 (N_21147,N_14121,N_14577);
or U21148 (N_21148,N_14541,N_12515);
and U21149 (N_21149,N_15943,N_17918);
or U21150 (N_21150,N_17589,N_17599);
nand U21151 (N_21151,N_13220,N_17866);
or U21152 (N_21152,N_16477,N_14729);
nand U21153 (N_21153,N_17337,N_14546);
xnor U21154 (N_21154,N_16046,N_15151);
nor U21155 (N_21155,N_16206,N_14978);
and U21156 (N_21156,N_17183,N_15796);
or U21157 (N_21157,N_14244,N_12390);
or U21158 (N_21158,N_17809,N_17102);
nor U21159 (N_21159,N_15454,N_13836);
and U21160 (N_21160,N_17710,N_12760);
xnor U21161 (N_21161,N_14838,N_16772);
and U21162 (N_21162,N_16979,N_14320);
nand U21163 (N_21163,N_12425,N_17758);
xnor U21164 (N_21164,N_17121,N_14380);
and U21165 (N_21165,N_14501,N_13521);
xor U21166 (N_21166,N_12809,N_12985);
and U21167 (N_21167,N_14583,N_13990);
nor U21168 (N_21168,N_12072,N_13456);
nand U21169 (N_21169,N_12316,N_15200);
nor U21170 (N_21170,N_12301,N_13558);
nand U21171 (N_21171,N_16066,N_12783);
nand U21172 (N_21172,N_15034,N_16090);
nor U21173 (N_21173,N_13082,N_13407);
and U21174 (N_21174,N_15892,N_14242);
nand U21175 (N_21175,N_13056,N_17752);
or U21176 (N_21176,N_14800,N_12657);
xor U21177 (N_21177,N_12847,N_17986);
xor U21178 (N_21178,N_13066,N_16972);
and U21179 (N_21179,N_16406,N_15868);
and U21180 (N_21180,N_17932,N_13338);
nand U21181 (N_21181,N_13972,N_17946);
nor U21182 (N_21182,N_15234,N_16219);
xor U21183 (N_21183,N_15075,N_17992);
xnor U21184 (N_21184,N_14668,N_16508);
xor U21185 (N_21185,N_14157,N_13154);
nand U21186 (N_21186,N_15948,N_12943);
nand U21187 (N_21187,N_17962,N_14293);
xor U21188 (N_21188,N_12252,N_16681);
or U21189 (N_21189,N_15596,N_12189);
or U21190 (N_21190,N_14582,N_12210);
and U21191 (N_21191,N_15584,N_15852);
or U21192 (N_21192,N_17632,N_15754);
and U21193 (N_21193,N_12886,N_15440);
and U21194 (N_21194,N_16876,N_16232);
xnor U21195 (N_21195,N_12978,N_12838);
nor U21196 (N_21196,N_17082,N_17914);
nand U21197 (N_21197,N_15753,N_15579);
xor U21198 (N_21198,N_15636,N_12240);
xor U21199 (N_21199,N_16986,N_17248);
nor U21200 (N_21200,N_15038,N_15567);
nand U21201 (N_21201,N_16322,N_17639);
and U21202 (N_21202,N_12363,N_12464);
or U21203 (N_21203,N_12456,N_14865);
nor U21204 (N_21204,N_16547,N_15191);
and U21205 (N_21205,N_17017,N_15181);
and U21206 (N_21206,N_14962,N_17791);
or U21207 (N_21207,N_13283,N_15812);
nand U21208 (N_21208,N_14282,N_14845);
or U21209 (N_21209,N_12524,N_16376);
or U21210 (N_21210,N_16819,N_13406);
nor U21211 (N_21211,N_17645,N_13168);
and U21212 (N_21212,N_13537,N_17017);
nand U21213 (N_21213,N_15610,N_17680);
xor U21214 (N_21214,N_15359,N_16295);
nor U21215 (N_21215,N_15819,N_16271);
nand U21216 (N_21216,N_17754,N_13332);
or U21217 (N_21217,N_16427,N_12950);
nor U21218 (N_21218,N_12803,N_14142);
nand U21219 (N_21219,N_14329,N_16480);
nand U21220 (N_21220,N_13953,N_13359);
and U21221 (N_21221,N_12772,N_12113);
and U21222 (N_21222,N_14201,N_15906);
nand U21223 (N_21223,N_13278,N_14765);
or U21224 (N_21224,N_14255,N_16825);
and U21225 (N_21225,N_15319,N_12680);
or U21226 (N_21226,N_13353,N_12193);
xnor U21227 (N_21227,N_14247,N_13349);
or U21228 (N_21228,N_17704,N_16051);
nand U21229 (N_21229,N_15346,N_12889);
nand U21230 (N_21230,N_14052,N_17265);
xnor U21231 (N_21231,N_15570,N_12681);
and U21232 (N_21232,N_12413,N_16494);
nand U21233 (N_21233,N_17763,N_12170);
nand U21234 (N_21234,N_12112,N_13116);
nor U21235 (N_21235,N_15536,N_16907);
and U21236 (N_21236,N_14265,N_15050);
or U21237 (N_21237,N_16137,N_16717);
nand U21238 (N_21238,N_15495,N_15054);
or U21239 (N_21239,N_13500,N_16492);
and U21240 (N_21240,N_17085,N_13744);
nor U21241 (N_21241,N_15716,N_15216);
or U21242 (N_21242,N_13833,N_14672);
nor U21243 (N_21243,N_15874,N_12652);
or U21244 (N_21244,N_13830,N_13684);
nand U21245 (N_21245,N_15644,N_14472);
xnor U21246 (N_21246,N_12762,N_17587);
and U21247 (N_21247,N_13652,N_16605);
and U21248 (N_21248,N_12585,N_16046);
xnor U21249 (N_21249,N_16367,N_15410);
and U21250 (N_21250,N_17238,N_13547);
nand U21251 (N_21251,N_16327,N_16685);
nor U21252 (N_21252,N_13147,N_14851);
xnor U21253 (N_21253,N_14132,N_13939);
or U21254 (N_21254,N_17096,N_16739);
nand U21255 (N_21255,N_15556,N_17196);
xnor U21256 (N_21256,N_15234,N_15665);
nor U21257 (N_21257,N_16855,N_12891);
nand U21258 (N_21258,N_14435,N_17788);
or U21259 (N_21259,N_15404,N_13228);
nor U21260 (N_21260,N_15283,N_12047);
and U21261 (N_21261,N_14843,N_12775);
or U21262 (N_21262,N_13408,N_17246);
nor U21263 (N_21263,N_15783,N_17877);
nor U21264 (N_21264,N_14489,N_17098);
and U21265 (N_21265,N_16078,N_14847);
nor U21266 (N_21266,N_12303,N_15432);
and U21267 (N_21267,N_15673,N_13520);
nor U21268 (N_21268,N_16770,N_15628);
xnor U21269 (N_21269,N_12304,N_16877);
xor U21270 (N_21270,N_15214,N_13619);
nand U21271 (N_21271,N_14882,N_14337);
xnor U21272 (N_21272,N_17623,N_12444);
nand U21273 (N_21273,N_15011,N_17157);
nor U21274 (N_21274,N_16561,N_16433);
nand U21275 (N_21275,N_14391,N_13187);
xor U21276 (N_21276,N_16916,N_13026);
or U21277 (N_21277,N_15579,N_14712);
and U21278 (N_21278,N_15798,N_16388);
nand U21279 (N_21279,N_15247,N_16565);
nand U21280 (N_21280,N_17297,N_17394);
or U21281 (N_21281,N_12537,N_14797);
or U21282 (N_21282,N_17094,N_14842);
nor U21283 (N_21283,N_13538,N_16416);
nand U21284 (N_21284,N_13536,N_15155);
nand U21285 (N_21285,N_16070,N_16701);
and U21286 (N_21286,N_13319,N_14207);
and U21287 (N_21287,N_16504,N_16708);
xnor U21288 (N_21288,N_17218,N_17901);
or U21289 (N_21289,N_16129,N_17188);
nand U21290 (N_21290,N_17024,N_17733);
nor U21291 (N_21291,N_12605,N_13506);
or U21292 (N_21292,N_14035,N_16689);
nor U21293 (N_21293,N_15262,N_16487);
nor U21294 (N_21294,N_17932,N_12320);
nand U21295 (N_21295,N_13990,N_13219);
xor U21296 (N_21296,N_12334,N_13811);
and U21297 (N_21297,N_16737,N_16361);
xnor U21298 (N_21298,N_15303,N_15565);
nand U21299 (N_21299,N_13271,N_13768);
xnor U21300 (N_21300,N_14529,N_14701);
xor U21301 (N_21301,N_13960,N_16527);
and U21302 (N_21302,N_16737,N_14543);
nor U21303 (N_21303,N_15117,N_17131);
or U21304 (N_21304,N_16579,N_14393);
xor U21305 (N_21305,N_13264,N_14653);
xnor U21306 (N_21306,N_16978,N_16951);
or U21307 (N_21307,N_13737,N_14264);
xnor U21308 (N_21308,N_17817,N_13204);
xor U21309 (N_21309,N_12611,N_13557);
xnor U21310 (N_21310,N_13043,N_13204);
xor U21311 (N_21311,N_13451,N_16829);
and U21312 (N_21312,N_15851,N_12968);
or U21313 (N_21313,N_13122,N_13686);
nor U21314 (N_21314,N_13726,N_16012);
and U21315 (N_21315,N_15186,N_15555);
nand U21316 (N_21316,N_14254,N_12158);
nand U21317 (N_21317,N_13883,N_12737);
nand U21318 (N_21318,N_12485,N_12863);
and U21319 (N_21319,N_15363,N_14245);
and U21320 (N_21320,N_13421,N_13140);
nor U21321 (N_21321,N_17151,N_16132);
nand U21322 (N_21322,N_13074,N_12466);
or U21323 (N_21323,N_13991,N_12329);
nand U21324 (N_21324,N_12134,N_14087);
and U21325 (N_21325,N_12934,N_17590);
nor U21326 (N_21326,N_17148,N_16740);
and U21327 (N_21327,N_16892,N_17815);
xor U21328 (N_21328,N_13111,N_13580);
nand U21329 (N_21329,N_16610,N_14371);
nor U21330 (N_21330,N_12125,N_15774);
xor U21331 (N_21331,N_13749,N_12376);
xor U21332 (N_21332,N_13216,N_12067);
xor U21333 (N_21333,N_16493,N_17616);
nand U21334 (N_21334,N_12609,N_15317);
and U21335 (N_21335,N_14785,N_17434);
nor U21336 (N_21336,N_14609,N_16570);
or U21337 (N_21337,N_12787,N_13171);
or U21338 (N_21338,N_17777,N_12119);
nand U21339 (N_21339,N_16733,N_16836);
or U21340 (N_21340,N_15314,N_13736);
or U21341 (N_21341,N_12287,N_16656);
nor U21342 (N_21342,N_13349,N_16709);
or U21343 (N_21343,N_17758,N_17932);
xnor U21344 (N_21344,N_15410,N_16261);
and U21345 (N_21345,N_13736,N_17867);
nand U21346 (N_21346,N_16299,N_16899);
or U21347 (N_21347,N_17647,N_16596);
nor U21348 (N_21348,N_14749,N_16032);
nand U21349 (N_21349,N_14347,N_12631);
nor U21350 (N_21350,N_13532,N_16444);
or U21351 (N_21351,N_12072,N_13138);
or U21352 (N_21352,N_12014,N_14522);
or U21353 (N_21353,N_14810,N_13600);
xnor U21354 (N_21354,N_16591,N_14285);
nand U21355 (N_21355,N_17599,N_13911);
or U21356 (N_21356,N_16414,N_15184);
nor U21357 (N_21357,N_17920,N_15199);
nand U21358 (N_21358,N_15680,N_13456);
nand U21359 (N_21359,N_14323,N_13786);
and U21360 (N_21360,N_17406,N_15448);
nor U21361 (N_21361,N_16832,N_15422);
nor U21362 (N_21362,N_12156,N_15161);
xnor U21363 (N_21363,N_12827,N_17656);
nor U21364 (N_21364,N_14867,N_15741);
or U21365 (N_21365,N_14280,N_17274);
nand U21366 (N_21366,N_16681,N_16810);
nor U21367 (N_21367,N_16122,N_13475);
or U21368 (N_21368,N_13489,N_15673);
nor U21369 (N_21369,N_16062,N_15418);
xor U21370 (N_21370,N_12744,N_14568);
xnor U21371 (N_21371,N_16040,N_14309);
nand U21372 (N_21372,N_13429,N_13633);
xor U21373 (N_21373,N_16192,N_12227);
nor U21374 (N_21374,N_15746,N_17885);
or U21375 (N_21375,N_14370,N_14398);
nor U21376 (N_21376,N_17463,N_14476);
xor U21377 (N_21377,N_15831,N_14967);
nand U21378 (N_21378,N_12700,N_14773);
nand U21379 (N_21379,N_14453,N_16906);
or U21380 (N_21380,N_13634,N_12023);
nor U21381 (N_21381,N_16635,N_12684);
xor U21382 (N_21382,N_17216,N_16469);
xnor U21383 (N_21383,N_16884,N_12353);
nor U21384 (N_21384,N_14473,N_13263);
and U21385 (N_21385,N_15526,N_13738);
and U21386 (N_21386,N_13006,N_14788);
or U21387 (N_21387,N_17345,N_17721);
or U21388 (N_21388,N_15749,N_15081);
nand U21389 (N_21389,N_12887,N_12914);
and U21390 (N_21390,N_17626,N_15226);
or U21391 (N_21391,N_14621,N_13227);
nor U21392 (N_21392,N_15714,N_13920);
or U21393 (N_21393,N_15378,N_16299);
and U21394 (N_21394,N_12516,N_14307);
nor U21395 (N_21395,N_12572,N_12493);
xor U21396 (N_21396,N_15870,N_13660);
nor U21397 (N_21397,N_15766,N_17758);
nand U21398 (N_21398,N_15631,N_12613);
xnor U21399 (N_21399,N_14531,N_16843);
and U21400 (N_21400,N_13865,N_16642);
nand U21401 (N_21401,N_13778,N_16229);
and U21402 (N_21402,N_14909,N_14899);
or U21403 (N_21403,N_14777,N_13097);
or U21404 (N_21404,N_15318,N_13617);
nor U21405 (N_21405,N_16861,N_15580);
xor U21406 (N_21406,N_17727,N_15645);
or U21407 (N_21407,N_16960,N_12304);
and U21408 (N_21408,N_17608,N_16173);
nor U21409 (N_21409,N_16771,N_13199);
or U21410 (N_21410,N_14519,N_17247);
or U21411 (N_21411,N_12592,N_14752);
xor U21412 (N_21412,N_16307,N_12896);
xnor U21413 (N_21413,N_13507,N_12967);
nand U21414 (N_21414,N_15643,N_16896);
nor U21415 (N_21415,N_12559,N_16288);
and U21416 (N_21416,N_15412,N_12189);
nor U21417 (N_21417,N_14709,N_13237);
xnor U21418 (N_21418,N_14355,N_13540);
nand U21419 (N_21419,N_16014,N_13181);
xnor U21420 (N_21420,N_16432,N_14917);
and U21421 (N_21421,N_12402,N_13260);
and U21422 (N_21422,N_16538,N_17369);
nand U21423 (N_21423,N_13768,N_13659);
xnor U21424 (N_21424,N_15189,N_16148);
nand U21425 (N_21425,N_12925,N_14660);
xor U21426 (N_21426,N_13743,N_17082);
nor U21427 (N_21427,N_15052,N_16751);
and U21428 (N_21428,N_12214,N_12373);
nor U21429 (N_21429,N_16998,N_13996);
nor U21430 (N_21430,N_12796,N_12933);
nor U21431 (N_21431,N_15867,N_15727);
xnor U21432 (N_21432,N_12984,N_13030);
nand U21433 (N_21433,N_17065,N_12960);
nand U21434 (N_21434,N_13815,N_15868);
nor U21435 (N_21435,N_12996,N_15948);
nand U21436 (N_21436,N_17550,N_13882);
xor U21437 (N_21437,N_12352,N_17969);
or U21438 (N_21438,N_14161,N_17106);
and U21439 (N_21439,N_14000,N_13827);
or U21440 (N_21440,N_16361,N_12629);
xnor U21441 (N_21441,N_17023,N_13424);
nand U21442 (N_21442,N_14842,N_16321);
nand U21443 (N_21443,N_16536,N_15824);
nor U21444 (N_21444,N_16586,N_15324);
nand U21445 (N_21445,N_15315,N_12370);
or U21446 (N_21446,N_17954,N_15258);
or U21447 (N_21447,N_12780,N_13259);
and U21448 (N_21448,N_16918,N_16002);
nor U21449 (N_21449,N_14031,N_14279);
and U21450 (N_21450,N_16455,N_13776);
or U21451 (N_21451,N_15719,N_13796);
nand U21452 (N_21452,N_15982,N_13340);
and U21453 (N_21453,N_13163,N_12824);
xnor U21454 (N_21454,N_14706,N_12849);
xnor U21455 (N_21455,N_12497,N_17318);
and U21456 (N_21456,N_13770,N_17904);
and U21457 (N_21457,N_12035,N_15781);
and U21458 (N_21458,N_17353,N_14766);
and U21459 (N_21459,N_14458,N_16103);
nor U21460 (N_21460,N_14249,N_15387);
or U21461 (N_21461,N_15221,N_17095);
nand U21462 (N_21462,N_12025,N_14657);
and U21463 (N_21463,N_14381,N_16702);
and U21464 (N_21464,N_16071,N_17632);
nand U21465 (N_21465,N_16033,N_12634);
nand U21466 (N_21466,N_16327,N_16578);
nand U21467 (N_21467,N_13935,N_15018);
and U21468 (N_21468,N_16277,N_17679);
nor U21469 (N_21469,N_15004,N_17706);
nor U21470 (N_21470,N_16690,N_12234);
nand U21471 (N_21471,N_12659,N_16280);
or U21472 (N_21472,N_14454,N_12389);
nor U21473 (N_21473,N_16225,N_13765);
and U21474 (N_21474,N_12084,N_12171);
nand U21475 (N_21475,N_16504,N_16900);
or U21476 (N_21476,N_16958,N_14252);
and U21477 (N_21477,N_13330,N_12871);
nand U21478 (N_21478,N_12750,N_14874);
nand U21479 (N_21479,N_15155,N_17456);
or U21480 (N_21480,N_17331,N_12377);
nor U21481 (N_21481,N_17140,N_17854);
and U21482 (N_21482,N_16225,N_16734);
xor U21483 (N_21483,N_12115,N_12320);
and U21484 (N_21484,N_12741,N_13240);
or U21485 (N_21485,N_14003,N_13222);
nor U21486 (N_21486,N_17465,N_13149);
or U21487 (N_21487,N_16209,N_15143);
or U21488 (N_21488,N_13069,N_17673);
or U21489 (N_21489,N_14736,N_14078);
nand U21490 (N_21490,N_12648,N_14140);
and U21491 (N_21491,N_12418,N_16713);
xor U21492 (N_21492,N_17787,N_14371);
and U21493 (N_21493,N_16298,N_13331);
and U21494 (N_21494,N_16192,N_17840);
and U21495 (N_21495,N_15872,N_14180);
or U21496 (N_21496,N_16495,N_17196);
xnor U21497 (N_21497,N_12520,N_14364);
or U21498 (N_21498,N_14005,N_17397);
nor U21499 (N_21499,N_12968,N_12259);
nor U21500 (N_21500,N_12621,N_15007);
xor U21501 (N_21501,N_14529,N_14011);
nor U21502 (N_21502,N_14928,N_15348);
nor U21503 (N_21503,N_12747,N_12599);
or U21504 (N_21504,N_12652,N_13996);
nor U21505 (N_21505,N_15535,N_12843);
or U21506 (N_21506,N_14180,N_15220);
nand U21507 (N_21507,N_16396,N_12749);
xor U21508 (N_21508,N_13040,N_13790);
and U21509 (N_21509,N_14867,N_15434);
xnor U21510 (N_21510,N_15962,N_12162);
or U21511 (N_21511,N_14723,N_12420);
nor U21512 (N_21512,N_15456,N_14876);
xnor U21513 (N_21513,N_14216,N_15903);
xor U21514 (N_21514,N_16534,N_13665);
or U21515 (N_21515,N_13001,N_14438);
nor U21516 (N_21516,N_16753,N_16896);
nor U21517 (N_21517,N_15835,N_15010);
and U21518 (N_21518,N_13964,N_12623);
nand U21519 (N_21519,N_12247,N_13472);
or U21520 (N_21520,N_15336,N_16481);
or U21521 (N_21521,N_14158,N_13159);
or U21522 (N_21522,N_13175,N_15340);
and U21523 (N_21523,N_16849,N_15910);
and U21524 (N_21524,N_15098,N_17098);
or U21525 (N_21525,N_13024,N_13509);
or U21526 (N_21526,N_15314,N_13218);
or U21527 (N_21527,N_16175,N_12662);
or U21528 (N_21528,N_16340,N_16522);
nand U21529 (N_21529,N_13854,N_13201);
and U21530 (N_21530,N_12620,N_13748);
and U21531 (N_21531,N_15889,N_12077);
nand U21532 (N_21532,N_12728,N_15756);
nor U21533 (N_21533,N_15833,N_16304);
nand U21534 (N_21534,N_16791,N_15769);
and U21535 (N_21535,N_16073,N_12111);
or U21536 (N_21536,N_13758,N_17823);
and U21537 (N_21537,N_13918,N_16997);
or U21538 (N_21538,N_16275,N_17437);
or U21539 (N_21539,N_16502,N_12844);
nor U21540 (N_21540,N_12208,N_12154);
nor U21541 (N_21541,N_12494,N_13933);
nor U21542 (N_21542,N_15621,N_14701);
xnor U21543 (N_21543,N_17601,N_13141);
nand U21544 (N_21544,N_12254,N_15687);
and U21545 (N_21545,N_17921,N_15475);
nor U21546 (N_21546,N_13067,N_12848);
nor U21547 (N_21547,N_17645,N_15529);
and U21548 (N_21548,N_14242,N_16792);
nand U21549 (N_21549,N_12740,N_14918);
xor U21550 (N_21550,N_15502,N_15650);
xor U21551 (N_21551,N_15314,N_12782);
xor U21552 (N_21552,N_12303,N_14573);
and U21553 (N_21553,N_15015,N_14996);
or U21554 (N_21554,N_15498,N_14379);
xor U21555 (N_21555,N_12343,N_12473);
xor U21556 (N_21556,N_16397,N_13146);
nand U21557 (N_21557,N_16086,N_15697);
nand U21558 (N_21558,N_16687,N_15504);
nor U21559 (N_21559,N_12134,N_14759);
and U21560 (N_21560,N_14591,N_16652);
nor U21561 (N_21561,N_14252,N_12063);
xor U21562 (N_21562,N_16392,N_17762);
xor U21563 (N_21563,N_12390,N_14947);
nor U21564 (N_21564,N_16574,N_13514);
and U21565 (N_21565,N_17484,N_14121);
nor U21566 (N_21566,N_16541,N_13186);
nand U21567 (N_21567,N_17618,N_16122);
and U21568 (N_21568,N_17531,N_14121);
nor U21569 (N_21569,N_13979,N_17030);
nand U21570 (N_21570,N_14978,N_13320);
nor U21571 (N_21571,N_13931,N_13789);
nor U21572 (N_21572,N_16561,N_16816);
nand U21573 (N_21573,N_14293,N_14839);
or U21574 (N_21574,N_12307,N_12255);
and U21575 (N_21575,N_12004,N_17480);
xnor U21576 (N_21576,N_14251,N_15926);
xnor U21577 (N_21577,N_16996,N_13072);
nor U21578 (N_21578,N_13323,N_13690);
or U21579 (N_21579,N_14123,N_13343);
nor U21580 (N_21580,N_13982,N_13462);
or U21581 (N_21581,N_13673,N_14185);
nor U21582 (N_21582,N_12628,N_14837);
nand U21583 (N_21583,N_17893,N_17053);
and U21584 (N_21584,N_16899,N_14547);
or U21585 (N_21585,N_13281,N_14955);
or U21586 (N_21586,N_13426,N_15965);
nand U21587 (N_21587,N_15174,N_17011);
and U21588 (N_21588,N_16798,N_13235);
xnor U21589 (N_21589,N_13777,N_15182);
and U21590 (N_21590,N_17735,N_14936);
or U21591 (N_21591,N_16288,N_15575);
xnor U21592 (N_21592,N_15390,N_14459);
and U21593 (N_21593,N_12599,N_15901);
and U21594 (N_21594,N_15984,N_13478);
nand U21595 (N_21595,N_12762,N_14031);
and U21596 (N_21596,N_13534,N_16867);
nand U21597 (N_21597,N_16380,N_12024);
nand U21598 (N_21598,N_12490,N_14046);
xnor U21599 (N_21599,N_17391,N_15732);
nand U21600 (N_21600,N_15901,N_12812);
xor U21601 (N_21601,N_14000,N_17666);
nand U21602 (N_21602,N_17257,N_14554);
xnor U21603 (N_21603,N_12774,N_17008);
nand U21604 (N_21604,N_14713,N_14869);
nand U21605 (N_21605,N_14604,N_13218);
and U21606 (N_21606,N_16742,N_17495);
nand U21607 (N_21607,N_16681,N_14123);
and U21608 (N_21608,N_13062,N_14918);
nor U21609 (N_21609,N_17875,N_13859);
nor U21610 (N_21610,N_14790,N_17187);
nand U21611 (N_21611,N_16969,N_13320);
and U21612 (N_21612,N_17475,N_17408);
nand U21613 (N_21613,N_12897,N_15662);
nand U21614 (N_21614,N_13269,N_16869);
nor U21615 (N_21615,N_14932,N_15644);
nor U21616 (N_21616,N_15919,N_16667);
and U21617 (N_21617,N_12748,N_15483);
and U21618 (N_21618,N_12031,N_14028);
nor U21619 (N_21619,N_12718,N_12429);
xnor U21620 (N_21620,N_12038,N_14260);
or U21621 (N_21621,N_15033,N_17565);
or U21622 (N_21622,N_14579,N_14613);
and U21623 (N_21623,N_14583,N_16158);
xor U21624 (N_21624,N_17016,N_12112);
or U21625 (N_21625,N_16267,N_15278);
nand U21626 (N_21626,N_14034,N_13493);
nor U21627 (N_21627,N_15750,N_17681);
nor U21628 (N_21628,N_15630,N_14152);
nor U21629 (N_21629,N_13729,N_14161);
or U21630 (N_21630,N_17786,N_12777);
xor U21631 (N_21631,N_13668,N_14864);
or U21632 (N_21632,N_14561,N_14798);
xor U21633 (N_21633,N_15982,N_15270);
or U21634 (N_21634,N_16756,N_13771);
xnor U21635 (N_21635,N_13273,N_16452);
nor U21636 (N_21636,N_16602,N_12398);
xnor U21637 (N_21637,N_17648,N_16235);
and U21638 (N_21638,N_16235,N_15091);
xor U21639 (N_21639,N_14830,N_16468);
and U21640 (N_21640,N_12541,N_16605);
and U21641 (N_21641,N_15614,N_17159);
xor U21642 (N_21642,N_12050,N_15486);
xnor U21643 (N_21643,N_17801,N_13129);
or U21644 (N_21644,N_13075,N_17388);
and U21645 (N_21645,N_12105,N_17832);
xor U21646 (N_21646,N_13028,N_12211);
or U21647 (N_21647,N_12412,N_13736);
and U21648 (N_21648,N_16796,N_15599);
and U21649 (N_21649,N_12935,N_12239);
nor U21650 (N_21650,N_13630,N_16714);
nand U21651 (N_21651,N_14437,N_15023);
xor U21652 (N_21652,N_14269,N_17569);
nand U21653 (N_21653,N_16266,N_12389);
and U21654 (N_21654,N_12211,N_12384);
or U21655 (N_21655,N_15266,N_16150);
nor U21656 (N_21656,N_16688,N_16214);
xor U21657 (N_21657,N_17303,N_17481);
xor U21658 (N_21658,N_12945,N_16676);
nor U21659 (N_21659,N_17106,N_17820);
xnor U21660 (N_21660,N_13257,N_12918);
nor U21661 (N_21661,N_17813,N_15652);
or U21662 (N_21662,N_14830,N_17937);
nand U21663 (N_21663,N_12359,N_13737);
nand U21664 (N_21664,N_14489,N_16856);
and U21665 (N_21665,N_16937,N_14071);
and U21666 (N_21666,N_12843,N_13587);
and U21667 (N_21667,N_13521,N_16596);
nand U21668 (N_21668,N_17684,N_14530);
or U21669 (N_21669,N_12465,N_15955);
or U21670 (N_21670,N_14099,N_14133);
xnor U21671 (N_21671,N_15857,N_12759);
nor U21672 (N_21672,N_16470,N_15196);
xor U21673 (N_21673,N_16961,N_13103);
nor U21674 (N_21674,N_12916,N_12853);
or U21675 (N_21675,N_14382,N_14154);
xor U21676 (N_21676,N_12701,N_16738);
nor U21677 (N_21677,N_13600,N_15490);
nand U21678 (N_21678,N_16412,N_16469);
or U21679 (N_21679,N_16338,N_14875);
or U21680 (N_21680,N_16263,N_16123);
and U21681 (N_21681,N_15089,N_13811);
nor U21682 (N_21682,N_14155,N_15931);
nand U21683 (N_21683,N_13138,N_17947);
nand U21684 (N_21684,N_16054,N_16944);
nand U21685 (N_21685,N_12951,N_16217);
nor U21686 (N_21686,N_16055,N_14225);
and U21687 (N_21687,N_15622,N_12391);
or U21688 (N_21688,N_13523,N_17078);
nand U21689 (N_21689,N_16959,N_15186);
nand U21690 (N_21690,N_17299,N_17005);
or U21691 (N_21691,N_16370,N_14642);
nor U21692 (N_21692,N_16077,N_15501);
nand U21693 (N_21693,N_16677,N_12562);
nor U21694 (N_21694,N_14097,N_15917);
nand U21695 (N_21695,N_17536,N_16050);
nor U21696 (N_21696,N_13027,N_13544);
and U21697 (N_21697,N_17323,N_17838);
nand U21698 (N_21698,N_16969,N_17607);
or U21699 (N_21699,N_17290,N_13789);
nand U21700 (N_21700,N_14340,N_12655);
nand U21701 (N_21701,N_17763,N_15712);
and U21702 (N_21702,N_13699,N_13238);
or U21703 (N_21703,N_14322,N_14788);
and U21704 (N_21704,N_16625,N_17211);
xnor U21705 (N_21705,N_15375,N_16243);
nand U21706 (N_21706,N_13646,N_16667);
nand U21707 (N_21707,N_16599,N_16825);
or U21708 (N_21708,N_15729,N_13395);
nand U21709 (N_21709,N_17605,N_16723);
or U21710 (N_21710,N_12391,N_15977);
or U21711 (N_21711,N_16615,N_16673);
nor U21712 (N_21712,N_17549,N_17420);
nand U21713 (N_21713,N_15442,N_17256);
xnor U21714 (N_21714,N_14418,N_14588);
and U21715 (N_21715,N_15119,N_12932);
or U21716 (N_21716,N_12746,N_14323);
nor U21717 (N_21717,N_15174,N_14160);
and U21718 (N_21718,N_16693,N_14540);
nor U21719 (N_21719,N_15058,N_16008);
nand U21720 (N_21720,N_17647,N_14195);
nor U21721 (N_21721,N_14458,N_17895);
and U21722 (N_21722,N_17281,N_15393);
nor U21723 (N_21723,N_14639,N_16025);
or U21724 (N_21724,N_12169,N_14199);
nand U21725 (N_21725,N_17944,N_15276);
xor U21726 (N_21726,N_13864,N_16124);
xnor U21727 (N_21727,N_13905,N_15006);
or U21728 (N_21728,N_13035,N_12281);
and U21729 (N_21729,N_17474,N_17908);
and U21730 (N_21730,N_13783,N_14692);
xor U21731 (N_21731,N_16249,N_15147);
and U21732 (N_21732,N_12845,N_12051);
nor U21733 (N_21733,N_17078,N_15806);
nor U21734 (N_21734,N_13939,N_13515);
xor U21735 (N_21735,N_13902,N_16283);
nor U21736 (N_21736,N_16236,N_17188);
or U21737 (N_21737,N_13759,N_14283);
xnor U21738 (N_21738,N_14277,N_16705);
nor U21739 (N_21739,N_13002,N_12258);
or U21740 (N_21740,N_14450,N_15245);
nor U21741 (N_21741,N_15530,N_12871);
nand U21742 (N_21742,N_17579,N_15043);
nand U21743 (N_21743,N_16715,N_13647);
or U21744 (N_21744,N_16043,N_15364);
and U21745 (N_21745,N_15689,N_13185);
nor U21746 (N_21746,N_17473,N_16343);
nor U21747 (N_21747,N_16257,N_15588);
nand U21748 (N_21748,N_14414,N_16454);
and U21749 (N_21749,N_14021,N_15304);
xor U21750 (N_21750,N_15661,N_17719);
xnor U21751 (N_21751,N_17156,N_14181);
xnor U21752 (N_21752,N_16042,N_12606);
xor U21753 (N_21753,N_12759,N_14099);
nor U21754 (N_21754,N_13561,N_16853);
nor U21755 (N_21755,N_17882,N_12957);
nand U21756 (N_21756,N_13225,N_13051);
and U21757 (N_21757,N_15691,N_15578);
nor U21758 (N_21758,N_12068,N_13387);
nor U21759 (N_21759,N_15666,N_15322);
and U21760 (N_21760,N_14341,N_16362);
xor U21761 (N_21761,N_17056,N_16499);
xnor U21762 (N_21762,N_12466,N_13529);
xnor U21763 (N_21763,N_12722,N_14997);
xor U21764 (N_21764,N_13103,N_14519);
and U21765 (N_21765,N_12893,N_17469);
and U21766 (N_21766,N_15579,N_13951);
nor U21767 (N_21767,N_13891,N_16291);
xor U21768 (N_21768,N_14459,N_13783);
or U21769 (N_21769,N_13493,N_12026);
nor U21770 (N_21770,N_15957,N_13444);
xor U21771 (N_21771,N_13164,N_16437);
xor U21772 (N_21772,N_14730,N_14678);
nor U21773 (N_21773,N_12549,N_16163);
nor U21774 (N_21774,N_16358,N_13533);
nor U21775 (N_21775,N_17934,N_16759);
nor U21776 (N_21776,N_14059,N_14572);
and U21777 (N_21777,N_15953,N_15217);
xnor U21778 (N_21778,N_16452,N_14634);
or U21779 (N_21779,N_13627,N_17585);
nand U21780 (N_21780,N_15759,N_15050);
or U21781 (N_21781,N_12581,N_14385);
and U21782 (N_21782,N_12968,N_17590);
nor U21783 (N_21783,N_15894,N_12640);
nand U21784 (N_21784,N_15675,N_16904);
xnor U21785 (N_21785,N_17500,N_15179);
nor U21786 (N_21786,N_16994,N_15508);
nor U21787 (N_21787,N_16868,N_14811);
nor U21788 (N_21788,N_13522,N_15633);
nor U21789 (N_21789,N_14301,N_13501);
xor U21790 (N_21790,N_16960,N_14022);
and U21791 (N_21791,N_14107,N_12774);
nor U21792 (N_21792,N_12800,N_16278);
nor U21793 (N_21793,N_15006,N_16755);
xnor U21794 (N_21794,N_17813,N_16932);
nor U21795 (N_21795,N_13926,N_17846);
and U21796 (N_21796,N_12578,N_15616);
and U21797 (N_21797,N_13737,N_16686);
and U21798 (N_21798,N_14934,N_13015);
xor U21799 (N_21799,N_13895,N_14246);
and U21800 (N_21800,N_16315,N_12621);
xor U21801 (N_21801,N_15609,N_16544);
nand U21802 (N_21802,N_17485,N_16305);
nor U21803 (N_21803,N_14401,N_17908);
or U21804 (N_21804,N_13806,N_16294);
nor U21805 (N_21805,N_17215,N_17903);
and U21806 (N_21806,N_15269,N_12173);
and U21807 (N_21807,N_13714,N_17706);
nand U21808 (N_21808,N_13529,N_12882);
xor U21809 (N_21809,N_12580,N_16401);
xnor U21810 (N_21810,N_14550,N_16573);
xor U21811 (N_21811,N_14172,N_13925);
and U21812 (N_21812,N_12069,N_15245);
nor U21813 (N_21813,N_15423,N_12393);
nand U21814 (N_21814,N_17225,N_17448);
and U21815 (N_21815,N_13413,N_16383);
and U21816 (N_21816,N_17026,N_14877);
nor U21817 (N_21817,N_17843,N_15313);
and U21818 (N_21818,N_15258,N_17771);
and U21819 (N_21819,N_16121,N_16905);
xnor U21820 (N_21820,N_12903,N_15776);
xor U21821 (N_21821,N_16761,N_15421);
nand U21822 (N_21822,N_13532,N_17480);
or U21823 (N_21823,N_15518,N_15922);
and U21824 (N_21824,N_17482,N_12835);
or U21825 (N_21825,N_12456,N_17966);
or U21826 (N_21826,N_16340,N_13017);
nand U21827 (N_21827,N_15229,N_17953);
or U21828 (N_21828,N_16635,N_14105);
nor U21829 (N_21829,N_13993,N_15640);
and U21830 (N_21830,N_12239,N_12211);
nor U21831 (N_21831,N_12309,N_16322);
and U21832 (N_21832,N_16670,N_16552);
or U21833 (N_21833,N_17497,N_12554);
xnor U21834 (N_21834,N_14313,N_16967);
xor U21835 (N_21835,N_16187,N_12561);
nand U21836 (N_21836,N_12994,N_15957);
nand U21837 (N_21837,N_12712,N_12975);
or U21838 (N_21838,N_14304,N_14798);
and U21839 (N_21839,N_16519,N_14412);
or U21840 (N_21840,N_12024,N_12974);
xor U21841 (N_21841,N_14578,N_12562);
xor U21842 (N_21842,N_17079,N_15270);
nand U21843 (N_21843,N_13469,N_13662);
nand U21844 (N_21844,N_13488,N_12587);
nor U21845 (N_21845,N_17387,N_15644);
nor U21846 (N_21846,N_13848,N_15103);
nor U21847 (N_21847,N_14170,N_13173);
and U21848 (N_21848,N_17839,N_17091);
xor U21849 (N_21849,N_13942,N_13406);
or U21850 (N_21850,N_13992,N_17145);
nor U21851 (N_21851,N_17622,N_17185);
nand U21852 (N_21852,N_17026,N_16063);
nand U21853 (N_21853,N_17644,N_14509);
nor U21854 (N_21854,N_16548,N_17723);
xnor U21855 (N_21855,N_14331,N_17072);
xor U21856 (N_21856,N_14274,N_16687);
xor U21857 (N_21857,N_16839,N_13896);
nand U21858 (N_21858,N_16132,N_14160);
nand U21859 (N_21859,N_17011,N_16915);
xor U21860 (N_21860,N_12536,N_12899);
nor U21861 (N_21861,N_15508,N_12266);
xnor U21862 (N_21862,N_13968,N_13811);
nand U21863 (N_21863,N_15117,N_13186);
nor U21864 (N_21864,N_17633,N_15654);
xnor U21865 (N_21865,N_14055,N_16077);
xor U21866 (N_21866,N_14981,N_13181);
xnor U21867 (N_21867,N_15582,N_15172);
or U21868 (N_21868,N_17471,N_14777);
xnor U21869 (N_21869,N_14987,N_14024);
xnor U21870 (N_21870,N_13487,N_14517);
xor U21871 (N_21871,N_15437,N_17641);
and U21872 (N_21872,N_12740,N_15765);
and U21873 (N_21873,N_17990,N_16796);
or U21874 (N_21874,N_16777,N_15243);
nor U21875 (N_21875,N_16546,N_14601);
xor U21876 (N_21876,N_12321,N_14886);
and U21877 (N_21877,N_12346,N_13128);
nand U21878 (N_21878,N_13501,N_17359);
nor U21879 (N_21879,N_16299,N_13284);
or U21880 (N_21880,N_15056,N_14738);
nand U21881 (N_21881,N_12278,N_15971);
nand U21882 (N_21882,N_17724,N_12607);
xor U21883 (N_21883,N_13909,N_12392);
or U21884 (N_21884,N_12691,N_15425);
nand U21885 (N_21885,N_15673,N_14405);
or U21886 (N_21886,N_17741,N_17812);
or U21887 (N_21887,N_17481,N_17652);
nand U21888 (N_21888,N_16798,N_13551);
nand U21889 (N_21889,N_16636,N_17433);
and U21890 (N_21890,N_12155,N_15811);
and U21891 (N_21891,N_17283,N_12493);
nand U21892 (N_21892,N_14897,N_16632);
and U21893 (N_21893,N_17002,N_14665);
xnor U21894 (N_21894,N_12422,N_13807);
or U21895 (N_21895,N_16499,N_15916);
nand U21896 (N_21896,N_17768,N_12899);
nand U21897 (N_21897,N_12808,N_16251);
nand U21898 (N_21898,N_13422,N_17927);
nor U21899 (N_21899,N_13266,N_14176);
nand U21900 (N_21900,N_13596,N_17405);
xor U21901 (N_21901,N_13118,N_14253);
xor U21902 (N_21902,N_16949,N_13402);
nor U21903 (N_21903,N_15810,N_16540);
xor U21904 (N_21904,N_16008,N_13990);
xnor U21905 (N_21905,N_17392,N_15385);
and U21906 (N_21906,N_15543,N_14207);
and U21907 (N_21907,N_16900,N_16919);
and U21908 (N_21908,N_15811,N_13545);
xnor U21909 (N_21909,N_14440,N_17115);
xnor U21910 (N_21910,N_13252,N_14546);
nor U21911 (N_21911,N_13493,N_13599);
and U21912 (N_21912,N_14284,N_14384);
nand U21913 (N_21913,N_17137,N_13317);
nor U21914 (N_21914,N_16567,N_12981);
nor U21915 (N_21915,N_14094,N_13589);
nand U21916 (N_21916,N_12072,N_15288);
nor U21917 (N_21917,N_12144,N_17127);
nor U21918 (N_21918,N_17830,N_14894);
and U21919 (N_21919,N_15532,N_13464);
xnor U21920 (N_21920,N_14015,N_14702);
nand U21921 (N_21921,N_14606,N_14880);
or U21922 (N_21922,N_14759,N_13364);
and U21923 (N_21923,N_17147,N_12942);
or U21924 (N_21924,N_12915,N_14435);
or U21925 (N_21925,N_12983,N_12363);
nor U21926 (N_21926,N_14780,N_13075);
and U21927 (N_21927,N_16547,N_15338);
and U21928 (N_21928,N_17610,N_15193);
nand U21929 (N_21929,N_12733,N_17705);
nand U21930 (N_21930,N_17712,N_13688);
and U21931 (N_21931,N_16925,N_14761);
and U21932 (N_21932,N_14500,N_13510);
or U21933 (N_21933,N_16974,N_15905);
and U21934 (N_21934,N_16302,N_12874);
xor U21935 (N_21935,N_14966,N_14126);
or U21936 (N_21936,N_12458,N_15252);
or U21937 (N_21937,N_17393,N_13751);
nand U21938 (N_21938,N_16777,N_15265);
xnor U21939 (N_21939,N_16375,N_13069);
or U21940 (N_21940,N_15343,N_14163);
or U21941 (N_21941,N_14398,N_14692);
xor U21942 (N_21942,N_15776,N_12485);
nand U21943 (N_21943,N_14693,N_12255);
nand U21944 (N_21944,N_16427,N_13653);
and U21945 (N_21945,N_16696,N_15976);
nor U21946 (N_21946,N_12137,N_17449);
or U21947 (N_21947,N_12163,N_14788);
nand U21948 (N_21948,N_13006,N_12372);
nor U21949 (N_21949,N_17666,N_12833);
nor U21950 (N_21950,N_14624,N_13474);
or U21951 (N_21951,N_14568,N_13394);
nor U21952 (N_21952,N_13857,N_17084);
or U21953 (N_21953,N_16506,N_14559);
nor U21954 (N_21954,N_16818,N_12830);
nor U21955 (N_21955,N_12783,N_16740);
nor U21956 (N_21956,N_13974,N_16728);
or U21957 (N_21957,N_12809,N_12913);
nor U21958 (N_21958,N_13030,N_14034);
nand U21959 (N_21959,N_14205,N_14837);
nand U21960 (N_21960,N_15440,N_17009);
nand U21961 (N_21961,N_14924,N_17752);
and U21962 (N_21962,N_17176,N_14907);
xnor U21963 (N_21963,N_17043,N_12005);
nor U21964 (N_21964,N_15758,N_17141);
or U21965 (N_21965,N_12778,N_13215);
nand U21966 (N_21966,N_12515,N_12192);
xnor U21967 (N_21967,N_15009,N_14059);
xnor U21968 (N_21968,N_17188,N_12407);
or U21969 (N_21969,N_13840,N_13468);
and U21970 (N_21970,N_15154,N_15368);
xor U21971 (N_21971,N_16855,N_16985);
xnor U21972 (N_21972,N_13333,N_16746);
or U21973 (N_21973,N_13765,N_13205);
xnor U21974 (N_21974,N_15999,N_15894);
nor U21975 (N_21975,N_15637,N_14926);
and U21976 (N_21976,N_15725,N_15139);
and U21977 (N_21977,N_13079,N_13427);
nand U21978 (N_21978,N_16607,N_16202);
or U21979 (N_21979,N_16380,N_15231);
nand U21980 (N_21980,N_14687,N_16688);
nand U21981 (N_21981,N_12188,N_15967);
and U21982 (N_21982,N_17594,N_15942);
nor U21983 (N_21983,N_15794,N_16985);
nand U21984 (N_21984,N_16586,N_14543);
xnor U21985 (N_21985,N_15857,N_14580);
and U21986 (N_21986,N_14514,N_14334);
nor U21987 (N_21987,N_13216,N_13627);
nand U21988 (N_21988,N_16990,N_16775);
or U21989 (N_21989,N_15477,N_13117);
xnor U21990 (N_21990,N_17909,N_12052);
nor U21991 (N_21991,N_12288,N_14661);
xor U21992 (N_21992,N_17742,N_16015);
nand U21993 (N_21993,N_15577,N_15092);
and U21994 (N_21994,N_17984,N_17484);
and U21995 (N_21995,N_15385,N_17070);
nand U21996 (N_21996,N_14578,N_16870);
nor U21997 (N_21997,N_16630,N_13996);
nor U21998 (N_21998,N_16222,N_16366);
and U21999 (N_21999,N_12231,N_17250);
xnor U22000 (N_22000,N_17402,N_14059);
nand U22001 (N_22001,N_15566,N_16960);
and U22002 (N_22002,N_17357,N_15009);
or U22003 (N_22003,N_15870,N_16028);
and U22004 (N_22004,N_15195,N_16506);
and U22005 (N_22005,N_17702,N_14817);
xnor U22006 (N_22006,N_17944,N_12741);
or U22007 (N_22007,N_12479,N_16703);
nand U22008 (N_22008,N_16878,N_14516);
xor U22009 (N_22009,N_12198,N_12330);
and U22010 (N_22010,N_17292,N_13624);
and U22011 (N_22011,N_12546,N_12206);
or U22012 (N_22012,N_17470,N_12945);
nand U22013 (N_22013,N_13514,N_16140);
and U22014 (N_22014,N_14875,N_14190);
nand U22015 (N_22015,N_13294,N_17525);
or U22016 (N_22016,N_14110,N_14104);
nor U22017 (N_22017,N_14702,N_13586);
xor U22018 (N_22018,N_16118,N_13577);
xor U22019 (N_22019,N_13888,N_16839);
and U22020 (N_22020,N_14622,N_13173);
nand U22021 (N_22021,N_15409,N_14507);
and U22022 (N_22022,N_14538,N_16649);
nand U22023 (N_22023,N_17852,N_16453);
nor U22024 (N_22024,N_12476,N_17092);
or U22025 (N_22025,N_12025,N_12945);
nand U22026 (N_22026,N_16418,N_16899);
or U22027 (N_22027,N_16571,N_16493);
xnor U22028 (N_22028,N_13949,N_17980);
xor U22029 (N_22029,N_16380,N_17735);
or U22030 (N_22030,N_14596,N_16670);
and U22031 (N_22031,N_12656,N_12829);
xnor U22032 (N_22032,N_15300,N_15181);
or U22033 (N_22033,N_14592,N_14513);
or U22034 (N_22034,N_15104,N_16458);
xor U22035 (N_22035,N_15277,N_17954);
nand U22036 (N_22036,N_13889,N_14167);
nand U22037 (N_22037,N_12577,N_16752);
nor U22038 (N_22038,N_14974,N_15119);
nor U22039 (N_22039,N_13913,N_12906);
nor U22040 (N_22040,N_17492,N_12445);
nand U22041 (N_22041,N_13796,N_14182);
and U22042 (N_22042,N_13181,N_12659);
or U22043 (N_22043,N_13048,N_12896);
xnor U22044 (N_22044,N_13385,N_12913);
xor U22045 (N_22045,N_16434,N_12207);
xnor U22046 (N_22046,N_16899,N_14308);
and U22047 (N_22047,N_12155,N_13291);
nor U22048 (N_22048,N_17507,N_15573);
nor U22049 (N_22049,N_12961,N_17042);
and U22050 (N_22050,N_13178,N_16798);
nor U22051 (N_22051,N_16846,N_15621);
or U22052 (N_22052,N_12036,N_14755);
nor U22053 (N_22053,N_17436,N_13641);
nor U22054 (N_22054,N_13582,N_17805);
nor U22055 (N_22055,N_16635,N_14945);
nand U22056 (N_22056,N_14164,N_17439);
or U22057 (N_22057,N_13192,N_12206);
nor U22058 (N_22058,N_12962,N_16861);
and U22059 (N_22059,N_12372,N_16761);
xnor U22060 (N_22060,N_12362,N_17400);
and U22061 (N_22061,N_13825,N_14830);
and U22062 (N_22062,N_12138,N_14762);
nor U22063 (N_22063,N_17853,N_12980);
nand U22064 (N_22064,N_16677,N_12347);
nand U22065 (N_22065,N_14962,N_12066);
nor U22066 (N_22066,N_15143,N_12771);
or U22067 (N_22067,N_12217,N_17624);
nand U22068 (N_22068,N_13633,N_15732);
xor U22069 (N_22069,N_16443,N_15319);
xnor U22070 (N_22070,N_14535,N_14315);
nor U22071 (N_22071,N_15503,N_14609);
nand U22072 (N_22072,N_17593,N_12799);
nor U22073 (N_22073,N_14793,N_14910);
or U22074 (N_22074,N_17884,N_14500);
xor U22075 (N_22075,N_13556,N_14308);
or U22076 (N_22076,N_12437,N_16591);
or U22077 (N_22077,N_15728,N_12986);
xor U22078 (N_22078,N_15721,N_16623);
xor U22079 (N_22079,N_16747,N_16779);
nor U22080 (N_22080,N_14613,N_17802);
xor U22081 (N_22081,N_16603,N_17565);
nor U22082 (N_22082,N_17065,N_13139);
or U22083 (N_22083,N_16655,N_17831);
xor U22084 (N_22084,N_14876,N_12585);
and U22085 (N_22085,N_16613,N_16328);
nor U22086 (N_22086,N_15140,N_16135);
and U22087 (N_22087,N_13689,N_12908);
and U22088 (N_22088,N_16545,N_14984);
nor U22089 (N_22089,N_17469,N_17913);
nand U22090 (N_22090,N_14017,N_12806);
and U22091 (N_22091,N_15754,N_17057);
nand U22092 (N_22092,N_17458,N_13475);
or U22093 (N_22093,N_13232,N_13803);
and U22094 (N_22094,N_17750,N_12486);
nor U22095 (N_22095,N_13255,N_15409);
nor U22096 (N_22096,N_13163,N_14722);
nand U22097 (N_22097,N_14027,N_17063);
or U22098 (N_22098,N_13977,N_15452);
or U22099 (N_22099,N_14184,N_16808);
xnor U22100 (N_22100,N_12692,N_17646);
nand U22101 (N_22101,N_13464,N_12880);
nand U22102 (N_22102,N_16410,N_17977);
or U22103 (N_22103,N_13681,N_15788);
and U22104 (N_22104,N_14862,N_13456);
or U22105 (N_22105,N_16505,N_16199);
nor U22106 (N_22106,N_13039,N_15337);
nand U22107 (N_22107,N_16655,N_12911);
nand U22108 (N_22108,N_14205,N_15496);
nand U22109 (N_22109,N_17890,N_13774);
nand U22110 (N_22110,N_15511,N_15832);
and U22111 (N_22111,N_13278,N_15798);
nand U22112 (N_22112,N_14818,N_16423);
nand U22113 (N_22113,N_16929,N_16857);
xnor U22114 (N_22114,N_13099,N_12584);
and U22115 (N_22115,N_13483,N_17980);
nor U22116 (N_22116,N_15176,N_16183);
and U22117 (N_22117,N_12006,N_14039);
nor U22118 (N_22118,N_12426,N_14139);
or U22119 (N_22119,N_16583,N_12528);
and U22120 (N_22120,N_12342,N_13717);
nand U22121 (N_22121,N_12222,N_13608);
nor U22122 (N_22122,N_14946,N_12153);
nand U22123 (N_22123,N_12815,N_17512);
nand U22124 (N_22124,N_12820,N_13115);
and U22125 (N_22125,N_17520,N_16672);
nand U22126 (N_22126,N_15099,N_15129);
nand U22127 (N_22127,N_14116,N_14253);
or U22128 (N_22128,N_13203,N_13795);
or U22129 (N_22129,N_14131,N_15745);
nand U22130 (N_22130,N_14786,N_16945);
xnor U22131 (N_22131,N_14244,N_13521);
and U22132 (N_22132,N_17903,N_12689);
xnor U22133 (N_22133,N_16160,N_12648);
nand U22134 (N_22134,N_14703,N_15499);
or U22135 (N_22135,N_17425,N_15719);
nor U22136 (N_22136,N_16292,N_12989);
or U22137 (N_22137,N_16013,N_12848);
or U22138 (N_22138,N_14304,N_14620);
nand U22139 (N_22139,N_13271,N_12308);
or U22140 (N_22140,N_13149,N_12390);
nand U22141 (N_22141,N_16572,N_15688);
or U22142 (N_22142,N_17546,N_14045);
xor U22143 (N_22143,N_16663,N_12891);
nand U22144 (N_22144,N_12006,N_14535);
and U22145 (N_22145,N_14655,N_16578);
nor U22146 (N_22146,N_15110,N_15194);
xor U22147 (N_22147,N_14818,N_15170);
nor U22148 (N_22148,N_15116,N_14864);
nor U22149 (N_22149,N_12581,N_16554);
xor U22150 (N_22150,N_13471,N_17839);
nor U22151 (N_22151,N_14918,N_13965);
or U22152 (N_22152,N_17884,N_14416);
or U22153 (N_22153,N_16411,N_16040);
and U22154 (N_22154,N_12038,N_15643);
or U22155 (N_22155,N_16443,N_16029);
or U22156 (N_22156,N_17381,N_14803);
nand U22157 (N_22157,N_17398,N_12818);
or U22158 (N_22158,N_13008,N_17048);
nand U22159 (N_22159,N_12691,N_17599);
nor U22160 (N_22160,N_12046,N_13701);
and U22161 (N_22161,N_14163,N_13519);
nand U22162 (N_22162,N_16882,N_17426);
or U22163 (N_22163,N_16049,N_13506);
or U22164 (N_22164,N_15254,N_12353);
and U22165 (N_22165,N_13717,N_14956);
nand U22166 (N_22166,N_16242,N_16192);
or U22167 (N_22167,N_15040,N_15542);
nand U22168 (N_22168,N_14739,N_17609);
nand U22169 (N_22169,N_13404,N_13326);
nand U22170 (N_22170,N_12268,N_15404);
nand U22171 (N_22171,N_14257,N_17679);
xnor U22172 (N_22172,N_13634,N_17601);
nor U22173 (N_22173,N_16902,N_15802);
nor U22174 (N_22174,N_14881,N_12552);
nand U22175 (N_22175,N_13131,N_16412);
or U22176 (N_22176,N_17826,N_14728);
xnor U22177 (N_22177,N_13421,N_15539);
xor U22178 (N_22178,N_12366,N_15108);
nor U22179 (N_22179,N_15757,N_14239);
xnor U22180 (N_22180,N_16105,N_12716);
xnor U22181 (N_22181,N_14873,N_14633);
nand U22182 (N_22182,N_12823,N_15393);
or U22183 (N_22183,N_12939,N_16557);
nor U22184 (N_22184,N_13708,N_14357);
nand U22185 (N_22185,N_17048,N_13536);
xnor U22186 (N_22186,N_17774,N_15850);
or U22187 (N_22187,N_14641,N_12249);
or U22188 (N_22188,N_12163,N_15681);
nand U22189 (N_22189,N_16723,N_16478);
or U22190 (N_22190,N_17124,N_16168);
nor U22191 (N_22191,N_17203,N_14291);
nand U22192 (N_22192,N_16035,N_14549);
nand U22193 (N_22193,N_12544,N_17465);
or U22194 (N_22194,N_16161,N_16926);
nand U22195 (N_22195,N_16146,N_17467);
nor U22196 (N_22196,N_13710,N_13418);
xnor U22197 (N_22197,N_15627,N_12191);
and U22198 (N_22198,N_15379,N_16424);
or U22199 (N_22199,N_16910,N_16056);
nand U22200 (N_22200,N_17113,N_12006);
nand U22201 (N_22201,N_17978,N_13971);
or U22202 (N_22202,N_13928,N_12612);
xnor U22203 (N_22203,N_14181,N_17914);
or U22204 (N_22204,N_17934,N_14010);
nor U22205 (N_22205,N_13179,N_12957);
xnor U22206 (N_22206,N_15410,N_12171);
and U22207 (N_22207,N_15706,N_15728);
nor U22208 (N_22208,N_14515,N_13991);
nand U22209 (N_22209,N_15896,N_13307);
and U22210 (N_22210,N_13789,N_14655);
or U22211 (N_22211,N_17107,N_12687);
and U22212 (N_22212,N_15557,N_14754);
xor U22213 (N_22213,N_14952,N_13525);
xnor U22214 (N_22214,N_15988,N_13066);
xnor U22215 (N_22215,N_16660,N_13397);
xnor U22216 (N_22216,N_14780,N_16061);
and U22217 (N_22217,N_16608,N_12921);
xnor U22218 (N_22218,N_15374,N_16826);
and U22219 (N_22219,N_15302,N_13156);
nor U22220 (N_22220,N_12407,N_14974);
and U22221 (N_22221,N_12642,N_15618);
nand U22222 (N_22222,N_12630,N_13386);
and U22223 (N_22223,N_13693,N_12515);
nor U22224 (N_22224,N_15859,N_16461);
nand U22225 (N_22225,N_15382,N_13188);
nand U22226 (N_22226,N_13816,N_15352);
and U22227 (N_22227,N_17368,N_17161);
and U22228 (N_22228,N_15390,N_16461);
and U22229 (N_22229,N_15503,N_12853);
and U22230 (N_22230,N_16841,N_16806);
or U22231 (N_22231,N_12695,N_12374);
and U22232 (N_22232,N_16132,N_17912);
nor U22233 (N_22233,N_17831,N_15142);
nand U22234 (N_22234,N_16876,N_13070);
and U22235 (N_22235,N_15204,N_16622);
or U22236 (N_22236,N_12400,N_17150);
and U22237 (N_22237,N_17408,N_17448);
or U22238 (N_22238,N_16236,N_14251);
or U22239 (N_22239,N_16912,N_12546);
and U22240 (N_22240,N_14518,N_16684);
nor U22241 (N_22241,N_15987,N_16304);
or U22242 (N_22242,N_14534,N_16425);
nand U22243 (N_22243,N_17064,N_16263);
nor U22244 (N_22244,N_17209,N_16727);
nor U22245 (N_22245,N_15969,N_17304);
or U22246 (N_22246,N_17081,N_16284);
or U22247 (N_22247,N_14186,N_12284);
nand U22248 (N_22248,N_16486,N_15500);
and U22249 (N_22249,N_14590,N_13904);
nor U22250 (N_22250,N_14177,N_15236);
xor U22251 (N_22251,N_15230,N_16880);
xnor U22252 (N_22252,N_14706,N_16886);
nor U22253 (N_22253,N_14884,N_16290);
or U22254 (N_22254,N_14496,N_17691);
xor U22255 (N_22255,N_12113,N_12391);
nor U22256 (N_22256,N_15184,N_16698);
nand U22257 (N_22257,N_16790,N_13838);
and U22258 (N_22258,N_15819,N_12501);
nand U22259 (N_22259,N_14006,N_13735);
and U22260 (N_22260,N_13171,N_14382);
nor U22261 (N_22261,N_12287,N_17326);
and U22262 (N_22262,N_15512,N_13477);
and U22263 (N_22263,N_16071,N_17638);
nor U22264 (N_22264,N_17681,N_16684);
or U22265 (N_22265,N_15096,N_15928);
nor U22266 (N_22266,N_15409,N_12240);
and U22267 (N_22267,N_15401,N_15769);
or U22268 (N_22268,N_13056,N_13522);
or U22269 (N_22269,N_12166,N_12041);
nor U22270 (N_22270,N_17770,N_15241);
nor U22271 (N_22271,N_13536,N_14586);
nand U22272 (N_22272,N_15314,N_13800);
and U22273 (N_22273,N_16490,N_17764);
and U22274 (N_22274,N_12009,N_13978);
and U22275 (N_22275,N_15000,N_14577);
and U22276 (N_22276,N_14115,N_12892);
or U22277 (N_22277,N_17521,N_12983);
or U22278 (N_22278,N_15711,N_16595);
nand U22279 (N_22279,N_15990,N_14271);
nand U22280 (N_22280,N_13506,N_14747);
xor U22281 (N_22281,N_13971,N_17422);
and U22282 (N_22282,N_14392,N_17396);
xnor U22283 (N_22283,N_16620,N_17365);
nand U22284 (N_22284,N_14137,N_12297);
or U22285 (N_22285,N_12989,N_15059);
and U22286 (N_22286,N_13532,N_14613);
and U22287 (N_22287,N_16886,N_13788);
nand U22288 (N_22288,N_13296,N_15954);
or U22289 (N_22289,N_16692,N_12967);
or U22290 (N_22290,N_16859,N_16929);
nand U22291 (N_22291,N_12728,N_15013);
nand U22292 (N_22292,N_15807,N_15137);
nor U22293 (N_22293,N_12753,N_12705);
and U22294 (N_22294,N_17215,N_16428);
xnor U22295 (N_22295,N_16695,N_17866);
nor U22296 (N_22296,N_15001,N_14304);
nand U22297 (N_22297,N_12929,N_13166);
xnor U22298 (N_22298,N_14688,N_17787);
nand U22299 (N_22299,N_13933,N_17327);
nor U22300 (N_22300,N_15022,N_14483);
or U22301 (N_22301,N_16299,N_17006);
xor U22302 (N_22302,N_17066,N_12900);
and U22303 (N_22303,N_13000,N_17374);
nor U22304 (N_22304,N_14901,N_12327);
or U22305 (N_22305,N_12181,N_13924);
and U22306 (N_22306,N_13996,N_12897);
nor U22307 (N_22307,N_17231,N_13795);
xnor U22308 (N_22308,N_15534,N_17383);
or U22309 (N_22309,N_17394,N_15497);
nand U22310 (N_22310,N_15582,N_15885);
nand U22311 (N_22311,N_13250,N_13715);
and U22312 (N_22312,N_17898,N_14063);
or U22313 (N_22313,N_12056,N_15888);
and U22314 (N_22314,N_15281,N_16539);
nor U22315 (N_22315,N_17161,N_12701);
or U22316 (N_22316,N_17456,N_15539);
or U22317 (N_22317,N_12318,N_14625);
nand U22318 (N_22318,N_12091,N_12156);
and U22319 (N_22319,N_13096,N_17071);
and U22320 (N_22320,N_17457,N_12333);
and U22321 (N_22321,N_16733,N_15876);
and U22322 (N_22322,N_13861,N_15177);
and U22323 (N_22323,N_16313,N_14925);
or U22324 (N_22324,N_15604,N_16502);
or U22325 (N_22325,N_14981,N_16075);
nor U22326 (N_22326,N_12674,N_17981);
xnor U22327 (N_22327,N_17671,N_15480);
nand U22328 (N_22328,N_16692,N_14920);
nor U22329 (N_22329,N_12329,N_16869);
or U22330 (N_22330,N_13162,N_14305);
nor U22331 (N_22331,N_15430,N_14025);
or U22332 (N_22332,N_16750,N_13724);
nand U22333 (N_22333,N_14443,N_14258);
xor U22334 (N_22334,N_15755,N_17806);
nand U22335 (N_22335,N_13009,N_16569);
or U22336 (N_22336,N_12348,N_17600);
or U22337 (N_22337,N_16163,N_12522);
nand U22338 (N_22338,N_13192,N_17721);
and U22339 (N_22339,N_16010,N_14360);
nand U22340 (N_22340,N_14597,N_17690);
or U22341 (N_22341,N_17067,N_14531);
and U22342 (N_22342,N_15228,N_12744);
nor U22343 (N_22343,N_16193,N_12766);
or U22344 (N_22344,N_17232,N_12495);
xnor U22345 (N_22345,N_12952,N_17555);
xnor U22346 (N_22346,N_13024,N_13028);
nand U22347 (N_22347,N_14907,N_14727);
nor U22348 (N_22348,N_15907,N_16708);
or U22349 (N_22349,N_13760,N_15592);
nor U22350 (N_22350,N_14287,N_14074);
nand U22351 (N_22351,N_13157,N_14277);
nand U22352 (N_22352,N_12518,N_14249);
or U22353 (N_22353,N_15089,N_16239);
or U22354 (N_22354,N_12567,N_14777);
nor U22355 (N_22355,N_13877,N_17979);
nand U22356 (N_22356,N_12121,N_17347);
xnor U22357 (N_22357,N_12880,N_16917);
nand U22358 (N_22358,N_16404,N_12737);
or U22359 (N_22359,N_17158,N_15439);
and U22360 (N_22360,N_17828,N_16399);
xor U22361 (N_22361,N_15801,N_15102);
nor U22362 (N_22362,N_12155,N_17680);
and U22363 (N_22363,N_14272,N_12606);
or U22364 (N_22364,N_14787,N_13365);
nand U22365 (N_22365,N_15213,N_13693);
nand U22366 (N_22366,N_16482,N_17364);
or U22367 (N_22367,N_13979,N_16902);
and U22368 (N_22368,N_17061,N_12216);
and U22369 (N_22369,N_12798,N_12961);
or U22370 (N_22370,N_13571,N_15116);
or U22371 (N_22371,N_16169,N_15766);
nand U22372 (N_22372,N_16141,N_12674);
or U22373 (N_22373,N_15379,N_12939);
nand U22374 (N_22374,N_14514,N_17104);
xor U22375 (N_22375,N_17262,N_16819);
xnor U22376 (N_22376,N_13120,N_14625);
and U22377 (N_22377,N_12112,N_17045);
nand U22378 (N_22378,N_15200,N_14354);
and U22379 (N_22379,N_12682,N_15121);
or U22380 (N_22380,N_15531,N_13716);
nor U22381 (N_22381,N_13504,N_12254);
or U22382 (N_22382,N_16801,N_16951);
xor U22383 (N_22383,N_16621,N_13160);
nand U22384 (N_22384,N_13246,N_15457);
nand U22385 (N_22385,N_16848,N_15976);
or U22386 (N_22386,N_13901,N_17370);
xor U22387 (N_22387,N_16339,N_15185);
nor U22388 (N_22388,N_17172,N_15209);
xnor U22389 (N_22389,N_16955,N_13505);
or U22390 (N_22390,N_17392,N_13345);
nor U22391 (N_22391,N_17670,N_17102);
or U22392 (N_22392,N_17379,N_16441);
nand U22393 (N_22393,N_14446,N_16443);
nand U22394 (N_22394,N_16679,N_13668);
nor U22395 (N_22395,N_13196,N_14417);
nand U22396 (N_22396,N_16365,N_14896);
nand U22397 (N_22397,N_12619,N_17189);
nor U22398 (N_22398,N_16013,N_12856);
and U22399 (N_22399,N_13723,N_13060);
nand U22400 (N_22400,N_12530,N_12348);
nor U22401 (N_22401,N_17829,N_15484);
and U22402 (N_22402,N_16233,N_16985);
xor U22403 (N_22403,N_14064,N_13108);
or U22404 (N_22404,N_17223,N_12160);
nand U22405 (N_22405,N_17813,N_16701);
xnor U22406 (N_22406,N_16352,N_15049);
and U22407 (N_22407,N_15683,N_14450);
or U22408 (N_22408,N_16251,N_17547);
or U22409 (N_22409,N_13606,N_12046);
xor U22410 (N_22410,N_13309,N_14652);
and U22411 (N_22411,N_14081,N_15678);
and U22412 (N_22412,N_13785,N_15993);
xnor U22413 (N_22413,N_16227,N_14369);
nand U22414 (N_22414,N_15813,N_12242);
and U22415 (N_22415,N_14884,N_16700);
or U22416 (N_22416,N_17191,N_13266);
xnor U22417 (N_22417,N_17812,N_17928);
or U22418 (N_22418,N_12095,N_14683);
nand U22419 (N_22419,N_12459,N_17800);
and U22420 (N_22420,N_13161,N_14445);
and U22421 (N_22421,N_15214,N_13661);
and U22422 (N_22422,N_13960,N_12558);
or U22423 (N_22423,N_16521,N_17859);
nand U22424 (N_22424,N_17544,N_12053);
and U22425 (N_22425,N_14083,N_15929);
nor U22426 (N_22426,N_17562,N_13637);
nor U22427 (N_22427,N_15083,N_15931);
or U22428 (N_22428,N_13060,N_12966);
nand U22429 (N_22429,N_12360,N_13030);
nor U22430 (N_22430,N_14462,N_14161);
and U22431 (N_22431,N_15804,N_13816);
nand U22432 (N_22432,N_14802,N_14521);
and U22433 (N_22433,N_15198,N_12308);
and U22434 (N_22434,N_15816,N_13908);
xor U22435 (N_22435,N_13133,N_13085);
or U22436 (N_22436,N_15301,N_12028);
and U22437 (N_22437,N_12902,N_14020);
and U22438 (N_22438,N_17399,N_13930);
and U22439 (N_22439,N_15742,N_13102);
xnor U22440 (N_22440,N_12914,N_16547);
and U22441 (N_22441,N_17891,N_13992);
xor U22442 (N_22442,N_16958,N_14947);
and U22443 (N_22443,N_16529,N_14698);
xor U22444 (N_22444,N_13484,N_13260);
or U22445 (N_22445,N_14196,N_13422);
xnor U22446 (N_22446,N_14687,N_15597);
xnor U22447 (N_22447,N_17568,N_12453);
nand U22448 (N_22448,N_17828,N_13667);
xnor U22449 (N_22449,N_17312,N_14985);
and U22450 (N_22450,N_16634,N_12563);
xnor U22451 (N_22451,N_17565,N_13950);
and U22452 (N_22452,N_13902,N_14331);
or U22453 (N_22453,N_14540,N_12849);
nand U22454 (N_22454,N_13843,N_13588);
and U22455 (N_22455,N_12444,N_13446);
nand U22456 (N_22456,N_16811,N_14220);
or U22457 (N_22457,N_12560,N_13035);
xor U22458 (N_22458,N_16030,N_15217);
xnor U22459 (N_22459,N_15202,N_14406);
xnor U22460 (N_22460,N_16429,N_12448);
xnor U22461 (N_22461,N_16385,N_13553);
or U22462 (N_22462,N_16809,N_12649);
nand U22463 (N_22463,N_16251,N_12888);
or U22464 (N_22464,N_13376,N_15749);
xnor U22465 (N_22465,N_13924,N_17742);
nor U22466 (N_22466,N_16416,N_17260);
and U22467 (N_22467,N_15400,N_12183);
or U22468 (N_22468,N_12924,N_17283);
nand U22469 (N_22469,N_12061,N_14113);
nor U22470 (N_22470,N_12556,N_15572);
and U22471 (N_22471,N_14553,N_17983);
xor U22472 (N_22472,N_15014,N_14027);
nor U22473 (N_22473,N_15432,N_16054);
nand U22474 (N_22474,N_14557,N_17719);
nand U22475 (N_22475,N_14047,N_17224);
and U22476 (N_22476,N_17891,N_13622);
nand U22477 (N_22477,N_13769,N_17284);
or U22478 (N_22478,N_12927,N_13641);
xnor U22479 (N_22479,N_14599,N_12985);
nand U22480 (N_22480,N_12187,N_16432);
nand U22481 (N_22481,N_14295,N_14638);
or U22482 (N_22482,N_16987,N_13196);
nand U22483 (N_22483,N_16670,N_12021);
nor U22484 (N_22484,N_15625,N_12147);
or U22485 (N_22485,N_15667,N_15620);
or U22486 (N_22486,N_14036,N_16289);
and U22487 (N_22487,N_14808,N_14079);
nand U22488 (N_22488,N_17666,N_17779);
nand U22489 (N_22489,N_16518,N_13342);
and U22490 (N_22490,N_14591,N_13277);
and U22491 (N_22491,N_13999,N_17594);
nor U22492 (N_22492,N_14921,N_14629);
nor U22493 (N_22493,N_16253,N_14210);
nand U22494 (N_22494,N_16544,N_13726);
xnor U22495 (N_22495,N_13692,N_16210);
and U22496 (N_22496,N_12534,N_13508);
nand U22497 (N_22497,N_13917,N_16858);
xnor U22498 (N_22498,N_16887,N_13112);
xor U22499 (N_22499,N_16087,N_15369);
xnor U22500 (N_22500,N_17120,N_14462);
and U22501 (N_22501,N_13485,N_14555);
and U22502 (N_22502,N_15156,N_14699);
xnor U22503 (N_22503,N_12539,N_15862);
and U22504 (N_22504,N_15216,N_15234);
nand U22505 (N_22505,N_17128,N_12751);
xnor U22506 (N_22506,N_16425,N_12704);
xor U22507 (N_22507,N_14032,N_16504);
nor U22508 (N_22508,N_17991,N_15727);
xor U22509 (N_22509,N_15222,N_16328);
nor U22510 (N_22510,N_16447,N_13708);
nor U22511 (N_22511,N_16075,N_15763);
nand U22512 (N_22512,N_14429,N_13001);
and U22513 (N_22513,N_16767,N_13465);
nand U22514 (N_22514,N_17953,N_13721);
and U22515 (N_22515,N_15664,N_13262);
and U22516 (N_22516,N_14039,N_16959);
and U22517 (N_22517,N_17403,N_12411);
or U22518 (N_22518,N_16596,N_14464);
and U22519 (N_22519,N_15620,N_15884);
nand U22520 (N_22520,N_14075,N_17884);
nor U22521 (N_22521,N_14040,N_14807);
nand U22522 (N_22522,N_14139,N_17533);
nor U22523 (N_22523,N_14720,N_13372);
nand U22524 (N_22524,N_15270,N_17199);
nand U22525 (N_22525,N_16789,N_12919);
nor U22526 (N_22526,N_16841,N_15601);
nor U22527 (N_22527,N_15948,N_17606);
and U22528 (N_22528,N_17020,N_12201);
and U22529 (N_22529,N_14126,N_17065);
or U22530 (N_22530,N_12250,N_17874);
and U22531 (N_22531,N_16942,N_14238);
nor U22532 (N_22532,N_14649,N_14808);
and U22533 (N_22533,N_16812,N_13493);
and U22534 (N_22534,N_14578,N_15307);
nor U22535 (N_22535,N_17405,N_14428);
xor U22536 (N_22536,N_14601,N_16352);
nand U22537 (N_22537,N_16359,N_14265);
xor U22538 (N_22538,N_13038,N_15047);
nor U22539 (N_22539,N_12649,N_15998);
xnor U22540 (N_22540,N_12477,N_13578);
or U22541 (N_22541,N_17073,N_17228);
and U22542 (N_22542,N_16158,N_17366);
nor U22543 (N_22543,N_16662,N_16114);
or U22544 (N_22544,N_15267,N_16435);
nand U22545 (N_22545,N_17073,N_15051);
or U22546 (N_22546,N_12453,N_17675);
nor U22547 (N_22547,N_14206,N_14165);
nor U22548 (N_22548,N_13256,N_16919);
xor U22549 (N_22549,N_17573,N_15312);
nand U22550 (N_22550,N_15882,N_17301);
nor U22551 (N_22551,N_14083,N_16664);
nand U22552 (N_22552,N_16014,N_16490);
nor U22553 (N_22553,N_15333,N_17538);
nor U22554 (N_22554,N_12232,N_13039);
xor U22555 (N_22555,N_12019,N_14197);
xnor U22556 (N_22556,N_14406,N_14401);
and U22557 (N_22557,N_17715,N_13756);
xor U22558 (N_22558,N_13932,N_13781);
and U22559 (N_22559,N_14703,N_12615);
xnor U22560 (N_22560,N_14120,N_12677);
and U22561 (N_22561,N_15961,N_14126);
xor U22562 (N_22562,N_12659,N_12347);
nand U22563 (N_22563,N_13277,N_14053);
xor U22564 (N_22564,N_14872,N_12816);
or U22565 (N_22565,N_16881,N_13282);
and U22566 (N_22566,N_13608,N_12692);
xnor U22567 (N_22567,N_12210,N_12031);
nor U22568 (N_22568,N_16215,N_16778);
and U22569 (N_22569,N_12750,N_17993);
and U22570 (N_22570,N_14873,N_13594);
or U22571 (N_22571,N_17170,N_13392);
nand U22572 (N_22572,N_12256,N_14027);
or U22573 (N_22573,N_17732,N_14034);
nand U22574 (N_22574,N_16640,N_15633);
or U22575 (N_22575,N_17116,N_15210);
nor U22576 (N_22576,N_15547,N_12576);
and U22577 (N_22577,N_17410,N_15215);
and U22578 (N_22578,N_17460,N_17456);
nor U22579 (N_22579,N_16009,N_14625);
nor U22580 (N_22580,N_17524,N_13209);
xnor U22581 (N_22581,N_15999,N_17420);
and U22582 (N_22582,N_17911,N_14637);
and U22583 (N_22583,N_14494,N_12774);
nor U22584 (N_22584,N_17853,N_15899);
xor U22585 (N_22585,N_12666,N_14577);
or U22586 (N_22586,N_14757,N_13645);
nor U22587 (N_22587,N_14676,N_13873);
xor U22588 (N_22588,N_12325,N_13905);
or U22589 (N_22589,N_13111,N_14139);
nor U22590 (N_22590,N_13819,N_13830);
xor U22591 (N_22591,N_13180,N_13557);
and U22592 (N_22592,N_13522,N_15211);
xor U22593 (N_22593,N_13384,N_13939);
xor U22594 (N_22594,N_17860,N_13067);
xor U22595 (N_22595,N_12894,N_13521);
or U22596 (N_22596,N_13644,N_15307);
or U22597 (N_22597,N_12182,N_12551);
nand U22598 (N_22598,N_17599,N_13092);
or U22599 (N_22599,N_17309,N_12777);
or U22600 (N_22600,N_13674,N_17627);
nor U22601 (N_22601,N_17273,N_13073);
nand U22602 (N_22602,N_14145,N_15115);
and U22603 (N_22603,N_12688,N_14476);
nor U22604 (N_22604,N_13397,N_13497);
nor U22605 (N_22605,N_14914,N_12229);
nor U22606 (N_22606,N_14253,N_13677);
nor U22607 (N_22607,N_12790,N_17406);
nand U22608 (N_22608,N_17367,N_12325);
nor U22609 (N_22609,N_14427,N_17243);
or U22610 (N_22610,N_17204,N_14236);
or U22611 (N_22611,N_12995,N_14684);
nor U22612 (N_22612,N_17925,N_13682);
and U22613 (N_22613,N_14816,N_16352);
and U22614 (N_22614,N_15329,N_13446);
and U22615 (N_22615,N_16662,N_15153);
and U22616 (N_22616,N_13473,N_17573);
nand U22617 (N_22617,N_13954,N_14500);
nand U22618 (N_22618,N_17196,N_12679);
and U22619 (N_22619,N_14849,N_12042);
and U22620 (N_22620,N_15328,N_17978);
nand U22621 (N_22621,N_12670,N_15402);
nand U22622 (N_22622,N_14783,N_15249);
xnor U22623 (N_22623,N_12928,N_16902);
xor U22624 (N_22624,N_12253,N_17472);
nor U22625 (N_22625,N_17829,N_15146);
or U22626 (N_22626,N_15821,N_16543);
and U22627 (N_22627,N_14682,N_13600);
nor U22628 (N_22628,N_17961,N_17052);
nor U22629 (N_22629,N_16839,N_17377);
and U22630 (N_22630,N_16791,N_17986);
and U22631 (N_22631,N_15584,N_12478);
nor U22632 (N_22632,N_12191,N_15170);
xor U22633 (N_22633,N_16730,N_15918);
nor U22634 (N_22634,N_14368,N_15462);
nand U22635 (N_22635,N_12217,N_16794);
and U22636 (N_22636,N_12251,N_13623);
or U22637 (N_22637,N_13509,N_17951);
nor U22638 (N_22638,N_13671,N_12462);
xnor U22639 (N_22639,N_12350,N_16981);
nor U22640 (N_22640,N_17164,N_14754);
xnor U22641 (N_22641,N_13550,N_12011);
and U22642 (N_22642,N_12049,N_12524);
xnor U22643 (N_22643,N_13714,N_16579);
and U22644 (N_22644,N_16618,N_12712);
nor U22645 (N_22645,N_14609,N_17401);
nand U22646 (N_22646,N_15237,N_17305);
and U22647 (N_22647,N_15433,N_15355);
nand U22648 (N_22648,N_13478,N_15259);
nor U22649 (N_22649,N_17762,N_15524);
or U22650 (N_22650,N_14098,N_14705);
and U22651 (N_22651,N_15738,N_15606);
or U22652 (N_22652,N_13133,N_17077);
and U22653 (N_22653,N_13912,N_17630);
nor U22654 (N_22654,N_12645,N_17066);
or U22655 (N_22655,N_12217,N_13187);
nor U22656 (N_22656,N_16418,N_13569);
or U22657 (N_22657,N_16853,N_13428);
nor U22658 (N_22658,N_12195,N_13464);
xnor U22659 (N_22659,N_16112,N_14417);
or U22660 (N_22660,N_13283,N_16250);
xor U22661 (N_22661,N_16514,N_12053);
and U22662 (N_22662,N_15656,N_12725);
and U22663 (N_22663,N_12937,N_14128);
nand U22664 (N_22664,N_14577,N_15947);
or U22665 (N_22665,N_15067,N_14932);
nor U22666 (N_22666,N_15904,N_15378);
nand U22667 (N_22667,N_14775,N_16271);
or U22668 (N_22668,N_12872,N_12452);
and U22669 (N_22669,N_13641,N_15091);
nor U22670 (N_22670,N_15297,N_14351);
or U22671 (N_22671,N_16277,N_12410);
nor U22672 (N_22672,N_15334,N_15518);
xnor U22673 (N_22673,N_13683,N_16934);
xnor U22674 (N_22674,N_14460,N_12528);
xnor U22675 (N_22675,N_12655,N_12813);
or U22676 (N_22676,N_13855,N_14968);
or U22677 (N_22677,N_13723,N_14783);
nand U22678 (N_22678,N_12957,N_17720);
nor U22679 (N_22679,N_14163,N_13600);
or U22680 (N_22680,N_14021,N_16820);
nand U22681 (N_22681,N_13022,N_16833);
or U22682 (N_22682,N_17251,N_17776);
or U22683 (N_22683,N_14635,N_14697);
xor U22684 (N_22684,N_12554,N_14114);
nand U22685 (N_22685,N_14096,N_14310);
nand U22686 (N_22686,N_12908,N_14166);
nand U22687 (N_22687,N_14547,N_16260);
xor U22688 (N_22688,N_13925,N_16537);
nand U22689 (N_22689,N_16135,N_12425);
and U22690 (N_22690,N_16273,N_16593);
or U22691 (N_22691,N_17672,N_16957);
nor U22692 (N_22692,N_15104,N_17827);
xnor U22693 (N_22693,N_13222,N_17344);
and U22694 (N_22694,N_13729,N_14467);
and U22695 (N_22695,N_13477,N_14706);
and U22696 (N_22696,N_14353,N_17982);
xor U22697 (N_22697,N_14663,N_17160);
xor U22698 (N_22698,N_15433,N_17496);
and U22699 (N_22699,N_17274,N_17408);
xnor U22700 (N_22700,N_13401,N_17924);
nor U22701 (N_22701,N_17169,N_13446);
nor U22702 (N_22702,N_16716,N_13378);
nand U22703 (N_22703,N_14883,N_12785);
nand U22704 (N_22704,N_14127,N_12379);
nand U22705 (N_22705,N_15554,N_14244);
xor U22706 (N_22706,N_12518,N_14497);
nor U22707 (N_22707,N_14994,N_16504);
nor U22708 (N_22708,N_13098,N_15353);
nor U22709 (N_22709,N_16245,N_13488);
nand U22710 (N_22710,N_16422,N_16839);
xnor U22711 (N_22711,N_12562,N_15036);
and U22712 (N_22712,N_15815,N_14653);
and U22713 (N_22713,N_15808,N_15841);
xnor U22714 (N_22714,N_12072,N_14860);
xor U22715 (N_22715,N_14383,N_16215);
nand U22716 (N_22716,N_15422,N_12499);
nor U22717 (N_22717,N_16785,N_16833);
nand U22718 (N_22718,N_15149,N_13042);
xnor U22719 (N_22719,N_14131,N_12436);
nand U22720 (N_22720,N_14888,N_13964);
nor U22721 (N_22721,N_14615,N_13959);
nand U22722 (N_22722,N_17798,N_16516);
or U22723 (N_22723,N_13103,N_16824);
and U22724 (N_22724,N_17596,N_16145);
xor U22725 (N_22725,N_15709,N_12274);
and U22726 (N_22726,N_14356,N_12685);
or U22727 (N_22727,N_15632,N_12287);
or U22728 (N_22728,N_17241,N_13010);
or U22729 (N_22729,N_14641,N_12471);
or U22730 (N_22730,N_13714,N_13106);
or U22731 (N_22731,N_12624,N_16615);
nor U22732 (N_22732,N_16600,N_12447);
nor U22733 (N_22733,N_13799,N_16889);
and U22734 (N_22734,N_17480,N_13634);
or U22735 (N_22735,N_13803,N_12335);
xnor U22736 (N_22736,N_16454,N_14020);
nand U22737 (N_22737,N_12842,N_13325);
and U22738 (N_22738,N_17070,N_16006);
and U22739 (N_22739,N_12166,N_15505);
or U22740 (N_22740,N_14078,N_13517);
nor U22741 (N_22741,N_15618,N_13746);
and U22742 (N_22742,N_14669,N_17310);
or U22743 (N_22743,N_13227,N_15032);
xnor U22744 (N_22744,N_13617,N_14471);
or U22745 (N_22745,N_15452,N_15345);
nor U22746 (N_22746,N_15832,N_14374);
nor U22747 (N_22747,N_13458,N_13529);
xnor U22748 (N_22748,N_13622,N_16712);
nor U22749 (N_22749,N_15229,N_14730);
or U22750 (N_22750,N_16670,N_14594);
nor U22751 (N_22751,N_12486,N_15626);
and U22752 (N_22752,N_14904,N_14348);
xor U22753 (N_22753,N_17553,N_17763);
xor U22754 (N_22754,N_15523,N_17076);
nor U22755 (N_22755,N_16194,N_12183);
and U22756 (N_22756,N_17461,N_16904);
xnor U22757 (N_22757,N_13882,N_13893);
xnor U22758 (N_22758,N_17616,N_12933);
xnor U22759 (N_22759,N_12025,N_14720);
xnor U22760 (N_22760,N_15397,N_15607);
nand U22761 (N_22761,N_17374,N_14759);
nand U22762 (N_22762,N_15760,N_17167);
xor U22763 (N_22763,N_14413,N_16517);
or U22764 (N_22764,N_16037,N_15277);
xor U22765 (N_22765,N_14483,N_17919);
nor U22766 (N_22766,N_13103,N_16840);
nand U22767 (N_22767,N_13187,N_15128);
or U22768 (N_22768,N_13195,N_14689);
nor U22769 (N_22769,N_16982,N_12981);
nor U22770 (N_22770,N_16822,N_16550);
xor U22771 (N_22771,N_13294,N_17916);
or U22772 (N_22772,N_13967,N_15877);
nor U22773 (N_22773,N_12363,N_13080);
and U22774 (N_22774,N_16747,N_16475);
and U22775 (N_22775,N_17756,N_13424);
or U22776 (N_22776,N_12218,N_14381);
nor U22777 (N_22777,N_17779,N_12526);
and U22778 (N_22778,N_13496,N_15517);
and U22779 (N_22779,N_14616,N_12789);
nand U22780 (N_22780,N_13010,N_12928);
nor U22781 (N_22781,N_16885,N_16746);
and U22782 (N_22782,N_16094,N_17299);
nand U22783 (N_22783,N_15547,N_16776);
nand U22784 (N_22784,N_17362,N_15847);
and U22785 (N_22785,N_15764,N_13999);
nand U22786 (N_22786,N_15058,N_16277);
nand U22787 (N_22787,N_12512,N_17636);
or U22788 (N_22788,N_16771,N_15564);
xnor U22789 (N_22789,N_16615,N_12512);
or U22790 (N_22790,N_12098,N_12324);
xnor U22791 (N_22791,N_17890,N_15330);
nor U22792 (N_22792,N_13044,N_12041);
nor U22793 (N_22793,N_17982,N_14030);
and U22794 (N_22794,N_17972,N_17527);
xor U22795 (N_22795,N_17253,N_13571);
xnor U22796 (N_22796,N_12427,N_15810);
nand U22797 (N_22797,N_17063,N_13134);
nand U22798 (N_22798,N_15535,N_14715);
nor U22799 (N_22799,N_16464,N_14605);
xnor U22800 (N_22800,N_15139,N_17699);
or U22801 (N_22801,N_13486,N_12933);
nor U22802 (N_22802,N_14387,N_17975);
or U22803 (N_22803,N_13903,N_14861);
and U22804 (N_22804,N_14745,N_12397);
and U22805 (N_22805,N_16097,N_16531);
and U22806 (N_22806,N_12284,N_17306);
or U22807 (N_22807,N_17888,N_16855);
and U22808 (N_22808,N_16678,N_15839);
or U22809 (N_22809,N_15057,N_12144);
or U22810 (N_22810,N_17074,N_15430);
nand U22811 (N_22811,N_13558,N_17332);
nand U22812 (N_22812,N_15490,N_14035);
nand U22813 (N_22813,N_12934,N_12958);
nor U22814 (N_22814,N_14780,N_12461);
and U22815 (N_22815,N_15813,N_13457);
nor U22816 (N_22816,N_14494,N_13933);
nand U22817 (N_22817,N_15619,N_17739);
xnor U22818 (N_22818,N_15556,N_14882);
nand U22819 (N_22819,N_14106,N_12678);
nor U22820 (N_22820,N_12787,N_17534);
and U22821 (N_22821,N_17830,N_14758);
nand U22822 (N_22822,N_17268,N_14390);
and U22823 (N_22823,N_17580,N_16567);
nand U22824 (N_22824,N_13939,N_13473);
and U22825 (N_22825,N_13562,N_12514);
nand U22826 (N_22826,N_17921,N_17522);
xnor U22827 (N_22827,N_13994,N_16956);
nand U22828 (N_22828,N_16613,N_14972);
nor U22829 (N_22829,N_14570,N_15123);
nor U22830 (N_22830,N_13628,N_17871);
nand U22831 (N_22831,N_17229,N_14162);
xnor U22832 (N_22832,N_16882,N_13376);
nand U22833 (N_22833,N_12611,N_17427);
nand U22834 (N_22834,N_16117,N_15706);
nand U22835 (N_22835,N_17819,N_15716);
nor U22836 (N_22836,N_15971,N_16021);
xor U22837 (N_22837,N_17363,N_12603);
xor U22838 (N_22838,N_12984,N_15030);
and U22839 (N_22839,N_16191,N_13352);
and U22840 (N_22840,N_12387,N_13826);
xnor U22841 (N_22841,N_12803,N_13970);
nor U22842 (N_22842,N_13346,N_17227);
nand U22843 (N_22843,N_13960,N_14781);
nor U22844 (N_22844,N_16982,N_13578);
or U22845 (N_22845,N_16401,N_12420);
nor U22846 (N_22846,N_14543,N_16304);
and U22847 (N_22847,N_12076,N_12429);
nand U22848 (N_22848,N_13144,N_17307);
and U22849 (N_22849,N_16104,N_15894);
xor U22850 (N_22850,N_12933,N_14267);
xnor U22851 (N_22851,N_16519,N_17937);
or U22852 (N_22852,N_15000,N_16312);
nor U22853 (N_22853,N_14380,N_17118);
nor U22854 (N_22854,N_17373,N_15817);
or U22855 (N_22855,N_15929,N_14790);
nand U22856 (N_22856,N_13945,N_17299);
or U22857 (N_22857,N_15786,N_17217);
nor U22858 (N_22858,N_17545,N_14082);
xor U22859 (N_22859,N_15635,N_13534);
xor U22860 (N_22860,N_17185,N_17034);
nand U22861 (N_22861,N_14155,N_14536);
or U22862 (N_22862,N_17599,N_16177);
or U22863 (N_22863,N_17050,N_12078);
and U22864 (N_22864,N_15769,N_17107);
and U22865 (N_22865,N_14209,N_15677);
nand U22866 (N_22866,N_17774,N_15684);
and U22867 (N_22867,N_17070,N_15644);
nand U22868 (N_22868,N_13722,N_17034);
and U22869 (N_22869,N_14409,N_16203);
or U22870 (N_22870,N_17050,N_14999);
or U22871 (N_22871,N_15257,N_13729);
xnor U22872 (N_22872,N_13631,N_12112);
nor U22873 (N_22873,N_17395,N_12270);
nand U22874 (N_22874,N_14676,N_12055);
nor U22875 (N_22875,N_16128,N_16902);
and U22876 (N_22876,N_14399,N_16429);
xnor U22877 (N_22877,N_12649,N_13668);
nor U22878 (N_22878,N_13065,N_14474);
nor U22879 (N_22879,N_17788,N_17104);
or U22880 (N_22880,N_14390,N_17062);
nand U22881 (N_22881,N_13580,N_16865);
xnor U22882 (N_22882,N_17191,N_15603);
nor U22883 (N_22883,N_12592,N_16965);
or U22884 (N_22884,N_16385,N_17597);
and U22885 (N_22885,N_15828,N_13473);
nor U22886 (N_22886,N_16681,N_14137);
xor U22887 (N_22887,N_14932,N_14130);
xor U22888 (N_22888,N_12490,N_17176);
or U22889 (N_22889,N_12477,N_16956);
nand U22890 (N_22890,N_16039,N_16146);
and U22891 (N_22891,N_17941,N_17665);
nand U22892 (N_22892,N_14119,N_16518);
or U22893 (N_22893,N_13642,N_16146);
nand U22894 (N_22894,N_14514,N_16269);
nand U22895 (N_22895,N_15371,N_12113);
or U22896 (N_22896,N_12059,N_16334);
and U22897 (N_22897,N_15195,N_14618);
nor U22898 (N_22898,N_14295,N_12600);
and U22899 (N_22899,N_12141,N_12919);
nand U22900 (N_22900,N_13866,N_16549);
nand U22901 (N_22901,N_16462,N_17291);
nor U22902 (N_22902,N_12798,N_16174);
nand U22903 (N_22903,N_12582,N_12122);
or U22904 (N_22904,N_15161,N_17710);
nor U22905 (N_22905,N_16954,N_17935);
nor U22906 (N_22906,N_15225,N_17425);
nand U22907 (N_22907,N_13306,N_17082);
xor U22908 (N_22908,N_14282,N_12286);
or U22909 (N_22909,N_15438,N_16652);
xor U22910 (N_22910,N_17418,N_17796);
nand U22911 (N_22911,N_16581,N_17788);
or U22912 (N_22912,N_16556,N_15723);
or U22913 (N_22913,N_16261,N_16619);
nand U22914 (N_22914,N_17414,N_12238);
nand U22915 (N_22915,N_13379,N_15432);
xnor U22916 (N_22916,N_14332,N_12442);
and U22917 (N_22917,N_12826,N_13959);
or U22918 (N_22918,N_12843,N_17299);
nor U22919 (N_22919,N_15564,N_16847);
xnor U22920 (N_22920,N_14495,N_12527);
nor U22921 (N_22921,N_15133,N_17407);
nor U22922 (N_22922,N_13572,N_17678);
nand U22923 (N_22923,N_12385,N_15750);
nand U22924 (N_22924,N_13375,N_15862);
or U22925 (N_22925,N_15761,N_12260);
xor U22926 (N_22926,N_15894,N_16616);
nand U22927 (N_22927,N_14296,N_14331);
nor U22928 (N_22928,N_17985,N_12031);
or U22929 (N_22929,N_13172,N_12650);
nand U22930 (N_22930,N_14901,N_13538);
or U22931 (N_22931,N_14141,N_16625);
nand U22932 (N_22932,N_15337,N_16687);
xor U22933 (N_22933,N_14253,N_16202);
and U22934 (N_22934,N_16288,N_15076);
or U22935 (N_22935,N_13312,N_13126);
nor U22936 (N_22936,N_17191,N_16932);
xor U22937 (N_22937,N_14026,N_14334);
nor U22938 (N_22938,N_16066,N_17366);
xnor U22939 (N_22939,N_13932,N_17138);
xor U22940 (N_22940,N_16201,N_17293);
or U22941 (N_22941,N_15546,N_14614);
xor U22942 (N_22942,N_13315,N_17973);
nand U22943 (N_22943,N_16364,N_15320);
nor U22944 (N_22944,N_16563,N_15589);
and U22945 (N_22945,N_16265,N_12065);
nor U22946 (N_22946,N_15396,N_14167);
nand U22947 (N_22947,N_13814,N_16907);
and U22948 (N_22948,N_17491,N_14607);
nor U22949 (N_22949,N_15178,N_12618);
nor U22950 (N_22950,N_14976,N_15119);
or U22951 (N_22951,N_16353,N_13318);
xnor U22952 (N_22952,N_12389,N_17572);
or U22953 (N_22953,N_17562,N_17713);
xor U22954 (N_22954,N_17438,N_17879);
or U22955 (N_22955,N_14511,N_14217);
nor U22956 (N_22956,N_12130,N_17957);
xor U22957 (N_22957,N_16017,N_16256);
and U22958 (N_22958,N_16039,N_16119);
xnor U22959 (N_22959,N_13156,N_17160);
nor U22960 (N_22960,N_16722,N_13828);
or U22961 (N_22961,N_13834,N_16023);
and U22962 (N_22962,N_16822,N_13176);
nand U22963 (N_22963,N_17004,N_12800);
nand U22964 (N_22964,N_13177,N_13157);
xnor U22965 (N_22965,N_16291,N_12000);
or U22966 (N_22966,N_16652,N_17084);
and U22967 (N_22967,N_15788,N_12385);
nor U22968 (N_22968,N_12346,N_15847);
or U22969 (N_22969,N_14484,N_16230);
nand U22970 (N_22970,N_17810,N_13557);
or U22971 (N_22971,N_13035,N_13239);
nor U22972 (N_22972,N_16561,N_14202);
or U22973 (N_22973,N_16391,N_15133);
xor U22974 (N_22974,N_16686,N_12583);
nor U22975 (N_22975,N_14506,N_17120);
and U22976 (N_22976,N_12105,N_14739);
nor U22977 (N_22977,N_15711,N_16904);
xor U22978 (N_22978,N_13957,N_17765);
nand U22979 (N_22979,N_13451,N_13409);
nor U22980 (N_22980,N_13692,N_16674);
nor U22981 (N_22981,N_12849,N_12872);
nand U22982 (N_22982,N_13394,N_17647);
or U22983 (N_22983,N_15432,N_17665);
and U22984 (N_22984,N_17855,N_12925);
nand U22985 (N_22985,N_17263,N_13408);
nand U22986 (N_22986,N_15062,N_13691);
nor U22987 (N_22987,N_14707,N_14782);
or U22988 (N_22988,N_17097,N_15304);
and U22989 (N_22989,N_17444,N_16952);
or U22990 (N_22990,N_13458,N_12820);
xnor U22991 (N_22991,N_14662,N_12179);
nand U22992 (N_22992,N_15576,N_15859);
or U22993 (N_22993,N_15508,N_15361);
and U22994 (N_22994,N_17935,N_14192);
nand U22995 (N_22995,N_16491,N_17645);
xor U22996 (N_22996,N_13102,N_12861);
nor U22997 (N_22997,N_15091,N_14608);
and U22998 (N_22998,N_14076,N_13437);
and U22999 (N_22999,N_16789,N_14218);
and U23000 (N_23000,N_16539,N_14375);
and U23001 (N_23001,N_15595,N_14313);
nor U23002 (N_23002,N_16647,N_12543);
xor U23003 (N_23003,N_15775,N_12516);
nor U23004 (N_23004,N_15255,N_13239);
xnor U23005 (N_23005,N_14960,N_16469);
nor U23006 (N_23006,N_15965,N_13609);
xnor U23007 (N_23007,N_17787,N_14350);
nor U23008 (N_23008,N_14410,N_15706);
nand U23009 (N_23009,N_13302,N_16410);
or U23010 (N_23010,N_12666,N_14363);
or U23011 (N_23011,N_12427,N_14727);
nor U23012 (N_23012,N_14047,N_13535);
xor U23013 (N_23013,N_12599,N_16944);
nor U23014 (N_23014,N_12679,N_16992);
nor U23015 (N_23015,N_16605,N_14105);
nor U23016 (N_23016,N_13983,N_12596);
xor U23017 (N_23017,N_14800,N_14137);
xnor U23018 (N_23018,N_13306,N_14319);
and U23019 (N_23019,N_15102,N_15478);
nand U23020 (N_23020,N_16330,N_13589);
and U23021 (N_23021,N_17278,N_15981);
and U23022 (N_23022,N_13066,N_12367);
or U23023 (N_23023,N_16092,N_14145);
or U23024 (N_23024,N_14773,N_12704);
nor U23025 (N_23025,N_16777,N_16275);
or U23026 (N_23026,N_16923,N_17929);
and U23027 (N_23027,N_15493,N_17440);
xor U23028 (N_23028,N_12866,N_13012);
or U23029 (N_23029,N_17676,N_16436);
and U23030 (N_23030,N_16561,N_14047);
nor U23031 (N_23031,N_14644,N_14761);
or U23032 (N_23032,N_15886,N_16138);
and U23033 (N_23033,N_13062,N_14957);
and U23034 (N_23034,N_16712,N_15452);
and U23035 (N_23035,N_15607,N_15971);
or U23036 (N_23036,N_17157,N_15893);
nand U23037 (N_23037,N_12876,N_12453);
and U23038 (N_23038,N_17057,N_13814);
nor U23039 (N_23039,N_17611,N_14621);
nand U23040 (N_23040,N_12399,N_12193);
and U23041 (N_23041,N_13450,N_15553);
nor U23042 (N_23042,N_14323,N_12333);
or U23043 (N_23043,N_16404,N_15561);
xor U23044 (N_23044,N_13886,N_14820);
and U23045 (N_23045,N_15238,N_16042);
nand U23046 (N_23046,N_17258,N_17522);
nand U23047 (N_23047,N_15410,N_12554);
xor U23048 (N_23048,N_16184,N_17485);
nand U23049 (N_23049,N_15741,N_14408);
and U23050 (N_23050,N_15551,N_13432);
and U23051 (N_23051,N_14156,N_13646);
and U23052 (N_23052,N_16932,N_17918);
and U23053 (N_23053,N_12896,N_16610);
and U23054 (N_23054,N_14538,N_14691);
and U23055 (N_23055,N_15394,N_15223);
nand U23056 (N_23056,N_15508,N_15405);
nor U23057 (N_23057,N_12770,N_17399);
xnor U23058 (N_23058,N_12982,N_16831);
nor U23059 (N_23059,N_17417,N_13293);
and U23060 (N_23060,N_14838,N_15396);
nor U23061 (N_23061,N_16242,N_12563);
xnor U23062 (N_23062,N_15075,N_16732);
nand U23063 (N_23063,N_15394,N_12575);
nand U23064 (N_23064,N_17775,N_15219);
xnor U23065 (N_23065,N_16760,N_12938);
or U23066 (N_23066,N_15435,N_15659);
nor U23067 (N_23067,N_17586,N_13176);
and U23068 (N_23068,N_16048,N_17785);
nor U23069 (N_23069,N_12266,N_13736);
xor U23070 (N_23070,N_17979,N_14015);
nor U23071 (N_23071,N_14387,N_15144);
or U23072 (N_23072,N_15173,N_15375);
xnor U23073 (N_23073,N_16141,N_17541);
or U23074 (N_23074,N_17177,N_12298);
xor U23075 (N_23075,N_12104,N_15353);
and U23076 (N_23076,N_12402,N_17813);
and U23077 (N_23077,N_15921,N_14441);
or U23078 (N_23078,N_14576,N_12726);
or U23079 (N_23079,N_15789,N_12135);
or U23080 (N_23080,N_13656,N_16444);
nor U23081 (N_23081,N_15285,N_15580);
and U23082 (N_23082,N_16509,N_13476);
or U23083 (N_23083,N_15211,N_17138);
nor U23084 (N_23084,N_15047,N_15479);
or U23085 (N_23085,N_15851,N_13976);
and U23086 (N_23086,N_13461,N_16810);
or U23087 (N_23087,N_17922,N_16093);
nand U23088 (N_23088,N_12010,N_13099);
or U23089 (N_23089,N_12759,N_16973);
or U23090 (N_23090,N_13622,N_15148);
nand U23091 (N_23091,N_17511,N_14706);
nor U23092 (N_23092,N_13250,N_12076);
xor U23093 (N_23093,N_17145,N_17587);
or U23094 (N_23094,N_15849,N_14995);
xnor U23095 (N_23095,N_15899,N_17170);
or U23096 (N_23096,N_13742,N_13437);
nor U23097 (N_23097,N_15447,N_16751);
xnor U23098 (N_23098,N_13366,N_15981);
and U23099 (N_23099,N_17933,N_14539);
nor U23100 (N_23100,N_14747,N_14707);
nand U23101 (N_23101,N_14994,N_14767);
or U23102 (N_23102,N_14085,N_14483);
nor U23103 (N_23103,N_13655,N_12385);
nor U23104 (N_23104,N_13841,N_16187);
xnor U23105 (N_23105,N_15894,N_16235);
or U23106 (N_23106,N_14809,N_15056);
nor U23107 (N_23107,N_13948,N_14315);
or U23108 (N_23108,N_12292,N_12922);
or U23109 (N_23109,N_15097,N_12217);
or U23110 (N_23110,N_17823,N_14289);
nand U23111 (N_23111,N_12301,N_16277);
nor U23112 (N_23112,N_12166,N_17290);
nor U23113 (N_23113,N_17216,N_17535);
xor U23114 (N_23114,N_12059,N_14220);
or U23115 (N_23115,N_12926,N_15624);
xor U23116 (N_23116,N_14137,N_15123);
or U23117 (N_23117,N_15210,N_14788);
or U23118 (N_23118,N_17539,N_12026);
xor U23119 (N_23119,N_17081,N_13616);
xnor U23120 (N_23120,N_12645,N_14148);
or U23121 (N_23121,N_17056,N_16285);
nor U23122 (N_23122,N_14851,N_13132);
or U23123 (N_23123,N_12779,N_16256);
nand U23124 (N_23124,N_12220,N_13670);
nor U23125 (N_23125,N_17607,N_16987);
or U23126 (N_23126,N_17141,N_14269);
nor U23127 (N_23127,N_17925,N_14907);
nand U23128 (N_23128,N_14469,N_15078);
nor U23129 (N_23129,N_16025,N_14545);
xnor U23130 (N_23130,N_17203,N_17783);
or U23131 (N_23131,N_14789,N_17093);
or U23132 (N_23132,N_17510,N_14154);
nor U23133 (N_23133,N_15906,N_12406);
nor U23134 (N_23134,N_17263,N_15096);
and U23135 (N_23135,N_13660,N_13100);
or U23136 (N_23136,N_16809,N_12902);
nor U23137 (N_23137,N_15653,N_16367);
nor U23138 (N_23138,N_15770,N_15667);
or U23139 (N_23139,N_15942,N_13208);
and U23140 (N_23140,N_16217,N_13528);
nor U23141 (N_23141,N_12012,N_14718);
or U23142 (N_23142,N_14869,N_12973);
xor U23143 (N_23143,N_14544,N_14856);
or U23144 (N_23144,N_12284,N_13465);
nor U23145 (N_23145,N_13308,N_14036);
or U23146 (N_23146,N_16770,N_17517);
nand U23147 (N_23147,N_17348,N_14336);
or U23148 (N_23148,N_14062,N_17253);
nor U23149 (N_23149,N_17840,N_13258);
xnor U23150 (N_23150,N_14175,N_12831);
and U23151 (N_23151,N_13428,N_15385);
nand U23152 (N_23152,N_17032,N_17316);
nor U23153 (N_23153,N_12362,N_16563);
and U23154 (N_23154,N_12425,N_16803);
nand U23155 (N_23155,N_16406,N_12259);
and U23156 (N_23156,N_16375,N_13553);
nand U23157 (N_23157,N_14783,N_13299);
or U23158 (N_23158,N_12267,N_12382);
xor U23159 (N_23159,N_15209,N_17341);
and U23160 (N_23160,N_14245,N_16362);
and U23161 (N_23161,N_17846,N_14963);
or U23162 (N_23162,N_14871,N_16057);
nand U23163 (N_23163,N_14578,N_12064);
and U23164 (N_23164,N_15356,N_12238);
nand U23165 (N_23165,N_17872,N_14882);
or U23166 (N_23166,N_15672,N_17800);
or U23167 (N_23167,N_13334,N_15073);
xor U23168 (N_23168,N_17781,N_15425);
or U23169 (N_23169,N_16392,N_14189);
nor U23170 (N_23170,N_17015,N_16483);
nand U23171 (N_23171,N_12957,N_17970);
or U23172 (N_23172,N_17741,N_13033);
nand U23173 (N_23173,N_12122,N_14726);
nor U23174 (N_23174,N_17078,N_17630);
or U23175 (N_23175,N_12639,N_14628);
nor U23176 (N_23176,N_14221,N_13802);
and U23177 (N_23177,N_16274,N_17133);
nand U23178 (N_23178,N_15192,N_15460);
or U23179 (N_23179,N_14430,N_16076);
xnor U23180 (N_23180,N_15052,N_17653);
and U23181 (N_23181,N_14615,N_13960);
nand U23182 (N_23182,N_13325,N_14617);
nor U23183 (N_23183,N_13246,N_13057);
nor U23184 (N_23184,N_16392,N_12549);
nand U23185 (N_23185,N_17551,N_17636);
nor U23186 (N_23186,N_12359,N_16658);
or U23187 (N_23187,N_17497,N_17580);
or U23188 (N_23188,N_15981,N_17859);
nor U23189 (N_23189,N_14329,N_15713);
or U23190 (N_23190,N_14823,N_15676);
or U23191 (N_23191,N_12017,N_16187);
nor U23192 (N_23192,N_12934,N_14666);
nor U23193 (N_23193,N_12963,N_13131);
or U23194 (N_23194,N_15291,N_17643);
nand U23195 (N_23195,N_14261,N_13845);
nor U23196 (N_23196,N_15748,N_15410);
and U23197 (N_23197,N_15134,N_15993);
nand U23198 (N_23198,N_12220,N_12853);
and U23199 (N_23199,N_12319,N_13932);
or U23200 (N_23200,N_15785,N_15564);
nor U23201 (N_23201,N_14782,N_15933);
and U23202 (N_23202,N_13496,N_17287);
nand U23203 (N_23203,N_15765,N_16412);
and U23204 (N_23204,N_13639,N_16078);
nand U23205 (N_23205,N_16890,N_17100);
or U23206 (N_23206,N_12291,N_15046);
nor U23207 (N_23207,N_16409,N_17115);
nor U23208 (N_23208,N_16101,N_15383);
nand U23209 (N_23209,N_17014,N_15188);
nor U23210 (N_23210,N_16689,N_15166);
nand U23211 (N_23211,N_16590,N_13102);
nor U23212 (N_23212,N_17458,N_15749);
nand U23213 (N_23213,N_12778,N_14981);
and U23214 (N_23214,N_14481,N_12703);
nand U23215 (N_23215,N_15681,N_16104);
or U23216 (N_23216,N_17833,N_17332);
nor U23217 (N_23217,N_16862,N_16605);
xor U23218 (N_23218,N_12297,N_15022);
nor U23219 (N_23219,N_12953,N_15354);
nor U23220 (N_23220,N_16213,N_14141);
and U23221 (N_23221,N_17166,N_14827);
and U23222 (N_23222,N_14014,N_17276);
and U23223 (N_23223,N_12951,N_16074);
and U23224 (N_23224,N_12188,N_15814);
nor U23225 (N_23225,N_12905,N_16797);
nand U23226 (N_23226,N_14062,N_15952);
or U23227 (N_23227,N_13622,N_12014);
nand U23228 (N_23228,N_13387,N_15202);
nor U23229 (N_23229,N_15069,N_12647);
nand U23230 (N_23230,N_14192,N_15071);
nand U23231 (N_23231,N_12296,N_14639);
nand U23232 (N_23232,N_13883,N_15504);
nor U23233 (N_23233,N_16287,N_12102);
xnor U23234 (N_23234,N_13682,N_12581);
and U23235 (N_23235,N_17868,N_16181);
xor U23236 (N_23236,N_16670,N_16478);
nor U23237 (N_23237,N_15437,N_17164);
nor U23238 (N_23238,N_14541,N_13462);
or U23239 (N_23239,N_13011,N_12718);
nor U23240 (N_23240,N_17482,N_17759);
and U23241 (N_23241,N_16145,N_12471);
nor U23242 (N_23242,N_13108,N_16344);
xor U23243 (N_23243,N_16595,N_13805);
nand U23244 (N_23244,N_12034,N_14677);
xnor U23245 (N_23245,N_14150,N_15335);
xor U23246 (N_23246,N_12163,N_17560);
and U23247 (N_23247,N_12129,N_14732);
nand U23248 (N_23248,N_12977,N_16174);
and U23249 (N_23249,N_15157,N_15604);
xnor U23250 (N_23250,N_15358,N_16892);
nand U23251 (N_23251,N_12353,N_16382);
xor U23252 (N_23252,N_15952,N_12230);
xnor U23253 (N_23253,N_17616,N_15154);
nand U23254 (N_23254,N_15000,N_15589);
or U23255 (N_23255,N_16116,N_17793);
nand U23256 (N_23256,N_14964,N_12251);
nand U23257 (N_23257,N_15275,N_14656);
xor U23258 (N_23258,N_15205,N_13961);
or U23259 (N_23259,N_15381,N_14327);
xor U23260 (N_23260,N_14855,N_15346);
and U23261 (N_23261,N_13545,N_12656);
or U23262 (N_23262,N_12835,N_12302);
or U23263 (N_23263,N_12975,N_12724);
and U23264 (N_23264,N_12192,N_16179);
or U23265 (N_23265,N_14025,N_16335);
nor U23266 (N_23266,N_15004,N_14258);
nor U23267 (N_23267,N_16681,N_12894);
nand U23268 (N_23268,N_17064,N_14087);
xnor U23269 (N_23269,N_14319,N_14378);
or U23270 (N_23270,N_14056,N_16518);
and U23271 (N_23271,N_13669,N_16537);
and U23272 (N_23272,N_13761,N_13290);
nor U23273 (N_23273,N_17000,N_16324);
nand U23274 (N_23274,N_14834,N_17910);
and U23275 (N_23275,N_14554,N_13032);
nand U23276 (N_23276,N_16847,N_14657);
and U23277 (N_23277,N_12652,N_13775);
xor U23278 (N_23278,N_14724,N_13954);
xnor U23279 (N_23279,N_16972,N_16937);
xnor U23280 (N_23280,N_14643,N_15424);
nor U23281 (N_23281,N_12727,N_15810);
nand U23282 (N_23282,N_15524,N_15388);
and U23283 (N_23283,N_13381,N_17453);
xnor U23284 (N_23284,N_12078,N_15736);
and U23285 (N_23285,N_12844,N_14372);
and U23286 (N_23286,N_16321,N_12506);
or U23287 (N_23287,N_17794,N_15105);
nor U23288 (N_23288,N_14178,N_14811);
and U23289 (N_23289,N_13600,N_15860);
or U23290 (N_23290,N_13697,N_14406);
xor U23291 (N_23291,N_14975,N_15662);
nor U23292 (N_23292,N_16089,N_17081);
nand U23293 (N_23293,N_16806,N_16629);
nor U23294 (N_23294,N_12312,N_14167);
nor U23295 (N_23295,N_16690,N_14626);
or U23296 (N_23296,N_13897,N_12754);
nand U23297 (N_23297,N_14151,N_12402);
and U23298 (N_23298,N_17812,N_15202);
nor U23299 (N_23299,N_12515,N_15083);
nand U23300 (N_23300,N_16789,N_13294);
and U23301 (N_23301,N_13322,N_15911);
and U23302 (N_23302,N_14542,N_15816);
nor U23303 (N_23303,N_14502,N_16479);
and U23304 (N_23304,N_15168,N_17686);
xor U23305 (N_23305,N_15304,N_13343);
xor U23306 (N_23306,N_14217,N_14685);
and U23307 (N_23307,N_17764,N_16846);
nand U23308 (N_23308,N_17546,N_13063);
or U23309 (N_23309,N_14367,N_15991);
or U23310 (N_23310,N_15417,N_13674);
nand U23311 (N_23311,N_16094,N_13211);
or U23312 (N_23312,N_12813,N_15494);
nand U23313 (N_23313,N_13457,N_12545);
nand U23314 (N_23314,N_17990,N_14100);
nor U23315 (N_23315,N_12839,N_16038);
nor U23316 (N_23316,N_16533,N_17673);
and U23317 (N_23317,N_15023,N_14612);
nor U23318 (N_23318,N_16357,N_13650);
nor U23319 (N_23319,N_15839,N_12363);
nand U23320 (N_23320,N_13129,N_15899);
xnor U23321 (N_23321,N_17478,N_14147);
and U23322 (N_23322,N_12492,N_12704);
nor U23323 (N_23323,N_14390,N_16647);
nor U23324 (N_23324,N_15270,N_15099);
or U23325 (N_23325,N_17540,N_13936);
xor U23326 (N_23326,N_16996,N_16013);
xnor U23327 (N_23327,N_14888,N_15202);
nand U23328 (N_23328,N_15962,N_15978);
nor U23329 (N_23329,N_13095,N_14722);
or U23330 (N_23330,N_14670,N_13169);
and U23331 (N_23331,N_15153,N_15691);
or U23332 (N_23332,N_12447,N_13515);
or U23333 (N_23333,N_14773,N_16729);
or U23334 (N_23334,N_12348,N_14551);
nor U23335 (N_23335,N_15943,N_14522);
nand U23336 (N_23336,N_17054,N_15798);
nand U23337 (N_23337,N_13523,N_13530);
or U23338 (N_23338,N_16690,N_12106);
nand U23339 (N_23339,N_17357,N_12650);
or U23340 (N_23340,N_14746,N_17240);
nand U23341 (N_23341,N_16998,N_12950);
or U23342 (N_23342,N_15178,N_17300);
nand U23343 (N_23343,N_14442,N_17748);
or U23344 (N_23344,N_17372,N_15306);
and U23345 (N_23345,N_13888,N_17083);
xnor U23346 (N_23346,N_16635,N_16685);
xnor U23347 (N_23347,N_17841,N_13521);
and U23348 (N_23348,N_14967,N_12004);
nand U23349 (N_23349,N_13440,N_15082);
xor U23350 (N_23350,N_13674,N_17020);
and U23351 (N_23351,N_17910,N_16980);
nor U23352 (N_23352,N_17299,N_17881);
nor U23353 (N_23353,N_13084,N_16618);
nor U23354 (N_23354,N_15279,N_13334);
or U23355 (N_23355,N_12896,N_15111);
or U23356 (N_23356,N_14533,N_14555);
xor U23357 (N_23357,N_16065,N_16277);
xor U23358 (N_23358,N_15989,N_14778);
xor U23359 (N_23359,N_12918,N_13379);
and U23360 (N_23360,N_16906,N_15279);
or U23361 (N_23361,N_12827,N_15864);
nor U23362 (N_23362,N_15755,N_14284);
or U23363 (N_23363,N_17627,N_14997);
nand U23364 (N_23364,N_16184,N_16898);
and U23365 (N_23365,N_12327,N_14550);
and U23366 (N_23366,N_12022,N_16286);
nand U23367 (N_23367,N_17927,N_16647);
and U23368 (N_23368,N_16270,N_17846);
and U23369 (N_23369,N_15690,N_12543);
nand U23370 (N_23370,N_14796,N_14702);
nand U23371 (N_23371,N_12900,N_14504);
nand U23372 (N_23372,N_16237,N_15616);
nand U23373 (N_23373,N_15791,N_15611);
nand U23374 (N_23374,N_14443,N_15074);
or U23375 (N_23375,N_14705,N_13416);
or U23376 (N_23376,N_14197,N_17401);
nor U23377 (N_23377,N_15041,N_15230);
xor U23378 (N_23378,N_13185,N_17071);
nor U23379 (N_23379,N_12308,N_17505);
or U23380 (N_23380,N_15903,N_13016);
or U23381 (N_23381,N_12856,N_17883);
nor U23382 (N_23382,N_14405,N_14904);
or U23383 (N_23383,N_13182,N_16008);
nor U23384 (N_23384,N_12140,N_17749);
xnor U23385 (N_23385,N_12368,N_17148);
nand U23386 (N_23386,N_17225,N_17209);
and U23387 (N_23387,N_13208,N_13366);
and U23388 (N_23388,N_13620,N_17717);
nor U23389 (N_23389,N_13101,N_14428);
and U23390 (N_23390,N_13518,N_14555);
nand U23391 (N_23391,N_14079,N_12063);
and U23392 (N_23392,N_14413,N_13535);
nor U23393 (N_23393,N_17643,N_13709);
and U23394 (N_23394,N_12047,N_15884);
nand U23395 (N_23395,N_12587,N_17240);
nand U23396 (N_23396,N_17832,N_17419);
nor U23397 (N_23397,N_13218,N_16765);
xor U23398 (N_23398,N_17440,N_15389);
and U23399 (N_23399,N_16996,N_13346);
or U23400 (N_23400,N_12979,N_17129);
nor U23401 (N_23401,N_12871,N_17655);
or U23402 (N_23402,N_16439,N_13543);
xnor U23403 (N_23403,N_12227,N_14095);
or U23404 (N_23404,N_12706,N_14370);
nand U23405 (N_23405,N_16374,N_16188);
and U23406 (N_23406,N_13300,N_14983);
and U23407 (N_23407,N_13355,N_13224);
or U23408 (N_23408,N_14422,N_14602);
nand U23409 (N_23409,N_13017,N_14882);
and U23410 (N_23410,N_14463,N_15446);
nand U23411 (N_23411,N_12139,N_13065);
and U23412 (N_23412,N_15257,N_15910);
nand U23413 (N_23413,N_14543,N_16353);
and U23414 (N_23414,N_13693,N_14843);
nor U23415 (N_23415,N_17560,N_13413);
xnor U23416 (N_23416,N_13707,N_16181);
xor U23417 (N_23417,N_14974,N_16021);
nor U23418 (N_23418,N_15236,N_13006);
nand U23419 (N_23419,N_14548,N_17829);
nor U23420 (N_23420,N_17359,N_17863);
and U23421 (N_23421,N_15769,N_17200);
xnor U23422 (N_23422,N_13709,N_13901);
nand U23423 (N_23423,N_14087,N_16996);
and U23424 (N_23424,N_14603,N_14609);
xor U23425 (N_23425,N_16223,N_16863);
and U23426 (N_23426,N_14567,N_17871);
nor U23427 (N_23427,N_16673,N_16218);
xnor U23428 (N_23428,N_16656,N_14046);
nand U23429 (N_23429,N_13793,N_17345);
or U23430 (N_23430,N_12395,N_14707);
xnor U23431 (N_23431,N_14620,N_17696);
and U23432 (N_23432,N_14075,N_16290);
and U23433 (N_23433,N_12707,N_16076);
nor U23434 (N_23434,N_14488,N_13891);
and U23435 (N_23435,N_17911,N_16804);
nor U23436 (N_23436,N_16531,N_17933);
nand U23437 (N_23437,N_15679,N_17859);
or U23438 (N_23438,N_14507,N_13498);
xnor U23439 (N_23439,N_12576,N_17127);
nand U23440 (N_23440,N_16093,N_16037);
or U23441 (N_23441,N_15902,N_14072);
nor U23442 (N_23442,N_15341,N_15892);
nand U23443 (N_23443,N_16222,N_16692);
xor U23444 (N_23444,N_14312,N_17055);
xnor U23445 (N_23445,N_17775,N_17618);
and U23446 (N_23446,N_14415,N_16711);
and U23447 (N_23447,N_15341,N_15553);
or U23448 (N_23448,N_12327,N_17936);
or U23449 (N_23449,N_16841,N_12121);
xor U23450 (N_23450,N_13454,N_15192);
xnor U23451 (N_23451,N_14992,N_17133);
xor U23452 (N_23452,N_14391,N_12494);
nor U23453 (N_23453,N_15612,N_13760);
nand U23454 (N_23454,N_14830,N_15377);
or U23455 (N_23455,N_14996,N_15758);
nor U23456 (N_23456,N_16654,N_12947);
xor U23457 (N_23457,N_15195,N_16764);
and U23458 (N_23458,N_12869,N_12291);
or U23459 (N_23459,N_12460,N_15179);
or U23460 (N_23460,N_12552,N_14039);
and U23461 (N_23461,N_14422,N_17916);
xnor U23462 (N_23462,N_13234,N_15784);
or U23463 (N_23463,N_14199,N_12524);
or U23464 (N_23464,N_15219,N_14942);
or U23465 (N_23465,N_16255,N_15913);
and U23466 (N_23466,N_13804,N_13821);
nor U23467 (N_23467,N_15670,N_17681);
and U23468 (N_23468,N_17151,N_17556);
nor U23469 (N_23469,N_16553,N_12814);
nor U23470 (N_23470,N_12822,N_15245);
and U23471 (N_23471,N_15385,N_12841);
or U23472 (N_23472,N_17054,N_12094);
or U23473 (N_23473,N_17493,N_14301);
nand U23474 (N_23474,N_12191,N_16892);
xnor U23475 (N_23475,N_14867,N_12593);
or U23476 (N_23476,N_12517,N_15295);
xor U23477 (N_23477,N_12196,N_15038);
nand U23478 (N_23478,N_16184,N_15194);
nand U23479 (N_23479,N_16281,N_14852);
or U23480 (N_23480,N_17172,N_15519);
nor U23481 (N_23481,N_12603,N_12828);
nor U23482 (N_23482,N_15008,N_15788);
and U23483 (N_23483,N_14815,N_15744);
and U23484 (N_23484,N_13283,N_15749);
nand U23485 (N_23485,N_14107,N_14371);
and U23486 (N_23486,N_12738,N_17595);
nor U23487 (N_23487,N_15831,N_12191);
nand U23488 (N_23488,N_15101,N_13147);
xnor U23489 (N_23489,N_14083,N_16498);
nand U23490 (N_23490,N_15127,N_15383);
nand U23491 (N_23491,N_16218,N_13897);
xor U23492 (N_23492,N_14203,N_12050);
xnor U23493 (N_23493,N_17043,N_15933);
nand U23494 (N_23494,N_15862,N_16206);
and U23495 (N_23495,N_16777,N_13740);
nor U23496 (N_23496,N_17925,N_12350);
or U23497 (N_23497,N_15564,N_14144);
or U23498 (N_23498,N_15756,N_15379);
xor U23499 (N_23499,N_17872,N_14805);
xnor U23500 (N_23500,N_14093,N_12959);
nand U23501 (N_23501,N_17196,N_14180);
or U23502 (N_23502,N_17302,N_16988);
nor U23503 (N_23503,N_16347,N_12461);
or U23504 (N_23504,N_12611,N_15474);
xnor U23505 (N_23505,N_14972,N_12710);
nor U23506 (N_23506,N_16353,N_16389);
or U23507 (N_23507,N_13057,N_14361);
xor U23508 (N_23508,N_12825,N_12355);
and U23509 (N_23509,N_13997,N_13565);
xnor U23510 (N_23510,N_15690,N_15329);
nand U23511 (N_23511,N_12281,N_14001);
xnor U23512 (N_23512,N_14041,N_12898);
and U23513 (N_23513,N_13002,N_14408);
nor U23514 (N_23514,N_14443,N_16792);
nor U23515 (N_23515,N_15441,N_15328);
nand U23516 (N_23516,N_16449,N_13647);
xnor U23517 (N_23517,N_13290,N_15783);
or U23518 (N_23518,N_17303,N_13597);
xnor U23519 (N_23519,N_14874,N_15379);
nor U23520 (N_23520,N_15078,N_12951);
or U23521 (N_23521,N_13595,N_14430);
and U23522 (N_23522,N_13206,N_12376);
or U23523 (N_23523,N_12698,N_13860);
nor U23524 (N_23524,N_16390,N_12101);
nor U23525 (N_23525,N_12523,N_14935);
and U23526 (N_23526,N_16944,N_12869);
or U23527 (N_23527,N_13581,N_16260);
or U23528 (N_23528,N_12592,N_17934);
or U23529 (N_23529,N_14283,N_15637);
and U23530 (N_23530,N_13261,N_16097);
nor U23531 (N_23531,N_12265,N_17066);
or U23532 (N_23532,N_16255,N_12644);
nor U23533 (N_23533,N_17881,N_16539);
nand U23534 (N_23534,N_13824,N_12321);
nand U23535 (N_23535,N_12553,N_14648);
xor U23536 (N_23536,N_17447,N_16212);
xnor U23537 (N_23537,N_17587,N_14191);
or U23538 (N_23538,N_13072,N_17163);
xnor U23539 (N_23539,N_17363,N_13074);
nand U23540 (N_23540,N_16291,N_16286);
and U23541 (N_23541,N_12457,N_16254);
xnor U23542 (N_23542,N_12907,N_17664);
xnor U23543 (N_23543,N_12570,N_15046);
or U23544 (N_23544,N_13983,N_13306);
and U23545 (N_23545,N_13215,N_17038);
xnor U23546 (N_23546,N_16197,N_14913);
and U23547 (N_23547,N_16258,N_16787);
and U23548 (N_23548,N_15338,N_17292);
xnor U23549 (N_23549,N_12201,N_15375);
and U23550 (N_23550,N_14530,N_15899);
or U23551 (N_23551,N_17305,N_17003);
and U23552 (N_23552,N_13183,N_12910);
nand U23553 (N_23553,N_17363,N_15732);
or U23554 (N_23554,N_16786,N_13204);
or U23555 (N_23555,N_16858,N_12318);
nor U23556 (N_23556,N_16939,N_12519);
xor U23557 (N_23557,N_15277,N_16375);
or U23558 (N_23558,N_13151,N_13544);
nand U23559 (N_23559,N_15199,N_12026);
nand U23560 (N_23560,N_17826,N_17701);
xor U23561 (N_23561,N_13966,N_15374);
or U23562 (N_23562,N_13691,N_17423);
and U23563 (N_23563,N_14073,N_12030);
or U23564 (N_23564,N_17016,N_17709);
nand U23565 (N_23565,N_14505,N_15725);
nand U23566 (N_23566,N_12243,N_14594);
nand U23567 (N_23567,N_13987,N_15820);
xor U23568 (N_23568,N_12757,N_15688);
or U23569 (N_23569,N_17242,N_17299);
nor U23570 (N_23570,N_13419,N_16780);
or U23571 (N_23571,N_17545,N_13995);
nor U23572 (N_23572,N_12816,N_16611);
or U23573 (N_23573,N_12274,N_13785);
or U23574 (N_23574,N_15739,N_12873);
or U23575 (N_23575,N_13573,N_17103);
nand U23576 (N_23576,N_13251,N_15625);
nand U23577 (N_23577,N_13749,N_17667);
nor U23578 (N_23578,N_17483,N_14772);
nor U23579 (N_23579,N_15068,N_14474);
and U23580 (N_23580,N_17917,N_12779);
nor U23581 (N_23581,N_13460,N_15079);
and U23582 (N_23582,N_14516,N_15111);
and U23583 (N_23583,N_14911,N_16316);
nand U23584 (N_23584,N_14691,N_16513);
xnor U23585 (N_23585,N_14732,N_14387);
xnor U23586 (N_23586,N_14779,N_12434);
nand U23587 (N_23587,N_16297,N_13460);
or U23588 (N_23588,N_12132,N_17591);
or U23589 (N_23589,N_12998,N_14170);
and U23590 (N_23590,N_12742,N_16007);
nand U23591 (N_23591,N_15935,N_13696);
nor U23592 (N_23592,N_14961,N_14486);
and U23593 (N_23593,N_16680,N_14060);
xor U23594 (N_23594,N_13501,N_17334);
nor U23595 (N_23595,N_15011,N_17331);
nor U23596 (N_23596,N_13090,N_13246);
and U23597 (N_23597,N_17643,N_16822);
and U23598 (N_23598,N_15578,N_15954);
xor U23599 (N_23599,N_12234,N_13777);
and U23600 (N_23600,N_13485,N_12244);
and U23601 (N_23601,N_16030,N_12790);
nand U23602 (N_23602,N_12413,N_14604);
xor U23603 (N_23603,N_12558,N_16899);
nand U23604 (N_23604,N_16244,N_17825);
or U23605 (N_23605,N_16401,N_16101);
nor U23606 (N_23606,N_12416,N_17078);
or U23607 (N_23607,N_14934,N_15112);
nor U23608 (N_23608,N_16485,N_16783);
xnor U23609 (N_23609,N_14588,N_15188);
and U23610 (N_23610,N_17829,N_17016);
or U23611 (N_23611,N_17840,N_14291);
or U23612 (N_23612,N_17135,N_14475);
nand U23613 (N_23613,N_15017,N_17773);
nor U23614 (N_23614,N_12470,N_15910);
xor U23615 (N_23615,N_15368,N_14422);
xnor U23616 (N_23616,N_13083,N_15682);
or U23617 (N_23617,N_16141,N_12909);
xnor U23618 (N_23618,N_14541,N_12206);
nand U23619 (N_23619,N_17252,N_14169);
nand U23620 (N_23620,N_16190,N_13802);
nor U23621 (N_23621,N_17582,N_13906);
xnor U23622 (N_23622,N_12987,N_16317);
xor U23623 (N_23623,N_16197,N_12613);
nand U23624 (N_23624,N_12368,N_14608);
or U23625 (N_23625,N_14832,N_13225);
and U23626 (N_23626,N_12680,N_12464);
nor U23627 (N_23627,N_15672,N_17366);
or U23628 (N_23628,N_16363,N_16366);
xnor U23629 (N_23629,N_17942,N_13525);
and U23630 (N_23630,N_13987,N_17952);
or U23631 (N_23631,N_12239,N_16551);
nand U23632 (N_23632,N_16227,N_13335);
nand U23633 (N_23633,N_16848,N_14997);
and U23634 (N_23634,N_12891,N_12500);
or U23635 (N_23635,N_15970,N_12417);
nor U23636 (N_23636,N_17506,N_16864);
nand U23637 (N_23637,N_17136,N_14466);
and U23638 (N_23638,N_17781,N_15614);
and U23639 (N_23639,N_16038,N_15771);
or U23640 (N_23640,N_17852,N_15701);
or U23641 (N_23641,N_17287,N_15292);
or U23642 (N_23642,N_16555,N_13942);
nor U23643 (N_23643,N_15811,N_15021);
xnor U23644 (N_23644,N_16399,N_15154);
xnor U23645 (N_23645,N_13656,N_15336);
xor U23646 (N_23646,N_16610,N_13612);
and U23647 (N_23647,N_12713,N_14229);
xor U23648 (N_23648,N_15881,N_13025);
and U23649 (N_23649,N_17048,N_12246);
nor U23650 (N_23650,N_16489,N_15614);
nor U23651 (N_23651,N_17559,N_17852);
xor U23652 (N_23652,N_12009,N_13604);
and U23653 (N_23653,N_16700,N_17738);
and U23654 (N_23654,N_14364,N_12011);
or U23655 (N_23655,N_16734,N_15629);
xor U23656 (N_23656,N_13776,N_12112);
or U23657 (N_23657,N_12840,N_15425);
or U23658 (N_23658,N_16528,N_16939);
nor U23659 (N_23659,N_14080,N_12336);
nor U23660 (N_23660,N_12320,N_17347);
nand U23661 (N_23661,N_12028,N_17016);
nand U23662 (N_23662,N_12655,N_16104);
nand U23663 (N_23663,N_16652,N_15849);
xnor U23664 (N_23664,N_13251,N_13195);
xnor U23665 (N_23665,N_16061,N_14188);
or U23666 (N_23666,N_14120,N_17161);
or U23667 (N_23667,N_17527,N_15427);
or U23668 (N_23668,N_12360,N_17695);
or U23669 (N_23669,N_13058,N_15988);
xnor U23670 (N_23670,N_14296,N_12700);
and U23671 (N_23671,N_16353,N_16652);
and U23672 (N_23672,N_12704,N_14506);
and U23673 (N_23673,N_13128,N_12229);
and U23674 (N_23674,N_16915,N_14793);
and U23675 (N_23675,N_12543,N_15655);
and U23676 (N_23676,N_16695,N_17396);
or U23677 (N_23677,N_16656,N_14453);
and U23678 (N_23678,N_17486,N_17382);
nand U23679 (N_23679,N_15392,N_14731);
nor U23680 (N_23680,N_17087,N_17873);
xor U23681 (N_23681,N_13668,N_17015);
xor U23682 (N_23682,N_17948,N_16932);
and U23683 (N_23683,N_14087,N_12764);
and U23684 (N_23684,N_13614,N_17796);
or U23685 (N_23685,N_13777,N_16349);
or U23686 (N_23686,N_15339,N_14218);
xnor U23687 (N_23687,N_15446,N_13773);
and U23688 (N_23688,N_12563,N_14248);
nand U23689 (N_23689,N_16507,N_12251);
xnor U23690 (N_23690,N_16667,N_15143);
and U23691 (N_23691,N_14097,N_17485);
nor U23692 (N_23692,N_12865,N_12776);
nor U23693 (N_23693,N_15834,N_14252);
or U23694 (N_23694,N_17958,N_16000);
nand U23695 (N_23695,N_13360,N_17822);
xor U23696 (N_23696,N_12924,N_13438);
nor U23697 (N_23697,N_17665,N_12796);
xnor U23698 (N_23698,N_14782,N_14646);
xor U23699 (N_23699,N_14938,N_16482);
nand U23700 (N_23700,N_14831,N_16289);
or U23701 (N_23701,N_15835,N_13487);
xor U23702 (N_23702,N_16136,N_17019);
nand U23703 (N_23703,N_15139,N_15981);
nor U23704 (N_23704,N_12393,N_13537);
nand U23705 (N_23705,N_16869,N_17693);
xnor U23706 (N_23706,N_17803,N_16558);
and U23707 (N_23707,N_15286,N_16138);
and U23708 (N_23708,N_12384,N_13962);
nor U23709 (N_23709,N_17974,N_12253);
nor U23710 (N_23710,N_13568,N_12986);
nand U23711 (N_23711,N_17374,N_17075);
or U23712 (N_23712,N_16463,N_15285);
or U23713 (N_23713,N_15598,N_12106);
or U23714 (N_23714,N_17175,N_13038);
xnor U23715 (N_23715,N_14994,N_14973);
or U23716 (N_23716,N_16900,N_15301);
or U23717 (N_23717,N_14853,N_15770);
nor U23718 (N_23718,N_13841,N_13573);
and U23719 (N_23719,N_16715,N_16598);
or U23720 (N_23720,N_17356,N_16427);
or U23721 (N_23721,N_15795,N_16102);
nor U23722 (N_23722,N_14364,N_17924);
xnor U23723 (N_23723,N_15737,N_14802);
or U23724 (N_23724,N_14776,N_15666);
and U23725 (N_23725,N_15680,N_16506);
xnor U23726 (N_23726,N_16140,N_16488);
nor U23727 (N_23727,N_17917,N_14715);
nand U23728 (N_23728,N_13487,N_16404);
and U23729 (N_23729,N_16550,N_14562);
nand U23730 (N_23730,N_14869,N_16840);
nor U23731 (N_23731,N_16652,N_17783);
or U23732 (N_23732,N_14707,N_15968);
or U23733 (N_23733,N_12874,N_17234);
xnor U23734 (N_23734,N_15970,N_17404);
or U23735 (N_23735,N_16127,N_16486);
nor U23736 (N_23736,N_14926,N_13750);
xnor U23737 (N_23737,N_17476,N_17272);
nor U23738 (N_23738,N_14866,N_15112);
nor U23739 (N_23739,N_13433,N_12319);
or U23740 (N_23740,N_12610,N_12648);
or U23741 (N_23741,N_16396,N_12019);
nor U23742 (N_23742,N_12768,N_16485);
xnor U23743 (N_23743,N_13172,N_17132);
nor U23744 (N_23744,N_13849,N_16676);
or U23745 (N_23745,N_16441,N_12074);
nand U23746 (N_23746,N_12492,N_16595);
or U23747 (N_23747,N_12520,N_15713);
or U23748 (N_23748,N_16886,N_12563);
nor U23749 (N_23749,N_17657,N_14314);
and U23750 (N_23750,N_14874,N_15949);
nand U23751 (N_23751,N_13646,N_17665);
nor U23752 (N_23752,N_15581,N_12856);
and U23753 (N_23753,N_12841,N_14385);
or U23754 (N_23754,N_13330,N_17265);
nand U23755 (N_23755,N_12288,N_15673);
or U23756 (N_23756,N_15410,N_12235);
and U23757 (N_23757,N_16421,N_14547);
and U23758 (N_23758,N_17682,N_12146);
nand U23759 (N_23759,N_17792,N_16465);
and U23760 (N_23760,N_17779,N_14534);
xnor U23761 (N_23761,N_12992,N_13254);
nand U23762 (N_23762,N_17819,N_12943);
nand U23763 (N_23763,N_14913,N_12124);
nor U23764 (N_23764,N_14945,N_13193);
or U23765 (N_23765,N_15507,N_12637);
nor U23766 (N_23766,N_16058,N_17890);
or U23767 (N_23767,N_17817,N_13398);
xnor U23768 (N_23768,N_12990,N_12073);
or U23769 (N_23769,N_14021,N_17286);
xor U23770 (N_23770,N_16006,N_17686);
and U23771 (N_23771,N_15855,N_15477);
and U23772 (N_23772,N_14832,N_14565);
nand U23773 (N_23773,N_15941,N_16935);
nor U23774 (N_23774,N_16951,N_12901);
nor U23775 (N_23775,N_16004,N_14065);
and U23776 (N_23776,N_14692,N_15836);
nor U23777 (N_23777,N_17137,N_12809);
nor U23778 (N_23778,N_16916,N_13276);
nand U23779 (N_23779,N_13222,N_14469);
nand U23780 (N_23780,N_15175,N_12035);
nand U23781 (N_23781,N_12304,N_16140);
xnor U23782 (N_23782,N_12138,N_16639);
and U23783 (N_23783,N_15965,N_15488);
nor U23784 (N_23784,N_12426,N_13961);
or U23785 (N_23785,N_12491,N_13019);
or U23786 (N_23786,N_17859,N_13514);
and U23787 (N_23787,N_12799,N_15438);
or U23788 (N_23788,N_16424,N_13003);
and U23789 (N_23789,N_15545,N_17428);
nor U23790 (N_23790,N_16056,N_13265);
xor U23791 (N_23791,N_16543,N_12381);
nand U23792 (N_23792,N_16718,N_16692);
xor U23793 (N_23793,N_15296,N_15392);
and U23794 (N_23794,N_15654,N_13883);
xor U23795 (N_23795,N_13730,N_17532);
or U23796 (N_23796,N_14906,N_15536);
and U23797 (N_23797,N_15870,N_13963);
xor U23798 (N_23798,N_12434,N_15852);
xnor U23799 (N_23799,N_12222,N_15177);
xor U23800 (N_23800,N_13838,N_14033);
or U23801 (N_23801,N_17377,N_13901);
nand U23802 (N_23802,N_17700,N_15964);
nor U23803 (N_23803,N_15407,N_14454);
or U23804 (N_23804,N_15967,N_17050);
nand U23805 (N_23805,N_12056,N_16110);
and U23806 (N_23806,N_17270,N_15220);
nor U23807 (N_23807,N_17037,N_13185);
nand U23808 (N_23808,N_17297,N_17968);
nor U23809 (N_23809,N_16290,N_13321);
and U23810 (N_23810,N_15710,N_12602);
and U23811 (N_23811,N_15827,N_14062);
nor U23812 (N_23812,N_12293,N_16125);
nand U23813 (N_23813,N_17384,N_14967);
and U23814 (N_23814,N_13228,N_17679);
and U23815 (N_23815,N_13555,N_13386);
or U23816 (N_23816,N_15393,N_13214);
nand U23817 (N_23817,N_14811,N_17596);
nand U23818 (N_23818,N_12565,N_15492);
and U23819 (N_23819,N_15319,N_17973);
and U23820 (N_23820,N_15511,N_17966);
and U23821 (N_23821,N_14744,N_14958);
xor U23822 (N_23822,N_16096,N_15072);
nor U23823 (N_23823,N_16667,N_14352);
nor U23824 (N_23824,N_13403,N_13140);
or U23825 (N_23825,N_13293,N_16546);
xnor U23826 (N_23826,N_16004,N_12329);
xnor U23827 (N_23827,N_15147,N_12446);
or U23828 (N_23828,N_13254,N_14658);
and U23829 (N_23829,N_13000,N_15144);
xor U23830 (N_23830,N_17097,N_17954);
xnor U23831 (N_23831,N_15385,N_12855);
nand U23832 (N_23832,N_14197,N_15623);
and U23833 (N_23833,N_12744,N_13467);
and U23834 (N_23834,N_16206,N_13046);
or U23835 (N_23835,N_14272,N_12215);
nor U23836 (N_23836,N_16474,N_14961);
xor U23837 (N_23837,N_13655,N_13177);
or U23838 (N_23838,N_15788,N_14078);
nand U23839 (N_23839,N_12938,N_17204);
xnor U23840 (N_23840,N_14568,N_13906);
and U23841 (N_23841,N_17732,N_13752);
and U23842 (N_23842,N_12746,N_14961);
and U23843 (N_23843,N_17060,N_17480);
nand U23844 (N_23844,N_17437,N_17739);
nand U23845 (N_23845,N_16316,N_12102);
nor U23846 (N_23846,N_12868,N_13650);
nand U23847 (N_23847,N_17330,N_14873);
nand U23848 (N_23848,N_14510,N_17567);
nand U23849 (N_23849,N_16193,N_15210);
and U23850 (N_23850,N_17887,N_14802);
nor U23851 (N_23851,N_17669,N_16147);
xnor U23852 (N_23852,N_14174,N_12279);
nor U23853 (N_23853,N_17643,N_16914);
nor U23854 (N_23854,N_13065,N_13882);
and U23855 (N_23855,N_14599,N_17667);
xnor U23856 (N_23856,N_17241,N_13170);
xor U23857 (N_23857,N_16884,N_13656);
nor U23858 (N_23858,N_16575,N_17150);
and U23859 (N_23859,N_12167,N_17993);
nor U23860 (N_23860,N_13176,N_12430);
or U23861 (N_23861,N_15096,N_12485);
xnor U23862 (N_23862,N_16170,N_12616);
nand U23863 (N_23863,N_12888,N_17113);
and U23864 (N_23864,N_16506,N_17505);
nor U23865 (N_23865,N_15317,N_14664);
or U23866 (N_23866,N_15291,N_17120);
nor U23867 (N_23867,N_13458,N_16866);
and U23868 (N_23868,N_13908,N_13554);
or U23869 (N_23869,N_16136,N_14575);
xor U23870 (N_23870,N_17759,N_16902);
and U23871 (N_23871,N_12976,N_16299);
and U23872 (N_23872,N_16447,N_16865);
and U23873 (N_23873,N_15107,N_15563);
nor U23874 (N_23874,N_17248,N_15539);
nand U23875 (N_23875,N_13949,N_14883);
xnor U23876 (N_23876,N_14643,N_12277);
nor U23877 (N_23877,N_17828,N_17411);
nand U23878 (N_23878,N_15990,N_15177);
xor U23879 (N_23879,N_14515,N_14617);
xor U23880 (N_23880,N_16798,N_13804);
or U23881 (N_23881,N_15155,N_15258);
or U23882 (N_23882,N_14709,N_17380);
xnor U23883 (N_23883,N_13408,N_15474);
and U23884 (N_23884,N_17895,N_16481);
nor U23885 (N_23885,N_17534,N_16187);
nand U23886 (N_23886,N_12767,N_13163);
xor U23887 (N_23887,N_15730,N_17196);
nand U23888 (N_23888,N_16055,N_15663);
and U23889 (N_23889,N_14573,N_16898);
and U23890 (N_23890,N_13024,N_13225);
xor U23891 (N_23891,N_17305,N_12650);
xnor U23892 (N_23892,N_12885,N_12209);
or U23893 (N_23893,N_15558,N_13795);
nand U23894 (N_23894,N_12773,N_15258);
and U23895 (N_23895,N_14331,N_16093);
or U23896 (N_23896,N_15331,N_15168);
and U23897 (N_23897,N_13343,N_16431);
nand U23898 (N_23898,N_14941,N_15711);
or U23899 (N_23899,N_14107,N_13533);
nor U23900 (N_23900,N_12129,N_14576);
nand U23901 (N_23901,N_13194,N_17741);
xor U23902 (N_23902,N_16890,N_12825);
and U23903 (N_23903,N_13090,N_15281);
nor U23904 (N_23904,N_12196,N_12155);
or U23905 (N_23905,N_17753,N_13022);
or U23906 (N_23906,N_15334,N_16144);
or U23907 (N_23907,N_12210,N_17054);
or U23908 (N_23908,N_14917,N_12328);
nor U23909 (N_23909,N_17379,N_15133);
or U23910 (N_23910,N_14868,N_16360);
xor U23911 (N_23911,N_14816,N_13970);
or U23912 (N_23912,N_15694,N_17706);
nand U23913 (N_23913,N_15976,N_12431);
and U23914 (N_23914,N_15951,N_14202);
nand U23915 (N_23915,N_15715,N_15924);
nand U23916 (N_23916,N_13605,N_13580);
nand U23917 (N_23917,N_16380,N_13319);
nand U23918 (N_23918,N_17821,N_14440);
or U23919 (N_23919,N_12743,N_16120);
or U23920 (N_23920,N_13557,N_15917);
nor U23921 (N_23921,N_13194,N_15881);
nor U23922 (N_23922,N_13350,N_16160);
and U23923 (N_23923,N_13660,N_17786);
xor U23924 (N_23924,N_14232,N_13588);
xor U23925 (N_23925,N_13059,N_15124);
nor U23926 (N_23926,N_12565,N_17770);
nor U23927 (N_23927,N_15819,N_14095);
nand U23928 (N_23928,N_17706,N_14419);
nand U23929 (N_23929,N_13463,N_14664);
nor U23930 (N_23930,N_13328,N_16896);
xor U23931 (N_23931,N_14862,N_16543);
and U23932 (N_23932,N_16208,N_14171);
or U23933 (N_23933,N_13216,N_13507);
or U23934 (N_23934,N_16043,N_12333);
or U23935 (N_23935,N_12003,N_12493);
xor U23936 (N_23936,N_12902,N_17627);
and U23937 (N_23937,N_13920,N_16933);
nand U23938 (N_23938,N_13647,N_13274);
nor U23939 (N_23939,N_16913,N_12165);
nand U23940 (N_23940,N_17929,N_12633);
nand U23941 (N_23941,N_13630,N_16946);
nor U23942 (N_23942,N_13101,N_15310);
nand U23943 (N_23943,N_15504,N_17281);
or U23944 (N_23944,N_16902,N_16725);
nand U23945 (N_23945,N_17348,N_13274);
nand U23946 (N_23946,N_14737,N_16743);
nor U23947 (N_23947,N_13351,N_13792);
nand U23948 (N_23948,N_15683,N_17791);
or U23949 (N_23949,N_14798,N_17388);
xnor U23950 (N_23950,N_17291,N_15802);
xnor U23951 (N_23951,N_15017,N_16794);
xnor U23952 (N_23952,N_12848,N_17761);
nand U23953 (N_23953,N_17733,N_14666);
nor U23954 (N_23954,N_14399,N_16854);
or U23955 (N_23955,N_13645,N_12483);
and U23956 (N_23956,N_13157,N_16003);
nand U23957 (N_23957,N_17862,N_12769);
xnor U23958 (N_23958,N_16475,N_16759);
nand U23959 (N_23959,N_15215,N_13997);
xor U23960 (N_23960,N_17094,N_17732);
or U23961 (N_23961,N_14844,N_16135);
nand U23962 (N_23962,N_16803,N_17337);
or U23963 (N_23963,N_13779,N_15818);
or U23964 (N_23964,N_16878,N_17169);
nor U23965 (N_23965,N_17765,N_17993);
nor U23966 (N_23966,N_16453,N_15516);
nand U23967 (N_23967,N_16144,N_12295);
and U23968 (N_23968,N_13741,N_17928);
nor U23969 (N_23969,N_16189,N_12103);
or U23970 (N_23970,N_14753,N_16190);
and U23971 (N_23971,N_16154,N_13693);
and U23972 (N_23972,N_17524,N_17981);
nand U23973 (N_23973,N_14896,N_17488);
xor U23974 (N_23974,N_12398,N_12153);
xnor U23975 (N_23975,N_12341,N_15183);
nor U23976 (N_23976,N_16863,N_14075);
nor U23977 (N_23977,N_14859,N_15957);
or U23978 (N_23978,N_14412,N_17335);
and U23979 (N_23979,N_12187,N_17985);
and U23980 (N_23980,N_12901,N_17186);
nand U23981 (N_23981,N_13867,N_14404);
and U23982 (N_23982,N_12411,N_15402);
or U23983 (N_23983,N_12997,N_15597);
and U23984 (N_23984,N_16786,N_15726);
and U23985 (N_23985,N_17725,N_17308);
nor U23986 (N_23986,N_14392,N_13510);
nor U23987 (N_23987,N_15792,N_12572);
nor U23988 (N_23988,N_12090,N_14736);
xor U23989 (N_23989,N_13876,N_12435);
nand U23990 (N_23990,N_13215,N_17908);
and U23991 (N_23991,N_17906,N_12677);
and U23992 (N_23992,N_14653,N_15546);
or U23993 (N_23993,N_17528,N_16806);
xor U23994 (N_23994,N_17243,N_13125);
or U23995 (N_23995,N_17949,N_13918);
xnor U23996 (N_23996,N_17987,N_13413);
nor U23997 (N_23997,N_15948,N_14151);
or U23998 (N_23998,N_17079,N_13302);
nand U23999 (N_23999,N_16458,N_17656);
xnor U24000 (N_24000,N_18205,N_22047);
nand U24001 (N_24001,N_20035,N_21852);
or U24002 (N_24002,N_21170,N_19815);
and U24003 (N_24003,N_22197,N_23841);
nor U24004 (N_24004,N_21654,N_20537);
and U24005 (N_24005,N_22703,N_23543);
xnor U24006 (N_24006,N_18040,N_20010);
and U24007 (N_24007,N_19629,N_22586);
and U24008 (N_24008,N_20141,N_18630);
xnor U24009 (N_24009,N_22323,N_22301);
xnor U24010 (N_24010,N_20558,N_20873);
nand U24011 (N_24011,N_21776,N_19306);
and U24012 (N_24012,N_18828,N_20988);
nand U24013 (N_24013,N_21155,N_21977);
nand U24014 (N_24014,N_22438,N_23711);
or U24015 (N_24015,N_20439,N_22713);
or U24016 (N_24016,N_19543,N_20438);
nor U24017 (N_24017,N_22901,N_18925);
nand U24018 (N_24018,N_22730,N_23830);
or U24019 (N_24019,N_18006,N_22045);
nor U24020 (N_24020,N_21373,N_21433);
nand U24021 (N_24021,N_19180,N_18854);
nand U24022 (N_24022,N_19279,N_21163);
or U24023 (N_24023,N_18015,N_20581);
nor U24024 (N_24024,N_20163,N_22238);
nor U24025 (N_24025,N_22255,N_22284);
and U24026 (N_24026,N_19513,N_20591);
xor U24027 (N_24027,N_21764,N_21955);
nor U24028 (N_24028,N_20629,N_21631);
and U24029 (N_24029,N_22254,N_21933);
or U24030 (N_24030,N_21080,N_19136);
nand U24031 (N_24031,N_21385,N_21168);
nand U24032 (N_24032,N_20370,N_18566);
and U24033 (N_24033,N_18818,N_19985);
and U24034 (N_24034,N_20703,N_21138);
or U24035 (N_24035,N_19716,N_19025);
nand U24036 (N_24036,N_19503,N_21021);
nand U24037 (N_24037,N_23719,N_19208);
and U24038 (N_24038,N_21970,N_20274);
xnor U24039 (N_24039,N_21516,N_19921);
nand U24040 (N_24040,N_22220,N_21626);
or U24041 (N_24041,N_21335,N_20321);
or U24042 (N_24042,N_22972,N_20584);
nand U24043 (N_24043,N_21334,N_23089);
nor U24044 (N_24044,N_23201,N_21740);
or U24045 (N_24045,N_21087,N_21622);
xnor U24046 (N_24046,N_19825,N_21183);
nand U24047 (N_24047,N_18954,N_22479);
and U24048 (N_24048,N_20418,N_20011);
or U24049 (N_24049,N_22804,N_22240);
nor U24050 (N_24050,N_18826,N_18491);
nor U24051 (N_24051,N_22552,N_22020);
nand U24052 (N_24052,N_19528,N_22485);
xor U24053 (N_24053,N_22691,N_21417);
and U24054 (N_24054,N_19017,N_22705);
or U24055 (N_24055,N_20769,N_23413);
nor U24056 (N_24056,N_21054,N_20243);
and U24057 (N_24057,N_21046,N_19016);
and U24058 (N_24058,N_18486,N_22232);
and U24059 (N_24059,N_23786,N_19874);
and U24060 (N_24060,N_22398,N_21503);
xor U24061 (N_24061,N_21827,N_18938);
or U24062 (N_24062,N_18268,N_22328);
or U24063 (N_24063,N_20901,N_20775);
xnor U24064 (N_24064,N_23821,N_21092);
nor U24065 (N_24065,N_22982,N_19442);
and U24066 (N_24066,N_21634,N_21440);
xnor U24067 (N_24067,N_21070,N_21041);
nor U24068 (N_24068,N_22570,N_18649);
and U24069 (N_24069,N_18127,N_19858);
xnor U24070 (N_24070,N_20313,N_19781);
xor U24071 (N_24071,N_19769,N_19797);
and U24072 (N_24072,N_23883,N_23899);
and U24073 (N_24073,N_18937,N_18669);
nor U24074 (N_24074,N_21632,N_23735);
nand U24075 (N_24075,N_23073,N_22203);
nor U24076 (N_24076,N_19057,N_18347);
xor U24077 (N_24077,N_23502,N_21913);
xor U24078 (N_24078,N_18216,N_23355);
xnor U24079 (N_24079,N_23902,N_22511);
and U24080 (N_24080,N_21450,N_19758);
nand U24081 (N_24081,N_18408,N_21361);
nand U24082 (N_24082,N_20115,N_23006);
nand U24083 (N_24083,N_21627,N_22355);
and U24084 (N_24084,N_21297,N_20518);
nor U24085 (N_24085,N_20360,N_18373);
nor U24086 (N_24086,N_19586,N_21754);
nor U24087 (N_24087,N_18034,N_19979);
and U24088 (N_24088,N_22661,N_19474);
and U24089 (N_24089,N_18454,N_18188);
xor U24090 (N_24090,N_22787,N_20031);
nor U24091 (N_24091,N_21712,N_23927);
and U24092 (N_24092,N_18733,N_23866);
or U24093 (N_24093,N_23244,N_22354);
or U24094 (N_24094,N_19893,N_20477);
xor U24095 (N_24095,N_18775,N_23570);
xnor U24096 (N_24096,N_23546,N_18855);
nor U24097 (N_24097,N_19746,N_20950);
xor U24098 (N_24098,N_20738,N_21310);
and U24099 (N_24099,N_22537,N_18088);
and U24100 (N_24100,N_18354,N_23583);
xor U24101 (N_24101,N_18580,N_23731);
nor U24102 (N_24102,N_19414,N_19524);
nand U24103 (N_24103,N_19691,N_23196);
and U24104 (N_24104,N_20139,N_21427);
xor U24105 (N_24105,N_23634,N_20932);
or U24106 (N_24106,N_21796,N_23028);
nand U24107 (N_24107,N_19976,N_18880);
xor U24108 (N_24108,N_18716,N_19157);
or U24109 (N_24109,N_23998,N_18067);
and U24110 (N_24110,N_19191,N_21120);
nor U24111 (N_24111,N_23056,N_21483);
nand U24112 (N_24112,N_20917,N_19896);
or U24113 (N_24113,N_21069,N_20421);
nor U24114 (N_24114,N_21062,N_23331);
nor U24115 (N_24115,N_18583,N_20131);
nor U24116 (N_24116,N_18328,N_19268);
nand U24117 (N_24117,N_19164,N_21071);
and U24118 (N_24118,N_18461,N_19996);
and U24119 (N_24119,N_23441,N_18129);
xor U24120 (N_24120,N_22802,N_23525);
and U24121 (N_24121,N_23567,N_22739);
and U24122 (N_24122,N_23014,N_23052);
xor U24123 (N_24123,N_19271,N_23511);
and U24124 (N_24124,N_19201,N_22711);
nor U24125 (N_24125,N_22602,N_20691);
xor U24126 (N_24126,N_23924,N_22720);
or U24127 (N_24127,N_22628,N_20836);
nand U24128 (N_24128,N_23415,N_18315);
nand U24129 (N_24129,N_20788,N_22967);
and U24130 (N_24130,N_20546,N_18248);
xor U24131 (N_24131,N_20616,N_23746);
and U24132 (N_24132,N_21783,N_19661);
xnor U24133 (N_24133,N_23578,N_19723);
xnor U24134 (N_24134,N_21262,N_22187);
or U24135 (N_24135,N_20797,N_20534);
and U24136 (N_24136,N_19370,N_18675);
nor U24137 (N_24137,N_20527,N_18529);
and U24138 (N_24138,N_19476,N_22286);
nor U24139 (N_24139,N_18276,N_23231);
and U24140 (N_24140,N_22824,N_19491);
nand U24141 (N_24141,N_23433,N_22388);
nor U24142 (N_24142,N_23519,N_18996);
nand U24143 (N_24143,N_21969,N_21469);
xnor U24144 (N_24144,N_22662,N_19798);
xnor U24145 (N_24145,N_22578,N_21719);
nand U24146 (N_24146,N_23799,N_21676);
xnor U24147 (N_24147,N_19789,N_20772);
nor U24148 (N_24148,N_19071,N_18707);
and U24149 (N_24149,N_20297,N_23234);
nor U24150 (N_24150,N_21322,N_21937);
and U24151 (N_24151,N_22403,N_20771);
or U24152 (N_24152,N_18052,N_23862);
xor U24153 (N_24153,N_22743,N_22084);
xor U24154 (N_24154,N_23532,N_22140);
nor U24155 (N_24155,N_21714,N_23467);
nand U24156 (N_24156,N_22776,N_23263);
nand U24157 (N_24157,N_22077,N_23982);
and U24158 (N_24158,N_23309,N_20080);
and U24159 (N_24159,N_20663,N_23167);
nand U24160 (N_24160,N_20883,N_18555);
or U24161 (N_24161,N_23470,N_22626);
or U24162 (N_24162,N_21090,N_18693);
xnor U24163 (N_24163,N_18965,N_22740);
xnor U24164 (N_24164,N_22075,N_20083);
nand U24165 (N_24165,N_21329,N_22441);
and U24166 (N_24166,N_19533,N_18252);
nand U24167 (N_24167,N_20942,N_21761);
xnor U24168 (N_24168,N_19492,N_23586);
xnor U24169 (N_24169,N_22501,N_23638);
and U24170 (N_24170,N_22549,N_20577);
xor U24171 (N_24171,N_21823,N_23401);
nor U24172 (N_24172,N_23933,N_23100);
nor U24173 (N_24173,N_19568,N_23615);
xor U24174 (N_24174,N_23689,N_18064);
xor U24175 (N_24175,N_22550,N_20713);
and U24176 (N_24176,N_19888,N_19674);
nor U24177 (N_24177,N_20453,N_22619);
nor U24178 (N_24178,N_23725,N_19981);
nand U24179 (N_24179,N_20575,N_23417);
nand U24180 (N_24180,N_19160,N_19406);
xor U24181 (N_24181,N_22593,N_19504);
nor U24182 (N_24182,N_21699,N_20081);
and U24183 (N_24183,N_22091,N_21501);
xnor U24184 (N_24184,N_21957,N_19968);
or U24185 (N_24185,N_21481,N_21906);
and U24186 (N_24186,N_20768,N_22087);
nor U24187 (N_24187,N_18969,N_18763);
and U24188 (N_24188,N_22491,N_21193);
or U24189 (N_24189,N_19579,N_22569);
nand U24190 (N_24190,N_23487,N_23227);
nor U24191 (N_24191,N_18392,N_18189);
nand U24192 (N_24192,N_22031,N_21103);
nor U24193 (N_24193,N_22182,N_19448);
nor U24194 (N_24194,N_21221,N_21927);
or U24195 (N_24195,N_22684,N_22893);
or U24196 (N_24196,N_20432,N_19530);
and U24197 (N_24197,N_18109,N_22110);
nand U24198 (N_24198,N_23255,N_20200);
nor U24199 (N_24199,N_18961,N_22443);
and U24200 (N_24200,N_20258,N_20820);
nand U24201 (N_24201,N_19034,N_23350);
and U24202 (N_24202,N_22565,N_22474);
nand U24203 (N_24203,N_23642,N_20921);
nor U24204 (N_24204,N_20059,N_22099);
nor U24205 (N_24205,N_20981,N_23134);
or U24206 (N_24206,N_19879,N_20340);
nand U24207 (N_24207,N_18919,N_22811);
nand U24208 (N_24208,N_22794,N_20113);
xor U24209 (N_24209,N_21064,N_20995);
nor U24210 (N_24210,N_22295,N_23684);
nor U24211 (N_24211,N_21822,N_23647);
xnor U24212 (N_24212,N_18297,N_18776);
xnor U24213 (N_24213,N_23595,N_20716);
nor U24214 (N_24214,N_18719,N_23714);
xnor U24215 (N_24215,N_21930,N_18889);
and U24216 (N_24216,N_23284,N_20112);
or U24217 (N_24217,N_22483,N_20962);
or U24218 (N_24218,N_19375,N_23276);
xnor U24219 (N_24219,N_22715,N_23754);
xor U24220 (N_24220,N_21410,N_18947);
nand U24221 (N_24221,N_19141,N_22963);
or U24222 (N_24222,N_20322,N_21419);
nand U24223 (N_24223,N_23903,N_19464);
nand U24224 (N_24224,N_18728,N_23741);
xor U24225 (N_24225,N_20918,N_21086);
xnor U24226 (N_24226,N_20374,N_18406);
or U24227 (N_24227,N_19767,N_18869);
and U24228 (N_24228,N_21033,N_19235);
nand U24229 (N_24229,N_22104,N_20282);
nand U24230 (N_24230,N_20645,N_21404);
xnor U24231 (N_24231,N_18682,N_23437);
nor U24232 (N_24232,N_19473,N_23379);
xnor U24233 (N_24233,N_18738,N_23537);
nand U24234 (N_24234,N_18367,N_21106);
nand U24235 (N_24235,N_23592,N_23439);
or U24236 (N_24236,N_19876,N_20920);
and U24237 (N_24237,N_21313,N_23091);
and U24238 (N_24238,N_23337,N_21562);
nand U24239 (N_24239,N_20466,N_18255);
nor U24240 (N_24240,N_18635,N_20777);
or U24241 (N_24241,N_18332,N_18986);
nor U24242 (N_24242,N_23356,N_23846);
or U24243 (N_24243,N_18972,N_23608);
and U24244 (N_24244,N_22588,N_18398);
nand U24245 (N_24245,N_21771,N_23017);
or U24246 (N_24246,N_21416,N_23604);
and U24247 (N_24247,N_21078,N_21848);
nand U24248 (N_24248,N_22222,N_18732);
and U24249 (N_24249,N_22946,N_19582);
nand U24250 (N_24250,N_19840,N_20268);
xnor U24251 (N_24251,N_23010,N_23188);
xnor U24252 (N_24252,N_21066,N_23914);
and U24253 (N_24253,N_18514,N_20568);
and U24254 (N_24254,N_23249,N_19621);
nand U24255 (N_24255,N_23116,N_20504);
or U24256 (N_24256,N_19786,N_22025);
or U24257 (N_24257,N_20643,N_23823);
nand U24258 (N_24258,N_23357,N_21035);
nor U24259 (N_24259,N_22381,N_22952);
and U24260 (N_24260,N_18598,N_18816);
xnor U24261 (N_24261,N_21019,N_18209);
nand U24262 (N_24262,N_21871,N_20667);
xor U24263 (N_24263,N_18565,N_18208);
nand U24264 (N_24264,N_21040,N_23972);
nand U24265 (N_24265,N_19747,N_21294);
and U24266 (N_24266,N_19889,N_23645);
nor U24267 (N_24267,N_19713,N_23093);
and U24268 (N_24268,N_18845,N_21910);
xnor U24269 (N_24269,N_19842,N_18870);
and U24270 (N_24270,N_22094,N_19993);
and U24271 (N_24271,N_19174,N_19771);
nor U24272 (N_24272,N_20232,N_21047);
xor U24273 (N_24273,N_19429,N_23287);
and U24274 (N_24274,N_22379,N_18358);
or U24275 (N_24275,N_21794,N_18157);
nand U24276 (N_24276,N_19199,N_19760);
nor U24277 (N_24277,N_23890,N_21574);
xor U24278 (N_24278,N_18678,N_21475);
or U24279 (N_24279,N_18231,N_18631);
nor U24280 (N_24280,N_21721,N_22613);
nand U24281 (N_24281,N_23328,N_21301);
and U24282 (N_24282,N_23959,N_23917);
or U24283 (N_24283,N_21458,N_21662);
and U24284 (N_24284,N_22410,N_23784);
or U24285 (N_24285,N_18512,N_23538);
and U24286 (N_24286,N_20120,N_20092);
or U24287 (N_24287,N_22192,N_22627);
nor U24288 (N_24288,N_23698,N_21383);
xnor U24289 (N_24289,N_20044,N_22041);
xor U24290 (N_24290,N_22169,N_23336);
nand U24291 (N_24291,N_19881,N_23506);
xnor U24292 (N_24292,N_19950,N_19081);
nor U24293 (N_24293,N_19994,N_23226);
and U24294 (N_24294,N_23720,N_18547);
xnor U24295 (N_24295,N_21133,N_20467);
xor U24296 (N_24296,N_19850,N_22559);
nor U24297 (N_24297,N_18182,N_20613);
xor U24298 (N_24298,N_21032,N_19304);
xnor U24299 (N_24299,N_22945,N_18174);
and U24300 (N_24300,N_23974,N_22506);
or U24301 (N_24301,N_20850,N_20956);
nand U24302 (N_24302,N_19759,N_19008);
xor U24303 (N_24303,N_19142,N_21849);
and U24304 (N_24304,N_21462,N_23329);
nand U24305 (N_24305,N_23791,N_20114);
or U24306 (N_24306,N_23819,N_19363);
and U24307 (N_24307,N_23448,N_23870);
and U24308 (N_24308,N_23728,N_20676);
or U24309 (N_24309,N_18151,N_22180);
nand U24310 (N_24310,N_21303,N_18201);
and U24311 (N_24311,N_22716,N_19852);
or U24312 (N_24312,N_23335,N_22095);
nand U24313 (N_24313,N_23019,N_18743);
nor U24314 (N_24314,N_21247,N_22728);
or U24315 (N_24315,N_19820,N_22816);
or U24316 (N_24316,N_20034,N_21319);
nor U24317 (N_24317,N_22142,N_23076);
or U24318 (N_24318,N_22299,N_19772);
nor U24319 (N_24319,N_20763,N_23874);
xnor U24320 (N_24320,N_22562,N_22664);
or U24321 (N_24321,N_20578,N_23923);
and U24322 (N_24322,N_18298,N_19166);
and U24323 (N_24323,N_23531,N_23650);
or U24324 (N_24324,N_20036,N_22873);
and U24325 (N_24325,N_18557,N_18783);
xor U24326 (N_24326,N_22680,N_18051);
and U24327 (N_24327,N_18009,N_22729);
xnor U24328 (N_24328,N_18036,N_18541);
or U24329 (N_24329,N_20523,N_19787);
nand U24330 (N_24330,N_19824,N_22842);
xor U24331 (N_24331,N_19964,N_18829);
or U24332 (N_24332,N_20482,N_21279);
nand U24333 (N_24333,N_20690,N_21137);
nor U24334 (N_24334,N_21207,N_23579);
nor U24335 (N_24335,N_22541,N_23993);
nand U24336 (N_24336,N_18416,N_18588);
or U24337 (N_24337,N_19277,N_19452);
or U24338 (N_24338,N_20238,N_20641);
nand U24339 (N_24339,N_21661,N_20885);
xor U24340 (N_24340,N_19417,N_23750);
xnor U24341 (N_24341,N_20593,N_21002);
nor U24342 (N_24342,N_21760,N_23294);
and U24343 (N_24343,N_21763,N_19118);
xor U24344 (N_24344,N_21808,N_18668);
nand U24345 (N_24345,N_18037,N_21988);
xnor U24346 (N_24346,N_20125,N_21816);
nor U24347 (N_24347,N_20734,N_23140);
and U24348 (N_24348,N_20673,N_20302);
and U24349 (N_24349,N_18280,N_20580);
nor U24350 (N_24350,N_18116,N_20576);
and U24351 (N_24351,N_22693,N_20710);
nand U24352 (N_24352,N_18844,N_19387);
nor U24353 (N_24353,N_18300,N_21026);
and U24354 (N_24354,N_23649,N_19577);
nand U24355 (N_24355,N_20524,N_23189);
xor U24356 (N_24356,N_21922,N_22857);
or U24357 (N_24357,N_19111,N_21670);
or U24358 (N_24358,N_20368,N_18956);
and U24359 (N_24359,N_22464,N_23346);
and U24360 (N_24360,N_23476,N_22298);
and U24361 (N_24361,N_20373,N_23063);
nand U24362 (N_24362,N_22974,N_19773);
nand U24363 (N_24363,N_21874,N_21704);
nor U24364 (N_24364,N_23793,N_23932);
nor U24365 (N_24365,N_21148,N_19278);
or U24366 (N_24366,N_19428,N_19944);
nand U24367 (N_24367,N_19229,N_22940);
or U24368 (N_24368,N_19939,N_18318);
and U24369 (N_24369,N_19952,N_22175);
xnor U24370 (N_24370,N_19446,N_22887);
nor U24371 (N_24371,N_23706,N_19855);
and U24372 (N_24372,N_19354,N_22564);
or U24373 (N_24373,N_19703,N_22476);
nor U24374 (N_24374,N_18968,N_19222);
or U24375 (N_24375,N_19209,N_23773);
nor U24376 (N_24376,N_20300,N_21153);
and U24377 (N_24377,N_20460,N_20720);
nand U24378 (N_24378,N_22212,N_23146);
and U24379 (N_24379,N_22208,N_20413);
xnor U24380 (N_24380,N_23316,N_20084);
nand U24381 (N_24381,N_21954,N_23256);
and U24382 (N_24382,N_23099,N_19733);
or U24383 (N_24383,N_19079,N_22599);
nor U24384 (N_24384,N_21130,N_20972);
xor U24385 (N_24385,N_19433,N_18703);
nor U24386 (N_24386,N_22995,N_21594);
or U24387 (N_24387,N_21999,N_20602);
nor U24388 (N_24388,N_19987,N_23863);
or U24389 (N_24389,N_22168,N_22271);
and U24390 (N_24390,N_19378,N_21528);
xor U24391 (N_24391,N_21174,N_23241);
nor U24392 (N_24392,N_18991,N_19575);
or U24393 (N_24393,N_21536,N_21864);
nand U24394 (N_24394,N_21030,N_23934);
xor U24395 (N_24395,N_23956,N_18907);
nand U24396 (N_24396,N_18169,N_19757);
and U24397 (N_24397,N_23718,N_18281);
nor U24398 (N_24398,N_23756,N_18835);
nor U24399 (N_24399,N_22000,N_22067);
nand U24400 (N_24400,N_22353,N_19693);
nand U24401 (N_24401,N_18639,N_22459);
nand U24402 (N_24402,N_23755,N_18955);
xnor U24403 (N_24403,N_22674,N_18381);
nor U24404 (N_24404,N_23760,N_19335);
or U24405 (N_24405,N_22707,N_20615);
nand U24406 (N_24406,N_23553,N_21010);
and U24407 (N_24407,N_22415,N_20687);
or U24408 (N_24408,N_22832,N_18660);
and U24409 (N_24409,N_18149,N_23632);
or U24410 (N_24410,N_19257,N_22587);
nand U24411 (N_24411,N_22756,N_23047);
and U24412 (N_24412,N_22477,N_22640);
and U24413 (N_24413,N_23965,N_21278);
nor U24414 (N_24414,N_21394,N_23266);
and U24415 (N_24415,N_19927,N_19726);
or U24416 (N_24416,N_18591,N_22665);
and U24417 (N_24417,N_23858,N_22418);
or U24418 (N_24418,N_18705,N_19313);
nand U24419 (N_24419,N_20564,N_21520);
nand U24420 (N_24420,N_18752,N_22130);
xnor U24421 (N_24421,N_18847,N_19512);
nand U24422 (N_24422,N_23143,N_23674);
xor U24423 (N_24423,N_21336,N_23472);
nand U24424 (N_24424,N_19743,N_20181);
nor U24425 (N_24425,N_20528,N_19652);
and U24426 (N_24426,N_22058,N_23853);
nand U24427 (N_24427,N_18412,N_20063);
or U24428 (N_24428,N_21154,N_18739);
xor U24429 (N_24429,N_22008,N_19104);
and U24430 (N_24430,N_20475,N_18082);
or U24431 (N_24431,N_21800,N_22216);
xnor U24432 (N_24432,N_23901,N_22827);
or U24433 (N_24433,N_23440,N_18960);
nor U24434 (N_24434,N_19907,N_20903);
or U24435 (N_24435,N_20062,N_19766);
nand U24436 (N_24436,N_21473,N_19567);
and U24437 (N_24437,N_19346,N_21577);
or U24438 (N_24438,N_18105,N_21756);
and U24439 (N_24439,N_23407,N_22539);
nor U24440 (N_24440,N_22400,N_19617);
nor U24441 (N_24441,N_21141,N_23889);
nand U24442 (N_24442,N_19975,N_23051);
nand U24443 (N_24443,N_19688,N_21869);
nor U24444 (N_24444,N_21146,N_20866);
nand U24445 (N_24445,N_22527,N_20553);
nand U24446 (N_24446,N_21560,N_23208);
xnor U24447 (N_24447,N_21352,N_20497);
and U24448 (N_24448,N_20086,N_21879);
nand U24449 (N_24449,N_19546,N_19650);
nand U24450 (N_24450,N_22188,N_21291);
xnor U24451 (N_24451,N_22554,N_18294);
nand U24452 (N_24452,N_20304,N_22151);
or U24453 (N_24453,N_21268,N_20261);
and U24454 (N_24454,N_19906,N_18967);
nand U24455 (N_24455,N_19936,N_20134);
nand U24456 (N_24456,N_22147,N_22880);
nand U24457 (N_24457,N_22278,N_23111);
nor U24458 (N_24458,N_19938,N_23061);
xnor U24459 (N_24459,N_18124,N_18632);
xnor U24460 (N_24460,N_22746,N_20483);
xnor U24461 (N_24461,N_22772,N_23939);
xnor U24462 (N_24462,N_23318,N_22976);
nor U24463 (N_24463,N_19828,N_22871);
or U24464 (N_24464,N_18797,N_18028);
nor U24465 (N_24465,N_22144,N_21178);
nor U24466 (N_24466,N_21327,N_19897);
and U24467 (N_24467,N_23037,N_23005);
and U24468 (N_24468,N_20293,N_18794);
nor U24469 (N_24469,N_22059,N_19947);
nand U24470 (N_24470,N_22908,N_19422);
nand U24471 (N_24471,N_23097,N_20761);
nand U24472 (N_24472,N_21512,N_21083);
nor U24473 (N_24473,N_21555,N_22797);
nand U24474 (N_24474,N_23510,N_20241);
nor U24475 (N_24475,N_22856,N_20379);
or U24476 (N_24476,N_21945,N_22710);
or U24477 (N_24477,N_19409,N_22011);
or U24478 (N_24478,N_19343,N_21616);
nor U24479 (N_24479,N_20471,N_21576);
or U24480 (N_24480,N_20585,N_23852);
or U24481 (N_24481,N_23971,N_22193);
or U24482 (N_24482,N_19517,N_20779);
nor U24483 (N_24483,N_23721,N_20223);
and U24484 (N_24484,N_22048,N_22935);
xnor U24485 (N_24485,N_23573,N_21253);
xor U24486 (N_24486,N_19056,N_23045);
and U24487 (N_24487,N_19322,N_22927);
nand U24488 (N_24488,N_19144,N_18619);
and U24489 (N_24489,N_21194,N_23383);
and U24490 (N_24490,N_21687,N_21903);
and U24491 (N_24491,N_18987,N_22219);
nand U24492 (N_24492,N_20870,N_19673);
and U24493 (N_24493,N_23436,N_22548);
nor U24494 (N_24494,N_18862,N_21612);
nor U24495 (N_24495,N_18303,N_23640);
nor U24496 (N_24496,N_18019,N_19327);
or U24497 (N_24497,N_18361,N_23360);
nor U24498 (N_24498,N_19754,N_23693);
nand U24499 (N_24499,N_18133,N_23996);
or U24500 (N_24500,N_19469,N_23575);
nor U24501 (N_24501,N_18144,N_23794);
xnor U24502 (N_24502,N_19549,N_20057);
nor U24503 (N_24503,N_20993,N_20994);
and U24504 (N_24504,N_20457,N_21489);
nand U24505 (N_24505,N_20701,N_19527);
xnor U24506 (N_24506,N_22178,N_19072);
or U24507 (N_24507,N_18047,N_21039);
xnor U24508 (N_24508,N_20224,N_18267);
nor U24509 (N_24509,N_18200,N_21613);
and U24510 (N_24510,N_21109,N_20510);
nor U24511 (N_24511,N_18701,N_21640);
or U24512 (N_24512,N_22941,N_22289);
xor U24513 (N_24513,N_23079,N_23347);
nand U24514 (N_24514,N_22266,N_22057);
nor U24515 (N_24515,N_19402,N_22167);
nand U24516 (N_24516,N_23526,N_19788);
nor U24517 (N_24517,N_18544,N_22456);
xor U24518 (N_24518,N_20319,N_20680);
and U24519 (N_24519,N_23062,N_18382);
nand U24520 (N_24520,N_19138,N_23808);
and U24521 (N_24521,N_21308,N_22973);
nor U24522 (N_24522,N_19735,N_18138);
and U24523 (N_24523,N_18838,N_23055);
xnor U24524 (N_24524,N_20548,N_22645);
nand U24525 (N_24525,N_21688,N_20237);
and U24526 (N_24526,N_22198,N_22894);
or U24527 (N_24527,N_19901,N_23418);
and U24528 (N_24528,N_19813,N_20449);
or U24529 (N_24529,N_23136,N_23364);
nand U24530 (N_24530,N_18623,N_19214);
nor U24531 (N_24531,N_20746,N_20765);
nand U24532 (N_24532,N_19800,N_18236);
and U24533 (N_24533,N_23622,N_20631);
and U24534 (N_24534,N_18614,N_21388);
nor U24535 (N_24535,N_22512,N_18002);
xor U24536 (N_24536,N_18362,N_22405);
nor U24537 (N_24537,N_20740,N_19894);
and U24538 (N_24538,N_22959,N_18095);
and U24539 (N_24539,N_23142,N_23795);
nor U24540 (N_24540,N_19488,N_21605);
or U24541 (N_24541,N_21674,N_18503);
nand U24542 (N_24542,N_23715,N_19934);
xor U24543 (N_24543,N_21254,N_21454);
nor U24544 (N_24544,N_22322,N_19823);
nor U24545 (N_24545,N_22853,N_18872);
nor U24546 (N_24546,N_19564,N_21581);
or U24547 (N_24547,N_22916,N_21288);
xnor U24548 (N_24548,N_20742,N_21744);
nand U24549 (N_24549,N_22958,N_23928);
and U24550 (N_24550,N_19694,N_19371);
xnor U24551 (N_24551,N_23955,N_20852);
or U24552 (N_24552,N_20094,N_21669);
nand U24553 (N_24553,N_21751,N_20682);
nor U24554 (N_24554,N_23565,N_19251);
nor U24555 (N_24555,N_19720,N_21914);
and U24556 (N_24556,N_21490,N_19745);
or U24557 (N_24557,N_21691,N_20211);
or U24558 (N_24558,N_23204,N_18000);
xnor U24559 (N_24559,N_22540,N_20928);
xor U24560 (N_24560,N_20462,N_18433);
xor U24561 (N_24561,N_21609,N_22448);
nand U24562 (N_24562,N_23771,N_22076);
and U24563 (N_24563,N_22660,N_23157);
or U24564 (N_24564,N_23512,N_20842);
xnor U24565 (N_24565,N_23677,N_18888);
xor U24566 (N_24566,N_18065,N_20480);
or U24567 (N_24567,N_23303,N_22877);
nor U24568 (N_24568,N_23524,N_22287);
nand U24569 (N_24569,N_20328,N_18949);
nor U24570 (N_24570,N_18291,N_19731);
and U24571 (N_24571,N_18923,N_20542);
or U24572 (N_24572,N_18237,N_19027);
xnor U24573 (N_24573,N_22678,N_22028);
and U24574 (N_24574,N_20954,N_19296);
and U24575 (N_24575,N_21641,N_18851);
xnor U24576 (N_24576,N_23709,N_20512);
nand U24577 (N_24577,N_22581,N_22926);
or U24578 (N_24578,N_22806,N_19030);
nand U24579 (N_24579,N_22751,N_18641);
and U24580 (N_24580,N_20958,N_18998);
and U24581 (N_24581,N_18532,N_18288);
and U24582 (N_24582,N_20889,N_18785);
xnor U24583 (N_24583,N_23020,N_23172);
and U24584 (N_24584,N_19381,N_19356);
or U24585 (N_24585,N_19958,N_19969);
xor U24586 (N_24586,N_23549,N_18523);
xnor U24587 (N_24587,N_22864,N_22071);
nor U24588 (N_24588,N_18488,N_23197);
or U24589 (N_24589,N_18604,N_23710);
nor U24590 (N_24590,N_21305,N_23717);
nor U24591 (N_24591,N_18542,N_19641);
nand U24592 (N_24592,N_22225,N_22702);
and U24593 (N_24593,N_22563,N_19290);
xor U24594 (N_24594,N_19196,N_21619);
nor U24595 (N_24595,N_23240,N_23209);
nor U24596 (N_24596,N_20886,N_20395);
and U24597 (N_24597,N_22442,N_22851);
and U24598 (N_24598,N_23551,N_23326);
nand U24599 (N_24599,N_19383,N_18883);
or U24600 (N_24600,N_21953,N_19495);
xor U24601 (N_24601,N_18399,N_23597);
xor U24602 (N_24602,N_18612,N_21856);
and U24603 (N_24603,N_21203,N_18304);
nand U24604 (N_24604,N_23814,N_22490);
and U24605 (N_24605,N_23548,N_18066);
nand U24606 (N_24606,N_23212,N_19341);
xnor U24607 (N_24607,N_22249,N_19047);
or U24608 (N_24608,N_19796,N_23008);
nor U24609 (N_24609,N_22064,N_18522);
nor U24610 (N_24610,N_20828,N_20611);
nand U24611 (N_24611,N_19183,N_19014);
and U24612 (N_24612,N_18409,N_23738);
nand U24613 (N_24613,N_19004,N_21079);
xor U24614 (N_24614,N_22118,N_19247);
or U24615 (N_24615,N_20569,N_20822);
nand U24616 (N_24616,N_23690,N_23339);
nor U24617 (N_24617,N_22132,N_21876);
and U24618 (N_24618,N_19083,N_22319);
nand U24619 (N_24619,N_22482,N_23986);
nand U24620 (N_24620,N_22356,N_20521);
xnor U24621 (N_24621,N_23113,N_18781);
nand U24622 (N_24622,N_19344,N_22605);
and U24623 (N_24623,N_21558,N_21689);
nand U24624 (N_24624,N_20074,N_22060);
nor U24625 (N_24625,N_21739,N_22273);
nor U24626 (N_24626,N_19254,N_19419);
nor U24627 (N_24627,N_23520,N_19403);
nor U24628 (N_24628,N_21015,N_18606);
nor U24629 (N_24629,N_22001,N_22882);
nand U24630 (N_24630,N_21031,N_18269);
nand U24631 (N_24631,N_21273,N_18404);
or U24632 (N_24632,N_23454,N_23242);
xor U24633 (N_24633,N_22555,N_21233);
xor U24634 (N_24634,N_18808,N_19922);
nand U24635 (N_24635,N_18338,N_22732);
nor U24636 (N_24636,N_23628,N_20323);
xor U24637 (N_24637,N_19810,N_21565);
nor U24638 (N_24638,N_20884,N_22164);
and U24639 (N_24639,N_20799,N_20509);
and U24640 (N_24640,N_18094,N_20603);
xor U24641 (N_24641,N_18181,N_20169);
xnor U24642 (N_24642,N_22211,N_19563);
nor U24643 (N_24643,N_18762,N_20149);
nor U24644 (N_24644,N_21198,N_19168);
or U24645 (N_24645,N_22589,N_21684);
and U24646 (N_24646,N_22371,N_19920);
and U24647 (N_24647,N_22106,N_20549);
or U24648 (N_24648,N_22324,N_19099);
nand U24649 (N_24649,N_21877,N_19843);
nand U24650 (N_24650,N_18771,N_23660);
or U24651 (N_24651,N_23539,N_21431);
and U24652 (N_24652,N_20122,N_19259);
nor U24653 (N_24653,N_20451,N_19242);
or U24654 (N_24654,N_20252,N_18620);
nand U24655 (N_24655,N_23160,N_20590);
nor U24656 (N_24656,N_18995,N_21480);
nand U24657 (N_24657,N_18487,N_19521);
or U24658 (N_24658,N_19986,N_22687);
and U24659 (N_24659,N_23624,N_19230);
or U24660 (N_24660,N_19677,N_19737);
or U24661 (N_24661,N_18822,N_18437);
or U24662 (N_24662,N_18953,N_20203);
and U24663 (N_24663,N_18786,N_18110);
xor U24664 (N_24664,N_20649,N_21283);
or U24665 (N_24665,N_21965,N_19946);
or U24666 (N_24666,N_19280,N_18505);
xor U24667 (N_24667,N_19561,N_18092);
nand U24668 (N_24668,N_22828,N_22288);
or U24669 (N_24669,N_23931,N_19298);
and U24670 (N_24670,N_18245,N_18857);
xnor U24671 (N_24671,N_22643,N_21644);
nor U24672 (N_24672,N_18768,N_18539);
or U24673 (N_24673,N_23135,N_22265);
and U24674 (N_24674,N_20545,N_22480);
and U24675 (N_24675,N_20168,N_20144);
nor U24676 (N_24676,N_20515,N_23826);
and U24677 (N_24677,N_22836,N_20935);
nand U24678 (N_24678,N_20915,N_23777);
nor U24679 (N_24679,N_20289,N_23832);
nand U24680 (N_24680,N_19357,N_18563);
xor U24681 (N_24681,N_22899,N_19231);
xnor U24682 (N_24682,N_19244,N_22649);
nor U24683 (N_24683,N_19712,N_18759);
xor U24684 (N_24684,N_22432,N_18478);
nor U24685 (N_24685,N_21255,N_20277);
and U24686 (N_24686,N_19749,N_23787);
and U24687 (N_24687,N_18410,N_22103);
and U24688 (N_24688,N_22788,N_21711);
nand U24689 (N_24689,N_20032,N_23498);
xor U24690 (N_24690,N_18850,N_18372);
and U24691 (N_24691,N_21867,N_21709);
or U24692 (N_24692,N_20936,N_20435);
xnor U24693 (N_24693,N_20706,N_22458);
nor U24694 (N_24694,N_20025,N_19880);
nor U24695 (N_24695,N_20020,N_18787);
and U24696 (N_24696,N_18164,N_23384);
and U24697 (N_24697,N_22054,N_18913);
nand U24698 (N_24698,N_19498,N_20909);
nand U24699 (N_24699,N_23410,N_19910);
xnor U24700 (N_24700,N_22213,N_23257);
xor U24701 (N_24701,N_18994,N_19202);
nor U24702 (N_24702,N_19902,N_19995);
or U24703 (N_24703,N_21964,N_20782);
or U24704 (N_24704,N_20910,N_23458);
nor U24705 (N_24705,N_20448,N_21331);
xnor U24706 (N_24706,N_18622,N_23885);
nor U24707 (N_24707,N_22435,N_20106);
nor U24708 (N_24708,N_23824,N_22709);
nand U24709 (N_24709,N_22081,N_20583);
nand U24710 (N_24710,N_20320,N_19276);
nand U24711 (N_24711,N_19634,N_19315);
xnor U24712 (N_24712,N_23474,N_22497);
and U24713 (N_24713,N_19390,N_18875);
nand U24714 (N_24714,N_20249,N_18190);
xnor U24715 (N_24715,N_20301,N_21635);
nor U24716 (N_24716,N_23007,N_21446);
and U24717 (N_24717,N_20634,N_19817);
nor U24718 (N_24718,N_19831,N_22437);
and U24719 (N_24719,N_22431,N_20525);
nand U24720 (N_24720,N_23400,N_22195);
xor U24721 (N_24721,N_18599,N_19226);
nor U24722 (N_24722,N_23822,N_20638);
or U24723 (N_24723,N_19398,N_23781);
and U24724 (N_24724,N_22111,N_18966);
and U24725 (N_24725,N_19783,N_22777);
nor U24726 (N_24726,N_22594,N_22629);
nor U24727 (N_24727,N_20529,N_19046);
nor U24728 (N_24728,N_22395,N_18655);
or U24729 (N_24729,N_19614,N_18979);
nand U24730 (N_24730,N_21572,N_22812);
and U24731 (N_24731,N_19642,N_20427);
xor U24732 (N_24732,N_18993,N_23324);
nand U24733 (N_24733,N_22654,N_18976);
nand U24734 (N_24734,N_18766,N_19255);
xnor U24735 (N_24735,N_18407,N_21215);
xor U24736 (N_24736,N_22413,N_22492);
xnor U24737 (N_24737,N_18863,N_19779);
nor U24738 (N_24738,N_19394,N_20812);
or U24739 (N_24739,N_20479,N_20829);
nand U24740 (N_24740,N_21554,N_19983);
or U24741 (N_24741,N_23958,N_21210);
and U24742 (N_24742,N_20166,N_23884);
nor U24743 (N_24743,N_18898,N_23108);
or U24744 (N_24744,N_19618,N_23121);
or U24745 (N_24745,N_23536,N_21892);
or U24746 (N_24746,N_21552,N_22333);
nand U24747 (N_24747,N_18141,N_23225);
nand U24748 (N_24748,N_21959,N_18789);
and U24749 (N_24749,N_20040,N_18330);
nor U24750 (N_24750,N_21299,N_22263);
and U24751 (N_24751,N_19021,N_22809);
or U24752 (N_24752,N_22066,N_19534);
nor U24753 (N_24753,N_23789,N_18568);
and U24754 (N_24754,N_23999,N_23145);
nand U24755 (N_24755,N_20890,N_21774);
and U24756 (N_24756,N_22835,N_21873);
nor U24757 (N_24757,N_19438,N_20660);
nand U24758 (N_24758,N_18434,N_20982);
nand U24759 (N_24759,N_20679,N_21785);
nor U24760 (N_24760,N_23105,N_20654);
or U24761 (N_24761,N_18258,N_18214);
nor U24762 (N_24762,N_21620,N_19359);
xnor U24763 (N_24763,N_21220,N_22112);
nor U24764 (N_24764,N_23280,N_23653);
and U24765 (N_24765,N_23164,N_22024);
and U24766 (N_24766,N_22297,N_23026);
nand U24767 (N_24767,N_18447,N_21987);
xor U24768 (N_24768,N_21216,N_20003);
or U24769 (N_24769,N_18673,N_19848);
or U24770 (N_24770,N_19948,N_22795);
or U24771 (N_24771,N_23466,N_23406);
nand U24772 (N_24772,N_18840,N_21855);
and U24773 (N_24773,N_22755,N_20815);
xor U24774 (N_24774,N_23018,N_18904);
and U24775 (N_24775,N_23636,N_18948);
and U24776 (N_24776,N_21438,N_18615);
and U24777 (N_24777,N_21360,N_19878);
and U24778 (N_24778,N_20907,N_21981);
xnor U24779 (N_24779,N_22574,N_18411);
nand U24780 (N_24780,N_18154,N_18629);
nand U24781 (N_24781,N_21006,N_18020);
xor U24782 (N_24782,N_22051,N_19405);
and U24783 (N_24783,N_23408,N_20614);
or U24784 (N_24784,N_23405,N_18191);
or U24785 (N_24785,N_20531,N_23724);
and U24786 (N_24786,N_23229,N_22320);
or U24787 (N_24787,N_18546,N_20990);
nor U24788 (N_24788,N_19457,N_23540);
nand U24789 (N_24789,N_22931,N_19265);
nand U24790 (N_24790,N_19596,N_19109);
nand U24791 (N_24791,N_22838,N_21921);
nand U24792 (N_24792,N_19162,N_21199);
or U24793 (N_24793,N_19795,N_21589);
nor U24794 (N_24794,N_22822,N_21569);
nand U24795 (N_24795,N_18498,N_18353);
nor U24796 (N_24796,N_20061,N_21841);
nand U24797 (N_24797,N_18442,N_19937);
nand U24798 (N_24798,N_21177,N_18908);
nor U24799 (N_24799,N_19246,N_20179);
xnor U24800 (N_24800,N_22754,N_18643);
nor U24801 (N_24801,N_19139,N_23505);
or U24802 (N_24802,N_23605,N_22433);
and U24803 (N_24803,N_19633,N_22526);
xor U24804 (N_24804,N_22259,N_18286);
nand U24805 (N_24805,N_18724,N_22805);
nor U24806 (N_24806,N_22692,N_18270);
nor U24807 (N_24807,N_21306,N_20914);
and U24808 (N_24808,N_19124,N_23743);
nand U24809 (N_24809,N_23521,N_19929);
xnor U24810 (N_24810,N_19135,N_22642);
and U24811 (N_24811,N_18830,N_23295);
nand U24812 (N_24812,N_23868,N_18026);
or U24813 (N_24813,N_19369,N_20830);
xor U24814 (N_24814,N_21502,N_21321);
or U24815 (N_24815,N_22775,N_21518);
xnor U24816 (N_24816,N_23022,N_22598);
nand U24817 (N_24817,N_22698,N_22942);
or U24818 (N_24818,N_18091,N_19340);
nor U24819 (N_24819,N_20572,N_19185);
nand U24820 (N_24820,N_20739,N_22385);
or U24821 (N_24821,N_19701,N_20681);
and U24822 (N_24822,N_20239,N_20622);
nor U24823 (N_24823,N_23664,N_23535);
xor U24824 (N_24824,N_22349,N_23613);
nor U24825 (N_24825,N_19233,N_22447);
nor U24826 (N_24826,N_23453,N_22733);
and U24827 (N_24827,N_21386,N_18990);
or U24828 (N_24828,N_18530,N_23184);
or U24829 (N_24829,N_22372,N_22648);
nor U24830 (N_24830,N_23670,N_20834);
nor U24831 (N_24831,N_22810,N_18265);
and U24832 (N_24832,N_21843,N_23404);
nor U24833 (N_24833,N_23667,N_22773);
or U24834 (N_24834,N_23966,N_19833);
or U24835 (N_24835,N_20316,N_20022);
nand U24836 (N_24836,N_22327,N_19443);
or U24837 (N_24837,N_21337,N_20816);
or U24838 (N_24838,N_20766,N_21870);
xnor U24839 (N_24839,N_19220,N_22070);
xor U24840 (N_24840,N_19449,N_22215);
xor U24841 (N_24841,N_19500,N_22830);
xor U24842 (N_24842,N_21018,N_21912);
nor U24843 (N_24843,N_18031,N_21320);
xor U24844 (N_24844,N_18360,N_23412);
xor U24845 (N_24845,N_21980,N_18517);
and U24846 (N_24846,N_23447,N_21853);
or U24847 (N_24847,N_18753,N_23442);
nor U24848 (N_24848,N_22380,N_20973);
xnor U24849 (N_24849,N_22879,N_18575);
nand U24850 (N_24850,N_23477,N_18355);
or U24851 (N_24851,N_19334,N_23591);
nand U24852 (N_24852,N_18793,N_21375);
xor U24853 (N_24853,N_18556,N_20048);
nand U24854 (N_24854,N_19052,N_21344);
and U24855 (N_24855,N_19557,N_20400);
nand U24856 (N_24856,N_23288,N_23954);
and U24857 (N_24857,N_18645,N_22359);
and U24858 (N_24858,N_19216,N_18230);
and U24859 (N_24859,N_21531,N_22831);
or U24860 (N_24860,N_22161,N_18038);
nand U24861 (N_24861,N_19291,N_20441);
and U24862 (N_24862,N_23094,N_19623);
xnor U24863 (N_24863,N_20332,N_22870);
nand U24864 (N_24864,N_20132,N_18957);
nand U24865 (N_24865,N_18130,N_21878);
and U24866 (N_24866,N_21736,N_19068);
or U24867 (N_24867,N_22393,N_23530);
or U24868 (N_24868,N_20431,N_23092);
nand U24869 (N_24869,N_23200,N_20735);
nand U24870 (N_24870,N_23123,N_18698);
nor U24871 (N_24871,N_19489,N_18740);
and U24872 (N_24872,N_18597,N_19116);
nand U24873 (N_24873,N_22614,N_18590);
and U24874 (N_24874,N_21172,N_20212);
xor U24875 (N_24875,N_22294,N_19130);
and U24876 (N_24876,N_23190,N_23844);
xnor U24877 (N_24877,N_22468,N_23534);
xor U24878 (N_24878,N_20468,N_18930);
nor U24879 (N_24879,N_19999,N_21896);
or U24880 (N_24880,N_18895,N_22409);
or U24881 (N_24881,N_19096,N_20843);
nand U24882 (N_24882,N_22966,N_19272);
and U24883 (N_24883,N_21755,N_21598);
xnor U24884 (N_24884,N_21460,N_18909);
xnor U24885 (N_24885,N_18610,N_20727);
xor U24886 (N_24886,N_20143,N_23462);
or U24887 (N_24887,N_19651,N_23054);
or U24888 (N_24888,N_18950,N_21144);
nand U24889 (N_24889,N_21511,N_22399);
nor U24890 (N_24890,N_19974,N_18369);
and U24891 (N_24891,N_20156,N_20285);
nand U24892 (N_24892,N_22117,N_20689);
xnor U24893 (N_24893,N_23065,N_20097);
nand U24894 (N_24894,N_18254,N_22052);
nor U24895 (N_24895,N_21606,N_19739);
or U24896 (N_24896,N_23118,N_19486);
xor U24897 (N_24897,N_22428,N_19637);
nand U24898 (N_24898,N_19805,N_19856);
nor U24899 (N_24899,N_18016,N_18397);
and U24900 (N_24900,N_19511,N_18746);
nand U24901 (N_24901,N_19080,N_20651);
nor U24902 (N_24902,N_19425,N_22509);
xor U24903 (N_24903,N_20488,N_18694);
xor U24904 (N_24904,N_19898,N_22462);
nor U24905 (N_24905,N_22233,N_18594);
nor U24906 (N_24906,N_21356,N_22933);
nor U24907 (N_24907,N_19044,N_18374);
nor U24908 (N_24908,N_21000,N_21947);
xor U24909 (N_24909,N_19106,N_19933);
xor U24910 (N_24910,N_20174,N_21722);
and U24911 (N_24911,N_21436,N_22784);
nor U24912 (N_24912,N_18259,N_20872);
or U24913 (N_24913,N_22823,N_18760);
xor U24914 (N_24914,N_20317,N_22173);
and U24915 (N_24915,N_19156,N_19911);
xor U24916 (N_24916,N_23112,N_21986);
or U24917 (N_24917,N_20056,N_20947);
and U24918 (N_24918,N_21643,N_23301);
nand U24919 (N_24919,N_18805,N_20217);
xor U24920 (N_24920,N_18185,N_19374);
and U24921 (N_24921,N_21269,N_19355);
xor U24922 (N_24922,N_19537,N_20718);
or U24923 (N_24923,N_20762,N_22819);
xnor U24924 (N_24924,N_21807,N_18261);
and U24925 (N_24925,N_21909,N_19647);
and U24926 (N_24926,N_21835,N_21668);
or U24927 (N_24927,N_22484,N_18551);
or U24928 (N_24928,N_22685,N_19212);
and U24929 (N_24929,N_19376,N_23612);
xor U24930 (N_24930,N_23561,N_20219);
nand U24931 (N_24931,N_23847,N_20721);
xnor U24932 (N_24932,N_22030,N_18633);
nand U24933 (N_24933,N_18638,N_19655);
and U24934 (N_24934,N_22218,N_18881);
nor U24935 (N_24935,N_23273,N_21710);
nand U24936 (N_24936,N_23416,N_20209);
or U24937 (N_24937,N_19529,N_21088);
nand U24938 (N_24938,N_22583,N_21100);
or U24939 (N_24939,N_21152,N_19045);
and U24940 (N_24940,N_21888,N_19613);
or U24941 (N_24941,N_21459,N_22505);
and U24942 (N_24942,N_21099,N_19472);
or U24943 (N_24943,N_21094,N_21333);
and U24944 (N_24944,N_23004,N_19738);
xnor U24945 (N_24945,N_21678,N_20946);
nand U24946 (N_24946,N_21082,N_20117);
and U24947 (N_24947,N_18721,N_18126);
nand U24948 (N_24948,N_19719,N_23704);
and U24949 (N_24949,N_21453,N_18674);
or U24950 (N_24950,N_19636,N_23585);
and U24951 (N_24951,N_23414,N_18242);
and U24952 (N_24952,N_19262,N_19362);
xnor U24953 (N_24953,N_21549,N_21452);
nand U24954 (N_24954,N_19232,N_19967);
nand U24955 (N_24955,N_19811,N_20359);
or U24956 (N_24956,N_19161,N_19465);
xnor U24957 (N_24957,N_18217,N_19715);
and U24958 (N_24958,N_21673,N_21239);
nor U24959 (N_24959,N_20986,N_19925);
and U24960 (N_24960,N_18801,N_21839);
or U24961 (N_24961,N_23362,N_20342);
or U24962 (N_24962,N_20102,N_22790);
or U24963 (N_24963,N_20330,N_23644);
or U24964 (N_24964,N_20005,N_19790);
nand U24965 (N_24965,N_20733,N_19953);
nand U24966 (N_24966,N_22985,N_21919);
nor U24967 (N_24967,N_20409,N_18435);
nand U24968 (N_24968,N_22975,N_19120);
and U24969 (N_24969,N_22796,N_19710);
or U24970 (N_24970,N_18711,N_22672);
xor U24971 (N_24971,N_22750,N_23003);
or U24972 (N_24972,N_20952,N_18459);
and U24973 (N_24973,N_19463,N_20398);
xnor U24974 (N_24974,N_20906,N_23421);
nor U24975 (N_24975,N_18500,N_21441);
nor U24976 (N_24976,N_18042,N_20831);
xor U24977 (N_24977,N_18662,N_18656);
nor U24978 (N_24978,N_20640,N_19031);
or U24979 (N_24979,N_19602,N_20308);
nand U24980 (N_24980,N_21049,N_20623);
nor U24981 (N_24981,N_22165,N_19293);
or U24982 (N_24982,N_23871,N_19799);
or U24983 (N_24983,N_22108,N_23668);
nor U24984 (N_24984,N_18107,N_21252);
nand U24985 (N_24985,N_19364,N_22172);
and U24986 (N_24986,N_19006,N_19358);
xor U24987 (N_24987,N_21391,N_23839);
nor U24988 (N_24988,N_22160,N_20808);
nor U24989 (N_24989,N_22872,N_19971);
nor U24990 (N_24990,N_21979,N_18417);
xnor U24991 (N_24991,N_20789,N_21672);
xor U24992 (N_24992,N_19885,N_18582);
or U24993 (N_24993,N_20450,N_21370);
and U24994 (N_24994,N_23739,N_23067);
nor U24995 (N_24995,N_21570,N_19576);
nor U24996 (N_24996,N_22282,N_20714);
nand U24997 (N_24997,N_22135,N_23835);
nor U24998 (N_24998,N_18550,N_19875);
xor U24999 (N_24999,N_20595,N_19681);
xor U25000 (N_25000,N_21267,N_22032);
nand U25001 (N_25001,N_18394,N_22595);
or U25002 (N_25002,N_22360,N_18081);
and U25003 (N_25003,N_22516,N_23050);
nor U25004 (N_25004,N_21161,N_23596);
and U25005 (N_25005,N_22960,N_22006);
and U25006 (N_25006,N_21218,N_20055);
xnor U25007 (N_25007,N_19912,N_22651);
or U25008 (N_25008,N_18723,N_21804);
xor U25009 (N_25009,N_21093,N_20412);
and U25010 (N_25010,N_20183,N_22867);
and U25011 (N_25011,N_19342,N_21445);
xnor U25012 (N_25012,N_23911,N_20443);
and U25013 (N_25013,N_23349,N_22712);
nand U25014 (N_25014,N_20671,N_18681);
xor U25015 (N_25015,N_20096,N_21089);
nand U25016 (N_25016,N_21374,N_23203);
xor U25017 (N_25017,N_18516,N_23378);
nor U25018 (N_25018,N_22900,N_18569);
nand U25019 (N_25019,N_22936,N_20015);
xnor U25020 (N_25020,N_21195,N_20180);
xor U25021 (N_25021,N_18699,N_19672);
or U25022 (N_25022,N_20393,N_18139);
and U25023 (N_25023,N_19666,N_21139);
and U25024 (N_25024,N_21264,N_21399);
or U25025 (N_25025,N_19905,N_22015);
and U25026 (N_25026,N_23550,N_22283);
nor U25027 (N_25027,N_18370,N_21765);
or U25028 (N_25028,N_21044,N_22731);
nor U25029 (N_25029,N_20140,N_21545);
nand U25030 (N_25030,N_19101,N_18148);
nor U25031 (N_25031,N_23239,N_22079);
xor U25032 (N_25032,N_21962,N_19649);
or U25033 (N_25033,N_18686,N_19807);
xor U25034 (N_25034,N_21939,N_18772);
and U25035 (N_25035,N_20305,N_21596);
xnor U25036 (N_25036,N_23941,N_20290);
and U25037 (N_25037,N_20007,N_21716);
or U25038 (N_25038,N_21435,N_23627);
and U25039 (N_25039,N_19961,N_19319);
nor U25040 (N_25040,N_18172,N_19439);
and U25041 (N_25041,N_18376,N_21748);
or U25042 (N_25042,N_23352,N_18170);
or U25043 (N_25043,N_19329,N_18911);
nand U25044 (N_25044,N_21916,N_18710);
nand U25045 (N_25045,N_22677,N_23450);
nor U25046 (N_25046,N_18425,N_18325);
nor U25047 (N_25047,N_18166,N_18296);
and U25048 (N_25048,N_18131,N_20748);
nand U25049 (N_25049,N_21418,N_23260);
nor U25050 (N_25050,N_23635,N_18388);
nand U25051 (N_25051,N_21222,N_22267);
or U25052 (N_25052,N_18050,N_20609);
nand U25053 (N_25053,N_20744,N_18211);
nand U25054 (N_25054,N_22370,N_20489);
nor U25055 (N_25055,N_21211,N_18204);
xor U25056 (N_25056,N_20329,N_21261);
and U25057 (N_25057,N_23345,N_18893);
xor U25058 (N_25058,N_20275,N_19018);
xor U25059 (N_25059,N_22597,N_22097);
or U25060 (N_25060,N_18221,N_18560);
or U25061 (N_25061,N_22352,N_22256);
xnor U25062 (N_25062,N_22953,N_23921);
or U25063 (N_25063,N_22700,N_18039);
or U25064 (N_25064,N_20145,N_19133);
and U25065 (N_25065,N_19965,N_18238);
nand U25066 (N_25066,N_21380,N_19565);
or U25067 (N_25067,N_19077,N_22852);
and U25068 (N_25068,N_22274,N_21213);
or U25069 (N_25069,N_21250,N_18308);
nor U25070 (N_25070,N_22669,N_19399);
nand U25071 (N_25071,N_23330,N_19845);
and U25072 (N_25072,N_22078,N_22368);
and U25073 (N_25073,N_19763,N_20172);
nand U25074 (N_25074,N_22983,N_18894);
or U25075 (N_25075,N_22854,N_22793);
nand U25076 (N_25076,N_19945,N_21022);
nor U25077 (N_25077,N_19851,N_21341);
xnor U25078 (N_25078,N_21646,N_19325);
and U25079 (N_25079,N_18917,N_22514);
xor U25080 (N_25080,N_18810,N_19724);
xor U25081 (N_25081,N_18220,N_22699);
or U25082 (N_25082,N_23658,N_18260);
and U25083 (N_25083,N_22889,N_22450);
or U25084 (N_25084,N_21098,N_18223);
and U25085 (N_25085,N_20821,N_20150);
xor U25086 (N_25086,N_18680,N_23702);
nand U25087 (N_25087,N_18249,N_20047);
nor U25088 (N_25088,N_21393,N_21889);
or U25089 (N_25089,N_19264,N_22556);
nor U25090 (N_25090,N_21801,N_23896);
or U25091 (N_25091,N_23277,N_18900);
nand U25092 (N_25092,N_22620,N_20565);
xnor U25093 (N_25093,N_19705,N_18609);
nand U25094 (N_25094,N_22600,N_21802);
nor U25095 (N_25095,N_21196,N_22157);
nor U25096 (N_25096,N_18314,N_19832);
nand U25097 (N_25097,N_22416,N_22785);
or U25098 (N_25098,N_21131,N_23805);
xnor U25099 (N_25099,N_18846,N_18492);
nand U25100 (N_25100,N_20231,N_21806);
xor U25101 (N_25101,N_23995,N_20394);
or U25102 (N_25102,N_22502,N_21343);
and U25103 (N_25103,N_18471,N_20648);
or U25104 (N_25104,N_19857,N_18465);
or U25105 (N_25105,N_19943,N_23686);
xnor U25106 (N_25106,N_18363,N_22065);
nor U25107 (N_25107,N_19084,N_21593);
or U25108 (N_25108,N_20547,N_21420);
xor U25109 (N_25109,N_18043,N_18457);
nor U25110 (N_25110,N_20825,N_22229);
or U25111 (N_25111,N_18161,N_22309);
or U25112 (N_25112,N_21136,N_18985);
nand U25113 (N_25113,N_21692,N_22326);
nand U25114 (N_25114,N_20033,N_19887);
nor U25115 (N_25115,N_19653,N_20485);
xnor U25116 (N_25116,N_22174,N_18183);
nand U25117 (N_25117,N_19562,N_19454);
or U25118 (N_25118,N_22228,N_18534);
xor U25119 (N_25119,N_19620,N_23691);
and U25120 (N_25120,N_22630,N_23449);
xnor U25121 (N_25121,N_21582,N_23665);
nand U25122 (N_25122,N_19883,N_23963);
xor U25123 (N_25123,N_22042,N_20845);
nand U25124 (N_25124,N_21523,N_23485);
nand U25125 (N_25125,N_20049,N_20361);
and U25126 (N_25126,N_19931,N_22209);
xor U25127 (N_25127,N_22362,N_19012);
and U25128 (N_25128,N_23446,N_23304);
or U25129 (N_25129,N_19129,N_20182);
nand U25130 (N_25130,N_20668,N_22621);
and U25131 (N_25131,N_19697,N_23429);
nor U25132 (N_25132,N_19861,N_20708);
nor U25133 (N_25133,N_18415,N_23682);
or U25134 (N_25134,N_22592,N_21228);
nand U25135 (N_25135,N_22467,N_23042);
nand U25136 (N_25136,N_23875,N_22023);
nor U25137 (N_25137,N_20697,N_20655);
xnor U25138 (N_25138,N_18832,N_23465);
or U25139 (N_25139,N_22517,N_21633);
and U25140 (N_25140,N_22005,N_19895);
xnor U25141 (N_25141,N_22269,N_19434);
and U25142 (N_25142,N_20325,N_18229);
nor U25143 (N_25143,N_22083,N_23563);
and U25144 (N_25144,N_21725,N_22457);
or U25145 (N_25145,N_19043,N_18395);
xnor U25146 (N_25146,N_22863,N_20573);
nand U25147 (N_25147,N_22096,N_23181);
nand U25148 (N_25148,N_20123,N_18663);
nor U25149 (N_25149,N_23976,N_21607);
and U25150 (N_25150,N_18069,N_19846);
and U25151 (N_25151,N_22759,N_22911);
xnor U25152 (N_25152,N_23497,N_20164);
xnor U25153 (N_25153,N_23590,N_20254);
and U25154 (N_25154,N_19086,N_19601);
or U25155 (N_25155,N_19300,N_23035);
and U25156 (N_25156,N_22090,N_22813);
and U25157 (N_25157,N_19397,N_18078);
nor U25158 (N_25158,N_23363,N_18212);
nor U25159 (N_25159,N_22465,N_19727);
or U25160 (N_25160,N_23369,N_20796);
nand U25161 (N_25161,N_18243,N_21904);
nand U25162 (N_25162,N_22010,N_19103);
nand U25163 (N_25163,N_21121,N_21894);
nor U25164 (N_25164,N_19744,N_22036);
or U25165 (N_25165,N_19748,N_23424);
nor U25166 (N_25166,N_21471,N_22116);
nand U25167 (N_25167,N_20791,N_21232);
nand U25168 (N_25168,N_21538,N_22917);
nand U25169 (N_25169,N_20875,N_18773);
or U25170 (N_25170,N_23267,N_21603);
nor U25171 (N_25171,N_22744,N_18324);
nor U25172 (N_25172,N_23952,N_23130);
xnor U25173 (N_25173,N_23000,N_19692);
nor U25174 (N_25174,N_21241,N_23882);
and U25175 (N_25175,N_19218,N_22635);
xor U25176 (N_25176,N_21975,N_22137);
xor U25177 (N_25177,N_19471,N_21707);
or U25178 (N_25178,N_22199,N_20922);
or U25179 (N_25179,N_23984,N_22697);
nand U25180 (N_25180,N_23348,N_21016);
or U25181 (N_25181,N_21863,N_22138);
nor U25182 (N_25182,N_21023,N_20216);
nor U25183 (N_25183,N_23059,N_21024);
and U25184 (N_25184,N_18008,N_22929);
nor U25185 (N_25185,N_21860,N_20073);
nor U25186 (N_25186,N_21715,N_21926);
xor U25187 (N_25187,N_20632,N_19337);
or U25188 (N_25188,N_18439,N_23908);
nand U25189 (N_25189,N_21084,N_20838);
xor U25190 (N_25190,N_23325,N_18342);
or U25191 (N_25191,N_19784,N_22843);
or U25192 (N_25192,N_18173,N_21658);
nor U25193 (N_25193,N_21323,N_18055);
and U25194 (N_25194,N_23258,N_21467);
nand U25195 (N_25195,N_23639,N_19022);
nor U25196 (N_25196,N_18331,N_21048);
xor U25197 (N_25197,N_20037,N_20481);
xor U25198 (N_25198,N_19598,N_19571);
and U25199 (N_25199,N_19459,N_18611);
nor U25200 (N_25200,N_23705,N_18700);
nor U25201 (N_25201,N_23177,N_21315);
and U25202 (N_25202,N_20058,N_21231);
nand U25203 (N_25203,N_19466,N_18210);
nor U25204 (N_25204,N_21650,N_21184);
and U25205 (N_25205,N_23518,N_23989);
nor U25206 (N_25206,N_23245,N_22210);
or U25207 (N_25207,N_22303,N_22109);
nand U25208 (N_25208,N_18428,N_18970);
nor U25209 (N_25209,N_23804,N_20046);
and U25210 (N_25210,N_19863,N_19531);
nor U25211 (N_25211,N_22757,N_21395);
xnor U25212 (N_25212,N_20470,N_18943);
and U25213 (N_25213,N_18792,N_22343);
and U25214 (N_25214,N_20759,N_20941);
or U25215 (N_25215,N_20178,N_23662);
xor U25216 (N_25216,N_20192,N_18453);
xnor U25217 (N_25217,N_23169,N_21406);
and U25218 (N_25218,N_18978,N_22242);
xnor U25219 (N_25219,N_18306,N_22150);
and U25220 (N_25220,N_22460,N_22115);
or U25221 (N_25221,N_18393,N_23048);
nand U25222 (N_25222,N_19190,N_21893);
or U25223 (N_25223,N_19171,N_18932);
xnor U25224 (N_25224,N_23205,N_20743);
or U25225 (N_25225,N_23529,N_22420);
nand U25226 (N_25226,N_21474,N_18241);
nor U25227 (N_25227,N_23759,N_22551);
nor U25228 (N_25228,N_18777,N_20371);
nand U25229 (N_25229,N_18717,N_21951);
nor U25230 (N_25230,N_19415,N_23248);
and U25231 (N_25231,N_20945,N_20550);
or U25232 (N_25232,N_21470,N_18685);
nand U25233 (N_25233,N_21244,N_23566);
nor U25234 (N_25234,N_20724,N_22668);
xor U25235 (N_25235,N_19236,N_20053);
xor U25236 (N_25236,N_18552,N_19177);
or U25237 (N_25237,N_20490,N_18820);
and U25238 (N_25238,N_22667,N_23936);
or U25239 (N_25239,N_22579,N_21534);
xnor U25240 (N_25240,N_22650,N_23961);
or U25241 (N_25241,N_22367,N_20072);
and U25242 (N_25242,N_23514,N_22977);
nand U25243 (N_25243,N_21766,N_23802);
and U25244 (N_25244,N_22612,N_23066);
or U25245 (N_25245,N_19671,N_23633);
nor U25246 (N_25246,N_23616,N_18371);
xnor U25247 (N_25247,N_19181,N_21060);
nand U25248 (N_25248,N_21185,N_23120);
xor U25249 (N_25249,N_23182,N_23697);
xnor U25250 (N_25250,N_21591,N_21354);
or U25251 (N_25251,N_19385,N_19847);
nor U25252 (N_25252,N_23468,N_23831);
nand U25253 (N_25253,N_21586,N_22363);
or U25254 (N_25254,N_19956,N_18788);
nor U25255 (N_25255,N_20363,N_23967);
and U25256 (N_25256,N_19949,N_19260);
or U25257 (N_25257,N_20938,N_21971);
xnor U25258 (N_25258,N_19619,N_22547);
or U25259 (N_25259,N_20624,N_18558);
nand U25260 (N_25260,N_22314,N_21814);
and U25261 (N_25261,N_19581,N_22653);
nand U25262 (N_25262,N_23930,N_18774);
or U25263 (N_25263,N_22568,N_23305);
xor U25264 (N_25264,N_18476,N_21695);
or U25265 (N_25265,N_21257,N_23681);
and U25266 (N_25266,N_23168,N_23452);
and U25267 (N_25267,N_21068,N_21300);
xnor U25268 (N_25268,N_22250,N_20088);
and U25269 (N_25269,N_18891,N_19819);
xor U25270 (N_25270,N_23910,N_22609);
xnor U25271 (N_25271,N_18247,N_23907);
and U25272 (N_25272,N_22655,N_22683);
and U25273 (N_25273,N_23319,N_18063);
nand U25274 (N_25274,N_21587,N_19570);
xor U25275 (N_25275,N_19538,N_20588);
or U25276 (N_25276,N_20774,N_23153);
nor U25277 (N_25277,N_19430,N_23165);
and U25278 (N_25278,N_19566,N_23886);
nand U25279 (N_25279,N_23254,N_18601);
or U25280 (N_25280,N_19256,N_23872);
and U25281 (N_25281,N_18379,N_22239);
xor U25282 (N_25282,N_18821,N_20650);
nand U25283 (N_25283,N_22623,N_21557);
nor U25284 (N_25284,N_23766,N_21882);
nor U25285 (N_25285,N_22765,N_20598);
xnor U25286 (N_25286,N_20963,N_22171);
or U25287 (N_25287,N_20968,N_21217);
nor U25288 (N_25288,N_18049,N_23629);
xor U25289 (N_25289,N_21730,N_18337);
nand U25290 (N_25290,N_20341,N_19776);
nor U25291 (N_25291,N_20358,N_21550);
nand U25292 (N_25292,N_20075,N_23589);
and U25293 (N_25293,N_18696,N_19455);
xnor U25294 (N_25294,N_18803,N_19802);
xnor U25295 (N_25295,N_20913,N_23947);
xnor U25296 (N_25296,N_19972,N_22155);
xnor U25297 (N_25297,N_20292,N_21113);
and U25298 (N_25298,N_18984,N_21781);
nand U25299 (N_25299,N_18121,N_23043);
and U25300 (N_25300,N_21447,N_18658);
nor U25301 (N_25301,N_19635,N_21448);
nor U25302 (N_25302,N_23790,N_18384);
nor U25303 (N_25303,N_23475,N_18497);
and U25304 (N_25304,N_21602,N_23834);
nand U25305 (N_25305,N_23068,N_19900);
nand U25306 (N_25306,N_20197,N_20066);
nand U25307 (N_25307,N_23752,N_19991);
or U25308 (N_25308,N_23671,N_18951);
xnor U25309 (N_25309,N_21013,N_22850);
nand U25310 (N_25310,N_18884,N_23124);
and U25311 (N_25311,N_21108,N_20930);
nand U25312 (N_25312,N_20348,N_20248);
nor U25313 (N_25313,N_21034,N_19360);
xnor U25314 (N_25314,N_21052,N_22998);
nor U25315 (N_25315,N_20685,N_18046);
or U25316 (N_25316,N_20674,N_23659);
nor U25317 (N_25317,N_20709,N_22183);
and U25318 (N_25318,N_21797,N_22427);
nor U25319 (N_25319,N_19785,N_19923);
xor U25320 (N_25320,N_18827,N_18287);
and U25321 (N_25321,N_18177,N_21425);
xor U25322 (N_25322,N_23906,N_20594);
and U25323 (N_25323,N_23285,N_23186);
nor U25324 (N_25324,N_23110,N_22979);
and U25325 (N_25325,N_22376,N_20665);
or U25326 (N_25326,N_19051,N_20798);
and U25327 (N_25327,N_18853,N_23988);
or U25328 (N_25328,N_21826,N_18029);
xnor U25329 (N_25329,N_19332,N_20175);
xor U25330 (N_25330,N_22886,N_20737);
or U25331 (N_25331,N_20195,N_22606);
and U25332 (N_25332,N_19091,N_18791);
nand U25333 (N_25333,N_19395,N_21911);
and U25334 (N_25334,N_21150,N_18010);
or U25335 (N_25335,N_23385,N_22268);
or U25336 (N_25336,N_23464,N_23675);
xnor U25337 (N_25337,N_20728,N_21162);
nor U25338 (N_25338,N_19028,N_23461);
or U25339 (N_25339,N_21713,N_22166);
xor U25340 (N_25340,N_22073,N_21621);
nor U25341 (N_25341,N_20454,N_21384);
nor U25342 (N_25342,N_20347,N_23788);
and U25343 (N_25343,N_20111,N_22538);
or U25344 (N_25344,N_20855,N_18962);
nand U25345 (N_25345,N_21846,N_21101);
and U25346 (N_25346,N_22897,N_23292);
xnor U25347 (N_25347,N_21318,N_20444);
and U25348 (N_25348,N_22646,N_19224);
nor U25349 (N_25349,N_20811,N_21075);
nand U25350 (N_25350,N_19468,N_18340);
nor U25351 (N_25351,N_23058,N_23584);
or U25352 (N_25352,N_20362,N_18313);
nand U25353 (N_25353,N_21792,N_23887);
nor U25354 (N_25354,N_21293,N_20520);
nand U25355 (N_25355,N_21347,N_23281);
nand U25356 (N_25356,N_20503,N_22892);
nor U25357 (N_25357,N_23491,N_20240);
xor U25358 (N_25358,N_23552,N_18351);
nand U25359 (N_25359,N_19812,N_23342);
or U25360 (N_25360,N_19978,N_18179);
and U25361 (N_25361,N_18391,N_23626);
or U25362 (N_25362,N_20696,N_20355);
or U25363 (N_25363,N_22603,N_22496);
and U25364 (N_25364,N_20810,N_22452);
or U25365 (N_25365,N_18431,N_21499);
and U25366 (N_25366,N_19761,N_21115);
or U25367 (N_25367,N_23601,N_21553);
nand U25368 (N_25368,N_21905,N_20204);
or U25369 (N_25369,N_20064,N_21169);
or U25370 (N_25370,N_22417,N_18194);
and U25371 (N_25371,N_19314,N_18030);
nand U25372 (N_25372,N_22472,N_20635);
or U25373 (N_25373,N_19698,N_19508);
xor U25374 (N_25374,N_20424,N_19980);
or U25375 (N_25375,N_23133,N_20402);
nand U25376 (N_25376,N_20832,N_19207);
and U25377 (N_25377,N_18160,N_19203);
xor U25378 (N_25378,N_22817,N_21861);
xor U25379 (N_25379,N_23545,N_22493);
nand U25380 (N_25380,N_18458,N_23699);
xor U25381 (N_25381,N_18784,N_21584);
and U25382 (N_25382,N_18311,N_20824);
nor U25383 (N_25383,N_22344,N_20389);
xnor U25384 (N_25384,N_18356,N_18815);
or U25385 (N_25385,N_21200,N_18075);
and U25386 (N_25386,N_21522,N_20693);
xor U25387 (N_25387,N_21340,N_19839);
and U25388 (N_25388,N_19125,N_23011);
nand U25389 (N_25389,N_18617,N_19015);
nand U25390 (N_25390,N_23372,N_19973);
or U25391 (N_25391,N_18145,N_18722);
nor U25392 (N_25392,N_18099,N_22378);
and U25393 (N_25393,N_23555,N_20516);
or U25394 (N_25394,N_20158,N_20233);
nor U25395 (N_25395,N_23282,N_21891);
nand U25396 (N_25396,N_18227,N_18482);
nor U25397 (N_25397,N_22003,N_19427);
or U25398 (N_25398,N_23749,N_21599);
and U25399 (N_25399,N_18901,N_20445);
nand U25400 (N_25400,N_18683,N_21773);
and U25401 (N_25401,N_20784,N_18484);
nand U25402 (N_25402,N_18526,N_18664);
nor U25403 (N_25403,N_19134,N_20858);
and U25404 (N_25404,N_20295,N_20307);
or U25405 (N_25405,N_22895,N_20000);
nor U25406 (N_25406,N_18511,N_20664);
nor U25407 (N_25407,N_19184,N_21246);
nor U25408 (N_25408,N_21214,N_20496);
xnor U25409 (N_25409,N_19675,N_22018);
xnor U25410 (N_25410,N_18271,N_19483);
nor U25411 (N_25411,N_19215,N_20030);
xor U25412 (N_25412,N_21201,N_23701);
xor U25413 (N_25413,N_18945,N_18636);
nand U25414 (N_25414,N_21697,N_20692);
nand U25415 (N_25415,N_23577,N_21359);
nand U25416 (N_25416,N_23302,N_22224);
and U25417 (N_25417,N_20818,N_23334);
and U25418 (N_25418,N_22950,N_21884);
nor U25419 (N_25419,N_20021,N_23237);
xnor U25420 (N_25420,N_22719,N_21831);
and U25421 (N_25421,N_19437,N_23829);
and U25422 (N_25422,N_19269,N_22608);
xnor U25423 (N_25423,N_19844,N_22507);
xnor U25424 (N_25424,N_22829,N_19718);
xor U25425 (N_25425,N_21487,N_19587);
nand U25426 (N_25426,N_21983,N_21705);
nor U25427 (N_25427,N_20694,N_19211);
nor U25428 (N_25428,N_21338,N_18490);
and U25429 (N_25429,N_18897,N_20227);
nor U25430 (N_25430,N_20326,N_20902);
xor U25431 (N_25431,N_23032,N_19305);
and U25432 (N_25432,N_19683,N_18934);
nor U25433 (N_25433,N_22855,N_18377);
and U25434 (N_25434,N_22339,N_21902);
nand U25435 (N_25435,N_23815,N_21020);
or U25436 (N_25436,N_18576,N_22454);
and U25437 (N_25437,N_19679,N_21349);
xnor U25438 (N_25438,N_22170,N_23609);
xor U25439 (N_25439,N_19042,N_21664);
xor U25440 (N_25440,N_20781,N_19423);
or U25441 (N_25441,N_20089,N_23817);
or U25442 (N_25442,N_21259,N_23246);
nand U25443 (N_25443,N_23758,N_20199);
or U25444 (N_25444,N_19248,N_22365);
xor U25445 (N_25445,N_18657,N_19764);
and U25446 (N_25446,N_23179,N_19654);
nor U25447 (N_25447,N_20230,N_19066);
xnor U25448 (N_25448,N_21219,N_20051);
nand U25449 (N_25449,N_23488,N_21387);
or U25450 (N_25450,N_21307,N_18579);
or U25451 (N_25451,N_22542,N_22543);
xnor U25452 (N_25452,N_20353,N_19307);
xnor U25453 (N_25453,N_21412,N_21746);
xnor U25454 (N_25454,N_22285,N_22734);
nor U25455 (N_25455,N_19064,N_20552);
or U25456 (N_25456,N_19345,N_22176);
or U25457 (N_25457,N_19656,N_19610);
or U25458 (N_25458,N_20327,N_18334);
xnor U25459 (N_25459,N_23581,N_22423);
nand U25460 (N_25460,N_19413,N_22590);
nor U25461 (N_25461,N_19114,N_18427);
or U25462 (N_25462,N_20378,N_22246);
nand U25463 (N_25463,N_21429,N_22639);
xor U25464 (N_25464,N_20184,N_18779);
nand U25465 (N_25465,N_19094,N_19249);
nand U25466 (N_25466,N_19686,N_21556);
nor U25467 (N_25467,N_19860,N_21059);
and U25468 (N_25468,N_23390,N_21298);
nand U25469 (N_25469,N_18240,N_20898);
xor U25470 (N_25470,N_23374,N_22657);
nor U25471 (N_25471,N_20344,N_23297);
nand U25472 (N_25472,N_22727,N_21624);
or U25473 (N_25473,N_22748,N_18718);
xnor U25474 (N_25474,N_20895,N_19170);
or U25475 (N_25475,N_19273,N_20891);
and U25476 (N_25476,N_19041,N_20586);
or U25477 (N_25477,N_22791,N_19794);
nor U25478 (N_25478,N_19599,N_19223);
xnor U25479 (N_25479,N_21364,N_19299);
and U25480 (N_25480,N_22884,N_19526);
or U25481 (N_25481,N_21072,N_18085);
nand U25482 (N_25482,N_19918,N_18153);
or U25483 (N_25483,N_20173,N_19158);
nor U25484 (N_25484,N_22406,N_18329);
and U25485 (N_25485,N_20582,N_23768);
or U25486 (N_25486,N_18593,N_23312);
and U25487 (N_25487,N_18860,N_23646);
xor U25488 (N_25488,N_19837,N_20656);
or U25489 (N_25489,N_22885,N_22644);
nor U25490 (N_25490,N_18089,N_18295);
nor U25491 (N_25491,N_19151,N_20880);
nor U25492 (N_25492,N_18060,N_20826);
and U25493 (N_25493,N_23445,N_20924);
nand U25494 (N_25494,N_23753,N_20760);
or U25495 (N_25495,N_18571,N_19050);
xnor U25496 (N_25496,N_18278,N_22584);
nor U25497 (N_25497,N_18007,N_20294);
or U25498 (N_25498,N_23559,N_22681);
nor U25499 (N_25499,N_20967,N_20770);
nand U25500 (N_25500,N_22402,N_21917);
or U25501 (N_25501,N_19736,N_21197);
nor U25502 (N_25502,N_23238,N_22021);
nor U25503 (N_25503,N_21824,N_20647);
or U25504 (N_25504,N_18072,N_20461);
nor U25505 (N_25505,N_20601,N_21693);
and U25506 (N_25506,N_18559,N_21994);
or U25507 (N_25507,N_20833,N_19970);
nand U25508 (N_25508,N_20803,N_19913);
or U25509 (N_25509,N_21466,N_19137);
or U25510 (N_25510,N_18022,N_20805);
xor U25511 (N_25511,N_19178,N_20067);
and U25512 (N_25512,N_20446,N_19197);
and U25513 (N_25513,N_23270,N_21488);
nand U25514 (N_25514,N_22029,N_21014);
and U25515 (N_25515,N_21659,N_19678);
nor U25516 (N_25516,N_19059,N_18349);
and U25517 (N_25517,N_19324,N_18902);
nor U25518 (N_25518,N_23977,N_21732);
nor U25519 (N_25519,N_23544,N_19033);
nand U25520 (N_25520,N_23801,N_19631);
nand U25521 (N_25521,N_18735,N_21845);
xnor U25522 (N_25522,N_23471,N_22992);
xor U25523 (N_25523,N_19266,N_19604);
and U25524 (N_25524,N_18973,N_20376);
xor U25525 (N_25525,N_23012,N_23542);
nor U25526 (N_25526,N_21390,N_23997);
xor U25527 (N_25527,N_20429,N_21681);
or U25528 (N_25528,N_19742,N_23493);
nand U25529 (N_25529,N_20959,N_23588);
nand U25530 (N_25530,N_18927,N_18914);
nand U25531 (N_25531,N_18562,N_22350);
xnor U25532 (N_25532,N_18730,N_20017);
or U25533 (N_25533,N_20253,N_19962);
and U25534 (N_25534,N_19590,N_21525);
xor U25535 (N_25535,N_21027,N_23090);
xnor U25536 (N_25536,N_18650,N_19578);
and U25537 (N_25537,N_23851,N_21630);
and U25538 (N_25538,N_18317,N_19826);
nand U25539 (N_25539,N_21036,N_23001);
xnor U25540 (N_25540,N_20987,N_22969);
nor U25541 (N_25541,N_19036,N_19421);
nor U25542 (N_25542,N_20263,N_20023);
or U25543 (N_25543,N_23081,N_23879);
xor U25544 (N_25544,N_19523,N_21430);
nor U25545 (N_25545,N_23938,N_23127);
or U25546 (N_25546,N_20260,N_20964);
nand U25547 (N_25547,N_19640,N_19752);
nor U25548 (N_25548,N_19350,N_22258);
or U25549 (N_25549,N_18477,N_21767);
nor U25550 (N_25550,N_20076,N_23074);
or U25551 (N_25551,N_21703,N_23716);
xor U25552 (N_25552,N_21600,N_23283);
xnor U25553 (N_25553,N_20354,N_21798);
or U25554 (N_25554,N_23307,N_20899);
xnor U25555 (N_25555,N_18222,N_23496);
xor U25556 (N_25556,N_18813,N_20146);
or U25557 (N_25557,N_19303,N_23236);
or U25558 (N_25558,N_21328,N_21171);
nor U25559 (N_25559,N_21461,N_19213);
xnor U25560 (N_25560,N_21365,N_21784);
nor U25561 (N_25561,N_22888,N_19320);
xnor U25562 (N_25562,N_21053,N_21944);
or U25563 (N_25563,N_22686,N_21304);
nand U25564 (N_25564,N_20823,N_20608);
or U25565 (N_25565,N_21734,N_18456);
nor U25566 (N_25566,N_21056,N_22994);
nor U25567 (N_25567,N_23233,N_18959);
nor U25568 (N_25568,N_19173,N_22361);
xor U25569 (N_25569,N_18691,N_19548);
nor U25570 (N_25570,N_22764,N_19302);
and U25571 (N_25571,N_23129,N_21548);
or U25572 (N_25572,N_19988,N_23072);
and U25573 (N_25573,N_18926,N_18253);
nand U25574 (N_25574,N_21778,N_23141);
and U25575 (N_25575,N_20827,N_19808);
nor U25576 (N_25576,N_19670,N_22499);
nor U25577 (N_25577,N_21918,N_20416);
xnor U25578 (N_25578,N_21973,N_20700);
nand U25579 (N_25579,N_22521,N_20757);
or U25580 (N_25580,N_22068,N_19270);
or U25581 (N_25581,N_22961,N_19462);
xor U25582 (N_25582,N_22518,N_20154);
xnor U25583 (N_25583,N_23152,N_18207);
nand U25584 (N_25584,N_23394,N_19384);
or U25585 (N_25585,N_19055,N_19545);
and U25586 (N_25586,N_21517,N_20752);
nand U25587 (N_25587,N_22251,N_23895);
nand U25588 (N_25588,N_20070,N_22997);
nand U25589 (N_25589,N_23533,N_21274);
nand U25590 (N_25590,N_21642,N_23469);
and U25591 (N_25591,N_23968,N_21575);
and U25592 (N_25592,N_22964,N_22948);
nor U25593 (N_25593,N_22158,N_19506);
xor U25594 (N_25594,N_19087,N_18413);
and U25595 (N_25595,N_22837,N_22610);
nand U25596 (N_25596,N_21782,N_20118);
and U25597 (N_25597,N_18672,N_21055);
xnor U25598 (N_25598,N_18584,N_20892);
nand U25599 (N_25599,N_20079,N_21547);
xor U25600 (N_25600,N_21742,N_23806);
and U25601 (N_25601,N_22012,N_21777);
and U25602 (N_25602,N_19060,N_18589);
nand U25603 (N_25603,N_21478,N_22102);
nand U25604 (N_25604,N_19676,N_23859);
and U25605 (N_25605,N_18098,N_18596);
and U25606 (N_25606,N_19816,N_19023);
or U25607 (N_25607,N_21179,N_18385);
nor U25608 (N_25608,N_19755,N_18146);
xor U25609 (N_25609,N_18341,N_22883);
nor U25610 (N_25610,N_20657,N_21563);
or U25611 (N_25611,N_18852,N_22696);
nand U25612 (N_25612,N_18450,N_18025);
nor U25613 (N_25613,N_22411,N_20050);
xnor U25614 (N_25614,N_23096,N_22163);
nand U25615 (N_25615,N_19542,N_22991);
or U25616 (N_25616,N_23215,N_22404);
and U25617 (N_25617,N_18528,N_18549);
nor U25618 (N_25618,N_19032,N_22741);
xnor U25619 (N_25619,N_21859,N_19065);
nand U25620 (N_25620,N_19499,N_22996);
or U25621 (N_25621,N_23672,N_23836);
and U25622 (N_25622,N_21813,N_20315);
and U25623 (N_25623,N_19928,N_19955);
nor U25624 (N_25624,N_23978,N_22473);
nand U25625 (N_25625,N_21004,N_23098);
and U25626 (N_25626,N_22636,N_19553);
nor U25627 (N_25627,N_20953,N_22561);
xnor U25628 (N_25628,N_22532,N_21498);
xnor U25629 (N_25629,N_18128,N_19515);
nand U25630 (N_25630,N_23125,N_22300);
xnor U25631 (N_25631,N_21508,N_20259);
or U25632 (N_25632,N_22949,N_19122);
xor U25633 (N_25633,N_20142,N_21463);
and U25634 (N_25634,N_23683,N_23987);
or U25635 (N_25635,N_22272,N_20469);
xor U25636 (N_25636,N_23029,N_22774);
or U25637 (N_25637,N_21803,N_18882);
nand U25638 (N_25638,N_22391,N_23107);
xnor U25639 (N_25639,N_22970,N_19658);
and U25640 (N_25640,N_20214,N_21768);
nand U25641 (N_25641,N_21929,N_21645);
nand U25642 (N_25642,N_19193,N_22659);
xnor U25643 (N_25643,N_22808,N_19904);
xnor U25644 (N_25644,N_21204,N_20420);
xnor U25645 (N_25645,N_21409,N_19281);
and U25646 (N_25646,N_18111,N_20900);
nor U25647 (N_25647,N_19379,N_18964);
or U25648 (N_25648,N_22724,N_19877);
xnor U25649 (N_25649,N_23708,N_19536);
xor U25650 (N_25650,N_21309,N_18720);
xnor U25651 (N_25651,N_19228,N_23015);
and U25652 (N_25652,N_18195,N_18679);
nand U25653 (N_25653,N_18187,N_19793);
nor U25654 (N_25654,N_18068,N_19001);
nor U25655 (N_25655,N_23023,N_21065);
and U25656 (N_25656,N_19011,N_23560);
nor U25657 (N_25657,N_18226,N_22181);
nor U25658 (N_25658,N_20187,N_22227);
or U25659 (N_25659,N_20068,N_18292);
or U25660 (N_25660,N_19908,N_20617);
xnor U25661 (N_25661,N_18284,N_21960);
and U25662 (N_25662,N_19702,N_22002);
or U25663 (N_25663,N_23757,N_22100);
xnor U25664 (N_25664,N_23775,N_19401);
nand U25665 (N_25665,N_23557,N_20863);
xor U25666 (N_25666,N_19061,N_21423);
nor U25667 (N_25667,N_21597,N_19507);
nand U25668 (N_25668,N_20426,N_18018);
xor U25669 (N_25669,N_22419,N_23041);
xnor U25670 (N_25670,N_22206,N_22072);
nand U25671 (N_25671,N_18819,N_21281);
and U25672 (N_25672,N_23214,N_20989);
xnor U25673 (N_25673,N_21192,N_23973);
or U25674 (N_25674,N_23962,N_21311);
and U25675 (N_25675,N_22866,N_18262);
xnor U25676 (N_25676,N_22722,N_20160);
and U25677 (N_25677,N_19252,N_21514);
xnor U25678 (N_25678,N_19250,N_21366);
and U25679 (N_25679,N_22337,N_20511);
xor U25680 (N_25680,N_19997,N_22105);
or U25681 (N_25681,N_18421,N_23849);
xor U25682 (N_25682,N_20093,N_20807);
or U25683 (N_25683,N_21991,N_23732);
nor U25684 (N_25684,N_22818,N_18449);
nand U25685 (N_25685,N_21465,N_22063);
nand U25686 (N_25686,N_21110,N_18140);
nor U25687 (N_25687,N_21583,N_18405);
and U25688 (N_25688,N_20246,N_21984);
xnor U25689 (N_25689,N_19225,N_21679);
nor U25690 (N_25690,N_18339,N_20312);
nand U25691 (N_25691,N_20859,N_18289);
nand U25692 (N_25692,N_18470,N_23855);
nand U25693 (N_25693,N_23333,N_22847);
and U25694 (N_25694,N_18538,N_22235);
and U25695 (N_25695,N_23053,N_23727);
nand U25696 (N_25696,N_21111,N_22069);
xor U25697 (N_25697,N_18448,N_22190);
nand U25698 (N_25698,N_20736,N_20392);
nor U25699 (N_25699,N_18096,N_21314);
nor U25700 (N_25700,N_22408,N_18048);
or U25701 (N_25701,N_20874,N_23296);
and U25702 (N_25702,N_23232,N_18906);
or U25703 (N_25703,N_19297,N_20116);
xor U25704 (N_25704,N_21908,N_23064);
and U25705 (N_25705,N_23576,N_20234);
or U25706 (N_25706,N_19552,N_23271);
xnor U25707 (N_25707,N_22207,N_22033);
and U25708 (N_25708,N_23377,N_20813);
xnor U25709 (N_25709,N_18989,N_21437);
nor U25710 (N_25710,N_20069,N_19126);
nor U25711 (N_25711,N_23251,N_23161);
and U25712 (N_25712,N_18123,N_21188);
or U25713 (N_25713,N_23574,N_22401);
nand U25714 (N_25714,N_18244,N_21601);
and U25715 (N_25715,N_18446,N_20291);
and U25716 (N_25716,N_20205,N_20039);
xnor U25717 (N_25717,N_19445,N_20434);
and U25718 (N_25718,N_22749,N_21362);
nor U25719 (N_25719,N_23922,N_19132);
nor U25720 (N_25720,N_21982,N_21249);
xor U25721 (N_25721,N_18475,N_23587);
and U25722 (N_25722,N_23602,N_20029);
xor U25723 (N_25723,N_19198,N_22338);
nand U25724 (N_25724,N_20837,N_22905);
and U25725 (N_25725,N_18171,N_22840);
or U25726 (N_25726,N_23810,N_20666);
nor U25727 (N_25727,N_21683,N_20399);
nor U25728 (N_25728,N_23854,N_20787);
nor U25729 (N_25729,N_22184,N_18778);
xnor U25730 (N_25730,N_22436,N_20800);
and U25731 (N_25731,N_22891,N_20318);
xor U25732 (N_25732,N_20269,N_23877);
nand U25733 (N_25733,N_20541,N_18648);
xnor U25734 (N_25734,N_19502,N_18874);
and U25735 (N_25735,N_20090,N_22302);
or U25736 (N_25736,N_22082,N_19070);
nand U25737 (N_25737,N_19388,N_20296);
nor U25738 (N_25738,N_20136,N_23166);
nor U25739 (N_25739,N_23818,N_19721);
and U25740 (N_25740,N_20110,N_18452);
nor U25741 (N_25741,N_18322,N_23920);
or U25742 (N_25742,N_18856,N_18971);
and U25743 (N_25743,N_22373,N_23951);
and U25744 (N_25744,N_20281,N_20013);
nor U25745 (N_25745,N_19336,N_21817);
or U25746 (N_25746,N_23516,N_23044);
and U25747 (N_25747,N_21868,N_22237);
xor U25748 (N_25748,N_19075,N_21486);
xnor U25749 (N_25749,N_22714,N_21533);
nand U25750 (N_25750,N_18504,N_23798);
or U25751 (N_25751,N_19054,N_23459);
xor U25752 (N_25752,N_19461,N_20786);
or U25753 (N_25753,N_21698,N_19037);
or U25754 (N_25754,N_22453,N_20311);
and U25755 (N_25755,N_18600,N_18087);
and U25756 (N_25756,N_18734,N_19192);
nand U25757 (N_25757,N_22260,N_20303);
and U25758 (N_25758,N_19424,N_23656);
nor U25759 (N_25759,N_19386,N_18823);
and U25760 (N_25760,N_22347,N_18234);
xor U25761 (N_25761,N_19435,N_21151);
nor U25762 (N_25762,N_18024,N_23949);
nand U25763 (N_25763,N_21225,N_19627);
nand U25764 (N_25764,N_20008,N_23148);
or U25765 (N_25765,N_20244,N_23800);
nand U25766 (N_25766,N_21345,N_23631);
xor U25767 (N_25767,N_18167,N_20513);
or U25768 (N_25768,N_22987,N_18011);
or U25769 (N_25769,N_19585,N_18150);
and U25770 (N_25770,N_23913,N_18159);
xnor U25771 (N_25771,N_20170,N_20155);
and U25772 (N_25772,N_23426,N_21457);
and U25773 (N_25773,N_23983,N_23402);
nor U25774 (N_25774,N_20985,N_23864);
nand U25775 (N_25775,N_21206,N_20455);
and U25776 (N_25776,N_23764,N_22618);
nor U25777 (N_25777,N_20194,N_23382);
nor U25778 (N_25778,N_18090,N_21003);
nand U25779 (N_25779,N_18525,N_21312);
nor U25780 (N_25780,N_20213,N_22525);
xnor U25781 (N_25781,N_23856,N_23547);
and U25782 (N_25782,N_18924,N_22133);
and U25783 (N_25783,N_18184,N_20991);
and U25784 (N_25784,N_19470,N_20670);
nand U25785 (N_25785,N_21875,N_23163);
or U25786 (N_25786,N_22928,N_23114);
or U25787 (N_25787,N_23643,N_19204);
xnor U25788 (N_25788,N_20152,N_22792);
or U25789 (N_25789,N_21992,N_20492);
or U25790 (N_25790,N_23838,N_23002);
xor U25791 (N_25791,N_18432,N_23216);
or U25792 (N_25792,N_21972,N_18176);
or U25793 (N_25793,N_23663,N_20508);
nand U25794 (N_25794,N_19038,N_20790);
xnor U25795 (N_25795,N_19107,N_18627);
or U25796 (N_25796,N_21928,N_22544);
or U25797 (N_25797,N_18071,N_22134);
xnor U25798 (N_25798,N_23117,N_20276);
xnor U25799 (N_25799,N_23077,N_19078);
and U25800 (N_25800,N_21728,N_20236);
and U25801 (N_25801,N_20266,N_20085);
xor U25802 (N_25802,N_20278,N_21482);
and U25803 (N_25803,N_19935,N_21363);
and U25804 (N_25804,N_23679,N_21256);
or U25805 (N_25805,N_22107,N_23268);
or U25806 (N_25806,N_21061,N_23156);
nand U25807 (N_25807,N_22923,N_18206);
nand U25808 (N_25808,N_23033,N_18618);
xor U25809 (N_25809,N_18274,N_18197);
nor U25810 (N_25810,N_21223,N_22782);
or U25811 (N_25811,N_20335,N_23696);
and U25812 (N_25812,N_18727,N_18595);
xor U25813 (N_25813,N_19458,N_18122);
or U25814 (N_25814,N_22924,N_21282);
and U25815 (N_25815,N_22335,N_21166);
xor U25816 (N_25816,N_20147,N_21191);
or U25817 (N_25817,N_18807,N_21791);
nand U25818 (N_25818,N_22126,N_22752);
nand U25819 (N_25819,N_21559,N_23027);
and U25820 (N_25820,N_22092,N_23217);
and U25821 (N_25821,N_20929,N_18118);
nand U25822 (N_25822,N_23403,N_22786);
and U25823 (N_25823,N_18501,N_21825);
and U25824 (N_25824,N_21931,N_22576);
nand U25825 (N_25825,N_18218,N_19516);
and U25826 (N_25826,N_22508,N_18400);
nand U25827 (N_25827,N_18843,N_19076);
nand U25828 (N_25828,N_22904,N_22988);
nand U25829 (N_25829,N_20965,N_23737);
xnor U25830 (N_25830,N_19915,N_19100);
nand U25831 (N_25831,N_22807,N_18899);
nand U25832 (N_25832,N_22841,N_21788);
or U25833 (N_25833,N_22336,N_20566);
xor U25834 (N_25834,N_21277,N_18462);
nor U25835 (N_25835,N_20794,N_20848);
xnor U25836 (N_25836,N_20846,N_22194);
nand U25837 (N_25837,N_18706,N_18316);
or U25838 (N_25838,N_21157,N_20381);
nand U25839 (N_25839,N_19287,N_19505);
nand U25840 (N_25840,N_18929,N_21936);
xnor U25841 (N_25841,N_23707,N_18531);
nand U25842 (N_25842,N_21043,N_19960);
nand U25843 (N_25843,N_19660,N_22652);
and U25844 (N_25844,N_19573,N_21923);
xnor U25845 (N_25845,N_19522,N_21935);
and U25846 (N_25846,N_18430,N_20996);
nor U25847 (N_25847,N_22312,N_19330);
nand U25848 (N_25848,N_19951,N_23894);
xor U25849 (N_25849,N_23381,N_20758);
nor U25850 (N_25850,N_22498,N_18878);
xnor U25851 (N_25851,N_19589,N_21444);
xor U25852 (N_25852,N_19308,N_22308);
or U25853 (N_25853,N_23610,N_19309);
xnor U25854 (N_25854,N_21324,N_23085);
nand U25855 (N_25855,N_19834,N_21414);
nor U25856 (N_25856,N_21295,N_22088);
and U25857 (N_25857,N_22723,N_21479);
nand U25858 (N_25858,N_18769,N_20494);
and U25859 (N_25859,N_18637,N_22334);
nand U25860 (N_25860,N_18005,N_21112);
nor U25861 (N_25861,N_21008,N_18652);
xnor U25862 (N_25862,N_22185,N_20975);
nor U25863 (N_25863,N_20560,N_19982);
nor U25864 (N_25864,N_23892,N_22281);
nand U25865 (N_25865,N_18621,N_23150);
xnor U25866 (N_25866,N_18708,N_22136);
or U25867 (N_25867,N_22726,N_21974);
or U25868 (N_25868,N_20937,N_23185);
xnor U25869 (N_25869,N_21007,N_22317);
xnor U25870 (N_25870,N_20130,N_22845);
xnor U25871 (N_25871,N_18163,N_20279);
and U25872 (N_25872,N_20574,N_18764);
or U25873 (N_25873,N_20126,N_21167);
nor U25874 (N_25874,N_23460,N_18481);
xnor U25875 (N_25875,N_22632,N_22383);
nor U25876 (N_25876,N_19053,N_19525);
nand U25877 (N_25877,N_19774,N_19175);
xor U25878 (N_25878,N_19189,N_23195);
nand U25879 (N_25879,N_18905,N_19447);
nor U25880 (N_25880,N_18608,N_18061);
nand U25881 (N_25881,N_19219,N_23878);
and U25882 (N_25882,N_19098,N_19932);
or U25883 (N_25883,N_19584,N_18644);
xnor U25884 (N_25884,N_20433,N_23075);
and U25885 (N_25885,N_21114,N_23554);
nor U25886 (N_25886,N_20407,N_22912);
and U25887 (N_25887,N_21117,N_21899);
or U25888 (N_25888,N_22466,N_21750);
xnor U25889 (N_25889,N_21881,N_23290);
nor U25890 (N_25890,N_21539,N_19717);
or U25891 (N_25891,N_20916,N_20980);
xnor U25892 (N_25892,N_20107,N_22264);
xnor U25893 (N_25893,N_21530,N_20196);
or U25894 (N_25894,N_20630,N_22039);
nor U25895 (N_25895,N_22567,N_18335);
or U25896 (N_25896,N_20364,N_18044);
and U25897 (N_25897,N_20440,N_19977);
or U25898 (N_25898,N_18077,N_18767);
nor U25899 (N_25899,N_19638,N_23803);
nand U25900 (N_25900,N_21235,N_20620);
xor U25901 (N_25901,N_22695,N_23937);
or U25902 (N_25902,N_23173,N_21769);
and U25903 (N_25903,N_18836,N_18928);
or U25904 (N_25904,N_20817,N_18460);
nand U25905 (N_25905,N_19092,N_21880);
nor U25906 (N_25906,N_20408,N_19444);
nand U25907 (N_25907,N_22019,N_20868);
and U25908 (N_25908,N_22663,N_23969);
nand U25909 (N_25909,N_18749,N_23975);
and U25910 (N_25910,N_18849,N_22055);
nor U25911 (N_25911,N_21325,N_22231);
xnor U25912 (N_25912,N_19187,N_20343);
and U25913 (N_25913,N_23391,N_21477);
or U25914 (N_25914,N_23582,N_21696);
and U25915 (N_25915,N_23039,N_21493);
nand U25916 (N_25916,N_23210,N_22121);
nand U25917 (N_25917,N_20215,N_20283);
and U25918 (N_25918,N_23109,N_19791);
nor U25919 (N_25919,N_18736,N_23358);
or U25920 (N_25920,N_19572,N_20726);
or U25921 (N_25921,N_21302,N_21915);
xnor U25922 (N_25922,N_22149,N_22424);
and U25923 (N_25923,N_18754,N_23131);
xnor U25924 (N_25924,N_18346,N_19326);
or U25925 (N_25925,N_23594,N_18301);
nand U25926 (N_25926,N_22766,N_20661);
or U25927 (N_25927,N_23944,N_18084);
xor U25928 (N_25928,N_23946,N_23222);
or U25929 (N_25929,N_22214,N_23820);
xor U25930 (N_25930,N_23455,N_19849);
and U25931 (N_25931,N_18647,N_23916);
and U25932 (N_25932,N_22902,N_21275);
and U25933 (N_25933,N_19282,N_19909);
nor U25934 (N_25934,N_21050,N_20148);
nor U25935 (N_25935,N_19331,N_20045);
xor U25936 (N_25936,N_23828,N_19753);
nor U25937 (N_25937,N_18023,N_19989);
nand U25938 (N_25938,N_20159,N_18493);
and U25939 (N_25939,N_22520,N_23293);
nor U25940 (N_25940,N_20001,N_20306);
and U25941 (N_25941,N_20351,N_21377);
nor U25942 (N_25942,N_22881,N_22679);
or U25943 (N_25943,N_23833,N_23673);
xnor U25944 (N_25944,N_21680,N_19121);
nor U25945 (N_25945,N_20124,N_23353);
and U25946 (N_25946,N_23261,N_22938);
or U25947 (N_25947,N_19872,N_20383);
nand U25948 (N_25948,N_18646,N_18239);
xor U25949 (N_25949,N_22311,N_21286);
nand U25950 (N_25950,N_19338,N_20723);
xnor U25951 (N_25951,N_22947,N_20926);
nand U25952 (N_25952,N_21272,N_18574);
and U25953 (N_25953,N_19412,N_23031);
xnor U25954 (N_25954,N_19426,N_23641);
nand U25955 (N_25955,N_22955,N_21546);
xnor U25956 (N_25956,N_20324,N_22735);
nor U25957 (N_25957,N_20476,N_22504);
or U25958 (N_25958,N_20867,N_21838);
nand U25959 (N_25959,N_23807,N_19351);
or U25960 (N_25960,N_20452,N_22907);
or U25961 (N_25961,N_23957,N_18386);
and U25962 (N_25962,N_23428,N_21124);
xor U25963 (N_25963,N_23087,N_20948);
and U25964 (N_25964,N_23778,N_23680);
or U25965 (N_25965,N_22202,N_20264);
xnor U25966 (N_25966,N_19410,N_21401);
xnor U25967 (N_25967,N_19891,N_22580);
nor U25968 (N_25968,N_22634,N_22234);
nand U25969 (N_25969,N_22086,N_22315);
nand U25970 (N_25970,N_21743,N_18671);
nand U25971 (N_25971,N_23909,N_18108);
and U25972 (N_25972,N_22223,N_20198);
xor U25973 (N_25973,N_19583,N_20484);
nor U25974 (N_25974,N_19867,N_19841);
xnor U25975 (N_25975,N_20849,N_21156);
and U25976 (N_25976,N_23269,N_19917);
xnor U25977 (N_25977,N_23688,N_22535);
nor U25978 (N_25978,N_20098,N_20495);
nand U25979 (N_25979,N_19200,N_19149);
xor U25980 (N_25980,N_18132,N_23180);
or U25981 (N_25981,N_18533,N_20012);
xnor U25982 (N_25982,N_20391,N_18725);
nand U25983 (N_25983,N_20628,N_21400);
nand U25984 (N_25984,N_21372,N_21590);
nand U25985 (N_25985,N_22148,N_23991);
nor U25986 (N_25986,N_22444,N_21735);
nor U25987 (N_25987,N_19110,N_21242);
nand U25988 (N_25988,N_21451,N_22798);
and U25989 (N_25989,N_20971,N_20060);
and U25990 (N_25990,N_18305,N_23122);
or U25991 (N_25991,N_21353,N_21647);
or U25992 (N_25992,N_21230,N_18983);
nor U25993 (N_25993,N_20299,N_23740);
xnor U25994 (N_25994,N_23827,N_20804);
nand U25995 (N_25995,N_20151,N_20191);
xor U25996 (N_25996,N_19725,N_19550);
and U25997 (N_25997,N_23069,N_23016);
nand U25998 (N_25998,N_21276,N_18507);
nand U25999 (N_25999,N_20785,N_22382);
and U26000 (N_26000,N_22486,N_23154);
or U26001 (N_26001,N_21628,N_20646);
xor U26002 (N_26002,N_21067,N_20465);
xnor U26003 (N_26003,N_19870,N_22849);
nor U26004 (N_26004,N_22358,N_22890);
xor U26005 (N_26005,N_18607,N_23457);
nand U26006 (N_26006,N_22396,N_20517);
xor U26007 (N_26007,N_20387,N_18613);
or U26008 (N_26008,N_19416,N_19801);
nand U26009 (N_26009,N_21173,N_19460);
or U26010 (N_26010,N_21966,N_21685);
or U26011 (N_26011,N_20273,N_18156);
nand U26012 (N_26012,N_23308,N_22397);
nor U26013 (N_26013,N_18887,N_23762);
nand U26014 (N_26014,N_21238,N_21890);
or U26015 (N_26015,N_20911,N_20567);
xnor U26016 (N_26016,N_19150,N_23132);
nand U26017 (N_26017,N_21997,N_23286);
nand U26018 (N_26018,N_23669,N_22495);
nor U26019 (N_26019,N_19882,N_22848);
nor U26020 (N_26020,N_21836,N_21296);
and U26021 (N_26021,N_23279,N_18429);
and U26022 (N_26022,N_23371,N_18178);
nor U26023 (N_26023,N_18035,N_23478);
and U26024 (N_26024,N_21125,N_18383);
or U26025 (N_26025,N_23310,N_19714);
or U26026 (N_26026,N_18567,N_22865);
nor U26027 (N_26027,N_18758,N_23187);
nor U26028 (N_26028,N_23945,N_20027);
and U26029 (N_26029,N_18858,N_22736);
or U26030 (N_26030,N_22440,N_23655);
xor U26031 (N_26031,N_21077,N_18215);
xor U26032 (N_26032,N_22500,N_23370);
xor U26033 (N_26033,N_21745,N_23071);
nand U26034 (N_26034,N_21998,N_20587);
nand U26035 (N_26035,N_21346,N_20747);
nand U26036 (N_26036,N_20974,N_18120);
xnor U26037 (N_26037,N_21379,N_23770);
or U26038 (N_26038,N_18573,N_22098);
nor U26039 (N_26039,N_18097,N_21270);
or U26040 (N_26040,N_19484,N_23451);
nor U26041 (N_26041,N_23925,N_20636);
nand U26042 (N_26042,N_19803,N_19560);
or U26043 (N_26043,N_20414,N_18747);
and U26044 (N_26044,N_18831,N_23396);
nor U26045 (N_26045,N_22114,N_22708);
and U26046 (N_26046,N_18524,N_21968);
xor U26047 (N_26047,N_20201,N_18426);
and U26048 (N_26048,N_20871,N_23252);
xor U26049 (N_26049,N_20463,N_18695);
nand U26050 (N_26050,N_22981,N_22557);
xnor U26051 (N_26051,N_19085,N_18326);
and U26052 (N_26052,N_19024,N_20801);
xnor U26053 (N_26053,N_19377,N_22425);
xor U26054 (N_26054,N_23084,N_18312);
nand U26055 (N_26055,N_18257,N_18742);
xor U26056 (N_26056,N_19002,N_23119);
xor U26057 (N_26057,N_20436,N_18506);
and U26058 (N_26058,N_18561,N_19467);
and U26059 (N_26059,N_19622,N_21287);
nand U26060 (N_26060,N_18418,N_22760);
nand U26061 (N_26061,N_18521,N_20208);
or U26062 (N_26062,N_21507,N_20403);
nand U26063 (N_26063,N_23857,N_20939);
and U26064 (N_26064,N_18348,N_23897);
xnor U26065 (N_26065,N_22241,N_20103);
nand U26066 (N_26066,N_21702,N_22778);
nand U26067 (N_26067,N_21248,N_20776);
or U26068 (N_26068,N_23888,N_18859);
xor U26069 (N_26069,N_23300,N_18616);
xnor U26070 (N_26070,N_20095,N_20157);
nand U26071 (N_26071,N_23495,N_23338);
nand U26072 (N_26072,N_23625,N_18634);
and U26073 (N_26073,N_22962,N_21081);
or U26074 (N_26074,N_23992,N_21147);
and U26075 (N_26075,N_23482,N_18293);
nand U26076 (N_26076,N_19966,N_21961);
and U26077 (N_26077,N_23571,N_21202);
or U26078 (N_26078,N_22089,N_22120);
xor U26079 (N_26079,N_18977,N_18070);
and U26080 (N_26080,N_23375,N_20331);
xor U26081 (N_26081,N_21592,N_18586);
nor U26082 (N_26082,N_20225,N_20267);
xor U26083 (N_26083,N_20731,N_18468);
nand U26084 (N_26084,N_20310,N_22920);
nor U26085 (N_26085,N_18004,N_20976);
nor U26086 (N_26086,N_22004,N_21840);
or U26087 (N_26087,N_19088,N_20271);
or U26088 (N_26088,N_19765,N_23247);
and U26089 (N_26089,N_21527,N_23918);
nand U26090 (N_26090,N_19301,N_21190);
nand U26091 (N_26091,N_18799,N_23480);
nand U26092 (N_26092,N_23483,N_18527);
nand U26093 (N_26093,N_23580,N_18654);
nor U26094 (N_26094,N_23745,N_20835);
xnor U26095 (N_26095,N_18469,N_18518);
and U26096 (N_26096,N_20121,N_22706);
xnor U26097 (N_26097,N_22745,N_19821);
nand U26098 (N_26098,N_23104,N_22656);
nor U26099 (N_26099,N_22129,N_20500);
nor U26100 (N_26100,N_20793,N_20366);
and U26101 (N_26101,N_21116,N_22279);
or U26102 (N_26102,N_23049,N_21422);
and U26103 (N_26103,N_21637,N_21639);
xnor U26104 (N_26104,N_22478,N_21989);
xor U26105 (N_26105,N_21950,N_19481);
nand U26106 (N_26106,N_22387,N_23171);
xor U26107 (N_26107,N_21358,N_18726);
or U26108 (N_26108,N_21963,N_23088);
xor U26109 (N_26109,N_21265,N_18463);
xor U26110 (N_26110,N_18041,N_22694);
nand U26111 (N_26111,N_22922,N_21029);
or U26112 (N_26112,N_19195,N_22421);
or U26113 (N_26113,N_20561,N_20896);
or U26114 (N_26114,N_20563,N_18423);
xnor U26115 (N_26115,N_20247,N_18056);
xor U26116 (N_26116,N_21726,N_19597);
and U26117 (N_26117,N_19146,N_19003);
or U26118 (N_26118,N_18302,N_21588);
xor U26119 (N_26119,N_21854,N_20627);
or U26120 (N_26120,N_19361,N_23915);
or U26121 (N_26121,N_20128,N_19074);
xnor U26122 (N_26122,N_18748,N_18057);
nor U26123 (N_26123,N_20423,N_19569);
nor U26124 (N_26124,N_22113,N_22868);
and U26125 (N_26125,N_21234,N_21818);
and U26126 (N_26126,N_19829,N_18886);
nand U26127 (N_26127,N_21208,N_18054);
or U26128 (N_26128,N_22545,N_19035);
and U26129 (N_26129,N_21832,N_22131);
or U26130 (N_26130,N_22080,N_23024);
xor U26131 (N_26131,N_21729,N_21434);
and U26132 (N_26132,N_18667,N_18350);
or U26133 (N_26133,N_20105,N_22101);
nor U26134 (N_26134,N_19105,N_19740);
or U26135 (N_26135,N_22631,N_21901);
nor U26136 (N_26136,N_19869,N_18345);
and U26137 (N_26137,N_19886,N_18921);
xor U26138 (N_26138,N_19768,N_22560);
nand U26139 (N_26139,N_22523,N_23970);
and U26140 (N_26140,N_21752,N_20732);
nor U26141 (N_26141,N_23149,N_21339);
or U26142 (N_26142,N_18865,N_22035);
nand U26143 (N_26143,N_18113,N_22414);
nor U26144 (N_26144,N_21521,N_22633);
nor U26145 (N_26145,N_20505,N_18537);
xnor U26146 (N_26146,N_18321,N_18751);
nor U26147 (N_26147,N_21367,N_18731);
and U26148 (N_26148,N_23021,N_19294);
or U26149 (N_26149,N_19687,N_20977);
nor U26150 (N_26150,N_20486,N_19873);
xnor U26151 (N_26151,N_18709,N_20137);
and U26152 (N_26152,N_19365,N_18665);
or U26153 (N_26153,N_20535,N_21485);
and U26154 (N_26154,N_20998,N_19595);
or U26155 (N_26155,N_21181,N_18817);
nand U26156 (N_26156,N_22390,N_18359);
nand U26157 (N_26157,N_18440,N_21212);
and U26158 (N_26158,N_19668,N_22331);
and U26159 (N_26159,N_22244,N_23712);
nand U26160 (N_26160,N_20678,N_22330);
and U26161 (N_26161,N_22789,N_18811);
nor U26162 (N_26162,N_20802,N_23151);
and U26163 (N_26163,N_21652,N_22389);
or U26164 (N_26164,N_18175,N_19903);
nor U26165 (N_26165,N_18076,N_20619);
nand U26166 (N_26166,N_22582,N_19685);
nor U26167 (N_26167,N_22351,N_20579);
or U26168 (N_26168,N_21862,N_22122);
nor U26169 (N_26169,N_20653,N_21614);
or U26170 (N_26170,N_23742,N_18053);
nand U26171 (N_26171,N_18310,N_19684);
nand U26172 (N_26172,N_18804,N_20555);
nand U26173 (N_26173,N_18073,N_18152);
nand U26174 (N_26174,N_21096,N_21737);
and U26175 (N_26175,N_23224,N_20405);
nor U26176 (N_26176,N_18186,N_20865);
nand U26177 (N_26177,N_23703,N_19123);
nor U26178 (N_26178,N_21051,N_23744);
or U26179 (N_26179,N_21995,N_23837);
nor U26180 (N_26180,N_19206,N_23034);
xnor U26181 (N_26181,N_22159,N_19404);
nor U26182 (N_26182,N_20876,N_22513);
and U26183 (N_26183,N_20385,N_22342);
nor U26184 (N_26184,N_18444,N_20857);
and U26185 (N_26185,N_20127,N_23747);
xor U26186 (N_26186,N_22834,N_18988);
nand U26187 (N_26187,N_22463,N_21779);
xor U26188 (N_26188,N_18877,N_18602);
nor U26189 (N_26189,N_22978,N_23395);
or U26190 (N_26190,N_20695,N_22056);
xnor U26191 (N_26191,N_22522,N_20396);
nand U26192 (N_26192,N_23891,N_21741);
xor U26193 (N_26193,N_22701,N_22022);
xnor U26194 (N_26194,N_23102,N_20162);
nand U26195 (N_26195,N_18536,N_20430);
xor U26196 (N_26196,N_20314,N_21506);
xnor U26197 (N_26197,N_20943,N_22534);
nor U26198 (N_26198,N_18866,N_18577);
nor U26199 (N_26199,N_21738,N_21938);
and U26200 (N_26200,N_18916,N_23393);
xnor U26201 (N_26201,N_18333,N_19131);
nand U26202 (N_26202,N_20375,N_23869);
nor U26203 (N_26203,N_22768,N_22566);
xor U26204 (N_26204,N_19010,N_23782);
and U26205 (N_26205,N_22257,N_19163);
and U26206 (N_26206,N_20262,N_19626);
xnor U26207 (N_26207,N_20526,N_23175);
nor U26208 (N_26208,N_21129,N_20970);
or U26209 (N_26209,N_23095,N_23138);
and U26210 (N_26210,N_19643,N_20862);
xnor U26211 (N_26211,N_18402,N_23990);
nor U26212 (N_26212,N_21229,N_21005);
nor U26213 (N_26213,N_19263,N_23617);
nor U26214 (N_26214,N_18086,N_18106);
xnor U26215 (N_26215,N_23264,N_22053);
nand U26216 (N_26216,N_23443,N_23486);
and U26217 (N_26217,N_19392,N_21543);
or U26218 (N_26218,N_22310,N_19864);
xor U26219 (N_26219,N_22519,N_22014);
and U26220 (N_26220,N_22085,N_23598);
and U26221 (N_26221,N_23040,N_23726);
xnor U26222 (N_26222,N_23994,N_22780);
xor U26223 (N_26223,N_20242,N_21924);
and U26224 (N_26224,N_19400,N_21342);
xnor U26225 (N_26225,N_19127,N_22321);
or U26226 (N_26226,N_21571,N_18873);
or U26227 (N_26227,N_18800,N_20028);
or U26228 (N_26228,N_18570,N_20280);
or U26229 (N_26229,N_23228,N_23507);
or U26230 (N_26230,N_20745,N_23368);
nor U26231 (N_26231,N_18225,N_21405);
nand U26232 (N_26232,N_21564,N_18741);
or U26233 (N_26233,N_23207,N_20642);
nor U26234 (N_26234,N_22658,N_18117);
nand U26235 (N_26235,N_20442,N_19866);
and U26236 (N_26236,N_23657,N_19090);
nor U26237 (N_26237,N_18510,N_18879);
or U26238 (N_26238,N_20119,N_23250);
nor U26239 (N_26239,N_19368,N_19762);
xnor U26240 (N_26240,N_22999,N_21793);
and U26241 (N_26241,N_19926,N_19487);
nor U26242 (N_26242,N_21611,N_23289);
nor U26243 (N_26243,N_21128,N_18690);
nand U26244 (N_26244,N_23850,N_22154);
nand U26245 (N_26245,N_18199,N_20612);
xor U26246 (N_26246,N_18074,N_21708);
xnor U26247 (N_26247,N_21786,N_22253);
or U26248 (N_26248,N_20659,N_22531);
nor U26249 (N_26249,N_21266,N_22919);
nand U26250 (N_26250,N_19108,N_22875);
and U26251 (N_26251,N_22986,N_20397);
and U26252 (N_26252,N_21260,N_20004);
xor U26253 (N_26253,N_23904,N_20698);
nand U26254 (N_26254,N_18021,N_18093);
nor U26255 (N_26255,N_19509,N_18443);
xnor U26256 (N_26256,N_22801,N_22753);
xnor U26257 (N_26257,N_21326,N_18232);
and U26258 (N_26258,N_20966,N_18626);
and U26259 (N_26259,N_19159,N_18540);
or U26260 (N_26260,N_18366,N_21145);
and U26261 (N_26261,N_21733,N_22455);
or U26262 (N_26262,N_20464,N_18375);
and U26263 (N_26263,N_22762,N_23564);
nor U26264 (N_26264,N_23637,N_20357);
and U26265 (N_26265,N_21537,N_18080);
nor U26266 (N_26266,N_21897,N_20717);
nor U26267 (N_26267,N_21237,N_21657);
or U26268 (N_26268,N_20847,N_18485);
and U26269 (N_26269,N_21809,N_19310);
and U26270 (N_26270,N_19258,N_19544);
nand U26271 (N_26271,N_19963,N_23340);
or U26272 (N_26272,N_23541,N_18364);
xnor U26273 (N_26273,N_21389,N_22434);
and U26274 (N_26274,N_23611,N_18263);
nor U26275 (N_26275,N_19859,N_21580);
xor U26276 (N_26276,N_19128,N_21958);
nor U26277 (N_26277,N_21762,N_19775);
and U26278 (N_26278,N_23843,N_23881);
xor U26279 (N_26279,N_20514,N_22293);
nor U26280 (N_26280,N_20908,N_20904);
or U26281 (N_26281,N_19147,N_21747);
or U26282 (N_26282,N_19234,N_19734);
nor U26283 (N_26283,N_22189,N_22369);
nor U26284 (N_26284,N_23221,N_19186);
xor U26285 (N_26285,N_23774,N_18513);
xnor U26286 (N_26286,N_21284,N_21251);
and U26287 (N_26287,N_23137,N_22670);
nor U26288 (N_26288,N_21895,N_18666);
or U26289 (N_26289,N_20228,N_23797);
or U26290 (N_26290,N_21830,N_20854);
and U26291 (N_26291,N_23009,N_19188);
nand U26292 (N_26292,N_19827,N_21585);
nand U26293 (N_26293,N_20819,N_20041);
xnor U26294 (N_26294,N_21491,N_20662);
nor U26295 (N_26295,N_18100,N_20077);
nand U26296 (N_26296,N_22044,N_18824);
nand U26297 (N_26297,N_23522,N_22913);
nor U26298 (N_26298,N_18942,N_18833);
and U26299 (N_26299,N_19172,N_21464);
xor U26300 (N_26300,N_23785,N_23695);
and U26301 (N_26301,N_22374,N_20931);
nor U26302 (N_26302,N_21510,N_23772);
xnor U26303 (N_26303,N_20186,N_23867);
or U26304 (N_26304,N_21655,N_21186);
nand U26305 (N_26305,N_18419,N_19593);
nor U26306 (N_26306,N_20190,N_21135);
nand U26307 (N_26307,N_18689,N_18892);
nor U26308 (N_26308,N_22783,N_23376);
and U26309 (N_26309,N_20683,N_22861);
nor U26310 (N_26310,N_22896,N_23619);
and U26311 (N_26311,N_20386,N_20167);
nand U26312 (N_26312,N_19930,N_21074);
nor U26313 (N_26313,N_19194,N_19062);
nand U26314 (N_26314,N_22062,N_22718);
nand U26315 (N_26315,N_20639,N_22040);
xor U26316 (N_26316,N_22394,N_20597);
nand U26317 (N_26317,N_21073,N_18729);
or U26318 (N_26318,N_18903,N_22422);
nor U26319 (N_26319,N_18309,N_18837);
nor U26320 (N_26320,N_22471,N_21866);
nor U26321 (N_26321,N_23648,N_19884);
or U26322 (N_26322,N_23713,N_23422);
and U26323 (N_26323,N_18033,N_19289);
or U26324 (N_26324,N_20104,N_18982);
nand U26325 (N_26325,N_22291,N_22201);
xnor U26326 (N_26326,N_19592,N_20927);
and U26327 (N_26327,N_21532,N_18165);
nor U26328 (N_26328,N_23687,N_21396);
xor U26329 (N_26329,N_21258,N_19892);
xnor U26330 (N_26330,N_18952,N_18180);
or U26331 (N_26331,N_21542,N_23126);
or U26332 (N_26332,N_21578,N_23676);
and U26333 (N_26333,N_19205,N_22673);
nor U26334 (N_26334,N_20658,N_21012);
or U26335 (N_26335,N_21844,N_20338);
and U26336 (N_26336,N_19722,N_23503);
and U26337 (N_26337,N_19657,N_23607);
xor U26338 (N_26338,N_22717,N_20250);
xor U26339 (N_26339,N_18283,N_22826);
nor U26340 (N_26340,N_20491,N_23128);
nor U26341 (N_26341,N_18365,N_18436);
nor U26342 (N_26342,N_19984,N_23218);
nor U26343 (N_26343,N_19456,N_23147);
nor U26344 (N_26344,N_19148,N_21608);
or U26345 (N_26345,N_21976,N_20551);
xor U26346 (N_26346,N_23101,N_23192);
xnor U26347 (N_26347,N_22007,N_19097);
xor U26348 (N_26348,N_18380,N_19588);
and U26349 (N_26349,N_18136,N_23842);
or U26350 (N_26350,N_20109,N_22689);
nand U26351 (N_26351,N_21330,N_21505);
nand U26352 (N_26352,N_23492,N_21932);
xor U26353 (N_26353,N_22205,N_18545);
and U26354 (N_26354,N_18765,N_21526);
xnor U26355 (N_26355,N_20605,N_22607);
xnor U26356 (N_26356,N_19780,N_19373);
xnor U26357 (N_26357,N_21595,N_23344);
and U26358 (N_26358,N_22575,N_19777);
or U26359 (N_26359,N_18119,N_22461);
and U26360 (N_26360,N_20099,N_20767);
or U26361 (N_26361,N_18946,N_19540);
nand U26362 (N_26362,N_20493,N_23513);
nand U26363 (N_26363,N_20881,N_20428);
and U26364 (N_26364,N_20091,N_23796);
nand U26365 (N_26365,N_23456,N_21561);
and U26366 (N_26366,N_21519,N_19665);
xnor U26367 (N_26367,N_23265,N_19451);
xnor U26368 (N_26368,N_21017,N_18861);
xnor U26369 (N_26369,N_21292,N_18864);
and U26370 (N_26370,N_23070,N_19117);
or U26371 (N_26371,N_19941,N_19165);
and U26372 (N_26372,N_23162,N_20135);
xor U26373 (N_26373,N_18933,N_18737);
and U26374 (N_26374,N_21160,N_22937);
nand U26375 (N_26375,N_22993,N_21749);
nor U26376 (N_26376,N_21925,N_19594);
xor U26377 (N_26377,N_20677,N_23211);
and U26378 (N_26378,N_20530,N_18474);
nand U26379 (N_26379,N_21164,N_19475);
and U26380 (N_26380,N_22429,N_20778);
nor U26381 (N_26381,N_18935,N_20600);
and U26382 (N_26382,N_20502,N_20652);
or U26383 (N_26383,N_20042,N_19662);
or U26384 (N_26384,N_23912,N_22943);
xnor U26385 (N_26385,N_22186,N_20334);
nor U26386 (N_26386,N_21285,N_22721);
nand U26387 (N_26387,N_20705,N_23199);
or U26388 (N_26388,N_19095,N_22800);
and U26389 (N_26389,N_18390,N_23315);
nor U26390 (N_26390,N_21009,N_23935);
nand U26391 (N_26391,N_23733,N_19145);
and U26392 (N_26392,N_20607,N_19706);
or U26393 (N_26393,N_18782,N_19240);
or U26394 (N_26394,N_20388,N_23388);
nand U26395 (N_26395,N_23614,N_21127);
or U26396 (N_26396,N_20417,N_18676);
nor U26397 (N_26397,N_21123,N_20519);
xnor U26398 (N_26398,N_18958,N_19664);
nand U26399 (N_26399,N_21415,N_21497);
and U26400 (N_26400,N_20235,N_19644);
or U26401 (N_26401,N_21636,N_18651);
or U26402 (N_26402,N_20997,N_18422);
xnor U26403 (N_26403,N_21439,N_18999);
xnor U26404 (N_26404,N_18104,N_21421);
or U26405 (N_26405,N_21402,N_22874);
nor U26406 (N_26406,N_19924,N_20756);
nand U26407 (N_26407,N_18940,N_19853);
xnor U26408 (N_26408,N_23926,N_20887);
nand U26409 (N_26409,N_23367,N_20054);
xor U26410 (N_26410,N_18867,N_19176);
nand U26411 (N_26411,N_18508,N_20108);
nand U26412 (N_26412,N_19349,N_23950);
nand U26413 (N_26413,N_19814,N_19048);
or U26414 (N_26414,N_21126,N_21723);
and U26415 (N_26415,N_18802,N_20101);
and U26416 (N_26416,N_22487,N_21648);
nor U26417 (N_26417,N_22558,N_18581);
or U26418 (N_26418,N_22046,N_22407);
xnor U26419 (N_26419,N_20257,N_18387);
or U26420 (N_26420,N_20840,N_18344);
xnor U26421 (N_26421,N_22553,N_22585);
nor U26422 (N_26422,N_20773,N_22990);
xor U26423 (N_26423,N_22704,N_19323);
or U26424 (N_26424,N_21780,N_18192);
nor U26425 (N_26425,N_19418,N_18467);
nand U26426 (N_26426,N_22439,N_18137);
or U26427 (N_26427,N_20369,N_18389);
nor U26428 (N_26428,N_21694,N_18059);
xor U26429 (N_26429,N_19639,N_19274);
xor U26430 (N_26430,N_22262,N_21104);
and U26431 (N_26431,N_21815,N_21500);
or U26432 (N_26432,N_21289,N_19391);
or U26433 (N_26433,N_19478,N_23170);
and U26434 (N_26434,N_21865,N_18275);
nand U26435 (N_26435,N_22624,N_19311);
nand U26436 (N_26436,N_18806,N_23816);
and U26437 (N_26437,N_20839,N_22846);
nand U26438 (N_26438,N_19559,N_20707);
nor U26439 (N_26439,N_23736,N_21165);
nand U26440 (N_26440,N_20272,N_18605);
or U26441 (N_26441,N_18755,N_19574);
nand U26442 (N_26442,N_21378,N_23343);
and U26443 (N_26443,N_20365,N_22939);
xnor U26444 (N_26444,N_18233,N_20719);
xnor U26445 (N_26445,N_21118,N_19628);
nand U26446 (N_26446,N_20633,N_18017);
and U26447 (N_26447,N_20270,N_22876);
nor U26448 (N_26448,N_21243,N_18368);
xnor U26449 (N_26449,N_19732,N_22469);
nor U26450 (N_26450,N_18578,N_21720);
xor U26451 (N_26451,N_19431,N_19243);
nand U26452 (N_26452,N_20038,N_22503);
or U26453 (N_26453,N_21541,N_18825);
nand U26454 (N_26454,N_21789,N_21887);
nand U26455 (N_26455,N_20043,N_23723);
or U26456 (N_26456,N_20919,N_21001);
nor U26457 (N_26457,N_21967,N_19321);
xnor U26458 (N_26458,N_23365,N_19261);
xor U26459 (N_26459,N_22616,N_22313);
or U26460 (N_26460,N_22839,N_20401);
nand U26461 (N_26461,N_19580,N_20570);
or U26462 (N_26462,N_21376,N_18012);
or U26463 (N_26463,N_22915,N_18554);
nand U26464 (N_26464,N_19730,N_19333);
nand U26465 (N_26465,N_23311,N_23572);
nor U26466 (N_26466,N_20002,N_23082);
nor U26467 (N_26467,N_22366,N_18535);
nand U26468 (N_26468,N_19112,N_20024);
nand U26469 (N_26469,N_18101,N_18494);
xor U26470 (N_26470,N_18058,N_19682);
xor U26471 (N_26471,N_20265,N_18158);
and U26472 (N_26472,N_22742,N_21492);
and U26473 (N_26473,N_21122,N_18198);
or U26474 (N_26474,N_19009,N_22878);
nand U26475 (N_26475,N_19496,N_19436);
or U26476 (N_26476,N_23865,N_19518);
xor U26477 (N_26477,N_22611,N_19600);
nor U26478 (N_26478,N_19940,N_22820);
xnor U26479 (N_26479,N_22844,N_18677);
and U26480 (N_26480,N_20610,N_21690);
nor U26481 (N_26481,N_23159,N_23734);
nand U26482 (N_26482,N_20018,N_21759);
nor U26483 (N_26483,N_21629,N_22050);
or U26484 (N_26484,N_20557,N_19411);
nand U26485 (N_26485,N_18250,N_22247);
nor U26486 (N_26486,N_19606,N_20188);
nor U26487 (N_26487,N_20618,N_18653);
nand U26488 (N_26488,N_22604,N_20346);
or U26489 (N_26489,N_18327,N_18403);
and U26490 (N_26490,N_21424,N_19695);
nor U26491 (N_26491,N_19143,N_18213);
xor U26492 (N_26492,N_20556,N_20255);
and U26493 (N_26493,N_22528,N_23481);
and U26494 (N_26494,N_22934,N_22671);
nand U26495 (N_26495,N_21656,N_19865);
and U26496 (N_26496,N_22737,N_23313);
nor U26497 (N_26497,N_19382,N_22304);
nand U26498 (N_26498,N_21934,N_22676);
nand U26499 (N_26499,N_22348,N_23423);
nand U26500 (N_26500,N_23219,N_21095);
or U26501 (N_26501,N_22529,N_19005);
nand U26502 (N_26502,N_23692,N_23652);
nor U26503 (N_26503,N_18757,N_22799);
and U26504 (N_26504,N_19551,N_21159);
nor U26505 (N_26505,N_19630,N_23880);
and U26506 (N_26506,N_19285,N_23840);
nand U26507 (N_26507,N_21700,N_22957);
xnor U26508 (N_26508,N_23243,N_18814);
nand U26509 (N_26509,N_19868,N_20415);
or U26510 (N_26510,N_22771,N_18702);
and U26511 (N_26511,N_23434,N_21042);
xor U26512 (N_26512,N_22038,N_22236);
nor U26513 (N_26513,N_23651,N_21236);
xor U26514 (N_26514,N_18336,N_19239);
nand U26515 (N_26515,N_18918,N_22984);
and U26516 (N_26516,N_21025,N_19441);
nand U26517 (N_26517,N_23825,N_18841);
xnor U26518 (N_26518,N_18931,N_23985);
nand U26519 (N_26519,N_21985,N_20499);
or U26520 (N_26520,N_19482,N_19152);
nand U26521 (N_26521,N_22470,N_21057);
nor U26522 (N_26522,N_18014,N_23419);
nor U26523 (N_26523,N_23397,N_19830);
xnor U26524 (N_26524,N_20532,N_19450);
xor U26525 (N_26525,N_23813,N_18062);
and U26526 (N_26526,N_19063,N_18592);
and U26527 (N_26527,N_18890,N_20626);
nand U26528 (N_26528,N_19669,N_22204);
nand U26529 (N_26529,N_22377,N_18974);
nor U26530 (N_26530,N_20082,N_19648);
xnor U26531 (N_26531,N_20751,N_23661);
or U26532 (N_26532,N_21993,N_23943);
and U26533 (N_26533,N_22392,N_20951);
nor U26534 (N_26534,N_23430,N_21638);
nor U26535 (N_26535,N_22572,N_21119);
nor U26536 (N_26536,N_20333,N_22530);
and U26537 (N_26537,N_22049,N_18687);
nand U26538 (N_26538,N_22345,N_23425);
and U26539 (N_26539,N_18520,N_20856);
nand U26540 (N_26540,N_22666,N_23980);
xnor U26541 (N_26541,N_19029,N_18812);
xnor U26542 (N_26542,N_20533,N_22944);
or U26543 (N_26543,N_18027,N_19959);
or U26544 (N_26544,N_23306,N_23420);
and U26545 (N_26545,N_22292,N_23275);
nor U26546 (N_26546,N_23030,N_18125);
or U26547 (N_26547,N_18489,N_20065);
or U26548 (N_26548,N_19453,N_20478);
nor U26549 (N_26549,N_20715,N_21821);
and U26550 (N_26550,N_22200,N_23435);
xnor U26551 (N_26551,N_21045,N_23630);
or U26552 (N_26552,N_21857,N_20992);
xnor U26553 (N_26553,N_19432,N_19182);
or U26554 (N_26554,N_19871,N_20934);
xor U26555 (N_26555,N_20869,N_20206);
nand U26556 (N_26556,N_20284,N_20380);
nor U26557 (N_26557,N_21504,N_18115);
and U26558 (N_26558,N_21350,N_23359);
or U26559 (N_26559,N_23929,N_20540);
nor U26560 (N_26560,N_23767,N_23494);
or U26561 (N_26561,N_20882,N_23623);
xnor U26562 (N_26562,N_18045,N_22763);
and U26563 (N_26563,N_19609,N_19007);
nor U26564 (N_26564,N_22533,N_20722);
nand U26565 (N_26565,N_21942,N_21617);
xor U26566 (N_26566,N_21076,N_23025);
and U26567 (N_26567,N_19555,N_19408);
or U26568 (N_26568,N_18548,N_20377);
and U26569 (N_26569,N_18495,N_20309);
nand U26570 (N_26570,N_20019,N_20165);
or U26571 (N_26571,N_18796,N_19348);
or U26572 (N_26572,N_19919,N_23504);
nor U26573 (N_26573,N_22305,N_22821);
and U26574 (N_26574,N_22426,N_22738);
nand U26575 (N_26575,N_21706,N_23893);
nand U26576 (N_26576,N_18761,N_22980);
nand U26577 (N_26577,N_21665,N_22346);
xnor U26578 (N_26578,N_21675,N_18112);
xnor U26579 (N_26579,N_19420,N_20016);
and U26580 (N_26580,N_23361,N_23618);
xor U26581 (N_26581,N_21496,N_19916);
or U26582 (N_26582,N_19477,N_20287);
nand U26583 (N_26583,N_18975,N_20536);
nor U26584 (N_26584,N_20893,N_21063);
xor U26585 (N_26585,N_20352,N_21189);
or U26586 (N_26586,N_20877,N_23783);
or U26587 (N_26587,N_21946,N_18553);
nor U26588 (N_26588,N_19514,N_19756);
nor U26589 (N_26589,N_21290,N_23569);
xor U26590 (N_26590,N_23919,N_22803);
nand U26591 (N_26591,N_21812,N_21371);
and U26592 (N_26592,N_21850,N_22123);
or U26593 (N_26593,N_18543,N_22898);
xor U26594 (N_26594,N_21900,N_18193);
or U26595 (N_26595,N_20161,N_23183);
and U26596 (N_26596,N_18235,N_18155);
xnor U26597 (N_26597,N_22860,N_20625);
nor U26598 (N_26598,N_23432,N_22177);
or U26599 (N_26599,N_18203,N_22296);
and U26600 (N_26600,N_18147,N_19113);
xor U26601 (N_26601,N_18196,N_19119);
and U26602 (N_26602,N_19485,N_23769);
nand U26603 (N_26603,N_21770,N_22971);
nand U26604 (N_26604,N_22921,N_22573);
or U26605 (N_26605,N_19615,N_20336);
and U26606 (N_26606,N_23399,N_18625);
nor U26607 (N_26607,N_23332,N_21351);
nand U26608 (N_26608,N_23751,N_22601);
xnor U26609 (N_26609,N_19312,N_19497);
nand U26610 (N_26610,N_20189,N_23860);
nor U26611 (N_26611,N_18502,N_20411);
or U26612 (N_26612,N_21413,N_23444);
nor U26613 (N_26613,N_20009,N_18714);
or U26614 (N_26614,N_18692,N_18003);
nand U26615 (N_26615,N_20604,N_21653);
nand U26616 (N_26616,N_22226,N_20220);
nand U26617 (N_26617,N_23527,N_21085);
nor U26618 (N_26618,N_18910,N_22767);
or U26619 (N_26619,N_21943,N_23317);
nor U26620 (N_26620,N_22245,N_22758);
and U26621 (N_26621,N_21790,N_22306);
xor U26622 (N_26622,N_18684,N_18642);
xor U26623 (N_26623,N_18424,N_18103);
or U26624 (N_26624,N_21357,N_20621);
xnor U26625 (N_26625,N_18992,N_21263);
or U26626 (N_26626,N_22859,N_18282);
nand U26627 (N_26627,N_20979,N_18246);
nor U26628 (N_26628,N_21226,N_20984);
and U26629 (N_26629,N_20176,N_23387);
or U26630 (N_26630,N_21795,N_19990);
or U26631 (N_26631,N_22179,N_20014);
nor U26632 (N_26632,N_18790,N_20153);
xor U26633 (N_26633,N_21579,N_23603);
or U26634 (N_26634,N_23700,N_22494);
xor U26635 (N_26635,N_19020,N_23060);
or U26636 (N_26636,N_18143,N_20218);
and U26637 (N_26637,N_23942,N_22909);
nand U26638 (N_26638,N_21280,N_22833);
xnor U26639 (N_26639,N_23272,N_19535);
or U26640 (N_26640,N_21949,N_21920);
xnor U26641 (N_26641,N_19645,N_20923);
xnor U26642 (N_26642,N_22510,N_20222);
and U26643 (N_26643,N_20229,N_18936);
nand U26644 (N_26644,N_18277,N_22340);
xnor U26645 (N_26645,N_23873,N_19067);
nor U26646 (N_26646,N_20860,N_22248);
or U26647 (N_26647,N_23115,N_19389);
xor U26648 (N_26648,N_19480,N_18396);
xnor U26649 (N_26649,N_23038,N_23508);
or U26650 (N_26650,N_18162,N_21660);
nor U26651 (N_26651,N_22747,N_20905);
nand U26652 (N_26652,N_22318,N_19407);
or U26653 (N_26653,N_23489,N_22770);
and U26654 (N_26654,N_22412,N_20699);
xor U26655 (N_26655,N_20606,N_18624);
nand U26656 (N_26656,N_21757,N_23900);
nor U26657 (N_26657,N_23380,N_21811);
and U26658 (N_26658,N_23593,N_18307);
nor U26659 (N_26659,N_19039,N_22968);
nand U26660 (N_26660,N_22445,N_22128);
xor U26661 (N_26661,N_21149,N_19728);
nand U26662 (N_26662,N_23411,N_18564);
xnor U26663 (N_26663,N_23354,N_23792);
nor U26664 (N_26664,N_18997,N_21566);
nand U26665 (N_26665,N_19696,N_21568);
nor U26666 (N_26666,N_23861,N_20809);
xor U26667 (N_26667,N_19957,N_18713);
xor U26668 (N_26668,N_22261,N_21271);
xnor U26669 (N_26669,N_19093,N_19154);
nor U26670 (N_26670,N_22617,N_18756);
xnor U26671 (N_26671,N_19708,N_20356);
or U26672 (N_26672,N_22119,N_23083);
and U26673 (N_26673,N_21143,N_23811);
nor U26674 (N_26674,N_21828,N_22332);
and U26675 (N_26675,N_22146,N_20961);
xnor U26676 (N_26676,N_19501,N_20792);
nor U26677 (N_26677,N_23473,N_21472);
or U26678 (N_26678,N_22903,N_23960);
or U26679 (N_26679,N_21898,N_21134);
nand U26680 (N_26680,N_22781,N_21851);
nor U26681 (N_26681,N_20245,N_18628);
or U26682 (N_26682,N_18266,N_19155);
and U26683 (N_26683,N_23484,N_20006);
and U26684 (N_26684,N_22325,N_19539);
xor U26685 (N_26685,N_18603,N_21245);
and U26686 (N_26686,N_20955,N_18885);
nor U26687 (N_26687,N_20814,N_23220);
and U26688 (N_26688,N_21426,N_18509);
or U26689 (N_26689,N_22307,N_20522);
and U26690 (N_26690,N_20729,N_23080);
xor U26691 (N_26691,N_23776,N_21775);
or U26692 (N_26692,N_23278,N_18264);
xor U26693 (N_26693,N_19292,N_23174);
xor U26694 (N_26694,N_22357,N_21885);
xor U26695 (N_26695,N_22252,N_22156);
or U26696 (N_26696,N_22761,N_23366);
and U26697 (N_26697,N_18251,N_19040);
and U26698 (N_26698,N_20298,N_20672);
nand U26699 (N_26699,N_19318,N_23206);
or U26700 (N_26700,N_23730,N_23678);
nand U26701 (N_26701,N_20487,N_21091);
xnor U26702 (N_26702,N_22690,N_22141);
and U26703 (N_26703,N_18114,N_21663);
nor U26704 (N_26704,N_20350,N_22965);
and U26705 (N_26705,N_21948,N_21398);
nand U26706 (N_26706,N_23389,N_21332);
or U26707 (N_26707,N_20437,N_18587);
nand U26708 (N_26708,N_21180,N_21829);
or U26709 (N_26709,N_22221,N_18285);
nor U26710 (N_26710,N_20185,N_19899);
and U26711 (N_26711,N_19778,N_18455);
or U26712 (N_26712,N_19167,N_22925);
or U26713 (N_26713,N_23409,N_19115);
nor U26714 (N_26714,N_20256,N_18473);
nand U26715 (N_26715,N_23235,N_19667);
and U26716 (N_26716,N_23106,N_21105);
or U26717 (N_26717,N_20730,N_23013);
and U26718 (N_26718,N_18661,N_21227);
or U26719 (N_26719,N_18464,N_18480);
nand U26720 (N_26720,N_18572,N_19659);
nor U26721 (N_26721,N_19836,N_21551);
xnor U26722 (N_26722,N_22316,N_22034);
or U26723 (N_26723,N_22016,N_22230);
and U26724 (N_26724,N_23499,N_22191);
and U26725 (N_26725,N_23057,N_19490);
xor U26726 (N_26726,N_23621,N_20554);
xor U26727 (N_26727,N_22386,N_20806);
and U26728 (N_26728,N_22026,N_18142);
nand U26729 (N_26729,N_21686,N_23155);
and U26730 (N_26730,N_21468,N_19295);
nor U26731 (N_26731,N_19245,N_21407);
and U26732 (N_26732,N_20193,N_22451);
and U26733 (N_26733,N_21182,N_22341);
and U26734 (N_26734,N_20861,N_20339);
and U26735 (N_26735,N_18839,N_20543);
xor U26736 (N_26736,N_19554,N_21540);
and U26737 (N_26737,N_19317,N_19750);
nor U26738 (N_26738,N_22869,N_23905);
or U26739 (N_26739,N_22989,N_18871);
nor U26740 (N_26740,N_21515,N_21833);
or U26741 (N_26741,N_19663,N_22682);
nor U26742 (N_26742,N_21610,N_18688);
nand U26743 (N_26743,N_21432,N_18750);
nor U26744 (N_26744,N_23322,N_23320);
or U26745 (N_26745,N_21858,N_20688);
and U26746 (N_26746,N_21567,N_20864);
xor U26747 (N_26747,N_18780,N_21731);
or U26748 (N_26748,N_20422,N_23501);
and U26749 (N_26749,N_19605,N_18941);
and U26750 (N_26750,N_18083,N_18202);
nor U26751 (N_26751,N_18499,N_23194);
nand U26752 (N_26752,N_20783,N_22641);
or U26753 (N_26753,N_22280,N_21941);
or U26754 (N_26754,N_23848,N_22647);
and U26755 (N_26755,N_23600,N_19541);
or U26756 (N_26756,N_20404,N_21158);
xor U26757 (N_26757,N_22196,N_23323);
or U26758 (N_26758,N_21348,N_20138);
nand U26759 (N_26759,N_21392,N_21701);
nor U26760 (N_26760,N_22825,N_23809);
nand U26761 (N_26761,N_18834,N_21907);
nand U26762 (N_26762,N_18912,N_20559);
xor U26763 (N_26763,N_21102,N_18451);
xnor U26764 (N_26764,N_22290,N_21753);
xnor U26765 (N_26765,N_19603,N_22430);
nand U26766 (N_26766,N_21037,N_20456);
nand U26767 (N_26767,N_20459,N_19704);
and U26768 (N_26768,N_22546,N_23341);
nand U26769 (N_26769,N_20390,N_22862);
nand U26770 (N_26770,N_23517,N_22622);
nand U26771 (N_26771,N_21097,N_19616);
nor U26772 (N_26772,N_22364,N_18256);
xnor U26773 (N_26773,N_23964,N_19558);
nor U26774 (N_26774,N_18228,N_19089);
xor U26775 (N_26775,N_19000,N_22061);
or U26776 (N_26776,N_20940,N_21411);
nand U26777 (N_26777,N_23262,N_19140);
and U26778 (N_26778,N_18876,N_20345);
xnor U26779 (N_26779,N_21187,N_18519);
and U26780 (N_26780,N_21978,N_20669);
nor U26781 (N_26781,N_23327,N_23438);
or U26782 (N_26782,N_20844,N_23213);
nand U26783 (N_26783,N_20712,N_22270);
xnor U26784 (N_26784,N_18219,N_23299);
and U26785 (N_26785,N_18896,N_21011);
or U26786 (N_26786,N_23953,N_21442);
and U26787 (N_26787,N_20226,N_19238);
xnor U26788 (N_26788,N_22615,N_21495);
xor U26789 (N_26789,N_18640,N_22481);
and U26790 (N_26790,N_20507,N_19612);
nand U26791 (N_26791,N_23509,N_19494);
nor U26792 (N_26792,N_18744,N_21799);
or U26793 (N_26793,N_18745,N_23176);
xor U26794 (N_26794,N_20684,N_23523);
xnor U26795 (N_26795,N_19835,N_21666);
xnor U26796 (N_26796,N_21529,N_20960);
nor U26797 (N_26797,N_21625,N_20337);
or U26798 (N_26798,N_23202,N_18922);
or U26799 (N_26799,N_21224,N_18585);
nor U26800 (N_26800,N_20851,N_18320);
and U26801 (N_26801,N_22625,N_23528);
nand U26802 (N_26802,N_23599,N_19221);
and U26803 (N_26803,N_20349,N_19782);
and U26804 (N_26804,N_19026,N_19283);
nor U26805 (N_26805,N_19396,N_20538);
nor U26806 (N_26806,N_21132,N_19366);
nand U26807 (N_26807,N_23558,N_23562);
nand U26808 (N_26808,N_19227,N_18441);
nand U26809 (N_26809,N_23490,N_20447);
nor U26810 (N_26810,N_19316,N_19611);
nor U26811 (N_26811,N_21476,N_20367);
nand U26812 (N_26812,N_18842,N_21142);
xnor U26813 (N_26813,N_22769,N_19608);
nand U26814 (N_26814,N_19479,N_23178);
nand U26815 (N_26815,N_20750,N_20372);
nand U26816 (N_26816,N_20410,N_18659);
or U26817 (N_26817,N_18715,N_23748);
nand U26818 (N_26818,N_22127,N_18224);
and U26819 (N_26819,N_22074,N_19253);
nor U26820 (N_26820,N_18472,N_19058);
xor U26821 (N_26821,N_22143,N_19339);
or U26822 (N_26822,N_21671,N_20592);
xnor U26823 (N_26823,N_23291,N_20725);
xnor U26824 (N_26824,N_21819,N_22596);
or U26825 (N_26825,N_21996,N_23144);
and U26826 (N_26826,N_21397,N_19179);
nor U26827 (N_26827,N_23812,N_22153);
nand U26828 (N_26828,N_22910,N_19729);
or U26829 (N_26829,N_19862,N_19689);
xor U26830 (N_26830,N_22488,N_19547);
and U26831 (N_26831,N_23779,N_18135);
and U26832 (N_26832,N_19372,N_19700);
nor U26833 (N_26833,N_22013,N_18515);
or U26834 (N_26834,N_20286,N_20704);
or U26835 (N_26835,N_20544,N_20052);
nand U26836 (N_26836,N_20795,N_23193);
nand U26837 (N_26837,N_21956,N_19707);
nor U26838 (N_26838,N_19804,N_19954);
nand U26839 (N_26839,N_22139,N_20425);
nor U26840 (N_26840,N_22638,N_23722);
or U26841 (N_26841,N_23876,N_21677);
nor U26842 (N_26842,N_23427,N_21456);
xor U26843 (N_26843,N_20753,N_19711);
and U26844 (N_26844,N_22093,N_21758);
and U26845 (N_26845,N_21886,N_22489);
xor U26846 (N_26846,N_20853,N_23981);
nor U26847 (N_26847,N_20472,N_20288);
and U26848 (N_26848,N_21535,N_21834);
nand U26849 (N_26849,N_19520,N_23654);
nor U26850 (N_26850,N_19680,N_21727);
or U26851 (N_26851,N_21872,N_23298);
and U26852 (N_26852,N_22027,N_18915);
and U26853 (N_26853,N_22571,N_18670);
and U26854 (N_26854,N_21618,N_18032);
nor U26855 (N_26855,N_20129,N_19210);
nor U26856 (N_26856,N_23198,N_19709);
and U26857 (N_26857,N_22145,N_19992);
or U26858 (N_26858,N_21382,N_20894);
and U26859 (N_26859,N_21724,N_19013);
nor U26860 (N_26860,N_23515,N_19217);
nand U26861 (N_26861,N_23314,N_21952);
xor U26862 (N_26862,N_19069,N_21810);
nor U26863 (N_26863,N_18466,N_21140);
nor U26864 (N_26864,N_21317,N_23940);
xor U26865 (N_26865,N_19998,N_18420);
and U26866 (N_26866,N_20999,N_20177);
xnor U26867 (N_26867,N_23321,N_20888);
nand U26868 (N_26868,N_19380,N_19153);
nand U26869 (N_26869,N_19353,N_20711);
nand U26870 (N_26870,N_23685,N_18697);
and U26871 (N_26871,N_21842,N_18299);
nor U26872 (N_26872,N_20384,N_20078);
and U26873 (N_26873,N_19275,N_18102);
and U26874 (N_26874,N_19624,N_20749);
nor U26875 (N_26875,N_21028,N_22536);
nor U26876 (N_26876,N_20754,N_20897);
and U26877 (N_26877,N_19082,N_20539);
nand U26878 (N_26878,N_19328,N_20949);
nor U26879 (N_26879,N_21428,N_23274);
nand U26880 (N_26880,N_22446,N_20944);
nand U26881 (N_26881,N_18770,N_22914);
nand U26882 (N_26882,N_23223,N_23046);
nand U26883 (N_26883,N_21940,N_20702);
nand U26884 (N_26884,N_18479,N_22152);
nand U26885 (N_26885,N_21509,N_18378);
or U26886 (N_26886,N_21883,N_20571);
or U26887 (N_26887,N_22906,N_19806);
xnor U26888 (N_26888,N_20644,N_20501);
xnor U26889 (N_26889,N_22449,N_20589);
nand U26890 (N_26890,N_19102,N_21355);
or U26891 (N_26891,N_20133,N_22275);
xnor U26892 (N_26892,N_23556,N_23979);
nand U26893 (N_26893,N_22277,N_21651);
nor U26894 (N_26894,N_18795,N_21443);
and U26895 (N_26895,N_19237,N_21667);
xor U26896 (N_26896,N_21455,N_18445);
or U26897 (N_26897,N_20675,N_22475);
or U26898 (N_26898,N_21369,N_20382);
or U26899 (N_26899,N_18134,N_21513);
xor U26900 (N_26900,N_19519,N_18939);
and U26901 (N_26901,N_22954,N_21176);
nor U26902 (N_26902,N_21403,N_19556);
and U26903 (N_26903,N_22043,N_23620);
or U26904 (N_26904,N_20251,N_19822);
nor U26905 (N_26905,N_18279,N_20780);
nand U26906 (N_26906,N_18944,N_18868);
xnor U26907 (N_26907,N_23763,N_20221);
nand U26908 (N_26908,N_22009,N_20841);
or U26909 (N_26909,N_22815,N_21107);
nand U26910 (N_26910,N_18920,N_22918);
nor U26911 (N_26911,N_19019,N_18848);
and U26912 (N_26912,N_18712,N_23500);
xnor U26913 (N_26913,N_20912,N_23103);
xor U26914 (N_26914,N_22930,N_19241);
or U26915 (N_26915,N_22017,N_20202);
nand U26916 (N_26916,N_21544,N_22637);
or U26917 (N_26917,N_21408,N_22675);
nor U26918 (N_26918,N_21175,N_23259);
and U26919 (N_26919,N_19049,N_20406);
nand U26920 (N_26920,N_18290,N_19510);
and U26921 (N_26921,N_20764,N_19532);
xor U26922 (N_26922,N_22217,N_18323);
and U26923 (N_26923,N_20473,N_23845);
nor U26924 (N_26924,N_22384,N_18414);
xor U26925 (N_26925,N_18798,N_20933);
xnor U26926 (N_26926,N_21494,N_20596);
or U26927 (N_26927,N_23479,N_22858);
or U26928 (N_26928,N_20506,N_18352);
nand U26929 (N_26929,N_23139,N_22276);
nand U26930 (N_26930,N_18013,N_23398);
nor U26931 (N_26931,N_19942,N_23086);
nand U26932 (N_26932,N_20637,N_19073);
nor U26933 (N_26933,N_19818,N_19367);
xor U26934 (N_26934,N_18319,N_19792);
or U26935 (N_26935,N_22125,N_23694);
and U26936 (N_26936,N_22243,N_19352);
nand U26937 (N_26937,N_21649,N_22591);
nor U26938 (N_26938,N_23373,N_20474);
xnor U26939 (N_26939,N_19591,N_19751);
and U26940 (N_26940,N_19267,N_20207);
nor U26941 (N_26941,N_22932,N_20879);
and U26942 (N_26942,N_21038,N_18483);
and U26943 (N_26943,N_20741,N_22524);
xor U26944 (N_26944,N_23392,N_20171);
and U26945 (N_26945,N_18273,N_20969);
xor U26946 (N_26946,N_19493,N_21772);
nand U26947 (N_26947,N_20755,N_21316);
and U26948 (N_26948,N_21449,N_22162);
or U26949 (N_26949,N_18079,N_19607);
nand U26950 (N_26950,N_19770,N_20925);
nand U26951 (N_26951,N_23948,N_18401);
nor U26952 (N_26952,N_23463,N_23898);
nand U26953 (N_26953,N_21604,N_21623);
nor U26954 (N_26954,N_21615,N_19741);
nor U26955 (N_26955,N_21682,N_19288);
and U26956 (N_26956,N_20458,N_21847);
xnor U26957 (N_26957,N_20686,N_21381);
nor U26958 (N_26958,N_21240,N_20419);
and U26959 (N_26959,N_21484,N_21805);
nor U26960 (N_26960,N_19690,N_19169);
or U26961 (N_26961,N_23253,N_19284);
or U26962 (N_26962,N_19699,N_23729);
and U26963 (N_26963,N_22688,N_19890);
and U26964 (N_26964,N_22725,N_22124);
nor U26965 (N_26965,N_22951,N_18980);
and U26966 (N_26966,N_20983,N_22329);
nor U26967 (N_26967,N_18001,N_20957);
nand U26968 (N_26968,N_23606,N_20026);
and U26969 (N_26969,N_18168,N_19625);
xnor U26970 (N_26970,N_19286,N_22814);
nor U26971 (N_26971,N_21718,N_23666);
or U26972 (N_26972,N_23351,N_18438);
nand U26973 (N_26973,N_23761,N_21837);
xor U26974 (N_26974,N_18496,N_20878);
xnor U26975 (N_26975,N_19646,N_21368);
nor U26976 (N_26976,N_18343,N_21820);
and U26977 (N_26977,N_22037,N_22956);
xnor U26978 (N_26978,N_22515,N_19838);
or U26979 (N_26979,N_23036,N_20599);
and U26980 (N_26980,N_18704,N_21990);
nand U26981 (N_26981,N_21524,N_20562);
nand U26982 (N_26982,N_23158,N_22577);
and U26983 (N_26983,N_23431,N_21573);
nand U26984 (N_26984,N_20071,N_19914);
nand U26985 (N_26985,N_18809,N_19632);
and U26986 (N_26986,N_23386,N_23780);
nand U26987 (N_26987,N_21209,N_20210);
xor U26988 (N_26988,N_23568,N_18963);
nor U26989 (N_26989,N_21787,N_23078);
and U26990 (N_26990,N_23230,N_18272);
or U26991 (N_26991,N_19347,N_18981);
and U26992 (N_26992,N_19854,N_19809);
nand U26993 (N_26993,N_23191,N_21717);
nor U26994 (N_26994,N_21205,N_20978);
xnor U26995 (N_26995,N_19393,N_20498);
and U26996 (N_26996,N_21058,N_22375);
nand U26997 (N_26997,N_22779,N_23765);
nand U26998 (N_26998,N_19440,N_20100);
and U26999 (N_26999,N_18357,N_20087);
xnor U27000 (N_27000,N_21573,N_21276);
nor U27001 (N_27001,N_22023,N_21349);
nand U27002 (N_27002,N_23454,N_18994);
xor U27003 (N_27003,N_22043,N_23949);
and U27004 (N_27004,N_21763,N_20041);
and U27005 (N_27005,N_22168,N_18757);
nand U27006 (N_27006,N_23108,N_20101);
or U27007 (N_27007,N_23507,N_22726);
nor U27008 (N_27008,N_18461,N_19875);
nor U27009 (N_27009,N_20541,N_21229);
or U27010 (N_27010,N_21285,N_23084);
or U27011 (N_27011,N_19831,N_20816);
and U27012 (N_27012,N_20638,N_22167);
nor U27013 (N_27013,N_19441,N_18301);
and U27014 (N_27014,N_22852,N_20908);
xnor U27015 (N_27015,N_18346,N_23189);
nor U27016 (N_27016,N_23701,N_22468);
nor U27017 (N_27017,N_18863,N_19566);
nor U27018 (N_27018,N_23006,N_19310);
nand U27019 (N_27019,N_22714,N_22168);
xnor U27020 (N_27020,N_21497,N_23631);
or U27021 (N_27021,N_20486,N_19071);
nand U27022 (N_27022,N_18825,N_20218);
and U27023 (N_27023,N_18158,N_19254);
and U27024 (N_27024,N_23518,N_23008);
xnor U27025 (N_27025,N_21210,N_19677);
nand U27026 (N_27026,N_20042,N_20104);
nand U27027 (N_27027,N_19400,N_21009);
or U27028 (N_27028,N_18010,N_21744);
and U27029 (N_27029,N_22212,N_19606);
and U27030 (N_27030,N_22983,N_23421);
and U27031 (N_27031,N_21825,N_18295);
nor U27032 (N_27032,N_20762,N_19450);
and U27033 (N_27033,N_18393,N_23794);
and U27034 (N_27034,N_19338,N_18069);
nor U27035 (N_27035,N_22360,N_21358);
or U27036 (N_27036,N_18559,N_20162);
and U27037 (N_27037,N_19255,N_18752);
nor U27038 (N_27038,N_20745,N_21485);
or U27039 (N_27039,N_18444,N_18335);
xor U27040 (N_27040,N_23778,N_23346);
xnor U27041 (N_27041,N_21444,N_22983);
nor U27042 (N_27042,N_23505,N_23518);
and U27043 (N_27043,N_18244,N_21078);
nand U27044 (N_27044,N_19422,N_18917);
xor U27045 (N_27045,N_20771,N_19097);
nand U27046 (N_27046,N_20121,N_19126);
nor U27047 (N_27047,N_23968,N_22005);
or U27048 (N_27048,N_18446,N_21696);
nor U27049 (N_27049,N_22977,N_21601);
nand U27050 (N_27050,N_18099,N_20844);
or U27051 (N_27051,N_18213,N_20948);
nand U27052 (N_27052,N_21567,N_20002);
or U27053 (N_27053,N_22318,N_20025);
xnor U27054 (N_27054,N_20372,N_23552);
and U27055 (N_27055,N_20303,N_21189);
and U27056 (N_27056,N_23214,N_23420);
nor U27057 (N_27057,N_20923,N_20212);
and U27058 (N_27058,N_21633,N_19116);
or U27059 (N_27059,N_20135,N_23551);
and U27060 (N_27060,N_22899,N_18851);
xor U27061 (N_27061,N_23651,N_18337);
xnor U27062 (N_27062,N_18545,N_21155);
and U27063 (N_27063,N_19694,N_23430);
or U27064 (N_27064,N_23497,N_21702);
nor U27065 (N_27065,N_21957,N_19300);
or U27066 (N_27066,N_21569,N_19640);
nor U27067 (N_27067,N_23923,N_21686);
nand U27068 (N_27068,N_20121,N_23006);
and U27069 (N_27069,N_23058,N_18396);
xor U27070 (N_27070,N_19880,N_19966);
and U27071 (N_27071,N_23534,N_18049);
nand U27072 (N_27072,N_21354,N_23752);
xor U27073 (N_27073,N_18387,N_19959);
and U27074 (N_27074,N_20148,N_21670);
or U27075 (N_27075,N_21474,N_19383);
nand U27076 (N_27076,N_21720,N_21484);
nor U27077 (N_27077,N_23216,N_19706);
nand U27078 (N_27078,N_23854,N_23705);
and U27079 (N_27079,N_18913,N_18771);
nand U27080 (N_27080,N_21018,N_18917);
or U27081 (N_27081,N_18816,N_20764);
xor U27082 (N_27082,N_20042,N_18166);
xor U27083 (N_27083,N_23499,N_22918);
nor U27084 (N_27084,N_20324,N_18600);
or U27085 (N_27085,N_20795,N_19365);
xor U27086 (N_27086,N_22965,N_21975);
nand U27087 (N_27087,N_18002,N_22903);
or U27088 (N_27088,N_19401,N_19059);
nand U27089 (N_27089,N_23298,N_22004);
or U27090 (N_27090,N_20923,N_23791);
nor U27091 (N_27091,N_23566,N_21112);
nand U27092 (N_27092,N_18201,N_18738);
nor U27093 (N_27093,N_19130,N_18356);
or U27094 (N_27094,N_22318,N_19679);
and U27095 (N_27095,N_20469,N_23398);
nor U27096 (N_27096,N_18039,N_18273);
xor U27097 (N_27097,N_18760,N_19015);
nand U27098 (N_27098,N_22927,N_20504);
and U27099 (N_27099,N_21723,N_18780);
xor U27100 (N_27100,N_23940,N_22630);
xnor U27101 (N_27101,N_23164,N_21830);
nor U27102 (N_27102,N_19882,N_21381);
nor U27103 (N_27103,N_21997,N_18438);
or U27104 (N_27104,N_23841,N_21157);
nor U27105 (N_27105,N_21068,N_21378);
nand U27106 (N_27106,N_21973,N_19040);
nand U27107 (N_27107,N_22517,N_22383);
nor U27108 (N_27108,N_19673,N_19370);
or U27109 (N_27109,N_22572,N_19467);
xnor U27110 (N_27110,N_22890,N_19865);
nand U27111 (N_27111,N_22517,N_21853);
or U27112 (N_27112,N_19299,N_18538);
or U27113 (N_27113,N_19054,N_21267);
xor U27114 (N_27114,N_19740,N_23511);
and U27115 (N_27115,N_19416,N_18731);
xnor U27116 (N_27116,N_20496,N_23920);
nand U27117 (N_27117,N_18681,N_22996);
nor U27118 (N_27118,N_23971,N_18808);
nor U27119 (N_27119,N_23811,N_18412);
nand U27120 (N_27120,N_19775,N_22917);
nand U27121 (N_27121,N_22822,N_18150);
and U27122 (N_27122,N_19973,N_20406);
or U27123 (N_27123,N_22847,N_20774);
xnor U27124 (N_27124,N_22728,N_22428);
or U27125 (N_27125,N_22705,N_23631);
or U27126 (N_27126,N_18487,N_19703);
xnor U27127 (N_27127,N_20302,N_22541);
nor U27128 (N_27128,N_23803,N_19760);
or U27129 (N_27129,N_20813,N_21391);
xor U27130 (N_27130,N_22268,N_21756);
nand U27131 (N_27131,N_23656,N_22965);
nor U27132 (N_27132,N_21647,N_23930);
or U27133 (N_27133,N_23923,N_18374);
or U27134 (N_27134,N_21148,N_22484);
and U27135 (N_27135,N_21574,N_19941);
xor U27136 (N_27136,N_21297,N_22131);
nand U27137 (N_27137,N_23427,N_19672);
nand U27138 (N_27138,N_21878,N_22877);
nor U27139 (N_27139,N_23172,N_18808);
and U27140 (N_27140,N_19069,N_20507);
nand U27141 (N_27141,N_21107,N_19329);
nor U27142 (N_27142,N_21265,N_19426);
and U27143 (N_27143,N_21497,N_21910);
nand U27144 (N_27144,N_18158,N_22469);
and U27145 (N_27145,N_21834,N_19047);
or U27146 (N_27146,N_20265,N_22465);
nor U27147 (N_27147,N_19040,N_22154);
and U27148 (N_27148,N_20646,N_22166);
nand U27149 (N_27149,N_20582,N_18544);
xor U27150 (N_27150,N_20874,N_20370);
nor U27151 (N_27151,N_19432,N_19610);
xnor U27152 (N_27152,N_18161,N_20410);
xnor U27153 (N_27153,N_21668,N_18070);
or U27154 (N_27154,N_21208,N_20668);
xor U27155 (N_27155,N_18060,N_20548);
and U27156 (N_27156,N_19651,N_22430);
xnor U27157 (N_27157,N_21038,N_19731);
or U27158 (N_27158,N_21789,N_23572);
xor U27159 (N_27159,N_23898,N_20642);
nand U27160 (N_27160,N_22957,N_21896);
or U27161 (N_27161,N_23673,N_23813);
xor U27162 (N_27162,N_20096,N_22598);
xor U27163 (N_27163,N_19988,N_22218);
or U27164 (N_27164,N_18565,N_18219);
nor U27165 (N_27165,N_19028,N_20878);
nand U27166 (N_27166,N_21509,N_22710);
xnor U27167 (N_27167,N_19181,N_19200);
nor U27168 (N_27168,N_20912,N_18253);
or U27169 (N_27169,N_22099,N_20037);
and U27170 (N_27170,N_19139,N_18681);
nand U27171 (N_27171,N_20540,N_18669);
and U27172 (N_27172,N_21161,N_22390);
nor U27173 (N_27173,N_23912,N_18308);
and U27174 (N_27174,N_22803,N_19536);
xnor U27175 (N_27175,N_21695,N_23620);
nand U27176 (N_27176,N_23484,N_18409);
or U27177 (N_27177,N_23497,N_22379);
or U27178 (N_27178,N_20344,N_19031);
nand U27179 (N_27179,N_18914,N_23587);
or U27180 (N_27180,N_18831,N_21519);
nand U27181 (N_27181,N_22433,N_20562);
or U27182 (N_27182,N_22041,N_23858);
and U27183 (N_27183,N_23040,N_22700);
or U27184 (N_27184,N_22868,N_20041);
and U27185 (N_27185,N_22172,N_20381);
and U27186 (N_27186,N_21404,N_18738);
or U27187 (N_27187,N_22900,N_20367);
and U27188 (N_27188,N_18201,N_22131);
nand U27189 (N_27189,N_19420,N_19396);
nor U27190 (N_27190,N_21519,N_19061);
xor U27191 (N_27191,N_19135,N_21223);
nand U27192 (N_27192,N_20833,N_23208);
xnor U27193 (N_27193,N_22015,N_19599);
nor U27194 (N_27194,N_23772,N_23600);
xnor U27195 (N_27195,N_18492,N_19201);
or U27196 (N_27196,N_23661,N_20314);
nand U27197 (N_27197,N_23298,N_18174);
nand U27198 (N_27198,N_18310,N_22209);
or U27199 (N_27199,N_20241,N_20112);
xnor U27200 (N_27200,N_19177,N_20321);
nor U27201 (N_27201,N_23130,N_22994);
nor U27202 (N_27202,N_21655,N_22649);
and U27203 (N_27203,N_22956,N_21199);
and U27204 (N_27204,N_21238,N_23829);
xnor U27205 (N_27205,N_23353,N_19651);
nand U27206 (N_27206,N_20489,N_21665);
or U27207 (N_27207,N_22472,N_18245);
and U27208 (N_27208,N_22822,N_18279);
nor U27209 (N_27209,N_23587,N_19096);
and U27210 (N_27210,N_20783,N_21677);
xnor U27211 (N_27211,N_19499,N_20205);
nand U27212 (N_27212,N_19583,N_18609);
nor U27213 (N_27213,N_19313,N_18150);
nor U27214 (N_27214,N_18510,N_22857);
nor U27215 (N_27215,N_21195,N_20253);
nor U27216 (N_27216,N_20695,N_20120);
nor U27217 (N_27217,N_21280,N_21808);
nor U27218 (N_27218,N_23523,N_22104);
or U27219 (N_27219,N_20442,N_19031);
nand U27220 (N_27220,N_20970,N_18922);
and U27221 (N_27221,N_20055,N_21498);
nand U27222 (N_27222,N_22619,N_23942);
xor U27223 (N_27223,N_22197,N_20112);
xnor U27224 (N_27224,N_22470,N_23304);
nand U27225 (N_27225,N_18611,N_22034);
nor U27226 (N_27226,N_23502,N_18838);
and U27227 (N_27227,N_20900,N_20039);
or U27228 (N_27228,N_20838,N_23628);
nand U27229 (N_27229,N_21446,N_22887);
xnor U27230 (N_27230,N_18102,N_21151);
or U27231 (N_27231,N_23408,N_20671);
and U27232 (N_27232,N_20489,N_21130);
or U27233 (N_27233,N_21387,N_18347);
nor U27234 (N_27234,N_21065,N_22033);
xnor U27235 (N_27235,N_18174,N_22403);
xnor U27236 (N_27236,N_23762,N_21361);
xor U27237 (N_27237,N_21799,N_22438);
or U27238 (N_27238,N_18755,N_19581);
nor U27239 (N_27239,N_23753,N_23945);
and U27240 (N_27240,N_18619,N_22428);
xor U27241 (N_27241,N_23584,N_19546);
and U27242 (N_27242,N_20293,N_20128);
or U27243 (N_27243,N_21462,N_18080);
nand U27244 (N_27244,N_18973,N_22685);
xnor U27245 (N_27245,N_21323,N_18006);
nand U27246 (N_27246,N_18699,N_22060);
nand U27247 (N_27247,N_21367,N_18537);
xor U27248 (N_27248,N_20689,N_20996);
or U27249 (N_27249,N_21214,N_20802);
and U27250 (N_27250,N_19316,N_21013);
nand U27251 (N_27251,N_21642,N_19670);
or U27252 (N_27252,N_21841,N_23334);
nand U27253 (N_27253,N_19706,N_23556);
nor U27254 (N_27254,N_23707,N_19082);
nand U27255 (N_27255,N_21443,N_19340);
xnor U27256 (N_27256,N_18449,N_23302);
or U27257 (N_27257,N_23824,N_23533);
nor U27258 (N_27258,N_23151,N_23635);
xor U27259 (N_27259,N_19588,N_23346);
and U27260 (N_27260,N_19424,N_21210);
nand U27261 (N_27261,N_18386,N_20839);
nand U27262 (N_27262,N_18790,N_20015);
nor U27263 (N_27263,N_23514,N_22088);
xor U27264 (N_27264,N_23512,N_20307);
and U27265 (N_27265,N_22319,N_20081);
xor U27266 (N_27266,N_23668,N_23542);
and U27267 (N_27267,N_18729,N_21951);
nand U27268 (N_27268,N_19311,N_18709);
xor U27269 (N_27269,N_22479,N_19582);
or U27270 (N_27270,N_18181,N_20898);
xnor U27271 (N_27271,N_23500,N_22369);
xnor U27272 (N_27272,N_21613,N_19060);
nand U27273 (N_27273,N_22018,N_23392);
and U27274 (N_27274,N_18139,N_18941);
xor U27275 (N_27275,N_22975,N_19714);
nor U27276 (N_27276,N_18205,N_18974);
and U27277 (N_27277,N_20604,N_23380);
nor U27278 (N_27278,N_19231,N_23581);
nand U27279 (N_27279,N_21574,N_18989);
nor U27280 (N_27280,N_22451,N_23318);
and U27281 (N_27281,N_19788,N_20047);
and U27282 (N_27282,N_18183,N_21302);
and U27283 (N_27283,N_20716,N_22292);
or U27284 (N_27284,N_22566,N_23137);
nor U27285 (N_27285,N_22936,N_19980);
and U27286 (N_27286,N_22488,N_18999);
nor U27287 (N_27287,N_21026,N_19816);
or U27288 (N_27288,N_20492,N_20550);
nor U27289 (N_27289,N_18098,N_19370);
or U27290 (N_27290,N_21527,N_23828);
nand U27291 (N_27291,N_22995,N_22570);
and U27292 (N_27292,N_22091,N_21963);
and U27293 (N_27293,N_20539,N_21637);
nor U27294 (N_27294,N_20331,N_21123);
and U27295 (N_27295,N_23183,N_20277);
xor U27296 (N_27296,N_23694,N_18317);
xor U27297 (N_27297,N_22604,N_19349);
nand U27298 (N_27298,N_20495,N_21184);
nor U27299 (N_27299,N_21833,N_20253);
nor U27300 (N_27300,N_19459,N_18090);
or U27301 (N_27301,N_20137,N_18807);
nor U27302 (N_27302,N_21994,N_20820);
and U27303 (N_27303,N_21577,N_22454);
and U27304 (N_27304,N_23124,N_22524);
and U27305 (N_27305,N_18542,N_20794);
nand U27306 (N_27306,N_20875,N_23300);
nor U27307 (N_27307,N_19694,N_19276);
and U27308 (N_27308,N_19249,N_18672);
xnor U27309 (N_27309,N_18969,N_19556);
nor U27310 (N_27310,N_20746,N_21905);
and U27311 (N_27311,N_21016,N_21882);
or U27312 (N_27312,N_18793,N_22677);
or U27313 (N_27313,N_19304,N_18698);
or U27314 (N_27314,N_20668,N_22996);
or U27315 (N_27315,N_19260,N_22238);
xor U27316 (N_27316,N_20217,N_19570);
nor U27317 (N_27317,N_20314,N_19604);
nor U27318 (N_27318,N_18146,N_19923);
xnor U27319 (N_27319,N_22110,N_19301);
or U27320 (N_27320,N_21275,N_22793);
nor U27321 (N_27321,N_20219,N_23863);
xnor U27322 (N_27322,N_23742,N_23080);
nand U27323 (N_27323,N_22955,N_23407);
or U27324 (N_27324,N_19053,N_18659);
xnor U27325 (N_27325,N_23090,N_20588);
or U27326 (N_27326,N_21134,N_20221);
and U27327 (N_27327,N_22568,N_21927);
or U27328 (N_27328,N_21861,N_18372);
nand U27329 (N_27329,N_21847,N_21330);
nor U27330 (N_27330,N_21346,N_23518);
nand U27331 (N_27331,N_21218,N_22363);
nand U27332 (N_27332,N_20510,N_18683);
xor U27333 (N_27333,N_22498,N_19145);
nand U27334 (N_27334,N_19119,N_21632);
and U27335 (N_27335,N_20761,N_22228);
nor U27336 (N_27336,N_23425,N_18735);
xnor U27337 (N_27337,N_20026,N_22765);
and U27338 (N_27338,N_18190,N_18253);
nor U27339 (N_27339,N_19302,N_23653);
and U27340 (N_27340,N_23531,N_23332);
nor U27341 (N_27341,N_20493,N_18268);
or U27342 (N_27342,N_22779,N_18420);
nand U27343 (N_27343,N_18088,N_21725);
nand U27344 (N_27344,N_20826,N_22216);
nand U27345 (N_27345,N_21280,N_20229);
nand U27346 (N_27346,N_19273,N_23753);
nand U27347 (N_27347,N_20235,N_23256);
or U27348 (N_27348,N_22443,N_20625);
and U27349 (N_27349,N_20438,N_19510);
xor U27350 (N_27350,N_20284,N_22974);
xnor U27351 (N_27351,N_19508,N_23929);
nand U27352 (N_27352,N_18542,N_19144);
and U27353 (N_27353,N_23127,N_18818);
nor U27354 (N_27354,N_23727,N_23665);
nor U27355 (N_27355,N_18587,N_18746);
nor U27356 (N_27356,N_21022,N_21821);
nand U27357 (N_27357,N_23582,N_21662);
nand U27358 (N_27358,N_23782,N_19646);
or U27359 (N_27359,N_19625,N_21917);
nor U27360 (N_27360,N_18528,N_22528);
nand U27361 (N_27361,N_19769,N_23840);
nand U27362 (N_27362,N_23892,N_18048);
nor U27363 (N_27363,N_21507,N_22513);
or U27364 (N_27364,N_23444,N_21599);
xor U27365 (N_27365,N_22684,N_18996);
and U27366 (N_27366,N_18012,N_20694);
nand U27367 (N_27367,N_21527,N_19695);
and U27368 (N_27368,N_23793,N_21417);
xnor U27369 (N_27369,N_18788,N_21309);
nor U27370 (N_27370,N_23096,N_18267);
xor U27371 (N_27371,N_18875,N_19736);
nor U27372 (N_27372,N_21224,N_21302);
or U27373 (N_27373,N_21032,N_23768);
xnor U27374 (N_27374,N_20276,N_19920);
xnor U27375 (N_27375,N_22157,N_21434);
xnor U27376 (N_27376,N_20300,N_20937);
or U27377 (N_27377,N_22405,N_23931);
xnor U27378 (N_27378,N_23898,N_19705);
and U27379 (N_27379,N_21426,N_21013);
or U27380 (N_27380,N_23379,N_20069);
nor U27381 (N_27381,N_20817,N_19357);
and U27382 (N_27382,N_19322,N_20882);
nor U27383 (N_27383,N_20963,N_19841);
nand U27384 (N_27384,N_21844,N_20492);
and U27385 (N_27385,N_22008,N_18175);
xor U27386 (N_27386,N_21800,N_20208);
nand U27387 (N_27387,N_19874,N_18656);
and U27388 (N_27388,N_20859,N_19152);
nor U27389 (N_27389,N_23650,N_20577);
xor U27390 (N_27390,N_22793,N_20803);
and U27391 (N_27391,N_20727,N_22068);
xor U27392 (N_27392,N_18672,N_22641);
or U27393 (N_27393,N_19672,N_22061);
xnor U27394 (N_27394,N_19317,N_22324);
nand U27395 (N_27395,N_23963,N_20477);
or U27396 (N_27396,N_22658,N_19577);
xnor U27397 (N_27397,N_18827,N_19513);
nand U27398 (N_27398,N_22918,N_22398);
xor U27399 (N_27399,N_19077,N_18307);
nand U27400 (N_27400,N_21675,N_21710);
nor U27401 (N_27401,N_19658,N_19763);
nor U27402 (N_27402,N_22917,N_19839);
nand U27403 (N_27403,N_21660,N_23250);
xnor U27404 (N_27404,N_19586,N_23723);
or U27405 (N_27405,N_18541,N_23301);
or U27406 (N_27406,N_21029,N_22138);
xnor U27407 (N_27407,N_20825,N_23195);
and U27408 (N_27408,N_21865,N_19006);
and U27409 (N_27409,N_23843,N_19395);
xnor U27410 (N_27410,N_22691,N_20601);
or U27411 (N_27411,N_18639,N_23709);
and U27412 (N_27412,N_22278,N_23326);
and U27413 (N_27413,N_23041,N_23327);
and U27414 (N_27414,N_20573,N_22459);
nor U27415 (N_27415,N_19461,N_20245);
xnor U27416 (N_27416,N_21241,N_23805);
and U27417 (N_27417,N_20171,N_20734);
or U27418 (N_27418,N_18766,N_20350);
or U27419 (N_27419,N_22432,N_23521);
nor U27420 (N_27420,N_18276,N_20396);
nor U27421 (N_27421,N_19009,N_20213);
nand U27422 (N_27422,N_18213,N_19998);
or U27423 (N_27423,N_19324,N_22729);
or U27424 (N_27424,N_20082,N_19845);
and U27425 (N_27425,N_20619,N_19328);
or U27426 (N_27426,N_23183,N_21537);
nor U27427 (N_27427,N_22882,N_21059);
nand U27428 (N_27428,N_23165,N_21295);
or U27429 (N_27429,N_21325,N_20851);
xor U27430 (N_27430,N_22773,N_18567);
and U27431 (N_27431,N_21893,N_22504);
xnor U27432 (N_27432,N_19328,N_21645);
and U27433 (N_27433,N_22600,N_22958);
or U27434 (N_27434,N_23960,N_21120);
xnor U27435 (N_27435,N_18187,N_22918);
nor U27436 (N_27436,N_18429,N_19719);
and U27437 (N_27437,N_23149,N_22554);
nand U27438 (N_27438,N_18949,N_18555);
or U27439 (N_27439,N_21643,N_23083);
or U27440 (N_27440,N_23130,N_20591);
nand U27441 (N_27441,N_23221,N_22294);
or U27442 (N_27442,N_22422,N_23912);
nand U27443 (N_27443,N_20838,N_21811);
xnor U27444 (N_27444,N_21860,N_19870);
xor U27445 (N_27445,N_21940,N_19697);
xnor U27446 (N_27446,N_19470,N_21387);
nand U27447 (N_27447,N_23661,N_21136);
or U27448 (N_27448,N_19587,N_23832);
nand U27449 (N_27449,N_21725,N_23270);
xnor U27450 (N_27450,N_20860,N_19534);
xnor U27451 (N_27451,N_21828,N_20288);
xor U27452 (N_27452,N_21204,N_20558);
xor U27453 (N_27453,N_20103,N_23801);
xor U27454 (N_27454,N_19863,N_18390);
xor U27455 (N_27455,N_22758,N_23727);
and U27456 (N_27456,N_20638,N_20455);
nor U27457 (N_27457,N_20579,N_21382);
and U27458 (N_27458,N_18411,N_19631);
xor U27459 (N_27459,N_23960,N_21658);
and U27460 (N_27460,N_18729,N_18236);
nand U27461 (N_27461,N_19483,N_21961);
and U27462 (N_27462,N_20467,N_21097);
or U27463 (N_27463,N_18140,N_19474);
xor U27464 (N_27464,N_19262,N_22336);
nand U27465 (N_27465,N_20713,N_23856);
nor U27466 (N_27466,N_20751,N_21837);
xor U27467 (N_27467,N_21515,N_18651);
nor U27468 (N_27468,N_23796,N_19773);
nor U27469 (N_27469,N_20477,N_19567);
nand U27470 (N_27470,N_20854,N_22503);
xor U27471 (N_27471,N_23280,N_18741);
nand U27472 (N_27472,N_18428,N_22907);
nor U27473 (N_27473,N_22382,N_23826);
and U27474 (N_27474,N_18552,N_20713);
nand U27475 (N_27475,N_20197,N_22952);
xnor U27476 (N_27476,N_18625,N_20836);
nand U27477 (N_27477,N_20412,N_20195);
xor U27478 (N_27478,N_21065,N_22262);
nand U27479 (N_27479,N_22056,N_19365);
nand U27480 (N_27480,N_19345,N_23396);
nand U27481 (N_27481,N_21129,N_21493);
or U27482 (N_27482,N_21934,N_22728);
and U27483 (N_27483,N_23846,N_23374);
xor U27484 (N_27484,N_23606,N_22567);
or U27485 (N_27485,N_18995,N_23442);
nor U27486 (N_27486,N_20739,N_20506);
nor U27487 (N_27487,N_19806,N_21453);
xnor U27488 (N_27488,N_18256,N_22019);
xor U27489 (N_27489,N_18178,N_20721);
nand U27490 (N_27490,N_21538,N_23808);
nor U27491 (N_27491,N_23500,N_23370);
and U27492 (N_27492,N_20493,N_22452);
xnor U27493 (N_27493,N_20828,N_22306);
nor U27494 (N_27494,N_23064,N_22913);
nor U27495 (N_27495,N_19498,N_19569);
xnor U27496 (N_27496,N_20670,N_22511);
or U27497 (N_27497,N_18099,N_19602);
xor U27498 (N_27498,N_23838,N_23497);
xor U27499 (N_27499,N_18029,N_18593);
or U27500 (N_27500,N_20154,N_18799);
or U27501 (N_27501,N_21118,N_19738);
nor U27502 (N_27502,N_19537,N_22094);
xnor U27503 (N_27503,N_18643,N_21997);
nand U27504 (N_27504,N_19313,N_19528);
and U27505 (N_27505,N_21336,N_19944);
or U27506 (N_27506,N_23587,N_20594);
or U27507 (N_27507,N_21036,N_23956);
xnor U27508 (N_27508,N_18969,N_19410);
nor U27509 (N_27509,N_23250,N_19336);
and U27510 (N_27510,N_19193,N_18612);
xnor U27511 (N_27511,N_20428,N_20222);
nand U27512 (N_27512,N_22969,N_22851);
or U27513 (N_27513,N_20736,N_18900);
and U27514 (N_27514,N_18928,N_23539);
xnor U27515 (N_27515,N_19717,N_19611);
or U27516 (N_27516,N_23581,N_18825);
xnor U27517 (N_27517,N_23321,N_23625);
or U27518 (N_27518,N_20918,N_18998);
nor U27519 (N_27519,N_22991,N_21269);
nor U27520 (N_27520,N_18819,N_21458);
or U27521 (N_27521,N_23725,N_18645);
xnor U27522 (N_27522,N_18026,N_23169);
nor U27523 (N_27523,N_21778,N_21152);
nor U27524 (N_27524,N_18787,N_19242);
or U27525 (N_27525,N_23816,N_20115);
nand U27526 (N_27526,N_19780,N_19200);
nand U27527 (N_27527,N_18146,N_23853);
nand U27528 (N_27528,N_19851,N_21402);
xnor U27529 (N_27529,N_23626,N_22060);
nor U27530 (N_27530,N_19940,N_23687);
or U27531 (N_27531,N_21256,N_20849);
and U27532 (N_27532,N_19924,N_22789);
nor U27533 (N_27533,N_21726,N_18761);
or U27534 (N_27534,N_20989,N_19681);
nor U27535 (N_27535,N_23814,N_18360);
xor U27536 (N_27536,N_18984,N_20061);
and U27537 (N_27537,N_19650,N_23540);
nand U27538 (N_27538,N_20389,N_20847);
and U27539 (N_27539,N_18317,N_21102);
nor U27540 (N_27540,N_20036,N_18265);
xor U27541 (N_27541,N_21705,N_22406);
xnor U27542 (N_27542,N_23367,N_22028);
and U27543 (N_27543,N_19649,N_20288);
nand U27544 (N_27544,N_20787,N_19946);
and U27545 (N_27545,N_18926,N_18793);
or U27546 (N_27546,N_23969,N_19006);
nand U27547 (N_27547,N_18099,N_23339);
or U27548 (N_27548,N_19277,N_18722);
nor U27549 (N_27549,N_22026,N_21014);
and U27550 (N_27550,N_20091,N_20178);
or U27551 (N_27551,N_23470,N_22052);
nor U27552 (N_27552,N_23126,N_20212);
or U27553 (N_27553,N_18281,N_20704);
and U27554 (N_27554,N_19377,N_23404);
nand U27555 (N_27555,N_21971,N_22174);
nand U27556 (N_27556,N_20945,N_23190);
nand U27557 (N_27557,N_20963,N_22209);
and U27558 (N_27558,N_19774,N_19311);
nand U27559 (N_27559,N_19566,N_22593);
or U27560 (N_27560,N_20165,N_22870);
or U27561 (N_27561,N_21496,N_20128);
nand U27562 (N_27562,N_20418,N_19230);
or U27563 (N_27563,N_18538,N_23192);
xor U27564 (N_27564,N_23964,N_18921);
or U27565 (N_27565,N_19703,N_23425);
and U27566 (N_27566,N_19878,N_20781);
nor U27567 (N_27567,N_20735,N_23255);
or U27568 (N_27568,N_22014,N_22259);
and U27569 (N_27569,N_21596,N_18646);
xnor U27570 (N_27570,N_21285,N_21240);
nand U27571 (N_27571,N_21570,N_21797);
or U27572 (N_27572,N_21191,N_21228);
nor U27573 (N_27573,N_20381,N_23839);
and U27574 (N_27574,N_21147,N_23310);
nor U27575 (N_27575,N_22373,N_20289);
xnor U27576 (N_27576,N_18863,N_18108);
nand U27577 (N_27577,N_18240,N_21736);
or U27578 (N_27578,N_18871,N_22954);
or U27579 (N_27579,N_19113,N_18925);
xnor U27580 (N_27580,N_22799,N_18140);
or U27581 (N_27581,N_20821,N_19942);
nor U27582 (N_27582,N_18536,N_18890);
xor U27583 (N_27583,N_19462,N_19179);
xnor U27584 (N_27584,N_23181,N_19941);
or U27585 (N_27585,N_22591,N_23657);
and U27586 (N_27586,N_23181,N_20127);
and U27587 (N_27587,N_19149,N_20026);
nor U27588 (N_27588,N_19672,N_21077);
nor U27589 (N_27589,N_22432,N_20810);
nand U27590 (N_27590,N_23654,N_18286);
or U27591 (N_27591,N_21942,N_20183);
nand U27592 (N_27592,N_22086,N_21060);
and U27593 (N_27593,N_21933,N_19016);
nor U27594 (N_27594,N_23212,N_18008);
and U27595 (N_27595,N_20824,N_22294);
or U27596 (N_27596,N_23960,N_19715);
and U27597 (N_27597,N_19464,N_21305);
and U27598 (N_27598,N_23304,N_20696);
nand U27599 (N_27599,N_18729,N_22608);
nor U27600 (N_27600,N_23454,N_21085);
or U27601 (N_27601,N_21489,N_20466);
and U27602 (N_27602,N_20826,N_20578);
nor U27603 (N_27603,N_18110,N_22178);
and U27604 (N_27604,N_23460,N_20192);
nand U27605 (N_27605,N_21359,N_19599);
or U27606 (N_27606,N_23996,N_20594);
and U27607 (N_27607,N_18306,N_22285);
xnor U27608 (N_27608,N_21280,N_19197);
xor U27609 (N_27609,N_21228,N_21068);
nand U27610 (N_27610,N_18790,N_19531);
xnor U27611 (N_27611,N_18692,N_23813);
nor U27612 (N_27612,N_21769,N_18830);
or U27613 (N_27613,N_21296,N_21437);
or U27614 (N_27614,N_18524,N_23917);
or U27615 (N_27615,N_19916,N_22156);
xor U27616 (N_27616,N_19441,N_22214);
xnor U27617 (N_27617,N_18720,N_20634);
nand U27618 (N_27618,N_23478,N_23064);
nand U27619 (N_27619,N_19598,N_22995);
or U27620 (N_27620,N_19066,N_22119);
and U27621 (N_27621,N_18107,N_22502);
and U27622 (N_27622,N_22910,N_22475);
or U27623 (N_27623,N_18986,N_22120);
and U27624 (N_27624,N_22379,N_20391);
or U27625 (N_27625,N_23405,N_21151);
xnor U27626 (N_27626,N_19157,N_23181);
xnor U27627 (N_27627,N_18724,N_20310);
or U27628 (N_27628,N_23658,N_21623);
nand U27629 (N_27629,N_22345,N_23049);
and U27630 (N_27630,N_20532,N_22622);
or U27631 (N_27631,N_23519,N_20516);
nand U27632 (N_27632,N_21698,N_20874);
nand U27633 (N_27633,N_23805,N_21481);
nand U27634 (N_27634,N_19868,N_19251);
xor U27635 (N_27635,N_19047,N_21727);
nand U27636 (N_27636,N_22806,N_23671);
and U27637 (N_27637,N_18052,N_22093);
nor U27638 (N_27638,N_22715,N_21196);
xnor U27639 (N_27639,N_19321,N_23901);
nand U27640 (N_27640,N_22368,N_21801);
nor U27641 (N_27641,N_18951,N_23194);
xnor U27642 (N_27642,N_23299,N_19542);
or U27643 (N_27643,N_19048,N_23166);
and U27644 (N_27644,N_19889,N_20837);
nand U27645 (N_27645,N_20260,N_19481);
or U27646 (N_27646,N_20550,N_22224);
and U27647 (N_27647,N_22137,N_23227);
or U27648 (N_27648,N_22230,N_23099);
nor U27649 (N_27649,N_21922,N_21256);
nor U27650 (N_27650,N_20008,N_20316);
nand U27651 (N_27651,N_20929,N_22948);
or U27652 (N_27652,N_20409,N_19228);
nor U27653 (N_27653,N_22113,N_20823);
nand U27654 (N_27654,N_21505,N_20045);
nor U27655 (N_27655,N_18532,N_19666);
nor U27656 (N_27656,N_20293,N_18185);
and U27657 (N_27657,N_21669,N_18048);
or U27658 (N_27658,N_21189,N_18051);
nand U27659 (N_27659,N_19553,N_23641);
xor U27660 (N_27660,N_23395,N_20404);
xor U27661 (N_27661,N_22368,N_21008);
and U27662 (N_27662,N_23132,N_23996);
xnor U27663 (N_27663,N_23576,N_21251);
nand U27664 (N_27664,N_18312,N_20712);
or U27665 (N_27665,N_21190,N_19543);
nand U27666 (N_27666,N_18389,N_19243);
xnor U27667 (N_27667,N_22095,N_20872);
and U27668 (N_27668,N_20554,N_23318);
nor U27669 (N_27669,N_21541,N_22128);
nand U27670 (N_27670,N_23355,N_20245);
xor U27671 (N_27671,N_22422,N_21158);
nand U27672 (N_27672,N_21379,N_21707);
xnor U27673 (N_27673,N_18626,N_23237);
nor U27674 (N_27674,N_18901,N_23869);
and U27675 (N_27675,N_20831,N_23991);
nand U27676 (N_27676,N_20073,N_19087);
nor U27677 (N_27677,N_23552,N_19438);
or U27678 (N_27678,N_22963,N_23508);
nand U27679 (N_27679,N_19322,N_18586);
xor U27680 (N_27680,N_20907,N_23237);
or U27681 (N_27681,N_19179,N_19702);
nand U27682 (N_27682,N_20251,N_19276);
nor U27683 (N_27683,N_19164,N_21053);
nor U27684 (N_27684,N_23859,N_19370);
or U27685 (N_27685,N_22660,N_23335);
xnor U27686 (N_27686,N_19567,N_19419);
and U27687 (N_27687,N_22566,N_18031);
xor U27688 (N_27688,N_18580,N_18222);
nor U27689 (N_27689,N_23802,N_23254);
and U27690 (N_27690,N_19599,N_19811);
nor U27691 (N_27691,N_20473,N_21565);
and U27692 (N_27692,N_19233,N_23507);
xor U27693 (N_27693,N_23885,N_23140);
nor U27694 (N_27694,N_21165,N_19583);
and U27695 (N_27695,N_23739,N_21355);
and U27696 (N_27696,N_19385,N_23117);
and U27697 (N_27697,N_20633,N_18593);
nand U27698 (N_27698,N_18910,N_20211);
xnor U27699 (N_27699,N_22653,N_20663);
or U27700 (N_27700,N_23699,N_23093);
or U27701 (N_27701,N_22871,N_20488);
nor U27702 (N_27702,N_18491,N_18403);
nor U27703 (N_27703,N_22501,N_23876);
nor U27704 (N_27704,N_21472,N_21887);
or U27705 (N_27705,N_22042,N_18718);
nand U27706 (N_27706,N_21119,N_22789);
or U27707 (N_27707,N_18684,N_22619);
and U27708 (N_27708,N_20805,N_21932);
and U27709 (N_27709,N_18260,N_22917);
nand U27710 (N_27710,N_18337,N_19566);
xnor U27711 (N_27711,N_18994,N_21991);
and U27712 (N_27712,N_21736,N_19662);
nand U27713 (N_27713,N_23128,N_18812);
and U27714 (N_27714,N_20768,N_22969);
nand U27715 (N_27715,N_21938,N_20425);
or U27716 (N_27716,N_20630,N_21089);
xor U27717 (N_27717,N_23162,N_21902);
and U27718 (N_27718,N_18646,N_20131);
nor U27719 (N_27719,N_19939,N_19917);
or U27720 (N_27720,N_21651,N_19790);
xor U27721 (N_27721,N_18909,N_22936);
xor U27722 (N_27722,N_18985,N_18620);
xor U27723 (N_27723,N_18474,N_20172);
and U27724 (N_27724,N_19396,N_19099);
or U27725 (N_27725,N_23248,N_23138);
xor U27726 (N_27726,N_20532,N_23294);
and U27727 (N_27727,N_23280,N_21797);
xor U27728 (N_27728,N_20200,N_21449);
xor U27729 (N_27729,N_22075,N_19285);
or U27730 (N_27730,N_21843,N_21457);
or U27731 (N_27731,N_18593,N_22606);
nand U27732 (N_27732,N_23931,N_19513);
nand U27733 (N_27733,N_21021,N_21913);
nand U27734 (N_27734,N_19113,N_19137);
or U27735 (N_27735,N_22583,N_20731);
or U27736 (N_27736,N_18234,N_20886);
and U27737 (N_27737,N_21696,N_23056);
xor U27738 (N_27738,N_19461,N_23155);
xnor U27739 (N_27739,N_22763,N_18679);
and U27740 (N_27740,N_19545,N_20865);
nor U27741 (N_27741,N_23828,N_23429);
nand U27742 (N_27742,N_19024,N_19437);
and U27743 (N_27743,N_20505,N_20807);
and U27744 (N_27744,N_21815,N_18065);
xnor U27745 (N_27745,N_22686,N_19212);
and U27746 (N_27746,N_21973,N_18351);
nor U27747 (N_27747,N_21159,N_20632);
nand U27748 (N_27748,N_18490,N_21658);
and U27749 (N_27749,N_18163,N_20747);
xor U27750 (N_27750,N_20590,N_18181);
nor U27751 (N_27751,N_20343,N_21496);
xor U27752 (N_27752,N_22169,N_20293);
xor U27753 (N_27753,N_20730,N_23757);
xnor U27754 (N_27754,N_20501,N_22709);
nor U27755 (N_27755,N_19524,N_23733);
nand U27756 (N_27756,N_18949,N_21772);
nor U27757 (N_27757,N_18293,N_22782);
and U27758 (N_27758,N_21015,N_22757);
or U27759 (N_27759,N_18061,N_19234);
nand U27760 (N_27760,N_22329,N_19786);
and U27761 (N_27761,N_20696,N_19710);
and U27762 (N_27762,N_19774,N_18041);
or U27763 (N_27763,N_18723,N_23183);
or U27764 (N_27764,N_19681,N_23079);
or U27765 (N_27765,N_19185,N_23170);
nand U27766 (N_27766,N_19089,N_20515);
or U27767 (N_27767,N_21014,N_23424);
nor U27768 (N_27768,N_20761,N_19847);
xnor U27769 (N_27769,N_22688,N_18412);
nor U27770 (N_27770,N_18147,N_22979);
nor U27771 (N_27771,N_20714,N_22966);
xnor U27772 (N_27772,N_19264,N_22138);
or U27773 (N_27773,N_20684,N_20577);
nand U27774 (N_27774,N_20319,N_21194);
xnor U27775 (N_27775,N_22045,N_20695);
and U27776 (N_27776,N_20653,N_19557);
nand U27777 (N_27777,N_20918,N_20224);
nor U27778 (N_27778,N_21629,N_23025);
or U27779 (N_27779,N_21002,N_23653);
and U27780 (N_27780,N_22139,N_20840);
nor U27781 (N_27781,N_23839,N_19267);
xnor U27782 (N_27782,N_18957,N_22532);
nand U27783 (N_27783,N_18871,N_22587);
nand U27784 (N_27784,N_23793,N_20774);
nor U27785 (N_27785,N_23942,N_21278);
xnor U27786 (N_27786,N_22623,N_23471);
or U27787 (N_27787,N_22019,N_20927);
and U27788 (N_27788,N_20026,N_20122);
nand U27789 (N_27789,N_21479,N_22975);
xor U27790 (N_27790,N_19759,N_20823);
nor U27791 (N_27791,N_21500,N_21724);
nand U27792 (N_27792,N_19539,N_22067);
nor U27793 (N_27793,N_20008,N_22369);
and U27794 (N_27794,N_22416,N_19074);
xnor U27795 (N_27795,N_23993,N_23552);
or U27796 (N_27796,N_21730,N_18604);
nor U27797 (N_27797,N_18589,N_18830);
or U27798 (N_27798,N_21671,N_22450);
and U27799 (N_27799,N_22679,N_23196);
xor U27800 (N_27800,N_22372,N_23263);
and U27801 (N_27801,N_20187,N_20472);
and U27802 (N_27802,N_19839,N_19222);
xor U27803 (N_27803,N_20135,N_19911);
or U27804 (N_27804,N_22032,N_21667);
nand U27805 (N_27805,N_19490,N_21146);
xnor U27806 (N_27806,N_20304,N_22787);
and U27807 (N_27807,N_23769,N_23952);
xor U27808 (N_27808,N_20658,N_21809);
nor U27809 (N_27809,N_22852,N_21808);
nand U27810 (N_27810,N_21866,N_19087);
or U27811 (N_27811,N_21941,N_20842);
nand U27812 (N_27812,N_21205,N_19022);
or U27813 (N_27813,N_22461,N_18341);
nor U27814 (N_27814,N_23855,N_21055);
or U27815 (N_27815,N_18050,N_22911);
nand U27816 (N_27816,N_22389,N_22486);
nand U27817 (N_27817,N_18106,N_20467);
nand U27818 (N_27818,N_18331,N_20143);
and U27819 (N_27819,N_19366,N_19561);
nor U27820 (N_27820,N_20115,N_21028);
or U27821 (N_27821,N_20835,N_22190);
xnor U27822 (N_27822,N_18614,N_22425);
nor U27823 (N_27823,N_19459,N_19537);
xor U27824 (N_27824,N_23809,N_18079);
nor U27825 (N_27825,N_20509,N_18206);
nor U27826 (N_27826,N_23514,N_20457);
and U27827 (N_27827,N_23054,N_22956);
or U27828 (N_27828,N_21347,N_18673);
and U27829 (N_27829,N_22416,N_23380);
nor U27830 (N_27830,N_18410,N_19492);
or U27831 (N_27831,N_23309,N_23576);
nand U27832 (N_27832,N_23129,N_20141);
xnor U27833 (N_27833,N_21880,N_19282);
or U27834 (N_27834,N_18087,N_19294);
nor U27835 (N_27835,N_21009,N_23918);
or U27836 (N_27836,N_21187,N_23722);
nand U27837 (N_27837,N_19361,N_19562);
nor U27838 (N_27838,N_23905,N_22393);
or U27839 (N_27839,N_21075,N_21875);
nor U27840 (N_27840,N_18350,N_20776);
or U27841 (N_27841,N_23729,N_22802);
xnor U27842 (N_27842,N_20772,N_18567);
nor U27843 (N_27843,N_20225,N_18418);
nor U27844 (N_27844,N_22443,N_18349);
or U27845 (N_27845,N_22946,N_22219);
nand U27846 (N_27846,N_19810,N_21834);
and U27847 (N_27847,N_21273,N_20173);
xor U27848 (N_27848,N_19352,N_22019);
and U27849 (N_27849,N_22576,N_20602);
and U27850 (N_27850,N_23814,N_20873);
nand U27851 (N_27851,N_18305,N_22481);
nor U27852 (N_27852,N_19214,N_18361);
nand U27853 (N_27853,N_20989,N_18210);
and U27854 (N_27854,N_19163,N_22393);
nor U27855 (N_27855,N_22558,N_22723);
nand U27856 (N_27856,N_23556,N_20958);
nor U27857 (N_27857,N_22217,N_20489);
xnor U27858 (N_27858,N_23285,N_18203);
nand U27859 (N_27859,N_20429,N_19399);
and U27860 (N_27860,N_22259,N_23075);
nand U27861 (N_27861,N_21033,N_19257);
or U27862 (N_27862,N_20671,N_23879);
nor U27863 (N_27863,N_21582,N_21520);
nor U27864 (N_27864,N_21673,N_20839);
nand U27865 (N_27865,N_19587,N_22096);
xor U27866 (N_27866,N_20615,N_20560);
nor U27867 (N_27867,N_21020,N_21813);
nor U27868 (N_27868,N_22805,N_18418);
or U27869 (N_27869,N_18543,N_20863);
nor U27870 (N_27870,N_18836,N_22107);
or U27871 (N_27871,N_21258,N_19016);
xnor U27872 (N_27872,N_21237,N_19960);
xnor U27873 (N_27873,N_18225,N_22415);
or U27874 (N_27874,N_23805,N_22190);
nor U27875 (N_27875,N_21117,N_22888);
or U27876 (N_27876,N_18946,N_23451);
nand U27877 (N_27877,N_21375,N_19352);
and U27878 (N_27878,N_23212,N_22301);
and U27879 (N_27879,N_21299,N_19758);
xnor U27880 (N_27880,N_20596,N_21382);
xor U27881 (N_27881,N_18181,N_23081);
nand U27882 (N_27882,N_19936,N_18872);
nand U27883 (N_27883,N_22236,N_18567);
and U27884 (N_27884,N_23930,N_18192);
or U27885 (N_27885,N_20273,N_20523);
xor U27886 (N_27886,N_19117,N_18134);
and U27887 (N_27887,N_21496,N_21969);
nor U27888 (N_27888,N_19273,N_20120);
nor U27889 (N_27889,N_23595,N_18977);
or U27890 (N_27890,N_18700,N_22854);
nor U27891 (N_27891,N_22331,N_19762);
or U27892 (N_27892,N_22520,N_20176);
nand U27893 (N_27893,N_18796,N_18254);
xnor U27894 (N_27894,N_21218,N_23690);
xor U27895 (N_27895,N_23766,N_19699);
nand U27896 (N_27896,N_18565,N_18887);
and U27897 (N_27897,N_18816,N_19028);
nor U27898 (N_27898,N_19336,N_19699);
xor U27899 (N_27899,N_23895,N_18545);
nor U27900 (N_27900,N_21959,N_20203);
or U27901 (N_27901,N_18859,N_21619);
nand U27902 (N_27902,N_19693,N_18158);
nor U27903 (N_27903,N_23954,N_19566);
and U27904 (N_27904,N_22126,N_22428);
and U27905 (N_27905,N_18335,N_18430);
nand U27906 (N_27906,N_18155,N_23935);
xor U27907 (N_27907,N_23166,N_21630);
nand U27908 (N_27908,N_19137,N_20904);
nor U27909 (N_27909,N_23800,N_23135);
nand U27910 (N_27910,N_18371,N_22549);
nand U27911 (N_27911,N_21062,N_23643);
and U27912 (N_27912,N_21869,N_22298);
and U27913 (N_27913,N_19930,N_20495);
nand U27914 (N_27914,N_20170,N_21192);
nand U27915 (N_27915,N_23924,N_21317);
and U27916 (N_27916,N_22461,N_22208);
and U27917 (N_27917,N_18696,N_19799);
nor U27918 (N_27918,N_19578,N_21260);
nor U27919 (N_27919,N_20357,N_21795);
nor U27920 (N_27920,N_19826,N_22254);
and U27921 (N_27921,N_20453,N_23461);
and U27922 (N_27922,N_20739,N_20540);
and U27923 (N_27923,N_21740,N_22739);
xnor U27924 (N_27924,N_22163,N_21647);
xor U27925 (N_27925,N_18742,N_20112);
nand U27926 (N_27926,N_22392,N_22716);
and U27927 (N_27927,N_23416,N_20171);
xor U27928 (N_27928,N_20762,N_23937);
or U27929 (N_27929,N_23648,N_23024);
nor U27930 (N_27930,N_19252,N_20249);
and U27931 (N_27931,N_23307,N_21065);
and U27932 (N_27932,N_21566,N_20294);
xor U27933 (N_27933,N_22073,N_18718);
or U27934 (N_27934,N_23057,N_23145);
or U27935 (N_27935,N_20723,N_21042);
nand U27936 (N_27936,N_21370,N_19858);
xor U27937 (N_27937,N_18880,N_19890);
xnor U27938 (N_27938,N_19275,N_21373);
xnor U27939 (N_27939,N_22038,N_21744);
nand U27940 (N_27940,N_18830,N_20104);
nor U27941 (N_27941,N_18999,N_23826);
and U27942 (N_27942,N_23621,N_21396);
and U27943 (N_27943,N_23629,N_18271);
or U27944 (N_27944,N_21129,N_22649);
nand U27945 (N_27945,N_18205,N_22706);
xor U27946 (N_27946,N_19830,N_21327);
nand U27947 (N_27947,N_21161,N_18938);
nor U27948 (N_27948,N_20394,N_23534);
or U27949 (N_27949,N_21309,N_23816);
nand U27950 (N_27950,N_18448,N_22601);
xor U27951 (N_27951,N_21559,N_21515);
and U27952 (N_27952,N_18134,N_18221);
nand U27953 (N_27953,N_22888,N_21116);
or U27954 (N_27954,N_18158,N_23187);
nor U27955 (N_27955,N_23778,N_19357);
nor U27956 (N_27956,N_23712,N_23677);
and U27957 (N_27957,N_19553,N_20557);
xor U27958 (N_27958,N_23155,N_21812);
nand U27959 (N_27959,N_22289,N_21241);
nor U27960 (N_27960,N_22147,N_18405);
or U27961 (N_27961,N_23251,N_20114);
nor U27962 (N_27962,N_18664,N_19034);
nand U27963 (N_27963,N_18902,N_18069);
and U27964 (N_27964,N_22799,N_19848);
xnor U27965 (N_27965,N_22711,N_20342);
xor U27966 (N_27966,N_21039,N_21706);
nand U27967 (N_27967,N_21275,N_20392);
xor U27968 (N_27968,N_22180,N_18610);
or U27969 (N_27969,N_18066,N_18774);
xnor U27970 (N_27970,N_21669,N_18839);
or U27971 (N_27971,N_22654,N_22359);
or U27972 (N_27972,N_20483,N_21180);
xnor U27973 (N_27973,N_20547,N_21424);
and U27974 (N_27974,N_22786,N_23467);
nor U27975 (N_27975,N_19542,N_21330);
xor U27976 (N_27976,N_22536,N_21688);
and U27977 (N_27977,N_20872,N_22503);
and U27978 (N_27978,N_19530,N_21903);
or U27979 (N_27979,N_18983,N_22560);
or U27980 (N_27980,N_19753,N_19357);
nand U27981 (N_27981,N_20823,N_22603);
nand U27982 (N_27982,N_21907,N_21513);
nor U27983 (N_27983,N_23331,N_22919);
xor U27984 (N_27984,N_19171,N_18206);
nand U27985 (N_27985,N_22251,N_21485);
or U27986 (N_27986,N_19471,N_20614);
xor U27987 (N_27987,N_23695,N_20263);
or U27988 (N_27988,N_19416,N_23354);
xnor U27989 (N_27989,N_21797,N_18936);
and U27990 (N_27990,N_20449,N_18349);
and U27991 (N_27991,N_19402,N_21158);
or U27992 (N_27992,N_19990,N_22931);
nand U27993 (N_27993,N_20898,N_19690);
nand U27994 (N_27994,N_21230,N_18788);
nand U27995 (N_27995,N_20980,N_21999);
or U27996 (N_27996,N_23271,N_23760);
nand U27997 (N_27997,N_21697,N_21468);
nand U27998 (N_27998,N_21616,N_23317);
xor U27999 (N_27999,N_20750,N_20254);
nor U28000 (N_28000,N_18607,N_21681);
nand U28001 (N_28001,N_23115,N_21499);
and U28002 (N_28002,N_18763,N_23329);
xnor U28003 (N_28003,N_23844,N_21559);
nand U28004 (N_28004,N_19296,N_22555);
or U28005 (N_28005,N_21568,N_20080);
nand U28006 (N_28006,N_21533,N_20064);
nor U28007 (N_28007,N_18269,N_23522);
and U28008 (N_28008,N_23935,N_19921);
nand U28009 (N_28009,N_18676,N_19768);
or U28010 (N_28010,N_22689,N_22834);
or U28011 (N_28011,N_23332,N_23298);
or U28012 (N_28012,N_22379,N_20166);
nand U28013 (N_28013,N_19176,N_21283);
nand U28014 (N_28014,N_23520,N_20189);
and U28015 (N_28015,N_23785,N_18787);
nor U28016 (N_28016,N_20658,N_21127);
or U28017 (N_28017,N_21001,N_20740);
nor U28018 (N_28018,N_21321,N_22201);
nand U28019 (N_28019,N_21652,N_21905);
xnor U28020 (N_28020,N_22979,N_21336);
nand U28021 (N_28021,N_20139,N_20216);
nand U28022 (N_28022,N_19746,N_21142);
or U28023 (N_28023,N_18970,N_19428);
nand U28024 (N_28024,N_19041,N_23429);
nand U28025 (N_28025,N_21303,N_23952);
nand U28026 (N_28026,N_20780,N_21329);
and U28027 (N_28027,N_20269,N_20331);
nand U28028 (N_28028,N_21765,N_20979);
and U28029 (N_28029,N_22576,N_23352);
xor U28030 (N_28030,N_20127,N_20838);
and U28031 (N_28031,N_19761,N_23522);
nor U28032 (N_28032,N_19701,N_22794);
xnor U28033 (N_28033,N_23232,N_19869);
or U28034 (N_28034,N_18927,N_23778);
nand U28035 (N_28035,N_19697,N_22738);
nor U28036 (N_28036,N_23240,N_21483);
xor U28037 (N_28037,N_23043,N_23523);
nor U28038 (N_28038,N_20162,N_19323);
xor U28039 (N_28039,N_21396,N_23267);
or U28040 (N_28040,N_19189,N_18672);
and U28041 (N_28041,N_23306,N_23114);
or U28042 (N_28042,N_18032,N_23334);
and U28043 (N_28043,N_23533,N_23565);
nor U28044 (N_28044,N_18097,N_19971);
or U28045 (N_28045,N_20233,N_21004);
and U28046 (N_28046,N_23261,N_19315);
nor U28047 (N_28047,N_21584,N_19568);
xnor U28048 (N_28048,N_18812,N_18973);
nand U28049 (N_28049,N_18793,N_23975);
or U28050 (N_28050,N_23396,N_22133);
xnor U28051 (N_28051,N_21625,N_19199);
nor U28052 (N_28052,N_22520,N_21066);
nand U28053 (N_28053,N_19663,N_22197);
nor U28054 (N_28054,N_19295,N_19372);
xnor U28055 (N_28055,N_22557,N_19929);
xor U28056 (N_28056,N_18486,N_22423);
nand U28057 (N_28057,N_19558,N_23744);
nor U28058 (N_28058,N_22752,N_22651);
xor U28059 (N_28059,N_18457,N_23042);
xnor U28060 (N_28060,N_21600,N_23619);
nor U28061 (N_28061,N_19193,N_21357);
and U28062 (N_28062,N_19126,N_22409);
nor U28063 (N_28063,N_21080,N_20891);
nand U28064 (N_28064,N_22379,N_22559);
nor U28065 (N_28065,N_21103,N_18371);
nor U28066 (N_28066,N_20031,N_19415);
nor U28067 (N_28067,N_22104,N_19266);
or U28068 (N_28068,N_22876,N_20069);
nor U28069 (N_28069,N_20275,N_22398);
and U28070 (N_28070,N_22497,N_19971);
nor U28071 (N_28071,N_20022,N_23588);
nand U28072 (N_28072,N_22756,N_23055);
nand U28073 (N_28073,N_21664,N_23490);
and U28074 (N_28074,N_22719,N_23216);
nand U28075 (N_28075,N_21944,N_20946);
nand U28076 (N_28076,N_23130,N_23815);
nand U28077 (N_28077,N_22061,N_22272);
and U28078 (N_28078,N_22116,N_20331);
nand U28079 (N_28079,N_23657,N_21112);
xor U28080 (N_28080,N_18363,N_19735);
xor U28081 (N_28081,N_18388,N_22733);
or U28082 (N_28082,N_23014,N_23501);
or U28083 (N_28083,N_20725,N_22179);
nand U28084 (N_28084,N_20742,N_22727);
nand U28085 (N_28085,N_23608,N_23255);
nand U28086 (N_28086,N_22712,N_19153);
nand U28087 (N_28087,N_23654,N_23320);
or U28088 (N_28088,N_19016,N_21650);
nor U28089 (N_28089,N_20135,N_19032);
nor U28090 (N_28090,N_22411,N_21284);
nor U28091 (N_28091,N_22950,N_19677);
and U28092 (N_28092,N_19159,N_23464);
xor U28093 (N_28093,N_19248,N_21031);
nand U28094 (N_28094,N_19604,N_22726);
xnor U28095 (N_28095,N_20533,N_22405);
nor U28096 (N_28096,N_20438,N_19888);
xnor U28097 (N_28097,N_23504,N_19883);
nand U28098 (N_28098,N_22486,N_23538);
nor U28099 (N_28099,N_19271,N_20317);
xnor U28100 (N_28100,N_19127,N_18015);
and U28101 (N_28101,N_20326,N_19770);
xor U28102 (N_28102,N_19665,N_19667);
or U28103 (N_28103,N_22291,N_22007);
or U28104 (N_28104,N_18118,N_23362);
xnor U28105 (N_28105,N_18066,N_20128);
nand U28106 (N_28106,N_20009,N_20849);
nor U28107 (N_28107,N_19782,N_23105);
xnor U28108 (N_28108,N_21156,N_22105);
or U28109 (N_28109,N_19884,N_18250);
xnor U28110 (N_28110,N_22276,N_23582);
or U28111 (N_28111,N_20104,N_18608);
nand U28112 (N_28112,N_18501,N_18905);
or U28113 (N_28113,N_22171,N_23496);
nor U28114 (N_28114,N_21738,N_20988);
and U28115 (N_28115,N_21689,N_19891);
nor U28116 (N_28116,N_19083,N_18399);
and U28117 (N_28117,N_18710,N_19169);
nor U28118 (N_28118,N_21465,N_19114);
nor U28119 (N_28119,N_18140,N_22616);
nand U28120 (N_28120,N_23153,N_21325);
and U28121 (N_28121,N_19080,N_23656);
xnor U28122 (N_28122,N_19053,N_18055);
and U28123 (N_28123,N_22337,N_19422);
nor U28124 (N_28124,N_19112,N_23825);
nand U28125 (N_28125,N_21539,N_18225);
nand U28126 (N_28126,N_18220,N_22782);
and U28127 (N_28127,N_23843,N_18568);
and U28128 (N_28128,N_22468,N_19236);
nor U28129 (N_28129,N_23865,N_20407);
and U28130 (N_28130,N_23677,N_21817);
and U28131 (N_28131,N_23734,N_22524);
and U28132 (N_28132,N_21269,N_20476);
nor U28133 (N_28133,N_18713,N_19569);
xor U28134 (N_28134,N_21075,N_19638);
nor U28135 (N_28135,N_22697,N_19568);
or U28136 (N_28136,N_22774,N_20232);
nand U28137 (N_28137,N_20096,N_23675);
xnor U28138 (N_28138,N_21633,N_23773);
or U28139 (N_28139,N_20129,N_19719);
nand U28140 (N_28140,N_21768,N_18768);
xor U28141 (N_28141,N_22254,N_21596);
nand U28142 (N_28142,N_23504,N_18435);
xor U28143 (N_28143,N_18619,N_23784);
xor U28144 (N_28144,N_21484,N_22497);
xor U28145 (N_28145,N_22671,N_19488);
xor U28146 (N_28146,N_23091,N_21366);
nand U28147 (N_28147,N_23658,N_23568);
nand U28148 (N_28148,N_18323,N_18974);
xor U28149 (N_28149,N_21642,N_18741);
xor U28150 (N_28150,N_20747,N_22352);
xnor U28151 (N_28151,N_20283,N_22569);
xor U28152 (N_28152,N_20552,N_23830);
and U28153 (N_28153,N_22028,N_22534);
nor U28154 (N_28154,N_20472,N_18357);
nor U28155 (N_28155,N_19536,N_18919);
nand U28156 (N_28156,N_20827,N_19364);
and U28157 (N_28157,N_21075,N_19722);
nand U28158 (N_28158,N_20291,N_21092);
and U28159 (N_28159,N_22080,N_18020);
or U28160 (N_28160,N_20803,N_18812);
or U28161 (N_28161,N_22784,N_20575);
and U28162 (N_28162,N_20317,N_22327);
and U28163 (N_28163,N_22156,N_20478);
xor U28164 (N_28164,N_21925,N_18624);
or U28165 (N_28165,N_22032,N_22320);
and U28166 (N_28166,N_23073,N_21143);
or U28167 (N_28167,N_20815,N_18861);
and U28168 (N_28168,N_19380,N_21876);
or U28169 (N_28169,N_19189,N_18698);
nor U28170 (N_28170,N_21579,N_21957);
and U28171 (N_28171,N_23073,N_19447);
and U28172 (N_28172,N_18004,N_18295);
nand U28173 (N_28173,N_21774,N_19910);
and U28174 (N_28174,N_20691,N_23125);
or U28175 (N_28175,N_22898,N_21575);
and U28176 (N_28176,N_18657,N_22215);
nor U28177 (N_28177,N_21589,N_20344);
and U28178 (N_28178,N_22677,N_22545);
xor U28179 (N_28179,N_19642,N_20961);
or U28180 (N_28180,N_20049,N_20745);
xor U28181 (N_28181,N_19125,N_21810);
nor U28182 (N_28182,N_22541,N_23581);
and U28183 (N_28183,N_18952,N_22154);
xnor U28184 (N_28184,N_20417,N_18480);
nor U28185 (N_28185,N_19851,N_20618);
and U28186 (N_28186,N_22333,N_19578);
xnor U28187 (N_28187,N_21712,N_22098);
nand U28188 (N_28188,N_18721,N_20044);
or U28189 (N_28189,N_19888,N_18666);
nor U28190 (N_28190,N_18254,N_22547);
or U28191 (N_28191,N_19075,N_21689);
xor U28192 (N_28192,N_21830,N_21199);
xnor U28193 (N_28193,N_18879,N_20702);
nor U28194 (N_28194,N_18049,N_18510);
xor U28195 (N_28195,N_22637,N_20555);
nand U28196 (N_28196,N_21127,N_23645);
xnor U28197 (N_28197,N_23669,N_21882);
or U28198 (N_28198,N_22077,N_21839);
and U28199 (N_28199,N_23967,N_18580);
nor U28200 (N_28200,N_22777,N_19648);
or U28201 (N_28201,N_22988,N_23159);
nor U28202 (N_28202,N_20909,N_20787);
or U28203 (N_28203,N_19583,N_22277);
nand U28204 (N_28204,N_19226,N_20975);
and U28205 (N_28205,N_19115,N_20340);
xnor U28206 (N_28206,N_21109,N_18247);
xnor U28207 (N_28207,N_23079,N_18561);
or U28208 (N_28208,N_23544,N_23526);
and U28209 (N_28209,N_22387,N_18892);
or U28210 (N_28210,N_20410,N_19817);
nand U28211 (N_28211,N_18907,N_20657);
or U28212 (N_28212,N_19147,N_20095);
and U28213 (N_28213,N_18177,N_21173);
xor U28214 (N_28214,N_22988,N_20720);
nand U28215 (N_28215,N_23525,N_18919);
xor U28216 (N_28216,N_22387,N_18911);
nand U28217 (N_28217,N_21196,N_21733);
nor U28218 (N_28218,N_21716,N_21437);
nor U28219 (N_28219,N_21952,N_23592);
and U28220 (N_28220,N_18522,N_19740);
xnor U28221 (N_28221,N_22075,N_22626);
nor U28222 (N_28222,N_19938,N_20004);
xnor U28223 (N_28223,N_18777,N_20478);
nand U28224 (N_28224,N_23925,N_22741);
nand U28225 (N_28225,N_22419,N_23225);
and U28226 (N_28226,N_21990,N_18542);
xnor U28227 (N_28227,N_22591,N_20749);
nand U28228 (N_28228,N_19994,N_19281);
nand U28229 (N_28229,N_21688,N_18491);
and U28230 (N_28230,N_19217,N_23198);
nand U28231 (N_28231,N_21130,N_18553);
xnor U28232 (N_28232,N_20279,N_20335);
and U28233 (N_28233,N_20660,N_19698);
xor U28234 (N_28234,N_18142,N_19356);
or U28235 (N_28235,N_22186,N_18611);
xor U28236 (N_28236,N_18120,N_21713);
or U28237 (N_28237,N_22726,N_20012);
nand U28238 (N_28238,N_20729,N_20350);
nor U28239 (N_28239,N_20248,N_20484);
and U28240 (N_28240,N_23330,N_21490);
nand U28241 (N_28241,N_20982,N_21131);
or U28242 (N_28242,N_22522,N_22421);
nand U28243 (N_28243,N_23724,N_19688);
nor U28244 (N_28244,N_21127,N_18554);
xnor U28245 (N_28245,N_19471,N_18395);
or U28246 (N_28246,N_22947,N_22311);
or U28247 (N_28247,N_20234,N_23597);
xnor U28248 (N_28248,N_19062,N_21529);
and U28249 (N_28249,N_19496,N_21326);
nand U28250 (N_28250,N_22704,N_20223);
or U28251 (N_28251,N_21130,N_20191);
nand U28252 (N_28252,N_21677,N_23720);
nand U28253 (N_28253,N_18652,N_20815);
nor U28254 (N_28254,N_22718,N_22812);
nor U28255 (N_28255,N_21148,N_23145);
or U28256 (N_28256,N_20210,N_22068);
xnor U28257 (N_28257,N_20301,N_22234);
nand U28258 (N_28258,N_18887,N_23506);
nand U28259 (N_28259,N_21584,N_18395);
or U28260 (N_28260,N_20050,N_18398);
or U28261 (N_28261,N_22341,N_21432);
xnor U28262 (N_28262,N_23389,N_19534);
nor U28263 (N_28263,N_23303,N_21313);
xor U28264 (N_28264,N_20819,N_18249);
xnor U28265 (N_28265,N_18824,N_22082);
nand U28266 (N_28266,N_22658,N_22294);
nand U28267 (N_28267,N_23410,N_22140);
nor U28268 (N_28268,N_18622,N_23822);
nor U28269 (N_28269,N_18391,N_23533);
xnor U28270 (N_28270,N_18085,N_19705);
or U28271 (N_28271,N_23107,N_21488);
or U28272 (N_28272,N_19768,N_22852);
or U28273 (N_28273,N_23422,N_19801);
xnor U28274 (N_28274,N_20750,N_18651);
nand U28275 (N_28275,N_18462,N_20023);
xor U28276 (N_28276,N_23010,N_20532);
or U28277 (N_28277,N_22285,N_19541);
xor U28278 (N_28278,N_21633,N_18184);
nand U28279 (N_28279,N_23686,N_20611);
xnor U28280 (N_28280,N_19254,N_18854);
nand U28281 (N_28281,N_20848,N_23946);
nor U28282 (N_28282,N_23024,N_20475);
or U28283 (N_28283,N_23256,N_22208);
xor U28284 (N_28284,N_21076,N_20163);
xnor U28285 (N_28285,N_18116,N_18795);
nand U28286 (N_28286,N_22775,N_20285);
xnor U28287 (N_28287,N_22222,N_20031);
and U28288 (N_28288,N_20677,N_21472);
nand U28289 (N_28289,N_20556,N_22273);
or U28290 (N_28290,N_18240,N_21235);
and U28291 (N_28291,N_19958,N_19615);
nand U28292 (N_28292,N_22635,N_21274);
or U28293 (N_28293,N_21329,N_18354);
or U28294 (N_28294,N_21171,N_23853);
xnor U28295 (N_28295,N_19831,N_20690);
nor U28296 (N_28296,N_23264,N_18897);
and U28297 (N_28297,N_20591,N_20538);
and U28298 (N_28298,N_19617,N_21988);
or U28299 (N_28299,N_20585,N_20231);
nand U28300 (N_28300,N_21567,N_23937);
nand U28301 (N_28301,N_20434,N_20466);
nor U28302 (N_28302,N_23026,N_19331);
xnor U28303 (N_28303,N_22729,N_20011);
nor U28304 (N_28304,N_21079,N_23401);
and U28305 (N_28305,N_21439,N_20029);
and U28306 (N_28306,N_19709,N_21025);
xor U28307 (N_28307,N_19252,N_21492);
xnor U28308 (N_28308,N_19213,N_20574);
or U28309 (N_28309,N_19445,N_20333);
nor U28310 (N_28310,N_23495,N_21664);
and U28311 (N_28311,N_21137,N_20332);
xor U28312 (N_28312,N_21568,N_22931);
xnor U28313 (N_28313,N_22779,N_22823);
nor U28314 (N_28314,N_23012,N_21897);
nor U28315 (N_28315,N_23670,N_21826);
xor U28316 (N_28316,N_20606,N_20052);
or U28317 (N_28317,N_20128,N_19480);
or U28318 (N_28318,N_21711,N_23322);
and U28319 (N_28319,N_23441,N_19716);
and U28320 (N_28320,N_23032,N_18490);
or U28321 (N_28321,N_19586,N_21336);
nor U28322 (N_28322,N_19226,N_18695);
or U28323 (N_28323,N_21025,N_20719);
or U28324 (N_28324,N_20641,N_23516);
and U28325 (N_28325,N_22860,N_20999);
xor U28326 (N_28326,N_18600,N_21249);
nand U28327 (N_28327,N_22490,N_18322);
nor U28328 (N_28328,N_22083,N_21432);
or U28329 (N_28329,N_20007,N_23235);
nand U28330 (N_28330,N_19543,N_22096);
xnor U28331 (N_28331,N_19113,N_23790);
nand U28332 (N_28332,N_21714,N_19563);
or U28333 (N_28333,N_20783,N_23933);
nor U28334 (N_28334,N_23287,N_19632);
xor U28335 (N_28335,N_19604,N_19587);
or U28336 (N_28336,N_21944,N_22057);
or U28337 (N_28337,N_23860,N_18041);
and U28338 (N_28338,N_23017,N_20337);
or U28339 (N_28339,N_18345,N_23000);
xor U28340 (N_28340,N_22099,N_22161);
xor U28341 (N_28341,N_22448,N_20390);
xor U28342 (N_28342,N_18267,N_20607);
nor U28343 (N_28343,N_18511,N_23833);
or U28344 (N_28344,N_20263,N_20578);
xnor U28345 (N_28345,N_18592,N_20251);
nor U28346 (N_28346,N_21030,N_19576);
nand U28347 (N_28347,N_22504,N_21453);
or U28348 (N_28348,N_20178,N_19015);
xor U28349 (N_28349,N_23482,N_19958);
xnor U28350 (N_28350,N_22521,N_18227);
nand U28351 (N_28351,N_22985,N_22930);
nand U28352 (N_28352,N_23757,N_21138);
nor U28353 (N_28353,N_18833,N_19334);
nand U28354 (N_28354,N_21491,N_21125);
and U28355 (N_28355,N_20101,N_19043);
or U28356 (N_28356,N_20494,N_22281);
xor U28357 (N_28357,N_19338,N_21681);
nand U28358 (N_28358,N_20477,N_21146);
or U28359 (N_28359,N_18881,N_19682);
nand U28360 (N_28360,N_22373,N_22315);
nor U28361 (N_28361,N_21905,N_23237);
and U28362 (N_28362,N_20522,N_18998);
xor U28363 (N_28363,N_22491,N_18720);
xnor U28364 (N_28364,N_23560,N_18094);
and U28365 (N_28365,N_23160,N_22552);
xnor U28366 (N_28366,N_22555,N_22739);
nor U28367 (N_28367,N_22778,N_21858);
xnor U28368 (N_28368,N_21080,N_22796);
or U28369 (N_28369,N_23343,N_22404);
nand U28370 (N_28370,N_18082,N_21490);
xor U28371 (N_28371,N_20318,N_18600);
nand U28372 (N_28372,N_22669,N_19042);
xnor U28373 (N_28373,N_18559,N_21600);
nand U28374 (N_28374,N_20612,N_23537);
or U28375 (N_28375,N_23974,N_19763);
xor U28376 (N_28376,N_23109,N_18664);
nand U28377 (N_28377,N_19519,N_19085);
nand U28378 (N_28378,N_19727,N_19159);
or U28379 (N_28379,N_18071,N_18049);
nor U28380 (N_28380,N_20837,N_21082);
nor U28381 (N_28381,N_22368,N_19121);
nand U28382 (N_28382,N_21897,N_20392);
xnor U28383 (N_28383,N_23454,N_19665);
nor U28384 (N_28384,N_23232,N_20537);
and U28385 (N_28385,N_19095,N_18593);
xor U28386 (N_28386,N_22466,N_18949);
or U28387 (N_28387,N_22075,N_22929);
and U28388 (N_28388,N_21403,N_20574);
xor U28389 (N_28389,N_21003,N_23868);
and U28390 (N_28390,N_18648,N_18382);
xnor U28391 (N_28391,N_19149,N_21741);
xor U28392 (N_28392,N_20865,N_18250);
xnor U28393 (N_28393,N_20844,N_19368);
and U28394 (N_28394,N_23588,N_20131);
nand U28395 (N_28395,N_23176,N_20453);
nand U28396 (N_28396,N_20840,N_23934);
nand U28397 (N_28397,N_20955,N_21340);
xor U28398 (N_28398,N_20309,N_19301);
or U28399 (N_28399,N_18400,N_22563);
or U28400 (N_28400,N_21666,N_19377);
xor U28401 (N_28401,N_23556,N_19458);
xor U28402 (N_28402,N_23015,N_23052);
nor U28403 (N_28403,N_22204,N_20381);
xor U28404 (N_28404,N_19708,N_23154);
xor U28405 (N_28405,N_23492,N_23683);
or U28406 (N_28406,N_21190,N_23247);
nor U28407 (N_28407,N_23400,N_20281);
nor U28408 (N_28408,N_21045,N_20822);
nand U28409 (N_28409,N_18606,N_20534);
or U28410 (N_28410,N_21885,N_20105);
and U28411 (N_28411,N_20642,N_18178);
nor U28412 (N_28412,N_21823,N_21290);
xor U28413 (N_28413,N_20196,N_20756);
and U28414 (N_28414,N_23219,N_21170);
nor U28415 (N_28415,N_19828,N_21039);
or U28416 (N_28416,N_19044,N_22348);
xor U28417 (N_28417,N_19571,N_20099);
and U28418 (N_28418,N_19726,N_23539);
nand U28419 (N_28419,N_23849,N_23539);
xor U28420 (N_28420,N_19497,N_22943);
and U28421 (N_28421,N_21633,N_23347);
nand U28422 (N_28422,N_19021,N_22025);
xor U28423 (N_28423,N_22314,N_19380);
and U28424 (N_28424,N_20195,N_21731);
nor U28425 (N_28425,N_23014,N_18182);
nor U28426 (N_28426,N_19541,N_18522);
nand U28427 (N_28427,N_22613,N_20216);
nand U28428 (N_28428,N_21199,N_19732);
and U28429 (N_28429,N_21628,N_19960);
nand U28430 (N_28430,N_21174,N_18516);
and U28431 (N_28431,N_23525,N_23101);
and U28432 (N_28432,N_22939,N_20074);
or U28433 (N_28433,N_21223,N_19635);
nand U28434 (N_28434,N_23660,N_20214);
and U28435 (N_28435,N_23956,N_19082);
or U28436 (N_28436,N_18618,N_20200);
nand U28437 (N_28437,N_20612,N_21210);
nand U28438 (N_28438,N_22579,N_19259);
xor U28439 (N_28439,N_19038,N_23561);
nor U28440 (N_28440,N_23367,N_23427);
nand U28441 (N_28441,N_18478,N_18193);
and U28442 (N_28442,N_21148,N_18992);
xnor U28443 (N_28443,N_20158,N_22513);
and U28444 (N_28444,N_22964,N_21427);
or U28445 (N_28445,N_22764,N_20225);
nand U28446 (N_28446,N_18314,N_20672);
nand U28447 (N_28447,N_20764,N_23325);
nor U28448 (N_28448,N_21372,N_21860);
nand U28449 (N_28449,N_18891,N_20799);
nor U28450 (N_28450,N_20735,N_19455);
and U28451 (N_28451,N_21319,N_20551);
or U28452 (N_28452,N_23939,N_23132);
nand U28453 (N_28453,N_23317,N_23510);
or U28454 (N_28454,N_19820,N_20516);
nand U28455 (N_28455,N_18814,N_23825);
and U28456 (N_28456,N_19361,N_20311);
and U28457 (N_28457,N_22602,N_22190);
nand U28458 (N_28458,N_18433,N_23526);
nand U28459 (N_28459,N_22991,N_21411);
nor U28460 (N_28460,N_18917,N_18697);
and U28461 (N_28461,N_19724,N_18488);
xnor U28462 (N_28462,N_18889,N_18962);
xor U28463 (N_28463,N_18947,N_19280);
xor U28464 (N_28464,N_19355,N_20480);
xnor U28465 (N_28465,N_19360,N_21903);
nand U28466 (N_28466,N_19988,N_22908);
and U28467 (N_28467,N_21041,N_22456);
nand U28468 (N_28468,N_21114,N_21912);
or U28469 (N_28469,N_22070,N_23308);
nor U28470 (N_28470,N_23510,N_20732);
xor U28471 (N_28471,N_20604,N_21992);
nor U28472 (N_28472,N_21022,N_23678);
xnor U28473 (N_28473,N_18320,N_20647);
or U28474 (N_28474,N_20149,N_21039);
nor U28475 (N_28475,N_19199,N_22426);
and U28476 (N_28476,N_19648,N_18601);
xnor U28477 (N_28477,N_18818,N_22728);
nor U28478 (N_28478,N_19522,N_23836);
and U28479 (N_28479,N_18076,N_20615);
nand U28480 (N_28480,N_23530,N_20469);
nor U28481 (N_28481,N_22217,N_19773);
nor U28482 (N_28482,N_21018,N_19926);
and U28483 (N_28483,N_23369,N_21830);
nor U28484 (N_28484,N_23054,N_23961);
nor U28485 (N_28485,N_22349,N_20238);
nor U28486 (N_28486,N_19310,N_18553);
nand U28487 (N_28487,N_22869,N_19978);
nor U28488 (N_28488,N_19964,N_23770);
nor U28489 (N_28489,N_19969,N_22514);
and U28490 (N_28490,N_19009,N_21456);
xnor U28491 (N_28491,N_23295,N_19309);
nand U28492 (N_28492,N_19321,N_22342);
xnor U28493 (N_28493,N_19653,N_20105);
nand U28494 (N_28494,N_20602,N_23824);
nor U28495 (N_28495,N_20833,N_19087);
xnor U28496 (N_28496,N_22474,N_21960);
nor U28497 (N_28497,N_19747,N_20808);
and U28498 (N_28498,N_22246,N_22613);
nand U28499 (N_28499,N_21531,N_22936);
or U28500 (N_28500,N_22977,N_23165);
nor U28501 (N_28501,N_20486,N_21311);
or U28502 (N_28502,N_23766,N_22543);
nand U28503 (N_28503,N_21511,N_23615);
xor U28504 (N_28504,N_23095,N_23788);
nor U28505 (N_28505,N_20187,N_21913);
and U28506 (N_28506,N_23641,N_21298);
nor U28507 (N_28507,N_22063,N_22707);
nand U28508 (N_28508,N_19014,N_21482);
nor U28509 (N_28509,N_20117,N_20534);
xor U28510 (N_28510,N_23441,N_20206);
and U28511 (N_28511,N_21232,N_18513);
nand U28512 (N_28512,N_22016,N_22322);
xnor U28513 (N_28513,N_19406,N_18507);
and U28514 (N_28514,N_20064,N_19499);
or U28515 (N_28515,N_18712,N_22778);
or U28516 (N_28516,N_23084,N_23519);
and U28517 (N_28517,N_20668,N_23617);
xnor U28518 (N_28518,N_22221,N_21143);
nand U28519 (N_28519,N_22755,N_22792);
or U28520 (N_28520,N_19444,N_19107);
or U28521 (N_28521,N_21989,N_19853);
xor U28522 (N_28522,N_22795,N_23351);
xnor U28523 (N_28523,N_19968,N_23461);
or U28524 (N_28524,N_21753,N_23192);
and U28525 (N_28525,N_21462,N_19918);
nor U28526 (N_28526,N_23739,N_21258);
nor U28527 (N_28527,N_23217,N_20591);
xnor U28528 (N_28528,N_22560,N_20418);
xor U28529 (N_28529,N_21851,N_22179);
nand U28530 (N_28530,N_18447,N_23018);
nor U28531 (N_28531,N_21612,N_21654);
nand U28532 (N_28532,N_22335,N_21928);
or U28533 (N_28533,N_22835,N_22734);
nand U28534 (N_28534,N_21812,N_19219);
xnor U28535 (N_28535,N_19159,N_23871);
nor U28536 (N_28536,N_22173,N_19273);
nand U28537 (N_28537,N_21052,N_22821);
nand U28538 (N_28538,N_22676,N_22246);
nand U28539 (N_28539,N_22133,N_21748);
xor U28540 (N_28540,N_21399,N_21367);
nand U28541 (N_28541,N_21361,N_23996);
xnor U28542 (N_28542,N_19729,N_19106);
or U28543 (N_28543,N_23920,N_20196);
nor U28544 (N_28544,N_18403,N_23082);
xnor U28545 (N_28545,N_22406,N_23397);
or U28546 (N_28546,N_23658,N_21055);
nand U28547 (N_28547,N_21242,N_21002);
and U28548 (N_28548,N_18935,N_21305);
nor U28549 (N_28549,N_18119,N_20666);
nor U28550 (N_28550,N_21405,N_19641);
and U28551 (N_28551,N_22927,N_22226);
or U28552 (N_28552,N_18144,N_21430);
nand U28553 (N_28553,N_19912,N_19868);
or U28554 (N_28554,N_21044,N_22909);
xor U28555 (N_28555,N_20469,N_20942);
nand U28556 (N_28556,N_21588,N_20668);
xnor U28557 (N_28557,N_20017,N_20110);
nor U28558 (N_28558,N_22140,N_21093);
and U28559 (N_28559,N_20322,N_18707);
nor U28560 (N_28560,N_21812,N_23931);
xnor U28561 (N_28561,N_20903,N_22669);
xnor U28562 (N_28562,N_20128,N_20631);
xnor U28563 (N_28563,N_21930,N_18234);
nor U28564 (N_28564,N_18904,N_21568);
and U28565 (N_28565,N_22356,N_23317);
xnor U28566 (N_28566,N_22053,N_19805);
and U28567 (N_28567,N_21345,N_23348);
nor U28568 (N_28568,N_18763,N_19508);
or U28569 (N_28569,N_21445,N_21347);
nor U28570 (N_28570,N_20262,N_19398);
nor U28571 (N_28571,N_18248,N_19204);
and U28572 (N_28572,N_18624,N_20862);
nor U28573 (N_28573,N_23358,N_21496);
xnor U28574 (N_28574,N_21388,N_22192);
and U28575 (N_28575,N_21860,N_18076);
and U28576 (N_28576,N_19317,N_18804);
and U28577 (N_28577,N_23318,N_21537);
xor U28578 (N_28578,N_23636,N_21133);
xnor U28579 (N_28579,N_23566,N_19519);
nor U28580 (N_28580,N_19249,N_23225);
xnor U28581 (N_28581,N_19901,N_21875);
nand U28582 (N_28582,N_22768,N_18610);
or U28583 (N_28583,N_18501,N_23054);
nand U28584 (N_28584,N_20822,N_19068);
nand U28585 (N_28585,N_20138,N_18257);
nand U28586 (N_28586,N_20078,N_20232);
nand U28587 (N_28587,N_18872,N_18392);
or U28588 (N_28588,N_23655,N_18037);
nand U28589 (N_28589,N_23321,N_20532);
nand U28590 (N_28590,N_22724,N_23484);
or U28591 (N_28591,N_23085,N_18426);
nand U28592 (N_28592,N_23088,N_20261);
and U28593 (N_28593,N_23656,N_20415);
and U28594 (N_28594,N_21032,N_23784);
nand U28595 (N_28595,N_20699,N_23478);
nand U28596 (N_28596,N_19439,N_18895);
and U28597 (N_28597,N_20040,N_20478);
and U28598 (N_28598,N_19766,N_22022);
xnor U28599 (N_28599,N_20895,N_21468);
xnor U28600 (N_28600,N_21145,N_23356);
nand U28601 (N_28601,N_19611,N_22428);
xnor U28602 (N_28602,N_21386,N_18179);
xnor U28603 (N_28603,N_21078,N_20246);
nand U28604 (N_28604,N_22430,N_19604);
and U28605 (N_28605,N_19207,N_21407);
nand U28606 (N_28606,N_23454,N_18271);
nor U28607 (N_28607,N_20287,N_22095);
or U28608 (N_28608,N_19757,N_19086);
or U28609 (N_28609,N_23722,N_23581);
or U28610 (N_28610,N_22164,N_21212);
or U28611 (N_28611,N_19561,N_23242);
nor U28612 (N_28612,N_19175,N_18936);
or U28613 (N_28613,N_21781,N_22122);
nor U28614 (N_28614,N_19692,N_21722);
nand U28615 (N_28615,N_20726,N_18527);
xor U28616 (N_28616,N_21065,N_18184);
nand U28617 (N_28617,N_19082,N_22233);
nor U28618 (N_28618,N_18694,N_21685);
nand U28619 (N_28619,N_19959,N_21687);
nand U28620 (N_28620,N_19675,N_23145);
or U28621 (N_28621,N_20700,N_21266);
or U28622 (N_28622,N_18846,N_22554);
xnor U28623 (N_28623,N_18422,N_22516);
nor U28624 (N_28624,N_21958,N_19038);
xnor U28625 (N_28625,N_18573,N_20039);
and U28626 (N_28626,N_21354,N_23417);
nor U28627 (N_28627,N_21397,N_19630);
xor U28628 (N_28628,N_22588,N_20322);
nand U28629 (N_28629,N_22570,N_23527);
or U28630 (N_28630,N_18263,N_22972);
or U28631 (N_28631,N_20201,N_19340);
and U28632 (N_28632,N_22875,N_18326);
or U28633 (N_28633,N_23926,N_18964);
nand U28634 (N_28634,N_22680,N_18710);
and U28635 (N_28635,N_23066,N_23611);
xnor U28636 (N_28636,N_21195,N_18982);
or U28637 (N_28637,N_20309,N_19629);
or U28638 (N_28638,N_22277,N_19653);
or U28639 (N_28639,N_21872,N_23142);
nand U28640 (N_28640,N_23133,N_23837);
nand U28641 (N_28641,N_23106,N_20239);
xor U28642 (N_28642,N_23963,N_23973);
or U28643 (N_28643,N_20219,N_21706);
xnor U28644 (N_28644,N_21029,N_21469);
or U28645 (N_28645,N_23054,N_22497);
nand U28646 (N_28646,N_20195,N_20060);
nor U28647 (N_28647,N_21964,N_20083);
nor U28648 (N_28648,N_18663,N_22431);
nand U28649 (N_28649,N_22826,N_18666);
nor U28650 (N_28650,N_23105,N_22781);
xor U28651 (N_28651,N_18192,N_23387);
nand U28652 (N_28652,N_23474,N_20725);
nor U28653 (N_28653,N_23018,N_20594);
nand U28654 (N_28654,N_21737,N_23005);
or U28655 (N_28655,N_18391,N_22804);
or U28656 (N_28656,N_20416,N_18316);
and U28657 (N_28657,N_19421,N_20827);
or U28658 (N_28658,N_19009,N_21889);
nor U28659 (N_28659,N_19344,N_21026);
and U28660 (N_28660,N_23438,N_22127);
and U28661 (N_28661,N_23066,N_19760);
xor U28662 (N_28662,N_23340,N_21077);
xnor U28663 (N_28663,N_19661,N_19429);
nand U28664 (N_28664,N_20285,N_21667);
nor U28665 (N_28665,N_22756,N_18764);
or U28666 (N_28666,N_21582,N_21474);
and U28667 (N_28667,N_23098,N_19624);
nand U28668 (N_28668,N_19420,N_21047);
and U28669 (N_28669,N_18082,N_20566);
and U28670 (N_28670,N_20880,N_22184);
and U28671 (N_28671,N_18973,N_19686);
nor U28672 (N_28672,N_19239,N_23276);
or U28673 (N_28673,N_21484,N_21298);
xnor U28674 (N_28674,N_21055,N_20253);
nand U28675 (N_28675,N_21377,N_21128);
or U28676 (N_28676,N_21330,N_19424);
nand U28677 (N_28677,N_22407,N_18213);
nor U28678 (N_28678,N_18732,N_19255);
nand U28679 (N_28679,N_21089,N_23250);
nor U28680 (N_28680,N_21014,N_19818);
xor U28681 (N_28681,N_23988,N_23343);
or U28682 (N_28682,N_18799,N_21632);
or U28683 (N_28683,N_22368,N_22661);
and U28684 (N_28684,N_23057,N_21398);
nor U28685 (N_28685,N_21164,N_23542);
or U28686 (N_28686,N_20322,N_22135);
nor U28687 (N_28687,N_22064,N_21535);
xnor U28688 (N_28688,N_18408,N_22938);
or U28689 (N_28689,N_20080,N_23028);
nand U28690 (N_28690,N_18160,N_19698);
or U28691 (N_28691,N_20580,N_23810);
nor U28692 (N_28692,N_21163,N_19142);
xor U28693 (N_28693,N_22154,N_20619);
and U28694 (N_28694,N_18804,N_18199);
nor U28695 (N_28695,N_20421,N_19892);
and U28696 (N_28696,N_19591,N_23721);
and U28697 (N_28697,N_19161,N_19106);
and U28698 (N_28698,N_21113,N_22703);
nand U28699 (N_28699,N_20542,N_20332);
xnor U28700 (N_28700,N_20675,N_18964);
or U28701 (N_28701,N_21595,N_20249);
or U28702 (N_28702,N_20575,N_23635);
or U28703 (N_28703,N_18264,N_22925);
nand U28704 (N_28704,N_21744,N_23573);
and U28705 (N_28705,N_22451,N_21028);
and U28706 (N_28706,N_23998,N_20927);
and U28707 (N_28707,N_19453,N_22955);
nor U28708 (N_28708,N_21839,N_22976);
and U28709 (N_28709,N_20952,N_23001);
or U28710 (N_28710,N_19010,N_22488);
nand U28711 (N_28711,N_18083,N_22055);
and U28712 (N_28712,N_23330,N_18635);
xor U28713 (N_28713,N_22496,N_21601);
xnor U28714 (N_28714,N_23867,N_21649);
nand U28715 (N_28715,N_23422,N_18194);
xnor U28716 (N_28716,N_22010,N_23017);
or U28717 (N_28717,N_20252,N_23425);
nor U28718 (N_28718,N_21125,N_22409);
xor U28719 (N_28719,N_19888,N_19571);
and U28720 (N_28720,N_19575,N_18160);
and U28721 (N_28721,N_21778,N_18234);
nor U28722 (N_28722,N_18335,N_20052);
or U28723 (N_28723,N_18293,N_19904);
nand U28724 (N_28724,N_22784,N_19811);
xor U28725 (N_28725,N_20190,N_18440);
nor U28726 (N_28726,N_22735,N_18433);
or U28727 (N_28727,N_22145,N_23529);
and U28728 (N_28728,N_21206,N_20889);
and U28729 (N_28729,N_21926,N_20125);
nand U28730 (N_28730,N_23150,N_20590);
or U28731 (N_28731,N_18847,N_22641);
nand U28732 (N_28732,N_23930,N_20428);
nor U28733 (N_28733,N_23354,N_23967);
nand U28734 (N_28734,N_19606,N_23388);
or U28735 (N_28735,N_23017,N_21521);
nand U28736 (N_28736,N_18574,N_19751);
or U28737 (N_28737,N_23354,N_18421);
nand U28738 (N_28738,N_23389,N_19280);
xnor U28739 (N_28739,N_22599,N_18378);
xor U28740 (N_28740,N_22359,N_22714);
nand U28741 (N_28741,N_21355,N_21315);
and U28742 (N_28742,N_18346,N_18054);
nand U28743 (N_28743,N_19768,N_20271);
nand U28744 (N_28744,N_20388,N_19848);
and U28745 (N_28745,N_18400,N_21491);
nand U28746 (N_28746,N_20328,N_18950);
nor U28747 (N_28747,N_22281,N_23596);
nor U28748 (N_28748,N_20294,N_18587);
or U28749 (N_28749,N_21136,N_20450);
nand U28750 (N_28750,N_23439,N_23650);
nand U28751 (N_28751,N_18084,N_19074);
xnor U28752 (N_28752,N_18392,N_22082);
and U28753 (N_28753,N_18406,N_18180);
nand U28754 (N_28754,N_19495,N_18295);
and U28755 (N_28755,N_21113,N_19473);
nand U28756 (N_28756,N_20523,N_19676);
or U28757 (N_28757,N_20121,N_22604);
nand U28758 (N_28758,N_20833,N_23270);
and U28759 (N_28759,N_18963,N_22386);
xor U28760 (N_28760,N_22732,N_18012);
nand U28761 (N_28761,N_22419,N_18923);
nand U28762 (N_28762,N_19622,N_23859);
nor U28763 (N_28763,N_19498,N_23874);
and U28764 (N_28764,N_23724,N_23024);
nor U28765 (N_28765,N_23205,N_20882);
nand U28766 (N_28766,N_19365,N_20950);
or U28767 (N_28767,N_19108,N_23209);
nand U28768 (N_28768,N_20832,N_18796);
xor U28769 (N_28769,N_18837,N_20470);
nor U28770 (N_28770,N_23805,N_18187);
or U28771 (N_28771,N_18186,N_18878);
and U28772 (N_28772,N_18317,N_19579);
nor U28773 (N_28773,N_22432,N_22157);
or U28774 (N_28774,N_19204,N_20512);
nor U28775 (N_28775,N_18569,N_20181);
or U28776 (N_28776,N_23524,N_22936);
nor U28777 (N_28777,N_21215,N_18713);
or U28778 (N_28778,N_22375,N_19682);
xnor U28779 (N_28779,N_19988,N_22978);
and U28780 (N_28780,N_20025,N_22416);
and U28781 (N_28781,N_21865,N_20343);
nand U28782 (N_28782,N_23290,N_23716);
nand U28783 (N_28783,N_21393,N_20808);
and U28784 (N_28784,N_19649,N_20698);
or U28785 (N_28785,N_18315,N_21353);
and U28786 (N_28786,N_18729,N_23220);
or U28787 (N_28787,N_22050,N_19477);
nor U28788 (N_28788,N_21221,N_21564);
nor U28789 (N_28789,N_20451,N_20282);
and U28790 (N_28790,N_23178,N_22767);
and U28791 (N_28791,N_20793,N_19226);
and U28792 (N_28792,N_19473,N_20960);
or U28793 (N_28793,N_18044,N_19844);
nor U28794 (N_28794,N_19007,N_18971);
xnor U28795 (N_28795,N_22007,N_22126);
or U28796 (N_28796,N_18929,N_20241);
nor U28797 (N_28797,N_21786,N_19668);
nand U28798 (N_28798,N_20030,N_20814);
nor U28799 (N_28799,N_18862,N_20659);
xnor U28800 (N_28800,N_20518,N_23567);
nand U28801 (N_28801,N_22849,N_20530);
or U28802 (N_28802,N_20473,N_21800);
xor U28803 (N_28803,N_20869,N_22324);
or U28804 (N_28804,N_23068,N_21446);
and U28805 (N_28805,N_21171,N_23998);
xor U28806 (N_28806,N_18328,N_20780);
and U28807 (N_28807,N_18824,N_18112);
nand U28808 (N_28808,N_19455,N_20812);
nand U28809 (N_28809,N_23229,N_21043);
or U28810 (N_28810,N_21241,N_18688);
nor U28811 (N_28811,N_21578,N_22877);
nor U28812 (N_28812,N_20413,N_19895);
nand U28813 (N_28813,N_18030,N_18121);
nor U28814 (N_28814,N_18122,N_21145);
nor U28815 (N_28815,N_18175,N_20738);
or U28816 (N_28816,N_19598,N_21128);
or U28817 (N_28817,N_20520,N_22841);
xor U28818 (N_28818,N_22125,N_18195);
nand U28819 (N_28819,N_18391,N_20163);
xnor U28820 (N_28820,N_19035,N_22723);
and U28821 (N_28821,N_18665,N_20743);
xnor U28822 (N_28822,N_20400,N_23359);
xor U28823 (N_28823,N_18909,N_18798);
nand U28824 (N_28824,N_18471,N_23219);
nand U28825 (N_28825,N_23230,N_21115);
or U28826 (N_28826,N_22403,N_22536);
nor U28827 (N_28827,N_20764,N_21581);
nand U28828 (N_28828,N_19805,N_21974);
and U28829 (N_28829,N_18411,N_20348);
and U28830 (N_28830,N_22626,N_22820);
and U28831 (N_28831,N_23218,N_20640);
or U28832 (N_28832,N_19054,N_20349);
nor U28833 (N_28833,N_21579,N_21240);
or U28834 (N_28834,N_18032,N_19383);
xnor U28835 (N_28835,N_20288,N_22829);
nor U28836 (N_28836,N_20777,N_21308);
xor U28837 (N_28837,N_18599,N_19491);
or U28838 (N_28838,N_21592,N_21170);
xnor U28839 (N_28839,N_22829,N_23964);
and U28840 (N_28840,N_19865,N_21407);
and U28841 (N_28841,N_20902,N_21822);
or U28842 (N_28842,N_20756,N_19266);
and U28843 (N_28843,N_22307,N_22555);
and U28844 (N_28844,N_20182,N_23119);
and U28845 (N_28845,N_18780,N_20056);
nand U28846 (N_28846,N_22186,N_21672);
xor U28847 (N_28847,N_19164,N_20401);
nor U28848 (N_28848,N_18275,N_23227);
or U28849 (N_28849,N_21337,N_22538);
nor U28850 (N_28850,N_21221,N_22507);
and U28851 (N_28851,N_22642,N_18119);
xor U28852 (N_28852,N_23519,N_22435);
and U28853 (N_28853,N_18414,N_21856);
xor U28854 (N_28854,N_20972,N_20426);
or U28855 (N_28855,N_23144,N_22575);
and U28856 (N_28856,N_23377,N_19814);
and U28857 (N_28857,N_18250,N_22288);
nor U28858 (N_28858,N_19825,N_21252);
or U28859 (N_28859,N_22590,N_19753);
and U28860 (N_28860,N_18287,N_21785);
or U28861 (N_28861,N_21949,N_19902);
nor U28862 (N_28862,N_22803,N_22767);
and U28863 (N_28863,N_21218,N_21945);
xnor U28864 (N_28864,N_18093,N_22782);
and U28865 (N_28865,N_23576,N_21831);
xor U28866 (N_28866,N_23239,N_20472);
xor U28867 (N_28867,N_23211,N_21742);
xor U28868 (N_28868,N_23433,N_21916);
xor U28869 (N_28869,N_23100,N_21915);
nand U28870 (N_28870,N_23172,N_21392);
nand U28871 (N_28871,N_18417,N_18638);
nand U28872 (N_28872,N_18542,N_20744);
nor U28873 (N_28873,N_22858,N_18444);
nor U28874 (N_28874,N_20700,N_18430);
and U28875 (N_28875,N_21600,N_18527);
xnor U28876 (N_28876,N_21346,N_18165);
xnor U28877 (N_28877,N_23266,N_19776);
xnor U28878 (N_28878,N_19570,N_18152);
nor U28879 (N_28879,N_20676,N_20138);
and U28880 (N_28880,N_22437,N_18151);
or U28881 (N_28881,N_19628,N_18930);
xor U28882 (N_28882,N_22848,N_21287);
or U28883 (N_28883,N_20557,N_22395);
or U28884 (N_28884,N_21791,N_19629);
or U28885 (N_28885,N_21656,N_21488);
nor U28886 (N_28886,N_22324,N_23034);
xnor U28887 (N_28887,N_21743,N_22811);
nand U28888 (N_28888,N_21432,N_22665);
xnor U28889 (N_28889,N_19567,N_18394);
nor U28890 (N_28890,N_21913,N_23599);
xor U28891 (N_28891,N_18314,N_22779);
nand U28892 (N_28892,N_20338,N_22105);
nor U28893 (N_28893,N_18131,N_21870);
nand U28894 (N_28894,N_22892,N_19643);
and U28895 (N_28895,N_19067,N_21290);
xnor U28896 (N_28896,N_23679,N_22907);
xnor U28897 (N_28897,N_20068,N_18160);
nand U28898 (N_28898,N_19309,N_22817);
nand U28899 (N_28899,N_20048,N_19690);
xnor U28900 (N_28900,N_18538,N_22356);
and U28901 (N_28901,N_21242,N_20847);
xnor U28902 (N_28902,N_23770,N_19310);
xor U28903 (N_28903,N_21054,N_19653);
or U28904 (N_28904,N_19577,N_22705);
or U28905 (N_28905,N_22385,N_23248);
and U28906 (N_28906,N_20013,N_18110);
nor U28907 (N_28907,N_20094,N_22046);
nand U28908 (N_28908,N_21396,N_18466);
nor U28909 (N_28909,N_22467,N_20690);
nor U28910 (N_28910,N_22835,N_18528);
nand U28911 (N_28911,N_19697,N_22033);
nor U28912 (N_28912,N_19267,N_22407);
nor U28913 (N_28913,N_23722,N_18213);
or U28914 (N_28914,N_18202,N_22880);
and U28915 (N_28915,N_19859,N_22854);
nor U28916 (N_28916,N_19057,N_20228);
nand U28917 (N_28917,N_19402,N_23615);
or U28918 (N_28918,N_21568,N_23104);
and U28919 (N_28919,N_20816,N_19362);
nand U28920 (N_28920,N_23042,N_20275);
nand U28921 (N_28921,N_23779,N_22581);
nand U28922 (N_28922,N_18025,N_19775);
xor U28923 (N_28923,N_22377,N_23819);
nand U28924 (N_28924,N_21550,N_23632);
and U28925 (N_28925,N_20908,N_18555);
or U28926 (N_28926,N_18499,N_19699);
and U28927 (N_28927,N_22543,N_21802);
nor U28928 (N_28928,N_21354,N_21301);
nand U28929 (N_28929,N_18289,N_19769);
nand U28930 (N_28930,N_20611,N_20049);
nor U28931 (N_28931,N_22667,N_21262);
xor U28932 (N_28932,N_21144,N_23181);
xor U28933 (N_28933,N_23710,N_20640);
nor U28934 (N_28934,N_21358,N_23121);
or U28935 (N_28935,N_22895,N_21573);
nor U28936 (N_28936,N_20543,N_23572);
xor U28937 (N_28937,N_19703,N_20508);
nor U28938 (N_28938,N_18111,N_19929);
nor U28939 (N_28939,N_21451,N_21523);
or U28940 (N_28940,N_23709,N_22447);
and U28941 (N_28941,N_22729,N_18786);
or U28942 (N_28942,N_22482,N_23146);
or U28943 (N_28943,N_22673,N_21525);
nor U28944 (N_28944,N_22252,N_18590);
nor U28945 (N_28945,N_18938,N_20114);
nand U28946 (N_28946,N_20199,N_23135);
xor U28947 (N_28947,N_19893,N_21407);
and U28948 (N_28948,N_23657,N_21736);
or U28949 (N_28949,N_20988,N_20246);
nor U28950 (N_28950,N_23717,N_19872);
nor U28951 (N_28951,N_22351,N_23545);
nor U28952 (N_28952,N_21293,N_23280);
and U28953 (N_28953,N_23038,N_23860);
xor U28954 (N_28954,N_18517,N_18224);
nor U28955 (N_28955,N_23434,N_23473);
or U28956 (N_28956,N_19815,N_20014);
xor U28957 (N_28957,N_21873,N_19323);
or U28958 (N_28958,N_23522,N_18524);
xnor U28959 (N_28959,N_19289,N_22120);
xor U28960 (N_28960,N_20215,N_18113);
xnor U28961 (N_28961,N_19747,N_20610);
xnor U28962 (N_28962,N_21261,N_19654);
or U28963 (N_28963,N_18502,N_23382);
and U28964 (N_28964,N_23387,N_22762);
or U28965 (N_28965,N_22641,N_22735);
or U28966 (N_28966,N_19550,N_21577);
and U28967 (N_28967,N_19963,N_20136);
nand U28968 (N_28968,N_21390,N_18125);
xor U28969 (N_28969,N_22405,N_20955);
and U28970 (N_28970,N_20233,N_20253);
or U28971 (N_28971,N_18872,N_19341);
and U28972 (N_28972,N_20499,N_19388);
xor U28973 (N_28973,N_23615,N_18573);
xor U28974 (N_28974,N_21826,N_21754);
xnor U28975 (N_28975,N_19894,N_19351);
or U28976 (N_28976,N_22141,N_18081);
xnor U28977 (N_28977,N_23195,N_18134);
nand U28978 (N_28978,N_21521,N_21219);
and U28979 (N_28979,N_18406,N_22753);
nand U28980 (N_28980,N_21770,N_21894);
nor U28981 (N_28981,N_19754,N_23155);
and U28982 (N_28982,N_18329,N_20991);
and U28983 (N_28983,N_19634,N_22165);
nor U28984 (N_28984,N_20287,N_18671);
nand U28985 (N_28985,N_22937,N_19960);
or U28986 (N_28986,N_20073,N_19573);
xor U28987 (N_28987,N_23880,N_22371);
or U28988 (N_28988,N_19693,N_23800);
xor U28989 (N_28989,N_19481,N_18503);
xnor U28990 (N_28990,N_20047,N_21658);
nor U28991 (N_28991,N_21709,N_21127);
xnor U28992 (N_28992,N_18115,N_22916);
xor U28993 (N_28993,N_23886,N_18587);
nor U28994 (N_28994,N_20620,N_19803);
nand U28995 (N_28995,N_19026,N_21699);
or U28996 (N_28996,N_20331,N_23867);
nand U28997 (N_28997,N_21835,N_22353);
or U28998 (N_28998,N_20706,N_19121);
or U28999 (N_28999,N_22823,N_18110);
xor U29000 (N_29000,N_23695,N_20551);
and U29001 (N_29001,N_20511,N_19819);
nor U29002 (N_29002,N_22376,N_21892);
xnor U29003 (N_29003,N_23840,N_20907);
nand U29004 (N_29004,N_22685,N_21089);
and U29005 (N_29005,N_18342,N_23185);
and U29006 (N_29006,N_22823,N_20106);
xnor U29007 (N_29007,N_20111,N_20789);
and U29008 (N_29008,N_21552,N_18102);
xnor U29009 (N_29009,N_21334,N_23874);
xor U29010 (N_29010,N_23373,N_22053);
nand U29011 (N_29011,N_18097,N_20137);
or U29012 (N_29012,N_20498,N_20787);
nor U29013 (N_29013,N_19773,N_22629);
nand U29014 (N_29014,N_18879,N_19045);
and U29015 (N_29015,N_20823,N_19956);
xnor U29016 (N_29016,N_22002,N_21125);
or U29017 (N_29017,N_21350,N_21757);
nand U29018 (N_29018,N_18675,N_18582);
xor U29019 (N_29019,N_18150,N_21409);
and U29020 (N_29020,N_23233,N_19669);
nand U29021 (N_29021,N_20647,N_20584);
nand U29022 (N_29022,N_23901,N_21534);
nand U29023 (N_29023,N_20144,N_18492);
nand U29024 (N_29024,N_22412,N_22163);
or U29025 (N_29025,N_23506,N_20615);
or U29026 (N_29026,N_21210,N_23924);
nor U29027 (N_29027,N_22556,N_20905);
or U29028 (N_29028,N_20518,N_21061);
and U29029 (N_29029,N_23221,N_19157);
xor U29030 (N_29030,N_22139,N_22737);
nor U29031 (N_29031,N_22919,N_18024);
nand U29032 (N_29032,N_23809,N_20592);
nand U29033 (N_29033,N_18730,N_20451);
and U29034 (N_29034,N_23015,N_23573);
xor U29035 (N_29035,N_19232,N_21127);
and U29036 (N_29036,N_22616,N_21724);
xnor U29037 (N_29037,N_23966,N_21140);
or U29038 (N_29038,N_21250,N_22534);
xor U29039 (N_29039,N_20010,N_23192);
xor U29040 (N_29040,N_22835,N_19562);
and U29041 (N_29041,N_22666,N_23605);
nand U29042 (N_29042,N_22026,N_21813);
or U29043 (N_29043,N_23535,N_21950);
and U29044 (N_29044,N_21975,N_20366);
nor U29045 (N_29045,N_18456,N_19080);
and U29046 (N_29046,N_19775,N_18867);
nand U29047 (N_29047,N_18010,N_19186);
nor U29048 (N_29048,N_19480,N_20924);
or U29049 (N_29049,N_20719,N_23612);
nand U29050 (N_29050,N_18889,N_20991);
xor U29051 (N_29051,N_20247,N_22390);
nor U29052 (N_29052,N_20109,N_21791);
and U29053 (N_29053,N_18302,N_23258);
nor U29054 (N_29054,N_19880,N_18508);
or U29055 (N_29055,N_21501,N_20080);
xnor U29056 (N_29056,N_21597,N_19924);
nor U29057 (N_29057,N_23107,N_21850);
or U29058 (N_29058,N_21293,N_23452);
and U29059 (N_29059,N_18497,N_18653);
or U29060 (N_29060,N_20689,N_21077);
nand U29061 (N_29061,N_19864,N_22186);
or U29062 (N_29062,N_22818,N_18258);
xor U29063 (N_29063,N_20564,N_20304);
and U29064 (N_29064,N_21484,N_19398);
xor U29065 (N_29065,N_23851,N_21014);
and U29066 (N_29066,N_19976,N_18913);
or U29067 (N_29067,N_23048,N_20430);
and U29068 (N_29068,N_21460,N_18444);
or U29069 (N_29069,N_20447,N_18804);
and U29070 (N_29070,N_18235,N_22217);
and U29071 (N_29071,N_22110,N_18126);
or U29072 (N_29072,N_23170,N_18183);
and U29073 (N_29073,N_18276,N_19093);
and U29074 (N_29074,N_22922,N_23835);
nand U29075 (N_29075,N_22307,N_22871);
xnor U29076 (N_29076,N_20791,N_21540);
or U29077 (N_29077,N_19010,N_19288);
or U29078 (N_29078,N_23881,N_19194);
nand U29079 (N_29079,N_20870,N_23221);
nor U29080 (N_29080,N_22499,N_18761);
nor U29081 (N_29081,N_19046,N_22109);
xnor U29082 (N_29082,N_23011,N_23876);
nor U29083 (N_29083,N_20486,N_18594);
nor U29084 (N_29084,N_21415,N_20168);
xnor U29085 (N_29085,N_23937,N_20154);
and U29086 (N_29086,N_23385,N_19087);
or U29087 (N_29087,N_22851,N_20818);
nand U29088 (N_29088,N_23139,N_22875);
and U29089 (N_29089,N_19145,N_23538);
nand U29090 (N_29090,N_22866,N_21420);
and U29091 (N_29091,N_19252,N_18547);
and U29092 (N_29092,N_22918,N_22657);
or U29093 (N_29093,N_22882,N_21454);
nand U29094 (N_29094,N_20314,N_23500);
nor U29095 (N_29095,N_23111,N_18435);
and U29096 (N_29096,N_21474,N_21395);
nand U29097 (N_29097,N_20351,N_21907);
nand U29098 (N_29098,N_19026,N_22905);
nor U29099 (N_29099,N_23903,N_19605);
xnor U29100 (N_29100,N_18097,N_18897);
nand U29101 (N_29101,N_21290,N_21607);
or U29102 (N_29102,N_21546,N_21048);
xnor U29103 (N_29103,N_18712,N_19328);
and U29104 (N_29104,N_23614,N_23599);
xor U29105 (N_29105,N_23671,N_19653);
nand U29106 (N_29106,N_23675,N_18628);
xor U29107 (N_29107,N_23911,N_20562);
nand U29108 (N_29108,N_21059,N_21805);
nor U29109 (N_29109,N_19316,N_23330);
nand U29110 (N_29110,N_22556,N_22207);
and U29111 (N_29111,N_18235,N_23416);
and U29112 (N_29112,N_19227,N_22327);
nor U29113 (N_29113,N_18859,N_23929);
and U29114 (N_29114,N_22429,N_18753);
or U29115 (N_29115,N_18284,N_21815);
nand U29116 (N_29116,N_19106,N_22154);
and U29117 (N_29117,N_19588,N_20310);
or U29118 (N_29118,N_19034,N_20202);
nor U29119 (N_29119,N_21072,N_21489);
and U29120 (N_29120,N_21628,N_18871);
or U29121 (N_29121,N_23861,N_19666);
and U29122 (N_29122,N_23889,N_23576);
or U29123 (N_29123,N_21664,N_19684);
xor U29124 (N_29124,N_22715,N_19928);
xor U29125 (N_29125,N_19638,N_22651);
or U29126 (N_29126,N_23782,N_23256);
or U29127 (N_29127,N_20238,N_23620);
nor U29128 (N_29128,N_22696,N_19091);
nor U29129 (N_29129,N_23871,N_23690);
or U29130 (N_29130,N_18895,N_23053);
nor U29131 (N_29131,N_20819,N_18047);
xor U29132 (N_29132,N_19277,N_23456);
or U29133 (N_29133,N_18935,N_21052);
nor U29134 (N_29134,N_23698,N_18145);
nand U29135 (N_29135,N_21472,N_21869);
nor U29136 (N_29136,N_23740,N_19268);
or U29137 (N_29137,N_22484,N_22480);
nand U29138 (N_29138,N_19667,N_22800);
or U29139 (N_29139,N_20993,N_18726);
or U29140 (N_29140,N_18191,N_18505);
nor U29141 (N_29141,N_22427,N_18121);
or U29142 (N_29142,N_21379,N_20896);
nor U29143 (N_29143,N_21346,N_18610);
xor U29144 (N_29144,N_21765,N_18744);
xor U29145 (N_29145,N_20865,N_19728);
or U29146 (N_29146,N_22892,N_18542);
or U29147 (N_29147,N_19624,N_23871);
xor U29148 (N_29148,N_22242,N_20056);
xnor U29149 (N_29149,N_18689,N_19488);
nor U29150 (N_29150,N_21508,N_19270);
or U29151 (N_29151,N_23572,N_22630);
or U29152 (N_29152,N_20350,N_19378);
or U29153 (N_29153,N_19845,N_22827);
nand U29154 (N_29154,N_23086,N_22470);
xnor U29155 (N_29155,N_18252,N_23722);
nor U29156 (N_29156,N_20876,N_21432);
and U29157 (N_29157,N_19947,N_22692);
nand U29158 (N_29158,N_23939,N_19302);
and U29159 (N_29159,N_22104,N_21000);
nor U29160 (N_29160,N_23188,N_23469);
and U29161 (N_29161,N_23443,N_18804);
and U29162 (N_29162,N_23908,N_21912);
nor U29163 (N_29163,N_18484,N_21137);
xor U29164 (N_29164,N_18522,N_19201);
xor U29165 (N_29165,N_21562,N_23000);
nor U29166 (N_29166,N_23238,N_20306);
and U29167 (N_29167,N_23316,N_22665);
nor U29168 (N_29168,N_20810,N_22124);
xor U29169 (N_29169,N_21440,N_18256);
xor U29170 (N_29170,N_19588,N_21583);
xor U29171 (N_29171,N_22888,N_19603);
xor U29172 (N_29172,N_19428,N_21475);
or U29173 (N_29173,N_19614,N_23750);
or U29174 (N_29174,N_19146,N_18231);
or U29175 (N_29175,N_19340,N_18242);
nand U29176 (N_29176,N_19344,N_21489);
nor U29177 (N_29177,N_22713,N_21199);
nor U29178 (N_29178,N_18522,N_22721);
or U29179 (N_29179,N_19835,N_20944);
nor U29180 (N_29180,N_21784,N_18617);
nor U29181 (N_29181,N_18575,N_23883);
nor U29182 (N_29182,N_21544,N_18654);
and U29183 (N_29183,N_22641,N_18718);
nor U29184 (N_29184,N_20654,N_20039);
nor U29185 (N_29185,N_23003,N_20659);
and U29186 (N_29186,N_23139,N_23692);
and U29187 (N_29187,N_18768,N_23320);
nor U29188 (N_29188,N_23646,N_23407);
and U29189 (N_29189,N_23753,N_21560);
nand U29190 (N_29190,N_23414,N_19192);
xor U29191 (N_29191,N_21083,N_19107);
and U29192 (N_29192,N_18594,N_20054);
nand U29193 (N_29193,N_19479,N_19617);
or U29194 (N_29194,N_19919,N_20339);
and U29195 (N_29195,N_20300,N_23488);
xnor U29196 (N_29196,N_22088,N_19889);
and U29197 (N_29197,N_19148,N_20959);
nand U29198 (N_29198,N_22419,N_20079);
nand U29199 (N_29199,N_23940,N_19338);
and U29200 (N_29200,N_23808,N_22265);
and U29201 (N_29201,N_19397,N_22058);
and U29202 (N_29202,N_20294,N_21501);
nand U29203 (N_29203,N_19010,N_19715);
nor U29204 (N_29204,N_23795,N_20141);
nor U29205 (N_29205,N_19353,N_21531);
or U29206 (N_29206,N_20956,N_20002);
nand U29207 (N_29207,N_18725,N_22217);
or U29208 (N_29208,N_23237,N_19615);
xnor U29209 (N_29209,N_23063,N_20166);
nand U29210 (N_29210,N_21921,N_20145);
xor U29211 (N_29211,N_22443,N_18848);
nand U29212 (N_29212,N_21060,N_22896);
nor U29213 (N_29213,N_22776,N_22535);
xnor U29214 (N_29214,N_20781,N_18863);
nand U29215 (N_29215,N_21497,N_18990);
nand U29216 (N_29216,N_19417,N_19203);
nor U29217 (N_29217,N_21187,N_19779);
xnor U29218 (N_29218,N_22053,N_22308);
nand U29219 (N_29219,N_18399,N_23642);
or U29220 (N_29220,N_21334,N_21001);
xnor U29221 (N_29221,N_18185,N_21356);
nand U29222 (N_29222,N_19672,N_19948);
nor U29223 (N_29223,N_22524,N_21246);
nand U29224 (N_29224,N_19290,N_23970);
nor U29225 (N_29225,N_22601,N_19441);
or U29226 (N_29226,N_18474,N_19320);
nor U29227 (N_29227,N_20072,N_21953);
and U29228 (N_29228,N_22250,N_20921);
xor U29229 (N_29229,N_23725,N_20774);
or U29230 (N_29230,N_21084,N_22661);
and U29231 (N_29231,N_21309,N_22178);
and U29232 (N_29232,N_18602,N_18383);
nor U29233 (N_29233,N_19210,N_23339);
xor U29234 (N_29234,N_20297,N_22228);
or U29235 (N_29235,N_19504,N_19608);
nor U29236 (N_29236,N_21063,N_19914);
xor U29237 (N_29237,N_23948,N_20188);
nand U29238 (N_29238,N_20578,N_21097);
nor U29239 (N_29239,N_19230,N_18136);
nor U29240 (N_29240,N_20391,N_23378);
nand U29241 (N_29241,N_18810,N_20351);
xor U29242 (N_29242,N_22202,N_23686);
and U29243 (N_29243,N_19701,N_19077);
and U29244 (N_29244,N_19969,N_21158);
or U29245 (N_29245,N_19475,N_20001);
or U29246 (N_29246,N_21103,N_22318);
nor U29247 (N_29247,N_23402,N_21929);
xor U29248 (N_29248,N_20926,N_18954);
xor U29249 (N_29249,N_18383,N_18055);
and U29250 (N_29250,N_23409,N_19711);
nor U29251 (N_29251,N_21949,N_20306);
or U29252 (N_29252,N_23131,N_23053);
nand U29253 (N_29253,N_18101,N_21595);
or U29254 (N_29254,N_22456,N_20548);
nand U29255 (N_29255,N_19418,N_18714);
or U29256 (N_29256,N_22396,N_20802);
and U29257 (N_29257,N_19310,N_21570);
nand U29258 (N_29258,N_22296,N_23609);
nor U29259 (N_29259,N_18690,N_23779);
nand U29260 (N_29260,N_21158,N_18155);
and U29261 (N_29261,N_23419,N_18369);
nand U29262 (N_29262,N_20297,N_18134);
xor U29263 (N_29263,N_21113,N_19195);
and U29264 (N_29264,N_21957,N_22883);
nor U29265 (N_29265,N_22575,N_23558);
or U29266 (N_29266,N_19195,N_21030);
and U29267 (N_29267,N_20114,N_23802);
xnor U29268 (N_29268,N_21460,N_23435);
nor U29269 (N_29269,N_18041,N_20098);
or U29270 (N_29270,N_21859,N_19378);
or U29271 (N_29271,N_23560,N_23269);
xnor U29272 (N_29272,N_23039,N_20373);
nor U29273 (N_29273,N_23837,N_20871);
nand U29274 (N_29274,N_18248,N_23201);
or U29275 (N_29275,N_20483,N_20265);
and U29276 (N_29276,N_18812,N_19186);
xnor U29277 (N_29277,N_20197,N_18026);
or U29278 (N_29278,N_20536,N_19976);
xor U29279 (N_29279,N_19113,N_22249);
and U29280 (N_29280,N_23163,N_23386);
and U29281 (N_29281,N_20947,N_22221);
or U29282 (N_29282,N_20493,N_20948);
xor U29283 (N_29283,N_19889,N_22892);
and U29284 (N_29284,N_19139,N_23695);
nor U29285 (N_29285,N_19657,N_19793);
nor U29286 (N_29286,N_23596,N_20063);
nand U29287 (N_29287,N_21355,N_18152);
and U29288 (N_29288,N_18407,N_21325);
nor U29289 (N_29289,N_20826,N_23254);
nor U29290 (N_29290,N_20123,N_18697);
nand U29291 (N_29291,N_20024,N_21236);
and U29292 (N_29292,N_22745,N_20379);
or U29293 (N_29293,N_18946,N_18537);
or U29294 (N_29294,N_22127,N_20524);
xor U29295 (N_29295,N_19194,N_20557);
and U29296 (N_29296,N_19965,N_21719);
xnor U29297 (N_29297,N_23372,N_18761);
nand U29298 (N_29298,N_18660,N_21916);
xor U29299 (N_29299,N_22929,N_21567);
and U29300 (N_29300,N_20274,N_21966);
nand U29301 (N_29301,N_22005,N_22010);
xor U29302 (N_29302,N_22200,N_21577);
nand U29303 (N_29303,N_21283,N_18886);
and U29304 (N_29304,N_22508,N_22760);
or U29305 (N_29305,N_18711,N_22451);
nand U29306 (N_29306,N_18413,N_20364);
xor U29307 (N_29307,N_22923,N_21054);
nand U29308 (N_29308,N_19691,N_20974);
or U29309 (N_29309,N_23297,N_23022);
nand U29310 (N_29310,N_18470,N_22019);
nand U29311 (N_29311,N_22428,N_22975);
nor U29312 (N_29312,N_22715,N_21494);
nor U29313 (N_29313,N_21988,N_19661);
or U29314 (N_29314,N_23429,N_19269);
xnor U29315 (N_29315,N_22197,N_19071);
nor U29316 (N_29316,N_18036,N_23500);
and U29317 (N_29317,N_19195,N_23840);
xnor U29318 (N_29318,N_20030,N_20565);
nand U29319 (N_29319,N_18283,N_19953);
and U29320 (N_29320,N_21045,N_19694);
xor U29321 (N_29321,N_23312,N_20871);
nand U29322 (N_29322,N_21613,N_18026);
xor U29323 (N_29323,N_22134,N_20316);
nor U29324 (N_29324,N_18220,N_22637);
nand U29325 (N_29325,N_21770,N_18461);
or U29326 (N_29326,N_21012,N_19780);
and U29327 (N_29327,N_23972,N_21953);
or U29328 (N_29328,N_21164,N_20407);
nand U29329 (N_29329,N_20767,N_19012);
and U29330 (N_29330,N_21136,N_19947);
xor U29331 (N_29331,N_18772,N_21260);
nor U29332 (N_29332,N_22971,N_18609);
nor U29333 (N_29333,N_23921,N_22555);
nand U29334 (N_29334,N_20091,N_22900);
and U29335 (N_29335,N_21834,N_23779);
or U29336 (N_29336,N_21769,N_23288);
xnor U29337 (N_29337,N_19013,N_18307);
xor U29338 (N_29338,N_18236,N_22097);
nand U29339 (N_29339,N_18277,N_22206);
nand U29340 (N_29340,N_21669,N_19215);
nand U29341 (N_29341,N_21700,N_21424);
and U29342 (N_29342,N_22769,N_19430);
xnor U29343 (N_29343,N_19701,N_23570);
xnor U29344 (N_29344,N_22906,N_20108);
and U29345 (N_29345,N_22648,N_22575);
nand U29346 (N_29346,N_20874,N_23615);
or U29347 (N_29347,N_20765,N_20369);
nor U29348 (N_29348,N_21023,N_23219);
xnor U29349 (N_29349,N_19184,N_19215);
nand U29350 (N_29350,N_21743,N_18204);
nor U29351 (N_29351,N_22390,N_18514);
xnor U29352 (N_29352,N_21761,N_20350);
nor U29353 (N_29353,N_18856,N_19273);
nor U29354 (N_29354,N_23396,N_22792);
xor U29355 (N_29355,N_23610,N_20417);
nor U29356 (N_29356,N_23283,N_18029);
and U29357 (N_29357,N_22693,N_21929);
nand U29358 (N_29358,N_19527,N_23773);
and U29359 (N_29359,N_21563,N_21881);
or U29360 (N_29360,N_22689,N_18379);
nand U29361 (N_29361,N_18964,N_18096);
nand U29362 (N_29362,N_21635,N_19378);
nand U29363 (N_29363,N_20194,N_21652);
nand U29364 (N_29364,N_20707,N_18626);
and U29365 (N_29365,N_18309,N_21630);
nor U29366 (N_29366,N_22906,N_20827);
nand U29367 (N_29367,N_19133,N_20360);
or U29368 (N_29368,N_19610,N_20593);
xor U29369 (N_29369,N_18334,N_19493);
and U29370 (N_29370,N_20636,N_20252);
and U29371 (N_29371,N_20486,N_23915);
and U29372 (N_29372,N_23907,N_18691);
and U29373 (N_29373,N_23027,N_20920);
xor U29374 (N_29374,N_20098,N_21789);
and U29375 (N_29375,N_21091,N_23422);
and U29376 (N_29376,N_22126,N_19451);
nor U29377 (N_29377,N_19502,N_19614);
and U29378 (N_29378,N_22995,N_21300);
nand U29379 (N_29379,N_20537,N_20136);
nor U29380 (N_29380,N_22998,N_22966);
or U29381 (N_29381,N_21956,N_18739);
and U29382 (N_29382,N_19596,N_22547);
nand U29383 (N_29383,N_20703,N_19588);
or U29384 (N_29384,N_23105,N_18760);
nand U29385 (N_29385,N_23790,N_19953);
xnor U29386 (N_29386,N_22594,N_23978);
or U29387 (N_29387,N_21512,N_22968);
nand U29388 (N_29388,N_23618,N_20834);
and U29389 (N_29389,N_21369,N_23092);
and U29390 (N_29390,N_18973,N_23498);
nor U29391 (N_29391,N_19821,N_18131);
nor U29392 (N_29392,N_18129,N_18838);
and U29393 (N_29393,N_20452,N_19008);
and U29394 (N_29394,N_19999,N_19573);
and U29395 (N_29395,N_20369,N_20600);
and U29396 (N_29396,N_21739,N_21466);
nor U29397 (N_29397,N_23759,N_20330);
or U29398 (N_29398,N_18924,N_23994);
nand U29399 (N_29399,N_18776,N_23717);
nand U29400 (N_29400,N_19889,N_19638);
nand U29401 (N_29401,N_18360,N_23512);
nand U29402 (N_29402,N_18922,N_22912);
xnor U29403 (N_29403,N_20538,N_21287);
nor U29404 (N_29404,N_20854,N_19609);
nor U29405 (N_29405,N_21009,N_19790);
and U29406 (N_29406,N_20024,N_18060);
nor U29407 (N_29407,N_18840,N_23270);
nand U29408 (N_29408,N_20698,N_18792);
nand U29409 (N_29409,N_21960,N_23402);
nand U29410 (N_29410,N_19213,N_19260);
and U29411 (N_29411,N_19168,N_22755);
and U29412 (N_29412,N_18044,N_20051);
xor U29413 (N_29413,N_19296,N_23993);
nand U29414 (N_29414,N_22423,N_21790);
or U29415 (N_29415,N_18686,N_22443);
xnor U29416 (N_29416,N_20008,N_22889);
and U29417 (N_29417,N_22663,N_18798);
or U29418 (N_29418,N_21796,N_21845);
and U29419 (N_29419,N_19326,N_20402);
nand U29420 (N_29420,N_18866,N_22687);
or U29421 (N_29421,N_20940,N_22072);
xnor U29422 (N_29422,N_22292,N_21080);
or U29423 (N_29423,N_22675,N_18330);
nor U29424 (N_29424,N_19175,N_19927);
nand U29425 (N_29425,N_19122,N_23260);
nor U29426 (N_29426,N_21076,N_20729);
xor U29427 (N_29427,N_23771,N_19497);
nand U29428 (N_29428,N_19371,N_18764);
and U29429 (N_29429,N_22722,N_18700);
or U29430 (N_29430,N_23468,N_19017);
xnor U29431 (N_29431,N_23784,N_22512);
or U29432 (N_29432,N_22861,N_23485);
xor U29433 (N_29433,N_22706,N_18020);
nand U29434 (N_29434,N_19957,N_23625);
nor U29435 (N_29435,N_21451,N_19522);
or U29436 (N_29436,N_22788,N_22868);
nor U29437 (N_29437,N_22072,N_19902);
and U29438 (N_29438,N_19190,N_21280);
nand U29439 (N_29439,N_19209,N_23125);
and U29440 (N_29440,N_23738,N_20410);
or U29441 (N_29441,N_22604,N_22081);
nor U29442 (N_29442,N_18246,N_18079);
xor U29443 (N_29443,N_23979,N_19560);
nand U29444 (N_29444,N_23684,N_21319);
xor U29445 (N_29445,N_18683,N_18016);
or U29446 (N_29446,N_19834,N_18816);
and U29447 (N_29447,N_21731,N_23584);
nand U29448 (N_29448,N_20370,N_20859);
nand U29449 (N_29449,N_21956,N_20677);
or U29450 (N_29450,N_21935,N_22961);
or U29451 (N_29451,N_18640,N_23640);
and U29452 (N_29452,N_23356,N_21575);
and U29453 (N_29453,N_23712,N_23750);
and U29454 (N_29454,N_23247,N_20938);
or U29455 (N_29455,N_23195,N_19124);
or U29456 (N_29456,N_20960,N_20348);
nor U29457 (N_29457,N_19451,N_22879);
nand U29458 (N_29458,N_19719,N_23997);
or U29459 (N_29459,N_18276,N_23537);
xor U29460 (N_29460,N_18879,N_22150);
nor U29461 (N_29461,N_18487,N_20507);
nand U29462 (N_29462,N_21909,N_22672);
nand U29463 (N_29463,N_22831,N_22622);
nand U29464 (N_29464,N_18461,N_20852);
nand U29465 (N_29465,N_18361,N_21206);
nor U29466 (N_29466,N_19895,N_21480);
xnor U29467 (N_29467,N_23783,N_22711);
or U29468 (N_29468,N_18554,N_21426);
nand U29469 (N_29469,N_18393,N_18358);
nand U29470 (N_29470,N_20168,N_20176);
xor U29471 (N_29471,N_21371,N_22974);
nand U29472 (N_29472,N_22902,N_21248);
nor U29473 (N_29473,N_18815,N_18706);
nor U29474 (N_29474,N_19186,N_18337);
xnor U29475 (N_29475,N_19137,N_22628);
xor U29476 (N_29476,N_20190,N_23298);
nor U29477 (N_29477,N_21853,N_18891);
and U29478 (N_29478,N_20674,N_18017);
nand U29479 (N_29479,N_23903,N_21867);
and U29480 (N_29480,N_22105,N_19265);
xnor U29481 (N_29481,N_22002,N_20605);
and U29482 (N_29482,N_19592,N_22262);
and U29483 (N_29483,N_18041,N_23465);
or U29484 (N_29484,N_23441,N_22069);
nand U29485 (N_29485,N_19771,N_19335);
nor U29486 (N_29486,N_22225,N_20635);
nor U29487 (N_29487,N_19595,N_21387);
or U29488 (N_29488,N_18757,N_21467);
xor U29489 (N_29489,N_21305,N_23227);
xor U29490 (N_29490,N_21084,N_21589);
and U29491 (N_29491,N_23235,N_19294);
nor U29492 (N_29492,N_23759,N_19894);
nor U29493 (N_29493,N_23389,N_23184);
and U29494 (N_29494,N_22323,N_20665);
nor U29495 (N_29495,N_19696,N_22117);
and U29496 (N_29496,N_18525,N_19240);
nand U29497 (N_29497,N_18823,N_23423);
nand U29498 (N_29498,N_22662,N_22359);
nor U29499 (N_29499,N_19521,N_22325);
or U29500 (N_29500,N_19157,N_23431);
and U29501 (N_29501,N_20121,N_19849);
xnor U29502 (N_29502,N_22452,N_18671);
and U29503 (N_29503,N_21428,N_21630);
or U29504 (N_29504,N_23701,N_20880);
xnor U29505 (N_29505,N_21787,N_21935);
and U29506 (N_29506,N_18855,N_23565);
and U29507 (N_29507,N_22115,N_19315);
nand U29508 (N_29508,N_18339,N_18737);
nand U29509 (N_29509,N_18198,N_21655);
or U29510 (N_29510,N_18393,N_18478);
and U29511 (N_29511,N_21163,N_18050);
and U29512 (N_29512,N_23964,N_20836);
nand U29513 (N_29513,N_20556,N_23388);
xor U29514 (N_29514,N_19596,N_22992);
nor U29515 (N_29515,N_22425,N_20169);
nand U29516 (N_29516,N_23627,N_19284);
xor U29517 (N_29517,N_21575,N_22597);
xor U29518 (N_29518,N_18103,N_21640);
nor U29519 (N_29519,N_20483,N_20988);
or U29520 (N_29520,N_22643,N_19168);
nand U29521 (N_29521,N_21279,N_23091);
nor U29522 (N_29522,N_21547,N_20200);
nand U29523 (N_29523,N_19282,N_20554);
xor U29524 (N_29524,N_22860,N_18924);
or U29525 (N_29525,N_20192,N_18418);
xor U29526 (N_29526,N_21592,N_21977);
nor U29527 (N_29527,N_22820,N_22331);
and U29528 (N_29528,N_20249,N_22075);
nor U29529 (N_29529,N_23681,N_20452);
xor U29530 (N_29530,N_23586,N_21546);
xor U29531 (N_29531,N_19693,N_18841);
nor U29532 (N_29532,N_21556,N_19372);
and U29533 (N_29533,N_23463,N_22249);
nor U29534 (N_29534,N_23221,N_23228);
nand U29535 (N_29535,N_22313,N_23406);
or U29536 (N_29536,N_21004,N_20077);
nand U29537 (N_29537,N_18645,N_20016);
or U29538 (N_29538,N_21983,N_18933);
xnor U29539 (N_29539,N_18882,N_22497);
or U29540 (N_29540,N_19781,N_21737);
nand U29541 (N_29541,N_23643,N_22318);
and U29542 (N_29542,N_18225,N_23528);
nor U29543 (N_29543,N_23294,N_20412);
xnor U29544 (N_29544,N_23038,N_22668);
nor U29545 (N_29545,N_19002,N_18528);
or U29546 (N_29546,N_22662,N_21473);
and U29547 (N_29547,N_19783,N_20001);
nand U29548 (N_29548,N_18006,N_20992);
and U29549 (N_29549,N_22832,N_23540);
nand U29550 (N_29550,N_22585,N_22715);
nand U29551 (N_29551,N_22818,N_19911);
nand U29552 (N_29552,N_23596,N_22125);
or U29553 (N_29553,N_21401,N_21236);
nand U29554 (N_29554,N_22585,N_20585);
nand U29555 (N_29555,N_23856,N_19511);
nor U29556 (N_29556,N_21120,N_22114);
nand U29557 (N_29557,N_19942,N_19695);
nor U29558 (N_29558,N_18473,N_22396);
or U29559 (N_29559,N_22083,N_19161);
and U29560 (N_29560,N_23294,N_20480);
and U29561 (N_29561,N_18518,N_23299);
and U29562 (N_29562,N_18133,N_23837);
nor U29563 (N_29563,N_21669,N_19675);
and U29564 (N_29564,N_22514,N_21458);
or U29565 (N_29565,N_18478,N_19451);
xor U29566 (N_29566,N_23173,N_19856);
and U29567 (N_29567,N_22126,N_18019);
xnor U29568 (N_29568,N_23076,N_19121);
xor U29569 (N_29569,N_21173,N_20409);
nand U29570 (N_29570,N_18729,N_18040);
and U29571 (N_29571,N_21490,N_22227);
or U29572 (N_29572,N_19994,N_22072);
or U29573 (N_29573,N_19871,N_21005);
or U29574 (N_29574,N_20956,N_22704);
xnor U29575 (N_29575,N_21415,N_20613);
and U29576 (N_29576,N_23278,N_19917);
nor U29577 (N_29577,N_19925,N_21542);
nand U29578 (N_29578,N_21765,N_23645);
or U29579 (N_29579,N_18218,N_18619);
nand U29580 (N_29580,N_20101,N_20486);
xor U29581 (N_29581,N_18092,N_18099);
or U29582 (N_29582,N_20015,N_23989);
or U29583 (N_29583,N_20094,N_21337);
and U29584 (N_29584,N_21376,N_23830);
xnor U29585 (N_29585,N_19984,N_19609);
and U29586 (N_29586,N_20306,N_20665);
nand U29587 (N_29587,N_19281,N_22100);
nor U29588 (N_29588,N_18029,N_19192);
nor U29589 (N_29589,N_21598,N_22281);
nand U29590 (N_29590,N_20645,N_21252);
or U29591 (N_29591,N_22674,N_23971);
and U29592 (N_29592,N_21505,N_23013);
xor U29593 (N_29593,N_22980,N_21664);
xor U29594 (N_29594,N_23896,N_19313);
nand U29595 (N_29595,N_19826,N_19417);
and U29596 (N_29596,N_20607,N_23687);
nand U29597 (N_29597,N_20448,N_22624);
or U29598 (N_29598,N_20034,N_23486);
nand U29599 (N_29599,N_20257,N_18608);
or U29600 (N_29600,N_23123,N_22164);
or U29601 (N_29601,N_18970,N_20171);
nor U29602 (N_29602,N_19140,N_19179);
nand U29603 (N_29603,N_20922,N_22953);
xor U29604 (N_29604,N_20754,N_21610);
nand U29605 (N_29605,N_23779,N_23978);
and U29606 (N_29606,N_19827,N_19805);
nand U29607 (N_29607,N_22052,N_20760);
nor U29608 (N_29608,N_21488,N_18945);
and U29609 (N_29609,N_18271,N_23326);
and U29610 (N_29610,N_18786,N_20505);
nor U29611 (N_29611,N_23872,N_19467);
xnor U29612 (N_29612,N_18230,N_19235);
or U29613 (N_29613,N_22269,N_23060);
and U29614 (N_29614,N_22792,N_20893);
nor U29615 (N_29615,N_23600,N_23597);
xor U29616 (N_29616,N_20747,N_21974);
nand U29617 (N_29617,N_20246,N_21144);
or U29618 (N_29618,N_22157,N_20461);
and U29619 (N_29619,N_20405,N_18952);
and U29620 (N_29620,N_22258,N_23569);
nand U29621 (N_29621,N_22144,N_20137);
or U29622 (N_29622,N_23056,N_18459);
xnor U29623 (N_29623,N_22626,N_18472);
nand U29624 (N_29624,N_22538,N_23689);
xnor U29625 (N_29625,N_23423,N_22920);
nor U29626 (N_29626,N_21428,N_20438);
or U29627 (N_29627,N_21247,N_22706);
or U29628 (N_29628,N_18938,N_21122);
xor U29629 (N_29629,N_20061,N_23363);
nand U29630 (N_29630,N_20693,N_19577);
nor U29631 (N_29631,N_19644,N_20749);
nor U29632 (N_29632,N_22898,N_19802);
and U29633 (N_29633,N_22222,N_20227);
xor U29634 (N_29634,N_20749,N_18504);
or U29635 (N_29635,N_21539,N_22480);
nor U29636 (N_29636,N_21001,N_23116);
and U29637 (N_29637,N_22958,N_19984);
nand U29638 (N_29638,N_18733,N_18044);
nor U29639 (N_29639,N_21522,N_22145);
or U29640 (N_29640,N_23386,N_21068);
nor U29641 (N_29641,N_22196,N_22580);
xnor U29642 (N_29642,N_20645,N_21785);
xnor U29643 (N_29643,N_20116,N_20677);
nor U29644 (N_29644,N_19092,N_22621);
or U29645 (N_29645,N_19893,N_22828);
nand U29646 (N_29646,N_19307,N_22581);
nor U29647 (N_29647,N_22417,N_21874);
nor U29648 (N_29648,N_20458,N_18079);
nor U29649 (N_29649,N_23768,N_21773);
nand U29650 (N_29650,N_19198,N_23718);
or U29651 (N_29651,N_19186,N_21578);
xor U29652 (N_29652,N_20923,N_22408);
nand U29653 (N_29653,N_18373,N_22652);
or U29654 (N_29654,N_21930,N_19556);
or U29655 (N_29655,N_18602,N_18996);
nand U29656 (N_29656,N_21453,N_22106);
xnor U29657 (N_29657,N_21690,N_22022);
nor U29658 (N_29658,N_23513,N_20931);
nor U29659 (N_29659,N_20363,N_22246);
nor U29660 (N_29660,N_20005,N_23366);
or U29661 (N_29661,N_21758,N_22786);
and U29662 (N_29662,N_20589,N_18124);
nand U29663 (N_29663,N_21508,N_21151);
nand U29664 (N_29664,N_23836,N_19466);
nor U29665 (N_29665,N_18768,N_18408);
nand U29666 (N_29666,N_19803,N_23435);
nor U29667 (N_29667,N_22410,N_18718);
or U29668 (N_29668,N_22714,N_22487);
nand U29669 (N_29669,N_20763,N_23439);
nand U29670 (N_29670,N_23878,N_20768);
xor U29671 (N_29671,N_22424,N_23833);
nor U29672 (N_29672,N_19404,N_21011);
nand U29673 (N_29673,N_19969,N_20152);
and U29674 (N_29674,N_18488,N_20378);
or U29675 (N_29675,N_18098,N_19797);
xnor U29676 (N_29676,N_20289,N_18519);
or U29677 (N_29677,N_22914,N_18895);
nor U29678 (N_29678,N_22549,N_19410);
nand U29679 (N_29679,N_18699,N_20560);
nor U29680 (N_29680,N_19284,N_22203);
xnor U29681 (N_29681,N_22146,N_21197);
nor U29682 (N_29682,N_22690,N_18246);
and U29683 (N_29683,N_21128,N_21950);
nand U29684 (N_29684,N_20062,N_23134);
xor U29685 (N_29685,N_19488,N_23069);
xor U29686 (N_29686,N_19748,N_21679);
nor U29687 (N_29687,N_21548,N_18850);
nand U29688 (N_29688,N_18593,N_19380);
nor U29689 (N_29689,N_21472,N_19316);
xnor U29690 (N_29690,N_23720,N_22849);
and U29691 (N_29691,N_20394,N_18699);
or U29692 (N_29692,N_19755,N_18671);
xor U29693 (N_29693,N_20032,N_19625);
and U29694 (N_29694,N_21843,N_19860);
or U29695 (N_29695,N_19918,N_20659);
nand U29696 (N_29696,N_19884,N_20361);
and U29697 (N_29697,N_20601,N_21036);
or U29698 (N_29698,N_22469,N_20983);
nand U29699 (N_29699,N_23170,N_21346);
and U29700 (N_29700,N_22091,N_21158);
nand U29701 (N_29701,N_23823,N_23888);
nor U29702 (N_29702,N_18683,N_21958);
and U29703 (N_29703,N_19159,N_19507);
nor U29704 (N_29704,N_21099,N_21283);
nor U29705 (N_29705,N_20577,N_21256);
nor U29706 (N_29706,N_18170,N_18637);
nor U29707 (N_29707,N_22009,N_21519);
nand U29708 (N_29708,N_20549,N_22655);
xor U29709 (N_29709,N_23422,N_21319);
xnor U29710 (N_29710,N_18523,N_20910);
nand U29711 (N_29711,N_18633,N_20530);
nor U29712 (N_29712,N_19074,N_20079);
nand U29713 (N_29713,N_21621,N_18916);
nand U29714 (N_29714,N_19195,N_22170);
xor U29715 (N_29715,N_19235,N_21757);
or U29716 (N_29716,N_18899,N_18792);
and U29717 (N_29717,N_23831,N_18581);
nand U29718 (N_29718,N_19283,N_18207);
xnor U29719 (N_29719,N_19451,N_20449);
and U29720 (N_29720,N_23424,N_18570);
xnor U29721 (N_29721,N_19454,N_19290);
xor U29722 (N_29722,N_21698,N_23508);
and U29723 (N_29723,N_18106,N_20210);
nor U29724 (N_29724,N_18916,N_20209);
and U29725 (N_29725,N_22377,N_22258);
and U29726 (N_29726,N_23973,N_20751);
and U29727 (N_29727,N_22938,N_18206);
nand U29728 (N_29728,N_18813,N_19029);
or U29729 (N_29729,N_20992,N_19937);
xnor U29730 (N_29730,N_20227,N_23367);
and U29731 (N_29731,N_21350,N_19950);
nand U29732 (N_29732,N_19462,N_20416);
nor U29733 (N_29733,N_20780,N_23364);
and U29734 (N_29734,N_20177,N_23822);
nand U29735 (N_29735,N_23454,N_18702);
nand U29736 (N_29736,N_21796,N_20613);
xnor U29737 (N_29737,N_18485,N_23394);
and U29738 (N_29738,N_21343,N_21366);
nor U29739 (N_29739,N_21725,N_21317);
and U29740 (N_29740,N_23388,N_18796);
or U29741 (N_29741,N_23347,N_22806);
nor U29742 (N_29742,N_18161,N_21663);
nor U29743 (N_29743,N_21002,N_20243);
xnor U29744 (N_29744,N_20982,N_21115);
nor U29745 (N_29745,N_22750,N_20913);
xnor U29746 (N_29746,N_19140,N_23739);
nand U29747 (N_29747,N_22504,N_21098);
xor U29748 (N_29748,N_21292,N_19911);
nand U29749 (N_29749,N_21102,N_23961);
and U29750 (N_29750,N_20271,N_23794);
nor U29751 (N_29751,N_22620,N_22631);
nand U29752 (N_29752,N_23069,N_21690);
nand U29753 (N_29753,N_21138,N_18535);
and U29754 (N_29754,N_19476,N_19790);
nor U29755 (N_29755,N_22426,N_23595);
nor U29756 (N_29756,N_18715,N_20371);
and U29757 (N_29757,N_19198,N_20103);
xor U29758 (N_29758,N_19300,N_19038);
nand U29759 (N_29759,N_19202,N_19150);
or U29760 (N_29760,N_19490,N_19276);
or U29761 (N_29761,N_18089,N_19335);
nor U29762 (N_29762,N_21003,N_22020);
or U29763 (N_29763,N_23450,N_22711);
or U29764 (N_29764,N_23822,N_22628);
and U29765 (N_29765,N_21447,N_21978);
nand U29766 (N_29766,N_23998,N_19145);
or U29767 (N_29767,N_19073,N_19918);
or U29768 (N_29768,N_20071,N_18163);
nor U29769 (N_29769,N_20522,N_20078);
xor U29770 (N_29770,N_18722,N_18047);
nand U29771 (N_29771,N_23679,N_23402);
and U29772 (N_29772,N_21994,N_22439);
and U29773 (N_29773,N_19741,N_22554);
nor U29774 (N_29774,N_21976,N_18931);
nor U29775 (N_29775,N_22597,N_23125);
xnor U29776 (N_29776,N_18316,N_20485);
xor U29777 (N_29777,N_22392,N_19354);
nand U29778 (N_29778,N_22988,N_22961);
and U29779 (N_29779,N_19257,N_20509);
and U29780 (N_29780,N_19603,N_23134);
and U29781 (N_29781,N_20767,N_19926);
and U29782 (N_29782,N_19317,N_19899);
nor U29783 (N_29783,N_21992,N_23934);
nand U29784 (N_29784,N_22278,N_21809);
xor U29785 (N_29785,N_23805,N_20523);
nor U29786 (N_29786,N_18653,N_23544);
or U29787 (N_29787,N_23582,N_19979);
xnor U29788 (N_29788,N_18472,N_19624);
and U29789 (N_29789,N_19260,N_19329);
or U29790 (N_29790,N_20925,N_22688);
nor U29791 (N_29791,N_20355,N_21477);
or U29792 (N_29792,N_23834,N_22796);
nor U29793 (N_29793,N_18752,N_21715);
nor U29794 (N_29794,N_18348,N_21064);
nand U29795 (N_29795,N_22633,N_19699);
nand U29796 (N_29796,N_23249,N_21093);
nor U29797 (N_29797,N_20411,N_21431);
or U29798 (N_29798,N_23900,N_18993);
or U29799 (N_29799,N_22357,N_19316);
xnor U29800 (N_29800,N_22556,N_18227);
and U29801 (N_29801,N_18594,N_19737);
nor U29802 (N_29802,N_19912,N_18333);
or U29803 (N_29803,N_22092,N_22818);
and U29804 (N_29804,N_22424,N_18724);
nor U29805 (N_29805,N_22993,N_21942);
xor U29806 (N_29806,N_23268,N_21438);
or U29807 (N_29807,N_21623,N_23367);
or U29808 (N_29808,N_21763,N_22803);
nor U29809 (N_29809,N_22352,N_22340);
nand U29810 (N_29810,N_22175,N_20482);
xnor U29811 (N_29811,N_21121,N_20198);
xor U29812 (N_29812,N_20233,N_18590);
or U29813 (N_29813,N_23708,N_21748);
nand U29814 (N_29814,N_20637,N_19553);
xor U29815 (N_29815,N_22808,N_23036);
nand U29816 (N_29816,N_19644,N_23667);
xnor U29817 (N_29817,N_21768,N_22800);
xor U29818 (N_29818,N_23215,N_21175);
or U29819 (N_29819,N_19471,N_20246);
xnor U29820 (N_29820,N_22499,N_21403);
xor U29821 (N_29821,N_21335,N_18601);
nor U29822 (N_29822,N_19443,N_20800);
and U29823 (N_29823,N_21048,N_19902);
nand U29824 (N_29824,N_19160,N_19275);
and U29825 (N_29825,N_20221,N_19361);
or U29826 (N_29826,N_20382,N_20524);
and U29827 (N_29827,N_20854,N_22869);
xnor U29828 (N_29828,N_23433,N_21299);
or U29829 (N_29829,N_20979,N_20348);
nor U29830 (N_29830,N_18613,N_21871);
nand U29831 (N_29831,N_18072,N_22454);
nor U29832 (N_29832,N_19372,N_18898);
xnor U29833 (N_29833,N_19616,N_21362);
or U29834 (N_29834,N_19582,N_20801);
nand U29835 (N_29835,N_22886,N_23939);
and U29836 (N_29836,N_20567,N_22101);
or U29837 (N_29837,N_20897,N_23189);
xor U29838 (N_29838,N_18728,N_18552);
nor U29839 (N_29839,N_19751,N_22762);
xor U29840 (N_29840,N_18916,N_20082);
nor U29841 (N_29841,N_19804,N_22499);
nor U29842 (N_29842,N_20989,N_23384);
nor U29843 (N_29843,N_21500,N_21255);
nor U29844 (N_29844,N_20719,N_19701);
nor U29845 (N_29845,N_20721,N_22476);
and U29846 (N_29846,N_23528,N_22435);
nand U29847 (N_29847,N_22492,N_21755);
and U29848 (N_29848,N_20384,N_23571);
nand U29849 (N_29849,N_22455,N_23515);
or U29850 (N_29850,N_19887,N_23649);
xnor U29851 (N_29851,N_20425,N_21388);
nor U29852 (N_29852,N_20762,N_22113);
xor U29853 (N_29853,N_21722,N_18710);
nand U29854 (N_29854,N_19201,N_18509);
xnor U29855 (N_29855,N_23377,N_22370);
xnor U29856 (N_29856,N_22964,N_22240);
or U29857 (N_29857,N_18309,N_21095);
and U29858 (N_29858,N_23265,N_20010);
xor U29859 (N_29859,N_22561,N_20681);
and U29860 (N_29860,N_21846,N_23974);
xnor U29861 (N_29861,N_20108,N_22304);
or U29862 (N_29862,N_18933,N_19095);
nand U29863 (N_29863,N_21021,N_23241);
and U29864 (N_29864,N_22541,N_19196);
or U29865 (N_29865,N_19850,N_18317);
nor U29866 (N_29866,N_20295,N_18246);
xnor U29867 (N_29867,N_23482,N_20341);
xor U29868 (N_29868,N_22667,N_19937);
nor U29869 (N_29869,N_23890,N_21738);
and U29870 (N_29870,N_22759,N_18842);
nor U29871 (N_29871,N_22733,N_20143);
and U29872 (N_29872,N_21724,N_23432);
xnor U29873 (N_29873,N_20205,N_19766);
or U29874 (N_29874,N_21219,N_18400);
and U29875 (N_29875,N_18687,N_21969);
and U29876 (N_29876,N_18219,N_21141);
and U29877 (N_29877,N_19957,N_20699);
xnor U29878 (N_29878,N_20105,N_21568);
xnor U29879 (N_29879,N_22294,N_23953);
nand U29880 (N_29880,N_21257,N_19223);
nand U29881 (N_29881,N_19250,N_21846);
nor U29882 (N_29882,N_22009,N_21377);
and U29883 (N_29883,N_18504,N_22912);
nand U29884 (N_29884,N_22726,N_22469);
nor U29885 (N_29885,N_21072,N_19391);
nand U29886 (N_29886,N_23444,N_21433);
nand U29887 (N_29887,N_21424,N_21678);
or U29888 (N_29888,N_23224,N_21307);
nor U29889 (N_29889,N_18925,N_18080);
xor U29890 (N_29890,N_23010,N_20596);
nor U29891 (N_29891,N_20113,N_18528);
or U29892 (N_29892,N_20054,N_18036);
xnor U29893 (N_29893,N_23872,N_19332);
nand U29894 (N_29894,N_23643,N_22645);
xor U29895 (N_29895,N_21061,N_18541);
nor U29896 (N_29896,N_19259,N_19204);
nor U29897 (N_29897,N_21109,N_20865);
or U29898 (N_29898,N_20056,N_18864);
nand U29899 (N_29899,N_19121,N_18191);
and U29900 (N_29900,N_18039,N_21198);
and U29901 (N_29901,N_23100,N_23334);
or U29902 (N_29902,N_23409,N_21029);
xnor U29903 (N_29903,N_18256,N_20890);
nand U29904 (N_29904,N_20313,N_22178);
xor U29905 (N_29905,N_22437,N_23796);
nand U29906 (N_29906,N_23586,N_22324);
xnor U29907 (N_29907,N_23202,N_19237);
or U29908 (N_29908,N_23965,N_20485);
and U29909 (N_29909,N_19455,N_23519);
or U29910 (N_29910,N_19258,N_23797);
xor U29911 (N_29911,N_19472,N_21293);
nor U29912 (N_29912,N_23239,N_18429);
and U29913 (N_29913,N_22055,N_22633);
or U29914 (N_29914,N_21148,N_18709);
nand U29915 (N_29915,N_19232,N_23545);
nand U29916 (N_29916,N_20577,N_23127);
nor U29917 (N_29917,N_20141,N_22462);
xor U29918 (N_29918,N_21799,N_20109);
nand U29919 (N_29919,N_23449,N_23640);
nor U29920 (N_29920,N_21664,N_21300);
or U29921 (N_29921,N_18031,N_21466);
nor U29922 (N_29922,N_20833,N_22505);
or U29923 (N_29923,N_22444,N_23015);
nand U29924 (N_29924,N_18118,N_18473);
or U29925 (N_29925,N_20204,N_18706);
nor U29926 (N_29926,N_22823,N_19089);
xor U29927 (N_29927,N_23757,N_22058);
nor U29928 (N_29928,N_18538,N_20283);
nor U29929 (N_29929,N_18356,N_23968);
and U29930 (N_29930,N_18116,N_19566);
and U29931 (N_29931,N_19142,N_21504);
and U29932 (N_29932,N_23872,N_23749);
xnor U29933 (N_29933,N_23657,N_21149);
or U29934 (N_29934,N_21969,N_23545);
xnor U29935 (N_29935,N_21814,N_18312);
xnor U29936 (N_29936,N_19509,N_22641);
and U29937 (N_29937,N_20188,N_23435);
nor U29938 (N_29938,N_20384,N_22680);
nand U29939 (N_29939,N_19689,N_20091);
or U29940 (N_29940,N_22213,N_21320);
or U29941 (N_29941,N_20245,N_18818);
and U29942 (N_29942,N_22899,N_21831);
nand U29943 (N_29943,N_22981,N_22404);
or U29944 (N_29944,N_19797,N_19366);
nor U29945 (N_29945,N_23606,N_19373);
and U29946 (N_29946,N_19299,N_21845);
nor U29947 (N_29947,N_18332,N_18763);
nand U29948 (N_29948,N_20792,N_20812);
or U29949 (N_29949,N_20692,N_18637);
nor U29950 (N_29950,N_20280,N_19689);
nand U29951 (N_29951,N_20765,N_19959);
xor U29952 (N_29952,N_20529,N_18488);
or U29953 (N_29953,N_18389,N_21342);
or U29954 (N_29954,N_21686,N_20818);
or U29955 (N_29955,N_20326,N_19182);
or U29956 (N_29956,N_22634,N_21558);
xor U29957 (N_29957,N_22566,N_18949);
nand U29958 (N_29958,N_18213,N_23116);
xnor U29959 (N_29959,N_23330,N_18085);
nor U29960 (N_29960,N_21555,N_21530);
nand U29961 (N_29961,N_22207,N_22582);
xor U29962 (N_29962,N_21633,N_19630);
xnor U29963 (N_29963,N_18283,N_20918);
and U29964 (N_29964,N_22528,N_19888);
or U29965 (N_29965,N_18223,N_22388);
or U29966 (N_29966,N_20862,N_20341);
xor U29967 (N_29967,N_20299,N_22499);
and U29968 (N_29968,N_19024,N_23308);
and U29969 (N_29969,N_19832,N_21202);
nor U29970 (N_29970,N_23113,N_21758);
nand U29971 (N_29971,N_18609,N_18244);
nor U29972 (N_29972,N_22227,N_18382);
nor U29973 (N_29973,N_23817,N_19919);
nand U29974 (N_29974,N_22186,N_19857);
xnor U29975 (N_29975,N_21800,N_21661);
nor U29976 (N_29976,N_23520,N_18221);
nor U29977 (N_29977,N_19288,N_18812);
nor U29978 (N_29978,N_19955,N_19982);
xnor U29979 (N_29979,N_23963,N_23668);
and U29980 (N_29980,N_23469,N_22797);
nand U29981 (N_29981,N_18264,N_23118);
xnor U29982 (N_29982,N_23227,N_18264);
and U29983 (N_29983,N_19700,N_19294);
or U29984 (N_29984,N_18689,N_19526);
nor U29985 (N_29985,N_18768,N_22834);
and U29986 (N_29986,N_19312,N_22509);
nor U29987 (N_29987,N_20497,N_21497);
xor U29988 (N_29988,N_23221,N_21284);
or U29989 (N_29989,N_19560,N_19168);
xor U29990 (N_29990,N_22572,N_21750);
and U29991 (N_29991,N_18640,N_20588);
and U29992 (N_29992,N_18346,N_21340);
or U29993 (N_29993,N_22011,N_18411);
xor U29994 (N_29994,N_21895,N_21833);
nand U29995 (N_29995,N_20144,N_19879);
or U29996 (N_29996,N_23597,N_18953);
nor U29997 (N_29997,N_21860,N_19232);
xnor U29998 (N_29998,N_20723,N_18732);
nand U29999 (N_29999,N_19226,N_19502);
nor UO_0 (O_0,N_28189,N_28511);
xnor UO_1 (O_1,N_26331,N_26309);
xor UO_2 (O_2,N_24731,N_26849);
nor UO_3 (O_3,N_24322,N_27853);
and UO_4 (O_4,N_28936,N_27957);
nand UO_5 (O_5,N_28210,N_27109);
and UO_6 (O_6,N_29590,N_27650);
nor UO_7 (O_7,N_24533,N_27653);
and UO_8 (O_8,N_28306,N_25328);
xnor UO_9 (O_9,N_28230,N_26984);
or UO_10 (O_10,N_25107,N_29558);
xnor UO_11 (O_11,N_27523,N_28024);
and UO_12 (O_12,N_26266,N_28538);
xnor UO_13 (O_13,N_27776,N_26550);
xor UO_14 (O_14,N_24430,N_27962);
nand UO_15 (O_15,N_26692,N_25426);
nand UO_16 (O_16,N_29873,N_26977);
xor UO_17 (O_17,N_24146,N_29276);
nand UO_18 (O_18,N_27795,N_27624);
nor UO_19 (O_19,N_29709,N_27455);
and UO_20 (O_20,N_29838,N_26393);
and UO_21 (O_21,N_25142,N_28676);
and UO_22 (O_22,N_25902,N_25489);
or UO_23 (O_23,N_25317,N_28435);
xor UO_24 (O_24,N_28274,N_25100);
nand UO_25 (O_25,N_24741,N_29400);
and UO_26 (O_26,N_26359,N_27718);
and UO_27 (O_27,N_27850,N_24798);
and UO_28 (O_28,N_24452,N_28046);
xor UO_29 (O_29,N_27179,N_28213);
or UO_30 (O_30,N_26219,N_28645);
nor UO_31 (O_31,N_28267,N_26509);
xnor UO_32 (O_32,N_28037,N_27929);
and UO_33 (O_33,N_24383,N_25806);
nand UO_34 (O_34,N_25395,N_25418);
xnor UO_35 (O_35,N_26882,N_27318);
and UO_36 (O_36,N_26942,N_28028);
and UO_37 (O_37,N_25858,N_29275);
or UO_38 (O_38,N_25597,N_24861);
xor UO_39 (O_39,N_29898,N_26188);
and UO_40 (O_40,N_29869,N_29040);
xnor UO_41 (O_41,N_24384,N_29807);
nor UO_42 (O_42,N_27324,N_27841);
and UO_43 (O_43,N_26850,N_29345);
or UO_44 (O_44,N_29199,N_25704);
xor UO_45 (O_45,N_24707,N_24259);
nand UO_46 (O_46,N_29226,N_27497);
and UO_47 (O_47,N_26385,N_28522);
nor UO_48 (O_48,N_29680,N_29739);
or UO_49 (O_49,N_24193,N_28412);
or UO_50 (O_50,N_24370,N_25094);
nor UO_51 (O_51,N_24000,N_24387);
nor UO_52 (O_52,N_27223,N_28455);
nand UO_53 (O_53,N_27117,N_27954);
and UO_54 (O_54,N_26362,N_28808);
and UO_55 (O_55,N_24374,N_27852);
xor UO_56 (O_56,N_26365,N_29190);
nand UO_57 (O_57,N_29086,N_25186);
and UO_58 (O_58,N_24411,N_25177);
nand UO_59 (O_59,N_24382,N_25075);
nor UO_60 (O_60,N_24875,N_27014);
nand UO_61 (O_61,N_25113,N_25706);
nand UO_62 (O_62,N_24845,N_25010);
xor UO_63 (O_63,N_26962,N_28359);
nand UO_64 (O_64,N_26286,N_28007);
or UO_65 (O_65,N_24795,N_26768);
nor UO_66 (O_66,N_28787,N_28151);
or UO_67 (O_67,N_27247,N_27142);
xor UO_68 (O_68,N_28913,N_29631);
nand UO_69 (O_69,N_27439,N_26319);
xor UO_70 (O_70,N_25125,N_24319);
and UO_71 (O_71,N_26391,N_29927);
xor UO_72 (O_72,N_27771,N_28652);
xnor UO_73 (O_73,N_26241,N_29989);
and UO_74 (O_74,N_26538,N_28835);
and UO_75 (O_75,N_24623,N_26593);
nor UO_76 (O_76,N_24584,N_29029);
or UO_77 (O_77,N_25590,N_29586);
or UO_78 (O_78,N_25735,N_27256);
nand UO_79 (O_79,N_26264,N_26552);
nand UO_80 (O_80,N_28017,N_28276);
and UO_81 (O_81,N_25988,N_24443);
nand UO_82 (O_82,N_25568,N_28141);
and UO_83 (O_83,N_27493,N_24982);
and UO_84 (O_84,N_27684,N_25859);
or UO_85 (O_85,N_28277,N_27446);
or UO_86 (O_86,N_28229,N_25141);
xor UO_87 (O_87,N_27531,N_25517);
nand UO_88 (O_88,N_27647,N_25624);
nor UO_89 (O_89,N_28216,N_28138);
nand UO_90 (O_90,N_26196,N_27281);
or UO_91 (O_91,N_27726,N_29777);
nor UO_92 (O_92,N_25534,N_27492);
nand UO_93 (O_93,N_29113,N_29445);
xor UO_94 (O_94,N_24094,N_28330);
and UO_95 (O_95,N_24328,N_28844);
nor UO_96 (O_96,N_25322,N_25938);
or UO_97 (O_97,N_26778,N_24925);
nor UO_98 (O_98,N_24519,N_26789);
xnor UO_99 (O_99,N_28980,N_28252);
and UO_100 (O_100,N_29726,N_25530);
or UO_101 (O_101,N_26719,N_24512);
and UO_102 (O_102,N_29691,N_29103);
or UO_103 (O_103,N_27143,N_27772);
nand UO_104 (O_104,N_28431,N_28419);
or UO_105 (O_105,N_26743,N_24460);
or UO_106 (O_106,N_26721,N_27222);
nor UO_107 (O_107,N_26884,N_26016);
or UO_108 (O_108,N_27111,N_26018);
nand UO_109 (O_109,N_29470,N_25648);
and UO_110 (O_110,N_24780,N_24294);
and UO_111 (O_111,N_26745,N_24763);
or UO_112 (O_112,N_25166,N_26676);
and UO_113 (O_113,N_28422,N_26132);
xnor UO_114 (O_114,N_27894,N_25847);
and UO_115 (O_115,N_28746,N_27000);
nor UO_116 (O_116,N_25430,N_29727);
nand UO_117 (O_117,N_25691,N_26926);
nand UO_118 (O_118,N_28405,N_28908);
nand UO_119 (O_119,N_25156,N_28702);
nor UO_120 (O_120,N_28919,N_26901);
nand UO_121 (O_121,N_26812,N_25413);
or UO_122 (O_122,N_28968,N_29167);
nand UO_123 (O_123,N_27651,N_29170);
nor UO_124 (O_124,N_28701,N_28956);
nor UO_125 (O_125,N_29532,N_28237);
xnor UO_126 (O_126,N_29817,N_28157);
or UO_127 (O_127,N_26049,N_25947);
nor UO_128 (O_128,N_26009,N_25538);
nand UO_129 (O_129,N_29320,N_24231);
xor UO_130 (O_130,N_24848,N_27180);
xor UO_131 (O_131,N_24622,N_29012);
nand UO_132 (O_132,N_24878,N_26269);
nand UO_133 (O_133,N_24559,N_26093);
nor UO_134 (O_134,N_25869,N_29014);
and UO_135 (O_135,N_25888,N_28887);
xor UO_136 (O_136,N_25742,N_25487);
xor UO_137 (O_137,N_26204,N_29616);
and UO_138 (O_138,N_29075,N_27886);
or UO_139 (O_139,N_24232,N_26140);
or UO_140 (O_140,N_25136,N_28019);
nand UO_141 (O_141,N_27182,N_28984);
nor UO_142 (O_142,N_24808,N_24029);
or UO_143 (O_143,N_26860,N_27075);
xnor UO_144 (O_144,N_29592,N_24479);
and UO_145 (O_145,N_27603,N_29706);
xnor UO_146 (O_146,N_26999,N_25975);
xnor UO_147 (O_147,N_29019,N_25604);
nand UO_148 (O_148,N_24826,N_27992);
nor UO_149 (O_149,N_24638,N_28148);
xor UO_150 (O_150,N_26311,N_28199);
or UO_151 (O_151,N_24569,N_26771);
nand UO_152 (O_152,N_25798,N_28211);
xor UO_153 (O_153,N_29372,N_26931);
or UO_154 (O_154,N_29987,N_28386);
nor UO_155 (O_155,N_27635,N_28066);
xor UO_156 (O_156,N_27609,N_26576);
or UO_157 (O_157,N_27203,N_26583);
or UO_158 (O_158,N_27924,N_28944);
or UO_159 (O_159,N_27141,N_27808);
or UO_160 (O_160,N_27269,N_24767);
nand UO_161 (O_161,N_26835,N_29135);
and UO_162 (O_162,N_25054,N_24675);
nor UO_163 (O_163,N_25133,N_25575);
and UO_164 (O_164,N_26810,N_28737);
xor UO_165 (O_165,N_26124,N_25327);
and UO_166 (O_166,N_28651,N_27414);
nor UO_167 (O_167,N_25443,N_24945);
or UO_168 (O_168,N_27326,N_29765);
and UO_169 (O_169,N_28029,N_29951);
xor UO_170 (O_170,N_29603,N_26099);
xor UO_171 (O_171,N_28396,N_28561);
nor UO_172 (O_172,N_25330,N_24132);
nand UO_173 (O_173,N_26031,N_27428);
xnor UO_174 (O_174,N_29172,N_27031);
nor UO_175 (O_175,N_26971,N_27390);
nor UO_176 (O_176,N_28454,N_28299);
nor UO_177 (O_177,N_26557,N_26117);
nor UO_178 (O_178,N_27548,N_28240);
nand UO_179 (O_179,N_27132,N_28067);
nor UO_180 (O_180,N_27791,N_28845);
and UO_181 (O_181,N_24646,N_24613);
nand UO_182 (O_182,N_28715,N_26037);
nor UO_183 (O_183,N_28491,N_28950);
nor UO_184 (O_184,N_27727,N_29140);
or UO_185 (O_185,N_26710,N_27385);
nand UO_186 (O_186,N_27987,N_29801);
and UO_187 (O_187,N_24561,N_29686);
and UO_188 (O_188,N_25268,N_29427);
or UO_189 (O_189,N_24988,N_29208);
nand UO_190 (O_190,N_25868,N_27519);
xnor UO_191 (O_191,N_29665,N_28177);
and UO_192 (O_192,N_27948,N_25215);
and UO_193 (O_193,N_29741,N_29679);
nor UO_194 (O_194,N_25466,N_26527);
nand UO_195 (O_195,N_25082,N_28933);
xnor UO_196 (O_196,N_29529,N_26980);
nand UO_197 (O_197,N_26974,N_24329);
xor UO_198 (O_198,N_24971,N_25004);
or UO_199 (O_199,N_29397,N_24380);
and UO_200 (O_200,N_24190,N_27283);
or UO_201 (O_201,N_25481,N_27836);
or UO_202 (O_202,N_29066,N_24385);
nand UO_203 (O_203,N_25863,N_26862);
nor UO_204 (O_204,N_25615,N_26453);
nand UO_205 (O_205,N_28162,N_26854);
nor UO_206 (O_206,N_25622,N_28384);
nor UO_207 (O_207,N_27129,N_27909);
and UO_208 (O_208,N_25793,N_28893);
nor UO_209 (O_209,N_26225,N_24568);
nand UO_210 (O_210,N_24158,N_28614);
xnor UO_211 (O_211,N_26275,N_24237);
nor UO_212 (O_212,N_26741,N_27242);
nor UO_213 (O_213,N_27865,N_29154);
or UO_214 (O_214,N_24333,N_29521);
xor UO_215 (O_215,N_28214,N_29497);
nor UO_216 (O_216,N_28172,N_29389);
nor UO_217 (O_217,N_29469,N_26905);
nor UO_218 (O_218,N_29522,N_29050);
nor UO_219 (O_219,N_29054,N_27513);
nor UO_220 (O_220,N_29753,N_28878);
or UO_221 (O_221,N_29660,N_28391);
nor UO_222 (O_222,N_24650,N_27566);
xor UO_223 (O_223,N_28127,N_26290);
nand UO_224 (O_224,N_24871,N_27122);
nor UO_225 (O_225,N_28866,N_24467);
nand UO_226 (O_226,N_26685,N_28732);
nand UO_227 (O_227,N_25705,N_28814);
nor UO_228 (O_228,N_27254,N_26891);
nand UO_229 (O_229,N_25972,N_25378);
and UO_230 (O_230,N_29045,N_27757);
xor UO_231 (O_231,N_25626,N_24641);
xnor UO_232 (O_232,N_25598,N_26279);
nor UO_233 (O_233,N_28823,N_24420);
nor UO_234 (O_234,N_29566,N_29303);
nand UO_235 (O_235,N_27309,N_29393);
and UO_236 (O_236,N_29857,N_26799);
and UO_237 (O_237,N_27662,N_25137);
or UO_238 (O_238,N_28343,N_29153);
xor UO_239 (O_239,N_24334,N_28730);
nand UO_240 (O_240,N_27646,N_25594);
nand UO_241 (O_241,N_24176,N_27690);
or UO_242 (O_242,N_26187,N_28855);
or UO_243 (O_243,N_27311,N_28429);
and UO_244 (O_244,N_24455,N_27691);
and UO_245 (O_245,N_25122,N_27748);
xor UO_246 (O_246,N_25767,N_27572);
or UO_247 (O_247,N_29827,N_24046);
nand UO_248 (O_248,N_26082,N_28088);
and UO_249 (O_249,N_25209,N_24700);
or UO_250 (O_250,N_29749,N_27370);
nand UO_251 (O_251,N_24256,N_26821);
xnor UO_252 (O_252,N_26885,N_26915);
nor UO_253 (O_253,N_26511,N_28225);
nand UO_254 (O_254,N_29635,N_28884);
or UO_255 (O_255,N_29772,N_29994);
nor UO_256 (O_256,N_24769,N_25901);
xor UO_257 (O_257,N_28508,N_29419);
and UO_258 (O_258,N_29251,N_29336);
or UO_259 (O_259,N_28310,N_26322);
xor UO_260 (O_260,N_26454,N_24099);
or UO_261 (O_261,N_27939,N_25008);
or UO_262 (O_262,N_27190,N_29923);
xor UO_263 (O_263,N_26804,N_26413);
nand UO_264 (O_264,N_25353,N_28914);
nand UO_265 (O_265,N_26736,N_25762);
and UO_266 (O_266,N_27374,N_27846);
nand UO_267 (O_267,N_26536,N_28659);
or UO_268 (O_268,N_24184,N_27154);
or UO_269 (O_269,N_28336,N_28228);
and UO_270 (O_270,N_24228,N_28793);
xnor UO_271 (O_271,N_28688,N_25173);
xor UO_272 (O_272,N_26801,N_26014);
nor UO_273 (O_273,N_27804,N_28929);
nand UO_274 (O_274,N_27536,N_26932);
xor UO_275 (O_275,N_29877,N_26348);
or UO_276 (O_276,N_27198,N_29974);
nor UO_277 (O_277,N_25049,N_29200);
nor UO_278 (O_278,N_25275,N_25952);
nor UO_279 (O_279,N_26571,N_28314);
nand UO_280 (O_280,N_27859,N_27689);
nand UO_281 (O_281,N_28945,N_29704);
nor UO_282 (O_282,N_26164,N_29152);
and UO_283 (O_283,N_25650,N_24394);
or UO_284 (O_284,N_29234,N_28828);
nor UO_285 (O_285,N_25198,N_24981);
xnor UO_286 (O_286,N_24412,N_29373);
or UO_287 (O_287,N_25830,N_28518);
and UO_288 (O_288,N_27342,N_26904);
or UO_289 (O_289,N_29952,N_24323);
nand UO_290 (O_290,N_29252,N_26062);
xor UO_291 (O_291,N_25323,N_25629);
nand UO_292 (O_292,N_27288,N_25039);
nand UO_293 (O_293,N_26080,N_29804);
or UO_294 (O_294,N_29625,N_29132);
nand UO_295 (O_295,N_24579,N_29241);
nand UO_296 (O_296,N_27972,N_29715);
or UO_297 (O_297,N_26339,N_26486);
xnor UO_298 (O_298,N_27366,N_25372);
nand UO_299 (O_299,N_28084,N_25657);
or UO_300 (O_300,N_28205,N_29426);
and UO_301 (O_301,N_27032,N_24896);
xor UO_302 (O_302,N_27049,N_28588);
nor UO_303 (O_303,N_25121,N_27160);
xnor UO_304 (O_304,N_26462,N_24835);
and UO_305 (O_305,N_26656,N_29614);
xnor UO_306 (O_306,N_24667,N_29297);
xnor UO_307 (O_307,N_26839,N_26913);
or UO_308 (O_308,N_25219,N_25021);
or UO_309 (O_309,N_29598,N_24143);
and UO_310 (O_310,N_24669,N_27863);
or UO_311 (O_311,N_25408,N_25846);
nor UO_312 (O_312,N_29123,N_26770);
xor UO_313 (O_313,N_27789,N_26421);
or UO_314 (O_314,N_29908,N_28865);
and UO_315 (O_315,N_25471,N_25612);
or UO_316 (O_316,N_24162,N_27970);
or UO_317 (O_317,N_24979,N_25060);
and UO_318 (O_318,N_29579,N_26960);
xor UO_319 (O_319,N_26883,N_26034);
nor UO_320 (O_320,N_24955,N_27565);
xor UO_321 (O_321,N_29893,N_27145);
and UO_322 (O_322,N_25526,N_29839);
or UO_323 (O_323,N_29093,N_24003);
or UO_324 (O_324,N_25759,N_26069);
and UO_325 (O_325,N_25843,N_29955);
or UO_326 (O_326,N_28358,N_25791);
or UO_327 (O_327,N_29349,N_29474);
or UO_328 (O_328,N_29279,N_29984);
nor UO_329 (O_329,N_28869,N_24629);
nor UO_330 (O_330,N_26975,N_28879);
nor UO_331 (O_331,N_25770,N_24873);
xnor UO_332 (O_332,N_24106,N_24537);
nor UO_333 (O_333,N_24214,N_25199);
or UO_334 (O_334,N_26243,N_28873);
xor UO_335 (O_335,N_27964,N_25690);
xor UO_336 (O_336,N_25143,N_27762);
nor UO_337 (O_337,N_28639,N_26531);
nand UO_338 (O_338,N_29482,N_26933);
and UO_339 (O_339,N_29022,N_26375);
nand UO_340 (O_340,N_26239,N_29229);
xnor UO_341 (O_341,N_24816,N_29929);
xor UO_342 (O_342,N_25112,N_24014);
nor UO_343 (O_343,N_29876,N_27818);
nand UO_344 (O_344,N_27080,N_26217);
xnor UO_345 (O_345,N_28517,N_27304);
nor UO_346 (O_346,N_26238,N_25250);
nor UO_347 (O_347,N_25725,N_25181);
and UO_348 (O_348,N_28939,N_26730);
or UO_349 (O_349,N_24618,N_25493);
nand UO_350 (O_350,N_24227,N_26227);
or UO_351 (O_351,N_24157,N_25549);
xor UO_352 (O_352,N_25535,N_29095);
xnor UO_353 (O_353,N_28691,N_25973);
nor UO_354 (O_354,N_26496,N_27538);
or UO_355 (O_355,N_26718,N_25776);
and UO_356 (O_356,N_29401,N_29041);
xnor UO_357 (O_357,N_25404,N_28365);
nand UO_358 (O_358,N_29463,N_26892);
nor UO_359 (O_359,N_28812,N_25043);
and UO_360 (O_360,N_28171,N_26325);
nor UO_361 (O_361,N_27549,N_24899);
and UO_362 (O_362,N_28272,N_27889);
nor UO_363 (O_363,N_26463,N_27404);
nand UO_364 (O_364,N_27996,N_25764);
xnor UO_365 (O_365,N_24814,N_28740);
nor UO_366 (O_366,N_25616,N_29479);
nand UO_367 (O_367,N_24092,N_25969);
and UO_368 (O_368,N_27765,N_28013);
or UO_369 (O_369,N_27167,N_26506);
and UO_370 (O_370,N_28091,N_24963);
nor UO_371 (O_371,N_24311,N_24514);
xnor UO_372 (O_372,N_27051,N_26178);
nor UO_373 (O_373,N_28040,N_28125);
or UO_374 (O_374,N_27120,N_27351);
nor UO_375 (O_375,N_29493,N_27403);
nor UO_376 (O_376,N_24822,N_29368);
or UO_377 (O_377,N_27039,N_27206);
or UO_378 (O_378,N_25392,N_29347);
xnor UO_379 (O_379,N_27755,N_29512);
xnor UO_380 (O_380,N_28262,N_25316);
and UO_381 (O_381,N_28313,N_29289);
xnor UO_382 (O_382,N_28729,N_25981);
xor UO_383 (O_383,N_27121,N_26629);
xnor UO_384 (O_384,N_28436,N_28990);
xnor UO_385 (O_385,N_27057,N_29774);
and UO_386 (O_386,N_24350,N_24160);
nand UO_387 (O_387,N_28801,N_26589);
nand UO_388 (O_388,N_26671,N_24859);
or UO_389 (O_389,N_27785,N_28898);
nor UO_390 (O_390,N_29581,N_28521);
nor UO_391 (O_391,N_24119,N_27272);
or UO_392 (O_392,N_27914,N_27583);
xor UO_393 (O_393,N_24892,N_24226);
and UO_394 (O_394,N_26759,N_29162);
or UO_395 (O_395,N_27817,N_26136);
or UO_396 (O_396,N_25723,N_26909);
nand UO_397 (O_397,N_25371,N_26208);
or UO_398 (O_398,N_28749,N_24199);
xnor UO_399 (O_399,N_29037,N_27289);
or UO_400 (O_400,N_29414,N_24564);
xor UO_401 (O_401,N_27613,N_26078);
and UO_402 (O_402,N_24761,N_25633);
nand UO_403 (O_403,N_26212,N_28619);
nand UO_404 (O_404,N_27930,N_25038);
nor UO_405 (O_405,N_26827,N_27163);
nor UO_406 (O_406,N_28383,N_24583);
or UO_407 (O_407,N_26711,N_26223);
nor UO_408 (O_408,N_29312,N_25427);
or UO_409 (O_409,N_27564,N_28051);
and UO_410 (O_410,N_28674,N_27052);
xor UO_411 (O_411,N_29783,N_28724);
xnor UO_412 (O_412,N_28297,N_29658);
nor UO_413 (O_413,N_28161,N_27730);
nor UO_414 (O_414,N_29648,N_26211);
or UO_415 (O_415,N_24931,N_28137);
nor UO_416 (O_416,N_24013,N_28147);
nor UO_417 (O_417,N_28438,N_27333);
nand UO_418 (O_418,N_29624,N_24487);
xnor UO_419 (O_419,N_25174,N_24023);
nor UO_420 (O_420,N_24451,N_26672);
and UO_421 (O_421,N_29295,N_25269);
nor UO_422 (O_422,N_27217,N_25341);
and UO_423 (O_423,N_27831,N_24694);
nand UO_424 (O_424,N_26541,N_27666);
or UO_425 (O_425,N_29387,N_28899);
or UO_426 (O_426,N_27199,N_26379);
or UO_427 (O_427,N_27923,N_28542);
and UO_428 (O_428,N_29773,N_24705);
and UO_429 (O_429,N_24539,N_27656);
nor UO_430 (O_430,N_26220,N_28603);
and UO_431 (O_431,N_25910,N_25029);
nand UO_432 (O_432,N_24096,N_25578);
or UO_433 (O_433,N_25312,N_28257);
nor UO_434 (O_434,N_28408,N_28699);
and UO_435 (O_435,N_26284,N_27926);
nand UO_436 (O_436,N_28209,N_29829);
nor UO_437 (O_437,N_24651,N_27018);
nor UO_438 (O_438,N_28525,N_29144);
nand UO_439 (O_439,N_27316,N_24484);
or UO_440 (O_440,N_25367,N_26865);
xor UO_441 (O_441,N_26395,N_29201);
nor UO_442 (O_442,N_24185,N_27262);
nor UO_443 (O_443,N_26330,N_28757);
and UO_444 (O_444,N_26332,N_26826);
and UO_445 (O_445,N_29067,N_26815);
nand UO_446 (O_446,N_26599,N_28070);
or UO_447 (O_447,N_24266,N_26600);
and UO_448 (O_448,N_29659,N_28905);
or UO_449 (O_449,N_26394,N_29287);
and UO_450 (O_450,N_24781,N_28786);
xor UO_451 (O_451,N_24052,N_26397);
and UO_452 (O_452,N_25571,N_25120);
or UO_453 (O_453,N_24563,N_24867);
nand UO_454 (O_454,N_26387,N_29439);
and UO_455 (O_455,N_24144,N_25479);
or UO_456 (O_456,N_24684,N_24865);
nand UO_457 (O_457,N_27606,N_25914);
or UO_458 (O_458,N_27136,N_27191);
or UO_459 (O_459,N_29429,N_27292);
or UO_460 (O_460,N_27149,N_29713);
or UO_461 (O_461,N_28545,N_28356);
nor UO_462 (O_462,N_25184,N_25270);
nand UO_463 (O_463,N_25354,N_27615);
nand UO_464 (O_464,N_27470,N_29443);
nand UO_465 (O_465,N_28567,N_25904);
xnor UO_466 (O_466,N_29420,N_29607);
nand UO_467 (O_467,N_28541,N_27241);
nand UO_468 (O_468,N_27685,N_25668);
xor UO_469 (O_469,N_29149,N_28414);
or UO_470 (O_470,N_24283,N_24620);
or UO_471 (O_471,N_28316,N_28625);
nor UO_472 (O_472,N_29793,N_27800);
nor UO_473 (O_473,N_28870,N_29990);
and UO_474 (O_474,N_26503,N_25949);
xnor UO_475 (O_475,N_25572,N_26030);
or UO_476 (O_476,N_25515,N_27275);
xor UO_477 (O_477,N_29130,N_26428);
nor UO_478 (O_478,N_24648,N_25452);
or UO_479 (O_479,N_29642,N_26235);
or UO_480 (O_480,N_24267,N_29995);
and UO_481 (O_481,N_25602,N_27979);
nand UO_482 (O_482,N_25216,N_29004);
xnor UO_483 (O_483,N_24125,N_27900);
and UO_484 (O_484,N_27728,N_24853);
xnor UO_485 (O_485,N_27001,N_27516);
nor UO_486 (O_486,N_28081,N_26459);
nand UO_487 (O_487,N_27761,N_26831);
xnor UO_488 (O_488,N_26853,N_24893);
xor UO_489 (O_489,N_26564,N_25414);
or UO_490 (O_490,N_29417,N_24191);
xnor UO_491 (O_491,N_27276,N_29227);
and UO_492 (O_492,N_28820,N_27661);
or UO_493 (O_493,N_24043,N_27530);
nand UO_494 (O_494,N_24765,N_27714);
xor UO_495 (O_495,N_24556,N_27479);
and UO_496 (O_496,N_27174,N_28390);
nor UO_497 (O_497,N_25309,N_26775);
or UO_498 (O_498,N_28174,N_25108);
xor UO_499 (O_499,N_26410,N_29001);
nor UO_500 (O_500,N_27216,N_24759);
and UO_501 (O_501,N_24607,N_25553);
xnor UO_502 (O_502,N_29612,N_25871);
nor UO_503 (O_503,N_27384,N_24168);
or UO_504 (O_504,N_27550,N_25611);
xor UO_505 (O_505,N_26414,N_24885);
xor UO_506 (O_506,N_26064,N_25297);
xnor UO_507 (O_507,N_29517,N_24983);
and UO_508 (O_508,N_25254,N_27193);
and UO_509 (O_509,N_26694,N_28876);
nand UO_510 (O_510,N_26688,N_29385);
nand UO_511 (O_511,N_27591,N_28339);
and UO_512 (O_512,N_26361,N_25772);
xor UO_513 (O_513,N_24140,N_24676);
xnor UO_514 (O_514,N_29997,N_28881);
nand UO_515 (O_515,N_27920,N_24277);
nand UO_516 (O_516,N_27208,N_29794);
or UO_517 (O_517,N_28983,N_26019);
nor UO_518 (O_518,N_25337,N_27412);
nand UO_519 (O_519,N_26824,N_28932);
or UO_520 (O_520,N_24686,N_26007);
xnor UO_521 (O_521,N_28097,N_27810);
or UO_522 (O_522,N_24726,N_25208);
nor UO_523 (O_523,N_26234,N_29525);
nor UO_524 (O_524,N_27074,N_29567);
nor UO_525 (O_525,N_24422,N_27540);
xnor UO_526 (O_526,N_25528,N_29290);
or UO_527 (O_527,N_28641,N_28816);
nor UO_528 (O_528,N_29495,N_26010);
nor UO_529 (O_529,N_26432,N_27864);
or UO_530 (O_530,N_25444,N_24447);
or UO_531 (O_531,N_27007,N_27814);
and UO_532 (O_532,N_27113,N_29830);
nor UO_533 (O_533,N_25324,N_28076);
or UO_534 (O_534,N_29311,N_25787);
nor UO_535 (O_535,N_29457,N_27994);
and UO_536 (O_536,N_27733,N_26720);
nand UO_537 (O_537,N_26300,N_27130);
and UO_538 (O_538,N_24503,N_29545);
or UO_539 (O_539,N_27286,N_24666);
xnor UO_540 (O_540,N_26179,N_26675);
xor UO_541 (O_541,N_26615,N_27745);
xnor UO_542 (O_542,N_29197,N_24950);
and UO_543 (O_543,N_26707,N_28735);
nand UO_544 (O_544,N_28510,N_27310);
or UO_545 (O_545,N_26598,N_25879);
nand UO_546 (O_546,N_27002,N_27619);
or UO_547 (O_547,N_28344,N_25920);
or UO_548 (O_548,N_27360,N_24720);
xnor UO_549 (O_549,N_27004,N_26524);
nand UO_550 (O_550,N_25631,N_28400);
and UO_551 (O_551,N_26859,N_27967);
xnor UO_552 (O_552,N_25700,N_29073);
nand UO_553 (O_553,N_28364,N_25024);
xnor UO_554 (O_554,N_27421,N_24693);
nand UO_555 (O_555,N_29613,N_26798);
nor UO_556 (O_556,N_25243,N_28411);
or UO_557 (O_557,N_28989,N_27192);
or UO_558 (O_558,N_29747,N_29183);
and UO_559 (O_559,N_29724,N_26844);
nor UO_560 (O_560,N_24086,N_26510);
and UO_561 (O_561,N_24944,N_26988);
xor UO_562 (O_562,N_27960,N_25290);
nor UO_563 (O_563,N_27234,N_28345);
nor UO_564 (O_564,N_25503,N_25931);
nor UO_565 (O_565,N_24634,N_25832);
nor UO_566 (O_566,N_28074,N_27503);
xnor UO_567 (O_567,N_29491,N_25609);
or UO_568 (O_568,N_26782,N_26021);
nor UO_569 (O_569,N_28327,N_24949);
nor UO_570 (O_570,N_29173,N_24342);
or UO_571 (O_571,N_27551,N_29632);
xnor UO_572 (O_572,N_29668,N_25228);
xnor UO_573 (O_573,N_25407,N_28481);
nor UO_574 (O_574,N_24524,N_27978);
nor UO_575 (O_575,N_24985,N_25398);
nand UO_576 (O_576,N_25302,N_25823);
or UO_577 (O_577,N_29334,N_24213);
or UO_578 (O_578,N_29106,N_27486);
nor UO_579 (O_579,N_28265,N_26785);
or UO_580 (O_580,N_25662,N_28063);
nand UO_581 (O_581,N_27911,N_25016);
nand UO_582 (O_582,N_29498,N_28264);
nor UO_583 (O_583,N_24482,N_24349);
xnor UO_584 (O_584,N_29575,N_24272);
xnor UO_585 (O_585,N_27759,N_29879);
and UO_586 (O_586,N_24987,N_28813);
and UO_587 (O_587,N_29020,N_26857);
and UO_588 (O_588,N_26426,N_29046);
nor UO_589 (O_589,N_25720,N_29629);
nand UO_590 (O_590,N_24252,N_28058);
nand UO_591 (O_591,N_24991,N_28885);
or UO_592 (O_592,N_24122,N_25329);
xnor UO_593 (O_593,N_28690,N_29175);
and UO_594 (O_594,N_28092,N_29109);
and UO_595 (O_595,N_25099,N_26472);
xnor UO_596 (O_596,N_26106,N_24105);
nand UO_597 (O_597,N_25247,N_24047);
or UO_598 (O_598,N_24485,N_26518);
and UO_599 (O_599,N_28445,N_26402);
and UO_600 (O_600,N_25391,N_28155);
or UO_601 (O_601,N_29578,N_24742);
and UO_602 (O_602,N_26948,N_29761);
or UO_603 (O_603,N_26105,N_25259);
and UO_604 (O_604,N_26923,N_26574);
nand UO_605 (O_605,N_27330,N_27096);
xnor UO_606 (O_606,N_26185,N_29950);
nor UO_607 (O_607,N_25350,N_29714);
xnor UO_608 (O_608,N_28920,N_29652);
nand UO_609 (O_609,N_25647,N_28271);
or UO_610 (O_610,N_29872,N_24254);
and UO_611 (O_611,N_27178,N_29315);
xnor UO_612 (O_612,N_24903,N_25027);
or UO_613 (O_613,N_25676,N_26992);
nand UO_614 (O_614,N_28570,N_26636);
and UO_615 (O_615,N_28890,N_28159);
and UO_616 (O_616,N_25817,N_28082);
or UO_617 (O_617,N_28236,N_24764);
or UO_618 (O_618,N_27392,N_25654);
or UO_619 (O_619,N_24797,N_29961);
and UO_620 (O_620,N_29993,N_29313);
xnor UO_621 (O_621,N_26540,N_24238);
and UO_622 (O_622,N_24296,N_27431);
xor UO_623 (O_623,N_24205,N_26956);
and UO_624 (O_624,N_25393,N_28407);
nor UO_625 (O_625,N_26200,N_26261);
xnor UO_626 (O_626,N_25491,N_29862);
or UO_627 (O_627,N_29245,N_27009);
xor UO_628 (O_628,N_24172,N_26701);
xor UO_629 (O_629,N_26317,N_29802);
and UO_630 (O_630,N_24643,N_29853);
nand UO_631 (O_631,N_25169,N_25939);
xor UO_632 (O_632,N_29228,N_27453);
and UO_633 (O_633,N_24103,N_25303);
or UO_634 (O_634,N_27418,N_24746);
or UO_635 (O_635,N_29527,N_25797);
and UO_636 (O_636,N_27017,N_28830);
or UO_637 (O_637,N_24400,N_26874);
xnor UO_638 (O_638,N_25390,N_29217);
xnor UO_639 (O_639,N_26278,N_24727);
or UO_640 (O_640,N_28725,N_27833);
xnor UO_641 (O_641,N_25664,N_26103);
nand UO_642 (O_642,N_26492,N_29165);
and UO_643 (O_643,N_24993,N_27869);
and UO_644 (O_644,N_27760,N_27362);
or UO_645 (O_645,N_25485,N_28026);
or UO_646 (O_646,N_29991,N_28317);
xnor UO_647 (O_647,N_24995,N_28041);
or UO_648 (O_648,N_26828,N_24264);
or UO_649 (O_649,N_25749,N_28819);
nand UO_650 (O_650,N_24457,N_24212);
xor UO_651 (O_651,N_26595,N_27672);
nand UO_652 (O_652,N_25033,N_28649);
and UO_653 (O_653,N_28498,N_24288);
and UO_654 (O_654,N_27692,N_28373);
nor UO_655 (O_655,N_27359,N_27072);
or UO_656 (O_656,N_28121,N_26640);
xor UO_657 (O_657,N_29634,N_28557);
nor UO_658 (O_658,N_25298,N_29936);
nand UO_659 (O_659,N_27895,N_26012);
xor UO_660 (O_660,N_25457,N_27466);
nor UO_661 (O_661,N_27176,N_29523);
nor UO_662 (O_662,N_24996,N_27697);
nor UO_663 (O_663,N_24668,N_27787);
or UO_664 (O_664,N_26752,N_27088);
nand UO_665 (O_665,N_29781,N_25319);
and UO_666 (O_666,N_25401,N_24462);
or UO_667 (O_667,N_26578,N_28556);
nand UO_668 (O_668,N_26781,N_26686);
nor UO_669 (O_669,N_27912,N_27477);
nand UO_670 (O_670,N_27673,N_26477);
nor UO_671 (O_671,N_25416,N_26986);
nor UO_672 (O_672,N_28987,N_25589);
or UO_673 (O_673,N_25084,N_29556);
or UO_674 (O_674,N_29571,N_26647);
nor UO_675 (O_675,N_24060,N_24773);
and UO_676 (O_676,N_24820,N_29515);
or UO_677 (O_677,N_28661,N_24067);
xnor UO_678 (O_678,N_28568,N_25511);
xnor UO_679 (O_679,N_24711,N_24215);
nand UO_680 (O_680,N_27876,N_28800);
nand UO_681 (O_681,N_24483,N_28840);
nor UO_682 (O_682,N_27378,N_28005);
and UO_683 (O_683,N_26700,N_26614);
and UO_684 (O_684,N_25875,N_25918);
nand UO_685 (O_685,N_27610,N_29430);
xor UO_686 (O_686,N_26581,N_26057);
nor UO_687 (O_687,N_25090,N_25741);
nand UO_688 (O_688,N_28582,N_27880);
xor UO_689 (O_689,N_24127,N_27778);
xnor UO_690 (O_690,N_27483,N_28827);
xnor UO_691 (O_691,N_28184,N_28969);
and UO_692 (O_692,N_28146,N_26713);
xor UO_693 (O_693,N_28633,N_26657);
and UO_694 (O_694,N_25738,N_27214);
nor UO_695 (O_695,N_27093,N_29379);
or UO_696 (O_696,N_28770,N_24100);
nor UO_697 (O_697,N_28326,N_29357);
xor UO_698 (O_698,N_27932,N_24309);
nand UO_699 (O_699,N_28794,N_27941);
nand UO_700 (O_700,N_24939,N_28578);
or UO_701 (O_701,N_27529,N_27062);
nand UO_702 (O_702,N_26959,N_24075);
nand UO_703 (O_703,N_28503,N_28428);
or UO_704 (O_704,N_24775,N_25519);
and UO_705 (O_705,N_29887,N_24585);
or UO_706 (O_706,N_26242,N_27595);
nand UO_707 (O_707,N_27467,N_29630);
nor UO_708 (O_708,N_28337,N_24042);
xor UO_709 (O_709,N_29353,N_28822);
or UO_710 (O_710,N_24026,N_25320);
xor UO_711 (O_711,N_26748,N_24416);
or UO_712 (O_712,N_25063,N_24839);
and UO_713 (O_713,N_25695,N_29939);
xnor UO_714 (O_714,N_25144,N_29587);
xnor UO_715 (O_715,N_25812,N_28083);
and UO_716 (O_716,N_27758,N_25160);
nand UO_717 (O_717,N_25527,N_29476);
xor UO_718 (O_718,N_24852,N_29117);
and UO_719 (O_719,N_24743,N_24178);
nand UO_720 (O_720,N_27561,N_25653);
or UO_721 (O_721,N_24281,N_24358);
nand UO_722 (O_722,N_28413,N_28075);
nand UO_723 (O_723,N_25206,N_25031);
nor UO_724 (O_724,N_29090,N_28404);
nand UO_725 (O_725,N_24747,N_28382);
or UO_726 (O_726,N_27828,N_24137);
or UO_727 (O_727,N_27416,N_24714);
or UO_728 (O_728,N_25809,N_27705);
nor UO_729 (O_729,N_26206,N_29903);
or UO_730 (O_730,N_29134,N_26250);
xor UO_731 (O_731,N_26197,N_27682);
or UO_732 (O_732,N_26714,N_24836);
nor UO_733 (O_733,N_27945,N_26158);
nand UO_734 (O_734,N_26654,N_29996);
nor UO_735 (O_735,N_27271,N_27719);
xnor UO_736 (O_736,N_26040,N_24977);
nand UO_737 (O_737,N_24766,N_24674);
nand UO_738 (O_738,N_24017,N_26484);
nand UO_739 (O_739,N_27915,N_26382);
xnor UO_740 (O_740,N_26568,N_25582);
or UO_741 (O_741,N_27963,N_28791);
nor UO_742 (O_742,N_24649,N_26054);
or UO_743 (O_743,N_29568,N_24135);
nand UO_744 (O_744,N_28902,N_24636);
xnor UO_745 (O_745,N_29053,N_24269);
xor UO_746 (O_746,N_28946,N_25760);
nor UO_747 (O_747,N_29407,N_29953);
nand UO_748 (O_748,N_28034,N_29268);
and UO_749 (O_749,N_28768,N_28672);
or UO_750 (O_750,N_29299,N_24113);
xnor UO_751 (O_751,N_29460,N_26447);
and UO_752 (O_752,N_24139,N_25380);
xnor UO_753 (O_753,N_24289,N_29465);
and UO_754 (O_754,N_25801,N_27473);
xnor UO_755 (O_755,N_29600,N_26095);
xor UO_756 (O_756,N_26569,N_28728);
nand UO_757 (O_757,N_29258,N_24582);
xnor UO_758 (O_758,N_27496,N_26102);
xnor UO_759 (O_759,N_27553,N_26617);
nand UO_760 (O_760,N_25850,N_29855);
nand UO_761 (O_761,N_27742,N_25557);
or UO_762 (O_762,N_24843,N_28621);
xor UO_763 (O_763,N_28668,N_26135);
nor UO_764 (O_764,N_28105,N_29341);
nor UO_765 (O_765,N_24126,N_28248);
and UO_766 (O_766,N_29155,N_29795);
nor UO_767 (O_767,N_27400,N_29231);
or UO_768 (O_768,N_28335,N_29859);
and UO_769 (O_769,N_25995,N_26146);
and UO_770 (O_770,N_25065,N_27660);
xor UO_771 (O_771,N_26360,N_26535);
and UO_772 (O_772,N_25114,N_26577);
nor UO_773 (O_773,N_28514,N_29888);
nand UO_774 (O_774,N_26157,N_25717);
nor UO_775 (O_775,N_29216,N_29366);
xnor UO_776 (O_776,N_24737,N_24580);
xor UO_777 (O_777,N_27928,N_25539);
nor UO_778 (O_778,N_28595,N_27287);
nor UO_779 (O_779,N_24332,N_28047);
xor UO_780 (O_780,N_29377,N_28874);
nand UO_781 (O_781,N_27335,N_24308);
or UO_782 (O_782,N_25193,N_27510);
nor UO_783 (O_783,N_29502,N_26822);
or UO_784 (O_784,N_28838,N_27569);
and UO_785 (O_785,N_27694,N_26138);
nand UO_786 (O_786,N_25061,N_28423);
or UO_787 (O_787,N_27604,N_28564);
nand UO_788 (O_788,N_26645,N_25516);
xnor UO_789 (O_789,N_24906,N_28288);
nand UO_790 (O_790,N_24010,N_26263);
and UO_791 (O_791,N_28634,N_28635);
or UO_792 (O_792,N_24909,N_29352);
nor UO_793 (O_793,N_29203,N_26175);
and UO_794 (O_794,N_27717,N_25507);
xnor UO_795 (O_795,N_26691,N_28982);
and UO_796 (O_796,N_26556,N_29141);
nand UO_797 (O_797,N_28860,N_28594);
nand UO_798 (O_798,N_28736,N_27925);
nand UO_799 (O_799,N_28903,N_26418);
xnor UO_800 (O_800,N_26293,N_24678);
xnor UO_801 (O_801,N_29171,N_27054);
or UO_802 (O_802,N_25896,N_25455);
and UO_803 (O_803,N_27675,N_24947);
nor UO_804 (O_804,N_25458,N_26562);
nor UO_805 (O_805,N_28329,N_28505);
and UO_806 (O_806,N_26609,N_27488);
nor UO_807 (O_807,N_28648,N_24624);
and UO_808 (O_808,N_29047,N_24225);
or UO_809 (O_809,N_29982,N_26706);
xnor UO_810 (O_810,N_29088,N_29849);
nor UO_811 (O_811,N_26072,N_25775);
xor UO_812 (O_812,N_27517,N_24535);
nand UO_813 (O_813,N_28290,N_29213);
and UO_814 (O_814,N_25153,N_29204);
or UO_815 (O_815,N_27209,N_28760);
and UO_816 (O_816,N_26520,N_25461);
nor UO_817 (O_817,N_29666,N_28615);
and UO_818 (O_818,N_29779,N_28054);
and UO_819 (O_819,N_28087,N_29915);
xor UO_820 (O_820,N_24427,N_25011);
nor UO_821 (O_821,N_29851,N_26214);
nand UO_822 (O_822,N_25893,N_28254);
nor UO_823 (O_823,N_27469,N_29637);
xor UO_824 (O_824,N_26215,N_24776);
or UO_825 (O_825,N_24786,N_25345);
nor UO_826 (O_826,N_25396,N_27332);
xnor UO_827 (O_827,N_25074,N_28283);
nand UO_828 (O_828,N_24224,N_27279);
and UO_829 (O_829,N_26644,N_26809);
xnor UO_830 (O_830,N_26174,N_28374);
nand UO_831 (O_831,N_29900,N_26594);
or UO_832 (O_832,N_26867,N_29418);
and UO_833 (O_833,N_29797,N_25865);
and UO_834 (O_834,N_24866,N_28108);
nor UO_835 (O_835,N_27458,N_26717);
or UO_836 (O_836,N_25502,N_29256);
xnor UO_837 (O_837,N_27041,N_26953);
xnor UO_838 (O_838,N_26342,N_28681);
and UO_839 (O_839,N_28124,N_27337);
xnor UO_840 (O_840,N_29376,N_26934);
or UO_841 (O_841,N_25282,N_24625);
xor UO_842 (O_842,N_26245,N_28464);
or UO_843 (O_843,N_28985,N_26323);
nor UO_844 (O_844,N_25703,N_26696);
and UO_845 (O_845,N_29550,N_29599);
xor UO_846 (O_846,N_28493,N_26130);
xnor UO_847 (O_847,N_25734,N_27617);
or UO_848 (O_848,N_25157,N_25707);
xnor UO_849 (O_849,N_24889,N_28424);
or UO_850 (O_850,N_25640,N_29608);
xor UO_851 (O_851,N_24827,N_25276);
and UO_852 (O_852,N_25628,N_26872);
xor UO_853 (O_853,N_27022,N_24658);
nand UO_854 (O_854,N_24324,N_28960);
and UO_855 (O_855,N_24847,N_25699);
nand UO_856 (O_856,N_29249,N_25877);
nand UO_857 (O_857,N_27383,N_29102);
nand UO_858 (O_858,N_29760,N_27518);
or UO_859 (O_859,N_29063,N_29237);
or UO_860 (O_860,N_26079,N_28839);
or UO_861 (O_861,N_28617,N_26852);
xor UO_862 (O_862,N_26790,N_26539);
nor UO_863 (O_863,N_26747,N_24953);
or UO_864 (O_864,N_28450,N_29656);
nand UO_865 (O_865,N_25332,N_25400);
xor UO_866 (O_866,N_27138,N_25293);
xor UO_867 (O_867,N_26807,N_29759);
xnor UO_868 (O_868,N_29560,N_26927);
xnor UO_869 (O_869,N_25389,N_26642);
or UO_870 (O_870,N_24870,N_29232);
and UO_871 (O_871,N_28015,N_28304);
xor UO_872 (O_872,N_29489,N_29413);
xnor UO_873 (O_873,N_29411,N_25718);
or UO_874 (O_874,N_25894,N_27640);
nor UO_875 (O_875,N_27998,N_29983);
and UO_876 (O_876,N_26522,N_28010);
nor UO_877 (O_877,N_28756,N_28862);
nor UO_878 (O_878,N_25349,N_29072);
nor UO_879 (O_879,N_28222,N_26004);
or UO_880 (O_880,N_25821,N_27126);
nand UO_881 (O_881,N_24230,N_25295);
xnor UO_882 (O_882,N_24446,N_27230);
or UO_883 (O_883,N_26356,N_25331);
nand UO_884 (O_884,N_26880,N_29628);
xnor UO_885 (O_885,N_29447,N_26690);
xnor UO_886 (O_886,N_25382,N_25451);
nand UO_887 (O_887,N_28049,N_24449);
and UO_888 (O_888,N_28817,N_24581);
nand UO_889 (O_889,N_28255,N_24612);
or UO_890 (O_890,N_26983,N_26658);
xor UO_891 (O_891,N_28996,N_27053);
and UO_892 (O_892,N_28821,N_28761);
and UO_893 (O_893,N_28892,N_27440);
or UO_894 (O_894,N_29118,N_29884);
and UO_895 (O_895,N_26941,N_28675);
or UO_896 (O_896,N_24220,N_29576);
and UO_897 (O_897,N_28758,N_25565);
and UO_898 (O_898,N_26283,N_25880);
xor UO_899 (O_899,N_28268,N_28463);
or UO_900 (O_900,N_24887,N_28771);
nor UO_901 (O_901,N_24216,N_28778);
nand UO_902 (O_902,N_25035,N_24734);
nor UO_903 (O_903,N_25460,N_24131);
and UO_904 (O_904,N_29555,N_26820);
xor UO_905 (O_905,N_24278,N_27848);
and UO_906 (O_906,N_26886,N_26625);
xnor UO_907 (O_907,N_27500,N_29559);
or UO_908 (O_908,N_27670,N_28340);
nor UO_909 (O_909,N_27382,N_26912);
xnor UO_910 (O_910,N_28624,N_24630);
and UO_911 (O_911,N_28096,N_27780);
or UO_912 (O_912,N_28457,N_26682);
xnor UO_913 (O_913,N_28922,N_27871);
nand UO_914 (O_914,N_28563,N_24793);
or UO_915 (O_915,N_26119,N_24219);
nand UO_916 (O_916,N_25051,N_28399);
xnor UO_917 (O_917,N_25432,N_29238);
or UO_918 (O_918,N_28640,N_29720);
nor UO_919 (O_919,N_28187,N_29112);
xnor UO_920 (O_920,N_29294,N_26715);
xor UO_921 (O_921,N_25249,N_25928);
or UO_922 (O_922,N_28585,N_28574);
or UO_923 (O_923,N_26712,N_25375);
nand UO_924 (O_924,N_24437,N_27050);
xor UO_925 (O_925,N_24932,N_29601);
nand UO_926 (O_926,N_27520,N_29142);
or UO_927 (O_927,N_27695,N_28163);
and UO_928 (O_928,N_27607,N_28176);
nor UO_929 (O_929,N_25780,N_26591);
xnor UO_930 (O_930,N_26159,N_29126);
and UO_931 (O_931,N_27560,N_29975);
nor UO_932 (O_932,N_24611,N_25960);
nand UO_933 (O_933,N_25056,N_27807);
nor UO_934 (O_934,N_25605,N_28942);
nand UO_935 (O_935,N_26318,N_25905);
nor UO_936 (O_936,N_28321,N_24194);
nor UO_937 (O_937,N_27732,N_24466);
nand UO_938 (O_938,N_24760,N_29078);
or UO_939 (O_939,N_27770,N_28694);
and UO_940 (O_940,N_28806,N_24829);
and UO_941 (O_941,N_27207,N_28589);
or UO_942 (O_942,N_29667,N_24340);
nand UO_943 (O_943,N_27159,N_25286);
or UO_944 (O_944,N_25313,N_29259);
xnor UO_945 (O_945,N_25415,N_29920);
nand UO_946 (O_946,N_25304,N_27919);
nand UO_947 (O_947,N_29776,N_26877);
or UO_948 (O_948,N_26695,N_24818);
or UO_949 (O_949,N_29771,N_28558);
nor UO_950 (O_950,N_26888,N_24515);
or UO_951 (O_951,N_26400,N_25621);
and UO_952 (O_952,N_27091,N_26674);
nor UO_953 (O_953,N_25899,N_25092);
and UO_954 (O_954,N_28591,N_28323);
nor UO_955 (O_955,N_27573,N_26246);
or UO_956 (O_956,N_25558,N_26949);
nand UO_957 (O_957,N_26773,N_29742);
or UO_958 (O_958,N_24039,N_27024);
or UO_959 (O_959,N_29186,N_24438);
xor UO_960 (O_960,N_26588,N_29074);
nand UO_961 (O_961,N_26683,N_29661);
xor UO_962 (O_962,N_25710,N_27094);
and UO_963 (O_963,N_26547,N_24154);
and UO_964 (O_964,N_24733,N_24748);
xnor UO_965 (O_965,N_28609,N_29331);
xnor UO_966 (O_966,N_26265,N_28851);
and UO_967 (O_967,N_27903,N_26856);
nand UO_968 (O_968,N_28604,N_29516);
and UO_969 (O_969,N_25071,N_26039);
and UO_970 (O_970,N_29224,N_28717);
nor UO_971 (O_971,N_26887,N_27562);
nor UO_972 (O_972,N_27687,N_25783);
nand UO_973 (O_973,N_25205,N_27734);
or UO_974 (O_974,N_27678,N_29958);
nor UO_975 (O_975,N_25435,N_25756);
nand UO_976 (O_976,N_26794,N_28149);
xnor UO_977 (O_977,N_29789,N_28951);
xnor UO_978 (O_978,N_26507,N_29338);
and UO_979 (O_979,N_26728,N_25613);
and UO_980 (O_980,N_25976,N_27891);
nand UO_981 (O_981,N_27922,N_27616);
or UO_982 (O_982,N_28831,N_27048);
nor UO_983 (O_983,N_29805,N_28590);
and UO_984 (O_984,N_24360,N_28023);
nand UO_985 (O_985,N_24545,N_26906);
and UO_986 (O_986,N_29828,N_24946);
nand UO_987 (O_987,N_25032,N_26795);
nor UO_988 (O_988,N_29021,N_28795);
and UO_989 (O_989,N_25306,N_29757);
nand UO_990 (O_990,N_29626,N_25050);
xor UO_991 (O_991,N_28038,N_24261);
and UO_992 (O_992,N_25889,N_26729);
nand UO_993 (O_993,N_26350,N_26734);
xnor UO_994 (O_994,N_25310,N_25494);
xor UO_995 (O_995,N_24560,N_24203);
nand UO_996 (O_996,N_29361,N_24397);
nor UO_997 (O_997,N_26586,N_29473);
nand UO_998 (O_998,N_25374,N_26663);
xor UO_999 (O_999,N_29092,N_28971);
xor UO_1000 (O_1000,N_28186,N_26560);
nand UO_1001 (O_1001,N_28064,N_26388);
or UO_1002 (O_1002,N_29133,N_25139);
or UO_1003 (O_1003,N_25020,N_27480);
xor UO_1004 (O_1004,N_28779,N_25970);
and UO_1005 (O_1005,N_29609,N_25000);
nor UO_1006 (O_1006,N_29310,N_26416);
and UO_1007 (O_1007,N_27060,N_26665);
nor UO_1008 (O_1008,N_25708,N_29390);
nand UO_1009 (O_1009,N_28346,N_24538);
nor UO_1010 (O_1010,N_28709,N_25222);
or UO_1011 (O_1011,N_24681,N_28955);
nor UO_1012 (O_1012,N_29025,N_28289);
and UO_1013 (O_1013,N_29719,N_24978);
and UO_1014 (O_1014,N_29641,N_28528);
xor UO_1015 (O_1015,N_26619,N_26366);
nand UO_1016 (O_1016,N_26111,N_24011);
and UO_1017 (O_1017,N_25822,N_25852);
xor UO_1018 (O_1018,N_29006,N_26991);
xnor UO_1019 (O_1019,N_27244,N_29189);
and UO_1020 (O_1020,N_29944,N_26134);
and UO_1021 (O_1021,N_27982,N_27767);
or UO_1022 (O_1022,N_24752,N_29921);
and UO_1023 (O_1023,N_26059,N_28577);
nand UO_1024 (O_1024,N_28952,N_24363);
or UO_1025 (O_1025,N_24081,N_27648);
nand UO_1026 (O_1026,N_29395,N_24803);
nand UO_1027 (O_1027,N_27940,N_25977);
and UO_1028 (O_1028,N_26473,N_29874);
nand UO_1029 (O_1029,N_28995,N_27586);
nand UO_1030 (O_1030,N_26744,N_27016);
or UO_1031 (O_1031,N_26455,N_29941);
xnor UO_1032 (O_1032,N_27341,N_28658);
nand UO_1033 (O_1033,N_29028,N_25475);
xnor UO_1034 (O_1034,N_29143,N_27168);
nor UO_1035 (O_1035,N_26145,N_27164);
and UO_1036 (O_1036,N_24033,N_25037);
nor UO_1037 (O_1037,N_26450,N_28192);
and UO_1038 (O_1038,N_27868,N_25012);
xor UO_1039 (O_1039,N_25045,N_28451);
xnor UO_1040 (O_1040,N_27856,N_24246);
xor UO_1041 (O_1041,N_26840,N_24481);
nand UO_1042 (O_1042,N_25721,N_29736);
nand UO_1043 (O_1043,N_26043,N_26036);
nor UO_1044 (O_1044,N_25862,N_27107);
nand UO_1045 (O_1045,N_27067,N_29247);
nor UO_1046 (O_1046,N_25150,N_24442);
nor UO_1047 (O_1047,N_27152,N_24600);
nand UO_1048 (O_1048,N_29962,N_28665);
or UO_1049 (O_1049,N_29332,N_28861);
nor UO_1050 (O_1050,N_29230,N_28854);
nor UO_1051 (O_1051,N_25449,N_24972);
nor UO_1052 (O_1052,N_27239,N_27693);
nor UO_1053 (O_1053,N_29381,N_28704);
xnor UO_1054 (O_1054,N_28065,N_24285);
nor UO_1055 (O_1055,N_25848,N_25217);
nor UO_1056 (O_1056,N_24774,N_24588);
and UO_1057 (O_1057,N_27786,N_27618);
nor UO_1058 (O_1058,N_25196,N_25419);
nor UO_1059 (O_1059,N_29007,N_25234);
nand UO_1060 (O_1060,N_28348,N_28975);
xnor UO_1061 (O_1061,N_26739,N_24574);
xor UO_1062 (O_1062,N_29378,N_24403);
nand UO_1063 (O_1063,N_28259,N_27033);
nor UO_1064 (O_1064,N_27997,N_27906);
nand UO_1065 (O_1065,N_25379,N_25524);
and UO_1066 (O_1066,N_26429,N_24197);
and UO_1067 (O_1067,N_28266,N_29800);
nor UO_1068 (O_1068,N_25870,N_26122);
nand UO_1069 (O_1069,N_29883,N_24458);
xnor UO_1070 (O_1070,N_24274,N_24108);
and UO_1071 (O_1071,N_28486,N_25567);
nor UO_1072 (O_1072,N_26505,N_29540);
xnor UO_1073 (O_1073,N_24750,N_24448);
xnor UO_1074 (O_1074,N_28759,N_26805);
and UO_1075 (O_1075,N_24777,N_26226);
nor UO_1076 (O_1076,N_25425,N_25339);
nor UO_1077 (O_1077,N_25636,N_27389);
xor UO_1078 (O_1078,N_29627,N_27943);
nor UO_1079 (O_1079,N_26508,N_24120);
or UO_1080 (O_1080,N_29840,N_28044);
and UO_1081 (O_1081,N_26190,N_28239);
nor UO_1082 (O_1082,N_24837,N_24599);
nor UO_1083 (O_1083,N_24507,N_28212);
and UO_1084 (O_1084,N_24118,N_28025);
xnor UO_1085 (O_1085,N_28261,N_26628);
nand UO_1086 (O_1086,N_25956,N_25218);
and UO_1087 (O_1087,N_25713,N_26530);
nor UO_1088 (O_1088,N_24085,N_29697);
nor UO_1089 (O_1089,N_25147,N_28291);
xnor UO_1090 (O_1090,N_29901,N_29392);
nand UO_1091 (O_1091,N_24640,N_25212);
nor UO_1092 (O_1092,N_29002,N_27056);
nand UO_1093 (O_1093,N_27578,N_28636);
and UO_1094 (O_1094,N_29728,N_26889);
or UO_1095 (O_1095,N_25803,N_25387);
nand UO_1096 (O_1096,N_29099,N_25903);
or UO_1097 (O_1097,N_29210,N_26334);
or UO_1098 (O_1098,N_27083,N_25357);
nand UO_1099 (O_1099,N_25955,N_26434);
and UO_1100 (O_1100,N_26013,N_28523);
xor UO_1101 (O_1101,N_29371,N_29111);
or UO_1102 (O_1102,N_26973,N_26512);
and UO_1103 (O_1103,N_29008,N_27588);
nor UO_1104 (O_1104,N_26442,N_24307);
or UO_1105 (O_1105,N_28492,N_26845);
nand UO_1106 (O_1106,N_26073,N_26476);
nand UO_1107 (O_1107,N_28410,N_29293);
and UO_1108 (O_1108,N_26349,N_28509);
nor UO_1109 (O_1109,N_27509,N_29992);
xor UO_1110 (O_1110,N_26425,N_28696);
nor UO_1111 (O_1111,N_29168,N_28220);
or UO_1112 (O_1112,N_25059,N_29163);
and UO_1113 (O_1113,N_28079,N_27887);
and UO_1114 (O_1114,N_28221,N_26076);
nand UO_1115 (O_1115,N_28565,N_25280);
xor UO_1116 (O_1116,N_26401,N_29335);
nand UO_1117 (O_1117,N_27334,N_28217);
nand UO_1118 (O_1118,N_25758,N_28703);
nand UO_1119 (O_1119,N_29506,N_29084);
and UO_1120 (O_1120,N_28420,N_25548);
or UO_1121 (O_1121,N_27059,N_25663);
and UO_1122 (O_1122,N_25652,N_25747);
and UO_1123 (O_1123,N_24221,N_26304);
nor UO_1124 (O_1124,N_27305,N_29384);
nand UO_1125 (O_1125,N_29490,N_24072);
xnor UO_1126 (O_1126,N_26899,N_25164);
xor UO_1127 (O_1127,N_26015,N_28195);
and UO_1128 (O_1128,N_26861,N_24722);
xor UO_1129 (O_1129,N_26149,N_28355);
or UO_1130 (O_1130,N_26277,N_26834);
nand UO_1131 (O_1131,N_27046,N_27219);
nor UO_1132 (O_1132,N_25962,N_29116);
or UO_1133 (O_1133,N_28679,N_25263);
nand UO_1134 (O_1134,N_29267,N_24952);
nor UO_1135 (O_1135,N_25273,N_25335);
nor UO_1136 (O_1136,N_27425,N_25473);
nand UO_1137 (O_1137,N_29274,N_24541);
nand UO_1138 (O_1138,N_27547,N_28198);
or UO_1139 (O_1139,N_28906,N_26846);
nand UO_1140 (O_1140,N_26621,N_28086);
and UO_1141 (O_1141,N_24495,N_25115);
and UO_1142 (O_1142,N_28052,N_26669);
nor UO_1143 (O_1143,N_24208,N_25658);
or UO_1144 (O_1144,N_29202,N_25110);
nand UO_1145 (O_1145,N_29943,N_26207);
nor UO_1146 (O_1146,N_29010,N_29535);
xnor UO_1147 (O_1147,N_29286,N_25627);
or UO_1148 (O_1148,N_26848,N_29548);
nand UO_1149 (O_1149,N_27638,N_29708);
nor UO_1150 (O_1150,N_25932,N_25834);
nand UO_1151 (O_1151,N_26116,N_26469);
and UO_1152 (O_1152,N_24111,N_24133);
nor UO_1153 (O_1153,N_25123,N_29544);
nand UO_1154 (O_1154,N_26237,N_26575);
nor UO_1155 (O_1155,N_29913,N_26087);
nor UO_1156 (O_1156,N_29448,N_26838);
and UO_1157 (O_1157,N_26422,N_24179);
nor UO_1158 (O_1158,N_24142,N_26989);
and UO_1159 (O_1159,N_25796,N_24801);
xor UO_1160 (O_1160,N_25933,N_25694);
xor UO_1161 (O_1161,N_26383,N_26071);
nand UO_1162 (O_1162,N_25260,N_29456);
nand UO_1163 (O_1163,N_28910,N_24372);
and UO_1164 (O_1164,N_29882,N_25737);
xor UO_1165 (O_1165,N_29057,N_27950);
or UO_1166 (O_1166,N_26664,N_29080);
xnor UO_1167 (O_1167,N_26635,N_28110);
xnor UO_1168 (O_1168,N_28745,N_24134);
or UO_1169 (O_1169,N_29431,N_24065);
or UO_1170 (O_1170,N_25917,N_25512);
xnor UO_1171 (O_1171,N_28555,N_24005);
xor UO_1172 (O_1172,N_25838,N_26653);
nand UO_1173 (O_1173,N_27437,N_27267);
and UO_1174 (O_1174,N_24530,N_28647);
and UO_1175 (O_1175,N_25913,N_24713);
nand UO_1176 (O_1176,N_25807,N_24785);
xnor UO_1177 (O_1177,N_25130,N_27369);
and UO_1178 (O_1178,N_25689,N_27803);
nand UO_1179 (O_1179,N_27599,N_28698);
and UO_1180 (O_1180,N_28918,N_27918);
nor UO_1181 (O_1181,N_27352,N_24290);
nor UO_1182 (O_1182,N_28825,N_29011);
xnor UO_1183 (O_1183,N_28078,N_27224);
nand UO_1184 (O_1184,N_25569,N_26515);
or UO_1185 (O_1185,N_25083,N_29159);
nor UO_1186 (O_1186,N_28353,N_24336);
and UO_1187 (O_1187,N_28093,N_24257);
nor UO_1188 (O_1188,N_29346,N_27444);
and UO_1189 (O_1189,N_25603,N_29860);
nand UO_1190 (O_1190,N_28123,N_24689);
nand UO_1191 (O_1191,N_24019,N_24171);
or UO_1192 (O_1192,N_27612,N_29889);
and UO_1193 (O_1193,N_25159,N_25999);
nor UO_1194 (O_1194,N_27063,N_24392);
xnor UO_1195 (O_1195,N_28646,N_27862);
nand UO_1196 (O_1196,N_29932,N_24838);
or UO_1197 (O_1197,N_29688,N_24123);
or UO_1198 (O_1198,N_27892,N_29981);
and UO_1199 (O_1199,N_28880,N_28964);
nor UO_1200 (O_1200,N_26836,N_29931);
nand UO_1201 (O_1201,N_24032,N_27112);
and UO_1202 (O_1202,N_26716,N_28573);
and UO_1203 (O_1203,N_24028,N_24088);
and UO_1204 (O_1204,N_24557,N_25909);
xor UO_1205 (O_1205,N_25294,N_29787);
and UO_1206 (O_1206,N_28797,N_25890);
nand UO_1207 (O_1207,N_26424,N_25779);
or UO_1208 (O_1208,N_24536,N_27103);
and UO_1209 (O_1209,N_29702,N_27541);
nand UO_1210 (O_1210,N_27375,N_26890);
and UO_1211 (O_1211,N_28487,N_28738);
nor UO_1212 (O_1212,N_25634,N_25358);
xnor UO_1213 (O_1213,N_27969,N_27409);
nand UO_1214 (O_1214,N_29543,N_27995);
or UO_1215 (O_1215,N_24919,N_25542);
nand UO_1216 (O_1216,N_28909,N_27766);
nor UO_1217 (O_1217,N_28488,N_28613);
or UO_1218 (O_1218,N_24369,N_26056);
nor UO_1219 (O_1219,N_29180,N_27592);
xnor UO_1220 (O_1220,N_24314,N_24591);
or UO_1221 (O_1221,N_27411,N_29375);
nand UO_1222 (O_1222,N_26910,N_27474);
xor UO_1223 (O_1223,N_24128,N_27563);
xnor UO_1224 (O_1224,N_26919,N_29065);
and UO_1225 (O_1225,N_27783,N_27589);
nand UO_1226 (O_1226,N_25782,N_29919);
and UO_1227 (O_1227,N_29169,N_25651);
and UO_1228 (O_1228,N_25053,N_24701);
nand UO_1229 (O_1229,N_28479,N_25883);
nand UO_1230 (O_1230,N_27364,N_26762);
xor UO_1231 (O_1231,N_29013,N_29270);
nand UO_1232 (O_1232,N_29904,N_29841);
xor UO_1233 (O_1233,N_29042,N_27465);
or UO_1234 (O_1234,N_26274,N_24863);
nor UO_1235 (O_1235,N_28938,N_28418);
and UO_1236 (O_1236,N_25411,N_26570);
or UO_1237 (O_1237,N_26776,N_28579);
xor UO_1238 (O_1238,N_28744,N_24783);
nor UO_1239 (O_1239,N_27301,N_25778);
xnor UO_1240 (O_1240,N_25237,N_28638);
or UO_1241 (O_1241,N_27977,N_27857);
nor UO_1242 (O_1242,N_24317,N_28815);
and UO_1243 (O_1243,N_29164,N_25854);
nor UO_1244 (O_1244,N_29509,N_27413);
nand UO_1245 (O_1245,N_26750,N_29949);
or UO_1246 (O_1246,N_29316,N_29940);
nand UO_1247 (O_1247,N_28292,N_26955);
xor UO_1248 (O_1248,N_27722,N_29326);
and UO_1249 (O_1249,N_25800,N_25815);
nand UO_1250 (O_1250,N_25436,N_25765);
nand UO_1251 (O_1251,N_28662,N_25773);
and UO_1252 (O_1252,N_28397,N_25543);
xnor UO_1253 (O_1253,N_24249,N_24594);
and UO_1254 (O_1254,N_26566,N_29700);
nand UO_1255 (O_1255,N_29875,N_29735);
nor UO_1256 (O_1256,N_29670,N_25926);
or UO_1257 (O_1257,N_25921,N_29906);
and UO_1258 (O_1258,N_27172,N_24670);
nand UO_1259 (O_1259,N_28475,N_24306);
xor UO_1260 (O_1260,N_29866,N_26559);
nor UO_1261 (O_1261,N_25235,N_27484);
or UO_1262 (O_1262,N_24153,N_29786);
nor UO_1263 (O_1263,N_29682,N_28278);
nor UO_1264 (O_1264,N_28443,N_26109);
nand UO_1265 (O_1265,N_28620,N_24351);
xor UO_1266 (O_1266,N_26580,N_24044);
nor UO_1267 (O_1267,N_25483,N_25802);
xor UO_1268 (O_1268,N_27406,N_24478);
or UO_1269 (O_1269,N_24076,N_29220);
or UO_1270 (O_1270,N_29674,N_25299);
xnor UO_1271 (O_1271,N_24526,N_29240);
nor UO_1272 (O_1272,N_26814,N_25399);
nor UO_1273 (O_1273,N_25980,N_28529);
nor UO_1274 (O_1274,N_24006,N_25178);
or UO_1275 (O_1275,N_26679,N_26448);
and UO_1276 (O_1276,N_28972,N_27426);
nand UO_1277 (O_1277,N_26205,N_26693);
nand UO_1278 (O_1278,N_24175,N_27799);
nand UO_1279 (O_1279,N_24015,N_26769);
or UO_1280 (O_1280,N_24426,N_24954);
and UO_1281 (O_1281,N_27468,N_25272);
and UO_1282 (O_1282,N_26514,N_28896);
and UO_1283 (O_1283,N_24251,N_28115);
or UO_1284 (O_1284,N_26534,N_25245);
and UO_1285 (O_1285,N_25911,N_27065);
and UO_1286 (O_1286,N_25967,N_24490);
and UO_1287 (O_1287,N_27356,N_29107);
nor UO_1288 (O_1288,N_28974,N_27285);
xor UO_1289 (O_1289,N_29101,N_25448);
and UO_1290 (O_1290,N_26601,N_27042);
nor UO_1291 (O_1291,N_29468,N_24461);
and UO_1292 (O_1292,N_24877,N_28685);
or UO_1293 (O_1293,N_25132,N_28050);
and UO_1294 (O_1294,N_26792,N_29422);
nand UO_1295 (O_1295,N_25474,N_27600);
and UO_1296 (O_1296,N_25073,N_26098);
xor UO_1297 (O_1297,N_29271,N_29137);
nand UO_1298 (O_1298,N_26280,N_26573);
xnor UO_1299 (O_1299,N_28363,N_28664);
and UO_1300 (O_1300,N_24361,N_26289);
and UO_1301 (O_1301,N_26965,N_26966);
or UO_1302 (O_1302,N_24077,N_24243);
nand UO_1303 (O_1303,N_27058,N_24465);
and UO_1304 (O_1304,N_28958,N_28104);
or UO_1305 (O_1305,N_25836,N_25957);
or UO_1306 (O_1306,N_24587,N_29255);
nand UO_1307 (O_1307,N_26632,N_26996);
nand UO_1308 (O_1308,N_28381,N_24090);
and UO_1309 (O_1309,N_26869,N_27456);
nand UO_1310 (O_1310,N_28393,N_24012);
nor UO_1311 (O_1311,N_29978,N_27037);
nor UO_1312 (O_1312,N_29318,N_25289);
and UO_1313 (O_1313,N_26914,N_28707);
or UO_1314 (O_1314,N_29435,N_25518);
xor UO_1315 (O_1315,N_27197,N_24572);
nor UO_1316 (O_1316,N_27654,N_27387);
nor UO_1317 (O_1317,N_28398,N_28280);
nor UO_1318 (O_1318,N_24592,N_25701);
nor UO_1319 (O_1319,N_28437,N_27211);
or UO_1320 (O_1320,N_29896,N_27593);
or UO_1321 (O_1321,N_28085,N_28610);
or UO_1322 (O_1322,N_26251,N_29815);
xnor UO_1323 (O_1323,N_29161,N_27195);
nor UO_1324 (O_1324,N_28333,N_28231);
nand UO_1325 (O_1325,N_26649,N_24567);
nor UO_1326 (O_1326,N_27988,N_24555);
and UO_1327 (O_1327,N_26753,N_26474);
and UO_1328 (O_1328,N_25853,N_28569);
and UO_1329 (O_1329,N_25541,N_26873);
xnor UO_1330 (O_1330,N_25456,N_29356);
and UO_1331 (O_1331,N_26970,N_28202);
nand UO_1332 (O_1332,N_28448,N_24616);
or UO_1333 (O_1333,N_27993,N_26273);
or UO_1334 (O_1334,N_25467,N_27026);
xor UO_1335 (O_1335,N_25600,N_28389);
nor UO_1336 (O_1336,N_29399,N_25670);
nand UO_1337 (O_1337,N_28605,N_25009);
or UO_1338 (O_1338,N_28994,N_25873);
and UO_1339 (O_1339,N_28833,N_26153);
and UO_1340 (O_1340,N_26740,N_28750);
or UO_1341 (O_1341,N_25958,N_26493);
nor UO_1342 (O_1342,N_29351,N_25826);
nor UO_1343 (O_1343,N_29205,N_27701);
and UO_1344 (O_1344,N_25438,N_26893);
nand UO_1345 (O_1345,N_25813,N_29524);
nor UO_1346 (O_1346,N_28935,N_24744);
nand UO_1347 (O_1347,N_29918,N_26823);
nand UO_1348 (O_1348,N_29845,N_26083);
and UO_1349 (O_1349,N_29364,N_26875);
and UO_1350 (O_1350,N_24884,N_27700);
xnor UO_1351 (O_1351,N_24181,N_29922);
nand UO_1352 (O_1352,N_28432,N_28721);
nand UO_1353 (O_1353,N_29486,N_26307);
xor UO_1354 (O_1354,N_28406,N_24211);
nor UO_1355 (O_1355,N_25497,N_29780);
nor UO_1356 (O_1356,N_24505,N_27652);
and UO_1357 (O_1357,N_29471,N_28031);
and UO_1358 (O_1358,N_24204,N_25079);
nor UO_1359 (O_1359,N_27081,N_27459);
nor UO_1360 (O_1360,N_25740,N_27379);
nor UO_1361 (O_1361,N_29121,N_26248);
xor UO_1362 (O_1362,N_28998,N_26726);
xnor UO_1363 (O_1363,N_27975,N_29825);
and UO_1364 (O_1364,N_28850,N_28062);
xnor UO_1365 (O_1365,N_24698,N_28045);
xor UO_1366 (O_1366,N_27106,N_27397);
xnor UO_1367 (O_1367,N_26011,N_24062);
or UO_1368 (O_1368,N_25257,N_29911);
nand UO_1369 (O_1369,N_29015,N_26380);
nand UO_1370 (O_1370,N_29907,N_24472);
nor UO_1371 (O_1371,N_25018,N_29125);
nor UO_1372 (O_1372,N_26045,N_24109);
or UO_1373 (O_1373,N_26727,N_26897);
xor UO_1374 (O_1374,N_26504,N_27432);
and UO_1375 (O_1375,N_29926,N_25412);
nand UO_1376 (O_1376,N_28324,N_26405);
or UO_1377 (O_1377,N_29207,N_25632);
nor UO_1378 (O_1378,N_25587,N_25296);
nor UO_1379 (O_1379,N_24680,N_25221);
and UO_1380 (O_1380,N_24217,N_24540);
nand UO_1381 (O_1381,N_28848,N_29698);
and UO_1382 (O_1382,N_26256,N_27809);
and UO_1383 (O_1383,N_24967,N_29032);
nand UO_1384 (O_1384,N_29960,N_26523);
nor UO_1385 (O_1385,N_28234,N_24445);
nor UO_1386 (O_1386,N_27021,N_26171);
nor UO_1387 (O_1387,N_26441,N_26481);
nor UO_1388 (O_1388,N_25422,N_26485);
and UO_1389 (O_1389,N_29048,N_25437);
nand UO_1390 (O_1390,N_24174,N_26435);
xor UO_1391 (O_1391,N_25659,N_29615);
xor UO_1392 (O_1392,N_24509,N_27587);
nor UO_1393 (O_1393,N_28032,N_29605);
nand UO_1394 (O_1394,N_26639,N_28925);
and UO_1395 (O_1395,N_26131,N_24940);
xor UO_1396 (O_1396,N_26612,N_29114);
and UO_1397 (O_1397,N_26166,N_27282);
and UO_1398 (O_1398,N_29291,N_26928);
and UO_1399 (O_1399,N_25520,N_28002);
nand UO_1400 (O_1400,N_24632,N_27462);
or UO_1401 (O_1401,N_26689,N_25266);
nand UO_1402 (O_1402,N_24087,N_28150);
nor UO_1403 (O_1403,N_28080,N_29740);
xor UO_1404 (O_1404,N_25158,N_25673);
nand UO_1405 (O_1405,N_26152,N_26249);
xor UO_1406 (O_1406,N_25138,N_25006);
xnor UO_1407 (O_1407,N_24917,N_27899);
nor UO_1408 (O_1408,N_27874,N_24402);
nand UO_1409 (O_1409,N_26177,N_28154);
xnor UO_1410 (O_1410,N_28751,N_29434);
and UO_1411 (O_1411,N_27263,N_29846);
xnor UO_1412 (O_1412,N_24652,N_26667);
or UO_1413 (O_1413,N_26833,N_29450);
xnor UO_1414 (O_1414,N_27668,N_24595);
xor UO_1415 (O_1415,N_29194,N_27099);
nand UO_1416 (O_1416,N_29689,N_26439);
or UO_1417 (O_1417,N_24059,N_27702);
xnor UO_1418 (O_1418,N_28572,N_24605);
nand UO_1419 (O_1419,N_28468,N_28611);
xnor UO_1420 (O_1420,N_25484,N_26025);
nor UO_1421 (O_1421,N_24672,N_25533);
nor UO_1422 (O_1422,N_26046,N_25255);
or UO_1423 (O_1423,N_29606,N_28012);
xor UO_1424 (O_1424,N_25239,N_29620);
nand UO_1425 (O_1425,N_26232,N_27704);
xor UO_1426 (O_1426,N_24856,N_27485);
nor UO_1427 (O_1427,N_27367,N_29178);
xnor UO_1428 (O_1428,N_24506,N_28897);
xnor UO_1429 (O_1429,N_29033,N_24589);
xnor UO_1430 (O_1430,N_25182,N_28245);
or UO_1431 (O_1431,N_27076,N_25402);
nand UO_1432 (O_1432,N_28482,N_24610);
or UO_1433 (O_1433,N_29269,N_25279);
or UO_1434 (O_1434,N_25148,N_26108);
and UO_1435 (O_1435,N_25908,N_25081);
nor UO_1436 (O_1436,N_25792,N_26746);
nand UO_1437 (O_1437,N_26678,N_24502);
or UO_1438 (O_1438,N_28208,N_26398);
nand UO_1439 (O_1439,N_29329,N_25459);
xor UO_1440 (O_1440,N_28705,N_27830);
xnor UO_1441 (O_1441,N_26529,N_26310);
or UO_1442 (O_1442,N_24073,N_27965);
nor UO_1443 (O_1443,N_27657,N_24305);
nand UO_1444 (O_1444,N_24738,N_29541);
xnor UO_1445 (O_1445,N_26498,N_24330);
and UO_1446 (O_1446,N_28539,N_24286);
xnor UO_1447 (O_1447,N_29831,N_29265);
or UO_1448 (O_1448,N_26961,N_28805);
nand UO_1449 (O_1449,N_25365,N_25161);
or UO_1450 (O_1450,N_24091,N_28551);
nor UO_1451 (O_1451,N_27415,N_25536);
and UO_1452 (O_1452,N_28338,N_24647);
and UO_1453 (O_1453,N_24359,N_29562);
or UO_1454 (O_1454,N_29582,N_24424);
xor UO_1455 (O_1455,N_28834,N_24355);
nand UO_1456 (O_1456,N_24522,N_24958);
or UO_1457 (O_1457,N_29446,N_24819);
and UO_1458 (O_1458,N_28677,N_25040);
xor UO_1459 (O_1459,N_25472,N_28550);
or UO_1460 (O_1460,N_25211,N_28376);
and UO_1461 (O_1461,N_25923,N_24778);
xor UO_1462 (O_1462,N_29854,N_24151);
or UO_1463 (O_1463,N_29711,N_27064);
and UO_1464 (O_1464,N_24928,N_27680);
nand UO_1465 (O_1465,N_27888,N_28036);
nor UO_1466 (O_1466,N_29850,N_26532);
nor UO_1467 (O_1467,N_27986,N_29821);
nand UO_1468 (O_1468,N_29244,N_26756);
and UO_1469 (O_1469,N_28165,N_25570);
and UO_1470 (O_1470,N_26112,N_28287);
nor UO_1471 (O_1471,N_28251,N_27084);
or UO_1472 (O_1472,N_26784,N_28433);
or UO_1473 (O_1473,N_24716,N_27233);
xnor UO_1474 (O_1474,N_25433,N_24456);
or UO_1475 (O_1475,N_29061,N_28894);
and UO_1476 (O_1476,N_27706,N_27794);
or UO_1477 (O_1477,N_24347,N_24475);
and UO_1478 (O_1478,N_24754,N_24513);
and UO_1479 (O_1479,N_28285,N_27393);
nor UO_1480 (O_1480,N_25882,N_24270);
xor UO_1481 (O_1481,N_24550,N_26681);
and UO_1482 (O_1482,N_28535,N_26749);
or UO_1483 (O_1483,N_29812,N_29026);
xnor UO_1484 (O_1484,N_28965,N_27649);
xor UO_1485 (O_1485,N_25876,N_26990);
and UO_1486 (O_1486,N_26358,N_26898);
xnor UO_1487 (O_1487,N_26590,N_28351);
and UO_1488 (O_1488,N_29965,N_28273);
or UO_1489 (O_1489,N_25884,N_28967);
nor UO_1490 (O_1490,N_25993,N_27567);
nand UO_1491 (O_1491,N_26475,N_28270);
and UO_1492 (O_1492,N_27200,N_25811);
nand UO_1493 (O_1493,N_27744,N_28923);
nand UO_1494 (O_1494,N_27235,N_26935);
and UO_1495 (O_1495,N_26296,N_28519);
nor UO_1496 (O_1496,N_24974,N_27038);
nand UO_1497 (O_1497,N_28193,N_29094);
and UO_1498 (O_1498,N_28167,N_29105);
or UO_1499 (O_1499,N_27793,N_24789);
and UO_1500 (O_1500,N_26216,N_24341);
or UO_1501 (O_1501,N_29350,N_24844);
nor UO_1502 (O_1502,N_27277,N_24961);
xor UO_1503 (O_1503,N_24811,N_25982);
and UO_1504 (O_1504,N_24240,N_29428);
nand UO_1505 (O_1505,N_28164,N_24606);
xnor UO_1506 (O_1506,N_29671,N_27596);
and UO_1507 (O_1507,N_27228,N_24501);
and UO_1508 (O_1508,N_28904,N_25258);
nand UO_1509 (O_1509,N_24523,N_28901);
and UO_1510 (O_1510,N_29055,N_28053);
nor UO_1511 (O_1511,N_25431,N_24736);
or UO_1512 (O_1512,N_27711,N_27085);
or UO_1513 (O_1513,N_26298,N_28530);
nor UO_1514 (O_1514,N_28632,N_28829);
and UO_1515 (O_1515,N_28132,N_25488);
and UO_1516 (O_1516,N_26755,N_26907);
xor UO_1517 (O_1517,N_24609,N_26757);
or UO_1518 (O_1518,N_27377,N_25971);
xnor UO_1519 (O_1519,N_25314,N_24593);
and UO_1520 (O_1520,N_29885,N_28244);
and UO_1521 (O_1521,N_25674,N_25111);
or UO_1522 (O_1522,N_26579,N_24915);
nand UO_1523 (O_1523,N_25248,N_29355);
and UO_1524 (O_1524,N_28767,N_29734);
and UO_1525 (O_1525,N_26023,N_28444);
or UO_1526 (O_1526,N_27147,N_27034);
or UO_1527 (O_1527,N_29998,N_26920);
xor UO_1528 (O_1528,N_27570,N_29386);
xnor UO_1529 (O_1529,N_29157,N_26808);
nor UO_1530 (O_1530,N_27433,N_27598);
and UO_1531 (O_1531,N_24860,N_25521);
or UO_1532 (O_1532,N_29692,N_27642);
nor UO_1533 (O_1533,N_26551,N_29596);
and UO_1534 (O_1534,N_25561,N_29467);
xnor UO_1535 (O_1535,N_28022,N_27043);
and UO_1536 (O_1536,N_27989,N_25022);
nor UO_1537 (O_1537,N_25711,N_24805);
and UO_1538 (O_1538,N_27347,N_26044);
and UO_1539 (O_1539,N_27422,N_25984);
xor UO_1540 (O_1540,N_27974,N_27165);
xnor UO_1541 (O_1541,N_24879,N_25201);
or UO_1542 (O_1542,N_25685,N_27355);
nor UO_1543 (O_1543,N_26516,N_29970);
nor UO_1544 (O_1544,N_26315,N_27327);
and UO_1545 (O_1545,N_25781,N_25790);
and UO_1546 (O_1546,N_29819,N_24371);
xnor UO_1547 (O_1547,N_29573,N_28930);
nor UO_1548 (O_1548,N_25963,N_27186);
xnor UO_1549 (O_1549,N_26553,N_28708);
or UO_1550 (O_1550,N_24037,N_27196);
or UO_1551 (O_1551,N_27270,N_29440);
nor UO_1552 (O_1552,N_29531,N_27665);
and UO_1553 (O_1553,N_29764,N_26150);
nor UO_1554 (O_1554,N_29076,N_24034);
nor UO_1555 (O_1555,N_29472,N_29174);
nor UO_1556 (O_1556,N_24933,N_29079);
nand UO_1557 (O_1557,N_25943,N_25804);
nand UO_1558 (O_1558,N_26203,N_27325);
xor UO_1559 (O_1559,N_25950,N_28368);
or UO_1560 (O_1560,N_27801,N_25623);
and UO_1561 (O_1561,N_25513,N_29653);
xnor UO_1562 (O_1562,N_25171,N_24002);
and UO_1563 (O_1563,N_26895,N_27750);
xnor UO_1564 (O_1564,N_26555,N_28826);
and UO_1565 (O_1565,N_26760,N_27315);
nor UO_1566 (O_1566,N_28061,N_28587);
nor UO_1567 (O_1567,N_26262,N_27495);
xnor UO_1568 (O_1568,N_27071,N_25351);
and UO_1569 (O_1569,N_26347,N_28372);
nor UO_1570 (O_1570,N_29499,N_25839);
or UO_1571 (O_1571,N_27866,N_29409);
or UO_1572 (O_1572,N_25596,N_24468);
and UO_1573 (O_1573,N_24596,N_27951);
or UO_1574 (O_1574,N_28660,N_28928);
or UO_1575 (O_1575,N_28183,N_28981);
nor UO_1576 (O_1576,N_26288,N_24115);
and UO_1577 (O_1577,N_28098,N_28295);
or UO_1578 (O_1578,N_26228,N_24510);
or UO_1579 (O_1579,N_28549,N_29223);
or UO_1580 (O_1580,N_27443,N_26411);
or UO_1581 (O_1581,N_29618,N_28303);
or UO_1582 (O_1582,N_28235,N_26460);
or UO_1583 (O_1583,N_27312,N_24124);
and UO_1584 (O_1584,N_28682,N_28490);
or UO_1585 (O_1585,N_25128,N_24779);
or UO_1586 (O_1586,N_28258,N_25739);
and UO_1587 (O_1587,N_28347,N_25162);
xnor UO_1588 (O_1588,N_26777,N_24558);
nand UO_1589 (O_1589,N_27579,N_28706);
or UO_1590 (O_1590,N_25892,N_28203);
or UO_1591 (O_1591,N_28832,N_25369);
or UO_1592 (O_1592,N_28992,N_28401);
nand UO_1593 (O_1593,N_28785,N_28409);
nand UO_1594 (O_1594,N_29453,N_24841);
nor UO_1595 (O_1595,N_26879,N_24910);
or UO_1596 (O_1596,N_28071,N_28200);
or UO_1597 (O_1597,N_24344,N_27175);
and UO_1598 (O_1598,N_24070,N_28926);
and UO_1599 (O_1599,N_29894,N_28711);
and UO_1600 (O_1600,N_27630,N_27716);
nand UO_1601 (O_1601,N_24927,N_28227);
or UO_1602 (O_1602,N_24842,N_25028);
or UO_1603 (O_1603,N_29646,N_26089);
or UO_1604 (O_1604,N_25964,N_24717);
or UO_1605 (O_1605,N_27148,N_25715);
nor UO_1606 (O_1606,N_27019,N_25066);
or UO_1607 (O_1607,N_26437,N_26075);
xor UO_1608 (O_1608,N_27290,N_24645);
and UO_1609 (O_1609,N_25644,N_25338);
and UO_1610 (O_1610,N_26444,N_24633);
and UO_1611 (O_1611,N_28663,N_29016);
or UO_1612 (O_1612,N_27740,N_27261);
nor UO_1613 (O_1613,N_27150,N_27534);
nand UO_1614 (O_1614,N_26722,N_24007);
nor UO_1615 (O_1615,N_25252,N_27835);
nand UO_1616 (O_1616,N_25146,N_26533);
or UO_1617 (O_1617,N_24642,N_28117);
and UO_1618 (O_1618,N_27170,N_27542);
xnor UO_1619 (O_1619,N_27544,N_28466);
xnor UO_1620 (O_1620,N_25118,N_27966);
nand UO_1621 (O_1621,N_26255,N_29864);
and UO_1622 (O_1622,N_24994,N_25987);
and UO_1623 (O_1623,N_25321,N_29959);
nor UO_1624 (O_1624,N_26972,N_28986);
nand UO_1625 (O_1625,N_24104,N_28863);
or UO_1626 (O_1626,N_26732,N_28425);
or UO_1627 (O_1627,N_24381,N_27030);
and UO_1628 (O_1628,N_27751,N_25630);
nor UO_1629 (O_1629,N_29179,N_24935);
or UO_1630 (O_1630,N_26199,N_28847);
or UO_1631 (O_1631,N_26544,N_25642);
nor UO_1632 (O_1632,N_27436,N_25643);
or UO_1633 (O_1633,N_26964,N_29272);
and UO_1634 (O_1634,N_28219,N_28949);
nor UO_1635 (O_1635,N_29823,N_26456);
nand UO_1636 (O_1636,N_29868,N_28021);
xnor UO_1637 (O_1637,N_29188,N_25752);
nand UO_1638 (O_1638,N_29977,N_27036);
and UO_1639 (O_1639,N_28781,N_26680);
and UO_1640 (O_1640,N_26951,N_29023);
nand UO_1641 (O_1641,N_27773,N_29038);
or UO_1642 (O_1642,N_27893,N_26606);
nor UO_1643 (O_1643,N_24951,N_24957);
nor UO_1644 (O_1644,N_28718,N_25771);
and UO_1645 (O_1645,N_29871,N_27012);
or UO_1646 (O_1646,N_28077,N_29552);
xnor UO_1647 (O_1647,N_25447,N_24202);
or UO_1648 (O_1648,N_29087,N_26139);
nand UO_1649 (O_1649,N_25895,N_26066);
or UO_1650 (O_1650,N_26407,N_29750);
or UO_1651 (O_1651,N_29891,N_25945);
and UO_1652 (O_1652,N_26626,N_27435);
xnor UO_1653 (O_1653,N_26126,N_24771);
nor UO_1654 (O_1654,N_29127,N_26048);
xnor UO_1655 (O_1655,N_29733,N_29323);
nor UO_1656 (O_1656,N_27294,N_27118);
nand UO_1657 (O_1657,N_25495,N_27999);
or UO_1658 (O_1658,N_24469,N_25508);
and UO_1659 (O_1659,N_28559,N_28576);
nand UO_1660 (O_1660,N_29036,N_24911);
xor UO_1661 (O_1661,N_26457,N_24022);
or UO_1662 (O_1662,N_27834,N_28727);
nor UO_1663 (O_1663,N_24890,N_29404);
or UO_1664 (O_1664,N_24164,N_28501);
xnor UO_1665 (O_1665,N_26938,N_28600);
xor UO_1666 (O_1666,N_26260,N_28385);
nand UO_1667 (O_1667,N_25047,N_26868);
nor UO_1668 (O_1668,N_25240,N_27628);
and UO_1669 (O_1669,N_27476,N_27822);
xnor UO_1670 (O_1670,N_29494,N_26878);
nand UO_1671 (O_1671,N_28524,N_27937);
nand UO_1672 (O_1672,N_24872,N_24891);
or UO_1673 (O_1673,N_27173,N_29834);
nand UO_1674 (O_1674,N_26436,N_29441);
or UO_1675 (O_1675,N_29792,N_24551);
and UO_1676 (O_1676,N_29663,N_24415);
or UO_1677 (O_1677,N_27255,N_28243);
nand UO_1678 (O_1678,N_28469,N_28446);
nor UO_1679 (O_1679,N_26616,N_28515);
nor UO_1680 (O_1680,N_28284,N_25264);
nand UO_1681 (O_1681,N_27952,N_28006);
nor UO_1682 (O_1682,N_25308,N_28325);
nand UO_1683 (O_1683,N_25523,N_25191);
and UO_1684 (O_1684,N_24914,N_24163);
or UO_1685 (O_1685,N_24054,N_26022);
or UO_1686 (O_1686,N_29743,N_28134);
nor UO_1687 (O_1687,N_25176,N_26092);
nand UO_1688 (O_1688,N_26090,N_25794);
and UO_1689 (O_1689,N_29425,N_24200);
nor UO_1690 (O_1690,N_28144,N_26412);
nand UO_1691 (O_1691,N_28777,N_24813);
and UO_1692 (O_1692,N_26024,N_25808);
and UO_1693 (O_1693,N_28033,N_29886);
and UO_1694 (O_1694,N_25638,N_27585);
nand UO_1695 (O_1695,N_27040,N_29563);
and UO_1696 (O_1696,N_27514,N_25253);
and UO_1697 (O_1697,N_25041,N_25985);
and UO_1698 (O_1698,N_24316,N_28782);
and UO_1699 (O_1699,N_25202,N_29151);
nor UO_1700 (O_1700,N_26650,N_26896);
or UO_1701 (O_1701,N_27321,N_25052);
nand UO_1702 (O_1702,N_26634,N_29703);
nor UO_1703 (O_1703,N_27140,N_27973);
and UO_1704 (O_1704,N_29060,N_29304);
or UO_1705 (O_1705,N_25953,N_24195);
and UO_1706 (O_1706,N_29309,N_24810);
nor UO_1707 (O_1707,N_27802,N_27890);
and UO_1708 (O_1708,N_26742,N_26813);
nand UO_1709 (O_1709,N_24850,N_24756);
or UO_1710 (O_1710,N_25941,N_27927);
nand UO_1711 (O_1711,N_29485,N_24187);
or UO_1712 (O_1712,N_29766,N_26191);
xnor UO_1713 (O_1713,N_26981,N_26758);
or UO_1714 (O_1714,N_29654,N_25814);
nand UO_1715 (O_1715,N_29412,N_24356);
and UO_1716 (O_1716,N_28120,N_28562);
and UO_1717 (O_1717,N_29538,N_28592);
nor UO_1718 (O_1718,N_27636,N_24263);
nand UO_1719 (O_1719,N_26329,N_28416);
xor UO_1720 (O_1720,N_24275,N_27394);
xnor UO_1721 (O_1721,N_26063,N_27069);
nor UO_1722 (O_1722,N_24715,N_24189);
and UO_1723 (O_1723,N_28190,N_24210);
and UO_1724 (O_1724,N_29138,N_24390);
xor UO_1725 (O_1725,N_29044,N_27376);
nand UO_1726 (O_1726,N_29333,N_26301);
xnor UO_1727 (O_1727,N_28452,N_27087);
xor UO_1728 (O_1728,N_29729,N_24206);
nor UO_1729 (O_1729,N_25584,N_25267);
nand UO_1730 (O_1730,N_25610,N_24699);
or UO_1731 (O_1731,N_29233,N_27225);
nand UO_1732 (O_1732,N_24975,N_28774);
xnor UO_1733 (O_1733,N_26842,N_25441);
xnor UO_1734 (O_1734,N_29343,N_26409);
nor UO_1735 (O_1735,N_27441,N_25545);
nor UO_1736 (O_1736,N_27419,N_26035);
nor UO_1737 (O_1737,N_28494,N_27840);
and UO_1738 (O_1738,N_24035,N_29064);
nand UO_1739 (O_1739,N_24517,N_27098);
or UO_1740 (O_1740,N_25935,N_29104);
nor UO_1741 (O_1741,N_29751,N_24223);
or UO_1742 (O_1742,N_25944,N_26148);
xnor UO_1743 (O_1743,N_25818,N_26467);
xor UO_1744 (O_1744,N_28599,N_26489);
nor UO_1745 (O_1745,N_29236,N_27696);
nand UO_1746 (O_1746,N_26943,N_27826);
nor UO_1747 (O_1747,N_28824,N_25058);
or UO_1748 (O_1748,N_29687,N_29031);
or UO_1749 (O_1749,N_27268,N_27601);
nand UO_1750 (O_1750,N_29604,N_25697);
xor UO_1751 (O_1751,N_24784,N_27629);
nor UO_1752 (O_1752,N_29110,N_29649);
nor UO_1753 (O_1753,N_25342,N_25919);
xnor UO_1754 (O_1754,N_24425,N_28133);
xor UO_1755 (O_1755,N_29669,N_28666);
or UO_1756 (O_1756,N_29423,N_24521);
or UO_1757 (O_1757,N_28057,N_25170);
or UO_1758 (O_1758,N_26081,N_24346);
nand UO_1759 (O_1759,N_24992,N_26061);
nand UO_1760 (O_1760,N_29363,N_25563);
nand UO_1761 (O_1761,N_24463,N_27110);
and UO_1762 (O_1762,N_28843,N_27867);
xnor UO_1763 (O_1763,N_26252,N_24310);
or UO_1764 (O_1764,N_26267,N_28875);
and UO_1765 (O_1765,N_24432,N_26186);
and UO_1766 (O_1766,N_28434,N_26446);
and UO_1767 (O_1767,N_25900,N_29514);
and UO_1768 (O_1768,N_27958,N_27185);
or UO_1769 (O_1769,N_26655,N_25948);
and UO_1770 (O_1770,N_26271,N_26306);
and UO_1771 (O_1771,N_29131,N_29261);
nor UO_1772 (O_1772,N_26638,N_28131);
or UO_1773 (O_1773,N_27532,N_26137);
or UO_1774 (O_1774,N_26259,N_28978);
xor UO_1775 (O_1775,N_28637,N_26572);
or UO_1776 (O_1776,N_25698,N_27991);
xnor UO_1777 (O_1777,N_28362,N_24331);
nor UO_1778 (O_1778,N_29280,N_26161);
nand UO_1779 (O_1779,N_29755,N_26791);
nor UO_1780 (O_1780,N_28895,N_27006);
nor UO_1781 (O_1781,N_25991,N_29799);
xor UO_1782 (O_1782,N_26218,N_27417);
nand UO_1783 (O_1783,N_28027,N_25440);
xor UO_1784 (O_1784,N_24049,N_27073);
nand UO_1785 (O_1785,N_29782,N_29089);
nand UO_1786 (O_1786,N_25849,N_24695);
xor UO_1787 (O_1787,N_24815,N_27921);
and UO_1788 (O_1788,N_29546,N_28973);
or UO_1789 (O_1789,N_27155,N_29595);
nor UO_1790 (O_1790,N_24637,N_24604);
and UO_1791 (O_1791,N_27104,N_27641);
or UO_1792 (O_1792,N_29365,N_24735);
or UO_1793 (O_1793,N_24083,N_26077);
nor UO_1794 (O_1794,N_28532,N_24665);
or UO_1795 (O_1795,N_29651,N_28584);
nand UO_1796 (O_1796,N_26047,N_25608);
nand UO_1797 (O_1797,N_27605,N_27344);
xnor UO_1798 (O_1798,N_28480,N_26085);
nor UO_1799 (O_1799,N_25334,N_25409);
xor UO_1800 (O_1800,N_27526,N_24659);
xor UO_1801 (O_1801,N_28441,N_24904);
nand UO_1802 (O_1802,N_29212,N_28692);
xor UO_1803 (O_1803,N_26086,N_27632);
and UO_1804 (O_1804,N_28807,N_25766);
nor UO_1805 (O_1805,N_29198,N_24562);
and UO_1806 (O_1806,N_24800,N_29791);
nor UO_1807 (O_1807,N_28716,N_25934);
nor UO_1808 (O_1808,N_29717,N_27320);
nand UO_1809 (O_1809,N_25646,N_27764);
nor UO_1810 (O_1810,N_25014,N_25087);
xnor UO_1811 (O_1811,N_28247,N_25285);
nand UO_1812 (O_1812,N_26053,N_26417);
nand UO_1813 (O_1813,N_28607,N_24327);
and UO_1814 (O_1814,N_24233,N_26997);
or UO_1815 (O_1815,N_25080,N_24718);
and UO_1816 (O_1816,N_29257,N_28328);
xnor UO_1817 (O_1817,N_24787,N_27243);
nand UO_1818 (O_1818,N_29082,N_27487);
nor UO_1819 (O_1819,N_28977,N_25867);
nand UO_1820 (O_1820,N_27134,N_29683);
nor UO_1821 (O_1821,N_24916,N_29024);
nor UO_1822 (O_1822,N_29844,N_25592);
nand UO_1823 (O_1823,N_26326,N_27340);
or UO_1824 (O_1824,N_26487,N_25262);
nor UO_1825 (O_1825,N_25992,N_27331);
nor UO_1826 (O_1826,N_24602,N_26787);
and UO_1827 (O_1827,N_24373,N_24631);
and UO_1828 (O_1828,N_26423,N_25961);
or UO_1829 (O_1829,N_25446,N_27796);
xnor UO_1830 (O_1830,N_29694,N_26697);
and UO_1831 (O_1831,N_26294,N_25886);
or UO_1832 (O_1832,N_24362,N_24697);
nor UO_1833 (O_1833,N_24291,N_28963);
nor UO_1834 (O_1834,N_26998,N_28546);
nor UO_1835 (O_1835,N_27774,N_26779);
or UO_1836 (O_1836,N_29685,N_24905);
or UO_1837 (O_1837,N_29322,N_28784);
xnor UO_1838 (O_1838,N_27102,N_25777);
or UO_1839 (O_1839,N_24473,N_27451);
nand UO_1840 (O_1840,N_24312,N_29438);
nand UO_1841 (O_1841,N_24692,N_29985);
xor UO_1842 (O_1842,N_25348,N_26528);
and UO_1843 (O_1843,N_25072,N_29814);
nand UO_1844 (O_1844,N_28116,N_28911);
nand UO_1845 (O_1845,N_26101,N_27777);
nand UO_1846 (O_1846,N_28686,N_25129);
or UO_1847 (O_1847,N_28207,N_25686);
and UO_1848 (O_1848,N_25986,N_26314);
nor UO_1849 (O_1849,N_26811,N_29784);
nor UO_1850 (O_1850,N_27671,N_26929);
and UO_1851 (O_1851,N_28298,N_29722);
or UO_1852 (O_1852,N_24936,N_24048);
xnor UO_1853 (O_1853,N_27245,N_28959);
xor UO_1854 (O_1854,N_25672,N_26646);
nor UO_1855 (O_1855,N_25388,N_29732);
and UO_1856 (O_1856,N_29933,N_29788);
xnor UO_1857 (O_1857,N_24376,N_28941);
or UO_1858 (O_1858,N_27300,N_24998);
nand UO_1859 (O_1859,N_29938,N_28947);
xnor UO_1860 (O_1860,N_27303,N_24710);
nand UO_1861 (O_1861,N_25620,N_28917);
nor UO_1862 (O_1862,N_25881,N_29934);
or UO_1863 (O_1863,N_29861,N_29191);
nand UO_1864 (O_1864,N_24441,N_24114);
or UO_1865 (O_1865,N_28055,N_27365);
nand UO_1866 (O_1866,N_24068,N_28596);
nor UO_1867 (O_1867,N_26802,N_29120);
xnor UO_1868 (O_1868,N_26430,N_29253);
xor UO_1869 (O_1869,N_26144,N_26607);
nand UO_1870 (O_1870,N_25429,N_26602);
nand UO_1871 (O_1871,N_26620,N_26291);
or UO_1872 (O_1872,N_25085,N_27749);
nand UO_1873 (O_1873,N_25151,N_28249);
nor UO_1874 (O_1874,N_27249,N_25714);
or UO_1875 (O_1875,N_28871,N_29206);
nand UO_1876 (O_1876,N_28626,N_25363);
nor UO_1877 (O_1877,N_24378,N_29374);
xnor UO_1878 (O_1878,N_26610,N_24708);
xor UO_1879 (O_1879,N_24973,N_28166);
and UO_1880 (O_1880,N_24271,N_29967);
and UO_1881 (O_1881,N_28670,N_27715);
nand UO_1882 (O_1882,N_26605,N_26937);
xnor UO_1883 (O_1883,N_28657,N_26786);
xor UO_1884 (O_1884,N_26930,N_24152);
or UO_1885 (O_1885,N_25833,N_27968);
xnor UO_1886 (O_1886,N_24315,N_24908);
xnor UO_1887 (O_1887,N_25837,N_26155);
xnor UO_1888 (O_1888,N_29701,N_27916);
and UO_1889 (O_1889,N_24966,N_24806);
xor UO_1890 (O_1890,N_24295,N_24531);
xnor UO_1891 (O_1891,N_24749,N_27424);
nor UO_1892 (O_1892,N_28307,N_25091);
or UO_1893 (O_1893,N_26661,N_27824);
nand UO_1894 (O_1894,N_27620,N_24621);
or UO_1895 (O_1895,N_27724,N_28349);
and UO_1896 (O_1896,N_26377,N_26372);
and UO_1897 (O_1897,N_28544,N_26950);
xnor UO_1898 (O_1898,N_26042,N_26479);
or UO_1899 (O_1899,N_26172,N_29000);
xnor UO_1900 (O_1900,N_24770,N_28537);
nand UO_1901 (O_1901,N_24824,N_26825);
xnor UO_1902 (O_1902,N_25095,N_25994);
nand UO_1903 (O_1903,N_24929,N_24846);
or UO_1904 (O_1904,N_26194,N_27902);
xor UO_1905 (O_1905,N_25453,N_27166);
xnor UO_1906 (O_1906,N_28379,N_25795);
nand UO_1907 (O_1907,N_28301,N_27851);
xor UO_1908 (O_1908,N_24518,N_27829);
xor UO_1909 (O_1909,N_27350,N_29758);
xor UO_1910 (O_1910,N_26438,N_26921);
xor UO_1911 (O_1911,N_27594,N_26490);
and UO_1912 (O_1912,N_26723,N_25537);
and UO_1913 (O_1913,N_29930,N_24428);
xnor UO_1914 (O_1914,N_26104,N_25861);
nand UO_1915 (O_1915,N_29150,N_28976);
and UO_1916 (O_1916,N_25649,N_25241);
and UO_1917 (O_1917,N_25403,N_25510);
nand UO_1918 (O_1918,N_28020,N_27363);
or UO_1919 (O_1919,N_27472,N_29039);
xnor UO_1920 (O_1920,N_25712,N_29973);
or UO_1921 (O_1921,N_25155,N_28937);
xor UO_1922 (O_1922,N_24753,N_24196);
nand UO_1923 (O_1923,N_24245,N_28489);
or UO_1924 (O_1924,N_28139,N_29027);
or UO_1925 (O_1925,N_25678,N_24234);
or UO_1926 (O_1926,N_28260,N_28130);
nand UO_1927 (O_1927,N_27885,N_26376);
nor UO_1928 (O_1928,N_29069,N_29181);
or UO_1929 (O_1929,N_26870,N_27597);
nor UO_1930 (O_1930,N_25002,N_29068);
nor UO_1931 (O_1931,N_29097,N_29100);
or UO_1932 (O_1932,N_25001,N_27669);
xor UO_1933 (O_1933,N_29647,N_26763);
nand UO_1934 (O_1934,N_24476,N_29243);
nand UO_1935 (O_1935,N_26002,N_25103);
xnor UO_1936 (O_1936,N_27232,N_25997);
nor UO_1937 (O_1937,N_25692,N_25872);
nor UO_1938 (O_1938,N_25385,N_25152);
nand UO_1939 (O_1939,N_27896,N_24644);
nor UO_1940 (O_1940,N_29324,N_26864);
xor UO_1941 (O_1941,N_24989,N_29124);
nand UO_1942 (O_1942,N_24938,N_24617);
nor UO_1943 (O_1943,N_27210,N_26443);
xnor UO_1944 (O_1944,N_29009,N_27805);
xnor UO_1945 (O_1945,N_27077,N_29610);
xor UO_1946 (O_1946,N_28536,N_24898);
and UO_1947 (O_1947,N_28859,N_25265);
or UO_1948 (O_1948,N_26253,N_25486);
and UO_1949 (O_1949,N_28714,N_28560);
and UO_1950 (O_1950,N_25588,N_27146);
or UO_1951 (O_1951,N_24431,N_24930);
nor UO_1952 (O_1952,N_24688,N_27768);
and UO_1953 (O_1953,N_24150,N_29677);
and UO_1954 (O_1954,N_25978,N_27306);
nor UO_1955 (O_1955,N_26624,N_28056);
xor UO_1956 (O_1956,N_26321,N_28269);
and UO_1957 (O_1957,N_25149,N_29081);
xnor UO_1958 (O_1958,N_28129,N_29969);
or UO_1959 (O_1959,N_26830,N_24706);
or UO_1960 (O_1960,N_29146,N_27237);
nand UO_1961 (O_1961,N_25025,N_26231);
xnor UO_1962 (O_1962,N_26168,N_24408);
xnor UO_1963 (O_1963,N_29185,N_24338);
nor UO_1964 (O_1964,N_25015,N_29710);
and UO_1965 (O_1965,N_25550,N_25576);
nor UO_1966 (O_1966,N_28185,N_28477);
and UO_1967 (O_1967,N_26946,N_26354);
nand UO_1968 (O_1968,N_26916,N_27135);
nor UO_1969 (O_1969,N_25755,N_24926);
or UO_1970 (O_1970,N_29881,N_25774);
xnor UO_1971 (O_1971,N_26180,N_24459);
xnor UO_1972 (O_1972,N_26302,N_24304);
and UO_1973 (O_1973,N_29979,N_29633);
or UO_1974 (O_1974,N_24352,N_24941);
nand UO_1975 (O_1975,N_24751,N_24888);
and UO_1976 (O_1976,N_24542,N_27522);
nand UO_1977 (O_1977,N_24110,N_24299);
nand UO_1978 (O_1978,N_24406,N_28126);
nor UO_1979 (O_1979,N_28754,N_24907);
xor UO_1980 (O_1980,N_26052,N_25086);
nand UO_1981 (O_1981,N_24117,N_26631);
nor UO_1982 (O_1982,N_26525,N_28927);
and UO_1983 (O_1983,N_25546,N_27944);
nor UO_1984 (O_1984,N_25410,N_24337);
or UO_1985 (O_1985,N_28415,N_29811);
nand UO_1986 (O_1986,N_26488,N_27329);
and UO_1987 (O_1987,N_25841,N_25744);
nand UO_1988 (O_1988,N_28242,N_28966);
xnor UO_1989 (O_1989,N_25492,N_24130);
nor UO_1990 (O_1990,N_28387,N_27683);
nor UO_1991 (O_1991,N_29239,N_29672);
nor UO_1992 (O_1992,N_24532,N_26803);
nor UO_1993 (O_1993,N_27539,N_25347);
nand UO_1994 (O_1994,N_25916,N_27343);
nor UO_1995 (O_1995,N_24302,N_29725);
nor UO_1996 (O_1996,N_28182,N_25442);
xor UO_1997 (O_1997,N_27278,N_26774);
or UO_1998 (O_1998,N_28726,N_24367);
or UO_1999 (O_1999,N_25768,N_28461);
or UO_2000 (O_2000,N_24690,N_26497);
and UO_2001 (O_2001,N_25829,N_24984);
or UO_2002 (O_2002,N_26281,N_24834);
and UO_2003 (O_2003,N_27707,N_29166);
or UO_2004 (O_2004,N_29091,N_29496);
nand UO_2005 (O_2005,N_27391,N_26911);
or UO_2006 (O_2006,N_27183,N_27797);
xnor UO_2007 (O_2007,N_27811,N_28361);
and UO_2008 (O_2008,N_24965,N_26303);
nor UO_2009 (O_2009,N_26969,N_25251);
and UO_2010 (O_2010,N_28775,N_27423);
xor UO_2011 (O_2011,N_28842,N_24004);
xnor UO_2012 (O_2012,N_26772,N_27842);
nor UO_2013 (O_2013,N_24685,N_25225);
xor UO_2014 (O_2014,N_29564,N_29176);
xor UO_2015 (O_2015,N_26918,N_28392);
nand UO_2016 (O_2016,N_24045,N_29518);
nor UO_2017 (O_2017,N_26210,N_28474);
or UO_2018 (O_2018,N_28030,N_24434);
nand UO_2019 (O_2019,N_26337,N_25068);
xor UO_2020 (O_2020,N_24662,N_27584);
or UO_2021 (O_2021,N_27491,N_28470);
nand UO_2022 (O_2022,N_27908,N_28180);
nand UO_2023 (O_2023,N_28140,N_26623);
xor UO_2024 (O_2024,N_25682,N_27681);
and UO_2025 (O_2025,N_24934,N_27250);
xor UO_2026 (O_2026,N_24121,N_26482);
and UO_2027 (O_2027,N_26603,N_25551);
nor UO_2028 (O_2028,N_28375,N_28246);
nand UO_2029 (O_2029,N_26788,N_28430);
nand UO_2030 (O_2030,N_28700,N_25724);
or UO_2031 (O_2031,N_24273,N_25968);
and UO_2032 (O_2032,N_26176,N_28858);
or UO_2033 (O_2033,N_28136,N_25878);
xnor UO_2034 (O_2034,N_25194,N_29085);
nor UO_2035 (O_2035,N_29707,N_24511);
nor UO_2036 (O_2036,N_25046,N_24298);
nand UO_2037 (O_2037,N_28783,N_24489);
or UO_2038 (O_2038,N_29650,N_25220);
nor UO_2039 (O_2039,N_29302,N_27554);
nand UO_2040 (O_2040,N_28602,N_26963);
nand UO_2041 (O_2041,N_26295,N_27372);
nor UO_2042 (O_2042,N_25666,N_26843);
nand UO_2043 (O_2043,N_28191,N_28792);
or UO_2044 (O_2044,N_29308,N_24297);
nor UO_2045 (O_2045,N_25499,N_26270);
and UO_2046 (O_2046,N_26491,N_27645);
nor UO_2047 (O_2047,N_27611,N_24440);
or UO_2048 (O_2048,N_27934,N_25233);
nand UO_2049 (O_2049,N_28377,N_25922);
nor UO_2050 (O_2050,N_24851,N_25007);
nor UO_2051 (O_2051,N_25464,N_24453);
nor UO_2052 (O_2052,N_27752,N_24833);
and UO_2053 (O_2053,N_28315,N_27264);
and UO_2054 (O_2054,N_27816,N_29096);
nor UO_2055 (O_2055,N_27153,N_24603);
nor UO_2056 (O_2056,N_27679,N_29160);
xor UO_2057 (O_2057,N_29569,N_27127);
nor UO_2058 (O_2058,N_26404,N_27015);
nand UO_2059 (O_2059,N_27571,N_28009);
xnor UO_2060 (O_2060,N_28748,N_25386);
xor UO_2061 (O_2061,N_24723,N_28628);
xor UO_2062 (O_2062,N_29139,N_28048);
nand UO_2063 (O_2063,N_27215,N_27361);
and UO_2064 (O_2064,N_26957,N_29380);
or UO_2065 (O_2065,N_24549,N_27238);
and UO_2066 (O_2066,N_27396,N_28954);
nor UO_2067 (O_2067,N_26738,N_28520);
nand UO_2068 (O_2068,N_28953,N_29296);
xor UO_2069 (O_2069,N_25117,N_29282);
nand UO_2070 (O_2070,N_27328,N_26978);
and UO_2071 (O_2071,N_24407,N_24388);
xnor UO_2072 (O_2072,N_25224,N_25394);
nand UO_2073 (O_2073,N_29398,N_27078);
xnor UO_2074 (O_2074,N_24236,N_29501);
nand UO_2075 (O_2075,N_29577,N_26029);
or UO_2076 (O_2076,N_28612,N_29892);
nor UO_2077 (O_2077,N_26209,N_29695);
nor UO_2078 (O_2078,N_28342,N_28720);
xnor UO_2079 (O_2079,N_28915,N_28458);
and UO_2080 (O_2080,N_24792,N_25189);
xnor UO_2081 (O_2081,N_27438,N_25203);
nand UO_2082 (O_2082,N_24590,N_29554);
nor UO_2083 (O_2083,N_27405,N_25192);
or UO_2084 (O_2084,N_27781,N_29946);
xnor UO_2085 (O_2085,N_26604,N_25428);
xnor UO_2086 (O_2086,N_26272,N_26684);
and UO_2087 (O_2087,N_28442,N_29820);
xor UO_2088 (O_2088,N_28499,N_25364);
nor UO_2089 (O_2089,N_24980,N_29306);
and UO_2090 (O_2090,N_24038,N_26107);
nand UO_2091 (O_2091,N_27537,N_26465);
xnor UO_2092 (O_2092,N_29756,N_27489);
nand UO_2093 (O_2093,N_29526,N_26502);
nor UO_2094 (O_2094,N_25034,N_27471);
nand UO_2095 (O_2095,N_27430,N_25465);
nand UO_2096 (O_2096,N_26114,N_24821);
xnor UO_2097 (O_2097,N_25292,N_25966);
nand UO_2098 (O_2098,N_25816,N_25377);
nand UO_2099 (O_2099,N_28993,N_29193);
or UO_2100 (O_2100,N_25940,N_27655);
and UO_2101 (O_2101,N_29639,N_26128);
or UO_2102 (O_2102,N_29148,N_27248);
nand UO_2103 (O_2103,N_29062,N_24180);
or UO_2104 (O_2104,N_28543,N_26633);
nor UO_2105 (O_2105,N_29712,N_24284);
nor UO_2106 (O_2106,N_24116,N_26495);
or UO_2107 (O_2107,N_28395,N_27427);
and UO_2108 (O_2108,N_27947,N_25925);
or UO_2109 (O_2109,N_25595,N_26328);
and UO_2110 (O_2110,N_29402,N_24626);
or UO_2111 (O_2111,N_27699,N_25857);
and UO_2112 (O_2112,N_25355,N_25005);
and UO_2113 (O_2113,N_27297,N_24959);
and UO_2114 (O_2114,N_29645,N_28497);
and UO_2115 (O_2115,N_29383,N_28218);
and UO_2116 (O_2116,N_24895,N_27395);
and UO_2117 (O_2117,N_24218,N_27284);
xor UO_2118 (O_2118,N_24470,N_28516);
nand UO_2119 (O_2119,N_26994,N_27980);
and UO_2120 (O_2120,N_24313,N_26567);
nor UO_2121 (O_2121,N_28223,N_26565);
xor UO_2122 (O_2122,N_25562,N_25709);
xor UO_2123 (O_2123,N_29461,N_25614);
nand UO_2124 (O_2124,N_29481,N_27574);
nand UO_2125 (O_2125,N_26100,N_24553);
and UO_2126 (O_2126,N_28811,N_29619);
nor UO_2127 (O_2127,N_27447,N_27119);
nand UO_2128 (O_2128,N_27735,N_26141);
xnor UO_2129 (O_2129,N_26182,N_27008);
nand UO_2130 (O_2130,N_25498,N_25540);
xor UO_2131 (O_2131,N_28101,N_25885);
xnor UO_2132 (O_2132,N_25301,N_28308);
and UO_2133 (O_2133,N_29833,N_29520);
xnor UO_2134 (O_2134,N_25819,N_25109);
nand UO_2135 (O_2135,N_26390,N_29513);
or UO_2136 (O_2136,N_27499,N_25274);
nor UO_2137 (O_2137,N_25915,N_29403);
nand UO_2138 (O_2138,N_26597,N_26944);
or UO_2139 (O_2139,N_24608,N_27688);
or UO_2140 (O_2140,N_24021,N_28796);
and UO_2141 (O_2141,N_27308,N_26451);
xor UO_2142 (O_2142,N_28962,N_28776);
nor UO_2143 (O_2143,N_28293,N_27257);
xor UO_2144 (O_2144,N_27220,N_26125);
or UO_2145 (O_2145,N_25019,N_26120);
xnor UO_2146 (O_2146,N_24477,N_29976);
xor UO_2147 (O_2147,N_27637,N_27061);
nand UO_2148 (O_2148,N_29156,N_25003);
nor UO_2149 (O_2149,N_27302,N_26452);
xnor UO_2150 (O_2150,N_26336,N_24279);
nand UO_2151 (O_2151,N_27798,N_27323);
or UO_2152 (O_2152,N_29585,N_25983);
nand UO_2153 (O_2153,N_27388,N_25078);
nor UO_2154 (O_2154,N_25585,N_29248);
xor UO_2155 (O_2155,N_24444,N_28948);
nor UO_2156 (O_2156,N_24719,N_24414);
xnor UO_2157 (O_2157,N_26193,N_25098);
and UO_2158 (O_2158,N_27336,N_24265);
nor UO_2159 (O_2159,N_24601,N_24173);
xnor UO_2160 (O_2160,N_26370,N_26698);
xnor UO_2161 (O_2161,N_25305,N_24886);
or UO_2162 (O_2162,N_28173,N_27511);
and UO_2163 (O_2163,N_29863,N_29536);
nor UO_2164 (O_2164,N_26662,N_29442);
or UO_2165 (O_2165,N_27307,N_29611);
nand UO_2166 (O_2166,N_28630,N_29477);
xnor UO_2167 (O_2167,N_26985,N_28456);
and UO_2168 (O_2168,N_27552,N_28943);
xnor UO_2169 (O_2169,N_25463,N_25702);
and UO_2170 (O_2170,N_24923,N_28667);
and UO_2171 (O_2171,N_24409,N_28394);
nor UO_2172 (O_2172,N_26041,N_28802);
nand UO_2173 (O_2173,N_29584,N_25898);
or UO_2174 (O_2174,N_26201,N_24791);
and UO_2175 (O_2175,N_26648,N_29957);
xor UO_2176 (O_2176,N_27713,N_27703);
nand UO_2177 (O_2177,N_26027,N_25679);
xor UO_2178 (O_2178,N_29459,N_24970);
xor UO_2179 (O_2179,N_27092,N_29136);
or UO_2180 (O_2180,N_28889,N_27349);
nand UO_2181 (O_2181,N_24498,N_27319);
and UO_2182 (O_2182,N_25359,N_26094);
and UO_2183 (O_2183,N_25586,N_25397);
and UO_2184 (O_2184,N_28586,N_29354);
xor UO_2185 (O_2185,N_24064,N_26408);
xnor UO_2186 (O_2186,N_29980,N_27501);
or UO_2187 (O_2187,N_25746,N_28764);
and UO_2188 (O_2188,N_25617,N_29878);
nor UO_2189 (O_2189,N_25381,N_27555);
nor UO_2190 (O_2190,N_27464,N_28472);
xnor UO_2191 (O_2191,N_25912,N_26458);
nor UO_2192 (O_2192,N_25750,N_29858);
nand UO_2193 (O_2193,N_25190,N_27131);
nand UO_2194 (O_2194,N_24386,N_24702);
nand UO_2195 (O_2195,N_25719,N_24999);
or UO_2196 (O_2196,N_27837,N_27339);
nor UO_2197 (O_2197,N_29432,N_27265);
and UO_2198 (O_2198,N_27806,N_26587);
nor UO_2199 (O_2199,N_26517,N_27047);
and UO_2200 (O_2200,N_25470,N_28039);
or UO_2201 (O_2201,N_26660,N_27020);
or UO_2202 (O_2202,N_24758,N_24325);
nor UO_2203 (O_2203,N_29487,N_24098);
nor UO_2204 (O_2204,N_26091,N_26369);
nand UO_2205 (O_2205,N_29391,N_29902);
xnor UO_2206 (O_2206,N_29664,N_27358);
nor UO_2207 (O_2207,N_28215,N_25131);
nand UO_2208 (O_2208,N_28181,N_28478);
or UO_2209 (O_2209,N_28836,N_29196);
xnor UO_2210 (O_2210,N_25116,N_27849);
nor UO_2211 (O_2211,N_27839,N_29017);
and UO_2212 (O_2212,N_28035,N_27246);
xnor UO_2213 (O_2213,N_24976,N_28319);
and UO_2214 (O_2214,N_25242,N_29836);
and UO_2215 (O_2215,N_25716,N_29458);
or UO_2216 (O_2216,N_25183,N_27913);
nor UO_2217 (O_2217,N_29071,N_28152);
xnor UO_2218 (O_2218,N_25154,N_25140);
xnor UO_2219 (O_2219,N_28089,N_29483);
or UO_2220 (O_2220,N_29890,N_29415);
or UO_2221 (O_2221,N_28597,N_25197);
or UO_2222 (O_2222,N_24141,N_24008);
xor UO_2223 (O_2223,N_24687,N_28867);
nor UO_2224 (O_2224,N_27494,N_25421);
and UO_2225 (O_2225,N_29681,N_26673);
or UO_2226 (O_2226,N_29988,N_26584);
and UO_2227 (O_2227,N_25343,N_24525);
or UO_2228 (O_2228,N_27910,N_25064);
nor UO_2229 (O_2229,N_28818,N_24740);
and UO_2230 (O_2230,N_28713,N_25824);
nor UO_2231 (O_2231,N_28118,N_24282);
nand UO_2232 (O_2232,N_26526,N_24040);
nand UO_2233 (O_2233,N_24486,N_29362);
xor UO_2234 (O_2234,N_24627,N_28886);
nor UO_2235 (O_2235,N_25126,N_25732);
xnor UO_2236 (O_2236,N_24293,N_28940);
nand UO_2237 (O_2237,N_28837,N_26751);
nor UO_2238 (O_2238,N_25017,N_24725);
nor UO_2239 (O_2239,N_29339,N_28554);
or UO_2240 (O_2240,N_24874,N_29813);
xor UO_2241 (O_2241,N_27942,N_29956);
and UO_2242 (O_2242,N_25368,N_25965);
nor UO_2243 (O_2243,N_28371,N_24375);
nor UO_2244 (O_2244,N_24491,N_27938);
nand UO_2245 (O_2245,N_29971,N_27879);
nand UO_2246 (O_2246,N_28421,N_25748);
nor UO_2247 (O_2247,N_24639,N_26151);
or UO_2248 (O_2248,N_28495,N_26677);
xor UO_2249 (O_2249,N_25936,N_26876);
or UO_2250 (O_2250,N_28846,N_24241);
nor UO_2251 (O_2251,N_29314,N_29454);
and UO_2252 (O_2252,N_26367,N_24830);
and UO_2253 (O_2253,N_27844,N_25352);
nand UO_2254 (O_2254,N_29192,N_29594);
xor UO_2255 (O_2255,N_25891,N_27739);
nand UO_2256 (O_2256,N_28485,N_29340);
xor UO_2257 (O_2257,N_25278,N_27218);
nor UO_2258 (O_2258,N_24790,N_29211);
and UO_2259 (O_2259,N_29848,N_26841);
nor UO_2260 (O_2260,N_24149,N_27955);
nor UO_2261 (O_2261,N_24566,N_29693);
xor UO_2262 (O_2262,N_24055,N_26764);
nand UO_2263 (O_2263,N_28145,N_25522);
and UO_2264 (O_2264,N_28241,N_27461);
nand UO_2265 (O_2265,N_25946,N_24165);
nor UO_2266 (O_2266,N_25230,N_25607);
nor UO_2267 (O_2267,N_27870,N_25232);
and UO_2268 (O_2268,N_26236,N_25693);
and UO_2269 (O_2269,N_27156,N_26480);
nor UO_2270 (O_2270,N_28366,N_28979);
nand UO_2271 (O_2271,N_29292,N_25547);
xor UO_2272 (O_2272,N_29806,N_27827);
and UO_2273 (O_2273,N_24138,N_29222);
nand UO_2274 (O_2274,N_27935,N_29655);
nor UO_2275 (O_2275,N_28719,N_29444);
or UO_2276 (O_2276,N_25555,N_26797);
xor UO_2277 (O_2277,N_27189,N_27528);
xnor UO_2278 (O_2278,N_28916,N_24755);
nor UO_2279 (O_2279,N_25660,N_26308);
xnor UO_2280 (O_2280,N_27946,N_28872);
xor UO_2281 (O_2281,N_25044,N_26233);
nand UO_2282 (O_2282,N_24554,N_24393);
or UO_2283 (O_2283,N_26967,N_28593);
and UO_2284 (O_2284,N_26058,N_25645);
xnor UO_2285 (O_2285,N_26343,N_26783);
or UO_2286 (O_2286,N_27602,N_27712);
nand UO_2287 (O_2287,N_27137,N_28090);
nor UO_2288 (O_2288,N_27066,N_25067);
or UO_2289 (O_2289,N_28921,N_27252);
or UO_2290 (O_2290,N_28655,N_25722);
and UO_2291 (O_2291,N_27434,N_25825);
or UO_2292 (O_2292,N_26074,N_24745);
and UO_2293 (O_2293,N_26254,N_28710);
xor UO_2294 (O_2294,N_29195,N_27976);
xnor UO_2295 (O_2295,N_27931,N_26123);
nor UO_2296 (O_2296,N_26419,N_28100);
or UO_2297 (O_2297,N_28934,N_24258);
or UO_2298 (O_2298,N_28296,N_27843);
nand UO_2299 (O_2299,N_25754,N_27971);
nand UO_2300 (O_2300,N_29184,N_29254);
xor UO_2301 (O_2301,N_25506,N_29570);
or UO_2302 (O_2302,N_26305,N_28762);
nor UO_2303 (O_2303,N_24577,N_24435);
or UO_2304 (O_2304,N_28286,N_29049);
or UO_2305 (O_2305,N_27729,N_25681);
and UO_2306 (O_2306,N_28790,N_25625);
nand UO_2307 (O_2307,N_28650,N_25214);
nand UO_2308 (O_2308,N_24809,N_27769);
or UO_2309 (O_2309,N_27410,N_28924);
nor UO_2310 (O_2310,N_27623,N_28733);
xnor UO_2311 (O_2311,N_26731,N_29768);
nand UO_2312 (O_2312,N_25036,N_27274);
or UO_2313 (O_2313,N_24429,N_28179);
nand UO_2314 (O_2314,N_25480,N_25088);
and UO_2315 (O_2315,N_25168,N_28427);
nor UO_2316 (O_2316,N_26500,N_26563);
or UO_2317 (O_2317,N_27260,N_27045);
nor UO_2318 (O_2318,N_25097,N_29369);
nand UO_2319 (O_2319,N_26643,N_28388);
xnor UO_2320 (O_2320,N_27027,N_24354);
nand UO_2321 (O_2321,N_29537,N_29410);
and UO_2322 (O_2322,N_25311,N_24924);
or UO_2323 (O_2323,N_24492,N_28004);
or UO_2324 (O_2324,N_29034,N_25579);
nand UO_2325 (O_2325,N_25042,N_29621);
nand UO_2326 (O_2326,N_26374,N_25284);
or UO_2327 (O_2327,N_26378,N_29507);
and UO_2328 (O_2328,N_26032,N_28380);
and UO_2329 (O_2329,N_24071,N_27011);
xnor UO_2330 (O_2330,N_24653,N_27872);
and UO_2331 (O_2331,N_26221,N_29796);
nand UO_2332 (O_2332,N_24318,N_29285);
nand UO_2333 (O_2333,N_27875,N_26464);
nand UO_2334 (O_2334,N_24292,N_25127);
or UO_2335 (O_2335,N_25226,N_24159);
and UO_2336 (O_2336,N_27736,N_27258);
nor UO_2337 (O_2337,N_27108,N_28502);
nor UO_2338 (O_2338,N_27905,N_25583);
xnor UO_2339 (O_2339,N_24573,N_27608);
nor UO_2340 (O_2340,N_28841,N_29870);
nor UO_2341 (O_2341,N_24496,N_29905);
and UO_2342 (O_2342,N_27273,N_25680);
nand UO_2343 (O_2343,N_28747,N_27070);
nand UO_2344 (O_2344,N_24365,N_26368);
nand UO_2345 (O_2345,N_24788,N_29574);
and UO_2346 (O_2346,N_24379,N_24436);
or UO_2347 (O_2347,N_25559,N_24421);
or UO_2348 (O_2348,N_24102,N_26871);
and UO_2349 (O_2349,N_27741,N_25175);
nand UO_2350 (O_2350,N_29098,N_24112);
and UO_2351 (O_2351,N_24222,N_27010);
nand UO_2352 (O_2352,N_29986,N_27507);
nand UO_2353 (O_2353,N_24832,N_24912);
nand UO_2354 (O_2354,N_29617,N_24757);
and UO_2355 (O_2355,N_25167,N_25271);
xor UO_2356 (O_2356,N_26461,N_24364);
nand UO_2357 (O_2357,N_27990,N_24260);
or UO_2358 (O_2358,N_25887,N_25469);
or UO_2359 (O_2359,N_28311,N_25261);
xor UO_2360 (O_2360,N_29480,N_27901);
nand UO_2361 (O_2361,N_27005,N_29790);
nand UO_2362 (O_2362,N_26940,N_24497);
and UO_2363 (O_2363,N_27371,N_29731);
or UO_2364 (O_2364,N_27709,N_24901);
and UO_2365 (O_2365,N_24335,N_27457);
nor UO_2366 (O_2366,N_26335,N_24057);
and UO_2367 (O_2367,N_26705,N_25439);
or UO_2368 (O_2368,N_27725,N_28102);
or UO_2369 (O_2369,N_26115,N_28473);
or UO_2370 (O_2370,N_28991,N_26922);
nand UO_2371 (O_2371,N_24825,N_27348);
nor UO_2372 (O_2372,N_28868,N_24063);
nand UO_2373 (O_2373,N_24494,N_25383);
xnor UO_2374 (O_2374,N_28318,N_29030);
and UO_2375 (O_2375,N_27723,N_26548);
and UO_2376 (O_2376,N_28370,N_26403);
nand UO_2377 (O_2377,N_25554,N_27614);
or UO_2378 (O_2378,N_28168,N_27090);
nand UO_2379 (O_2379,N_26313,N_27402);
and UO_2380 (O_2380,N_29818,N_24056);
xor UO_2381 (O_2381,N_29464,N_28403);
nor UO_2382 (O_2382,N_25639,N_29059);
xnor UO_2383 (O_2383,N_26761,N_26198);
nand UO_2384 (O_2384,N_24405,N_25641);
xor UO_2385 (O_2385,N_25906,N_25860);
and UO_2386 (O_2386,N_28496,N_24635);
nor UO_2387 (O_2387,N_26819,N_29337);
and UO_2388 (O_2388,N_27738,N_27025);
nor UO_2389 (O_2389,N_27151,N_25552);
xor UO_2390 (O_2390,N_29942,N_29214);
or UO_2391 (O_2391,N_25989,N_24894);
nor UO_2392 (O_2392,N_24186,N_29738);
nand UO_2393 (O_2393,N_24207,N_26735);
nor UO_2394 (O_2394,N_28253,N_27838);
nor UO_2395 (O_2395,N_24345,N_26806);
or UO_2396 (O_2396,N_29187,N_26320);
nand UO_2397 (O_2397,N_27720,N_27114);
nand UO_2398 (O_2398,N_25591,N_27481);
or UO_2399 (O_2399,N_28575,N_29298);
and UO_2400 (O_2400,N_28194,N_26608);
nand UO_2401 (O_2401,N_25661,N_25325);
nor UO_2402 (O_2402,N_24728,N_29035);
xnor UO_2403 (O_2403,N_28763,N_27627);
nand UO_2404 (O_2404,N_27581,N_24391);
xnor UO_2405 (O_2405,N_29597,N_27449);
xnor UO_2406 (O_2406,N_25669,N_29421);
nand UO_2407 (O_2407,N_25601,N_25874);
nor UO_2408 (O_2408,N_24276,N_27123);
xor UO_2409 (O_2409,N_25406,N_29328);
and UO_2410 (O_2410,N_29534,N_28143);
nor UO_2411 (O_2411,N_26005,N_25070);
nor UO_2412 (O_2412,N_28695,N_28627);
nand UO_2413 (O_2413,N_28891,N_24069);
and UO_2414 (O_2414,N_29348,N_28799);
nor UO_2415 (O_2415,N_29837,N_29721);
xor UO_2416 (O_2416,N_29640,N_28008);
nand UO_2417 (O_2417,N_28804,N_24504);
and UO_2418 (O_2418,N_28957,N_28449);
nor UO_2419 (O_2419,N_29018,N_28459);
xor UO_2420 (O_2420,N_24918,N_24303);
nor UO_2421 (O_2421,N_29824,N_24474);
and UO_2422 (O_2422,N_29145,N_28533);
or UO_2423 (O_2423,N_26543,N_27812);
or UO_2424 (O_2424,N_27756,N_29705);
nand UO_2425 (O_2425,N_29396,N_25424);
and UO_2426 (O_2426,N_24101,N_28618);
nand UO_2427 (O_2427,N_27521,N_27779);
and UO_2428 (O_2428,N_26863,N_29745);
xnor UO_2429 (O_2429,N_24960,N_26316);
nor UO_2430 (O_2430,N_29263,N_24855);
nand UO_2431 (O_2431,N_26917,N_29505);
nand UO_2432 (O_2432,N_28294,N_26363);
or UO_2433 (O_2433,N_29277,N_25573);
xor UO_2434 (O_2434,N_24235,N_25897);
and UO_2435 (O_2435,N_29327,N_24691);
xnor UO_2436 (O_2436,N_26097,N_24986);
or UO_2437 (O_2437,N_28302,N_27317);
nor UO_2438 (O_2438,N_26060,N_26096);
and UO_2439 (O_2439,N_26670,N_25763);
nand UO_2440 (O_2440,N_26592,N_25929);
xor UO_2441 (O_2441,N_26154,N_27644);
and UO_2442 (O_2442,N_29968,N_25057);
nand UO_2443 (O_2443,N_26287,N_24061);
xnor UO_2444 (O_2444,N_26173,N_26733);
xor UO_2445 (O_2445,N_27095,N_25185);
or UO_2446 (O_2446,N_25244,N_29622);
nor UO_2447 (O_2447,N_29455,N_26240);
xor UO_2448 (O_2448,N_25231,N_28417);
xor UO_2449 (O_2449,N_28332,N_27229);
xnor UO_2450 (O_2450,N_29242,N_24417);
nor UO_2451 (O_2451,N_28734,N_26900);
nor UO_2452 (O_2452,N_24058,N_24881);
and UO_2453 (O_2453,N_26257,N_25096);
and UO_2454 (O_2454,N_29250,N_27029);
and UO_2455 (O_2455,N_28534,N_26371);
xnor UO_2456 (O_2456,N_28367,N_24366);
nor UO_2457 (O_2457,N_25423,N_25172);
nor UO_2458 (O_2458,N_24817,N_24182);
and UO_2459 (O_2459,N_25514,N_27663);
or UO_2460 (O_2460,N_27746,N_25360);
nand UO_2461 (O_2461,N_24654,N_27512);
or UO_2462 (O_2462,N_28350,N_26519);
nor UO_2463 (O_2463,N_25532,N_26945);
or UO_2464 (O_2464,N_27543,N_24828);
and UO_2465 (O_2465,N_26561,N_29005);
or UO_2466 (O_2466,N_27399,N_26129);
nand UO_2467 (O_2467,N_28961,N_26708);
or UO_2468 (O_2468,N_27380,N_25618);
nor UO_2469 (O_2469,N_27212,N_29832);
xor UO_2470 (O_2470,N_25842,N_27055);
and UO_2471 (O_2471,N_26855,N_25835);
nand UO_2472 (O_2472,N_24897,N_24343);
nand UO_2473 (O_2473,N_25134,N_27825);
or UO_2474 (O_2474,N_28440,N_24433);
or UO_2475 (O_2475,N_26381,N_25501);
and UO_2476 (O_2476,N_25671,N_26979);
xnor UO_2477 (O_2477,N_28622,N_29437);
nor UO_2478 (O_2478,N_25336,N_27293);
xor UO_2479 (O_2479,N_25599,N_26351);
xnor UO_2480 (O_2480,N_28642,N_25656);
xnor UO_2481 (O_2481,N_26829,N_24543);
nand UO_2482 (O_2482,N_28069,N_27580);
xnor UO_2483 (O_2483,N_29416,N_25300);
xor UO_2484 (O_2484,N_29077,N_26192);
and UO_2485 (O_2485,N_29281,N_25745);
nand UO_2486 (O_2486,N_26903,N_24255);
and UO_2487 (O_2487,N_27897,N_28684);
nand UO_2488 (O_2488,N_28712,N_29083);
or UO_2489 (O_2489,N_26017,N_26958);
and UO_2490 (O_2490,N_28540,N_24244);
nor UO_2491 (O_2491,N_28689,N_26925);
nor UO_2492 (O_2492,N_26816,N_25277);
nand UO_2493 (O_2493,N_25204,N_24368);
nand UO_2494 (O_2494,N_24450,N_26668);
nand UO_2495 (O_2495,N_29177,N_26003);
xor UO_2496 (O_2496,N_28803,N_27898);
or UO_2497 (O_2497,N_24661,N_24922);
and UO_2498 (O_2498,N_28060,N_25683);
or UO_2499 (O_2499,N_24066,N_24849);
nor UO_2500 (O_2500,N_28512,N_26299);
nor UO_2501 (O_2501,N_25930,N_27621);
xnor UO_2502 (O_2502,N_24053,N_28107);
and UO_2503 (O_2503,N_28073,N_25165);
xor UO_2504 (O_2504,N_25845,N_25761);
xnor UO_2505 (O_2505,N_27086,N_28119);
xnor UO_2506 (O_2506,N_28153,N_29699);
nor UO_2507 (O_2507,N_25851,N_28857);
xnor UO_2508 (O_2508,N_25187,N_25104);
nor UO_2509 (O_2509,N_29770,N_24937);
and UO_2510 (O_2510,N_28849,N_24454);
nor UO_2511 (O_2511,N_28331,N_27201);
or UO_2512 (O_2512,N_29043,N_29528);
and UO_2513 (O_2513,N_24080,N_28907);
or UO_2514 (O_2514,N_27313,N_27506);
xor UO_2515 (O_2515,N_27295,N_29880);
nand UO_2516 (O_2516,N_24614,N_29542);
xnor UO_2517 (O_2517,N_25462,N_27667);
nand UO_2518 (O_2518,N_25482,N_24030);
nand UO_2519 (O_2519,N_29549,N_25089);
nand UO_2520 (O_2520,N_29947,N_25213);
and UO_2521 (O_2521,N_24664,N_29684);
nor UO_2522 (O_2522,N_24093,N_28780);
and UO_2523 (O_2523,N_29504,N_28504);
and UO_2524 (O_2524,N_29115,N_27251);
and UO_2525 (O_2525,N_27508,N_26939);
nand UO_2526 (O_2526,N_24357,N_25093);
nand UO_2527 (O_2527,N_27533,N_24913);
nand UO_2528 (O_2528,N_24145,N_26244);
and UO_2529 (O_2529,N_29056,N_26050);
xnor UO_2530 (O_2530,N_27213,N_24300);
or UO_2531 (O_2531,N_27505,N_29475);
and UO_2532 (O_2532,N_25287,N_27115);
xor UO_2533 (O_2533,N_26384,N_27753);
and UO_2534 (O_2534,N_25619,N_29937);
and UO_2535 (O_2535,N_29810,N_28697);
nand UO_2536 (O_2536,N_28142,N_29909);
nor UO_2537 (O_2537,N_28606,N_25478);
and UO_2538 (O_2538,N_24001,N_26837);
or UO_2539 (O_2539,N_27498,N_26546);
nor UO_2540 (O_2540,N_24546,N_25454);
nand UO_2541 (O_2541,N_28583,N_26357);
or UO_2542 (O_2542,N_24161,N_28188);
xnor UO_2543 (O_2543,N_28752,N_26651);
or UO_2544 (O_2544,N_27881,N_27984);
and UO_2545 (O_2545,N_27475,N_29928);
or UO_2546 (O_2546,N_25684,N_28178);
nand UO_2547 (O_2547,N_24520,N_29954);
or UO_2548 (O_2548,N_26399,N_28912);
nor UO_2549 (O_2549,N_24857,N_26127);
nor UO_2550 (O_2550,N_25736,N_24854);
and UO_2551 (O_2551,N_25346,N_26355);
xor UO_2552 (O_2552,N_29835,N_26440);
xor UO_2553 (O_2553,N_24794,N_28580);
and UO_2554 (O_2554,N_24183,N_29662);
nor UO_2555 (O_2555,N_26585,N_28309);
nand UO_2556 (O_2556,N_24410,N_28526);
and UO_2557 (O_2557,N_25784,N_27674);
nor UO_2558 (O_2558,N_29852,N_27883);
or UO_2559 (O_2559,N_28900,N_28094);
nand UO_2560 (O_2560,N_27639,N_27162);
nor UO_2561 (O_2561,N_28743,N_25855);
and UO_2562 (O_2562,N_25476,N_28099);
or UO_2563 (O_2563,N_26051,N_28531);
xnor UO_2564 (O_2564,N_25529,N_29867);
and UO_2565 (O_2565,N_26618,N_24418);
xnor UO_2566 (O_2566,N_27448,N_26008);
xnor UO_2567 (O_2567,N_27860,N_24732);
or UO_2568 (O_2568,N_26703,N_27079);
or UO_2569 (O_2569,N_26001,N_28357);
nor UO_2570 (O_2570,N_29762,N_28128);
nor UO_2571 (O_2571,N_28447,N_24253);
and UO_2572 (O_2572,N_28810,N_29503);
xnor UO_2573 (O_2573,N_25753,N_28014);
xor UO_2574 (O_2574,N_28378,N_26521);
or UO_2575 (O_2575,N_24250,N_27478);
or UO_2576 (O_2576,N_29051,N_24943);
or UO_2577 (O_2577,N_29488,N_27407);
or UO_2578 (O_2578,N_24339,N_28109);
or UO_2579 (O_2579,N_29737,N_27490);
nand UO_2580 (O_2580,N_24880,N_28623);
and UO_2581 (O_2581,N_29182,N_27184);
xnor UO_2582 (O_2582,N_28883,N_27450);
nor UO_2583 (O_2583,N_25840,N_27622);
xor UO_2584 (O_2584,N_26169,N_27576);
nor UO_2585 (O_2585,N_27205,N_27368);
and UO_2586 (O_2586,N_27731,N_27454);
nand UO_2587 (O_2587,N_25504,N_28224);
nand UO_2588 (O_2588,N_28483,N_28256);
xor UO_2589 (O_2589,N_27631,N_24287);
or UO_2590 (O_2590,N_27878,N_28552);
or UO_2591 (O_2591,N_28275,N_29058);
nand UO_2592 (O_2592,N_24969,N_24990);
xor UO_2593 (O_2593,N_26327,N_26433);
xor UO_2594 (O_2594,N_27460,N_24575);
nor UO_2595 (O_2595,N_28769,N_26666);
nand UO_2596 (O_2596,N_25124,N_27314);
xor UO_2597 (O_2597,N_24703,N_24682);
nand UO_2598 (O_2598,N_28000,N_29358);
nor UO_2599 (O_2599,N_25525,N_24508);
xor UO_2600 (O_2600,N_26483,N_26088);
xnor UO_2601 (O_2601,N_24628,N_24868);
and UO_2602 (O_2602,N_24321,N_26766);
xnor UO_2603 (O_2603,N_26333,N_25564);
nor UO_2604 (O_2604,N_24534,N_24799);
or UO_2605 (O_2605,N_24188,N_26345);
or UO_2606 (O_2606,N_28970,N_27847);
or UO_2607 (O_2607,N_29367,N_28453);
and UO_2608 (O_2608,N_25728,N_25531);
xnor UO_2609 (O_2609,N_27420,N_27983);
xnor UO_2610 (O_2610,N_28513,N_28643);
xnor UO_2611 (O_2611,N_25076,N_26163);
nor UO_2612 (O_2612,N_25101,N_27737);
and UO_2613 (O_2613,N_28114,N_27266);
nor UO_2614 (O_2614,N_27089,N_24883);
nor UO_2615 (O_2615,N_27788,N_28723);
nand UO_2616 (O_2616,N_26195,N_25959);
nand UO_2617 (O_2617,N_26353,N_24169);
and UO_2618 (O_2618,N_24036,N_29122);
nor UO_2619 (O_2619,N_29319,N_24942);
xor UO_2620 (O_2620,N_25866,N_28484);
or UO_2621 (O_2621,N_28206,N_24147);
or UO_2622 (O_2622,N_26065,N_26993);
nor UO_2623 (O_2623,N_27013,N_24499);
nor UO_2624 (O_2624,N_24041,N_29539);
or UO_2625 (O_2625,N_27820,N_24399);
and UO_2626 (O_2626,N_26230,N_27710);
or UO_2627 (O_2627,N_29591,N_29003);
or UO_2628 (O_2628,N_29452,N_29307);
xor UO_2629 (O_2629,N_25281,N_28305);
nor UO_2630 (O_2630,N_24709,N_27202);
nor UO_2631 (O_2631,N_26184,N_29912);
xnor UO_2632 (O_2632,N_26338,N_27959);
nor UO_2633 (O_2633,N_26637,N_28506);
xor UO_2634 (O_2634,N_28352,N_25326);
and UO_2635 (O_2635,N_28250,N_24804);
or UO_2636 (O_2636,N_29673,N_24389);
nor UO_2637 (O_2637,N_24395,N_26352);
nand UO_2638 (O_2638,N_25370,N_26229);
nor UO_2639 (O_2639,N_27784,N_29484);
xor UO_2640 (O_2640,N_25434,N_24840);
xor UO_2641 (O_2641,N_24320,N_26406);
and UO_2642 (O_2642,N_27338,N_26780);
nand UO_2643 (O_2643,N_25384,N_24404);
nand UO_2644 (O_2644,N_26026,N_25979);
xnor UO_2645 (O_2645,N_29638,N_24657);
or UO_2646 (O_2646,N_28798,N_24242);
and UO_2647 (O_2647,N_29808,N_27743);
and UO_2648 (O_2648,N_27559,N_24353);
or UO_2649 (O_2649,N_28201,N_27790);
nor UO_2650 (O_2650,N_25223,N_26630);
or UO_2651 (O_2651,N_29510,N_26687);
xor UO_2652 (O_2652,N_28369,N_25188);
nor UO_2653 (O_2653,N_28462,N_25288);
nor UO_2654 (O_2654,N_27626,N_26167);
nand UO_2655 (O_2655,N_28018,N_24107);
nor UO_2656 (O_2656,N_29266,N_29533);
xnor UO_2657 (O_2657,N_28765,N_25026);
or UO_2658 (O_2658,N_25769,N_24671);
xor UO_2659 (O_2659,N_27158,N_25236);
nor UO_2660 (O_2660,N_28170,N_26724);
nor UO_2661 (O_2661,N_27936,N_27452);
nand UO_2662 (O_2662,N_24721,N_28553);
nor UO_2663 (O_2663,N_24155,N_27204);
nor UO_2664 (O_2664,N_29305,N_28856);
xor UO_2665 (O_2665,N_28566,N_29676);
nor UO_2666 (O_2666,N_27884,N_24656);
nor UO_2667 (O_2667,N_24248,N_24079);
and UO_2668 (O_2668,N_24673,N_27556);
xor UO_2669 (O_2669,N_24129,N_25405);
nand UO_2670 (O_2670,N_29557,N_27855);
and UO_2671 (O_2671,N_29388,N_28043);
nand UO_2672 (O_2672,N_28160,N_24858);
nand UO_2673 (O_2673,N_28877,N_24962);
or UO_2674 (O_2674,N_28113,N_27854);
nor UO_2675 (O_2675,N_27177,N_28888);
xnor UO_2676 (O_2676,N_24529,N_27296);
nor UO_2677 (O_2677,N_27133,N_26494);
nand UO_2678 (O_2678,N_29551,N_28460);
xnor UO_2679 (O_2679,N_27003,N_27558);
and UO_2680 (O_2680,N_28312,N_26709);
and UO_2681 (O_2681,N_25566,N_28095);
or UO_2682 (O_2682,N_27345,N_27792);
and UO_2683 (O_2683,N_29128,N_29344);
nor UO_2684 (O_2684,N_26258,N_26162);
or UO_2685 (O_2685,N_26754,N_27187);
and UO_2686 (O_2686,N_29565,N_28673);
or UO_2687 (O_2687,N_24831,N_29636);
nand UO_2688 (O_2688,N_26268,N_26627);
nand UO_2689 (O_2689,N_26373,N_28175);
nor UO_2690 (O_2690,N_29718,N_29917);
or UO_2691 (O_2691,N_25805,N_27582);
or UO_2692 (O_2692,N_26147,N_29763);
nor UO_2693 (O_2693,N_25119,N_28016);
nand UO_2694 (O_2694,N_24578,N_26415);
and UO_2695 (O_2695,N_29406,N_24997);
nor UO_2696 (O_2696,N_29330,N_27823);
and UO_2697 (O_2697,N_26028,N_29966);
nand UO_2698 (O_2698,N_24552,N_24051);
and UO_2699 (O_2699,N_27194,N_27882);
nor UO_2700 (O_2700,N_27322,N_25030);
nor UO_2701 (O_2701,N_24968,N_24571);
xor UO_2702 (O_2702,N_25450,N_29847);
nand UO_2703 (O_2703,N_26936,N_25974);
or UO_2704 (O_2704,N_27956,N_27845);
xor UO_2705 (O_2705,N_27813,N_25179);
or UO_2706 (O_2706,N_26143,N_27357);
nor UO_2707 (O_2707,N_26866,N_27259);
nand UO_2708 (O_2708,N_25505,N_29260);
xnor UO_2709 (O_2709,N_26020,N_25733);
or UO_2710 (O_2710,N_25726,N_28864);
xnor UO_2711 (O_2711,N_28988,N_25291);
nand UO_2712 (O_2712,N_28722,N_26995);
and UO_2713 (O_2713,N_24020,N_25055);
xnor UO_2714 (O_2714,N_25924,N_29451);
or UO_2715 (O_2715,N_25606,N_26449);
xnor UO_2716 (O_2716,N_29972,N_24956);
or UO_2717 (O_2717,N_27821,N_25789);
nand UO_2718 (O_2718,N_28644,N_28439);
nand UO_2719 (O_2719,N_28322,N_29301);
nand UO_2720 (O_2720,N_25864,N_29643);
xor UO_2721 (O_2721,N_29070,N_25675);
and UO_2722 (O_2722,N_27082,N_24876);
xor UO_2723 (O_2723,N_27157,N_25105);
and UO_2724 (O_2724,N_26767,N_28629);
xor UO_2725 (O_2725,N_27676,N_28680);
or UO_2726 (O_2726,N_26976,N_27035);
xor UO_2727 (O_2727,N_29843,N_29752);
and UO_2728 (O_2728,N_29746,N_28608);
nor UO_2729 (O_2729,N_26545,N_25477);
and UO_2730 (O_2730,N_28282,N_24768);
nor UO_2731 (O_2731,N_26513,N_27100);
or UO_2732 (O_2732,N_28683,N_27463);
nor UO_2733 (O_2733,N_28072,N_25844);
nor UO_2734 (O_2734,N_27527,N_25246);
nand UO_2735 (O_2735,N_26858,N_28731);
xnor UO_2736 (O_2736,N_25340,N_29511);
and UO_2737 (O_2737,N_29589,N_27634);
nand UO_2738 (O_2738,N_24782,N_27291);
or UO_2739 (O_2739,N_27125,N_27698);
xnor UO_2740 (O_2740,N_24812,N_27525);
nor UO_2741 (O_2741,N_24882,N_27782);
xnor UO_2742 (O_2742,N_29964,N_25799);
xor UO_2743 (O_2743,N_29748,N_29262);
or UO_2744 (O_2744,N_26652,N_25927);
nand UO_2745 (O_2745,N_29826,N_28426);
and UO_2746 (O_2746,N_26213,N_24655);
nand UO_2747 (O_2747,N_29925,N_27299);
nor UO_2748 (O_2748,N_27023,N_27763);
xnor UO_2749 (O_2749,N_29424,N_25362);
nor UO_2750 (O_2750,N_26392,N_29278);
xor UO_2751 (O_2751,N_28158,N_24326);
xnor UO_2752 (O_2752,N_25667,N_24527);
nor UO_2753 (O_2753,N_27775,N_27557);
or UO_2754 (O_2754,N_24016,N_27832);
and UO_2755 (O_2755,N_29910,N_24948);
xnor UO_2756 (O_2756,N_29602,N_27568);
xor UO_2757 (O_2757,N_25907,N_26659);
or UO_2758 (O_2758,N_28598,N_24192);
nor UO_2759 (O_2759,N_26924,N_24696);
nand UO_2760 (O_2760,N_25135,N_26613);
and UO_2761 (O_2761,N_29593,N_29690);
nand UO_2762 (O_2762,N_28742,N_24576);
xor UO_2763 (O_2763,N_24544,N_26800);
nand UO_2764 (O_2764,N_28500,N_28279);
xor UO_2765 (O_2765,N_25468,N_29623);
nand UO_2766 (O_2766,N_29264,N_28852);
nand UO_2767 (O_2767,N_24423,N_25757);
nor UO_2768 (O_2768,N_25356,N_26033);
nand UO_2769 (O_2769,N_29342,N_25593);
nor UO_2770 (O_2770,N_26982,N_26466);
nand UO_2771 (O_2771,N_29895,N_29288);
xor UO_2772 (O_2772,N_26737,N_24027);
or UO_2773 (O_2773,N_24619,N_29492);
nor UO_2774 (O_2774,N_25062,N_27226);
xor UO_2775 (O_2775,N_28197,N_29580);
nand UO_2776 (O_2776,N_27445,N_28111);
xnor UO_2777 (O_2777,N_27101,N_25163);
nor UO_2778 (O_2778,N_27280,N_25490);
xnor UO_2779 (O_2779,N_24597,N_27504);
or UO_2780 (O_2780,N_24615,N_25574);
and UO_2781 (O_2781,N_28334,N_26038);
and UO_2782 (O_2782,N_25788,N_29283);
and UO_2783 (O_2783,N_29588,N_25786);
and UO_2784 (O_2784,N_27524,N_28402);
nand UO_2785 (O_2785,N_26796,N_29778);
xor UO_2786 (O_2786,N_26954,N_28169);
nand UO_2787 (O_2787,N_25655,N_28068);
or UO_2788 (O_2788,N_29775,N_28226);
nand UO_2789 (O_2789,N_24031,N_24586);
or UO_2790 (O_2790,N_24677,N_24439);
nor UO_2791 (O_2791,N_29129,N_29561);
or UO_2792 (O_2792,N_24823,N_25729);
or UO_2793 (O_2793,N_27633,N_27933);
xnor UO_2794 (O_2794,N_28471,N_28601);
or UO_2795 (O_2795,N_27643,N_29935);
nand UO_2796 (O_2796,N_25996,N_27917);
or UO_2797 (O_2797,N_28755,N_25560);
and UO_2798 (O_2798,N_25227,N_24964);
or UO_2799 (O_2799,N_28238,N_24547);
nor UO_2800 (O_2800,N_25077,N_25743);
nor UO_2801 (O_2801,N_27169,N_29218);
xnor UO_2802 (O_2802,N_26000,N_25942);
or UO_2803 (O_2803,N_27721,N_25069);
nor UO_2804 (O_2804,N_28654,N_25013);
and UO_2805 (O_2805,N_27171,N_25256);
nor UO_2806 (O_2806,N_29803,N_29856);
nand UO_2807 (O_2807,N_29785,N_25318);
or UO_2808 (O_2808,N_24772,N_25210);
nor UO_2809 (O_2809,N_26881,N_27028);
and UO_2810 (O_2810,N_24024,N_28354);
nor UO_2811 (O_2811,N_27754,N_29809);
nand UO_2812 (O_2812,N_27907,N_24301);
nand UO_2813 (O_2813,N_27097,N_25283);
nand UO_2814 (O_2814,N_24712,N_29553);
and UO_2815 (O_2815,N_25145,N_29215);
nor UO_2816 (O_2816,N_26224,N_29547);
xor UO_2817 (O_2817,N_29370,N_28882);
xor UO_2818 (O_2818,N_25828,N_24401);
nand UO_2819 (O_2819,N_28671,N_29219);
nand UO_2820 (O_2820,N_29899,N_25200);
xnor UO_2821 (O_2821,N_28112,N_26851);
or UO_2822 (O_2822,N_29914,N_25307);
nand UO_2823 (O_2823,N_26181,N_26344);
or UO_2824 (O_2824,N_25023,N_28011);
and UO_2825 (O_2825,N_24247,N_29405);
nand UO_2826 (O_2826,N_24471,N_28122);
xor UO_2827 (O_2827,N_28507,N_29436);
and UO_2828 (O_2828,N_27873,N_24348);
or UO_2829 (O_2829,N_27953,N_26396);
nor UO_2830 (O_2830,N_28196,N_28999);
or UO_2831 (O_2831,N_24796,N_26165);
and UO_2832 (O_2832,N_28631,N_24239);
and UO_2833 (O_2833,N_29822,N_27625);
and UO_2834 (O_2834,N_25361,N_28693);
nand UO_2835 (O_2835,N_24201,N_26160);
nor UO_2836 (O_2836,N_29321,N_29519);
and UO_2837 (O_2837,N_26276,N_29500);
and UO_2838 (O_2838,N_24704,N_24377);
nand UO_2839 (O_2839,N_27590,N_24136);
nor UO_2840 (O_2840,N_25730,N_28773);
and UO_2841 (O_2841,N_25106,N_24419);
nand UO_2842 (O_2842,N_29730,N_28204);
and UO_2843 (O_2843,N_25333,N_25180);
nor UO_2844 (O_2844,N_24516,N_28788);
nor UO_2845 (O_2845,N_27877,N_26987);
nand UO_2846 (O_2846,N_29147,N_27659);
and UO_2847 (O_2847,N_24528,N_27502);
and UO_2848 (O_2848,N_26341,N_28653);
nor UO_2849 (O_2849,N_28320,N_25937);
nor UO_2850 (O_2850,N_24724,N_28931);
xnor UO_2851 (O_2851,N_27353,N_27068);
or UO_2852 (O_2852,N_27181,N_25229);
nor UO_2853 (O_2853,N_29963,N_24729);
or UO_2854 (O_2854,N_27546,N_25500);
nand UO_2855 (O_2855,N_28103,N_27227);
or UO_2856 (O_2856,N_24280,N_29644);
nand UO_2857 (O_2857,N_28263,N_26894);
nand UO_2858 (O_2858,N_29235,N_24268);
nand UO_2859 (O_2859,N_24683,N_27575);
and UO_2860 (O_2860,N_25102,N_25238);
nand UO_2861 (O_2861,N_25373,N_27236);
or UO_2862 (O_2862,N_24209,N_25751);
nor UO_2863 (O_2863,N_28548,N_27577);
nand UO_2864 (O_2864,N_24900,N_29360);
nand UO_2865 (O_2865,N_27124,N_29225);
and UO_2866 (O_2866,N_29945,N_24082);
xor UO_2867 (O_2867,N_28766,N_26110);
nor UO_2868 (O_2868,N_25315,N_25727);
nor UO_2869 (O_2869,N_27116,N_26247);
or UO_2870 (O_2870,N_29924,N_25785);
xnor UO_2871 (O_2871,N_24869,N_24025);
or UO_2872 (O_2872,N_28741,N_28547);
xnor UO_2873 (O_2873,N_27815,N_24548);
nand UO_2874 (O_2874,N_24097,N_26817);
nand UO_2875 (O_2875,N_24660,N_29696);
xor UO_2876 (O_2876,N_28042,N_24078);
and UO_2877 (O_2877,N_28616,N_26952);
nand UO_2878 (O_2878,N_29052,N_28809);
and UO_2879 (O_2879,N_27677,N_29583);
nand UO_2880 (O_2880,N_29466,N_26170);
nand UO_2881 (O_2881,N_26596,N_27398);
nand UO_2882 (O_2882,N_27961,N_26818);
xnor UO_2883 (O_2883,N_26113,N_24480);
nor UO_2884 (O_2884,N_24802,N_27429);
nor UO_2885 (O_2885,N_29508,N_24500);
nor UO_2886 (O_2886,N_24413,N_25581);
nand UO_2887 (O_2887,N_26431,N_27105);
xnor UO_2888 (O_2888,N_27545,N_24084);
nand UO_2889 (O_2889,N_28789,N_26611);
xnor UO_2890 (O_2890,N_25954,N_28465);
or UO_2891 (O_2891,N_26558,N_26297);
or UO_2892 (O_2892,N_25417,N_27708);
or UO_2893 (O_2893,N_27221,N_24663);
or UO_2894 (O_2894,N_26340,N_29916);
nor UO_2895 (O_2895,N_24920,N_26902);
nor UO_2896 (O_2896,N_28135,N_24565);
and UO_2897 (O_2897,N_26202,N_26968);
nand UO_2898 (O_2898,N_24170,N_27044);
xor UO_2899 (O_2899,N_25951,N_26582);
xor UO_2900 (O_2900,N_27664,N_27401);
nor UO_2901 (O_2901,N_28467,N_26542);
xor UO_2902 (O_2902,N_24921,N_26702);
nand UO_2903 (O_2903,N_27139,N_28997);
nor UO_2904 (O_2904,N_27188,N_28360);
and UO_2905 (O_2905,N_24739,N_29754);
and UO_2906 (O_2906,N_29325,N_29449);
nand UO_2907 (O_2907,N_26832,N_26324);
nand UO_2908 (O_2908,N_26501,N_24762);
and UO_2909 (O_2909,N_29433,N_25048);
xor UO_2910 (O_2910,N_25677,N_26142);
xor UO_2911 (O_2911,N_29221,N_26067);
and UO_2912 (O_2912,N_27861,N_27354);
and UO_2913 (O_2913,N_29394,N_27482);
nand UO_2914 (O_2914,N_27949,N_26222);
nand UO_2915 (O_2915,N_24679,N_26389);
nor UO_2916 (O_2916,N_25990,N_29816);
xor UO_2917 (O_2917,N_28571,N_24148);
nor UO_2918 (O_2918,N_24488,N_24262);
xnor UO_2919 (O_2919,N_29284,N_29108);
or UO_2920 (O_2920,N_26471,N_27658);
nand UO_2921 (O_2921,N_27346,N_28156);
nand UO_2922 (O_2922,N_25831,N_28232);
or UO_2923 (O_2923,N_26549,N_26292);
nand UO_2924 (O_2924,N_26445,N_24009);
and UO_2925 (O_2925,N_24396,N_26055);
or UO_2926 (O_2926,N_25820,N_26189);
and UO_2927 (O_2927,N_25687,N_28687);
nor UO_2928 (O_2928,N_28739,N_29246);
xor UO_2929 (O_2929,N_28300,N_25195);
xnor UO_2930 (O_2930,N_26847,N_28001);
or UO_2931 (O_2931,N_24902,N_24177);
and UO_2932 (O_2932,N_24464,N_26765);
nor UO_2933 (O_2933,N_29865,N_24018);
or UO_2934 (O_2934,N_28003,N_27253);
xnor UO_2935 (O_2935,N_26006,N_29723);
nand UO_2936 (O_2936,N_28476,N_24156);
nand UO_2937 (O_2937,N_27298,N_24493);
and UO_2938 (O_2938,N_26068,N_25827);
nand UO_2939 (O_2939,N_26386,N_24862);
xnor UO_2940 (O_2940,N_26183,N_29767);
nand UO_2941 (O_2941,N_29209,N_27231);
and UO_2942 (O_2942,N_29678,N_24398);
nor UO_2943 (O_2943,N_27858,N_27381);
xor UO_2944 (O_2944,N_25731,N_28106);
or UO_2945 (O_2945,N_24864,N_28853);
xnor UO_2946 (O_2946,N_27240,N_27747);
and UO_2947 (O_2947,N_25580,N_26478);
nor UO_2948 (O_2948,N_24095,N_29948);
nor UO_2949 (O_2949,N_24198,N_24730);
and UO_2950 (O_2950,N_27408,N_27819);
and UO_2951 (O_2951,N_26364,N_29675);
and UO_2952 (O_2952,N_27161,N_25696);
nand UO_2953 (O_2953,N_24074,N_27515);
nand UO_2954 (O_2954,N_26641,N_26346);
nand UO_2955 (O_2955,N_25207,N_27373);
xor UO_2956 (O_2956,N_29769,N_27535);
or UO_2957 (O_2957,N_28059,N_24167);
or UO_2958 (O_2958,N_26070,N_29317);
xor UO_2959 (O_2959,N_25688,N_25635);
or UO_2960 (O_2960,N_28656,N_26470);
nand UO_2961 (O_2961,N_25376,N_27442);
xnor UO_2962 (O_2962,N_29382,N_24807);
nor UO_2963 (O_2963,N_24570,N_29462);
nor UO_2964 (O_2964,N_26121,N_26156);
xor UO_2965 (O_2965,N_26312,N_25556);
or UO_2966 (O_2966,N_29478,N_28753);
nand UO_2967 (O_2967,N_29359,N_26282);
and UO_2968 (O_2968,N_27386,N_29999);
nor UO_2969 (O_2969,N_27904,N_27128);
and UO_2970 (O_2970,N_26285,N_26725);
nor UO_2971 (O_2971,N_27686,N_29657);
nand UO_2972 (O_2972,N_27985,N_25544);
xor UO_2973 (O_2973,N_29798,N_25998);
nor UO_2974 (O_2974,N_26622,N_29842);
nor UO_2975 (O_2975,N_27981,N_24166);
xor UO_2976 (O_2976,N_29897,N_26420);
xor UO_2977 (O_2977,N_29744,N_28341);
nand UO_2978 (O_2978,N_26468,N_28281);
or UO_2979 (O_2979,N_26427,N_25509);
nand UO_2980 (O_2980,N_26699,N_25366);
nor UO_2981 (O_2981,N_26499,N_24229);
and UO_2982 (O_2982,N_29716,N_29273);
nand UO_2983 (O_2983,N_25344,N_28581);
nand UO_2984 (O_2984,N_26793,N_25445);
or UO_2985 (O_2985,N_25810,N_26537);
or UO_2986 (O_2986,N_26133,N_26084);
nand UO_2987 (O_2987,N_24050,N_28678);
and UO_2988 (O_2988,N_26908,N_28527);
or UO_2989 (O_2989,N_28772,N_29530);
or UO_2990 (O_2990,N_24598,N_26554);
nor UO_2991 (O_2991,N_25496,N_29119);
or UO_2992 (O_2992,N_24089,N_29408);
nand UO_2993 (O_2993,N_25637,N_26118);
nand UO_2994 (O_2994,N_29300,N_25420);
nand UO_2995 (O_2995,N_28233,N_29572);
nand UO_2996 (O_2996,N_29158,N_27144);
nand UO_2997 (O_2997,N_28669,N_25577);
nand UO_2998 (O_2998,N_26704,N_25856);
nand UO_2999 (O_2999,N_25665,N_26947);
nand UO_3000 (O_3000,N_25314,N_24416);
xor UO_3001 (O_3001,N_29426,N_29260);
nor UO_3002 (O_3002,N_28267,N_26049);
or UO_3003 (O_3003,N_25499,N_27435);
nor UO_3004 (O_3004,N_25066,N_24401);
nand UO_3005 (O_3005,N_29641,N_28403);
and UO_3006 (O_3006,N_26159,N_28786);
xnor UO_3007 (O_3007,N_26804,N_24157);
nand UO_3008 (O_3008,N_26931,N_29496);
nand UO_3009 (O_3009,N_28840,N_28863);
and UO_3010 (O_3010,N_29692,N_26648);
or UO_3011 (O_3011,N_27295,N_26771);
xnor UO_3012 (O_3012,N_27612,N_25407);
xnor UO_3013 (O_3013,N_28600,N_27912);
nor UO_3014 (O_3014,N_28197,N_26672);
or UO_3015 (O_3015,N_28612,N_27388);
nor UO_3016 (O_3016,N_28677,N_27628);
nor UO_3017 (O_3017,N_29739,N_25284);
nand UO_3018 (O_3018,N_25060,N_25100);
or UO_3019 (O_3019,N_25331,N_26717);
or UO_3020 (O_3020,N_27810,N_26953);
and UO_3021 (O_3021,N_28677,N_26338);
nand UO_3022 (O_3022,N_29915,N_27015);
nor UO_3023 (O_3023,N_27334,N_25146);
or UO_3024 (O_3024,N_26114,N_25511);
nand UO_3025 (O_3025,N_24500,N_26139);
nand UO_3026 (O_3026,N_24402,N_28196);
nand UO_3027 (O_3027,N_29044,N_28317);
nand UO_3028 (O_3028,N_25552,N_27459);
or UO_3029 (O_3029,N_27662,N_28593);
or UO_3030 (O_3030,N_24854,N_27606);
nand UO_3031 (O_3031,N_24768,N_26177);
nand UO_3032 (O_3032,N_27776,N_24886);
and UO_3033 (O_3033,N_27589,N_24623);
or UO_3034 (O_3034,N_24857,N_24792);
or UO_3035 (O_3035,N_29862,N_26633);
and UO_3036 (O_3036,N_28120,N_28061);
nor UO_3037 (O_3037,N_29481,N_25943);
nand UO_3038 (O_3038,N_29732,N_27583);
xor UO_3039 (O_3039,N_27066,N_27083);
nor UO_3040 (O_3040,N_27147,N_24698);
xnor UO_3041 (O_3041,N_28931,N_24455);
nand UO_3042 (O_3042,N_28295,N_24173);
or UO_3043 (O_3043,N_29641,N_24727);
or UO_3044 (O_3044,N_25397,N_29566);
nand UO_3045 (O_3045,N_29758,N_26799);
nand UO_3046 (O_3046,N_24639,N_29216);
or UO_3047 (O_3047,N_29643,N_28610);
xor UO_3048 (O_3048,N_26179,N_28442);
xnor UO_3049 (O_3049,N_28306,N_29300);
and UO_3050 (O_3050,N_24888,N_25299);
and UO_3051 (O_3051,N_25021,N_24978);
or UO_3052 (O_3052,N_26266,N_25183);
xnor UO_3053 (O_3053,N_27109,N_29734);
nand UO_3054 (O_3054,N_27719,N_29099);
nand UO_3055 (O_3055,N_25292,N_29943);
xor UO_3056 (O_3056,N_26402,N_24838);
nor UO_3057 (O_3057,N_26498,N_25336);
xnor UO_3058 (O_3058,N_26508,N_27208);
and UO_3059 (O_3059,N_26441,N_26550);
or UO_3060 (O_3060,N_28531,N_24344);
xor UO_3061 (O_3061,N_29955,N_24227);
and UO_3062 (O_3062,N_25954,N_28100);
nand UO_3063 (O_3063,N_27176,N_25167);
and UO_3064 (O_3064,N_24666,N_29094);
nand UO_3065 (O_3065,N_29853,N_24338);
nor UO_3066 (O_3066,N_29666,N_25636);
and UO_3067 (O_3067,N_25430,N_27049);
xor UO_3068 (O_3068,N_28658,N_25056);
nand UO_3069 (O_3069,N_25627,N_24135);
and UO_3070 (O_3070,N_24535,N_28002);
xor UO_3071 (O_3071,N_25261,N_29717);
and UO_3072 (O_3072,N_28085,N_25492);
xor UO_3073 (O_3073,N_24755,N_28671);
nand UO_3074 (O_3074,N_27026,N_27477);
and UO_3075 (O_3075,N_27086,N_28674);
nand UO_3076 (O_3076,N_29245,N_24439);
nand UO_3077 (O_3077,N_25697,N_28521);
xnor UO_3078 (O_3078,N_27729,N_28923);
xor UO_3079 (O_3079,N_24626,N_24836);
or UO_3080 (O_3080,N_24953,N_28610);
or UO_3081 (O_3081,N_28334,N_28501);
and UO_3082 (O_3082,N_24636,N_27322);
xor UO_3083 (O_3083,N_26241,N_27247);
nor UO_3084 (O_3084,N_24746,N_25650);
xor UO_3085 (O_3085,N_25604,N_28642);
or UO_3086 (O_3086,N_27705,N_25251);
xnor UO_3087 (O_3087,N_26467,N_28340);
and UO_3088 (O_3088,N_27323,N_25713);
and UO_3089 (O_3089,N_26536,N_29274);
xnor UO_3090 (O_3090,N_26771,N_28494);
or UO_3091 (O_3091,N_27469,N_26501);
and UO_3092 (O_3092,N_29311,N_26345);
nor UO_3093 (O_3093,N_29690,N_29479);
or UO_3094 (O_3094,N_29796,N_26592);
or UO_3095 (O_3095,N_29805,N_28246);
nor UO_3096 (O_3096,N_24635,N_26907);
or UO_3097 (O_3097,N_29562,N_27874);
xnor UO_3098 (O_3098,N_27140,N_24697);
nor UO_3099 (O_3099,N_26508,N_24950);
or UO_3100 (O_3100,N_29579,N_27872);
nor UO_3101 (O_3101,N_27224,N_25103);
nor UO_3102 (O_3102,N_29019,N_26618);
and UO_3103 (O_3103,N_29296,N_27736);
and UO_3104 (O_3104,N_25258,N_26485);
xnor UO_3105 (O_3105,N_26614,N_24571);
nor UO_3106 (O_3106,N_27916,N_28104);
or UO_3107 (O_3107,N_29560,N_27327);
and UO_3108 (O_3108,N_26934,N_29533);
nor UO_3109 (O_3109,N_27707,N_29150);
xor UO_3110 (O_3110,N_27875,N_24247);
nand UO_3111 (O_3111,N_26722,N_26275);
and UO_3112 (O_3112,N_25587,N_26121);
or UO_3113 (O_3113,N_28012,N_24185);
xnor UO_3114 (O_3114,N_27202,N_28782);
xor UO_3115 (O_3115,N_29117,N_29947);
nand UO_3116 (O_3116,N_25658,N_25147);
xnor UO_3117 (O_3117,N_29464,N_29668);
or UO_3118 (O_3118,N_25102,N_25059);
nand UO_3119 (O_3119,N_28959,N_24499);
nor UO_3120 (O_3120,N_25323,N_29458);
and UO_3121 (O_3121,N_26404,N_28521);
and UO_3122 (O_3122,N_28978,N_26046);
and UO_3123 (O_3123,N_25024,N_25620);
and UO_3124 (O_3124,N_29809,N_26004);
nand UO_3125 (O_3125,N_27487,N_28814);
or UO_3126 (O_3126,N_26159,N_27107);
or UO_3127 (O_3127,N_25353,N_26889);
nor UO_3128 (O_3128,N_24091,N_29414);
nor UO_3129 (O_3129,N_27278,N_27063);
and UO_3130 (O_3130,N_25851,N_24716);
or UO_3131 (O_3131,N_25086,N_26036);
xor UO_3132 (O_3132,N_29399,N_26808);
nand UO_3133 (O_3133,N_29894,N_26123);
nand UO_3134 (O_3134,N_25357,N_28943);
or UO_3135 (O_3135,N_24108,N_24247);
nand UO_3136 (O_3136,N_24021,N_28598);
or UO_3137 (O_3137,N_24702,N_28900);
and UO_3138 (O_3138,N_29123,N_25191);
nor UO_3139 (O_3139,N_26973,N_29687);
or UO_3140 (O_3140,N_24614,N_25377);
nor UO_3141 (O_3141,N_28463,N_28825);
nand UO_3142 (O_3142,N_24445,N_26059);
or UO_3143 (O_3143,N_26540,N_28122);
nor UO_3144 (O_3144,N_24974,N_24913);
xor UO_3145 (O_3145,N_25103,N_25887);
nand UO_3146 (O_3146,N_28697,N_24462);
nor UO_3147 (O_3147,N_25338,N_25860);
xor UO_3148 (O_3148,N_29725,N_28312);
and UO_3149 (O_3149,N_29157,N_24940);
and UO_3150 (O_3150,N_29683,N_27135);
or UO_3151 (O_3151,N_28808,N_27923);
nor UO_3152 (O_3152,N_24886,N_24881);
xor UO_3153 (O_3153,N_28596,N_28090);
nand UO_3154 (O_3154,N_27612,N_25133);
nor UO_3155 (O_3155,N_24411,N_24655);
and UO_3156 (O_3156,N_25402,N_29723);
nand UO_3157 (O_3157,N_26530,N_25108);
nor UO_3158 (O_3158,N_28270,N_25055);
xor UO_3159 (O_3159,N_24647,N_26957);
xor UO_3160 (O_3160,N_25648,N_29840);
nand UO_3161 (O_3161,N_25043,N_25951);
nand UO_3162 (O_3162,N_24998,N_25155);
or UO_3163 (O_3163,N_29171,N_25289);
xnor UO_3164 (O_3164,N_28229,N_25299);
nand UO_3165 (O_3165,N_24135,N_29389);
nor UO_3166 (O_3166,N_29119,N_27317);
nor UO_3167 (O_3167,N_27224,N_26953);
nand UO_3168 (O_3168,N_25875,N_24984);
and UO_3169 (O_3169,N_24594,N_24968);
or UO_3170 (O_3170,N_28369,N_29453);
nor UO_3171 (O_3171,N_25605,N_28610);
xnor UO_3172 (O_3172,N_26796,N_27665);
and UO_3173 (O_3173,N_26043,N_27911);
or UO_3174 (O_3174,N_25792,N_25875);
and UO_3175 (O_3175,N_26652,N_25269);
nand UO_3176 (O_3176,N_25290,N_28556);
and UO_3177 (O_3177,N_25821,N_24728);
and UO_3178 (O_3178,N_28556,N_24987);
nand UO_3179 (O_3179,N_28400,N_26165);
xnor UO_3180 (O_3180,N_29579,N_29270);
xor UO_3181 (O_3181,N_28916,N_29259);
nand UO_3182 (O_3182,N_29527,N_27730);
xnor UO_3183 (O_3183,N_26468,N_24367);
nand UO_3184 (O_3184,N_26726,N_28345);
nor UO_3185 (O_3185,N_29885,N_27086);
and UO_3186 (O_3186,N_28674,N_24881);
xnor UO_3187 (O_3187,N_25139,N_25607);
and UO_3188 (O_3188,N_27865,N_29042);
nor UO_3189 (O_3189,N_27014,N_27052);
and UO_3190 (O_3190,N_27267,N_26649);
nand UO_3191 (O_3191,N_28155,N_24592);
and UO_3192 (O_3192,N_26788,N_27152);
nand UO_3193 (O_3193,N_28621,N_26604);
or UO_3194 (O_3194,N_26843,N_29961);
and UO_3195 (O_3195,N_29790,N_28433);
nand UO_3196 (O_3196,N_27011,N_26085);
or UO_3197 (O_3197,N_26155,N_24411);
nor UO_3198 (O_3198,N_27035,N_29027);
and UO_3199 (O_3199,N_29694,N_26054);
xnor UO_3200 (O_3200,N_28708,N_28873);
xnor UO_3201 (O_3201,N_25767,N_24016);
nor UO_3202 (O_3202,N_27862,N_26361);
xor UO_3203 (O_3203,N_28605,N_24034);
or UO_3204 (O_3204,N_24786,N_28351);
nand UO_3205 (O_3205,N_24874,N_26266);
or UO_3206 (O_3206,N_27534,N_26670);
nor UO_3207 (O_3207,N_29890,N_27740);
nand UO_3208 (O_3208,N_25185,N_24058);
nor UO_3209 (O_3209,N_25309,N_29079);
nor UO_3210 (O_3210,N_24739,N_24568);
or UO_3211 (O_3211,N_29463,N_28931);
or UO_3212 (O_3212,N_28518,N_24441);
nand UO_3213 (O_3213,N_25456,N_25678);
and UO_3214 (O_3214,N_29648,N_27350);
and UO_3215 (O_3215,N_27332,N_27765);
and UO_3216 (O_3216,N_25600,N_29172);
xor UO_3217 (O_3217,N_28414,N_24740);
xor UO_3218 (O_3218,N_28952,N_28281);
and UO_3219 (O_3219,N_26011,N_27865);
nor UO_3220 (O_3220,N_25778,N_28201);
and UO_3221 (O_3221,N_29398,N_29466);
or UO_3222 (O_3222,N_29992,N_29702);
nand UO_3223 (O_3223,N_25907,N_26384);
xor UO_3224 (O_3224,N_28005,N_28242);
and UO_3225 (O_3225,N_24167,N_26354);
and UO_3226 (O_3226,N_25679,N_25729);
and UO_3227 (O_3227,N_24367,N_29196);
or UO_3228 (O_3228,N_24038,N_29000);
and UO_3229 (O_3229,N_29696,N_25580);
nor UO_3230 (O_3230,N_24308,N_25152);
or UO_3231 (O_3231,N_25248,N_24536);
nor UO_3232 (O_3232,N_24148,N_28120);
or UO_3233 (O_3233,N_28271,N_24553);
xor UO_3234 (O_3234,N_28663,N_25337);
xnor UO_3235 (O_3235,N_27980,N_26624);
xor UO_3236 (O_3236,N_25078,N_26083);
nand UO_3237 (O_3237,N_25508,N_28619);
xor UO_3238 (O_3238,N_26778,N_28834);
and UO_3239 (O_3239,N_24482,N_27965);
nor UO_3240 (O_3240,N_29879,N_24738);
xnor UO_3241 (O_3241,N_29791,N_29322);
and UO_3242 (O_3242,N_25438,N_28870);
or UO_3243 (O_3243,N_27414,N_25397);
or UO_3244 (O_3244,N_24465,N_27878);
and UO_3245 (O_3245,N_24366,N_28694);
or UO_3246 (O_3246,N_28547,N_25245);
xor UO_3247 (O_3247,N_27452,N_28649);
xnor UO_3248 (O_3248,N_26936,N_29550);
and UO_3249 (O_3249,N_28757,N_27376);
xor UO_3250 (O_3250,N_29527,N_29615);
and UO_3251 (O_3251,N_27183,N_24502);
xor UO_3252 (O_3252,N_28487,N_24678);
or UO_3253 (O_3253,N_26912,N_26259);
nand UO_3254 (O_3254,N_26680,N_29756);
xor UO_3255 (O_3255,N_26966,N_26220);
nor UO_3256 (O_3256,N_24476,N_27139);
or UO_3257 (O_3257,N_29242,N_29967);
xnor UO_3258 (O_3258,N_27111,N_26476);
and UO_3259 (O_3259,N_28395,N_27366);
nand UO_3260 (O_3260,N_25707,N_25197);
or UO_3261 (O_3261,N_26622,N_26538);
nor UO_3262 (O_3262,N_24452,N_27427);
nor UO_3263 (O_3263,N_27614,N_25786);
nor UO_3264 (O_3264,N_29655,N_28797);
or UO_3265 (O_3265,N_24053,N_29950);
xor UO_3266 (O_3266,N_26015,N_26854);
nand UO_3267 (O_3267,N_29406,N_24818);
or UO_3268 (O_3268,N_25272,N_29090);
and UO_3269 (O_3269,N_28119,N_25671);
xor UO_3270 (O_3270,N_27741,N_26967);
and UO_3271 (O_3271,N_29891,N_25902);
nor UO_3272 (O_3272,N_26669,N_24645);
or UO_3273 (O_3273,N_27741,N_24710);
and UO_3274 (O_3274,N_29175,N_24191);
nor UO_3275 (O_3275,N_25852,N_24891);
or UO_3276 (O_3276,N_27278,N_29778);
nor UO_3277 (O_3277,N_27117,N_29938);
or UO_3278 (O_3278,N_25670,N_27326);
and UO_3279 (O_3279,N_25318,N_24617);
or UO_3280 (O_3280,N_25301,N_25417);
nand UO_3281 (O_3281,N_25212,N_27402);
nand UO_3282 (O_3282,N_28929,N_26370);
nand UO_3283 (O_3283,N_28162,N_29748);
nand UO_3284 (O_3284,N_24112,N_25424);
xor UO_3285 (O_3285,N_24818,N_26368);
nor UO_3286 (O_3286,N_26197,N_29162);
nor UO_3287 (O_3287,N_26517,N_27067);
nor UO_3288 (O_3288,N_26815,N_26770);
xnor UO_3289 (O_3289,N_26567,N_25991);
nand UO_3290 (O_3290,N_27963,N_26510);
xnor UO_3291 (O_3291,N_29454,N_29479);
nor UO_3292 (O_3292,N_26969,N_27740);
nor UO_3293 (O_3293,N_24071,N_26875);
nand UO_3294 (O_3294,N_29885,N_26174);
xor UO_3295 (O_3295,N_28602,N_29123);
xnor UO_3296 (O_3296,N_24743,N_25515);
or UO_3297 (O_3297,N_28075,N_27736);
nor UO_3298 (O_3298,N_28402,N_29262);
and UO_3299 (O_3299,N_29035,N_26121);
xor UO_3300 (O_3300,N_29492,N_28117);
xor UO_3301 (O_3301,N_25757,N_29530);
xnor UO_3302 (O_3302,N_24193,N_25930);
and UO_3303 (O_3303,N_26416,N_28145);
nor UO_3304 (O_3304,N_24774,N_29412);
nor UO_3305 (O_3305,N_29253,N_29365);
or UO_3306 (O_3306,N_26839,N_26468);
nand UO_3307 (O_3307,N_28641,N_28276);
xnor UO_3308 (O_3308,N_28486,N_27951);
or UO_3309 (O_3309,N_27576,N_27676);
or UO_3310 (O_3310,N_29882,N_28575);
or UO_3311 (O_3311,N_29392,N_26177);
nand UO_3312 (O_3312,N_26916,N_26190);
xor UO_3313 (O_3313,N_25580,N_24920);
or UO_3314 (O_3314,N_28173,N_26760);
nor UO_3315 (O_3315,N_26726,N_25687);
xor UO_3316 (O_3316,N_25821,N_26506);
or UO_3317 (O_3317,N_28908,N_29051);
or UO_3318 (O_3318,N_27715,N_24979);
or UO_3319 (O_3319,N_27671,N_29865);
xor UO_3320 (O_3320,N_26295,N_24587);
nor UO_3321 (O_3321,N_27826,N_29614);
nor UO_3322 (O_3322,N_25357,N_26782);
xor UO_3323 (O_3323,N_25177,N_24491);
nand UO_3324 (O_3324,N_27741,N_29424);
nor UO_3325 (O_3325,N_27520,N_29558);
nand UO_3326 (O_3326,N_24768,N_27347);
xor UO_3327 (O_3327,N_26847,N_25807);
xnor UO_3328 (O_3328,N_26790,N_29425);
nand UO_3329 (O_3329,N_27729,N_27936);
xnor UO_3330 (O_3330,N_27296,N_24358);
nand UO_3331 (O_3331,N_29038,N_28382);
xnor UO_3332 (O_3332,N_25825,N_27247);
xor UO_3333 (O_3333,N_27361,N_25207);
nor UO_3334 (O_3334,N_29342,N_25047);
nor UO_3335 (O_3335,N_27901,N_28227);
nand UO_3336 (O_3336,N_26851,N_29657);
or UO_3337 (O_3337,N_25552,N_26770);
xor UO_3338 (O_3338,N_28207,N_25655);
xnor UO_3339 (O_3339,N_29048,N_27797);
nor UO_3340 (O_3340,N_24136,N_24713);
xor UO_3341 (O_3341,N_25644,N_24976);
and UO_3342 (O_3342,N_24222,N_27283);
nor UO_3343 (O_3343,N_29970,N_26719);
and UO_3344 (O_3344,N_24227,N_24275);
nand UO_3345 (O_3345,N_29893,N_26237);
nor UO_3346 (O_3346,N_24364,N_25554);
nor UO_3347 (O_3347,N_26993,N_28164);
and UO_3348 (O_3348,N_28248,N_26450);
nand UO_3349 (O_3349,N_26725,N_26190);
xor UO_3350 (O_3350,N_25360,N_25768);
or UO_3351 (O_3351,N_29330,N_26684);
or UO_3352 (O_3352,N_26396,N_29325);
nor UO_3353 (O_3353,N_29755,N_29714);
or UO_3354 (O_3354,N_27654,N_25405);
nor UO_3355 (O_3355,N_29706,N_25520);
nand UO_3356 (O_3356,N_28115,N_28488);
and UO_3357 (O_3357,N_29023,N_26186);
xor UO_3358 (O_3358,N_24696,N_27811);
and UO_3359 (O_3359,N_25726,N_29722);
xor UO_3360 (O_3360,N_28473,N_24337);
nor UO_3361 (O_3361,N_29169,N_29377);
nand UO_3362 (O_3362,N_27635,N_26563);
nor UO_3363 (O_3363,N_27335,N_27822);
xnor UO_3364 (O_3364,N_27079,N_28380);
and UO_3365 (O_3365,N_27129,N_27584);
xor UO_3366 (O_3366,N_24628,N_27239);
or UO_3367 (O_3367,N_24281,N_26608);
nor UO_3368 (O_3368,N_29406,N_28078);
xnor UO_3369 (O_3369,N_29416,N_27552);
and UO_3370 (O_3370,N_27393,N_27793);
xnor UO_3371 (O_3371,N_29113,N_25734);
and UO_3372 (O_3372,N_29150,N_24582);
or UO_3373 (O_3373,N_28739,N_26085);
and UO_3374 (O_3374,N_24726,N_25885);
nand UO_3375 (O_3375,N_26356,N_28993);
or UO_3376 (O_3376,N_25749,N_24937);
or UO_3377 (O_3377,N_29829,N_26225);
xor UO_3378 (O_3378,N_27622,N_25167);
and UO_3379 (O_3379,N_25418,N_29674);
nor UO_3380 (O_3380,N_28671,N_29463);
nand UO_3381 (O_3381,N_27261,N_24301);
or UO_3382 (O_3382,N_27510,N_24789);
nor UO_3383 (O_3383,N_28154,N_25292);
xor UO_3384 (O_3384,N_27026,N_27020);
nand UO_3385 (O_3385,N_28509,N_24554);
nor UO_3386 (O_3386,N_29909,N_29868);
xor UO_3387 (O_3387,N_26970,N_25568);
xor UO_3388 (O_3388,N_27624,N_27775);
and UO_3389 (O_3389,N_26935,N_24726);
and UO_3390 (O_3390,N_27987,N_26280);
and UO_3391 (O_3391,N_29515,N_29697);
or UO_3392 (O_3392,N_24032,N_27694);
nand UO_3393 (O_3393,N_25478,N_26120);
or UO_3394 (O_3394,N_24640,N_27308);
and UO_3395 (O_3395,N_25644,N_27056);
nand UO_3396 (O_3396,N_26010,N_26204);
and UO_3397 (O_3397,N_29046,N_24619);
nor UO_3398 (O_3398,N_29775,N_26150);
and UO_3399 (O_3399,N_29006,N_29002);
xor UO_3400 (O_3400,N_24617,N_25074);
or UO_3401 (O_3401,N_29717,N_29347);
or UO_3402 (O_3402,N_29448,N_27691);
and UO_3403 (O_3403,N_28160,N_29709);
and UO_3404 (O_3404,N_29945,N_25288);
and UO_3405 (O_3405,N_29905,N_24604);
and UO_3406 (O_3406,N_25983,N_25728);
xnor UO_3407 (O_3407,N_25191,N_25211);
and UO_3408 (O_3408,N_25568,N_28088);
and UO_3409 (O_3409,N_24787,N_25509);
and UO_3410 (O_3410,N_27472,N_26028);
and UO_3411 (O_3411,N_27105,N_29636);
nand UO_3412 (O_3412,N_29107,N_26703);
and UO_3413 (O_3413,N_24896,N_24876);
nand UO_3414 (O_3414,N_26550,N_24991);
nor UO_3415 (O_3415,N_26198,N_24641);
and UO_3416 (O_3416,N_29124,N_28673);
or UO_3417 (O_3417,N_26128,N_26062);
nand UO_3418 (O_3418,N_24495,N_29113);
xor UO_3419 (O_3419,N_25320,N_27324);
nor UO_3420 (O_3420,N_25749,N_25579);
or UO_3421 (O_3421,N_24556,N_26858);
xor UO_3422 (O_3422,N_28672,N_25522);
xnor UO_3423 (O_3423,N_27967,N_24786);
nor UO_3424 (O_3424,N_25734,N_24983);
or UO_3425 (O_3425,N_29255,N_27124);
and UO_3426 (O_3426,N_27029,N_27253);
nor UO_3427 (O_3427,N_29988,N_27550);
or UO_3428 (O_3428,N_29995,N_27026);
or UO_3429 (O_3429,N_27590,N_26427);
or UO_3430 (O_3430,N_27320,N_25488);
xor UO_3431 (O_3431,N_25983,N_25169);
and UO_3432 (O_3432,N_26364,N_26228);
nor UO_3433 (O_3433,N_24684,N_24669);
or UO_3434 (O_3434,N_28937,N_27415);
or UO_3435 (O_3435,N_29765,N_27583);
nor UO_3436 (O_3436,N_26169,N_26761);
nor UO_3437 (O_3437,N_25912,N_25392);
nand UO_3438 (O_3438,N_29763,N_24387);
xnor UO_3439 (O_3439,N_29050,N_27575);
or UO_3440 (O_3440,N_27457,N_25025);
or UO_3441 (O_3441,N_27081,N_27732);
xnor UO_3442 (O_3442,N_27793,N_27171);
nand UO_3443 (O_3443,N_27739,N_24024);
nor UO_3444 (O_3444,N_25006,N_28536);
nand UO_3445 (O_3445,N_26296,N_26514);
or UO_3446 (O_3446,N_28859,N_24424);
nor UO_3447 (O_3447,N_26129,N_24255);
xor UO_3448 (O_3448,N_25511,N_26032);
and UO_3449 (O_3449,N_28842,N_24217);
and UO_3450 (O_3450,N_27527,N_28653);
or UO_3451 (O_3451,N_24170,N_29714);
and UO_3452 (O_3452,N_27706,N_28885);
xor UO_3453 (O_3453,N_28544,N_24178);
nand UO_3454 (O_3454,N_28215,N_27459);
nor UO_3455 (O_3455,N_26890,N_25836);
nand UO_3456 (O_3456,N_24588,N_27783);
xor UO_3457 (O_3457,N_24150,N_26894);
nand UO_3458 (O_3458,N_27790,N_25008);
nor UO_3459 (O_3459,N_25237,N_27419);
nor UO_3460 (O_3460,N_29321,N_24726);
xor UO_3461 (O_3461,N_24967,N_24635);
nor UO_3462 (O_3462,N_29638,N_29574);
nor UO_3463 (O_3463,N_28755,N_26016);
nand UO_3464 (O_3464,N_27146,N_24202);
nor UO_3465 (O_3465,N_27467,N_24272);
nand UO_3466 (O_3466,N_26043,N_26727);
nand UO_3467 (O_3467,N_29700,N_28618);
xor UO_3468 (O_3468,N_28697,N_25003);
nor UO_3469 (O_3469,N_29937,N_27871);
nand UO_3470 (O_3470,N_26834,N_27267);
or UO_3471 (O_3471,N_28478,N_24959);
nor UO_3472 (O_3472,N_27026,N_29760);
or UO_3473 (O_3473,N_26852,N_24115);
nor UO_3474 (O_3474,N_24994,N_26825);
or UO_3475 (O_3475,N_27287,N_26972);
or UO_3476 (O_3476,N_25108,N_27876);
and UO_3477 (O_3477,N_29583,N_24284);
or UO_3478 (O_3478,N_29479,N_27716);
and UO_3479 (O_3479,N_29484,N_27984);
and UO_3480 (O_3480,N_28005,N_25732);
nand UO_3481 (O_3481,N_25453,N_25026);
nand UO_3482 (O_3482,N_24269,N_25645);
nor UO_3483 (O_3483,N_24239,N_29938);
nand UO_3484 (O_3484,N_26759,N_24535);
nand UO_3485 (O_3485,N_27087,N_27186);
xnor UO_3486 (O_3486,N_27935,N_26635);
nor UO_3487 (O_3487,N_27332,N_29215);
xnor UO_3488 (O_3488,N_27619,N_25097);
nor UO_3489 (O_3489,N_28202,N_24061);
nand UO_3490 (O_3490,N_24071,N_28869);
nand UO_3491 (O_3491,N_27905,N_25954);
or UO_3492 (O_3492,N_25591,N_29200);
nor UO_3493 (O_3493,N_25573,N_29773);
nor UO_3494 (O_3494,N_29033,N_28957);
xnor UO_3495 (O_3495,N_27425,N_29862);
nor UO_3496 (O_3496,N_25338,N_26874);
nor UO_3497 (O_3497,N_28469,N_25761);
nand UO_3498 (O_3498,N_28116,N_26428);
and UO_3499 (O_3499,N_25314,N_28623);
endmodule