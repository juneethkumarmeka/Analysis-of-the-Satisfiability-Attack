module basic_1000_10000_1500_5_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_358,In_214);
xor U1 (N_1,In_510,In_995);
or U2 (N_2,In_7,In_488);
nor U3 (N_3,In_897,In_245);
xor U4 (N_4,In_97,In_264);
or U5 (N_5,In_376,In_909);
xnor U6 (N_6,In_641,In_415);
xor U7 (N_7,In_262,In_514);
xnor U8 (N_8,In_311,In_340);
and U9 (N_9,In_492,In_568);
nor U10 (N_10,In_741,In_140);
nor U11 (N_11,In_533,In_852);
nand U12 (N_12,In_529,In_180);
and U13 (N_13,In_960,In_870);
nand U14 (N_14,In_189,In_696);
and U15 (N_15,In_699,In_932);
xnor U16 (N_16,In_320,In_829);
or U17 (N_17,In_94,In_871);
xnor U18 (N_18,In_885,In_495);
nor U19 (N_19,In_893,In_435);
or U20 (N_20,In_400,In_946);
nand U21 (N_21,In_344,In_153);
xnor U22 (N_22,In_839,In_198);
and U23 (N_23,In_923,In_194);
or U24 (N_24,In_319,In_802);
or U25 (N_25,In_539,In_117);
nand U26 (N_26,In_670,In_952);
nand U27 (N_27,In_184,In_123);
and U28 (N_28,In_112,In_700);
nor U29 (N_29,In_137,In_273);
xnor U30 (N_30,In_432,In_223);
or U31 (N_31,In_808,In_444);
xnor U32 (N_32,In_485,In_973);
xor U33 (N_33,In_797,In_76);
and U34 (N_34,In_305,In_980);
or U35 (N_35,In_385,In_567);
and U36 (N_36,In_902,In_398);
xor U37 (N_37,In_56,In_339);
and U38 (N_38,In_917,In_436);
or U39 (N_39,In_594,In_66);
or U40 (N_40,In_393,In_636);
or U41 (N_41,In_232,In_517);
or U42 (N_42,In_860,In_589);
nor U43 (N_43,In_763,In_477);
nor U44 (N_44,In_947,In_82);
nor U45 (N_45,In_145,In_32);
and U46 (N_46,In_186,In_507);
xor U47 (N_47,In_801,In_883);
nor U48 (N_48,In_226,In_269);
and U49 (N_49,In_61,In_570);
nor U50 (N_50,In_686,In_289);
xnor U51 (N_51,In_470,In_261);
nor U52 (N_52,In_343,In_12);
or U53 (N_53,In_683,In_614);
or U54 (N_54,In_820,In_668);
nand U55 (N_55,In_384,In_407);
or U56 (N_56,In_162,In_607);
nand U57 (N_57,In_855,In_388);
and U58 (N_58,In_325,In_411);
nand U59 (N_59,In_154,In_687);
and U60 (N_60,In_848,In_595);
and U61 (N_61,In_95,In_943);
or U62 (N_62,In_933,In_654);
and U63 (N_63,In_205,In_886);
or U64 (N_64,In_375,In_966);
xnor U65 (N_65,In_530,In_310);
nor U66 (N_66,In_743,In_134);
and U67 (N_67,In_287,In_793);
and U68 (N_68,In_945,In_337);
nor U69 (N_69,In_299,In_425);
xor U70 (N_70,In_366,In_838);
or U71 (N_71,In_88,In_677);
nand U72 (N_72,In_518,In_635);
nor U73 (N_73,In_833,In_901);
nand U74 (N_74,In_660,In_944);
nor U75 (N_75,In_612,In_212);
nand U76 (N_76,In_234,In_397);
and U77 (N_77,In_35,In_576);
and U78 (N_78,In_775,In_782);
nand U79 (N_79,In_899,In_867);
nand U80 (N_80,In_71,In_132);
xnor U81 (N_81,In_431,In_578);
or U82 (N_82,In_680,In_642);
and U83 (N_83,In_499,In_40);
xnor U84 (N_84,In_950,In_286);
or U85 (N_85,In_513,In_404);
and U86 (N_86,In_896,In_11);
and U87 (N_87,In_599,In_124);
or U88 (N_88,In_815,In_20);
nor U89 (N_89,In_242,In_129);
xor U90 (N_90,In_449,In_42);
or U91 (N_91,In_847,In_998);
nand U92 (N_92,In_949,In_334);
nand U93 (N_93,In_483,In_554);
and U94 (N_94,In_907,In_579);
nor U95 (N_95,In_948,In_955);
nor U96 (N_96,In_377,In_479);
nor U97 (N_97,In_4,In_900);
xnor U98 (N_98,In_715,In_600);
nand U99 (N_99,In_63,In_239);
and U100 (N_100,In_130,In_48);
nand U101 (N_101,In_523,In_742);
or U102 (N_102,In_928,In_993);
and U103 (N_103,In_260,In_355);
nand U104 (N_104,In_638,In_342);
nor U105 (N_105,In_586,In_288);
nand U106 (N_106,In_72,In_656);
nand U107 (N_107,In_231,In_988);
and U108 (N_108,In_942,In_758);
nand U109 (N_109,In_673,In_103);
or U110 (N_110,In_462,In_159);
and U111 (N_111,In_148,In_293);
or U112 (N_112,In_46,In_228);
xnor U113 (N_113,In_109,In_887);
xor U114 (N_114,In_409,In_751);
nor U115 (N_115,In_772,In_716);
nand U116 (N_116,In_224,In_827);
xor U117 (N_117,In_512,In_703);
or U118 (N_118,In_13,In_975);
nand U119 (N_119,In_718,In_633);
nor U120 (N_120,In_978,In_531);
nor U121 (N_121,In_448,In_6);
xor U122 (N_122,In_295,In_545);
nor U123 (N_123,In_329,In_611);
or U124 (N_124,In_433,In_122);
or U125 (N_125,In_596,In_296);
and U126 (N_126,In_753,In_185);
or U127 (N_127,In_606,In_649);
and U128 (N_128,In_965,In_707);
and U129 (N_129,In_27,In_104);
or U130 (N_130,In_18,In_877);
nor U131 (N_131,In_354,In_981);
xnor U132 (N_132,In_475,In_369);
or U133 (N_133,In_745,In_754);
or U134 (N_134,In_836,In_939);
and U135 (N_135,In_583,In_75);
xor U136 (N_136,In_892,In_647);
nand U137 (N_137,In_663,In_776);
nand U138 (N_138,In_328,In_956);
or U139 (N_139,In_556,In_546);
nand U140 (N_140,In_834,In_780);
or U141 (N_141,In_508,In_970);
and U142 (N_142,In_386,In_559);
nor U143 (N_143,In_733,In_868);
nand U144 (N_144,In_884,In_128);
nor U145 (N_145,In_240,In_613);
or U146 (N_146,In_940,In_694);
nand U147 (N_147,In_593,In_506);
or U148 (N_148,In_5,In_681);
nor U149 (N_149,In_958,In_762);
nor U150 (N_150,In_68,In_817);
xor U151 (N_151,In_314,In_674);
or U152 (N_152,In_267,In_915);
or U153 (N_153,In_265,In_620);
or U154 (N_154,In_527,In_637);
and U155 (N_155,In_102,In_62);
and U156 (N_156,In_504,In_29);
nand U157 (N_157,In_1,In_304);
nand U158 (N_158,In_221,In_746);
or U159 (N_159,In_769,In_252);
and U160 (N_160,In_255,In_478);
nor U161 (N_161,In_951,In_230);
xor U162 (N_162,In_350,In_165);
xor U163 (N_163,In_464,In_14);
or U164 (N_164,In_552,In_356);
nor U165 (N_165,In_47,In_617);
xor U166 (N_166,In_662,In_278);
nor U167 (N_167,In_627,In_98);
and U168 (N_168,In_936,In_509);
and U169 (N_169,In_710,In_985);
nand U170 (N_170,In_712,In_237);
nand U171 (N_171,In_428,In_106);
nand U172 (N_172,In_284,In_580);
or U173 (N_173,In_525,In_381);
or U174 (N_174,In_361,In_147);
xnor U175 (N_175,In_172,In_115);
and U176 (N_176,In_591,In_290);
nand U177 (N_177,In_93,In_351);
nor U178 (N_178,In_650,In_786);
or U179 (N_179,In_789,In_999);
nor U180 (N_180,In_891,In_630);
or U181 (N_181,In_968,In_73);
and U182 (N_182,In_77,In_417);
nand U183 (N_183,In_910,In_209);
and U184 (N_184,In_659,In_536);
xnor U185 (N_185,In_308,In_759);
or U186 (N_186,In_248,In_96);
and U187 (N_187,In_938,In_86);
and U188 (N_188,In_179,In_438);
nor U189 (N_189,In_442,In_496);
nor U190 (N_190,In_52,In_116);
and U191 (N_191,In_601,In_878);
or U192 (N_192,In_423,In_332);
or U193 (N_193,In_312,In_90);
nor U194 (N_194,In_53,In_626);
nor U195 (N_195,In_401,In_357);
and U196 (N_196,In_511,In_688);
xnor U197 (N_197,In_418,In_987);
or U198 (N_198,In_434,In_729);
nor U199 (N_199,In_930,In_564);
xnor U200 (N_200,In_806,In_441);
or U201 (N_201,In_822,In_502);
nor U202 (N_202,In_0,In_466);
xnor U203 (N_203,In_997,In_810);
and U204 (N_204,In_452,In_204);
xor U205 (N_205,In_816,In_698);
nand U206 (N_206,In_608,In_60);
nand U207 (N_207,In_675,In_439);
nor U208 (N_208,In_161,In_846);
nand U209 (N_209,In_655,In_830);
nor U210 (N_210,In_573,In_918);
nor U211 (N_211,In_330,In_459);
xor U212 (N_212,In_735,In_989);
nor U213 (N_213,In_31,In_487);
or U214 (N_214,In_74,In_872);
or U215 (N_215,In_168,In_363);
nand U216 (N_216,In_824,In_920);
or U217 (N_217,In_544,In_996);
or U218 (N_218,In_282,In_202);
or U219 (N_219,In_30,In_23);
xnor U220 (N_220,In_709,In_461);
xnor U221 (N_221,In_225,In_705);
and U222 (N_222,In_976,In_692);
nand U223 (N_223,In_904,In_790);
nand U224 (N_224,In_266,In_301);
nand U225 (N_225,In_218,In_349);
or U226 (N_226,In_131,In_322);
xnor U227 (N_227,In_163,In_338);
xor U228 (N_228,In_333,In_781);
nand U229 (N_229,In_445,In_164);
and U230 (N_230,In_535,In_602);
and U231 (N_231,In_991,In_203);
nand U232 (N_232,In_480,In_146);
nor U233 (N_233,In_831,In_176);
or U234 (N_234,In_538,In_645);
nor U235 (N_235,In_610,In_658);
or U236 (N_236,In_843,In_22);
nand U237 (N_237,In_292,In_542);
or U238 (N_238,In_133,In_992);
nor U239 (N_239,In_321,In_983);
nand U240 (N_240,In_135,In_156);
xor U241 (N_241,In_927,In_412);
nor U242 (N_242,In_721,In_577);
nand U243 (N_243,In_251,In_724);
nand U244 (N_244,In_263,In_138);
and U245 (N_245,In_934,In_813);
nor U246 (N_246,In_443,In_160);
or U247 (N_247,In_166,In_701);
nor U248 (N_248,In_51,In_279);
and U249 (N_249,In_585,In_874);
xnor U250 (N_250,In_640,In_661);
nor U251 (N_251,In_17,In_727);
xnor U252 (N_252,In_250,In_800);
nand U253 (N_253,In_362,In_736);
nor U254 (N_254,In_574,In_875);
and U255 (N_255,In_474,In_937);
or U256 (N_256,In_268,In_590);
nand U257 (N_257,In_54,In_757);
and U258 (N_258,In_520,In_791);
nor U259 (N_259,In_648,In_405);
nand U260 (N_260,In_121,In_64);
and U261 (N_261,In_318,In_201);
nor U262 (N_262,In_632,In_519);
nor U263 (N_263,In_811,In_276);
nand U264 (N_264,In_247,In_484);
xnor U265 (N_265,In_603,In_118);
nand U266 (N_266,In_587,In_812);
nand U267 (N_267,In_890,In_274);
nand U268 (N_268,In_684,In_748);
nand U269 (N_269,In_850,In_55);
and U270 (N_270,In_181,In_158);
or U271 (N_271,In_280,In_770);
nand U272 (N_272,In_561,In_395);
and U273 (N_273,In_458,In_380);
nor U274 (N_274,In_481,In_300);
nor U275 (N_275,In_430,In_560);
or U276 (N_276,In_313,In_895);
nor U277 (N_277,In_220,In_964);
xnor U278 (N_278,In_861,In_919);
xnor U279 (N_279,In_246,In_139);
xor U280 (N_280,In_720,In_534);
xor U281 (N_281,In_581,In_646);
xor U282 (N_282,In_200,In_555);
or U283 (N_283,In_714,In_653);
xor U284 (N_284,In_28,In_657);
xnor U285 (N_285,In_494,In_562);
xnor U286 (N_286,In_364,In_864);
or U287 (N_287,In_382,In_114);
nand U288 (N_288,In_717,In_229);
or U289 (N_289,In_550,In_490);
xor U290 (N_290,In_553,In_921);
and U291 (N_291,In_378,In_36);
and U292 (N_292,In_197,In_387);
or U293 (N_293,In_799,In_456);
xor U294 (N_294,In_592,In_854);
xor U295 (N_295,In_446,In_120);
or U296 (N_296,In_227,In_219);
and U297 (N_297,In_195,In_467);
xnor U298 (N_298,In_87,In_419);
nor U299 (N_299,In_678,In_935);
or U300 (N_300,In_243,In_368);
xor U301 (N_301,In_193,In_169);
or U302 (N_302,In_460,In_971);
and U303 (N_303,In_170,In_105);
nor U304 (N_304,In_190,In_241);
nor U305 (N_305,In_882,In_691);
xnor U306 (N_306,In_410,In_216);
nor U307 (N_307,In_768,In_739);
xor U308 (N_308,In_565,In_336);
and U309 (N_309,In_825,In_986);
and U310 (N_310,In_528,In_571);
xor U311 (N_311,In_814,In_497);
and U312 (N_312,In_651,In_152);
and U313 (N_313,In_713,In_522);
nand U314 (N_314,In_244,In_666);
nand U315 (N_315,In_621,In_315);
xnor U316 (N_316,In_25,In_360);
nor U317 (N_317,In_155,In_403);
xnor U318 (N_318,In_258,In_738);
or U319 (N_319,In_39,In_383);
nor U320 (N_320,In_233,In_916);
or U321 (N_321,In_803,In_119);
nor U322 (N_322,In_865,In_150);
xor U323 (N_323,In_175,In_747);
nor U324 (N_324,In_778,In_760);
or U325 (N_325,In_914,In_809);
nand U326 (N_326,In_188,In_211);
xor U327 (N_327,In_771,In_111);
and U328 (N_328,In_697,In_416);
and U329 (N_329,In_174,In_796);
nor U330 (N_330,In_457,In_347);
xnor U331 (N_331,In_540,In_957);
and U332 (N_332,In_889,In_862);
and U333 (N_333,In_183,In_644);
or U334 (N_334,In_44,In_110);
or U335 (N_335,In_327,In_906);
nand U336 (N_336,In_69,In_465);
nor U337 (N_337,In_424,In_414);
xnor U338 (N_338,In_9,In_515);
and U339 (N_339,In_563,In_421);
or U340 (N_340,In_851,In_543);
or U341 (N_341,In_99,In_259);
and U342 (N_342,In_547,In_679);
nor U343 (N_343,In_784,In_548);
nand U344 (N_344,In_489,In_961);
and U345 (N_345,In_764,In_766);
nand U346 (N_346,In_45,In_787);
or U347 (N_347,In_672,In_83);
nand U348 (N_348,In_429,In_500);
xor U349 (N_349,In_807,In_584);
xor U350 (N_350,In_631,In_501);
nor U351 (N_351,In_21,In_406);
nor U352 (N_352,In_24,In_222);
xor U353 (N_353,In_374,In_685);
nor U354 (N_354,In_217,In_210);
xor U355 (N_355,In_818,In_238);
nand U356 (N_356,In_732,In_972);
nand U357 (N_357,In_994,In_682);
or U358 (N_358,In_837,In_127);
nand U359 (N_359,In_622,In_756);
and U360 (N_360,In_307,In_59);
nor U361 (N_361,In_823,In_984);
and U362 (N_362,In_722,In_89);
or U363 (N_363,In_982,In_353);
xor U364 (N_364,In_725,In_624);
xor U365 (N_365,In_967,In_690);
nor U366 (N_366,In_609,In_371);
nand U367 (N_367,In_953,In_505);
xor U368 (N_368,In_881,In_521);
nor U369 (N_369,In_532,In_731);
nor U370 (N_370,In_297,In_941);
and U371 (N_371,In_167,In_486);
xor U372 (N_372,In_925,In_26);
xor U373 (N_373,In_929,In_619);
nor U374 (N_374,In_912,In_396);
and U375 (N_375,In_761,In_541);
and U376 (N_376,In_84,In_922);
and U377 (N_377,In_272,In_34);
xor U378 (N_378,In_779,In_671);
nand U379 (N_379,In_785,In_208);
nand U380 (N_380,In_863,In_664);
xnor U381 (N_381,In_41,In_558);
nand U382 (N_382,In_359,In_667);
nor U383 (N_383,In_33,In_298);
or U384 (N_384,In_737,In_346);
nand U385 (N_385,In_79,In_335);
or U386 (N_386,In_113,In_235);
or U387 (N_387,In_708,In_482);
nand U388 (N_388,In_750,In_605);
or U389 (N_389,In_783,In_926);
nand U390 (N_390,In_788,In_634);
nor U391 (N_391,In_575,In_394);
nand U392 (N_392,In_463,In_911);
or U393 (N_393,In_798,In_676);
nor U394 (N_394,In_693,In_873);
nor U395 (N_395,In_990,In_551);
nand U396 (N_396,In_572,In_271);
xnor U397 (N_397,In_136,In_367);
and U398 (N_398,In_468,In_171);
nor U399 (N_399,In_126,In_379);
and U400 (N_400,In_767,In_755);
and U401 (N_401,In_752,In_2);
or U402 (N_402,In_623,In_853);
or U403 (N_403,In_777,In_471);
nand U404 (N_404,In_866,In_426);
nor U405 (N_405,In_566,In_80);
or U406 (N_406,In_408,In_413);
xnor U407 (N_407,In_143,In_37);
and U408 (N_408,In_702,In_840);
nand U409 (N_409,In_931,In_142);
or U410 (N_410,In_604,In_794);
xnor U411 (N_411,In_744,In_805);
and U412 (N_412,In_78,In_979);
or U413 (N_413,In_749,In_447);
and U414 (N_414,In_859,In_476);
nor U415 (N_415,In_588,In_16);
nand U416 (N_416,In_841,In_954);
nand U417 (N_417,In_826,In_569);
nand U418 (N_418,In_913,In_723);
nor U419 (N_419,In_695,In_57);
xor U420 (N_420,In_108,In_391);
or U421 (N_421,In_628,In_832);
xor U422 (N_422,In_81,In_213);
xor U423 (N_423,In_19,In_389);
or U424 (N_424,In_730,In_191);
nand U425 (N_425,In_706,In_43);
and U426 (N_426,In_420,In_844);
or U427 (N_427,In_437,In_879);
nor U428 (N_428,In_50,In_85);
and U429 (N_429,In_792,In_549);
nor U430 (N_430,In_774,In_345);
or U431 (N_431,In_92,In_450);
nor U432 (N_432,In_173,In_291);
and U433 (N_433,In_157,In_669);
and U434 (N_434,In_473,In_894);
xor U435 (N_435,In_516,In_3);
nand U436 (N_436,In_773,In_719);
or U437 (N_437,In_652,In_107);
nand U438 (N_438,In_842,In_711);
or U439 (N_439,In_869,In_597);
and U440 (N_440,In_281,In_962);
or U441 (N_441,In_125,In_493);
nand U442 (N_442,In_643,In_306);
xnor U443 (N_443,In_856,In_65);
xor U444 (N_444,In_498,In_819);
nor U445 (N_445,In_275,In_196);
or U446 (N_446,In_38,In_629);
xor U447 (N_447,In_835,In_765);
or U448 (N_448,In_503,In_828);
nor U449 (N_449,In_491,In_323);
nor U450 (N_450,In_390,In_144);
xor U451 (N_451,In_302,In_324);
nor U452 (N_452,In_821,In_199);
nor U453 (N_453,In_903,In_91);
nand U454 (N_454,In_880,In_427);
nor U455 (N_455,In_728,In_192);
and U456 (N_456,In_348,In_303);
xnor U457 (N_457,In_15,In_618);
nand U458 (N_458,In_270,In_898);
nor U459 (N_459,In_149,In_326);
and U460 (N_460,In_100,In_402);
or U461 (N_461,In_10,In_141);
xnor U462 (N_462,In_455,In_963);
and U463 (N_463,In_876,In_58);
xor U464 (N_464,In_959,In_704);
or U465 (N_465,In_182,In_206);
or U466 (N_466,In_472,In_845);
or U467 (N_467,In_277,In_969);
and U468 (N_468,In_256,In_615);
or U469 (N_469,In_392,In_908);
nor U470 (N_470,In_454,In_317);
nor U471 (N_471,In_399,In_422);
nor U472 (N_472,In_453,In_352);
and U473 (N_473,In_207,In_598);
or U474 (N_474,In_101,In_370);
xnor U475 (N_475,In_70,In_236);
nor U476 (N_476,In_924,In_616);
and U477 (N_477,In_309,In_537);
nand U478 (N_478,In_557,In_215);
xor U479 (N_479,In_331,In_795);
nand U480 (N_480,In_888,In_294);
xor U481 (N_481,In_665,In_726);
or U482 (N_482,In_440,In_49);
or U483 (N_483,In_857,In_254);
and U484 (N_484,In_905,In_974);
or U485 (N_485,In_178,In_977);
or U486 (N_486,In_804,In_625);
nand U487 (N_487,In_689,In_285);
or U488 (N_488,In_849,In_151);
and U489 (N_489,In_257,In_582);
nand U490 (N_490,In_373,In_451);
and U491 (N_491,In_67,In_639);
nand U492 (N_492,In_858,In_283);
xor U493 (N_493,In_187,In_526);
nor U494 (N_494,In_177,In_253);
and U495 (N_495,In_734,In_8);
nor U496 (N_496,In_524,In_372);
xnor U497 (N_497,In_740,In_249);
nor U498 (N_498,In_469,In_316);
nand U499 (N_499,In_341,In_365);
nor U500 (N_500,In_198,In_192);
and U501 (N_501,In_647,In_956);
xnor U502 (N_502,In_444,In_603);
and U503 (N_503,In_563,In_365);
nor U504 (N_504,In_708,In_40);
xnor U505 (N_505,In_892,In_843);
xor U506 (N_506,In_633,In_657);
or U507 (N_507,In_620,In_565);
or U508 (N_508,In_22,In_613);
or U509 (N_509,In_4,In_629);
or U510 (N_510,In_529,In_868);
nor U511 (N_511,In_911,In_158);
or U512 (N_512,In_461,In_218);
nand U513 (N_513,In_244,In_984);
nor U514 (N_514,In_643,In_450);
nand U515 (N_515,In_193,In_661);
xor U516 (N_516,In_857,In_730);
or U517 (N_517,In_827,In_53);
nand U518 (N_518,In_204,In_727);
nand U519 (N_519,In_777,In_204);
or U520 (N_520,In_154,In_277);
or U521 (N_521,In_474,In_331);
or U522 (N_522,In_361,In_632);
or U523 (N_523,In_905,In_477);
nor U524 (N_524,In_955,In_162);
nand U525 (N_525,In_600,In_936);
and U526 (N_526,In_344,In_835);
nand U527 (N_527,In_147,In_125);
nand U528 (N_528,In_256,In_722);
xor U529 (N_529,In_137,In_956);
or U530 (N_530,In_920,In_460);
nor U531 (N_531,In_173,In_36);
and U532 (N_532,In_506,In_807);
and U533 (N_533,In_486,In_263);
nor U534 (N_534,In_967,In_882);
xor U535 (N_535,In_727,In_918);
xnor U536 (N_536,In_792,In_126);
nand U537 (N_537,In_292,In_54);
nor U538 (N_538,In_254,In_634);
xnor U539 (N_539,In_125,In_551);
and U540 (N_540,In_969,In_989);
nand U541 (N_541,In_162,In_104);
and U542 (N_542,In_465,In_910);
nand U543 (N_543,In_321,In_11);
nand U544 (N_544,In_553,In_923);
and U545 (N_545,In_496,In_529);
nand U546 (N_546,In_648,In_609);
nand U547 (N_547,In_206,In_223);
xnor U548 (N_548,In_705,In_347);
or U549 (N_549,In_697,In_578);
nor U550 (N_550,In_335,In_551);
nor U551 (N_551,In_232,In_839);
xor U552 (N_552,In_565,In_241);
and U553 (N_553,In_699,In_501);
xnor U554 (N_554,In_713,In_305);
nor U555 (N_555,In_449,In_138);
and U556 (N_556,In_987,In_292);
or U557 (N_557,In_14,In_435);
and U558 (N_558,In_35,In_739);
nand U559 (N_559,In_743,In_139);
or U560 (N_560,In_99,In_701);
or U561 (N_561,In_1,In_893);
nand U562 (N_562,In_264,In_561);
and U563 (N_563,In_134,In_190);
nor U564 (N_564,In_788,In_233);
xnor U565 (N_565,In_672,In_765);
or U566 (N_566,In_242,In_400);
nor U567 (N_567,In_638,In_78);
xnor U568 (N_568,In_700,In_943);
nand U569 (N_569,In_640,In_654);
or U570 (N_570,In_987,In_250);
and U571 (N_571,In_907,In_567);
nand U572 (N_572,In_177,In_48);
nand U573 (N_573,In_765,In_57);
nand U574 (N_574,In_173,In_963);
and U575 (N_575,In_452,In_584);
nand U576 (N_576,In_123,In_992);
nor U577 (N_577,In_676,In_745);
nor U578 (N_578,In_160,In_428);
nor U579 (N_579,In_391,In_886);
and U580 (N_580,In_195,In_184);
xnor U581 (N_581,In_840,In_423);
or U582 (N_582,In_15,In_13);
and U583 (N_583,In_344,In_543);
nor U584 (N_584,In_275,In_87);
nand U585 (N_585,In_287,In_240);
nor U586 (N_586,In_635,In_466);
and U587 (N_587,In_540,In_660);
or U588 (N_588,In_449,In_60);
xnor U589 (N_589,In_411,In_290);
nor U590 (N_590,In_111,In_540);
nor U591 (N_591,In_515,In_41);
nor U592 (N_592,In_599,In_580);
or U593 (N_593,In_227,In_287);
nand U594 (N_594,In_417,In_931);
and U595 (N_595,In_211,In_35);
nor U596 (N_596,In_210,In_271);
nor U597 (N_597,In_707,In_603);
xnor U598 (N_598,In_579,In_959);
nand U599 (N_599,In_344,In_864);
and U600 (N_600,In_694,In_883);
nor U601 (N_601,In_392,In_560);
or U602 (N_602,In_56,In_761);
nand U603 (N_603,In_461,In_162);
and U604 (N_604,In_979,In_86);
xnor U605 (N_605,In_119,In_299);
and U606 (N_606,In_682,In_578);
xnor U607 (N_607,In_597,In_749);
nand U608 (N_608,In_901,In_79);
or U609 (N_609,In_916,In_903);
nor U610 (N_610,In_419,In_25);
nand U611 (N_611,In_574,In_571);
nand U612 (N_612,In_205,In_356);
nor U613 (N_613,In_454,In_513);
and U614 (N_614,In_856,In_960);
nor U615 (N_615,In_168,In_797);
nand U616 (N_616,In_548,In_733);
xor U617 (N_617,In_441,In_966);
nor U618 (N_618,In_427,In_421);
nor U619 (N_619,In_575,In_329);
xnor U620 (N_620,In_812,In_627);
nand U621 (N_621,In_478,In_730);
or U622 (N_622,In_617,In_401);
nand U623 (N_623,In_280,In_752);
or U624 (N_624,In_867,In_884);
nor U625 (N_625,In_913,In_323);
nor U626 (N_626,In_927,In_925);
and U627 (N_627,In_333,In_492);
or U628 (N_628,In_355,In_915);
nand U629 (N_629,In_717,In_207);
and U630 (N_630,In_178,In_905);
and U631 (N_631,In_582,In_267);
xnor U632 (N_632,In_729,In_302);
and U633 (N_633,In_783,In_12);
nor U634 (N_634,In_638,In_315);
xnor U635 (N_635,In_265,In_615);
nor U636 (N_636,In_842,In_661);
nor U637 (N_637,In_655,In_720);
nand U638 (N_638,In_188,In_120);
nand U639 (N_639,In_860,In_423);
xor U640 (N_640,In_514,In_273);
xor U641 (N_641,In_323,In_146);
nor U642 (N_642,In_146,In_898);
nand U643 (N_643,In_972,In_567);
and U644 (N_644,In_427,In_515);
and U645 (N_645,In_11,In_932);
nor U646 (N_646,In_695,In_919);
or U647 (N_647,In_384,In_588);
and U648 (N_648,In_124,In_972);
nand U649 (N_649,In_408,In_738);
or U650 (N_650,In_763,In_393);
and U651 (N_651,In_932,In_269);
nor U652 (N_652,In_544,In_61);
nor U653 (N_653,In_869,In_281);
xor U654 (N_654,In_519,In_316);
and U655 (N_655,In_464,In_387);
nor U656 (N_656,In_735,In_713);
xnor U657 (N_657,In_620,In_548);
and U658 (N_658,In_160,In_695);
or U659 (N_659,In_723,In_410);
nor U660 (N_660,In_662,In_102);
and U661 (N_661,In_849,In_7);
or U662 (N_662,In_667,In_433);
or U663 (N_663,In_600,In_386);
or U664 (N_664,In_937,In_191);
or U665 (N_665,In_112,In_485);
or U666 (N_666,In_570,In_924);
nand U667 (N_667,In_723,In_39);
nor U668 (N_668,In_196,In_27);
nand U669 (N_669,In_532,In_884);
xnor U670 (N_670,In_453,In_959);
nor U671 (N_671,In_454,In_191);
or U672 (N_672,In_25,In_904);
nor U673 (N_673,In_861,In_476);
or U674 (N_674,In_192,In_594);
nor U675 (N_675,In_457,In_19);
nand U676 (N_676,In_497,In_417);
nand U677 (N_677,In_378,In_931);
xnor U678 (N_678,In_22,In_118);
nor U679 (N_679,In_691,In_853);
nand U680 (N_680,In_311,In_785);
or U681 (N_681,In_335,In_720);
xnor U682 (N_682,In_216,In_788);
and U683 (N_683,In_159,In_957);
xnor U684 (N_684,In_519,In_480);
and U685 (N_685,In_283,In_841);
nand U686 (N_686,In_865,In_258);
or U687 (N_687,In_952,In_72);
or U688 (N_688,In_591,In_991);
nor U689 (N_689,In_570,In_297);
and U690 (N_690,In_251,In_737);
nor U691 (N_691,In_998,In_86);
xnor U692 (N_692,In_702,In_719);
and U693 (N_693,In_919,In_535);
xnor U694 (N_694,In_5,In_731);
xnor U695 (N_695,In_974,In_909);
nand U696 (N_696,In_257,In_581);
or U697 (N_697,In_443,In_425);
nor U698 (N_698,In_924,In_906);
xor U699 (N_699,In_178,In_236);
nand U700 (N_700,In_787,In_50);
nand U701 (N_701,In_87,In_901);
nor U702 (N_702,In_128,In_974);
nand U703 (N_703,In_678,In_173);
and U704 (N_704,In_95,In_548);
and U705 (N_705,In_404,In_402);
nand U706 (N_706,In_693,In_935);
nor U707 (N_707,In_195,In_551);
and U708 (N_708,In_270,In_178);
nor U709 (N_709,In_775,In_816);
or U710 (N_710,In_302,In_461);
and U711 (N_711,In_901,In_761);
nand U712 (N_712,In_532,In_846);
xnor U713 (N_713,In_653,In_854);
nor U714 (N_714,In_9,In_872);
or U715 (N_715,In_89,In_569);
xnor U716 (N_716,In_117,In_394);
and U717 (N_717,In_995,In_506);
nand U718 (N_718,In_291,In_569);
or U719 (N_719,In_191,In_612);
nand U720 (N_720,In_79,In_25);
xor U721 (N_721,In_301,In_472);
xnor U722 (N_722,In_667,In_888);
nor U723 (N_723,In_308,In_654);
nand U724 (N_724,In_192,In_196);
or U725 (N_725,In_918,In_907);
or U726 (N_726,In_756,In_886);
nor U727 (N_727,In_838,In_841);
or U728 (N_728,In_2,In_472);
and U729 (N_729,In_490,In_773);
xor U730 (N_730,In_738,In_706);
xnor U731 (N_731,In_427,In_819);
nor U732 (N_732,In_765,In_913);
xor U733 (N_733,In_638,In_142);
nand U734 (N_734,In_947,In_196);
and U735 (N_735,In_299,In_255);
and U736 (N_736,In_97,In_682);
and U737 (N_737,In_721,In_924);
nand U738 (N_738,In_2,In_844);
xnor U739 (N_739,In_360,In_895);
nor U740 (N_740,In_395,In_18);
nand U741 (N_741,In_693,In_884);
xnor U742 (N_742,In_223,In_203);
and U743 (N_743,In_893,In_91);
or U744 (N_744,In_49,In_888);
xnor U745 (N_745,In_524,In_74);
nor U746 (N_746,In_520,In_779);
nand U747 (N_747,In_188,In_97);
nor U748 (N_748,In_507,In_253);
xor U749 (N_749,In_652,In_928);
xnor U750 (N_750,In_575,In_976);
xor U751 (N_751,In_725,In_867);
and U752 (N_752,In_722,In_806);
nor U753 (N_753,In_175,In_818);
xnor U754 (N_754,In_916,In_556);
nor U755 (N_755,In_319,In_629);
and U756 (N_756,In_420,In_186);
and U757 (N_757,In_174,In_295);
nor U758 (N_758,In_11,In_22);
or U759 (N_759,In_523,In_897);
or U760 (N_760,In_769,In_553);
and U761 (N_761,In_895,In_921);
and U762 (N_762,In_214,In_846);
xor U763 (N_763,In_172,In_644);
or U764 (N_764,In_274,In_164);
nand U765 (N_765,In_447,In_38);
or U766 (N_766,In_837,In_502);
xnor U767 (N_767,In_807,In_479);
xnor U768 (N_768,In_26,In_214);
nor U769 (N_769,In_414,In_547);
or U770 (N_770,In_49,In_70);
or U771 (N_771,In_274,In_633);
nand U772 (N_772,In_522,In_466);
xor U773 (N_773,In_813,In_605);
nand U774 (N_774,In_570,In_535);
and U775 (N_775,In_116,In_790);
xor U776 (N_776,In_541,In_360);
or U777 (N_777,In_343,In_452);
and U778 (N_778,In_242,In_489);
nor U779 (N_779,In_834,In_710);
xor U780 (N_780,In_209,In_962);
or U781 (N_781,In_189,In_73);
nor U782 (N_782,In_53,In_344);
nor U783 (N_783,In_358,In_261);
xor U784 (N_784,In_387,In_518);
xor U785 (N_785,In_662,In_49);
and U786 (N_786,In_808,In_945);
nor U787 (N_787,In_131,In_219);
xnor U788 (N_788,In_774,In_561);
xnor U789 (N_789,In_158,In_806);
and U790 (N_790,In_619,In_567);
and U791 (N_791,In_378,In_548);
xor U792 (N_792,In_257,In_402);
xnor U793 (N_793,In_150,In_79);
and U794 (N_794,In_520,In_511);
xor U795 (N_795,In_437,In_101);
or U796 (N_796,In_709,In_676);
and U797 (N_797,In_865,In_201);
and U798 (N_798,In_666,In_976);
nand U799 (N_799,In_225,In_537);
nand U800 (N_800,In_216,In_886);
and U801 (N_801,In_260,In_54);
nor U802 (N_802,In_149,In_935);
nor U803 (N_803,In_430,In_839);
nor U804 (N_804,In_923,In_431);
nor U805 (N_805,In_217,In_268);
nand U806 (N_806,In_393,In_161);
nor U807 (N_807,In_41,In_342);
and U808 (N_808,In_30,In_212);
xnor U809 (N_809,In_280,In_604);
xor U810 (N_810,In_41,In_193);
or U811 (N_811,In_298,In_149);
or U812 (N_812,In_880,In_642);
nand U813 (N_813,In_84,In_425);
and U814 (N_814,In_94,In_441);
or U815 (N_815,In_878,In_58);
xor U816 (N_816,In_201,In_886);
or U817 (N_817,In_662,In_863);
or U818 (N_818,In_56,In_563);
nor U819 (N_819,In_692,In_775);
or U820 (N_820,In_944,In_164);
xnor U821 (N_821,In_540,In_604);
nand U822 (N_822,In_479,In_529);
nand U823 (N_823,In_516,In_842);
nor U824 (N_824,In_906,In_578);
nand U825 (N_825,In_82,In_997);
and U826 (N_826,In_969,In_906);
or U827 (N_827,In_796,In_399);
xor U828 (N_828,In_116,In_134);
nand U829 (N_829,In_823,In_165);
xor U830 (N_830,In_63,In_315);
and U831 (N_831,In_559,In_624);
xnor U832 (N_832,In_257,In_810);
or U833 (N_833,In_200,In_893);
xnor U834 (N_834,In_35,In_150);
or U835 (N_835,In_843,In_26);
nor U836 (N_836,In_361,In_133);
nor U837 (N_837,In_156,In_280);
and U838 (N_838,In_711,In_750);
nand U839 (N_839,In_828,In_497);
or U840 (N_840,In_926,In_668);
nand U841 (N_841,In_921,In_564);
or U842 (N_842,In_955,In_279);
and U843 (N_843,In_770,In_894);
xnor U844 (N_844,In_94,In_417);
xor U845 (N_845,In_833,In_390);
nor U846 (N_846,In_91,In_42);
nand U847 (N_847,In_485,In_164);
nand U848 (N_848,In_413,In_72);
and U849 (N_849,In_52,In_922);
xnor U850 (N_850,In_788,In_677);
and U851 (N_851,In_903,In_67);
nand U852 (N_852,In_127,In_897);
xor U853 (N_853,In_685,In_756);
xor U854 (N_854,In_692,In_585);
and U855 (N_855,In_17,In_747);
nand U856 (N_856,In_471,In_597);
nand U857 (N_857,In_447,In_248);
and U858 (N_858,In_925,In_696);
xnor U859 (N_859,In_269,In_692);
nor U860 (N_860,In_637,In_738);
xor U861 (N_861,In_102,In_465);
xor U862 (N_862,In_19,In_894);
nand U863 (N_863,In_349,In_533);
nand U864 (N_864,In_957,In_832);
nand U865 (N_865,In_4,In_380);
or U866 (N_866,In_524,In_773);
nand U867 (N_867,In_848,In_13);
or U868 (N_868,In_745,In_284);
nand U869 (N_869,In_123,In_971);
nor U870 (N_870,In_20,In_318);
or U871 (N_871,In_191,In_766);
or U872 (N_872,In_331,In_850);
nor U873 (N_873,In_860,In_532);
xnor U874 (N_874,In_757,In_46);
xor U875 (N_875,In_978,In_19);
and U876 (N_876,In_779,In_343);
and U877 (N_877,In_793,In_829);
xnor U878 (N_878,In_69,In_794);
xnor U879 (N_879,In_545,In_763);
nand U880 (N_880,In_332,In_806);
xnor U881 (N_881,In_131,In_414);
nor U882 (N_882,In_583,In_854);
nand U883 (N_883,In_990,In_800);
nor U884 (N_884,In_233,In_58);
xor U885 (N_885,In_34,In_529);
xnor U886 (N_886,In_849,In_688);
xor U887 (N_887,In_987,In_368);
nor U888 (N_888,In_559,In_46);
or U889 (N_889,In_469,In_391);
or U890 (N_890,In_81,In_463);
or U891 (N_891,In_48,In_598);
and U892 (N_892,In_511,In_939);
nor U893 (N_893,In_993,In_493);
nor U894 (N_894,In_55,In_701);
nand U895 (N_895,In_417,In_381);
nor U896 (N_896,In_771,In_86);
and U897 (N_897,In_984,In_767);
nand U898 (N_898,In_431,In_54);
nor U899 (N_899,In_173,In_887);
nand U900 (N_900,In_389,In_678);
nand U901 (N_901,In_868,In_20);
nor U902 (N_902,In_338,In_27);
xor U903 (N_903,In_988,In_431);
nand U904 (N_904,In_885,In_149);
or U905 (N_905,In_109,In_665);
nor U906 (N_906,In_125,In_291);
nand U907 (N_907,In_578,In_903);
nor U908 (N_908,In_264,In_12);
and U909 (N_909,In_962,In_801);
nor U910 (N_910,In_528,In_567);
and U911 (N_911,In_172,In_370);
and U912 (N_912,In_257,In_635);
xor U913 (N_913,In_446,In_506);
nand U914 (N_914,In_811,In_822);
nand U915 (N_915,In_20,In_703);
xnor U916 (N_916,In_50,In_850);
and U917 (N_917,In_466,In_755);
nor U918 (N_918,In_512,In_490);
nor U919 (N_919,In_725,In_729);
nor U920 (N_920,In_909,In_311);
nand U921 (N_921,In_701,In_498);
and U922 (N_922,In_793,In_763);
and U923 (N_923,In_328,In_210);
or U924 (N_924,In_875,In_872);
xnor U925 (N_925,In_462,In_618);
and U926 (N_926,In_386,In_68);
nand U927 (N_927,In_917,In_642);
nand U928 (N_928,In_722,In_933);
xor U929 (N_929,In_291,In_11);
or U930 (N_930,In_41,In_968);
nand U931 (N_931,In_488,In_769);
or U932 (N_932,In_743,In_963);
and U933 (N_933,In_326,In_765);
and U934 (N_934,In_230,In_381);
and U935 (N_935,In_551,In_389);
and U936 (N_936,In_343,In_582);
and U937 (N_937,In_429,In_840);
xnor U938 (N_938,In_152,In_453);
or U939 (N_939,In_519,In_664);
or U940 (N_940,In_228,In_191);
or U941 (N_941,In_303,In_715);
or U942 (N_942,In_398,In_895);
nor U943 (N_943,In_685,In_909);
and U944 (N_944,In_22,In_383);
nand U945 (N_945,In_121,In_795);
xnor U946 (N_946,In_215,In_131);
nand U947 (N_947,In_567,In_854);
nand U948 (N_948,In_267,In_506);
or U949 (N_949,In_659,In_921);
xnor U950 (N_950,In_631,In_206);
and U951 (N_951,In_504,In_942);
xnor U952 (N_952,In_327,In_711);
or U953 (N_953,In_631,In_604);
nand U954 (N_954,In_542,In_376);
xnor U955 (N_955,In_332,In_979);
nor U956 (N_956,In_592,In_751);
or U957 (N_957,In_468,In_188);
or U958 (N_958,In_284,In_3);
or U959 (N_959,In_506,In_991);
or U960 (N_960,In_641,In_600);
or U961 (N_961,In_988,In_725);
or U962 (N_962,In_198,In_406);
xnor U963 (N_963,In_840,In_18);
nand U964 (N_964,In_353,In_430);
and U965 (N_965,In_568,In_231);
nor U966 (N_966,In_402,In_448);
xnor U967 (N_967,In_656,In_531);
xor U968 (N_968,In_817,In_643);
nor U969 (N_969,In_614,In_804);
nor U970 (N_970,In_478,In_68);
nor U971 (N_971,In_827,In_724);
or U972 (N_972,In_73,In_566);
nor U973 (N_973,In_929,In_184);
and U974 (N_974,In_34,In_478);
and U975 (N_975,In_566,In_141);
xnor U976 (N_976,In_5,In_240);
nor U977 (N_977,In_370,In_247);
or U978 (N_978,In_813,In_236);
nor U979 (N_979,In_360,In_386);
xnor U980 (N_980,In_381,In_993);
nor U981 (N_981,In_286,In_199);
xnor U982 (N_982,In_36,In_206);
nand U983 (N_983,In_333,In_587);
nor U984 (N_984,In_960,In_441);
and U985 (N_985,In_580,In_452);
nand U986 (N_986,In_277,In_495);
nand U987 (N_987,In_766,In_893);
or U988 (N_988,In_719,In_636);
nor U989 (N_989,In_195,In_7);
and U990 (N_990,In_389,In_920);
or U991 (N_991,In_256,In_999);
or U992 (N_992,In_254,In_497);
xor U993 (N_993,In_552,In_550);
xor U994 (N_994,In_173,In_663);
or U995 (N_995,In_387,In_706);
and U996 (N_996,In_364,In_499);
xor U997 (N_997,In_575,In_573);
and U998 (N_998,In_995,In_320);
nor U999 (N_999,In_299,In_684);
nand U1000 (N_1000,In_36,In_361);
nand U1001 (N_1001,In_452,In_412);
nand U1002 (N_1002,In_158,In_835);
or U1003 (N_1003,In_227,In_707);
or U1004 (N_1004,In_711,In_500);
nor U1005 (N_1005,In_815,In_761);
nand U1006 (N_1006,In_75,In_187);
nand U1007 (N_1007,In_118,In_253);
xor U1008 (N_1008,In_155,In_283);
nand U1009 (N_1009,In_706,In_109);
nor U1010 (N_1010,In_666,In_278);
nand U1011 (N_1011,In_160,In_431);
xor U1012 (N_1012,In_607,In_504);
and U1013 (N_1013,In_964,In_46);
and U1014 (N_1014,In_630,In_684);
and U1015 (N_1015,In_8,In_84);
or U1016 (N_1016,In_982,In_292);
nor U1017 (N_1017,In_283,In_661);
nand U1018 (N_1018,In_828,In_28);
and U1019 (N_1019,In_812,In_616);
and U1020 (N_1020,In_53,In_339);
xnor U1021 (N_1021,In_742,In_835);
and U1022 (N_1022,In_819,In_86);
nor U1023 (N_1023,In_823,In_967);
or U1024 (N_1024,In_627,In_274);
nor U1025 (N_1025,In_854,In_614);
or U1026 (N_1026,In_928,In_424);
nand U1027 (N_1027,In_780,In_226);
or U1028 (N_1028,In_275,In_159);
xnor U1029 (N_1029,In_112,In_363);
and U1030 (N_1030,In_977,In_902);
nand U1031 (N_1031,In_462,In_780);
and U1032 (N_1032,In_310,In_464);
xor U1033 (N_1033,In_720,In_600);
nor U1034 (N_1034,In_397,In_48);
nor U1035 (N_1035,In_786,In_810);
nor U1036 (N_1036,In_154,In_189);
nand U1037 (N_1037,In_928,In_400);
or U1038 (N_1038,In_35,In_18);
nor U1039 (N_1039,In_5,In_815);
and U1040 (N_1040,In_402,In_18);
nand U1041 (N_1041,In_359,In_238);
nor U1042 (N_1042,In_410,In_55);
and U1043 (N_1043,In_175,In_95);
nand U1044 (N_1044,In_451,In_363);
or U1045 (N_1045,In_929,In_842);
and U1046 (N_1046,In_127,In_514);
or U1047 (N_1047,In_755,In_134);
xnor U1048 (N_1048,In_601,In_538);
and U1049 (N_1049,In_225,In_752);
nand U1050 (N_1050,In_241,In_408);
and U1051 (N_1051,In_270,In_276);
nand U1052 (N_1052,In_597,In_692);
or U1053 (N_1053,In_465,In_674);
nor U1054 (N_1054,In_346,In_303);
nand U1055 (N_1055,In_714,In_46);
xor U1056 (N_1056,In_359,In_685);
or U1057 (N_1057,In_464,In_891);
or U1058 (N_1058,In_175,In_22);
or U1059 (N_1059,In_358,In_79);
nand U1060 (N_1060,In_381,In_292);
nor U1061 (N_1061,In_708,In_792);
or U1062 (N_1062,In_930,In_348);
nand U1063 (N_1063,In_577,In_953);
xor U1064 (N_1064,In_725,In_676);
or U1065 (N_1065,In_813,In_747);
nor U1066 (N_1066,In_332,In_972);
nor U1067 (N_1067,In_277,In_997);
nor U1068 (N_1068,In_792,In_969);
or U1069 (N_1069,In_850,In_233);
and U1070 (N_1070,In_271,In_397);
nand U1071 (N_1071,In_440,In_6);
xnor U1072 (N_1072,In_727,In_964);
or U1073 (N_1073,In_992,In_406);
and U1074 (N_1074,In_699,In_958);
and U1075 (N_1075,In_336,In_747);
nor U1076 (N_1076,In_855,In_599);
xor U1077 (N_1077,In_666,In_476);
or U1078 (N_1078,In_596,In_214);
nor U1079 (N_1079,In_877,In_442);
or U1080 (N_1080,In_707,In_40);
and U1081 (N_1081,In_511,In_591);
xnor U1082 (N_1082,In_770,In_199);
nand U1083 (N_1083,In_165,In_960);
nand U1084 (N_1084,In_913,In_382);
or U1085 (N_1085,In_821,In_791);
nor U1086 (N_1086,In_31,In_14);
nor U1087 (N_1087,In_222,In_374);
or U1088 (N_1088,In_661,In_844);
or U1089 (N_1089,In_589,In_677);
nand U1090 (N_1090,In_692,In_400);
and U1091 (N_1091,In_951,In_638);
nand U1092 (N_1092,In_209,In_871);
and U1093 (N_1093,In_586,In_303);
or U1094 (N_1094,In_641,In_40);
or U1095 (N_1095,In_287,In_412);
and U1096 (N_1096,In_64,In_103);
or U1097 (N_1097,In_907,In_657);
nor U1098 (N_1098,In_581,In_404);
and U1099 (N_1099,In_328,In_139);
or U1100 (N_1100,In_376,In_884);
or U1101 (N_1101,In_558,In_73);
and U1102 (N_1102,In_398,In_216);
xnor U1103 (N_1103,In_476,In_240);
nand U1104 (N_1104,In_322,In_103);
xnor U1105 (N_1105,In_698,In_193);
nor U1106 (N_1106,In_871,In_846);
and U1107 (N_1107,In_476,In_948);
xnor U1108 (N_1108,In_761,In_974);
xnor U1109 (N_1109,In_245,In_96);
nand U1110 (N_1110,In_841,In_549);
or U1111 (N_1111,In_158,In_215);
nand U1112 (N_1112,In_693,In_834);
and U1113 (N_1113,In_882,In_529);
xnor U1114 (N_1114,In_888,In_731);
xor U1115 (N_1115,In_190,In_207);
and U1116 (N_1116,In_823,In_971);
nand U1117 (N_1117,In_220,In_881);
nor U1118 (N_1118,In_1,In_286);
xnor U1119 (N_1119,In_140,In_527);
or U1120 (N_1120,In_47,In_1);
and U1121 (N_1121,In_125,In_959);
and U1122 (N_1122,In_410,In_856);
and U1123 (N_1123,In_556,In_312);
and U1124 (N_1124,In_228,In_27);
and U1125 (N_1125,In_22,In_865);
nand U1126 (N_1126,In_424,In_523);
or U1127 (N_1127,In_953,In_712);
or U1128 (N_1128,In_979,In_512);
xnor U1129 (N_1129,In_665,In_729);
nand U1130 (N_1130,In_0,In_929);
nor U1131 (N_1131,In_751,In_701);
nor U1132 (N_1132,In_482,In_378);
and U1133 (N_1133,In_582,In_111);
nor U1134 (N_1134,In_28,In_154);
and U1135 (N_1135,In_659,In_850);
or U1136 (N_1136,In_903,In_368);
and U1137 (N_1137,In_745,In_241);
nor U1138 (N_1138,In_979,In_845);
and U1139 (N_1139,In_595,In_101);
nor U1140 (N_1140,In_961,In_73);
or U1141 (N_1141,In_717,In_571);
nor U1142 (N_1142,In_199,In_499);
nand U1143 (N_1143,In_463,In_785);
xnor U1144 (N_1144,In_335,In_310);
or U1145 (N_1145,In_506,In_128);
xnor U1146 (N_1146,In_262,In_928);
and U1147 (N_1147,In_544,In_641);
nor U1148 (N_1148,In_886,In_530);
nor U1149 (N_1149,In_288,In_932);
nand U1150 (N_1150,In_70,In_118);
and U1151 (N_1151,In_204,In_296);
nand U1152 (N_1152,In_964,In_184);
nor U1153 (N_1153,In_863,In_256);
nor U1154 (N_1154,In_556,In_272);
xnor U1155 (N_1155,In_836,In_819);
nand U1156 (N_1156,In_718,In_683);
or U1157 (N_1157,In_580,In_188);
or U1158 (N_1158,In_962,In_446);
or U1159 (N_1159,In_433,In_707);
and U1160 (N_1160,In_234,In_171);
or U1161 (N_1161,In_710,In_532);
xnor U1162 (N_1162,In_211,In_613);
nor U1163 (N_1163,In_791,In_926);
nor U1164 (N_1164,In_990,In_447);
xor U1165 (N_1165,In_462,In_981);
and U1166 (N_1166,In_922,In_598);
nor U1167 (N_1167,In_811,In_360);
and U1168 (N_1168,In_779,In_477);
or U1169 (N_1169,In_35,In_368);
and U1170 (N_1170,In_83,In_575);
or U1171 (N_1171,In_719,In_541);
or U1172 (N_1172,In_544,In_581);
xnor U1173 (N_1173,In_122,In_256);
or U1174 (N_1174,In_224,In_274);
nor U1175 (N_1175,In_679,In_930);
nor U1176 (N_1176,In_4,In_278);
nand U1177 (N_1177,In_629,In_79);
and U1178 (N_1178,In_837,In_93);
xnor U1179 (N_1179,In_491,In_657);
or U1180 (N_1180,In_289,In_345);
nand U1181 (N_1181,In_393,In_42);
and U1182 (N_1182,In_568,In_782);
and U1183 (N_1183,In_274,In_157);
nand U1184 (N_1184,In_757,In_591);
and U1185 (N_1185,In_494,In_935);
or U1186 (N_1186,In_452,In_651);
nor U1187 (N_1187,In_460,In_143);
nand U1188 (N_1188,In_561,In_517);
nor U1189 (N_1189,In_776,In_464);
and U1190 (N_1190,In_268,In_129);
xnor U1191 (N_1191,In_719,In_235);
and U1192 (N_1192,In_740,In_773);
and U1193 (N_1193,In_941,In_255);
nand U1194 (N_1194,In_332,In_158);
nor U1195 (N_1195,In_589,In_928);
nand U1196 (N_1196,In_463,In_577);
xor U1197 (N_1197,In_600,In_652);
or U1198 (N_1198,In_834,In_969);
nor U1199 (N_1199,In_897,In_372);
nand U1200 (N_1200,In_932,In_534);
nor U1201 (N_1201,In_113,In_930);
nor U1202 (N_1202,In_223,In_368);
nand U1203 (N_1203,In_366,In_576);
xnor U1204 (N_1204,In_970,In_535);
and U1205 (N_1205,In_526,In_634);
nand U1206 (N_1206,In_803,In_756);
nand U1207 (N_1207,In_675,In_194);
xnor U1208 (N_1208,In_270,In_58);
nand U1209 (N_1209,In_331,In_198);
xnor U1210 (N_1210,In_994,In_468);
or U1211 (N_1211,In_866,In_65);
or U1212 (N_1212,In_114,In_86);
and U1213 (N_1213,In_117,In_82);
nor U1214 (N_1214,In_7,In_742);
xor U1215 (N_1215,In_246,In_704);
or U1216 (N_1216,In_976,In_294);
xnor U1217 (N_1217,In_291,In_422);
or U1218 (N_1218,In_875,In_961);
and U1219 (N_1219,In_434,In_920);
nor U1220 (N_1220,In_80,In_78);
xor U1221 (N_1221,In_368,In_503);
nor U1222 (N_1222,In_766,In_918);
and U1223 (N_1223,In_822,In_4);
and U1224 (N_1224,In_634,In_938);
nand U1225 (N_1225,In_239,In_171);
or U1226 (N_1226,In_435,In_737);
xnor U1227 (N_1227,In_744,In_443);
or U1228 (N_1228,In_253,In_682);
nor U1229 (N_1229,In_207,In_485);
and U1230 (N_1230,In_927,In_124);
xor U1231 (N_1231,In_844,In_241);
nand U1232 (N_1232,In_996,In_574);
and U1233 (N_1233,In_924,In_834);
nand U1234 (N_1234,In_850,In_599);
nor U1235 (N_1235,In_181,In_355);
xor U1236 (N_1236,In_156,In_450);
nand U1237 (N_1237,In_192,In_858);
and U1238 (N_1238,In_270,In_998);
xor U1239 (N_1239,In_194,In_540);
xor U1240 (N_1240,In_477,In_253);
xor U1241 (N_1241,In_291,In_617);
xnor U1242 (N_1242,In_96,In_809);
nor U1243 (N_1243,In_72,In_285);
nor U1244 (N_1244,In_775,In_288);
xor U1245 (N_1245,In_58,In_37);
or U1246 (N_1246,In_428,In_101);
nor U1247 (N_1247,In_691,In_803);
xor U1248 (N_1248,In_336,In_638);
nand U1249 (N_1249,In_121,In_679);
nor U1250 (N_1250,In_902,In_974);
nand U1251 (N_1251,In_769,In_137);
nor U1252 (N_1252,In_65,In_32);
nand U1253 (N_1253,In_914,In_46);
xnor U1254 (N_1254,In_104,In_257);
xnor U1255 (N_1255,In_329,In_767);
and U1256 (N_1256,In_376,In_826);
or U1257 (N_1257,In_658,In_748);
nor U1258 (N_1258,In_518,In_425);
xnor U1259 (N_1259,In_509,In_839);
nand U1260 (N_1260,In_45,In_578);
or U1261 (N_1261,In_396,In_537);
nand U1262 (N_1262,In_564,In_941);
and U1263 (N_1263,In_733,In_417);
nand U1264 (N_1264,In_405,In_349);
xor U1265 (N_1265,In_163,In_120);
nand U1266 (N_1266,In_810,In_916);
or U1267 (N_1267,In_477,In_724);
xor U1268 (N_1268,In_436,In_100);
and U1269 (N_1269,In_788,In_771);
or U1270 (N_1270,In_169,In_876);
and U1271 (N_1271,In_94,In_708);
nand U1272 (N_1272,In_928,In_116);
or U1273 (N_1273,In_808,In_72);
nand U1274 (N_1274,In_576,In_662);
xor U1275 (N_1275,In_195,In_858);
nand U1276 (N_1276,In_93,In_402);
nor U1277 (N_1277,In_716,In_342);
nor U1278 (N_1278,In_559,In_774);
xnor U1279 (N_1279,In_666,In_263);
nor U1280 (N_1280,In_717,In_405);
nand U1281 (N_1281,In_654,In_556);
nand U1282 (N_1282,In_196,In_588);
or U1283 (N_1283,In_939,In_370);
or U1284 (N_1284,In_292,In_506);
and U1285 (N_1285,In_439,In_728);
nand U1286 (N_1286,In_718,In_583);
and U1287 (N_1287,In_820,In_42);
xor U1288 (N_1288,In_31,In_505);
nor U1289 (N_1289,In_442,In_804);
nor U1290 (N_1290,In_870,In_319);
nand U1291 (N_1291,In_139,In_554);
or U1292 (N_1292,In_494,In_377);
nor U1293 (N_1293,In_10,In_52);
xor U1294 (N_1294,In_51,In_713);
or U1295 (N_1295,In_527,In_609);
nand U1296 (N_1296,In_168,In_322);
xor U1297 (N_1297,In_27,In_221);
xor U1298 (N_1298,In_629,In_632);
nor U1299 (N_1299,In_780,In_665);
nor U1300 (N_1300,In_1,In_172);
nor U1301 (N_1301,In_717,In_880);
nand U1302 (N_1302,In_844,In_858);
xor U1303 (N_1303,In_727,In_961);
or U1304 (N_1304,In_384,In_168);
or U1305 (N_1305,In_492,In_881);
and U1306 (N_1306,In_29,In_3);
nor U1307 (N_1307,In_226,In_914);
nand U1308 (N_1308,In_262,In_788);
nand U1309 (N_1309,In_872,In_518);
xnor U1310 (N_1310,In_647,In_359);
nor U1311 (N_1311,In_911,In_450);
or U1312 (N_1312,In_202,In_321);
nand U1313 (N_1313,In_863,In_997);
and U1314 (N_1314,In_224,In_301);
and U1315 (N_1315,In_850,In_601);
and U1316 (N_1316,In_724,In_646);
nor U1317 (N_1317,In_874,In_987);
nand U1318 (N_1318,In_405,In_63);
or U1319 (N_1319,In_477,In_381);
or U1320 (N_1320,In_383,In_509);
nand U1321 (N_1321,In_66,In_753);
nand U1322 (N_1322,In_799,In_120);
or U1323 (N_1323,In_26,In_945);
or U1324 (N_1324,In_367,In_854);
or U1325 (N_1325,In_684,In_627);
or U1326 (N_1326,In_498,In_974);
xor U1327 (N_1327,In_964,In_278);
and U1328 (N_1328,In_879,In_643);
or U1329 (N_1329,In_249,In_357);
nor U1330 (N_1330,In_371,In_839);
xor U1331 (N_1331,In_67,In_141);
nor U1332 (N_1332,In_786,In_370);
xnor U1333 (N_1333,In_288,In_436);
or U1334 (N_1334,In_807,In_966);
or U1335 (N_1335,In_329,In_235);
nand U1336 (N_1336,In_438,In_348);
or U1337 (N_1337,In_458,In_805);
nor U1338 (N_1338,In_419,In_136);
nor U1339 (N_1339,In_582,In_211);
nand U1340 (N_1340,In_162,In_159);
or U1341 (N_1341,In_394,In_2);
nand U1342 (N_1342,In_470,In_192);
or U1343 (N_1343,In_16,In_60);
or U1344 (N_1344,In_89,In_921);
nand U1345 (N_1345,In_863,In_66);
nand U1346 (N_1346,In_906,In_346);
xnor U1347 (N_1347,In_503,In_965);
nor U1348 (N_1348,In_780,In_785);
xnor U1349 (N_1349,In_562,In_142);
and U1350 (N_1350,In_986,In_34);
nand U1351 (N_1351,In_992,In_25);
xor U1352 (N_1352,In_207,In_348);
nor U1353 (N_1353,In_72,In_60);
and U1354 (N_1354,In_674,In_531);
nand U1355 (N_1355,In_955,In_515);
nand U1356 (N_1356,In_207,In_526);
and U1357 (N_1357,In_907,In_467);
xor U1358 (N_1358,In_762,In_190);
and U1359 (N_1359,In_699,In_34);
xor U1360 (N_1360,In_823,In_191);
xnor U1361 (N_1361,In_53,In_98);
and U1362 (N_1362,In_689,In_172);
xnor U1363 (N_1363,In_990,In_492);
xnor U1364 (N_1364,In_50,In_686);
or U1365 (N_1365,In_932,In_420);
nand U1366 (N_1366,In_741,In_272);
or U1367 (N_1367,In_732,In_332);
and U1368 (N_1368,In_58,In_955);
nand U1369 (N_1369,In_823,In_961);
or U1370 (N_1370,In_733,In_673);
or U1371 (N_1371,In_864,In_911);
and U1372 (N_1372,In_985,In_321);
xnor U1373 (N_1373,In_53,In_875);
xnor U1374 (N_1374,In_613,In_12);
nand U1375 (N_1375,In_516,In_73);
nor U1376 (N_1376,In_484,In_190);
nand U1377 (N_1377,In_736,In_797);
or U1378 (N_1378,In_888,In_430);
nor U1379 (N_1379,In_799,In_379);
xnor U1380 (N_1380,In_938,In_622);
nor U1381 (N_1381,In_464,In_448);
or U1382 (N_1382,In_936,In_337);
or U1383 (N_1383,In_678,In_429);
or U1384 (N_1384,In_828,In_737);
nor U1385 (N_1385,In_935,In_606);
nand U1386 (N_1386,In_696,In_247);
nor U1387 (N_1387,In_621,In_926);
xor U1388 (N_1388,In_323,In_553);
or U1389 (N_1389,In_353,In_270);
and U1390 (N_1390,In_166,In_322);
nand U1391 (N_1391,In_210,In_755);
or U1392 (N_1392,In_876,In_365);
nor U1393 (N_1393,In_797,In_469);
or U1394 (N_1394,In_691,In_748);
nor U1395 (N_1395,In_340,In_929);
or U1396 (N_1396,In_742,In_897);
or U1397 (N_1397,In_920,In_681);
nor U1398 (N_1398,In_599,In_530);
and U1399 (N_1399,In_589,In_675);
and U1400 (N_1400,In_373,In_325);
nor U1401 (N_1401,In_559,In_414);
xnor U1402 (N_1402,In_211,In_782);
or U1403 (N_1403,In_297,In_668);
xor U1404 (N_1404,In_618,In_221);
nand U1405 (N_1405,In_48,In_591);
xor U1406 (N_1406,In_687,In_401);
nor U1407 (N_1407,In_963,In_276);
nor U1408 (N_1408,In_622,In_481);
nor U1409 (N_1409,In_380,In_45);
nand U1410 (N_1410,In_953,In_445);
nor U1411 (N_1411,In_57,In_549);
nand U1412 (N_1412,In_555,In_348);
xnor U1413 (N_1413,In_98,In_578);
and U1414 (N_1414,In_277,In_270);
nor U1415 (N_1415,In_972,In_941);
or U1416 (N_1416,In_7,In_667);
xnor U1417 (N_1417,In_706,In_538);
and U1418 (N_1418,In_495,In_232);
xor U1419 (N_1419,In_886,In_813);
and U1420 (N_1420,In_648,In_310);
nand U1421 (N_1421,In_351,In_629);
nand U1422 (N_1422,In_913,In_718);
nand U1423 (N_1423,In_265,In_77);
nor U1424 (N_1424,In_926,In_777);
nand U1425 (N_1425,In_754,In_846);
and U1426 (N_1426,In_254,In_478);
xor U1427 (N_1427,In_976,In_704);
nand U1428 (N_1428,In_260,In_711);
xor U1429 (N_1429,In_646,In_704);
xor U1430 (N_1430,In_497,In_706);
and U1431 (N_1431,In_56,In_913);
or U1432 (N_1432,In_990,In_980);
or U1433 (N_1433,In_852,In_238);
and U1434 (N_1434,In_431,In_119);
or U1435 (N_1435,In_47,In_992);
and U1436 (N_1436,In_41,In_333);
or U1437 (N_1437,In_315,In_190);
nand U1438 (N_1438,In_980,In_787);
and U1439 (N_1439,In_242,In_31);
nand U1440 (N_1440,In_374,In_415);
or U1441 (N_1441,In_819,In_202);
and U1442 (N_1442,In_879,In_673);
nand U1443 (N_1443,In_561,In_27);
nand U1444 (N_1444,In_561,In_138);
nand U1445 (N_1445,In_969,In_466);
and U1446 (N_1446,In_911,In_119);
xnor U1447 (N_1447,In_41,In_241);
and U1448 (N_1448,In_496,In_388);
xnor U1449 (N_1449,In_272,In_820);
and U1450 (N_1450,In_310,In_928);
and U1451 (N_1451,In_829,In_247);
nand U1452 (N_1452,In_866,In_733);
xnor U1453 (N_1453,In_78,In_928);
nand U1454 (N_1454,In_299,In_157);
nand U1455 (N_1455,In_988,In_986);
or U1456 (N_1456,In_105,In_930);
and U1457 (N_1457,In_637,In_696);
or U1458 (N_1458,In_440,In_291);
xor U1459 (N_1459,In_980,In_410);
and U1460 (N_1460,In_979,In_286);
nor U1461 (N_1461,In_933,In_451);
or U1462 (N_1462,In_542,In_9);
or U1463 (N_1463,In_535,In_138);
nor U1464 (N_1464,In_46,In_823);
nand U1465 (N_1465,In_938,In_407);
nand U1466 (N_1466,In_368,In_442);
or U1467 (N_1467,In_30,In_675);
and U1468 (N_1468,In_422,In_492);
or U1469 (N_1469,In_981,In_360);
and U1470 (N_1470,In_324,In_989);
xnor U1471 (N_1471,In_930,In_369);
and U1472 (N_1472,In_690,In_952);
xor U1473 (N_1473,In_520,In_409);
or U1474 (N_1474,In_316,In_745);
xnor U1475 (N_1475,In_673,In_302);
and U1476 (N_1476,In_411,In_844);
and U1477 (N_1477,In_197,In_663);
and U1478 (N_1478,In_598,In_64);
xnor U1479 (N_1479,In_471,In_681);
xnor U1480 (N_1480,In_815,In_182);
nor U1481 (N_1481,In_457,In_796);
xnor U1482 (N_1482,In_961,In_47);
nor U1483 (N_1483,In_599,In_404);
nand U1484 (N_1484,In_227,In_438);
xnor U1485 (N_1485,In_825,In_806);
nand U1486 (N_1486,In_715,In_946);
nand U1487 (N_1487,In_103,In_489);
nor U1488 (N_1488,In_840,In_376);
xor U1489 (N_1489,In_371,In_108);
nor U1490 (N_1490,In_889,In_740);
nand U1491 (N_1491,In_545,In_397);
nand U1492 (N_1492,In_120,In_166);
and U1493 (N_1493,In_316,In_187);
nor U1494 (N_1494,In_341,In_839);
nand U1495 (N_1495,In_251,In_610);
and U1496 (N_1496,In_127,In_292);
xnor U1497 (N_1497,In_113,In_605);
nor U1498 (N_1498,In_263,In_324);
or U1499 (N_1499,In_589,In_133);
nand U1500 (N_1500,In_919,In_686);
and U1501 (N_1501,In_329,In_279);
or U1502 (N_1502,In_988,In_188);
xor U1503 (N_1503,In_985,In_393);
and U1504 (N_1504,In_278,In_335);
nor U1505 (N_1505,In_509,In_53);
nor U1506 (N_1506,In_242,In_696);
nand U1507 (N_1507,In_820,In_523);
or U1508 (N_1508,In_868,In_768);
or U1509 (N_1509,In_361,In_298);
or U1510 (N_1510,In_456,In_584);
nor U1511 (N_1511,In_46,In_548);
xnor U1512 (N_1512,In_704,In_472);
and U1513 (N_1513,In_517,In_835);
or U1514 (N_1514,In_891,In_362);
xnor U1515 (N_1515,In_200,In_303);
xnor U1516 (N_1516,In_442,In_371);
or U1517 (N_1517,In_973,In_958);
and U1518 (N_1518,In_128,In_188);
nor U1519 (N_1519,In_192,In_259);
nor U1520 (N_1520,In_384,In_632);
nand U1521 (N_1521,In_344,In_113);
xor U1522 (N_1522,In_178,In_528);
and U1523 (N_1523,In_274,In_898);
nand U1524 (N_1524,In_496,In_385);
and U1525 (N_1525,In_692,In_227);
nor U1526 (N_1526,In_774,In_159);
or U1527 (N_1527,In_414,In_240);
and U1528 (N_1528,In_262,In_398);
nor U1529 (N_1529,In_563,In_595);
nand U1530 (N_1530,In_492,In_271);
nand U1531 (N_1531,In_428,In_589);
nor U1532 (N_1532,In_880,In_826);
nor U1533 (N_1533,In_745,In_644);
or U1534 (N_1534,In_295,In_421);
nor U1535 (N_1535,In_230,In_152);
and U1536 (N_1536,In_334,In_422);
or U1537 (N_1537,In_504,In_70);
xor U1538 (N_1538,In_381,In_706);
nand U1539 (N_1539,In_971,In_367);
nor U1540 (N_1540,In_731,In_965);
nand U1541 (N_1541,In_667,In_326);
and U1542 (N_1542,In_67,In_287);
or U1543 (N_1543,In_759,In_133);
and U1544 (N_1544,In_874,In_924);
nand U1545 (N_1545,In_690,In_962);
xnor U1546 (N_1546,In_500,In_731);
and U1547 (N_1547,In_602,In_712);
and U1548 (N_1548,In_98,In_752);
xnor U1549 (N_1549,In_23,In_534);
and U1550 (N_1550,In_680,In_413);
nor U1551 (N_1551,In_87,In_269);
nand U1552 (N_1552,In_0,In_831);
and U1553 (N_1553,In_396,In_993);
and U1554 (N_1554,In_405,In_29);
nand U1555 (N_1555,In_496,In_387);
and U1556 (N_1556,In_986,In_23);
and U1557 (N_1557,In_440,In_11);
nand U1558 (N_1558,In_561,In_14);
nor U1559 (N_1559,In_849,In_363);
and U1560 (N_1560,In_518,In_704);
and U1561 (N_1561,In_865,In_368);
nand U1562 (N_1562,In_497,In_736);
or U1563 (N_1563,In_579,In_83);
nor U1564 (N_1564,In_439,In_846);
nand U1565 (N_1565,In_74,In_852);
and U1566 (N_1566,In_338,In_528);
nand U1567 (N_1567,In_177,In_620);
nand U1568 (N_1568,In_987,In_192);
xor U1569 (N_1569,In_78,In_116);
nand U1570 (N_1570,In_911,In_273);
nand U1571 (N_1571,In_545,In_950);
nand U1572 (N_1572,In_62,In_569);
xor U1573 (N_1573,In_803,In_319);
nor U1574 (N_1574,In_881,In_128);
nor U1575 (N_1575,In_192,In_288);
xnor U1576 (N_1576,In_170,In_466);
xnor U1577 (N_1577,In_475,In_821);
or U1578 (N_1578,In_428,In_394);
or U1579 (N_1579,In_852,In_428);
and U1580 (N_1580,In_46,In_142);
and U1581 (N_1581,In_158,In_838);
and U1582 (N_1582,In_289,In_451);
xor U1583 (N_1583,In_850,In_329);
nand U1584 (N_1584,In_357,In_750);
and U1585 (N_1585,In_55,In_50);
nand U1586 (N_1586,In_61,In_467);
nand U1587 (N_1587,In_141,In_736);
xnor U1588 (N_1588,In_241,In_858);
and U1589 (N_1589,In_470,In_132);
xnor U1590 (N_1590,In_520,In_721);
xnor U1591 (N_1591,In_376,In_882);
nor U1592 (N_1592,In_408,In_187);
and U1593 (N_1593,In_991,In_887);
and U1594 (N_1594,In_799,In_484);
nor U1595 (N_1595,In_583,In_794);
nor U1596 (N_1596,In_870,In_634);
nor U1597 (N_1597,In_270,In_935);
or U1598 (N_1598,In_900,In_866);
nor U1599 (N_1599,In_41,In_978);
xnor U1600 (N_1600,In_43,In_511);
nand U1601 (N_1601,In_289,In_372);
nor U1602 (N_1602,In_980,In_469);
xnor U1603 (N_1603,In_758,In_85);
xor U1604 (N_1604,In_709,In_38);
or U1605 (N_1605,In_40,In_857);
nor U1606 (N_1606,In_964,In_478);
xnor U1607 (N_1607,In_401,In_793);
nor U1608 (N_1608,In_630,In_664);
nand U1609 (N_1609,In_938,In_497);
nor U1610 (N_1610,In_515,In_853);
nor U1611 (N_1611,In_684,In_544);
and U1612 (N_1612,In_88,In_972);
and U1613 (N_1613,In_425,In_401);
nor U1614 (N_1614,In_399,In_141);
nor U1615 (N_1615,In_678,In_197);
or U1616 (N_1616,In_953,In_601);
or U1617 (N_1617,In_818,In_213);
or U1618 (N_1618,In_696,In_25);
and U1619 (N_1619,In_261,In_63);
nand U1620 (N_1620,In_319,In_251);
xnor U1621 (N_1621,In_502,In_820);
nand U1622 (N_1622,In_562,In_104);
and U1623 (N_1623,In_418,In_576);
nand U1624 (N_1624,In_829,In_962);
and U1625 (N_1625,In_785,In_845);
nor U1626 (N_1626,In_312,In_455);
xnor U1627 (N_1627,In_183,In_792);
nor U1628 (N_1628,In_860,In_939);
nand U1629 (N_1629,In_547,In_921);
nor U1630 (N_1630,In_134,In_99);
xnor U1631 (N_1631,In_694,In_763);
nand U1632 (N_1632,In_888,In_953);
nand U1633 (N_1633,In_58,In_722);
nand U1634 (N_1634,In_745,In_13);
or U1635 (N_1635,In_943,In_975);
and U1636 (N_1636,In_61,In_909);
xnor U1637 (N_1637,In_837,In_201);
xnor U1638 (N_1638,In_944,In_662);
or U1639 (N_1639,In_373,In_426);
xnor U1640 (N_1640,In_324,In_966);
or U1641 (N_1641,In_520,In_230);
xor U1642 (N_1642,In_157,In_675);
nor U1643 (N_1643,In_148,In_403);
or U1644 (N_1644,In_806,In_437);
nand U1645 (N_1645,In_403,In_329);
xnor U1646 (N_1646,In_657,In_365);
nand U1647 (N_1647,In_462,In_374);
or U1648 (N_1648,In_663,In_150);
nand U1649 (N_1649,In_450,In_432);
nor U1650 (N_1650,In_39,In_72);
xnor U1651 (N_1651,In_64,In_781);
or U1652 (N_1652,In_180,In_438);
xnor U1653 (N_1653,In_275,In_687);
nand U1654 (N_1654,In_149,In_631);
xor U1655 (N_1655,In_472,In_57);
and U1656 (N_1656,In_363,In_551);
or U1657 (N_1657,In_279,In_299);
and U1658 (N_1658,In_167,In_573);
nor U1659 (N_1659,In_407,In_593);
and U1660 (N_1660,In_517,In_346);
xor U1661 (N_1661,In_899,In_803);
nand U1662 (N_1662,In_253,In_462);
nor U1663 (N_1663,In_766,In_65);
xor U1664 (N_1664,In_910,In_749);
or U1665 (N_1665,In_190,In_856);
nand U1666 (N_1666,In_566,In_210);
and U1667 (N_1667,In_782,In_510);
or U1668 (N_1668,In_489,In_868);
xor U1669 (N_1669,In_295,In_500);
or U1670 (N_1670,In_177,In_448);
nand U1671 (N_1671,In_403,In_203);
nor U1672 (N_1672,In_131,In_280);
nor U1673 (N_1673,In_199,In_593);
or U1674 (N_1674,In_239,In_108);
xor U1675 (N_1675,In_605,In_371);
or U1676 (N_1676,In_298,In_382);
nand U1677 (N_1677,In_858,In_157);
xnor U1678 (N_1678,In_733,In_430);
xor U1679 (N_1679,In_34,In_751);
or U1680 (N_1680,In_414,In_724);
nand U1681 (N_1681,In_684,In_186);
or U1682 (N_1682,In_444,In_769);
xor U1683 (N_1683,In_543,In_644);
xnor U1684 (N_1684,In_607,In_203);
or U1685 (N_1685,In_945,In_987);
nand U1686 (N_1686,In_366,In_817);
nand U1687 (N_1687,In_755,In_926);
nor U1688 (N_1688,In_799,In_457);
xor U1689 (N_1689,In_301,In_662);
and U1690 (N_1690,In_120,In_976);
and U1691 (N_1691,In_478,In_104);
nor U1692 (N_1692,In_649,In_941);
and U1693 (N_1693,In_295,In_530);
xnor U1694 (N_1694,In_862,In_417);
or U1695 (N_1695,In_732,In_991);
and U1696 (N_1696,In_95,In_540);
or U1697 (N_1697,In_769,In_11);
nor U1698 (N_1698,In_531,In_186);
nand U1699 (N_1699,In_13,In_962);
nor U1700 (N_1700,In_989,In_690);
or U1701 (N_1701,In_965,In_686);
and U1702 (N_1702,In_789,In_34);
nand U1703 (N_1703,In_945,In_710);
nand U1704 (N_1704,In_486,In_540);
xor U1705 (N_1705,In_947,In_359);
or U1706 (N_1706,In_280,In_907);
or U1707 (N_1707,In_96,In_416);
nand U1708 (N_1708,In_158,In_194);
nand U1709 (N_1709,In_793,In_144);
and U1710 (N_1710,In_413,In_526);
or U1711 (N_1711,In_121,In_163);
xor U1712 (N_1712,In_658,In_401);
xor U1713 (N_1713,In_869,In_192);
or U1714 (N_1714,In_516,In_912);
nor U1715 (N_1715,In_959,In_192);
xor U1716 (N_1716,In_25,In_710);
or U1717 (N_1717,In_763,In_107);
nor U1718 (N_1718,In_937,In_449);
and U1719 (N_1719,In_657,In_81);
or U1720 (N_1720,In_189,In_283);
or U1721 (N_1721,In_520,In_406);
xnor U1722 (N_1722,In_448,In_11);
nand U1723 (N_1723,In_360,In_731);
or U1724 (N_1724,In_108,In_944);
nand U1725 (N_1725,In_382,In_592);
nand U1726 (N_1726,In_322,In_690);
xor U1727 (N_1727,In_775,In_719);
or U1728 (N_1728,In_518,In_632);
nand U1729 (N_1729,In_708,In_187);
and U1730 (N_1730,In_305,In_883);
nor U1731 (N_1731,In_261,In_854);
or U1732 (N_1732,In_127,In_487);
or U1733 (N_1733,In_775,In_250);
nor U1734 (N_1734,In_181,In_275);
nor U1735 (N_1735,In_462,In_359);
or U1736 (N_1736,In_292,In_753);
or U1737 (N_1737,In_694,In_150);
nor U1738 (N_1738,In_380,In_957);
or U1739 (N_1739,In_124,In_654);
xnor U1740 (N_1740,In_249,In_139);
or U1741 (N_1741,In_548,In_9);
or U1742 (N_1742,In_402,In_294);
and U1743 (N_1743,In_258,In_61);
and U1744 (N_1744,In_767,In_879);
nand U1745 (N_1745,In_900,In_610);
xor U1746 (N_1746,In_406,In_159);
nor U1747 (N_1747,In_875,In_505);
or U1748 (N_1748,In_499,In_316);
xor U1749 (N_1749,In_767,In_961);
and U1750 (N_1750,In_799,In_427);
nor U1751 (N_1751,In_96,In_973);
or U1752 (N_1752,In_685,In_328);
or U1753 (N_1753,In_729,In_769);
nor U1754 (N_1754,In_297,In_374);
nor U1755 (N_1755,In_566,In_120);
or U1756 (N_1756,In_150,In_845);
xnor U1757 (N_1757,In_310,In_735);
or U1758 (N_1758,In_206,In_602);
xor U1759 (N_1759,In_522,In_57);
and U1760 (N_1760,In_362,In_572);
xor U1761 (N_1761,In_479,In_587);
or U1762 (N_1762,In_574,In_757);
nand U1763 (N_1763,In_530,In_164);
nor U1764 (N_1764,In_486,In_402);
nand U1765 (N_1765,In_671,In_897);
and U1766 (N_1766,In_52,In_721);
nor U1767 (N_1767,In_89,In_789);
nor U1768 (N_1768,In_607,In_371);
nand U1769 (N_1769,In_451,In_313);
nand U1770 (N_1770,In_152,In_700);
or U1771 (N_1771,In_4,In_238);
and U1772 (N_1772,In_542,In_641);
and U1773 (N_1773,In_620,In_661);
or U1774 (N_1774,In_360,In_592);
xor U1775 (N_1775,In_157,In_62);
nand U1776 (N_1776,In_723,In_904);
xnor U1777 (N_1777,In_752,In_254);
or U1778 (N_1778,In_191,In_362);
and U1779 (N_1779,In_131,In_221);
xor U1780 (N_1780,In_411,In_114);
nor U1781 (N_1781,In_103,In_38);
and U1782 (N_1782,In_480,In_344);
nand U1783 (N_1783,In_805,In_19);
xnor U1784 (N_1784,In_508,In_141);
nand U1785 (N_1785,In_404,In_825);
nand U1786 (N_1786,In_64,In_999);
and U1787 (N_1787,In_379,In_85);
or U1788 (N_1788,In_179,In_617);
or U1789 (N_1789,In_99,In_616);
or U1790 (N_1790,In_248,In_13);
nand U1791 (N_1791,In_233,In_875);
or U1792 (N_1792,In_534,In_130);
and U1793 (N_1793,In_511,In_272);
nand U1794 (N_1794,In_946,In_559);
or U1795 (N_1795,In_413,In_864);
nor U1796 (N_1796,In_366,In_704);
and U1797 (N_1797,In_351,In_995);
xnor U1798 (N_1798,In_46,In_401);
nand U1799 (N_1799,In_122,In_341);
and U1800 (N_1800,In_710,In_892);
xor U1801 (N_1801,In_600,In_402);
and U1802 (N_1802,In_14,In_22);
nand U1803 (N_1803,In_68,In_497);
xor U1804 (N_1804,In_784,In_254);
or U1805 (N_1805,In_204,In_215);
and U1806 (N_1806,In_68,In_580);
nor U1807 (N_1807,In_918,In_228);
nor U1808 (N_1808,In_21,In_99);
or U1809 (N_1809,In_445,In_185);
and U1810 (N_1810,In_197,In_615);
and U1811 (N_1811,In_71,In_755);
nor U1812 (N_1812,In_745,In_960);
nor U1813 (N_1813,In_178,In_641);
nor U1814 (N_1814,In_664,In_302);
or U1815 (N_1815,In_657,In_658);
nor U1816 (N_1816,In_259,In_117);
or U1817 (N_1817,In_631,In_300);
and U1818 (N_1818,In_387,In_414);
or U1819 (N_1819,In_281,In_720);
nand U1820 (N_1820,In_496,In_139);
or U1821 (N_1821,In_523,In_575);
and U1822 (N_1822,In_447,In_374);
nand U1823 (N_1823,In_389,In_953);
nand U1824 (N_1824,In_517,In_767);
nor U1825 (N_1825,In_978,In_569);
and U1826 (N_1826,In_192,In_62);
xor U1827 (N_1827,In_249,In_987);
and U1828 (N_1828,In_18,In_113);
or U1829 (N_1829,In_87,In_204);
and U1830 (N_1830,In_301,In_912);
nor U1831 (N_1831,In_514,In_874);
and U1832 (N_1832,In_719,In_958);
nand U1833 (N_1833,In_721,In_327);
and U1834 (N_1834,In_614,In_587);
or U1835 (N_1835,In_564,In_426);
or U1836 (N_1836,In_520,In_748);
or U1837 (N_1837,In_274,In_243);
xnor U1838 (N_1838,In_763,In_768);
xnor U1839 (N_1839,In_39,In_654);
or U1840 (N_1840,In_422,In_772);
or U1841 (N_1841,In_107,In_320);
nor U1842 (N_1842,In_751,In_511);
or U1843 (N_1843,In_29,In_559);
nand U1844 (N_1844,In_847,In_908);
and U1845 (N_1845,In_701,In_29);
or U1846 (N_1846,In_598,In_383);
xnor U1847 (N_1847,In_690,In_61);
or U1848 (N_1848,In_384,In_81);
and U1849 (N_1849,In_837,In_663);
xor U1850 (N_1850,In_747,In_501);
xor U1851 (N_1851,In_813,In_46);
or U1852 (N_1852,In_503,In_479);
nor U1853 (N_1853,In_567,In_898);
nor U1854 (N_1854,In_333,In_804);
or U1855 (N_1855,In_848,In_319);
nand U1856 (N_1856,In_199,In_238);
nor U1857 (N_1857,In_746,In_145);
xnor U1858 (N_1858,In_46,In_134);
or U1859 (N_1859,In_297,In_701);
nor U1860 (N_1860,In_951,In_669);
or U1861 (N_1861,In_742,In_92);
nand U1862 (N_1862,In_451,In_237);
nand U1863 (N_1863,In_685,In_594);
nor U1864 (N_1864,In_917,In_163);
xnor U1865 (N_1865,In_121,In_299);
or U1866 (N_1866,In_571,In_56);
and U1867 (N_1867,In_201,In_579);
and U1868 (N_1868,In_454,In_804);
and U1869 (N_1869,In_457,In_397);
or U1870 (N_1870,In_896,In_101);
or U1871 (N_1871,In_215,In_123);
xor U1872 (N_1872,In_251,In_597);
nand U1873 (N_1873,In_389,In_666);
nor U1874 (N_1874,In_311,In_27);
and U1875 (N_1875,In_987,In_399);
xnor U1876 (N_1876,In_981,In_216);
nand U1877 (N_1877,In_527,In_78);
and U1878 (N_1878,In_969,In_907);
or U1879 (N_1879,In_960,In_156);
xnor U1880 (N_1880,In_800,In_311);
or U1881 (N_1881,In_332,In_368);
nand U1882 (N_1882,In_816,In_972);
xor U1883 (N_1883,In_340,In_628);
or U1884 (N_1884,In_766,In_468);
nor U1885 (N_1885,In_857,In_62);
xnor U1886 (N_1886,In_378,In_617);
xnor U1887 (N_1887,In_609,In_59);
or U1888 (N_1888,In_496,In_405);
nand U1889 (N_1889,In_835,In_209);
or U1890 (N_1890,In_991,In_111);
or U1891 (N_1891,In_4,In_489);
nor U1892 (N_1892,In_731,In_124);
and U1893 (N_1893,In_459,In_468);
xor U1894 (N_1894,In_555,In_645);
nor U1895 (N_1895,In_215,In_461);
xnor U1896 (N_1896,In_870,In_62);
and U1897 (N_1897,In_228,In_896);
and U1898 (N_1898,In_558,In_337);
xnor U1899 (N_1899,In_899,In_453);
nand U1900 (N_1900,In_866,In_496);
nand U1901 (N_1901,In_266,In_985);
nor U1902 (N_1902,In_988,In_907);
or U1903 (N_1903,In_367,In_963);
nor U1904 (N_1904,In_358,In_151);
and U1905 (N_1905,In_124,In_455);
nand U1906 (N_1906,In_763,In_23);
or U1907 (N_1907,In_651,In_864);
or U1908 (N_1908,In_995,In_816);
or U1909 (N_1909,In_17,In_741);
nor U1910 (N_1910,In_103,In_66);
and U1911 (N_1911,In_398,In_479);
and U1912 (N_1912,In_614,In_172);
xnor U1913 (N_1913,In_623,In_541);
nor U1914 (N_1914,In_483,In_617);
xor U1915 (N_1915,In_878,In_474);
or U1916 (N_1916,In_808,In_131);
nand U1917 (N_1917,In_220,In_965);
or U1918 (N_1918,In_100,In_542);
nor U1919 (N_1919,In_501,In_841);
and U1920 (N_1920,In_194,In_826);
or U1921 (N_1921,In_765,In_705);
and U1922 (N_1922,In_976,In_482);
xor U1923 (N_1923,In_658,In_535);
and U1924 (N_1924,In_214,In_987);
xor U1925 (N_1925,In_556,In_926);
nor U1926 (N_1926,In_257,In_533);
or U1927 (N_1927,In_666,In_72);
and U1928 (N_1928,In_573,In_703);
or U1929 (N_1929,In_101,In_523);
and U1930 (N_1930,In_903,In_420);
nor U1931 (N_1931,In_466,In_525);
xor U1932 (N_1932,In_536,In_874);
and U1933 (N_1933,In_222,In_496);
xor U1934 (N_1934,In_923,In_448);
nand U1935 (N_1935,In_526,In_720);
and U1936 (N_1936,In_361,In_644);
nor U1937 (N_1937,In_684,In_283);
and U1938 (N_1938,In_779,In_783);
and U1939 (N_1939,In_477,In_655);
and U1940 (N_1940,In_852,In_64);
nand U1941 (N_1941,In_978,In_675);
xor U1942 (N_1942,In_551,In_188);
nand U1943 (N_1943,In_678,In_138);
xnor U1944 (N_1944,In_8,In_65);
and U1945 (N_1945,In_740,In_353);
or U1946 (N_1946,In_292,In_730);
nor U1947 (N_1947,In_9,In_484);
xnor U1948 (N_1948,In_564,In_279);
or U1949 (N_1949,In_437,In_601);
nor U1950 (N_1950,In_323,In_922);
xnor U1951 (N_1951,In_545,In_486);
nand U1952 (N_1952,In_512,In_340);
and U1953 (N_1953,In_607,In_768);
nand U1954 (N_1954,In_108,In_220);
or U1955 (N_1955,In_76,In_36);
nand U1956 (N_1956,In_920,In_891);
nor U1957 (N_1957,In_985,In_930);
and U1958 (N_1958,In_544,In_493);
nor U1959 (N_1959,In_926,In_353);
nor U1960 (N_1960,In_320,In_24);
nor U1961 (N_1961,In_416,In_993);
xor U1962 (N_1962,In_586,In_796);
and U1963 (N_1963,In_781,In_628);
nand U1964 (N_1964,In_237,In_38);
xnor U1965 (N_1965,In_561,In_215);
nor U1966 (N_1966,In_777,In_522);
xnor U1967 (N_1967,In_300,In_843);
and U1968 (N_1968,In_168,In_521);
or U1969 (N_1969,In_485,In_994);
and U1970 (N_1970,In_497,In_560);
and U1971 (N_1971,In_655,In_718);
and U1972 (N_1972,In_938,In_40);
nand U1973 (N_1973,In_819,In_355);
nor U1974 (N_1974,In_997,In_116);
and U1975 (N_1975,In_684,In_614);
or U1976 (N_1976,In_64,In_914);
nor U1977 (N_1977,In_289,In_169);
nand U1978 (N_1978,In_917,In_716);
xnor U1979 (N_1979,In_124,In_843);
or U1980 (N_1980,In_493,In_428);
and U1981 (N_1981,In_648,In_207);
nor U1982 (N_1982,In_900,In_48);
or U1983 (N_1983,In_663,In_170);
and U1984 (N_1984,In_460,In_408);
or U1985 (N_1985,In_362,In_464);
nor U1986 (N_1986,In_711,In_209);
or U1987 (N_1987,In_944,In_924);
or U1988 (N_1988,In_730,In_230);
nand U1989 (N_1989,In_762,In_809);
and U1990 (N_1990,In_345,In_5);
nand U1991 (N_1991,In_906,In_400);
or U1992 (N_1992,In_510,In_843);
nor U1993 (N_1993,In_2,In_102);
or U1994 (N_1994,In_937,In_987);
or U1995 (N_1995,In_46,In_405);
and U1996 (N_1996,In_44,In_613);
nor U1997 (N_1997,In_970,In_903);
nor U1998 (N_1998,In_354,In_665);
and U1999 (N_1999,In_34,In_723);
and U2000 (N_2000,N_815,N_1550);
and U2001 (N_2001,N_922,N_1015);
or U2002 (N_2002,N_309,N_851);
nand U2003 (N_2003,N_935,N_1393);
xnor U2004 (N_2004,N_373,N_984);
xor U2005 (N_2005,N_813,N_1904);
nor U2006 (N_2006,N_872,N_1941);
nor U2007 (N_2007,N_1145,N_1533);
nand U2008 (N_2008,N_55,N_80);
nand U2009 (N_2009,N_1237,N_1355);
and U2010 (N_2010,N_212,N_431);
xor U2011 (N_2011,N_395,N_434);
or U2012 (N_2012,N_1195,N_23);
nor U2013 (N_2013,N_299,N_1526);
and U2014 (N_2014,N_121,N_1947);
nor U2015 (N_2015,N_168,N_1257);
or U2016 (N_2016,N_1586,N_1814);
or U2017 (N_2017,N_1809,N_961);
and U2018 (N_2018,N_707,N_356);
nor U2019 (N_2019,N_448,N_256);
nor U2020 (N_2020,N_642,N_1148);
nor U2021 (N_2021,N_369,N_891);
or U2022 (N_2022,N_1827,N_1133);
nand U2023 (N_2023,N_1522,N_492);
and U2024 (N_2024,N_731,N_52);
nor U2025 (N_2025,N_746,N_1160);
and U2026 (N_2026,N_788,N_177);
or U2027 (N_2027,N_1937,N_1092);
or U2028 (N_2028,N_1549,N_567);
nor U2029 (N_2029,N_1365,N_986);
nor U2030 (N_2030,N_1495,N_1175);
xnor U2031 (N_2031,N_215,N_463);
nor U2032 (N_2032,N_730,N_580);
or U2033 (N_2033,N_1073,N_592);
or U2034 (N_2034,N_1482,N_1464);
nor U2035 (N_2035,N_814,N_1130);
xnor U2036 (N_2036,N_1514,N_229);
xor U2037 (N_2037,N_693,N_482);
nor U2038 (N_2038,N_1595,N_971);
and U2039 (N_2039,N_1036,N_577);
or U2040 (N_2040,N_1174,N_105);
or U2041 (N_2041,N_651,N_724);
or U2042 (N_2042,N_1633,N_1587);
or U2043 (N_2043,N_669,N_1493);
and U2044 (N_2044,N_462,N_363);
or U2045 (N_2045,N_194,N_690);
nand U2046 (N_2046,N_1953,N_1731);
or U2047 (N_2047,N_1998,N_766);
and U2048 (N_2048,N_32,N_1326);
and U2049 (N_2049,N_1745,N_141);
nand U2050 (N_2050,N_655,N_1610);
xor U2051 (N_2051,N_728,N_1795);
nand U2052 (N_2052,N_786,N_833);
nand U2053 (N_2053,N_1119,N_613);
nand U2054 (N_2054,N_173,N_501);
xor U2055 (N_2055,N_1507,N_1016);
xor U2056 (N_2056,N_519,N_1616);
nand U2057 (N_2057,N_745,N_1887);
nor U2058 (N_2058,N_364,N_1375);
or U2059 (N_2059,N_257,N_1774);
nor U2060 (N_2060,N_1746,N_608);
or U2061 (N_2061,N_1339,N_1995);
xor U2062 (N_2062,N_609,N_439);
nor U2063 (N_2063,N_416,N_1655);
xor U2064 (N_2064,N_1151,N_1758);
and U2065 (N_2065,N_920,N_1222);
or U2066 (N_2066,N_1648,N_516);
and U2067 (N_2067,N_797,N_252);
and U2068 (N_2068,N_500,N_1697);
or U2069 (N_2069,N_1909,N_1836);
and U2070 (N_2070,N_251,N_1511);
or U2071 (N_2071,N_1753,N_1192);
or U2072 (N_2072,N_960,N_254);
nor U2073 (N_2073,N_1368,N_1422);
nand U2074 (N_2074,N_404,N_735);
nor U2075 (N_2075,N_1254,N_945);
or U2076 (N_2076,N_502,N_204);
xnor U2077 (N_2077,N_110,N_1806);
xor U2078 (N_2078,N_1409,N_205);
nor U2079 (N_2079,N_1670,N_456);
or U2080 (N_2080,N_1308,N_1129);
or U2081 (N_2081,N_1531,N_799);
xor U2082 (N_2082,N_1283,N_1162);
nor U2083 (N_2083,N_1793,N_143);
xor U2084 (N_2084,N_249,N_1699);
nor U2085 (N_2085,N_650,N_1630);
xnor U2086 (N_2086,N_532,N_1852);
nand U2087 (N_2087,N_1235,N_894);
nand U2088 (N_2088,N_331,N_487);
xnor U2089 (N_2089,N_713,N_524);
and U2090 (N_2090,N_1134,N_1004);
or U2091 (N_2091,N_1426,N_852);
or U2092 (N_2092,N_1741,N_1617);
xnor U2093 (N_2093,N_1197,N_1223);
nand U2094 (N_2094,N_1647,N_937);
nor U2095 (N_2095,N_1124,N_1345);
and U2096 (N_2096,N_1387,N_1496);
and U2097 (N_2097,N_403,N_1733);
xor U2098 (N_2098,N_1445,N_1009);
xnor U2099 (N_2099,N_1159,N_161);
nor U2100 (N_2100,N_183,N_1028);
or U2101 (N_2101,N_1501,N_1157);
and U2102 (N_2102,N_647,N_1144);
xor U2103 (N_2103,N_278,N_847);
xnor U2104 (N_2104,N_1529,N_1948);
xnor U2105 (N_2105,N_732,N_96);
nor U2106 (N_2106,N_1007,N_76);
nand U2107 (N_2107,N_758,N_347);
nor U2108 (N_2108,N_1994,N_1861);
and U2109 (N_2109,N_147,N_686);
and U2110 (N_2110,N_1959,N_791);
and U2111 (N_2111,N_1650,N_754);
or U2112 (N_2112,N_1581,N_550);
and U2113 (N_2113,N_515,N_972);
nor U2114 (N_2114,N_311,N_526);
nand U2115 (N_2115,N_1076,N_1320);
nand U2116 (N_2116,N_170,N_1220);
nor U2117 (N_2117,N_1938,N_339);
and U2118 (N_2118,N_545,N_372);
nand U2119 (N_2119,N_1245,N_1026);
nor U2120 (N_2120,N_536,N_598);
and U2121 (N_2121,N_901,N_185);
xor U2122 (N_2122,N_1463,N_209);
xor U2123 (N_2123,N_1819,N_1556);
nor U2124 (N_2124,N_602,N_523);
or U2125 (N_2125,N_546,N_645);
or U2126 (N_2126,N_997,N_1239);
xnor U2127 (N_2127,N_688,N_1182);
and U2128 (N_2128,N_910,N_468);
xor U2129 (N_2129,N_1961,N_1775);
xor U2130 (N_2130,N_135,N_368);
and U2131 (N_2131,N_1373,N_822);
and U2132 (N_2132,N_1504,N_981);
or U2133 (N_2133,N_140,N_1849);
nor U2134 (N_2134,N_530,N_1503);
xor U2135 (N_2135,N_1548,N_376);
or U2136 (N_2136,N_300,N_1611);
nand U2137 (N_2137,N_874,N_101);
nor U2138 (N_2138,N_1958,N_909);
and U2139 (N_2139,N_783,N_151);
nand U2140 (N_2140,N_190,N_321);
and U2141 (N_2141,N_1155,N_1113);
nand U2142 (N_2142,N_330,N_1848);
nor U2143 (N_2143,N_585,N_762);
xor U2144 (N_2144,N_1097,N_354);
xnor U2145 (N_2145,N_255,N_1810);
nor U2146 (N_2146,N_1893,N_1221);
and U2147 (N_2147,N_1046,N_112);
and U2148 (N_2148,N_1263,N_405);
xor U2149 (N_2149,N_1988,N_264);
nand U2150 (N_2150,N_558,N_294);
nand U2151 (N_2151,N_1767,N_1043);
or U2152 (N_2152,N_1030,N_438);
nand U2153 (N_2153,N_1191,N_411);
and U2154 (N_2154,N_623,N_952);
nand U2155 (N_2155,N_892,N_1108);
nor U2156 (N_2156,N_1189,N_1275);
xnor U2157 (N_2157,N_350,N_1930);
xor U2158 (N_2158,N_88,N_129);
nand U2159 (N_2159,N_186,N_1407);
and U2160 (N_2160,N_571,N_1540);
nand U2161 (N_2161,N_1804,N_1000);
nand U2162 (N_2162,N_1834,N_1984);
or U2163 (N_2163,N_1591,N_1613);
nor U2164 (N_2164,N_722,N_1544);
nor U2165 (N_2165,N_1226,N_370);
nand U2166 (N_2166,N_583,N_664);
and U2167 (N_2167,N_322,N_725);
xnor U2168 (N_2168,N_1681,N_914);
or U2169 (N_2169,N_683,N_305);
or U2170 (N_2170,N_646,N_634);
or U2171 (N_2171,N_1816,N_1011);
xor U2172 (N_2172,N_86,N_301);
xnor U2173 (N_2173,N_378,N_1094);
nand U2174 (N_2174,N_635,N_1341);
or U2175 (N_2175,N_342,N_1494);
xnor U2176 (N_2176,N_1208,N_1140);
xor U2177 (N_2177,N_1999,N_420);
nor U2178 (N_2178,N_1954,N_421);
nand U2179 (N_2179,N_594,N_1249);
or U2180 (N_2180,N_1762,N_235);
xnor U2181 (N_2181,N_648,N_139);
and U2182 (N_2182,N_887,N_1851);
and U2183 (N_2183,N_1408,N_628);
and U2184 (N_2184,N_1858,N_1715);
nand U2185 (N_2185,N_1776,N_599);
xnor U2186 (N_2186,N_181,N_1412);
xor U2187 (N_2187,N_1770,N_108);
and U2188 (N_2188,N_1059,N_216);
nand U2189 (N_2189,N_802,N_197);
nor U2190 (N_2190,N_1943,N_668);
or U2191 (N_2191,N_1637,N_845);
or U2192 (N_2192,N_1618,N_1825);
or U2193 (N_2193,N_1467,N_1693);
xor U2194 (N_2194,N_213,N_319);
or U2195 (N_2195,N_1318,N_834);
or U2196 (N_2196,N_315,N_1038);
or U2197 (N_2197,N_980,N_965);
and U2198 (N_2198,N_1530,N_261);
and U2199 (N_2199,N_663,N_162);
xor U2200 (N_2200,N_1362,N_1604);
and U2201 (N_2201,N_1465,N_352);
or U2202 (N_2202,N_1180,N_1356);
and U2203 (N_2203,N_308,N_678);
and U2204 (N_2204,N_63,N_593);
nor U2205 (N_2205,N_1997,N_1792);
nor U2206 (N_2206,N_942,N_46);
xnor U2207 (N_2207,N_780,N_1844);
or U2208 (N_2208,N_239,N_1781);
nor U2209 (N_2209,N_221,N_1319);
xnor U2210 (N_2210,N_1480,N_1115);
nor U2211 (N_2211,N_617,N_596);
xor U2212 (N_2212,N_581,N_611);
xor U2213 (N_2213,N_640,N_1612);
and U2214 (N_2214,N_698,N_964);
and U2215 (N_2215,N_1957,N_1456);
or U2216 (N_2216,N_1980,N_206);
nor U2217 (N_2217,N_572,N_1190);
nor U2218 (N_2218,N_1098,N_24);
or U2219 (N_2219,N_1603,N_1337);
and U2220 (N_2220,N_1993,N_1940);
nand U2221 (N_2221,N_1601,N_934);
and U2222 (N_2222,N_1569,N_184);
nand U2223 (N_2223,N_464,N_486);
or U2224 (N_2224,N_760,N_214);
nor U2225 (N_2225,N_1677,N_207);
or U2226 (N_2226,N_1925,N_20);
and U2227 (N_2227,N_1967,N_1923);
nor U2228 (N_2228,N_772,N_1256);
nor U2229 (N_2229,N_1786,N_131);
xnor U2230 (N_2230,N_1079,N_414);
and U2231 (N_2231,N_1489,N_970);
nor U2232 (N_2232,N_1935,N_259);
or U2233 (N_2233,N_1734,N_440);
or U2234 (N_2234,N_993,N_1684);
and U2235 (N_2235,N_1979,N_1454);
nand U2236 (N_2236,N_916,N_1484);
nor U2237 (N_2237,N_1846,N_1340);
nand U2238 (N_2238,N_11,N_1118);
or U2239 (N_2239,N_358,N_1588);
nor U2240 (N_2240,N_1748,N_1837);
nor U2241 (N_2241,N_1910,N_533);
or U2242 (N_2242,N_954,N_904);
or U2243 (N_2243,N_1668,N_361);
nand U2244 (N_2244,N_0,N_1262);
xor U2245 (N_2245,N_1759,N_1646);
nand U2246 (N_2246,N_1952,N_918);
nor U2247 (N_2247,N_1641,N_280);
and U2248 (N_2248,N_1334,N_461);
nor U2249 (N_2249,N_233,N_554);
xnor U2250 (N_2250,N_1607,N_1832);
and U2251 (N_2251,N_898,N_351);
or U2252 (N_2252,N_600,N_862);
nor U2253 (N_2253,N_1936,N_1900);
nor U2254 (N_2254,N_97,N_320);
nand U2255 (N_2255,N_1181,N_696);
nand U2256 (N_2256,N_832,N_324);
nor U2257 (N_2257,N_312,N_1333);
or U2258 (N_2258,N_557,N_908);
nor U2259 (N_2259,N_1578,N_41);
xor U2260 (N_2260,N_1344,N_304);
nand U2261 (N_2261,N_1778,N_427);
nor U2262 (N_2262,N_751,N_1605);
nor U2263 (N_2263,N_1512,N_1545);
nand U2264 (N_2264,N_1717,N_848);
nor U2265 (N_2265,N_1455,N_1201);
or U2266 (N_2266,N_303,N_1558);
nand U2267 (N_2267,N_1372,N_1638);
nor U2268 (N_2268,N_1777,N_19);
nand U2269 (N_2269,N_485,N_1424);
xor U2270 (N_2270,N_629,N_125);
nand U2271 (N_2271,N_787,N_283);
nor U2272 (N_2272,N_559,N_578);
and U2273 (N_2273,N_33,N_38);
nand U2274 (N_2274,N_1752,N_1877);
nand U2275 (N_2275,N_1070,N_475);
nor U2276 (N_2276,N_1669,N_1913);
nand U2277 (N_2277,N_969,N_889);
nor U2278 (N_2278,N_1662,N_727);
or U2279 (N_2279,N_1072,N_1765);
and U2280 (N_2280,N_1277,N_1782);
nand U2281 (N_2281,N_1672,N_1570);
nor U2282 (N_2282,N_17,N_1788);
or U2283 (N_2283,N_1905,N_784);
or U2284 (N_2284,N_1187,N_1213);
nand U2285 (N_2285,N_1866,N_1258);
nor U2286 (N_2286,N_1838,N_752);
or U2287 (N_2287,N_1659,N_1104);
xnor U2288 (N_2288,N_1560,N_313);
and U2289 (N_2289,N_1653,N_988);
xor U2290 (N_2290,N_286,N_389);
xnor U2291 (N_2291,N_953,N_1768);
nor U2292 (N_2292,N_477,N_743);
xor U2293 (N_2293,N_1944,N_262);
and U2294 (N_2294,N_525,N_145);
and U2295 (N_2295,N_494,N_1184);
and U2296 (N_2296,N_576,N_825);
nor U2297 (N_2297,N_708,N_807);
xor U2298 (N_2298,N_306,N_756);
or U2299 (N_2299,N_1582,N_142);
or U2300 (N_2300,N_203,N_614);
or U2301 (N_2301,N_619,N_77);
nor U2302 (N_2302,N_1423,N_98);
or U2303 (N_2303,N_1143,N_1583);
nand U2304 (N_2304,N_591,N_1307);
and U2305 (N_2305,N_946,N_137);
nor U2306 (N_2306,N_798,N_1721);
nand U2307 (N_2307,N_962,N_1101);
nor U2308 (N_2308,N_1619,N_1085);
nand U2309 (N_2309,N_15,N_705);
nand U2310 (N_2310,N_1719,N_882);
xor U2311 (N_2311,N_1709,N_36);
nor U2312 (N_2312,N_1272,N_1859);
xnor U2313 (N_2313,N_1391,N_1347);
and U2314 (N_2314,N_93,N_293);
and U2315 (N_2315,N_706,N_672);
xor U2316 (N_2316,N_408,N_134);
or U2317 (N_2317,N_560,N_1193);
or U2318 (N_2318,N_511,N_1413);
and U2319 (N_2319,N_1698,N_562);
and U2320 (N_2320,N_1666,N_1679);
nand U2321 (N_2321,N_1006,N_1614);
xnor U2322 (N_2322,N_169,N_1096);
and U2323 (N_2323,N_335,N_166);
nor U2324 (N_2324,N_907,N_779);
nor U2325 (N_2325,N_1688,N_1797);
nand U2326 (N_2326,N_146,N_1439);
or U2327 (N_2327,N_1282,N_1527);
nand U2328 (N_2328,N_747,N_610);
or U2329 (N_2329,N_1280,N_1627);
nand U2330 (N_2330,N_553,N_947);
nand U2331 (N_2331,N_1031,N_712);
and U2332 (N_2332,N_375,N_1546);
and U2333 (N_2333,N_653,N_450);
and U2334 (N_2334,N_1740,N_1176);
and U2335 (N_2335,N_1343,N_1831);
nor U2336 (N_2336,N_775,N_555);
xor U2337 (N_2337,N_1790,N_966);
and U2338 (N_2338,N_1125,N_1010);
nor U2339 (N_2339,N_1084,N_1657);
xor U2340 (N_2340,N_179,N_938);
nor U2341 (N_2341,N_79,N_89);
xor U2342 (N_2342,N_341,N_1390);
nand U2343 (N_2343,N_1346,N_451);
and U2344 (N_2344,N_710,N_1014);
nand U2345 (N_2345,N_398,N_429);
nand U2346 (N_2346,N_1402,N_1080);
and U2347 (N_2347,N_211,N_130);
and U2348 (N_2348,N_896,N_857);
or U2349 (N_2349,N_520,N_1898);
or U2350 (N_2350,N_344,N_87);
xor U2351 (N_2351,N_826,N_1968);
xnor U2352 (N_2352,N_824,N_1942);
nor U2353 (N_2353,N_679,N_157);
and U2354 (N_2354,N_1592,N_1596);
nand U2355 (N_2355,N_1105,N_460);
nand U2356 (N_2356,N_26,N_950);
xnor U2357 (N_2357,N_73,N_1142);
nor U2358 (N_2358,N_83,N_1298);
and U2359 (N_2359,N_1847,N_42);
or U2360 (N_2360,N_397,N_75);
nor U2361 (N_2361,N_1951,N_1172);
nor U2362 (N_2362,N_1285,N_178);
or U2363 (N_2363,N_1442,N_535);
xnor U2364 (N_2364,N_638,N_1845);
nand U2365 (N_2365,N_1394,N_191);
nor U2366 (N_2366,N_1219,N_879);
and U2367 (N_2367,N_71,N_821);
xor U2368 (N_2368,N_1652,N_1363);
and U2369 (N_2369,N_1695,N_1574);
or U2370 (N_2370,N_956,N_296);
xor U2371 (N_2371,N_192,N_1912);
nor U2372 (N_2372,N_1061,N_1117);
xnor U2373 (N_2373,N_1029,N_1626);
nand U2374 (N_2374,N_1723,N_1966);
and U2375 (N_2375,N_268,N_835);
nand U2376 (N_2376,N_801,N_878);
xnor U2377 (N_2377,N_1460,N_1982);
xnor U2378 (N_2378,N_329,N_337);
xor U2379 (N_2379,N_765,N_1446);
nand U2380 (N_2380,N_114,N_1764);
nand U2381 (N_2381,N_603,N_1559);
nand U2382 (N_2382,N_948,N_590);
or U2383 (N_2383,N_1317,N_1022);
and U2384 (N_2384,N_1327,N_867);
xor U2385 (N_2385,N_1542,N_940);
and U2386 (N_2386,N_926,N_377);
xnor U2387 (N_2387,N_155,N_871);
xnor U2388 (N_2388,N_54,N_85);
and U2389 (N_2389,N_1121,N_1449);
nand U2390 (N_2390,N_1732,N_1150);
and U2391 (N_2391,N_276,N_1903);
nand U2392 (N_2392,N_1801,N_1576);
nand U2393 (N_2393,N_810,N_466);
or U2394 (N_2394,N_1367,N_1458);
nor U2395 (N_2395,N_1056,N_458);
xnor U2396 (N_2396,N_677,N_153);
and U2397 (N_2397,N_345,N_1867);
or U2398 (N_2398,N_625,N_994);
xnor U2399 (N_2399,N_1138,N_837);
xnor U2400 (N_2400,N_1629,N_1236);
or U2401 (N_2401,N_1265,N_1515);
nor U2402 (N_2402,N_564,N_1137);
xnor U2403 (N_2403,N_1510,N_164);
and U2404 (N_2404,N_790,N_172);
nand U2405 (N_2405,N_445,N_1479);
and U2406 (N_2406,N_327,N_1939);
or U2407 (N_2407,N_921,N_855);
and U2408 (N_2408,N_269,N_764);
xnor U2409 (N_2409,N_1091,N_1013);
nand U2410 (N_2410,N_292,N_1579);
nor U2411 (N_2411,N_84,N_1521);
xor U2412 (N_2412,N_840,N_607);
nor U2413 (N_2413,N_467,N_829);
xor U2414 (N_2414,N_1815,N_503);
nand U2415 (N_2415,N_637,N_1154);
or U2416 (N_2416,N_1818,N_1297);
or U2417 (N_2417,N_1547,N_1054);
and U2418 (N_2418,N_1253,N_1976);
or U2419 (N_2419,N_497,N_685);
xor U2420 (N_2420,N_1163,N_1032);
xor U2421 (N_2421,N_180,N_490);
xnor U2422 (N_2422,N_1787,N_1396);
nor U2423 (N_2423,N_1131,N_1562);
or U2424 (N_2424,N_1983,N_1896);
xor U2425 (N_2425,N_1803,N_45);
nor U2426 (N_2426,N_39,N_1751);
or U2427 (N_2427,N_733,N_499);
and U2428 (N_2428,N_355,N_1293);
or U2429 (N_2429,N_6,N_428);
or U2430 (N_2430,N_778,N_1987);
and U2431 (N_2431,N_393,N_115);
and U2432 (N_2432,N_1873,N_923);
and U2433 (N_2433,N_265,N_1857);
xnor U2434 (N_2434,N_44,N_1917);
nand U2435 (N_2435,N_95,N_588);
and U2436 (N_2436,N_1399,N_1403);
or U2437 (N_2437,N_61,N_1821);
or U2438 (N_2438,N_1335,N_1499);
xnor U2439 (N_2439,N_1884,N_1735);
or U2440 (N_2440,N_449,N_1209);
or U2441 (N_2441,N_556,N_1794);
or U2442 (N_2442,N_808,N_1452);
xor U2443 (N_2443,N_1271,N_27);
xor U2444 (N_2444,N_694,N_1643);
or U2445 (N_2445,N_744,N_1490);
nor U2446 (N_2446,N_528,N_1383);
and U2447 (N_2447,N_384,N_94);
or U2448 (N_2448,N_543,N_267);
nand U2449 (N_2449,N_1382,N_1744);
and U2450 (N_2450,N_16,N_1349);
nor U2451 (N_2451,N_1784,N_888);
nand U2452 (N_2452,N_43,N_806);
and U2453 (N_2453,N_817,N_1702);
or U2454 (N_2454,N_1312,N_323);
nand U2455 (N_2455,N_446,N_1431);
xor U2456 (N_2456,N_156,N_82);
and U2457 (N_2457,N_413,N_1594);
and U2458 (N_2458,N_682,N_1664);
or U2459 (N_2459,N_1077,N_1811);
nor U2460 (N_2460,N_123,N_761);
nor U2461 (N_2461,N_903,N_452);
or U2462 (N_2462,N_1268,N_91);
nor U2463 (N_2463,N_298,N_1716);
or U2464 (N_2464,N_721,N_174);
and U2465 (N_2465,N_805,N_1754);
xor U2466 (N_2466,N_1651,N_1281);
or U2467 (N_2467,N_455,N_1164);
or U2468 (N_2468,N_28,N_1481);
and U2469 (N_2469,N_812,N_1761);
and U2470 (N_2470,N_1278,N_1992);
and U2471 (N_2471,N_1194,N_1516);
and U2472 (N_2472,N_990,N_703);
and U2473 (N_2473,N_366,N_402);
nand U2474 (N_2474,N_453,N_739);
or U2475 (N_2475,N_1828,N_1251);
xor U2476 (N_2476,N_444,N_1631);
nand U2477 (N_2477,N_816,N_1242);
nand U2478 (N_2478,N_447,N_1071);
or U2479 (N_2479,N_272,N_917);
xnor U2480 (N_2480,N_1950,N_493);
or U2481 (N_2481,N_160,N_622);
nor U2482 (N_2482,N_1380,N_804);
xor U2483 (N_2483,N_955,N_621);
or U2484 (N_2484,N_1156,N_1128);
nand U2485 (N_2485,N_1856,N_1524);
and U2486 (N_2486,N_1087,N_720);
or U2487 (N_2487,N_1667,N_1728);
xnor U2488 (N_2488,N_781,N_1060);
xor U2489 (N_2489,N_1921,N_218);
xor U2490 (N_2490,N_1429,N_512);
xnor U2491 (N_2491,N_326,N_729);
xnor U2492 (N_2492,N_1049,N_1020);
nand U2493 (N_2493,N_877,N_1276);
and U2494 (N_2494,N_1215,N_605);
xnor U2495 (N_2495,N_632,N_317);
and U2496 (N_2496,N_1720,N_542);
and U2497 (N_2497,N_106,N_187);
nand U2498 (N_2498,N_843,N_1042);
nand U2499 (N_2499,N_436,N_362);
nand U2500 (N_2500,N_1066,N_1287);
nor U2501 (N_2501,N_1963,N_1932);
nor U2502 (N_2502,N_277,N_291);
nor U2503 (N_2503,N_929,N_963);
xor U2504 (N_2504,N_1881,N_1685);
nand U2505 (N_2505,N_74,N_1990);
and U2506 (N_2506,N_457,N_674);
nor U2507 (N_2507,N_924,N_1435);
xor U2508 (N_2508,N_1024,N_1606);
and U2509 (N_2509,N_1807,N_1350);
nor U2510 (N_2510,N_521,N_1416);
nand U2511 (N_2511,N_1047,N_763);
or U2512 (N_2512,N_875,N_1185);
or U2513 (N_2513,N_367,N_1589);
nor U2514 (N_2514,N_1969,N_1323);
or U2515 (N_2515,N_1945,N_69);
nand U2516 (N_2516,N_531,N_1975);
nor U2517 (N_2517,N_1041,N_1977);
nor U2518 (N_2518,N_1267,N_1568);
nor U2519 (N_2519,N_736,N_868);
nor U2520 (N_2520,N_943,N_1019);
xor U2521 (N_2521,N_124,N_1120);
xor U2522 (N_2522,N_263,N_381);
xor U2523 (N_2523,N_1244,N_1878);
xnor U2524 (N_2524,N_1750,N_473);
and U2525 (N_2525,N_1475,N_400);
or U2526 (N_2526,N_1069,N_1301);
nand U2527 (N_2527,N_1949,N_1370);
or U2528 (N_2528,N_673,N_35);
and U2529 (N_2529,N_1502,N_1057);
nand U2530 (N_2530,N_1395,N_58);
nand U2531 (N_2531,N_508,N_510);
nand U2532 (N_2532,N_1956,N_476);
and U2533 (N_2533,N_1425,N_819);
or U2534 (N_2534,N_1227,N_1989);
xor U2535 (N_2535,N_1899,N_498);
xnor U2536 (N_2536,N_568,N_587);
xor U2537 (N_2537,N_565,N_767);
and U2538 (N_2538,N_893,N_1114);
or U2539 (N_2539,N_630,N_1141);
or U2540 (N_2540,N_1246,N_675);
nand U2541 (N_2541,N_1289,N_1434);
or U2542 (N_2542,N_1817,N_1722);
nor U2543 (N_2543,N_430,N_717);
or U2544 (N_2544,N_325,N_360);
or U2545 (N_2545,N_1188,N_979);
and U2546 (N_2546,N_1528,N_37);
or U2547 (N_2547,N_1152,N_332);
nand U2548 (N_2548,N_595,N_989);
or U2549 (N_2549,N_1321,N_195);
and U2550 (N_2550,N_1273,N_715);
nor U2551 (N_2551,N_1330,N_1712);
or U2552 (N_2552,N_47,N_870);
nor U2553 (N_2553,N_809,N_509);
and U2554 (N_2554,N_1432,N_1294);
nand U2555 (N_2555,N_936,N_925);
nor U2556 (N_2556,N_454,N_1771);
nand U2557 (N_2557,N_1525,N_1342);
nor U2558 (N_2558,N_225,N_1922);
nor U2559 (N_2559,N_232,N_253);
or U2560 (N_2560,N_1021,N_853);
nand U2561 (N_2561,N_1146,N_944);
xnor U2562 (N_2562,N_830,N_234);
xor U2563 (N_2563,N_68,N_246);
nand U2564 (N_2564,N_873,N_1371);
nand U2565 (N_2565,N_517,N_171);
or U2566 (N_2566,N_90,N_769);
and U2567 (N_2567,N_1214,N_1064);
nor U2568 (N_2568,N_1632,N_51);
nor U2569 (N_2569,N_1050,N_601);
and U2570 (N_2570,N_569,N_1218);
and U2571 (N_2571,N_1597,N_1);
nand U2572 (N_2572,N_514,N_1216);
or U2573 (N_2573,N_883,N_48);
xnor U2574 (N_2574,N_1683,N_927);
nor U2575 (N_2575,N_1749,N_12);
nand U2576 (N_2576,N_1443,N_1035);
xor U2577 (N_2577,N_803,N_982);
xnor U2578 (N_2578,N_1126,N_1931);
or U2579 (N_2579,N_1247,N_1829);
or U2580 (N_2580,N_5,N_1785);
and U2581 (N_2581,N_1971,N_1791);
xor U2582 (N_2582,N_859,N_275);
xor U2583 (N_2583,N_1170,N_1955);
nor U2584 (N_2584,N_1658,N_755);
nand U2585 (N_2585,N_711,N_227);
nand U2586 (N_2586,N_67,N_1924);
nor U2587 (N_2587,N_201,N_913);
nand U2588 (N_2588,N_863,N_1789);
and U2589 (N_2589,N_1635,N_1058);
xnor U2590 (N_2590,N_422,N_1295);
and U2591 (N_2591,N_618,N_1886);
xor U2592 (N_2592,N_1173,N_1691);
xnor U2593 (N_2593,N_597,N_1441);
nor U2594 (N_2594,N_549,N_1238);
nand U2595 (N_2595,N_1474,N_1902);
nor U2596 (N_2596,N_270,N_1168);
nand U2597 (N_2597,N_1665,N_552);
or U2598 (N_2598,N_379,N_890);
or U2599 (N_2599,N_1615,N_702);
nor U2600 (N_2600,N_1377,N_1880);
nor U2601 (N_2601,N_1075,N_1730);
or U2602 (N_2602,N_886,N_1427);
nand U2603 (N_2603,N_973,N_1398);
nor U2604 (N_2604,N_976,N_340);
nor U2605 (N_2605,N_1894,N_1973);
nand U2606 (N_2606,N_346,N_1034);
nor U2607 (N_2607,N_14,N_1306);
or U2608 (N_2608,N_1654,N_1478);
and U2609 (N_2609,N_1314,N_1483);
and U2610 (N_2610,N_1625,N_589);
and U2611 (N_2611,N_1692,N_175);
xnor U2612 (N_2612,N_995,N_884);
and U2613 (N_2613,N_1012,N_522);
nor U2614 (N_2614,N_1083,N_1366);
or U2615 (N_2615,N_406,N_1336);
and U2616 (N_2616,N_676,N_1850);
xor U2617 (N_2617,N_1266,N_1534);
nand U2618 (N_2618,N_1166,N_1561);
or U2619 (N_2619,N_1714,N_504);
and U2620 (N_2620,N_1300,N_1200);
and U2621 (N_2621,N_1211,N_1357);
xnor U2622 (N_2622,N_1139,N_1675);
or U2623 (N_2623,N_1401,N_1316);
nor U2624 (N_2624,N_176,N_1779);
and U2625 (N_2625,N_584,N_656);
xnor U2626 (N_2626,N_689,N_616);
nand U2627 (N_2627,N_1315,N_469);
and U2628 (N_2628,N_459,N_704);
and U2629 (N_2629,N_250,N_1727);
nor U2630 (N_2630,N_540,N_220);
and U2631 (N_2631,N_1565,N_8);
nand U2632 (N_2632,N_231,N_1112);
and U2633 (N_2633,N_302,N_1196);
xnor U2634 (N_2634,N_912,N_133);
or U2635 (N_2635,N_1946,N_1891);
or U2636 (N_2636,N_620,N_13);
nand U2637 (N_2637,N_1868,N_1081);
nor U2638 (N_2638,N_1225,N_1639);
xor U2639 (N_2639,N_1978,N_56);
and U2640 (N_2640,N_1167,N_1178);
or U2641 (N_2641,N_21,N_1299);
and U2642 (N_2642,N_958,N_701);
xor U2643 (N_2643,N_1555,N_737);
or U2644 (N_2644,N_1198,N_118);
xnor U2645 (N_2645,N_1261,N_714);
or U2646 (N_2646,N_1351,N_1885);
or U2647 (N_2647,N_750,N_50);
or U2648 (N_2648,N_489,N_230);
nor U2649 (N_2649,N_70,N_1202);
nand U2650 (N_2650,N_748,N_1532);
or U2651 (N_2651,N_1573,N_880);
and U2652 (N_2652,N_738,N_1906);
and U2653 (N_2653,N_1572,N_1487);
or U2654 (N_2654,N_1250,N_391);
nor U2655 (N_2655,N_1093,N_974);
nand U2656 (N_2656,N_537,N_548);
nor U2657 (N_2657,N_1352,N_465);
and U2658 (N_2658,N_1203,N_388);
and U2659 (N_2659,N_1325,N_314);
nor U2660 (N_2660,N_1313,N_2);
xor U2661 (N_2661,N_1763,N_777);
and U2662 (N_2662,N_1210,N_182);
nand U2663 (N_2663,N_1869,N_1147);
nand U2664 (N_2664,N_116,N_905);
nand U2665 (N_2665,N_759,N_1005);
xor U2666 (N_2666,N_1149,N_1418);
xor U2667 (N_2667,N_1824,N_266);
nand U2668 (N_2668,N_295,N_1102);
xor U2669 (N_2669,N_1882,N_671);
nand U2670 (N_2670,N_484,N_643);
nand U2671 (N_2671,N_1820,N_1563);
xnor U2672 (N_2672,N_1875,N_435);
and U2673 (N_2673,N_800,N_838);
and U2674 (N_2674,N_1498,N_1122);
or U2675 (N_2675,N_359,N_386);
xnor U2676 (N_2676,N_196,N_1996);
or U2677 (N_2677,N_998,N_1260);
or U2678 (N_2678,N_1437,N_794);
nand U2679 (N_2679,N_1310,N_606);
xnor U2680 (N_2680,N_1890,N_1243);
nand U2681 (N_2681,N_1742,N_307);
and U2682 (N_2682,N_1388,N_1364);
xor U2683 (N_2683,N_681,N_1008);
xor U2684 (N_2684,N_697,N_529);
nand U2685 (N_2685,N_749,N_1433);
or U2686 (N_2686,N_219,N_424);
xnor U2687 (N_2687,N_1381,N_776);
xor U2688 (N_2688,N_1468,N_915);
or U2689 (N_2689,N_1879,N_684);
xor U2690 (N_2690,N_1908,N_1447);
nor U2691 (N_2691,N_1331,N_165);
xor U2692 (N_2692,N_1466,N_1621);
and U2693 (N_2693,N_1862,N_544);
xnor U2694 (N_2694,N_338,N_495);
and U2695 (N_2695,N_1911,N_1165);
and U2696 (N_2696,N_1517,N_1798);
nor U2697 (N_2697,N_1045,N_1274);
xor U2698 (N_2698,N_1259,N_1593);
and U2699 (N_2699,N_1915,N_1703);
xnor U2700 (N_2700,N_1505,N_1835);
and U2701 (N_2701,N_692,N_999);
xnor U2702 (N_2702,N_1212,N_1205);
or U2703 (N_2703,N_959,N_1769);
nor U2704 (N_2704,N_282,N_1374);
nand U2705 (N_2705,N_1600,N_1230);
or U2706 (N_2706,N_1839,N_1676);
and U2707 (N_2707,N_238,N_279);
and U2708 (N_2708,N_1726,N_1324);
nor U2709 (N_2709,N_1415,N_1506);
nand U2710 (N_2710,N_59,N_518);
and U2711 (N_2711,N_1575,N_1384);
nand U2712 (N_2712,N_757,N_1055);
nor U2713 (N_2713,N_864,N_1737);
nand U2714 (N_2714,N_563,N_1711);
nand U2715 (N_2715,N_316,N_336);
xor U2716 (N_2716,N_1585,N_649);
or U2717 (N_2717,N_1379,N_1233);
or U2718 (N_2718,N_1500,N_773);
or U2719 (N_2719,N_472,N_1962);
nor U2720 (N_2720,N_1421,N_1116);
nand U2721 (N_2721,N_1609,N_1234);
nor U2722 (N_2722,N_854,N_245);
nor U2723 (N_2723,N_1461,N_792);
or U2724 (N_2724,N_860,N_1361);
and U2725 (N_2725,N_1017,N_1623);
xnor U2726 (N_2726,N_241,N_1311);
and U2727 (N_2727,N_1303,N_390);
or U2728 (N_2728,N_1123,N_1812);
and U2729 (N_2729,N_1037,N_1889);
nand U2730 (N_2730,N_1459,N_573);
nor U2731 (N_2731,N_771,N_654);
xnor U2732 (N_2732,N_1231,N_1883);
or U2733 (N_2733,N_774,N_1964);
and U2734 (N_2734,N_1736,N_876);
or U2735 (N_2735,N_1048,N_652);
nand U2736 (N_2736,N_1292,N_866);
or U2737 (N_2737,N_1661,N_491);
and U2738 (N_2738,N_1766,N_538);
xnor U2739 (N_2739,N_897,N_1538);
or U2740 (N_2740,N_442,N_65);
or U2741 (N_2741,N_861,N_1707);
and U2742 (N_2742,N_1100,N_968);
or U2743 (N_2743,N_1485,N_841);
and U2744 (N_2744,N_1927,N_1229);
or U2745 (N_2745,N_811,N_983);
xnor U2746 (N_2746,N_1204,N_1025);
or U2747 (N_2747,N_1566,N_1309);
nor U2748 (N_2748,N_1039,N_1823);
and U2749 (N_2749,N_1718,N_152);
and U2750 (N_2750,N_644,N_111);
nand U2751 (N_2751,N_1708,N_823);
or U2752 (N_2752,N_992,N_1062);
nand U2753 (N_2753,N_1183,N_163);
nor U2754 (N_2754,N_575,N_1929);
nor U2755 (N_2755,N_1359,N_836);
nand U2756 (N_2756,N_1796,N_831);
xor U2757 (N_2757,N_1640,N_1536);
or U2758 (N_2758,N_796,N_1584);
or U2759 (N_2759,N_1406,N_1934);
and U2760 (N_2760,N_789,N_1177);
nor U2761 (N_2761,N_1743,N_1696);
nand U2762 (N_2762,N_639,N_1981);
nor U2763 (N_2763,N_1892,N_1678);
or U2764 (N_2764,N_92,N_1420);
and U2765 (N_2765,N_885,N_1111);
and U2766 (N_2766,N_401,N_667);
and U2767 (N_2767,N_741,N_941);
nor U2768 (N_2768,N_719,N_858);
nand U2769 (N_2769,N_1539,N_1358);
or U2770 (N_2770,N_40,N_1783);
and U2771 (N_2771,N_410,N_478);
nand U2772 (N_2772,N_726,N_1473);
or U2773 (N_2773,N_734,N_1040);
nand U2774 (N_2774,N_1109,N_1296);
nand U2775 (N_2775,N_1338,N_1078);
nand U2776 (N_2776,N_818,N_399);
and U2777 (N_2777,N_856,N_1649);
nor U2778 (N_2778,N_1492,N_22);
and U2779 (N_2779,N_1674,N_247);
xnor U2780 (N_2780,N_310,N_483);
xor U2781 (N_2781,N_109,N_604);
xnor U2782 (N_2782,N_827,N_407);
and U2783 (N_2783,N_1110,N_1161);
xor U2784 (N_2784,N_1863,N_334);
nand U2785 (N_2785,N_1760,N_1199);
nand U2786 (N_2786,N_1870,N_1486);
or U2787 (N_2787,N_154,N_1304);
or U2788 (N_2788,N_1874,N_223);
or U2789 (N_2789,N_1169,N_1919);
nand U2790 (N_2790,N_1290,N_1724);
xnor U2791 (N_2791,N_991,N_513);
or U2792 (N_2792,N_1477,N_657);
nand U2793 (N_2793,N_1065,N_1067);
and U2794 (N_2794,N_412,N_470);
or U2795 (N_2795,N_18,N_1855);
and U2796 (N_2796,N_1513,N_1472);
and U2797 (N_2797,N_919,N_768);
or U2798 (N_2798,N_881,N_709);
nor U2799 (N_2799,N_1052,N_78);
or U2800 (N_2800,N_29,N_1417);
nand U2801 (N_2801,N_547,N_100);
nor U2802 (N_2802,N_931,N_1153);
or U2803 (N_2803,N_1830,N_1389);
nor U2804 (N_2804,N_236,N_66);
and U2805 (N_2805,N_1755,N_288);
xor U2806 (N_2806,N_1901,N_967);
or U2807 (N_2807,N_1888,N_158);
or U2808 (N_2808,N_1103,N_1965);
and U2809 (N_2809,N_1284,N_1800);
xor U2810 (N_2810,N_348,N_633);
and U2811 (N_2811,N_666,N_700);
or U2812 (N_2812,N_740,N_1088);
and U2813 (N_2813,N_687,N_1897);
and U2814 (N_2814,N_385,N_770);
and U2815 (N_2815,N_1003,N_850);
and U2816 (N_2816,N_1687,N_1636);
or U2817 (N_2817,N_1701,N_899);
or U2818 (N_2818,N_1491,N_1599);
and U2819 (N_2819,N_1876,N_260);
or U2820 (N_2820,N_1232,N_1332);
nand U2821 (N_2821,N_906,N_1224);
or U2822 (N_2822,N_1864,N_289);
or U2823 (N_2823,N_1264,N_189);
and U2824 (N_2824,N_1551,N_1772);
xnor U2825 (N_2825,N_723,N_285);
or U2826 (N_2826,N_1255,N_1386);
and U2827 (N_2827,N_1082,N_793);
nand U2828 (N_2828,N_1974,N_1557);
xor U2829 (N_2829,N_1378,N_911);
xor U2830 (N_2830,N_665,N_1813);
nand U2831 (N_2831,N_1354,N_895);
or U2832 (N_2832,N_1571,N_188);
nor U2833 (N_2833,N_394,N_1622);
nor U2834 (N_2834,N_662,N_271);
nand U2835 (N_2835,N_1132,N_49);
and U2836 (N_2836,N_820,N_349);
or U2837 (N_2837,N_1642,N_99);
nand U2838 (N_2838,N_1279,N_1462);
or U2839 (N_2839,N_928,N_328);
and U2840 (N_2840,N_695,N_1106);
nor U2841 (N_2841,N_1348,N_1302);
and U2842 (N_2842,N_113,N_1729);
nor U2843 (N_2843,N_1519,N_1704);
nor U2844 (N_2844,N_287,N_81);
nand U2845 (N_2845,N_842,N_273);
and U2846 (N_2846,N_1186,N_1694);
nor U2847 (N_2847,N_240,N_418);
or U2848 (N_2848,N_1002,N_1686);
and U2849 (N_2849,N_357,N_374);
nor U2850 (N_2850,N_1841,N_433);
nand U2851 (N_2851,N_1972,N_975);
nand U2852 (N_2852,N_670,N_1826);
xor U2853 (N_2853,N_1598,N_1833);
and U2854 (N_2854,N_1451,N_1710);
nor U2855 (N_2855,N_1228,N_658);
xor U2856 (N_2856,N_481,N_1051);
nor U2857 (N_2857,N_1288,N_1628);
xnor U2858 (N_2858,N_1895,N_570);
or U2859 (N_2859,N_1523,N_441);
nor U2860 (N_2860,N_1689,N_30);
or U2861 (N_2861,N_541,N_680);
nor U2862 (N_2862,N_128,N_333);
nor U2863 (N_2863,N_193,N_865);
xor U2864 (N_2864,N_1291,N_290);
nand U2865 (N_2865,N_167,N_426);
and U2866 (N_2866,N_1508,N_126);
or U2867 (N_2867,N_217,N_210);
and U2868 (N_2868,N_1706,N_561);
nand U2869 (N_2869,N_1063,N_1725);
xor U2870 (N_2870,N_1488,N_844);
xor U2871 (N_2871,N_660,N_432);
xor U2872 (N_2872,N_10,N_1660);
xnor U2873 (N_2873,N_1023,N_1469);
and U2874 (N_2874,N_1799,N_1780);
nor U2875 (N_2875,N_661,N_392);
nand U2876 (N_2876,N_415,N_4);
and U2877 (N_2877,N_949,N_1305);
or U2878 (N_2878,N_9,N_1033);
and U2879 (N_2879,N_1476,N_25);
xor U2880 (N_2880,N_1444,N_297);
or U2881 (N_2881,N_1543,N_1001);
nand U2882 (N_2882,N_902,N_471);
xnor U2883 (N_2883,N_828,N_1756);
nor U2884 (N_2884,N_1535,N_846);
nand U2885 (N_2885,N_148,N_284);
xor U2886 (N_2886,N_539,N_716);
nand U2887 (N_2887,N_7,N_1018);
nor U2888 (N_2888,N_1680,N_582);
nand U2889 (N_2889,N_1590,N_1353);
and U2890 (N_2890,N_127,N_978);
nand U2891 (N_2891,N_199,N_742);
nor U2892 (N_2892,N_987,N_1960);
or U2893 (N_2893,N_939,N_409);
and U2894 (N_2894,N_136,N_795);
xor U2895 (N_2895,N_479,N_208);
nand U2896 (N_2896,N_102,N_1644);
nand U2897 (N_2897,N_1553,N_1690);
nand U2898 (N_2898,N_957,N_1840);
nor U2899 (N_2899,N_318,N_1860);
and U2900 (N_2900,N_869,N_1552);
and U2901 (N_2901,N_1135,N_1564);
xnor U2902 (N_2902,N_566,N_104);
and U2903 (N_2903,N_1865,N_1369);
xnor U2904 (N_2904,N_353,N_380);
or U2905 (N_2905,N_753,N_1252);
nand U2906 (N_2906,N_527,N_1673);
nand U2907 (N_2907,N_699,N_1757);
or U2908 (N_2908,N_60,N_159);
or U2909 (N_2909,N_274,N_226);
xor U2910 (N_2910,N_1580,N_1385);
or U2911 (N_2911,N_1985,N_612);
nand U2912 (N_2912,N_117,N_574);
and U2913 (N_2913,N_371,N_659);
nand U2914 (N_2914,N_506,N_480);
nor U2915 (N_2915,N_1842,N_641);
and U2916 (N_2916,N_849,N_122);
nor U2917 (N_2917,N_1645,N_1918);
nor U2918 (N_2918,N_132,N_1671);
nor U2919 (N_2919,N_951,N_119);
or U2920 (N_2920,N_1554,N_1567);
nand U2921 (N_2921,N_1620,N_1537);
and U2922 (N_2922,N_1397,N_1376);
or U2923 (N_2923,N_1871,N_1329);
nand U2924 (N_2924,N_103,N_1991);
and U2925 (N_2925,N_1872,N_691);
and U2926 (N_2926,N_1328,N_1095);
or U2927 (N_2927,N_1470,N_615);
xor U2928 (N_2928,N_1854,N_248);
xnor U2929 (N_2929,N_1410,N_1248);
nor U2930 (N_2930,N_1440,N_507);
xnor U2931 (N_2931,N_200,N_243);
nand U2932 (N_2932,N_1808,N_1624);
nor U2933 (N_2933,N_281,N_1207);
xor U2934 (N_2934,N_488,N_1471);
or U2935 (N_2935,N_1802,N_1541);
and U2936 (N_2936,N_1520,N_985);
nor U2937 (N_2937,N_383,N_1970);
and U2938 (N_2938,N_107,N_144);
nor U2939 (N_2939,N_496,N_1705);
xnor U2940 (N_2940,N_120,N_636);
nand U2941 (N_2941,N_782,N_1086);
xor U2942 (N_2942,N_1107,N_202);
xor U2943 (N_2943,N_1497,N_586);
xnor U2944 (N_2944,N_1634,N_34);
xor U2945 (N_2945,N_1453,N_387);
nor U2946 (N_2946,N_718,N_1158);
nor U2947 (N_2947,N_237,N_1853);
nor U2948 (N_2948,N_417,N_1933);
nor U2949 (N_2949,N_1419,N_579);
xor U2950 (N_2950,N_1053,N_53);
nand U2951 (N_2951,N_1843,N_1907);
nor U2952 (N_2952,N_138,N_1322);
nor U2953 (N_2953,N_1928,N_1509);
or U2954 (N_2954,N_1099,N_382);
and U2955 (N_2955,N_1739,N_57);
nor U2956 (N_2956,N_365,N_996);
nand U2957 (N_2957,N_437,N_1682);
nand U2958 (N_2958,N_244,N_1286);
nor U2959 (N_2959,N_1400,N_1241);
and U2960 (N_2960,N_1240,N_551);
nand U2961 (N_2961,N_1700,N_1430);
nor U2962 (N_2962,N_1089,N_1405);
xnor U2963 (N_2963,N_1926,N_1090);
and U2964 (N_2964,N_785,N_3);
xor U2965 (N_2965,N_343,N_1206);
nor U2966 (N_2966,N_258,N_1360);
nand U2967 (N_2967,N_1436,N_1428);
nand U2968 (N_2968,N_1518,N_534);
and U2969 (N_2969,N_396,N_1136);
and U2970 (N_2970,N_222,N_1920);
nor U2971 (N_2971,N_1916,N_1450);
or U2972 (N_2972,N_1577,N_419);
nand U2973 (N_2973,N_1027,N_1414);
xnor U2974 (N_2974,N_198,N_423);
or U2975 (N_2975,N_624,N_930);
and U2976 (N_2976,N_1822,N_1404);
nor U2977 (N_2977,N_31,N_631);
nand U2978 (N_2978,N_474,N_1392);
nand U2979 (N_2979,N_1074,N_977);
nor U2980 (N_2980,N_1608,N_1914);
nor U2981 (N_2981,N_1663,N_1270);
nand U2982 (N_2982,N_900,N_1713);
nor U2983 (N_2983,N_626,N_1411);
or U2984 (N_2984,N_505,N_1457);
xor U2985 (N_2985,N_933,N_1068);
and U2986 (N_2986,N_150,N_1738);
nand U2987 (N_2987,N_839,N_1448);
and U2988 (N_2988,N_425,N_1986);
and U2989 (N_2989,N_224,N_1656);
and U2990 (N_2990,N_1171,N_1044);
nor U2991 (N_2991,N_1438,N_62);
or U2992 (N_2992,N_1747,N_1127);
nand U2993 (N_2993,N_1602,N_1773);
nand U2994 (N_2994,N_443,N_1179);
nor U2995 (N_2995,N_932,N_149);
or U2996 (N_2996,N_627,N_1269);
and U2997 (N_2997,N_1805,N_1217);
and U2998 (N_2998,N_72,N_242);
nand U2999 (N_2999,N_228,N_64);
or U3000 (N_3000,N_1191,N_557);
and U3001 (N_3001,N_538,N_620);
and U3002 (N_3002,N_1094,N_1372);
and U3003 (N_3003,N_708,N_1096);
or U3004 (N_3004,N_1583,N_717);
xnor U3005 (N_3005,N_174,N_1672);
or U3006 (N_3006,N_803,N_1640);
nand U3007 (N_3007,N_252,N_1374);
xnor U3008 (N_3008,N_1148,N_512);
nand U3009 (N_3009,N_827,N_1668);
nand U3010 (N_3010,N_95,N_1907);
nor U3011 (N_3011,N_1735,N_1631);
or U3012 (N_3012,N_1239,N_173);
nand U3013 (N_3013,N_1317,N_219);
nor U3014 (N_3014,N_1019,N_1120);
xor U3015 (N_3015,N_259,N_672);
and U3016 (N_3016,N_597,N_685);
nor U3017 (N_3017,N_939,N_1297);
and U3018 (N_3018,N_1304,N_363);
xnor U3019 (N_3019,N_1467,N_358);
nor U3020 (N_3020,N_456,N_1276);
and U3021 (N_3021,N_1823,N_500);
and U3022 (N_3022,N_1623,N_215);
nand U3023 (N_3023,N_627,N_492);
nand U3024 (N_3024,N_937,N_422);
nand U3025 (N_3025,N_1895,N_413);
or U3026 (N_3026,N_295,N_394);
nor U3027 (N_3027,N_1777,N_185);
and U3028 (N_3028,N_140,N_988);
nand U3029 (N_3029,N_1431,N_737);
and U3030 (N_3030,N_909,N_847);
nand U3031 (N_3031,N_284,N_1199);
or U3032 (N_3032,N_1688,N_522);
xnor U3033 (N_3033,N_1512,N_1810);
xor U3034 (N_3034,N_962,N_1404);
xor U3035 (N_3035,N_894,N_1446);
or U3036 (N_3036,N_1465,N_820);
nand U3037 (N_3037,N_540,N_1005);
nor U3038 (N_3038,N_1130,N_800);
or U3039 (N_3039,N_905,N_517);
and U3040 (N_3040,N_1649,N_558);
nand U3041 (N_3041,N_671,N_648);
and U3042 (N_3042,N_377,N_482);
and U3043 (N_3043,N_125,N_1507);
nand U3044 (N_3044,N_634,N_336);
nor U3045 (N_3045,N_1171,N_1061);
and U3046 (N_3046,N_47,N_1430);
nor U3047 (N_3047,N_1861,N_914);
or U3048 (N_3048,N_1798,N_1979);
or U3049 (N_3049,N_88,N_462);
xnor U3050 (N_3050,N_1664,N_582);
and U3051 (N_3051,N_1749,N_629);
or U3052 (N_3052,N_1628,N_1237);
nor U3053 (N_3053,N_1402,N_1074);
or U3054 (N_3054,N_1551,N_1888);
and U3055 (N_3055,N_1670,N_1397);
nor U3056 (N_3056,N_334,N_1420);
nor U3057 (N_3057,N_1729,N_1797);
xor U3058 (N_3058,N_1531,N_686);
and U3059 (N_3059,N_1184,N_1768);
nor U3060 (N_3060,N_1770,N_639);
nor U3061 (N_3061,N_1456,N_1451);
and U3062 (N_3062,N_253,N_1181);
nand U3063 (N_3063,N_282,N_1458);
or U3064 (N_3064,N_989,N_902);
nor U3065 (N_3065,N_1438,N_1382);
nand U3066 (N_3066,N_626,N_1271);
or U3067 (N_3067,N_1053,N_1252);
nor U3068 (N_3068,N_1884,N_100);
nand U3069 (N_3069,N_314,N_877);
and U3070 (N_3070,N_302,N_1143);
nand U3071 (N_3071,N_463,N_294);
and U3072 (N_3072,N_778,N_1760);
and U3073 (N_3073,N_710,N_393);
nor U3074 (N_3074,N_1968,N_1441);
nor U3075 (N_3075,N_605,N_1751);
nand U3076 (N_3076,N_1758,N_483);
nand U3077 (N_3077,N_1253,N_1019);
nor U3078 (N_3078,N_1207,N_817);
and U3079 (N_3079,N_427,N_678);
xnor U3080 (N_3080,N_1238,N_63);
xor U3081 (N_3081,N_456,N_1649);
or U3082 (N_3082,N_540,N_1374);
nor U3083 (N_3083,N_941,N_820);
nor U3084 (N_3084,N_937,N_338);
and U3085 (N_3085,N_866,N_1621);
or U3086 (N_3086,N_1232,N_1179);
nor U3087 (N_3087,N_169,N_1915);
or U3088 (N_3088,N_1911,N_1469);
xnor U3089 (N_3089,N_1611,N_291);
nand U3090 (N_3090,N_1532,N_1733);
and U3091 (N_3091,N_1515,N_1106);
or U3092 (N_3092,N_1118,N_885);
and U3093 (N_3093,N_1196,N_25);
nand U3094 (N_3094,N_125,N_796);
nand U3095 (N_3095,N_1884,N_406);
xor U3096 (N_3096,N_65,N_1747);
nor U3097 (N_3097,N_588,N_426);
xor U3098 (N_3098,N_1979,N_1916);
nor U3099 (N_3099,N_1266,N_800);
xor U3100 (N_3100,N_1042,N_809);
or U3101 (N_3101,N_219,N_501);
or U3102 (N_3102,N_833,N_1587);
or U3103 (N_3103,N_25,N_1223);
xnor U3104 (N_3104,N_75,N_1952);
nor U3105 (N_3105,N_1754,N_450);
or U3106 (N_3106,N_1579,N_1192);
nand U3107 (N_3107,N_113,N_943);
xnor U3108 (N_3108,N_806,N_1831);
nor U3109 (N_3109,N_1661,N_38);
or U3110 (N_3110,N_321,N_1712);
nand U3111 (N_3111,N_1977,N_1841);
xnor U3112 (N_3112,N_1118,N_591);
nor U3113 (N_3113,N_944,N_1661);
nand U3114 (N_3114,N_938,N_454);
and U3115 (N_3115,N_987,N_604);
nand U3116 (N_3116,N_856,N_1708);
nor U3117 (N_3117,N_1199,N_478);
or U3118 (N_3118,N_617,N_1674);
and U3119 (N_3119,N_1165,N_133);
nand U3120 (N_3120,N_1639,N_1788);
xnor U3121 (N_3121,N_442,N_295);
or U3122 (N_3122,N_1279,N_819);
nor U3123 (N_3123,N_1264,N_661);
nand U3124 (N_3124,N_1580,N_862);
xnor U3125 (N_3125,N_1810,N_543);
nor U3126 (N_3126,N_1647,N_1034);
xor U3127 (N_3127,N_297,N_365);
xor U3128 (N_3128,N_608,N_687);
or U3129 (N_3129,N_1597,N_403);
nand U3130 (N_3130,N_948,N_862);
xnor U3131 (N_3131,N_483,N_1661);
nand U3132 (N_3132,N_974,N_1265);
xor U3133 (N_3133,N_708,N_13);
nand U3134 (N_3134,N_994,N_803);
or U3135 (N_3135,N_1084,N_1273);
nor U3136 (N_3136,N_1873,N_1526);
nand U3137 (N_3137,N_1569,N_247);
nor U3138 (N_3138,N_250,N_873);
nand U3139 (N_3139,N_1952,N_1319);
or U3140 (N_3140,N_1162,N_1332);
or U3141 (N_3141,N_1213,N_1176);
xor U3142 (N_3142,N_1180,N_1959);
xor U3143 (N_3143,N_584,N_1323);
or U3144 (N_3144,N_1180,N_532);
nand U3145 (N_3145,N_141,N_539);
xor U3146 (N_3146,N_420,N_1867);
and U3147 (N_3147,N_1683,N_755);
nor U3148 (N_3148,N_189,N_1726);
and U3149 (N_3149,N_803,N_1106);
nand U3150 (N_3150,N_606,N_1275);
and U3151 (N_3151,N_1635,N_109);
and U3152 (N_3152,N_423,N_790);
and U3153 (N_3153,N_337,N_1518);
xor U3154 (N_3154,N_419,N_428);
xor U3155 (N_3155,N_342,N_790);
and U3156 (N_3156,N_1942,N_1697);
xor U3157 (N_3157,N_1181,N_1352);
and U3158 (N_3158,N_1210,N_338);
nor U3159 (N_3159,N_931,N_1415);
xnor U3160 (N_3160,N_152,N_91);
nand U3161 (N_3161,N_1274,N_1428);
nor U3162 (N_3162,N_873,N_1482);
xor U3163 (N_3163,N_411,N_593);
nor U3164 (N_3164,N_800,N_38);
and U3165 (N_3165,N_451,N_1875);
nor U3166 (N_3166,N_1785,N_594);
and U3167 (N_3167,N_1473,N_1828);
and U3168 (N_3168,N_1410,N_733);
nor U3169 (N_3169,N_1337,N_1926);
xnor U3170 (N_3170,N_74,N_588);
nor U3171 (N_3171,N_188,N_699);
and U3172 (N_3172,N_1344,N_1924);
nor U3173 (N_3173,N_1416,N_505);
xor U3174 (N_3174,N_628,N_699);
nand U3175 (N_3175,N_321,N_1916);
nand U3176 (N_3176,N_1602,N_61);
or U3177 (N_3177,N_1641,N_1736);
nor U3178 (N_3178,N_805,N_536);
nand U3179 (N_3179,N_111,N_898);
nand U3180 (N_3180,N_626,N_1611);
xnor U3181 (N_3181,N_699,N_798);
nand U3182 (N_3182,N_253,N_698);
and U3183 (N_3183,N_807,N_768);
xnor U3184 (N_3184,N_825,N_160);
and U3185 (N_3185,N_27,N_686);
nor U3186 (N_3186,N_171,N_1010);
nand U3187 (N_3187,N_267,N_787);
and U3188 (N_3188,N_877,N_288);
nand U3189 (N_3189,N_529,N_716);
nor U3190 (N_3190,N_994,N_863);
nor U3191 (N_3191,N_302,N_316);
nand U3192 (N_3192,N_1854,N_512);
or U3193 (N_3193,N_1417,N_560);
xor U3194 (N_3194,N_945,N_1308);
and U3195 (N_3195,N_311,N_932);
or U3196 (N_3196,N_980,N_192);
nor U3197 (N_3197,N_1986,N_1886);
xor U3198 (N_3198,N_1442,N_105);
nand U3199 (N_3199,N_347,N_703);
nor U3200 (N_3200,N_1029,N_1344);
nand U3201 (N_3201,N_1328,N_1807);
xor U3202 (N_3202,N_802,N_1561);
xnor U3203 (N_3203,N_58,N_1266);
xor U3204 (N_3204,N_734,N_948);
xor U3205 (N_3205,N_181,N_771);
nor U3206 (N_3206,N_1813,N_477);
or U3207 (N_3207,N_1317,N_1121);
nand U3208 (N_3208,N_266,N_375);
nand U3209 (N_3209,N_1463,N_630);
and U3210 (N_3210,N_1724,N_1347);
nand U3211 (N_3211,N_394,N_1667);
nor U3212 (N_3212,N_1475,N_1134);
xnor U3213 (N_3213,N_467,N_1352);
or U3214 (N_3214,N_266,N_202);
or U3215 (N_3215,N_1958,N_414);
nor U3216 (N_3216,N_1047,N_310);
or U3217 (N_3217,N_833,N_155);
and U3218 (N_3218,N_19,N_478);
xnor U3219 (N_3219,N_1968,N_901);
nor U3220 (N_3220,N_1941,N_1790);
xnor U3221 (N_3221,N_1115,N_1044);
nor U3222 (N_3222,N_1698,N_1261);
or U3223 (N_3223,N_752,N_638);
xor U3224 (N_3224,N_530,N_932);
nand U3225 (N_3225,N_387,N_1520);
and U3226 (N_3226,N_586,N_1823);
nor U3227 (N_3227,N_1023,N_532);
nand U3228 (N_3228,N_1013,N_1099);
nor U3229 (N_3229,N_1161,N_1227);
nand U3230 (N_3230,N_673,N_501);
xnor U3231 (N_3231,N_333,N_1421);
xor U3232 (N_3232,N_1386,N_623);
nor U3233 (N_3233,N_616,N_1052);
nor U3234 (N_3234,N_216,N_590);
or U3235 (N_3235,N_192,N_97);
and U3236 (N_3236,N_1288,N_888);
and U3237 (N_3237,N_260,N_1593);
or U3238 (N_3238,N_939,N_402);
nand U3239 (N_3239,N_1775,N_752);
xnor U3240 (N_3240,N_460,N_214);
and U3241 (N_3241,N_106,N_881);
and U3242 (N_3242,N_1392,N_739);
and U3243 (N_3243,N_139,N_501);
and U3244 (N_3244,N_9,N_973);
nand U3245 (N_3245,N_917,N_216);
or U3246 (N_3246,N_247,N_1158);
nand U3247 (N_3247,N_1324,N_1203);
or U3248 (N_3248,N_134,N_1698);
xnor U3249 (N_3249,N_323,N_1043);
nand U3250 (N_3250,N_1720,N_1450);
or U3251 (N_3251,N_324,N_411);
xnor U3252 (N_3252,N_1017,N_1668);
and U3253 (N_3253,N_1683,N_181);
or U3254 (N_3254,N_1934,N_1333);
and U3255 (N_3255,N_1436,N_1660);
nand U3256 (N_3256,N_149,N_300);
xor U3257 (N_3257,N_1189,N_1650);
or U3258 (N_3258,N_1689,N_196);
or U3259 (N_3259,N_1527,N_1540);
nor U3260 (N_3260,N_1926,N_1712);
nor U3261 (N_3261,N_65,N_1765);
or U3262 (N_3262,N_729,N_1683);
or U3263 (N_3263,N_517,N_511);
and U3264 (N_3264,N_374,N_1971);
and U3265 (N_3265,N_1060,N_209);
or U3266 (N_3266,N_389,N_1576);
nand U3267 (N_3267,N_1225,N_1314);
and U3268 (N_3268,N_923,N_806);
xor U3269 (N_3269,N_751,N_1292);
xnor U3270 (N_3270,N_1435,N_858);
nand U3271 (N_3271,N_93,N_1077);
xor U3272 (N_3272,N_1448,N_741);
nor U3273 (N_3273,N_464,N_287);
xor U3274 (N_3274,N_676,N_1119);
nand U3275 (N_3275,N_1779,N_1895);
nor U3276 (N_3276,N_1590,N_1605);
nor U3277 (N_3277,N_1699,N_824);
or U3278 (N_3278,N_689,N_142);
nand U3279 (N_3279,N_692,N_1743);
nand U3280 (N_3280,N_1406,N_924);
and U3281 (N_3281,N_643,N_433);
and U3282 (N_3282,N_449,N_1238);
xnor U3283 (N_3283,N_1428,N_712);
or U3284 (N_3284,N_504,N_240);
and U3285 (N_3285,N_1392,N_583);
and U3286 (N_3286,N_1716,N_1827);
nor U3287 (N_3287,N_1154,N_1918);
xnor U3288 (N_3288,N_660,N_1015);
nor U3289 (N_3289,N_355,N_808);
xnor U3290 (N_3290,N_1799,N_1715);
and U3291 (N_3291,N_28,N_831);
xor U3292 (N_3292,N_946,N_146);
nand U3293 (N_3293,N_1219,N_1183);
nor U3294 (N_3294,N_518,N_1320);
nand U3295 (N_3295,N_1298,N_1301);
and U3296 (N_3296,N_309,N_1699);
xor U3297 (N_3297,N_1722,N_1994);
nor U3298 (N_3298,N_390,N_1436);
and U3299 (N_3299,N_1946,N_730);
and U3300 (N_3300,N_1223,N_89);
xor U3301 (N_3301,N_1564,N_1415);
nor U3302 (N_3302,N_1990,N_588);
and U3303 (N_3303,N_140,N_1961);
and U3304 (N_3304,N_17,N_1935);
and U3305 (N_3305,N_1763,N_1683);
nor U3306 (N_3306,N_282,N_1094);
nor U3307 (N_3307,N_751,N_413);
and U3308 (N_3308,N_679,N_316);
or U3309 (N_3309,N_1212,N_1419);
and U3310 (N_3310,N_781,N_1319);
nor U3311 (N_3311,N_1094,N_366);
xor U3312 (N_3312,N_900,N_1466);
xnor U3313 (N_3313,N_847,N_1423);
nand U3314 (N_3314,N_617,N_1226);
nand U3315 (N_3315,N_994,N_853);
nand U3316 (N_3316,N_1443,N_147);
or U3317 (N_3317,N_1968,N_745);
or U3318 (N_3318,N_880,N_1882);
xnor U3319 (N_3319,N_1580,N_917);
xnor U3320 (N_3320,N_1508,N_194);
and U3321 (N_3321,N_815,N_1482);
nor U3322 (N_3322,N_1998,N_1371);
nand U3323 (N_3323,N_665,N_995);
and U3324 (N_3324,N_710,N_1716);
nand U3325 (N_3325,N_1880,N_1326);
and U3326 (N_3326,N_584,N_598);
and U3327 (N_3327,N_1676,N_1232);
nor U3328 (N_3328,N_478,N_256);
nand U3329 (N_3329,N_352,N_569);
nand U3330 (N_3330,N_1995,N_1750);
and U3331 (N_3331,N_1164,N_1159);
or U3332 (N_3332,N_51,N_453);
and U3333 (N_3333,N_989,N_1692);
nor U3334 (N_3334,N_122,N_1857);
xor U3335 (N_3335,N_665,N_786);
or U3336 (N_3336,N_15,N_1991);
and U3337 (N_3337,N_94,N_563);
and U3338 (N_3338,N_1537,N_1219);
and U3339 (N_3339,N_588,N_1956);
and U3340 (N_3340,N_1705,N_777);
nor U3341 (N_3341,N_1616,N_1857);
and U3342 (N_3342,N_1255,N_396);
nand U3343 (N_3343,N_1092,N_127);
and U3344 (N_3344,N_1264,N_196);
nor U3345 (N_3345,N_743,N_99);
nand U3346 (N_3346,N_1240,N_290);
nor U3347 (N_3347,N_1918,N_1696);
nand U3348 (N_3348,N_166,N_763);
or U3349 (N_3349,N_1831,N_1496);
or U3350 (N_3350,N_1980,N_1582);
nand U3351 (N_3351,N_1805,N_625);
and U3352 (N_3352,N_59,N_578);
or U3353 (N_3353,N_65,N_380);
nand U3354 (N_3354,N_1422,N_916);
and U3355 (N_3355,N_1548,N_1787);
nor U3356 (N_3356,N_692,N_1267);
nor U3357 (N_3357,N_670,N_1923);
nand U3358 (N_3358,N_1631,N_1269);
and U3359 (N_3359,N_1629,N_112);
nand U3360 (N_3360,N_523,N_893);
nor U3361 (N_3361,N_17,N_331);
xnor U3362 (N_3362,N_1113,N_1377);
and U3363 (N_3363,N_774,N_795);
or U3364 (N_3364,N_1772,N_387);
xor U3365 (N_3365,N_1086,N_1507);
or U3366 (N_3366,N_1470,N_934);
or U3367 (N_3367,N_268,N_160);
nand U3368 (N_3368,N_1716,N_1195);
or U3369 (N_3369,N_382,N_92);
or U3370 (N_3370,N_1742,N_1107);
xnor U3371 (N_3371,N_1261,N_1438);
xnor U3372 (N_3372,N_562,N_300);
and U3373 (N_3373,N_608,N_1571);
nor U3374 (N_3374,N_1911,N_620);
or U3375 (N_3375,N_1372,N_19);
and U3376 (N_3376,N_181,N_1635);
nor U3377 (N_3377,N_959,N_1925);
xnor U3378 (N_3378,N_1760,N_443);
nor U3379 (N_3379,N_1901,N_1202);
or U3380 (N_3380,N_1409,N_1254);
nor U3381 (N_3381,N_860,N_169);
or U3382 (N_3382,N_1036,N_1729);
nand U3383 (N_3383,N_850,N_331);
or U3384 (N_3384,N_162,N_456);
nor U3385 (N_3385,N_1293,N_947);
or U3386 (N_3386,N_250,N_719);
nand U3387 (N_3387,N_107,N_1795);
nor U3388 (N_3388,N_1973,N_206);
and U3389 (N_3389,N_19,N_148);
xnor U3390 (N_3390,N_1328,N_763);
or U3391 (N_3391,N_242,N_1656);
xnor U3392 (N_3392,N_1307,N_287);
xor U3393 (N_3393,N_548,N_1767);
nor U3394 (N_3394,N_1479,N_94);
or U3395 (N_3395,N_1984,N_1717);
and U3396 (N_3396,N_1834,N_968);
xor U3397 (N_3397,N_68,N_1092);
nand U3398 (N_3398,N_1391,N_1618);
nor U3399 (N_3399,N_1102,N_1645);
nand U3400 (N_3400,N_70,N_249);
and U3401 (N_3401,N_540,N_644);
xnor U3402 (N_3402,N_669,N_292);
nor U3403 (N_3403,N_1237,N_1833);
xor U3404 (N_3404,N_795,N_1689);
nor U3405 (N_3405,N_1815,N_822);
nor U3406 (N_3406,N_922,N_370);
xor U3407 (N_3407,N_1070,N_1469);
nand U3408 (N_3408,N_1393,N_101);
nand U3409 (N_3409,N_1291,N_1024);
nor U3410 (N_3410,N_1895,N_512);
nand U3411 (N_3411,N_362,N_1653);
nand U3412 (N_3412,N_1300,N_1637);
nand U3413 (N_3413,N_430,N_251);
nor U3414 (N_3414,N_890,N_1846);
and U3415 (N_3415,N_34,N_1715);
and U3416 (N_3416,N_511,N_57);
and U3417 (N_3417,N_1255,N_611);
or U3418 (N_3418,N_624,N_681);
nor U3419 (N_3419,N_712,N_904);
xor U3420 (N_3420,N_57,N_1147);
or U3421 (N_3421,N_492,N_1954);
and U3422 (N_3422,N_1234,N_1144);
nor U3423 (N_3423,N_1757,N_1773);
nor U3424 (N_3424,N_785,N_1507);
and U3425 (N_3425,N_1698,N_1342);
xor U3426 (N_3426,N_390,N_1018);
xnor U3427 (N_3427,N_1019,N_1156);
xor U3428 (N_3428,N_1467,N_763);
and U3429 (N_3429,N_1447,N_1155);
nor U3430 (N_3430,N_1406,N_1720);
nor U3431 (N_3431,N_1292,N_63);
and U3432 (N_3432,N_1218,N_1075);
nor U3433 (N_3433,N_1663,N_1656);
nor U3434 (N_3434,N_71,N_1846);
and U3435 (N_3435,N_1403,N_1555);
xor U3436 (N_3436,N_1046,N_882);
and U3437 (N_3437,N_1112,N_1002);
or U3438 (N_3438,N_1043,N_1644);
nand U3439 (N_3439,N_1035,N_744);
nor U3440 (N_3440,N_313,N_832);
xor U3441 (N_3441,N_558,N_343);
or U3442 (N_3442,N_647,N_1806);
nand U3443 (N_3443,N_251,N_1167);
and U3444 (N_3444,N_1495,N_1983);
nand U3445 (N_3445,N_668,N_30);
and U3446 (N_3446,N_660,N_940);
and U3447 (N_3447,N_364,N_488);
or U3448 (N_3448,N_1330,N_1757);
xnor U3449 (N_3449,N_149,N_1474);
or U3450 (N_3450,N_1748,N_1209);
nor U3451 (N_3451,N_1413,N_92);
and U3452 (N_3452,N_659,N_211);
nand U3453 (N_3453,N_513,N_1992);
nand U3454 (N_3454,N_810,N_499);
nor U3455 (N_3455,N_1417,N_766);
nor U3456 (N_3456,N_1574,N_1587);
nor U3457 (N_3457,N_1646,N_51);
or U3458 (N_3458,N_778,N_1230);
xor U3459 (N_3459,N_179,N_1221);
nand U3460 (N_3460,N_1621,N_715);
and U3461 (N_3461,N_471,N_839);
nand U3462 (N_3462,N_630,N_1367);
xnor U3463 (N_3463,N_1355,N_968);
nor U3464 (N_3464,N_1253,N_9);
and U3465 (N_3465,N_1782,N_439);
nor U3466 (N_3466,N_145,N_1026);
nand U3467 (N_3467,N_1858,N_1334);
and U3468 (N_3468,N_1649,N_976);
or U3469 (N_3469,N_1538,N_1106);
nand U3470 (N_3470,N_1900,N_1201);
or U3471 (N_3471,N_408,N_1850);
xor U3472 (N_3472,N_132,N_1760);
nand U3473 (N_3473,N_1113,N_1541);
nor U3474 (N_3474,N_1372,N_556);
and U3475 (N_3475,N_277,N_1353);
xnor U3476 (N_3476,N_118,N_480);
or U3477 (N_3477,N_243,N_56);
nor U3478 (N_3478,N_1153,N_1061);
or U3479 (N_3479,N_1444,N_1019);
xnor U3480 (N_3480,N_1407,N_872);
xor U3481 (N_3481,N_185,N_1826);
xor U3482 (N_3482,N_1488,N_883);
nand U3483 (N_3483,N_455,N_1119);
nor U3484 (N_3484,N_1830,N_1873);
or U3485 (N_3485,N_427,N_400);
nand U3486 (N_3486,N_502,N_849);
nor U3487 (N_3487,N_1647,N_1775);
or U3488 (N_3488,N_1572,N_681);
nand U3489 (N_3489,N_1400,N_1290);
nand U3490 (N_3490,N_1384,N_1786);
and U3491 (N_3491,N_732,N_805);
or U3492 (N_3492,N_738,N_1151);
and U3493 (N_3493,N_391,N_1003);
and U3494 (N_3494,N_375,N_1092);
nor U3495 (N_3495,N_748,N_752);
nand U3496 (N_3496,N_1135,N_346);
nand U3497 (N_3497,N_1146,N_1719);
and U3498 (N_3498,N_151,N_358);
nor U3499 (N_3499,N_1278,N_919);
nor U3500 (N_3500,N_1240,N_646);
xor U3501 (N_3501,N_2,N_1989);
or U3502 (N_3502,N_435,N_278);
xor U3503 (N_3503,N_97,N_428);
nor U3504 (N_3504,N_1439,N_511);
xnor U3505 (N_3505,N_145,N_879);
and U3506 (N_3506,N_363,N_793);
nand U3507 (N_3507,N_743,N_1144);
xor U3508 (N_3508,N_1734,N_459);
or U3509 (N_3509,N_1637,N_1002);
xor U3510 (N_3510,N_148,N_246);
or U3511 (N_3511,N_1202,N_1213);
nand U3512 (N_3512,N_1590,N_1715);
nand U3513 (N_3513,N_27,N_1577);
nand U3514 (N_3514,N_572,N_1947);
nand U3515 (N_3515,N_440,N_67);
nand U3516 (N_3516,N_451,N_799);
and U3517 (N_3517,N_691,N_836);
nor U3518 (N_3518,N_1627,N_736);
nand U3519 (N_3519,N_1790,N_1862);
xor U3520 (N_3520,N_1003,N_614);
or U3521 (N_3521,N_463,N_371);
nand U3522 (N_3522,N_281,N_1136);
xor U3523 (N_3523,N_1309,N_44);
or U3524 (N_3524,N_1367,N_1056);
or U3525 (N_3525,N_579,N_384);
nor U3526 (N_3526,N_992,N_1166);
xnor U3527 (N_3527,N_1612,N_365);
nand U3528 (N_3528,N_973,N_114);
nor U3529 (N_3529,N_1810,N_35);
nor U3530 (N_3530,N_1722,N_27);
nand U3531 (N_3531,N_606,N_89);
and U3532 (N_3532,N_632,N_800);
and U3533 (N_3533,N_1847,N_1674);
nor U3534 (N_3534,N_542,N_1277);
or U3535 (N_3535,N_105,N_681);
or U3536 (N_3536,N_1240,N_1464);
or U3537 (N_3537,N_484,N_1772);
nor U3538 (N_3538,N_781,N_1837);
xnor U3539 (N_3539,N_137,N_688);
nand U3540 (N_3540,N_780,N_1323);
and U3541 (N_3541,N_160,N_1478);
or U3542 (N_3542,N_282,N_1805);
nand U3543 (N_3543,N_1183,N_1669);
xnor U3544 (N_3544,N_1577,N_1506);
or U3545 (N_3545,N_354,N_1943);
nor U3546 (N_3546,N_1839,N_1345);
nor U3547 (N_3547,N_1751,N_776);
xnor U3548 (N_3548,N_1905,N_1225);
or U3549 (N_3549,N_1596,N_480);
xor U3550 (N_3550,N_897,N_1923);
nand U3551 (N_3551,N_911,N_1185);
nor U3552 (N_3552,N_1317,N_1329);
nor U3553 (N_3553,N_851,N_182);
or U3554 (N_3554,N_1545,N_431);
or U3555 (N_3555,N_84,N_1659);
nand U3556 (N_3556,N_1440,N_1664);
and U3557 (N_3557,N_1570,N_930);
and U3558 (N_3558,N_1043,N_1628);
nand U3559 (N_3559,N_1339,N_1329);
or U3560 (N_3560,N_471,N_1682);
xor U3561 (N_3561,N_1513,N_1086);
or U3562 (N_3562,N_939,N_1051);
and U3563 (N_3563,N_279,N_727);
nor U3564 (N_3564,N_1063,N_372);
nand U3565 (N_3565,N_1770,N_131);
nand U3566 (N_3566,N_140,N_1852);
nor U3567 (N_3567,N_673,N_1370);
nand U3568 (N_3568,N_681,N_1037);
nor U3569 (N_3569,N_1544,N_1406);
or U3570 (N_3570,N_1919,N_399);
or U3571 (N_3571,N_1776,N_1127);
and U3572 (N_3572,N_1646,N_616);
xor U3573 (N_3573,N_1789,N_1070);
nor U3574 (N_3574,N_1979,N_939);
and U3575 (N_3575,N_4,N_410);
and U3576 (N_3576,N_1559,N_649);
nor U3577 (N_3577,N_475,N_1484);
nor U3578 (N_3578,N_1345,N_778);
and U3579 (N_3579,N_135,N_234);
xor U3580 (N_3580,N_1554,N_526);
or U3581 (N_3581,N_1537,N_735);
xnor U3582 (N_3582,N_141,N_1563);
nor U3583 (N_3583,N_609,N_156);
or U3584 (N_3584,N_1398,N_870);
xnor U3585 (N_3585,N_1593,N_1438);
nor U3586 (N_3586,N_262,N_833);
xor U3587 (N_3587,N_1269,N_972);
and U3588 (N_3588,N_761,N_1570);
or U3589 (N_3589,N_191,N_631);
nor U3590 (N_3590,N_993,N_1082);
xnor U3591 (N_3591,N_1111,N_1015);
xnor U3592 (N_3592,N_130,N_1170);
or U3593 (N_3593,N_552,N_303);
and U3594 (N_3594,N_1186,N_775);
nand U3595 (N_3595,N_854,N_396);
or U3596 (N_3596,N_255,N_1753);
nor U3597 (N_3597,N_295,N_1182);
and U3598 (N_3598,N_1200,N_1733);
nand U3599 (N_3599,N_1350,N_1958);
or U3600 (N_3600,N_400,N_559);
and U3601 (N_3601,N_353,N_1322);
or U3602 (N_3602,N_21,N_1590);
nand U3603 (N_3603,N_1915,N_289);
or U3604 (N_3604,N_1074,N_116);
nand U3605 (N_3605,N_10,N_1838);
and U3606 (N_3606,N_644,N_1955);
nor U3607 (N_3607,N_583,N_1566);
or U3608 (N_3608,N_1267,N_1470);
and U3609 (N_3609,N_1856,N_92);
xor U3610 (N_3610,N_380,N_1769);
nor U3611 (N_3611,N_706,N_415);
nor U3612 (N_3612,N_1810,N_1497);
nand U3613 (N_3613,N_1548,N_474);
and U3614 (N_3614,N_295,N_1259);
xor U3615 (N_3615,N_1036,N_1937);
and U3616 (N_3616,N_1363,N_1064);
and U3617 (N_3617,N_1262,N_1385);
xnor U3618 (N_3618,N_1387,N_1964);
and U3619 (N_3619,N_1997,N_702);
or U3620 (N_3620,N_1717,N_1753);
or U3621 (N_3621,N_742,N_1795);
and U3622 (N_3622,N_679,N_1764);
nor U3623 (N_3623,N_1249,N_500);
xnor U3624 (N_3624,N_1587,N_997);
and U3625 (N_3625,N_1808,N_285);
nor U3626 (N_3626,N_459,N_445);
xnor U3627 (N_3627,N_234,N_1899);
nand U3628 (N_3628,N_1800,N_518);
and U3629 (N_3629,N_1575,N_984);
xnor U3630 (N_3630,N_1289,N_144);
nor U3631 (N_3631,N_864,N_96);
or U3632 (N_3632,N_555,N_1326);
nand U3633 (N_3633,N_1586,N_737);
and U3634 (N_3634,N_293,N_1586);
nand U3635 (N_3635,N_1889,N_384);
xor U3636 (N_3636,N_1504,N_425);
nand U3637 (N_3637,N_57,N_1557);
nor U3638 (N_3638,N_941,N_1106);
nand U3639 (N_3639,N_1412,N_539);
nand U3640 (N_3640,N_429,N_1561);
and U3641 (N_3641,N_1871,N_149);
xor U3642 (N_3642,N_830,N_258);
and U3643 (N_3643,N_20,N_1337);
nor U3644 (N_3644,N_909,N_475);
xor U3645 (N_3645,N_1486,N_191);
xnor U3646 (N_3646,N_1458,N_706);
and U3647 (N_3647,N_1526,N_205);
or U3648 (N_3648,N_855,N_1126);
or U3649 (N_3649,N_720,N_912);
or U3650 (N_3650,N_1747,N_1662);
xor U3651 (N_3651,N_1614,N_1618);
xor U3652 (N_3652,N_1698,N_1483);
and U3653 (N_3653,N_1301,N_1440);
and U3654 (N_3654,N_1803,N_1476);
nand U3655 (N_3655,N_295,N_290);
nor U3656 (N_3656,N_621,N_253);
xor U3657 (N_3657,N_355,N_1289);
nand U3658 (N_3658,N_1078,N_1691);
nand U3659 (N_3659,N_1627,N_629);
nor U3660 (N_3660,N_1531,N_51);
nand U3661 (N_3661,N_851,N_1988);
nor U3662 (N_3662,N_109,N_489);
xor U3663 (N_3663,N_390,N_890);
and U3664 (N_3664,N_1478,N_1365);
xnor U3665 (N_3665,N_671,N_39);
nand U3666 (N_3666,N_934,N_244);
xor U3667 (N_3667,N_1357,N_115);
xnor U3668 (N_3668,N_1121,N_825);
or U3669 (N_3669,N_596,N_1315);
or U3670 (N_3670,N_1206,N_1023);
nor U3671 (N_3671,N_441,N_1746);
or U3672 (N_3672,N_1609,N_951);
or U3673 (N_3673,N_1553,N_1973);
nand U3674 (N_3674,N_377,N_1719);
xnor U3675 (N_3675,N_1184,N_547);
nand U3676 (N_3676,N_1382,N_1929);
or U3677 (N_3677,N_1550,N_327);
and U3678 (N_3678,N_1751,N_574);
nand U3679 (N_3679,N_76,N_940);
or U3680 (N_3680,N_1178,N_522);
nor U3681 (N_3681,N_883,N_1682);
nand U3682 (N_3682,N_162,N_467);
xnor U3683 (N_3683,N_793,N_820);
and U3684 (N_3684,N_1412,N_1239);
and U3685 (N_3685,N_1709,N_1738);
or U3686 (N_3686,N_306,N_444);
and U3687 (N_3687,N_1187,N_1417);
nand U3688 (N_3688,N_721,N_1873);
nor U3689 (N_3689,N_407,N_1824);
nand U3690 (N_3690,N_1414,N_1713);
nor U3691 (N_3691,N_1189,N_300);
xor U3692 (N_3692,N_23,N_365);
and U3693 (N_3693,N_280,N_1547);
nand U3694 (N_3694,N_361,N_565);
nand U3695 (N_3695,N_1669,N_1180);
or U3696 (N_3696,N_1694,N_1692);
nand U3697 (N_3697,N_1067,N_422);
xnor U3698 (N_3698,N_243,N_1635);
nor U3699 (N_3699,N_228,N_1173);
nor U3700 (N_3700,N_1334,N_1250);
and U3701 (N_3701,N_356,N_111);
xor U3702 (N_3702,N_1572,N_833);
nor U3703 (N_3703,N_1855,N_488);
and U3704 (N_3704,N_1398,N_362);
nor U3705 (N_3705,N_320,N_1682);
or U3706 (N_3706,N_1491,N_1047);
and U3707 (N_3707,N_389,N_600);
nor U3708 (N_3708,N_854,N_1061);
nor U3709 (N_3709,N_585,N_1013);
and U3710 (N_3710,N_630,N_609);
nor U3711 (N_3711,N_1330,N_964);
and U3712 (N_3712,N_221,N_1002);
xor U3713 (N_3713,N_1538,N_1745);
nand U3714 (N_3714,N_454,N_1602);
nor U3715 (N_3715,N_1371,N_1308);
nand U3716 (N_3716,N_1580,N_1698);
nand U3717 (N_3717,N_648,N_305);
nand U3718 (N_3718,N_69,N_552);
nor U3719 (N_3719,N_234,N_1250);
and U3720 (N_3720,N_1789,N_1800);
nor U3721 (N_3721,N_1063,N_664);
nand U3722 (N_3722,N_714,N_438);
nand U3723 (N_3723,N_1278,N_1250);
nand U3724 (N_3724,N_1701,N_1918);
nor U3725 (N_3725,N_1883,N_426);
xor U3726 (N_3726,N_1161,N_1122);
or U3727 (N_3727,N_518,N_1143);
nand U3728 (N_3728,N_650,N_1479);
nor U3729 (N_3729,N_943,N_46);
xnor U3730 (N_3730,N_383,N_872);
or U3731 (N_3731,N_751,N_1345);
xnor U3732 (N_3732,N_1224,N_1832);
or U3733 (N_3733,N_927,N_692);
nor U3734 (N_3734,N_1235,N_119);
nor U3735 (N_3735,N_560,N_357);
nand U3736 (N_3736,N_1188,N_1533);
nand U3737 (N_3737,N_1984,N_914);
and U3738 (N_3738,N_595,N_1155);
nand U3739 (N_3739,N_193,N_1701);
nor U3740 (N_3740,N_537,N_205);
or U3741 (N_3741,N_845,N_378);
nor U3742 (N_3742,N_1472,N_333);
xor U3743 (N_3743,N_1252,N_469);
nand U3744 (N_3744,N_1868,N_1732);
nor U3745 (N_3745,N_832,N_519);
nor U3746 (N_3746,N_823,N_928);
or U3747 (N_3747,N_1385,N_1661);
and U3748 (N_3748,N_807,N_1538);
and U3749 (N_3749,N_1099,N_1846);
and U3750 (N_3750,N_680,N_892);
and U3751 (N_3751,N_1367,N_141);
nand U3752 (N_3752,N_1338,N_1403);
and U3753 (N_3753,N_1091,N_83);
or U3754 (N_3754,N_546,N_777);
or U3755 (N_3755,N_461,N_122);
nor U3756 (N_3756,N_407,N_628);
or U3757 (N_3757,N_1790,N_667);
or U3758 (N_3758,N_960,N_1206);
nand U3759 (N_3759,N_1615,N_138);
or U3760 (N_3760,N_696,N_1604);
and U3761 (N_3761,N_1643,N_364);
xnor U3762 (N_3762,N_1350,N_1663);
nand U3763 (N_3763,N_1684,N_487);
nand U3764 (N_3764,N_1684,N_739);
nor U3765 (N_3765,N_1040,N_1217);
and U3766 (N_3766,N_1975,N_1823);
or U3767 (N_3767,N_359,N_1370);
and U3768 (N_3768,N_1033,N_1568);
and U3769 (N_3769,N_858,N_1252);
nand U3770 (N_3770,N_134,N_1588);
and U3771 (N_3771,N_1015,N_509);
or U3772 (N_3772,N_886,N_979);
nor U3773 (N_3773,N_1523,N_421);
or U3774 (N_3774,N_1056,N_888);
and U3775 (N_3775,N_838,N_444);
nor U3776 (N_3776,N_1089,N_470);
or U3777 (N_3777,N_1204,N_954);
xor U3778 (N_3778,N_528,N_1323);
nor U3779 (N_3779,N_1107,N_1563);
nand U3780 (N_3780,N_1573,N_398);
nand U3781 (N_3781,N_727,N_576);
and U3782 (N_3782,N_680,N_1912);
nor U3783 (N_3783,N_763,N_832);
nand U3784 (N_3784,N_571,N_693);
and U3785 (N_3785,N_1789,N_10);
nor U3786 (N_3786,N_561,N_306);
or U3787 (N_3787,N_726,N_1275);
and U3788 (N_3788,N_1528,N_1186);
xor U3789 (N_3789,N_1823,N_944);
nor U3790 (N_3790,N_648,N_1551);
xnor U3791 (N_3791,N_1585,N_691);
or U3792 (N_3792,N_1681,N_1635);
nor U3793 (N_3793,N_177,N_1811);
nand U3794 (N_3794,N_677,N_57);
xor U3795 (N_3795,N_1870,N_713);
xor U3796 (N_3796,N_1567,N_408);
nor U3797 (N_3797,N_977,N_1220);
nand U3798 (N_3798,N_1344,N_1261);
nand U3799 (N_3799,N_354,N_157);
or U3800 (N_3800,N_133,N_79);
and U3801 (N_3801,N_455,N_73);
nand U3802 (N_3802,N_1936,N_776);
nor U3803 (N_3803,N_924,N_260);
nand U3804 (N_3804,N_1035,N_1750);
nand U3805 (N_3805,N_524,N_800);
or U3806 (N_3806,N_1748,N_827);
xor U3807 (N_3807,N_1836,N_1692);
or U3808 (N_3808,N_622,N_1190);
nand U3809 (N_3809,N_862,N_877);
or U3810 (N_3810,N_510,N_1932);
and U3811 (N_3811,N_340,N_784);
xnor U3812 (N_3812,N_147,N_10);
or U3813 (N_3813,N_881,N_1663);
xnor U3814 (N_3814,N_916,N_1743);
or U3815 (N_3815,N_178,N_1096);
nor U3816 (N_3816,N_1253,N_333);
and U3817 (N_3817,N_195,N_1017);
or U3818 (N_3818,N_548,N_1857);
xnor U3819 (N_3819,N_640,N_1095);
or U3820 (N_3820,N_1088,N_1967);
nor U3821 (N_3821,N_1468,N_1839);
nand U3822 (N_3822,N_935,N_1068);
and U3823 (N_3823,N_886,N_1826);
nand U3824 (N_3824,N_889,N_1244);
or U3825 (N_3825,N_62,N_994);
or U3826 (N_3826,N_1966,N_1804);
or U3827 (N_3827,N_1072,N_834);
or U3828 (N_3828,N_270,N_744);
and U3829 (N_3829,N_125,N_867);
and U3830 (N_3830,N_1983,N_550);
and U3831 (N_3831,N_434,N_1203);
xnor U3832 (N_3832,N_1688,N_1091);
xor U3833 (N_3833,N_1159,N_154);
nor U3834 (N_3834,N_344,N_1897);
nor U3835 (N_3835,N_1891,N_1609);
nand U3836 (N_3836,N_137,N_1448);
or U3837 (N_3837,N_1059,N_144);
and U3838 (N_3838,N_1354,N_1365);
nand U3839 (N_3839,N_1145,N_350);
or U3840 (N_3840,N_463,N_1589);
nand U3841 (N_3841,N_278,N_1535);
nor U3842 (N_3842,N_1824,N_1432);
xnor U3843 (N_3843,N_968,N_1742);
nand U3844 (N_3844,N_59,N_897);
xor U3845 (N_3845,N_1547,N_1410);
nor U3846 (N_3846,N_665,N_396);
xnor U3847 (N_3847,N_253,N_985);
or U3848 (N_3848,N_670,N_239);
or U3849 (N_3849,N_741,N_731);
or U3850 (N_3850,N_1826,N_1002);
or U3851 (N_3851,N_896,N_136);
nand U3852 (N_3852,N_1564,N_57);
nor U3853 (N_3853,N_156,N_1818);
nand U3854 (N_3854,N_1233,N_1591);
or U3855 (N_3855,N_1839,N_481);
or U3856 (N_3856,N_294,N_496);
and U3857 (N_3857,N_1543,N_960);
and U3858 (N_3858,N_412,N_1096);
and U3859 (N_3859,N_1883,N_1507);
xor U3860 (N_3860,N_248,N_116);
or U3861 (N_3861,N_94,N_1946);
nor U3862 (N_3862,N_995,N_327);
or U3863 (N_3863,N_1300,N_435);
or U3864 (N_3864,N_1663,N_1858);
or U3865 (N_3865,N_1599,N_177);
or U3866 (N_3866,N_518,N_683);
xor U3867 (N_3867,N_101,N_851);
or U3868 (N_3868,N_0,N_1465);
nand U3869 (N_3869,N_1854,N_303);
or U3870 (N_3870,N_1676,N_1752);
nor U3871 (N_3871,N_1859,N_1051);
nor U3872 (N_3872,N_1439,N_1236);
and U3873 (N_3873,N_404,N_326);
nor U3874 (N_3874,N_827,N_1103);
or U3875 (N_3875,N_31,N_1816);
or U3876 (N_3876,N_1282,N_653);
and U3877 (N_3877,N_1548,N_80);
and U3878 (N_3878,N_918,N_1229);
nand U3879 (N_3879,N_1756,N_1818);
or U3880 (N_3880,N_623,N_1260);
and U3881 (N_3881,N_1153,N_665);
or U3882 (N_3882,N_1851,N_515);
or U3883 (N_3883,N_1822,N_589);
nand U3884 (N_3884,N_1894,N_954);
xor U3885 (N_3885,N_1897,N_1461);
or U3886 (N_3886,N_26,N_1719);
and U3887 (N_3887,N_376,N_1927);
or U3888 (N_3888,N_1027,N_464);
nor U3889 (N_3889,N_1655,N_558);
or U3890 (N_3890,N_1130,N_1900);
and U3891 (N_3891,N_919,N_665);
nor U3892 (N_3892,N_1343,N_507);
nor U3893 (N_3893,N_600,N_82);
nand U3894 (N_3894,N_194,N_1922);
or U3895 (N_3895,N_730,N_671);
nand U3896 (N_3896,N_1036,N_1594);
nand U3897 (N_3897,N_289,N_878);
nor U3898 (N_3898,N_1843,N_892);
xor U3899 (N_3899,N_338,N_1260);
nand U3900 (N_3900,N_582,N_1438);
and U3901 (N_3901,N_608,N_353);
and U3902 (N_3902,N_1524,N_1906);
xor U3903 (N_3903,N_220,N_1072);
or U3904 (N_3904,N_1801,N_1182);
nand U3905 (N_3905,N_1715,N_516);
xor U3906 (N_3906,N_1461,N_670);
xnor U3907 (N_3907,N_947,N_457);
nor U3908 (N_3908,N_1447,N_34);
and U3909 (N_3909,N_1120,N_390);
nand U3910 (N_3910,N_502,N_1181);
and U3911 (N_3911,N_106,N_232);
nand U3912 (N_3912,N_674,N_1170);
and U3913 (N_3913,N_1301,N_433);
nand U3914 (N_3914,N_617,N_289);
nand U3915 (N_3915,N_618,N_1778);
nand U3916 (N_3916,N_900,N_632);
nor U3917 (N_3917,N_889,N_1349);
nand U3918 (N_3918,N_803,N_792);
nand U3919 (N_3919,N_421,N_1385);
nand U3920 (N_3920,N_264,N_464);
xnor U3921 (N_3921,N_285,N_1930);
nor U3922 (N_3922,N_1928,N_1035);
xnor U3923 (N_3923,N_985,N_1030);
nand U3924 (N_3924,N_1026,N_84);
xnor U3925 (N_3925,N_117,N_1829);
nor U3926 (N_3926,N_969,N_1089);
and U3927 (N_3927,N_1640,N_1050);
or U3928 (N_3928,N_686,N_909);
xor U3929 (N_3929,N_593,N_1601);
nor U3930 (N_3930,N_1584,N_760);
nand U3931 (N_3931,N_444,N_1330);
nand U3932 (N_3932,N_163,N_1879);
and U3933 (N_3933,N_1410,N_726);
nor U3934 (N_3934,N_1840,N_79);
nand U3935 (N_3935,N_91,N_1591);
xor U3936 (N_3936,N_76,N_56);
or U3937 (N_3937,N_1383,N_1526);
and U3938 (N_3938,N_1655,N_1033);
and U3939 (N_3939,N_796,N_1715);
or U3940 (N_3940,N_1545,N_324);
xor U3941 (N_3941,N_594,N_1074);
or U3942 (N_3942,N_1963,N_823);
or U3943 (N_3943,N_1782,N_1321);
or U3944 (N_3944,N_33,N_1757);
xor U3945 (N_3945,N_1725,N_713);
nor U3946 (N_3946,N_306,N_1060);
xnor U3947 (N_3947,N_1820,N_1020);
nand U3948 (N_3948,N_1762,N_1668);
nor U3949 (N_3949,N_470,N_361);
xor U3950 (N_3950,N_183,N_1195);
nor U3951 (N_3951,N_1475,N_1150);
xnor U3952 (N_3952,N_1029,N_14);
nand U3953 (N_3953,N_1920,N_671);
nand U3954 (N_3954,N_816,N_1636);
or U3955 (N_3955,N_380,N_1296);
nor U3956 (N_3956,N_529,N_1063);
nand U3957 (N_3957,N_1550,N_60);
nor U3958 (N_3958,N_1536,N_635);
and U3959 (N_3959,N_417,N_1407);
or U3960 (N_3960,N_206,N_1722);
nor U3961 (N_3961,N_1270,N_1237);
and U3962 (N_3962,N_17,N_434);
nor U3963 (N_3963,N_1724,N_661);
nand U3964 (N_3964,N_207,N_1296);
nand U3965 (N_3965,N_974,N_1614);
nor U3966 (N_3966,N_568,N_564);
or U3967 (N_3967,N_1559,N_986);
xor U3968 (N_3968,N_981,N_1284);
xnor U3969 (N_3969,N_1545,N_452);
or U3970 (N_3970,N_1158,N_962);
and U3971 (N_3971,N_1080,N_1266);
and U3972 (N_3972,N_618,N_512);
nor U3973 (N_3973,N_843,N_417);
and U3974 (N_3974,N_67,N_423);
and U3975 (N_3975,N_1801,N_1039);
xor U3976 (N_3976,N_1201,N_1970);
or U3977 (N_3977,N_959,N_1324);
and U3978 (N_3978,N_720,N_966);
nor U3979 (N_3979,N_38,N_763);
nand U3980 (N_3980,N_508,N_231);
and U3981 (N_3981,N_26,N_546);
nor U3982 (N_3982,N_1151,N_1277);
nor U3983 (N_3983,N_1907,N_1430);
nor U3984 (N_3984,N_810,N_950);
nor U3985 (N_3985,N_28,N_847);
nor U3986 (N_3986,N_852,N_1025);
nand U3987 (N_3987,N_640,N_354);
and U3988 (N_3988,N_901,N_167);
nor U3989 (N_3989,N_460,N_1128);
nand U3990 (N_3990,N_1187,N_196);
nor U3991 (N_3991,N_1141,N_1942);
or U3992 (N_3992,N_141,N_171);
or U3993 (N_3993,N_193,N_280);
xnor U3994 (N_3994,N_673,N_1130);
and U3995 (N_3995,N_1604,N_1374);
or U3996 (N_3996,N_1426,N_1745);
nor U3997 (N_3997,N_269,N_895);
nor U3998 (N_3998,N_447,N_324);
nor U3999 (N_3999,N_524,N_40);
and U4000 (N_4000,N_2798,N_2110);
and U4001 (N_4001,N_2840,N_3483);
nor U4002 (N_4002,N_3796,N_3987);
nand U4003 (N_4003,N_2395,N_2909);
xor U4004 (N_4004,N_3390,N_2932);
and U4005 (N_4005,N_3913,N_2913);
or U4006 (N_4006,N_2308,N_3960);
or U4007 (N_4007,N_3232,N_3793);
xor U4008 (N_4008,N_3735,N_3239);
nand U4009 (N_4009,N_2153,N_3554);
nand U4010 (N_4010,N_2648,N_3800);
nor U4011 (N_4011,N_2875,N_2499);
nor U4012 (N_4012,N_2267,N_2322);
nand U4013 (N_4013,N_2792,N_3714);
nand U4014 (N_4014,N_3967,N_2761);
or U4015 (N_4015,N_3475,N_3188);
and U4016 (N_4016,N_2524,N_2218);
and U4017 (N_4017,N_3296,N_3459);
nor U4018 (N_4018,N_2513,N_2626);
nand U4019 (N_4019,N_3241,N_2955);
nor U4020 (N_4020,N_2755,N_2887);
nor U4021 (N_4021,N_3910,N_2802);
nor U4022 (N_4022,N_3309,N_3036);
or U4023 (N_4023,N_2098,N_2115);
xnor U4024 (N_4024,N_3864,N_3210);
nand U4025 (N_4025,N_2476,N_2057);
or U4026 (N_4026,N_3692,N_2271);
xnor U4027 (N_4027,N_3731,N_3620);
and U4028 (N_4028,N_3738,N_2597);
and U4029 (N_4029,N_3784,N_3123);
and U4030 (N_4030,N_3672,N_3280);
and U4031 (N_4031,N_2140,N_2179);
nand U4032 (N_4032,N_2008,N_2893);
and U4033 (N_4033,N_2343,N_2034);
or U4034 (N_4034,N_2454,N_3785);
nor U4035 (N_4035,N_3596,N_3129);
nor U4036 (N_4036,N_2885,N_3988);
and U4037 (N_4037,N_3400,N_3387);
xor U4038 (N_4038,N_2611,N_3011);
nor U4039 (N_4039,N_2128,N_2192);
or U4040 (N_4040,N_2331,N_2073);
nor U4041 (N_4041,N_3328,N_2938);
xor U4042 (N_4042,N_2497,N_2441);
xor U4043 (N_4043,N_2920,N_2613);
nor U4044 (N_4044,N_2171,N_2534);
nand U4045 (N_4045,N_2634,N_3093);
xor U4046 (N_4046,N_3555,N_2667);
or U4047 (N_4047,N_2195,N_3087);
nor U4048 (N_4048,N_2064,N_3171);
xnor U4049 (N_4049,N_2815,N_3574);
and U4050 (N_4050,N_2656,N_3410);
nor U4051 (N_4051,N_2849,N_2004);
xor U4052 (N_4052,N_3030,N_2374);
nand U4053 (N_4053,N_2445,N_2075);
and U4054 (N_4054,N_3031,N_3366);
nand U4055 (N_4055,N_3331,N_2202);
nor U4056 (N_4056,N_3004,N_2463);
or U4057 (N_4057,N_2207,N_3329);
nor U4058 (N_4058,N_3112,N_2067);
xnor U4059 (N_4059,N_2472,N_2341);
nand U4060 (N_4060,N_3308,N_3393);
xor U4061 (N_4061,N_3628,N_2651);
nor U4062 (N_4062,N_2683,N_2049);
and U4063 (N_4063,N_3652,N_3952);
and U4064 (N_4064,N_3565,N_2041);
and U4065 (N_4065,N_3334,N_3127);
and U4066 (N_4066,N_3920,N_3580);
and U4067 (N_4067,N_2339,N_3655);
or U4068 (N_4068,N_2520,N_3552);
nor U4069 (N_4069,N_3000,N_3852);
nor U4070 (N_4070,N_2869,N_3613);
xnor U4071 (N_4071,N_3290,N_3423);
nor U4072 (N_4072,N_3931,N_2045);
or U4073 (N_4073,N_3950,N_2829);
or U4074 (N_4074,N_3181,N_3252);
nor U4075 (N_4075,N_3942,N_3279);
and U4076 (N_4076,N_3616,N_2591);
nand U4077 (N_4077,N_3072,N_3917);
xnor U4078 (N_4078,N_2797,N_3198);
or U4079 (N_4079,N_2163,N_2675);
xnor U4080 (N_4080,N_3395,N_3775);
nand U4081 (N_4081,N_3377,N_2738);
or U4082 (N_4082,N_2927,N_3227);
xnor U4083 (N_4083,N_3892,N_2154);
and U4084 (N_4084,N_3243,N_2354);
xnor U4085 (N_4085,N_3458,N_3570);
or U4086 (N_4086,N_2779,N_3592);
and U4087 (N_4087,N_3027,N_3343);
xor U4088 (N_4088,N_3765,N_3991);
nand U4089 (N_4089,N_3949,N_2165);
nand U4090 (N_4090,N_2631,N_2724);
nand U4091 (N_4091,N_3877,N_3396);
and U4092 (N_4092,N_2650,N_3638);
xnor U4093 (N_4093,N_2495,N_2372);
nand U4094 (N_4094,N_2337,N_2796);
xor U4095 (N_4095,N_3542,N_2100);
xnor U4096 (N_4096,N_2889,N_3195);
or U4097 (N_4097,N_2027,N_2997);
and U4098 (N_4098,N_2805,N_3148);
nor U4099 (N_4099,N_3818,N_2870);
xor U4100 (N_4100,N_2384,N_2733);
nor U4101 (N_4101,N_3223,N_2261);
nand U4102 (N_4102,N_3914,N_2795);
and U4103 (N_4103,N_3955,N_3984);
and U4104 (N_4104,N_2213,N_2223);
nand U4105 (N_4105,N_2949,N_2940);
nand U4106 (N_4106,N_2655,N_2572);
xnor U4107 (N_4107,N_2469,N_3741);
and U4108 (N_4108,N_2898,N_3016);
nand U4109 (N_4109,N_3451,N_2595);
and U4110 (N_4110,N_2297,N_2323);
or U4111 (N_4111,N_2984,N_2960);
or U4112 (N_4112,N_3420,N_2808);
and U4113 (N_4113,N_2915,N_2172);
or U4114 (N_4114,N_2208,N_2737);
or U4115 (N_4115,N_3314,N_3575);
and U4116 (N_4116,N_2155,N_3262);
nor U4117 (N_4117,N_3657,N_2127);
xor U4118 (N_4118,N_2676,N_3083);
and U4119 (N_4119,N_2684,N_2157);
nor U4120 (N_4120,N_3042,N_3189);
nand U4121 (N_4121,N_3907,N_3159);
nor U4122 (N_4122,N_3287,N_3375);
or U4123 (N_4123,N_2429,N_2446);
and U4124 (N_4124,N_2545,N_2905);
or U4125 (N_4125,N_2962,N_3249);
xnor U4126 (N_4126,N_3209,N_2068);
nor U4127 (N_4127,N_3855,N_3023);
nand U4128 (N_4128,N_3503,N_3677);
xnor U4129 (N_4129,N_2088,N_2828);
nor U4130 (N_4130,N_2824,N_3450);
and U4131 (N_4131,N_2943,N_2402);
xor U4132 (N_4132,N_3771,N_2780);
nand U4133 (N_4133,N_3763,N_2142);
nor U4134 (N_4134,N_2810,N_2229);
xnor U4135 (N_4135,N_2575,N_3637);
nor U4136 (N_4136,N_2831,N_3923);
nor U4137 (N_4137,N_2135,N_2566);
and U4138 (N_4138,N_3529,N_3369);
nand U4139 (N_4139,N_2000,N_2401);
xnor U4140 (N_4140,N_3240,N_3983);
or U4141 (N_4141,N_2183,N_3518);
nor U4142 (N_4142,N_3105,N_2149);
nor U4143 (N_4143,N_2874,N_2877);
and U4144 (N_4144,N_2602,N_3591);
xnor U4145 (N_4145,N_3065,N_3604);
and U4146 (N_4146,N_3037,N_2674);
nor U4147 (N_4147,N_2091,N_3218);
nand U4148 (N_4148,N_3624,N_3556);
nand U4149 (N_4149,N_2704,N_3557);
and U4150 (N_4150,N_2778,N_2348);
nand U4151 (N_4151,N_3102,N_2822);
nand U4152 (N_4152,N_3598,N_2070);
or U4153 (N_4153,N_2508,N_3835);
and U4154 (N_4154,N_2948,N_2661);
nor U4155 (N_4155,N_2406,N_2498);
nor U4156 (N_4156,N_2132,N_3075);
and U4157 (N_4157,N_2916,N_3891);
xnor U4158 (N_4158,N_3126,N_2911);
or U4159 (N_4159,N_2987,N_3664);
and U4160 (N_4160,N_3216,N_3999);
nand U4161 (N_4161,N_2031,N_2478);
nor U4162 (N_4162,N_3666,N_3959);
xor U4163 (N_4163,N_2090,N_3258);
nor U4164 (N_4164,N_2845,N_2934);
nor U4165 (N_4165,N_2579,N_2638);
xnor U4166 (N_4166,N_2825,N_2053);
or U4167 (N_4167,N_3339,N_3456);
or U4168 (N_4168,N_3968,N_3367);
nor U4169 (N_4169,N_3205,N_3662);
and U4170 (N_4170,N_2578,N_3663);
nand U4171 (N_4171,N_2584,N_3933);
nor U4172 (N_4172,N_3285,N_3379);
nor U4173 (N_4173,N_2505,N_2220);
and U4174 (N_4174,N_2443,N_2989);
or U4175 (N_4175,N_3405,N_3149);
nand U4176 (N_4176,N_3630,N_3494);
or U4177 (N_4177,N_2345,N_2865);
and U4178 (N_4178,N_2622,N_2671);
nand U4179 (N_4179,N_2488,N_3930);
or U4180 (N_4180,N_3866,N_3090);
nand U4181 (N_4181,N_2227,N_3193);
or U4182 (N_4182,N_2200,N_2537);
xnor U4183 (N_4183,N_3641,N_2158);
xor U4184 (N_4184,N_2921,N_2603);
xnor U4185 (N_4185,N_3550,N_2240);
and U4186 (N_4186,N_3535,N_3363);
and U4187 (N_4187,N_3301,N_3484);
nor U4188 (N_4188,N_3862,N_3789);
nand U4189 (N_4189,N_2108,N_3665);
nor U4190 (N_4190,N_3108,N_2025);
nand U4191 (N_4191,N_2936,N_3858);
or U4192 (N_4192,N_3745,N_2225);
and U4193 (N_4193,N_3059,N_2834);
nand U4194 (N_4194,N_3300,N_2050);
xnor U4195 (N_4195,N_3819,N_2769);
xor U4196 (N_4196,N_2884,N_3727);
nor U4197 (N_4197,N_2425,N_2470);
and U4198 (N_4198,N_2512,N_2658);
and U4199 (N_4199,N_3839,N_3602);
and U4200 (N_4200,N_2176,N_3337);
xor U4201 (N_4201,N_2460,N_3166);
or U4202 (N_4202,N_2727,N_2099);
xor U4203 (N_4203,N_3768,N_3512);
and U4204 (N_4204,N_3577,N_2363);
and U4205 (N_4205,N_3947,N_3773);
xnor U4206 (N_4206,N_2219,N_2596);
or U4207 (N_4207,N_2614,N_3926);
and U4208 (N_4208,N_2491,N_2526);
nor U4209 (N_4209,N_2616,N_3131);
and U4210 (N_4210,N_2882,N_3704);
xor U4211 (N_4211,N_3842,N_2121);
or U4212 (N_4212,N_3956,N_2479);
xor U4213 (N_4213,N_3817,N_3837);
nor U4214 (N_4214,N_2421,N_3725);
and U4215 (N_4215,N_3536,N_2935);
nor U4216 (N_4216,N_3180,N_2096);
nand U4217 (N_4217,N_3767,N_2419);
nand U4218 (N_4218,N_3951,N_2246);
and U4219 (N_4219,N_3432,N_3452);
and U4220 (N_4220,N_3614,N_2087);
or U4221 (N_4221,N_3815,N_2371);
or U4222 (N_4222,N_3764,N_2394);
xnor U4223 (N_4223,N_3691,N_2646);
xnor U4224 (N_4224,N_3203,N_3443);
nand U4225 (N_4225,N_3017,N_2799);
xnor U4226 (N_4226,N_2917,N_3305);
xnor U4227 (N_4227,N_3101,N_3809);
or U4228 (N_4228,N_3860,N_2642);
xor U4229 (N_4229,N_3215,N_3840);
or U4230 (N_4230,N_2409,N_3994);
or U4231 (N_4231,N_3272,N_2022);
nand U4232 (N_4232,N_2922,N_2999);
and U4233 (N_4233,N_3415,N_3573);
nor U4234 (N_4234,N_2423,N_2111);
xnor U4235 (N_4235,N_2293,N_3441);
or U4236 (N_4236,N_3632,N_2609);
xnor U4237 (N_4237,N_2599,N_2147);
nor U4238 (N_4238,N_2474,N_2500);
xor U4239 (N_4239,N_3022,N_2996);
or U4240 (N_4240,N_2690,N_3660);
nor U4241 (N_4241,N_2471,N_3754);
or U4242 (N_4242,N_3019,N_3060);
xnor U4243 (N_4243,N_3921,N_3546);
xnor U4244 (N_4244,N_2467,N_3797);
xnor U4245 (N_4245,N_2836,N_2329);
or U4246 (N_4246,N_2814,N_2092);
nand U4247 (N_4247,N_3394,N_2264);
or U4248 (N_4248,N_3121,N_3856);
nor U4249 (N_4249,N_2458,N_3590);
and U4250 (N_4250,N_2991,N_2427);
nand U4251 (N_4251,N_3470,N_3647);
nor U4252 (N_4252,N_3879,N_3317);
nor U4253 (N_4253,N_3242,N_2897);
nand U4254 (N_4254,N_3737,N_2803);
or U4255 (N_4255,N_3578,N_2003);
xnor U4256 (N_4256,N_3356,N_2527);
xnor U4257 (N_4257,N_3275,N_2490);
xnor U4258 (N_4258,N_2310,N_3461);
nor U4259 (N_4259,N_3878,N_2486);
nand U4260 (N_4260,N_3699,N_2017);
nand U4261 (N_4261,N_2693,N_2827);
xor U4262 (N_4262,N_2515,N_3289);
or U4263 (N_4263,N_2681,N_2744);
xnor U4264 (N_4264,N_3943,N_2871);
nor U4265 (N_4265,N_2785,N_2580);
nor U4266 (N_4266,N_3200,N_3116);
and U4267 (N_4267,N_3762,N_2782);
xnor U4268 (N_4268,N_2617,N_2259);
nor U4269 (N_4269,N_3712,N_3562);
nand U4270 (N_4270,N_2013,N_3003);
nor U4271 (N_4271,N_3235,N_2235);
nor U4272 (N_4272,N_2686,N_2324);
nand U4273 (N_4273,N_2946,N_3211);
and U4274 (N_4274,N_3327,N_2839);
or U4275 (N_4275,N_3498,N_3247);
xnor U4276 (N_4276,N_2494,N_2344);
nand U4277 (N_4277,N_2189,N_3045);
or U4278 (N_4278,N_3903,N_2481);
nand U4279 (N_4279,N_3125,N_2842);
nand U4280 (N_4280,N_2431,N_3120);
xor U4281 (N_4281,N_3689,N_3713);
xnor U4282 (N_4282,N_3905,N_2336);
nor U4283 (N_4283,N_2014,N_2790);
nor U4284 (N_4284,N_3306,N_3680);
or U4285 (N_4285,N_2995,N_2914);
xnor U4286 (N_4286,N_2417,N_3863);
and U4287 (N_4287,N_2024,N_2381);
nor U4288 (N_4288,N_3505,N_3832);
xor U4289 (N_4289,N_3154,N_3747);
xnor U4290 (N_4290,N_2206,N_3729);
nor U4291 (N_4291,N_3338,N_2411);
or U4292 (N_4292,N_3136,N_2872);
xnor U4293 (N_4293,N_3497,N_2403);
xnor U4294 (N_4294,N_2653,N_3260);
xnor U4295 (N_4295,N_3969,N_2282);
or U4296 (N_4296,N_2956,N_3576);
or U4297 (N_4297,N_2277,N_2789);
nor U4298 (N_4298,N_2464,N_3047);
nand U4299 (N_4299,N_2466,N_3640);
xor U4300 (N_4300,N_2424,N_2397);
and U4301 (N_4301,N_3890,N_3212);
or U4302 (N_4302,N_2151,N_3185);
nor U4303 (N_4303,N_2569,N_3281);
or U4304 (N_4304,N_2982,N_2120);
nor U4305 (N_4305,N_3579,N_2577);
xor U4306 (N_4306,N_2295,N_2585);
xnor U4307 (N_4307,N_2800,N_3612);
xor U4308 (N_4308,N_3902,N_3634);
or U4309 (N_4309,N_2433,N_2544);
and U4310 (N_4310,N_2391,N_2414);
or U4311 (N_4311,N_2055,N_3670);
or U4312 (N_4312,N_2573,N_2233);
nand U4313 (N_4313,N_3548,N_3124);
nor U4314 (N_4314,N_2986,N_3277);
and U4315 (N_4315,N_3511,N_2688);
and U4316 (N_4316,N_3474,N_2636);
or U4317 (N_4317,N_2838,N_3845);
or U4318 (N_4318,N_3990,N_3389);
and U4319 (N_4319,N_2722,N_2725);
and U4320 (N_4320,N_3897,N_3981);
xnor U4321 (N_4321,N_2813,N_2518);
nor U4322 (N_4322,N_2705,N_3373);
xor U4323 (N_4323,N_3304,N_2888);
nor U4324 (N_4324,N_2734,N_3276);
xor U4325 (N_4325,N_2489,N_2162);
and U4326 (N_4326,N_3791,N_3168);
xnor U4327 (N_4327,N_3111,N_3651);
nor U4328 (N_4328,N_3040,N_2863);
nand U4329 (N_4329,N_3523,N_3418);
nor U4330 (N_4330,N_2009,N_3977);
nor U4331 (N_4331,N_2112,N_3096);
and U4332 (N_4332,N_2104,N_3985);
or U4333 (N_4333,N_3954,N_2902);
and U4334 (N_4334,N_3748,N_2730);
nor U4335 (N_4335,N_3069,N_3774);
xor U4336 (N_4336,N_2496,N_2103);
and U4337 (N_4337,N_3122,N_3081);
or U4338 (N_4338,N_2383,N_2042);
or U4339 (N_4339,N_3700,N_2742);
nand U4340 (N_4340,N_3078,N_3001);
xor U4341 (N_4341,N_2747,N_3486);
or U4342 (N_4342,N_3872,N_3493);
xor U4343 (N_4343,N_3583,N_3833);
nand U4344 (N_4344,N_3046,N_2001);
and U4345 (N_4345,N_3739,N_3467);
and U4346 (N_4346,N_3318,N_3491);
xor U4347 (N_4347,N_3371,N_2855);
nor U4348 (N_4348,N_3757,N_2187);
and U4349 (N_4349,N_2663,N_2714);
or U4350 (N_4350,N_3468,N_2239);
nor U4351 (N_4351,N_2450,N_2307);
nand U4352 (N_4352,N_3399,N_2033);
nand U4353 (N_4353,N_2581,N_3229);
and U4354 (N_4354,N_2188,N_2380);
nand U4355 (N_4355,N_3867,N_3848);
nor U4356 (N_4356,N_3360,N_3939);
xnor U4357 (N_4357,N_3671,N_3052);
and U4358 (N_4358,N_3772,N_2198);
and U4359 (N_4359,N_3694,N_2783);
and U4360 (N_4360,N_3869,N_2359);
nor U4361 (N_4361,N_3411,N_2748);
nand U4362 (N_4362,N_2850,N_3345);
nor U4363 (N_4363,N_2468,N_2694);
nand U4364 (N_4364,N_3996,N_2807);
xor U4365 (N_4365,N_2150,N_3284);
and U4366 (N_4366,N_2501,N_3050);
xor U4367 (N_4367,N_2832,N_2720);
and U4368 (N_4368,N_2245,N_3071);
nand U4369 (N_4369,N_2657,N_3365);
nor U4370 (N_4370,N_3798,N_2018);
and U4371 (N_4371,N_3445,N_2444);
nor U4372 (N_4372,N_2502,N_3526);
and U4373 (N_4373,N_2951,N_2891);
nand U4374 (N_4374,N_3315,N_3353);
xnor U4375 (N_4375,N_3654,N_2028);
xnor U4376 (N_4376,N_2186,N_2767);
xnor U4377 (N_4377,N_3495,N_2482);
or U4378 (N_4378,N_2123,N_2843);
nand U4379 (N_4379,N_2878,N_2774);
nand U4380 (N_4380,N_2274,N_2131);
nor U4381 (N_4381,N_3457,N_2061);
nor U4382 (N_4382,N_3134,N_3898);
and U4383 (N_4383,N_3728,N_2304);
and U4384 (N_4384,N_3502,N_2258);
and U4385 (N_4385,N_3153,N_2228);
and U4386 (N_4386,N_2193,N_3979);
nor U4387 (N_4387,N_3310,N_2594);
and U4388 (N_4388,N_2238,N_2679);
or U4389 (N_4389,N_2553,N_3934);
and U4390 (N_4390,N_3292,N_2029);
or U4391 (N_4391,N_2032,N_3559);
or U4392 (N_4392,N_2939,N_2144);
nor U4393 (N_4393,N_2105,N_3246);
nand U4394 (N_4394,N_3534,N_3831);
or U4395 (N_4395,N_2990,N_3294);
or U4396 (N_4396,N_3909,N_3828);
and U4397 (N_4397,N_3342,N_2654);
nand U4398 (N_4398,N_2896,N_3717);
or U4399 (N_4399,N_3683,N_2568);
xor U4400 (N_4400,N_3421,N_2138);
and U4401 (N_4401,N_3874,N_2452);
nor U4402 (N_4402,N_2817,N_3513);
nor U4403 (N_4403,N_3135,N_3225);
or U4404 (N_4404,N_2360,N_2334);
and U4405 (N_4405,N_2196,N_3274);
xor U4406 (N_4406,N_2377,N_2992);
nand U4407 (N_4407,N_3732,N_2119);
or U4408 (N_4408,N_3409,N_2160);
or U4409 (N_4409,N_3182,N_2291);
and U4410 (N_4410,N_2130,N_3026);
nand U4411 (N_4411,N_3029,N_3253);
xnor U4412 (N_4412,N_2062,N_3650);
or U4413 (N_4413,N_2217,N_2528);
and U4414 (N_4414,N_3736,N_2361);
nor U4415 (N_4415,N_3092,N_3307);
and U4416 (N_4416,N_3783,N_2641);
nand U4417 (N_4417,N_2673,N_2630);
and U4418 (N_4418,N_3117,N_2185);
or U4419 (N_4419,N_2906,N_3838);
nor U4420 (N_4420,N_2574,N_2892);
nand U4421 (N_4421,N_3916,N_2637);
or U4422 (N_4422,N_3341,N_3521);
nor U4423 (N_4423,N_2289,N_3063);
or U4424 (N_4424,N_3433,N_3585);
nor U4425 (N_4425,N_3268,N_2036);
xor U4426 (N_4426,N_2645,N_2085);
xor U4427 (N_4427,N_2710,N_2369);
xnor U4428 (N_4428,N_3074,N_3416);
nor U4429 (N_4429,N_2290,N_3516);
nand U4430 (N_4430,N_3094,N_3678);
and U4431 (N_4431,N_3701,N_3463);
or U4432 (N_4432,N_3007,N_3077);
nor U4433 (N_4433,N_2919,N_2901);
and U4434 (N_4434,N_2804,N_2352);
and U4435 (N_4435,N_3806,N_3847);
nor U4436 (N_4436,N_2020,N_3465);
and U4437 (N_4437,N_2170,N_2947);
and U4438 (N_4438,N_3722,N_3312);
xor U4439 (N_4439,N_2776,N_3541);
nor U4440 (N_4440,N_2707,N_2094);
nor U4441 (N_4441,N_2485,N_3291);
and U4442 (N_4442,N_2434,N_2137);
nor U4443 (N_4443,N_3257,N_3582);
xor U4444 (N_4444,N_2538,N_2818);
or U4445 (N_4445,N_2442,N_2854);
and U4446 (N_4446,N_2101,N_2640);
nand U4447 (N_4447,N_3370,N_3619);
nand U4448 (N_4448,N_3133,N_3675);
and U4449 (N_4449,N_2081,N_3349);
nor U4450 (N_4450,N_2788,N_2672);
or U4451 (N_4451,N_2373,N_2270);
xor U4452 (N_4452,N_2841,N_3472);
and U4453 (N_4453,N_2350,N_3164);
nor U4454 (N_4454,N_3448,N_2766);
nor U4455 (N_4455,N_2677,N_3490);
and U4456 (N_4456,N_3015,N_3220);
nor U4457 (N_4457,N_2970,N_3412);
xnor U4458 (N_4458,N_3407,N_2953);
nor U4459 (N_4459,N_3928,N_3440);
or U4460 (N_4460,N_2392,N_3986);
or U4461 (N_4461,N_2719,N_2303);
nor U4462 (N_4462,N_2621,N_3519);
and U4463 (N_4463,N_3138,N_2660);
and U4464 (N_4464,N_2393,N_3567);
xnor U4465 (N_4465,N_2226,N_2076);
or U4466 (N_4466,N_3098,N_2422);
and U4467 (N_4467,N_3234,N_3270);
or U4468 (N_4468,N_2632,N_2124);
or U4469 (N_4469,N_3288,N_2950);
xor U4470 (N_4470,N_3237,N_3893);
nor U4471 (N_4471,N_2857,N_3147);
xnor U4472 (N_4472,N_2241,N_3836);
and U4473 (N_4473,N_3636,N_2060);
and U4474 (N_4474,N_3221,N_2317);
nand U4475 (N_4475,N_3733,N_3158);
nand U4476 (N_4476,N_2106,N_2601);
and U4477 (N_4477,N_2039,N_3068);
nor U4478 (N_4478,N_3401,N_3751);
nor U4479 (N_4479,N_3623,N_3615);
nor U4480 (N_4480,N_3621,N_3217);
and U4481 (N_4481,N_3611,N_2330);
xnor U4482 (N_4482,N_2963,N_2074);
and U4483 (N_4483,N_3130,N_3719);
and U4484 (N_4484,N_2907,N_3222);
nand U4485 (N_4485,N_3499,N_2629);
and U4486 (N_4486,N_3876,N_3661);
and U4487 (N_4487,N_2961,N_2399);
nor U4488 (N_4488,N_2968,N_2389);
and U4489 (N_4489,N_3896,N_3825);
nor U4490 (N_4490,N_3781,N_3478);
nor U4491 (N_4491,N_3659,N_2254);
xor U4492 (N_4492,N_3032,N_3794);
and U4493 (N_4493,N_3953,N_3392);
nand U4494 (N_4494,N_2558,N_3070);
or U4495 (N_4495,N_2449,N_3061);
or U4496 (N_4496,N_2430,N_2886);
and U4497 (N_4497,N_3199,N_3586);
nand U4498 (N_4498,N_2260,N_3788);
nor U4499 (N_4499,N_3254,N_3527);
xnor U4500 (N_4500,N_2556,N_2912);
nor U4501 (N_4501,N_2976,N_2619);
or U4502 (N_4502,N_3021,N_3089);
nand U4503 (N_4503,N_2318,N_2349);
nand U4504 (N_4504,N_2781,N_2844);
xnor U4505 (N_4505,N_2696,N_3230);
xor U4506 (N_4506,N_3740,N_3204);
nand U4507 (N_4507,N_2978,N_3350);
and U4508 (N_4508,N_2925,N_3020);
nand U4509 (N_4509,N_3311,N_3524);
xor U4510 (N_4510,N_3795,N_3018);
nand U4511 (N_4511,N_3476,N_3971);
or U4512 (N_4512,N_2689,N_2900);
and U4513 (N_4513,N_2715,N_2214);
and U4514 (N_4514,N_3803,N_3846);
and U4515 (N_4515,N_2590,N_2368);
xnor U4516 (N_4516,N_2881,N_3265);
or U4517 (N_4517,N_2570,N_2851);
xor U4518 (N_4518,N_3057,N_3496);
nand U4519 (N_4519,N_2164,N_3627);
or U4520 (N_4520,N_2005,N_2477);
nor U4521 (N_4521,N_3668,N_3790);
or U4522 (N_4522,N_2086,N_2952);
or U4523 (N_4523,N_3256,N_2199);
or U4524 (N_4524,N_3186,N_3635);
nor U4525 (N_4525,N_3264,N_3425);
nor U4526 (N_4526,N_2052,N_2903);
xnor U4527 (N_4527,N_3169,N_3201);
or U4528 (N_4528,N_3912,N_2294);
nor U4529 (N_4529,N_3698,N_2550);
and U4530 (N_4530,N_3500,N_3226);
nor U4531 (N_4531,N_3024,N_3174);
nand U4532 (N_4532,N_3989,N_2954);
nor U4533 (N_4533,N_3471,N_2669);
and U4534 (N_4534,N_3780,N_3469);
nor U4535 (N_4535,N_3946,N_2255);
nand U4536 (N_4536,N_3271,N_2625);
xor U4537 (N_4537,N_2412,N_2867);
or U4538 (N_4538,N_3162,N_2775);
or U4539 (N_4539,N_3572,N_3537);
nor U4540 (N_4540,N_3076,N_3183);
nand U4541 (N_4541,N_2521,N_2197);
nand U4542 (N_4542,N_3888,N_3384);
nand U4543 (N_4543,N_2750,N_3080);
and U4544 (N_4544,N_3477,N_3388);
nand U4545 (N_4545,N_2691,N_2316);
nand U4546 (N_4546,N_3859,N_3753);
and U4547 (N_4547,N_3854,N_3324);
and U4548 (N_4548,N_3267,N_3282);
and U4549 (N_4549,N_2139,N_2212);
or U4550 (N_4550,N_3173,N_2862);
and U4551 (N_4551,N_2211,N_3368);
nand U4552 (N_4552,N_3940,N_3853);
nor U4553 (N_4553,N_3648,N_3295);
or U4554 (N_4554,N_2387,N_3357);
nand U4555 (N_4555,N_3646,N_3581);
xnor U4556 (N_4556,N_2717,N_2205);
nor U4557 (N_4557,N_3901,N_2523);
and U4558 (N_4558,N_2510,N_3049);
nor U4559 (N_4559,N_3250,N_3900);
or U4560 (N_4560,N_3571,N_3008);
nor U4561 (N_4561,N_3397,N_2230);
xor U4562 (N_4562,N_2113,N_2746);
nand U4563 (N_4563,N_3894,N_2895);
nand U4564 (N_4564,N_2821,N_2152);
or U4565 (N_4565,N_2695,N_3383);
xor U4566 (N_4566,N_2335,N_3716);
and U4567 (N_4567,N_2847,N_2257);
or U4568 (N_4568,N_3255,N_3444);
nand U4569 (N_4569,N_3880,N_3937);
xor U4570 (N_4570,N_2701,N_2051);
nand U4571 (N_4571,N_2026,N_3233);
nand U4572 (N_4572,N_3653,N_3381);
nor U4573 (N_4573,N_3113,N_2066);
nor U4574 (N_4574,N_3455,N_2285);
nand U4575 (N_4575,N_3404,N_3028);
and U4576 (N_4576,N_3084,N_3179);
nand U4577 (N_4577,N_3889,N_2311);
nand U4578 (N_4578,N_3073,N_2593);
or U4579 (N_4579,N_2216,N_2107);
xnor U4580 (N_4580,N_3697,N_3553);
or U4581 (N_4581,N_3167,N_3427);
and U4582 (N_4582,N_2618,N_3629);
nor U4583 (N_4583,N_2784,N_2236);
and U4584 (N_4584,N_3643,N_2918);
and U4585 (N_4585,N_2483,N_2757);
and U4586 (N_4586,N_3938,N_3514);
nor U4587 (N_4587,N_3509,N_3278);
or U4588 (N_4588,N_2856,N_3196);
xnor U4589 (N_4589,N_3814,N_3742);
and U4590 (N_4590,N_3799,N_3165);
nand U4591 (N_4591,N_2256,N_2451);
nand U4592 (N_4592,N_2358,N_3447);
or U4593 (N_4593,N_2305,N_3231);
or U4594 (N_4594,N_2894,N_2347);
or U4595 (N_4595,N_3776,N_3091);
and U4596 (N_4596,N_2923,N_2077);
or U4597 (N_4597,N_3792,N_2125);
nor U4598 (N_4598,N_3066,N_2980);
xnor U4599 (N_4599,N_2635,N_2080);
and U4600 (N_4600,N_2519,N_3549);
nor U4601 (N_4601,N_3821,N_3316);
or U4602 (N_4602,N_2209,N_3283);
nand U4603 (N_4603,N_2168,N_3782);
nor U4604 (N_4604,N_3214,N_2969);
nor U4605 (N_4605,N_2242,N_3140);
xnor U4606 (N_4606,N_2959,N_2612);
nor U4607 (N_4607,N_3355,N_2148);
nand U4608 (N_4608,N_3376,N_2447);
or U4609 (N_4609,N_3568,N_3145);
xnor U4610 (N_4610,N_3473,N_3827);
nor U4611 (N_4611,N_2666,N_3726);
nor U4612 (N_4612,N_2286,N_2700);
or U4613 (N_4613,N_3813,N_2563);
nand U4614 (N_4614,N_2560,N_2351);
nand U4615 (N_4615,N_2487,N_2072);
or U4616 (N_4616,N_3925,N_3882);
nor U4617 (N_4617,N_2983,N_2548);
or U4618 (N_4618,N_2019,N_3600);
nand U4619 (N_4619,N_3885,N_2159);
nor U4620 (N_4620,N_2002,N_3302);
and U4621 (N_4621,N_3146,N_3434);
nand U4622 (N_4622,N_3208,N_3351);
nor U4623 (N_4623,N_3594,N_3013);
xnor U4624 (N_4624,N_2276,N_2231);
and U4625 (N_4625,N_2525,N_2035);
or U4626 (N_4626,N_2456,N_2977);
or U4627 (N_4627,N_2643,N_3333);
or U4628 (N_4628,N_3899,N_3436);
and U4629 (N_4629,N_2362,N_2278);
nand U4630 (N_4630,N_2732,N_2438);
xor U4631 (N_4631,N_3224,N_2222);
or U4632 (N_4632,N_3707,N_3099);
and U4633 (N_4633,N_2772,N_3431);
nor U4634 (N_4634,N_2114,N_3560);
or U4635 (N_4635,N_2794,N_3143);
and U4636 (N_4636,N_2448,N_3992);
and U4637 (N_4637,N_3446,N_3709);
nand U4638 (N_4638,N_2210,N_3644);
nand U4639 (N_4639,N_2492,N_3743);
nand U4640 (N_4640,N_3347,N_3177);
nand U4641 (N_4641,N_3163,N_3426);
and U4642 (N_4642,N_3033,N_2044);
nand U4643 (N_4643,N_3402,N_2702);
nand U4644 (N_4644,N_3358,N_2801);
nor U4645 (N_4645,N_2167,N_3348);
or U4646 (N_4646,N_2945,N_2268);
xnor U4647 (N_4647,N_2504,N_2866);
and U4648 (N_4648,N_2759,N_3501);
xor U4649 (N_4649,N_3944,N_2038);
xor U4650 (N_4650,N_2678,N_2820);
and U4651 (N_4651,N_3911,N_2899);
or U4652 (N_4652,N_2012,N_3686);
nand U4653 (N_4653,N_3403,N_3332);
or U4654 (N_4654,N_3682,N_2253);
nor U4655 (N_4655,N_2529,N_2342);
nor U4656 (N_4656,N_2752,N_2191);
and U4657 (N_4657,N_2682,N_3194);
or U4658 (N_4658,N_2607,N_3398);
or U4659 (N_4659,N_3352,N_2942);
xor U4660 (N_4660,N_2117,N_2215);
nand U4661 (N_4661,N_3335,N_2366);
or U4662 (N_4662,N_2583,N_2706);
or U4663 (N_4663,N_2861,N_3980);
nand U4664 (N_4664,N_2190,N_2514);
or U4665 (N_4665,N_2078,N_2567);
nor U4666 (N_4666,N_2516,N_3118);
xnor U4667 (N_4667,N_3479,N_3103);
and U4668 (N_4668,N_2390,N_3645);
nand U4669 (N_4669,N_2382,N_3929);
and U4670 (N_4670,N_2555,N_3034);
nor U4671 (N_4671,N_2649,N_2540);
nor U4672 (N_4672,N_3734,N_2326);
or U4673 (N_4673,N_2375,N_3964);
xor U4674 (N_4674,N_2941,N_3141);
nand U4675 (N_4675,N_3865,N_3850);
xor U4676 (N_4676,N_3067,N_3043);
or U4677 (N_4677,N_2770,N_3871);
and U4678 (N_4678,N_3064,N_2493);
or U4679 (N_4679,N_3808,N_3172);
and U4680 (N_4680,N_3695,N_3759);
nand U4681 (N_4681,N_3430,N_3758);
nand U4682 (N_4682,N_2204,N_3963);
nor U4683 (N_4683,N_2249,N_3012);
nand U4684 (N_4684,N_3128,N_3669);
nor U4685 (N_4685,N_2069,N_2340);
and U4686 (N_4686,N_3184,N_3540);
or U4687 (N_4687,N_3545,N_2332);
nor U4688 (N_4688,N_2541,N_2852);
xor U4689 (N_4689,N_3082,N_2811);
nand U4690 (N_4690,N_2309,N_2994);
xnor U4691 (N_4691,N_3155,N_2615);
nand U4692 (N_4692,N_2972,N_3462);
xnor U4693 (N_4693,N_3919,N_3051);
and U4694 (N_4694,N_2539,N_3010);
nand U4695 (N_4695,N_3533,N_2046);
or U4696 (N_4696,N_2079,N_2016);
or U4697 (N_4697,N_2272,N_2461);
and U4698 (N_4698,N_3547,N_2712);
nor U4699 (N_4699,N_3924,N_3685);
nor U4700 (N_4700,N_2740,N_2806);
nand U4701 (N_4701,N_3085,N_3972);
nor U4702 (N_4702,N_2175,N_2306);
nand U4703 (N_4703,N_2166,N_3192);
and U4704 (N_4704,N_2532,N_3693);
nor U4705 (N_4705,N_3606,N_2754);
and U4706 (N_4706,N_2731,N_2910);
and U4707 (N_4707,N_2095,N_2313);
nand U4708 (N_4708,N_3438,N_3236);
nor U4709 (N_4709,N_3551,N_3744);
nor U4710 (N_4710,N_3945,N_2530);
xnor U4711 (N_4711,N_2662,N_2944);
xnor U4712 (N_4712,N_2605,N_3419);
and U4713 (N_4713,N_3391,N_3626);
or U4714 (N_4714,N_2146,N_2762);
xnor U4715 (N_4715,N_2931,N_3908);
nor U4716 (N_4716,N_2302,N_3086);
nor U4717 (N_4717,N_2589,N_3107);
or U4718 (N_4718,N_2161,N_3152);
nor U4719 (N_4719,N_3320,N_2413);
or U4720 (N_4720,N_3750,N_2604);
xor U4721 (N_4721,N_3507,N_2007);
or U4722 (N_4722,N_3779,N_2040);
xnor U4723 (N_4723,N_3156,N_2753);
xnor U4724 (N_4724,N_3344,N_2559);
xor U4725 (N_4725,N_2102,N_2557);
and U4726 (N_4726,N_2484,N_2571);
and U4727 (N_4727,N_2439,N_2979);
or U4728 (N_4728,N_3609,N_3708);
or U4729 (N_4729,N_3110,N_2388);
xnor U4730 (N_4730,N_3492,N_3408);
and U4731 (N_4731,N_3439,N_2880);
xor U4732 (N_4732,N_2723,N_3385);
nand U4733 (N_4733,N_2184,N_3649);
or U4734 (N_4734,N_3566,N_3816);
nand U4735 (N_4735,N_3530,N_3025);
or U4736 (N_4736,N_3014,N_2554);
nand U4737 (N_4737,N_2418,N_2773);
xnor U4738 (N_4738,N_3690,N_3705);
nand U4739 (N_4739,N_2357,N_3993);
or U4740 (N_4740,N_3386,N_2549);
nand U4741 (N_4741,N_2312,N_2296);
or U4742 (N_4742,N_2252,N_3506);
or U4743 (N_4743,N_3730,N_2713);
nand U4744 (N_4744,N_3326,N_2244);
or U4745 (N_4745,N_2426,N_3104);
xor U4746 (N_4746,N_2864,N_2763);
and U4747 (N_4747,N_3058,N_2958);
nand U4748 (N_4748,N_2873,N_3406);
or U4749 (N_4749,N_2353,N_2535);
xnor U4750 (N_4750,N_3633,N_3362);
nor U4751 (N_4751,N_3702,N_2633);
nor U4752 (N_4752,N_3978,N_3176);
nand U4753 (N_4753,N_2587,N_3228);
xnor U4754 (N_4754,N_2685,N_2435);
and U4755 (N_4755,N_2974,N_2420);
xnor U4756 (N_4756,N_2288,N_2552);
nor U4757 (N_4757,N_3009,N_3610);
or U4758 (N_4758,N_2509,N_2812);
and U4759 (N_4759,N_2355,N_3824);
or U4760 (N_4760,N_3622,N_3721);
and U4761 (N_4761,N_3044,N_2030);
or U4762 (N_4762,N_3807,N_2365);
nand U4763 (N_4763,N_2680,N_2021);
and U4764 (N_4764,N_3487,N_2262);
or U4765 (N_4765,N_2760,N_3187);
or U4766 (N_4766,N_2181,N_3508);
nor U4767 (N_4767,N_2457,N_2728);
nand U4768 (N_4768,N_3039,N_2266);
and U4769 (N_4769,N_2315,N_3414);
nand U4770 (N_4770,N_3041,N_2396);
xnor U4771 (N_4771,N_2793,N_3881);
xnor U4772 (N_4772,N_3970,N_3711);
nand U4773 (N_4773,N_2858,N_2965);
nand U4774 (N_4774,N_3510,N_2967);
xnor U4775 (N_4775,N_2522,N_3595);
nor U4776 (N_4776,N_2071,N_2462);
or U4777 (N_4777,N_2201,N_3995);
and U4778 (N_4778,N_3895,N_3528);
nor U4779 (N_4779,N_2440,N_3973);
xor U4780 (N_4780,N_2835,N_2928);
nand U4781 (N_4781,N_2708,N_2321);
or U4782 (N_4782,N_2156,N_3787);
xnor U4783 (N_4783,N_2432,N_3770);
xor U4784 (N_4784,N_2665,N_2178);
and U4785 (N_4785,N_2385,N_2265);
xor U4786 (N_4786,N_3687,N_2973);
xor U4787 (N_4787,N_3532,N_3617);
nand U4788 (N_4788,N_2777,N_2600);
nor U4789 (N_4789,N_3587,N_2174);
xnor U4790 (N_4790,N_3340,N_2860);
nand U4791 (N_4791,N_3904,N_2287);
nand U4792 (N_4792,N_2791,N_2699);
xnor U4793 (N_4793,N_3688,N_2405);
nand U4794 (N_4794,N_3658,N_2063);
xnor U4795 (N_4795,N_2292,N_3829);
and U4796 (N_4796,N_2379,N_3273);
or U4797 (N_4797,N_2275,N_2023);
nand U4798 (N_4798,N_3696,N_3804);
or U4799 (N_4799,N_3957,N_3109);
and U4800 (N_4800,N_2169,N_3906);
or U4801 (N_4801,N_2981,N_2221);
nand U4802 (N_4802,N_2930,N_2764);
and U4803 (N_4803,N_2823,N_2826);
nor U4804 (N_4804,N_2415,N_3543);
xnor U4805 (N_4805,N_3170,N_2543);
xor U4806 (N_4806,N_3935,N_3361);
or U4807 (N_4807,N_2771,N_2765);
nor U4808 (N_4808,N_2768,N_2378);
nand U4809 (N_4809,N_3191,N_3724);
nand U4810 (N_4810,N_3038,N_3749);
and U4811 (N_4811,N_2065,N_2097);
xnor U4812 (N_4812,N_3142,N_3778);
nor U4813 (N_4813,N_3884,N_2507);
xnor U4814 (N_4814,N_2533,N_2904);
and U4815 (N_4815,N_2006,N_2056);
nand U4816 (N_4816,N_2756,N_3965);
nor U4817 (N_4817,N_2816,N_2346);
or U4818 (N_4818,N_3531,N_3380);
or U4819 (N_4819,N_3563,N_2370);
nor U4820 (N_4820,N_3710,N_3720);
xor U4821 (N_4821,N_2517,N_2089);
nor U4822 (N_4822,N_2143,N_2966);
nand U4823 (N_4823,N_2608,N_3599);
or U4824 (N_4824,N_2837,N_3207);
xnor U4825 (N_4825,N_2703,N_2404);
and U4826 (N_4826,N_2263,N_2251);
nand U4827 (N_4827,N_2933,N_2606);
nand U4828 (N_4828,N_3261,N_3417);
nor U4829 (N_4829,N_2015,N_2749);
nand U4830 (N_4830,N_3313,N_3482);
or U4831 (N_4831,N_3812,N_3197);
and U4832 (N_4832,N_3359,N_2926);
xnor U4833 (N_4833,N_2048,N_3976);
nor U4834 (N_4834,N_2506,N_3202);
nor U4835 (N_4835,N_2745,N_3830);
nor U4836 (N_4836,N_3303,N_3618);
and U4837 (N_4837,N_2644,N_3681);
xor U4838 (N_4838,N_3132,N_2542);
nor U4839 (N_4839,N_2624,N_3715);
nand U4840 (N_4840,N_2652,N_3589);
xor U4841 (N_4841,N_3870,N_2562);
or U4842 (N_4842,N_3883,N_3150);
xnor U4843 (N_4843,N_2237,N_2356);
and U4844 (N_4844,N_3752,N_2122);
and U4845 (N_4845,N_3564,N_3244);
xnor U4846 (N_4846,N_2592,N_2367);
nor U4847 (N_4847,N_2280,N_2546);
or U4848 (N_4848,N_3160,N_2830);
and U4849 (N_4849,N_3374,N_2299);
nand U4850 (N_4850,N_3525,N_2093);
nor U4851 (N_4851,N_3843,N_3263);
and U4852 (N_4852,N_2118,N_3826);
nor U4853 (N_4853,N_3756,N_3975);
or U4854 (N_4854,N_2809,N_3558);
nor U4855 (N_4855,N_3608,N_2751);
nor U4856 (N_4856,N_2536,N_2475);
nor U4857 (N_4857,N_3593,N_3372);
or U4858 (N_4858,N_2194,N_3062);
nor U4859 (N_4859,N_3259,N_3982);
nand U4860 (N_4860,N_2726,N_3539);
xnor U4861 (N_4861,N_2890,N_3106);
xnor U4862 (N_4862,N_3053,N_3139);
xor U4863 (N_4863,N_3449,N_2284);
nand U4864 (N_4864,N_3378,N_3437);
nor U4865 (N_4865,N_2988,N_3442);
or U4866 (N_4866,N_3642,N_3601);
nor U4867 (N_4867,N_3480,N_3178);
or U4868 (N_4868,N_2328,N_3515);
xnor U4869 (N_4869,N_3857,N_3517);
and U4870 (N_4870,N_3321,N_3625);
or U4871 (N_4871,N_3886,N_2084);
or U4872 (N_4872,N_2833,N_2043);
and U4873 (N_4873,N_2224,N_3035);
nor U4874 (N_4874,N_3841,N_3997);
nand U4875 (N_4875,N_2929,N_2846);
nand U4876 (N_4876,N_2819,N_2083);
and U4877 (N_4877,N_3849,N_2698);
nor U4878 (N_4878,N_2576,N_2243);
xnor U4879 (N_4879,N_3079,N_2588);
and U4880 (N_4880,N_3723,N_3213);
or U4881 (N_4881,N_2664,N_3998);
or U4882 (N_4882,N_3755,N_3175);
or U4883 (N_4883,N_3958,N_3238);
xor U4884 (N_4884,N_3656,N_2610);
xnor U4885 (N_4885,N_2993,N_2531);
and U4886 (N_4886,N_2924,N_3605);
nand U4887 (N_4887,N_3607,N_3769);
or U4888 (N_4888,N_3330,N_2459);
and U4889 (N_4889,N_2883,N_2848);
nor U4890 (N_4890,N_3157,N_3961);
nor U4891 (N_4891,N_2908,N_2547);
xnor U4892 (N_4892,N_3119,N_3097);
and U4893 (N_4893,N_2971,N_2659);
nand U4894 (N_4894,N_3429,N_2647);
nand U4895 (N_4895,N_2300,N_3676);
and U4896 (N_4896,N_3251,N_2786);
nand U4897 (N_4897,N_2037,N_3974);
nor U4898 (N_4898,N_3005,N_3703);
nor U4899 (N_4899,N_2697,N_2736);
or U4900 (N_4900,N_2234,N_2129);
and U4901 (N_4901,N_3056,N_3801);
xor U4902 (N_4902,N_3868,N_3746);
or U4903 (N_4903,N_3936,N_2455);
or U4904 (N_4904,N_2400,N_2059);
nand U4905 (N_4905,N_3927,N_2582);
nand U4906 (N_4906,N_3100,N_2408);
xor U4907 (N_4907,N_2116,N_3115);
nand U4908 (N_4908,N_3137,N_3319);
or U4909 (N_4909,N_3603,N_2687);
or U4910 (N_4910,N_2058,N_2109);
or U4911 (N_4911,N_3298,N_2551);
xnor U4912 (N_4912,N_3760,N_3674);
nor U4913 (N_4913,N_3639,N_2283);
nor U4914 (N_4914,N_2453,N_3597);
nor U4915 (N_4915,N_3428,N_2670);
nand U4916 (N_4916,N_3161,N_3054);
xnor U4917 (N_4917,N_2721,N_2269);
xnor U4918 (N_4918,N_2985,N_2126);
or U4919 (N_4919,N_3095,N_3048);
nor U4920 (N_4920,N_2333,N_2975);
xnor U4921 (N_4921,N_2203,N_2957);
nand U4922 (N_4922,N_2398,N_3873);
or U4923 (N_4923,N_2853,N_3544);
or U4924 (N_4924,N_3299,N_3802);
and U4925 (N_4925,N_3766,N_3805);
nand U4926 (N_4926,N_3293,N_2248);
or U4927 (N_4927,N_3706,N_2325);
or U4928 (N_4928,N_3822,N_2735);
xnor U4929 (N_4929,N_2628,N_3922);
xor U4930 (N_4930,N_2623,N_3834);
or U4931 (N_4931,N_3481,N_3588);
nand U4932 (N_4932,N_3875,N_3088);
nor U4933 (N_4933,N_2386,N_2620);
nor U4934 (N_4934,N_3488,N_3435);
or U4935 (N_4935,N_3520,N_3266);
nor U4936 (N_4936,N_2428,N_3325);
nor U4937 (N_4937,N_2561,N_3673);
nor U4938 (N_4938,N_2718,N_2437);
or U4939 (N_4939,N_2964,N_3966);
nor U4940 (N_4940,N_2319,N_2247);
nand U4941 (N_4941,N_3918,N_3584);
nand U4942 (N_4942,N_3962,N_3786);
nor U4943 (N_4943,N_2010,N_2711);
or U4944 (N_4944,N_2729,N_3932);
or U4945 (N_4945,N_2250,N_2741);
nand U4946 (N_4946,N_2134,N_2047);
nor U4947 (N_4947,N_2320,N_3887);
nand U4948 (N_4948,N_3002,N_2639);
nor U4949 (N_4949,N_3006,N_3941);
xnor U4950 (N_4950,N_2180,N_2565);
nor U4951 (N_4951,N_2868,N_3219);
and U4952 (N_4952,N_2937,N_2586);
or U4953 (N_4953,N_2416,N_2232);
or U4954 (N_4954,N_3522,N_2338);
nand U4955 (N_4955,N_3561,N_2327);
nand U4956 (N_4956,N_2314,N_3504);
and U4957 (N_4957,N_2376,N_3297);
xor U4958 (N_4958,N_2298,N_3424);
and U4959 (N_4959,N_3810,N_2709);
and U4960 (N_4960,N_2173,N_3245);
nor U4961 (N_4961,N_3364,N_2879);
or U4962 (N_4962,N_3948,N_3667);
or U4963 (N_4963,N_2465,N_3151);
nor U4964 (N_4964,N_2177,N_3422);
and U4965 (N_4965,N_3915,N_2281);
nand U4966 (N_4966,N_2182,N_3811);
or U4967 (N_4967,N_2407,N_3861);
and U4968 (N_4968,N_2133,N_3248);
nor U4969 (N_4969,N_3286,N_3190);
nor U4970 (N_4970,N_2564,N_2998);
and U4971 (N_4971,N_3453,N_3454);
and U4972 (N_4972,N_3844,N_3466);
nor U4973 (N_4973,N_3336,N_2141);
nand U4974 (N_4974,N_2011,N_2876);
nand U4975 (N_4975,N_3485,N_3322);
or U4976 (N_4976,N_3569,N_2627);
xor U4977 (N_4977,N_3718,N_2758);
or U4978 (N_4978,N_2273,N_2743);
nand U4979 (N_4979,N_3269,N_3144);
and U4980 (N_4980,N_2859,N_2668);
nand U4981 (N_4981,N_3114,N_3851);
xnor U4982 (N_4982,N_3538,N_3777);
nor U4983 (N_4983,N_2054,N_2301);
xnor U4984 (N_4984,N_3820,N_3464);
nand U4985 (N_4985,N_2279,N_2739);
or U4986 (N_4986,N_2716,N_2503);
nor U4987 (N_4987,N_2082,N_2410);
nand U4988 (N_4988,N_2511,N_3055);
and U4989 (N_4989,N_2598,N_2436);
or U4990 (N_4990,N_2692,N_2136);
and U4991 (N_4991,N_3489,N_3823);
or U4992 (N_4992,N_3631,N_2480);
nand U4993 (N_4993,N_3413,N_3761);
nor U4994 (N_4994,N_3346,N_3460);
or U4995 (N_4995,N_2787,N_3206);
and U4996 (N_4996,N_3679,N_2145);
nor U4997 (N_4997,N_3684,N_3323);
xnor U4998 (N_4998,N_3354,N_3382);
xnor U4999 (N_4999,N_2473,N_2364);
and U5000 (N_5000,N_2310,N_2051);
nand U5001 (N_5001,N_3814,N_2961);
nand U5002 (N_5002,N_3436,N_3968);
xnor U5003 (N_5003,N_3805,N_3711);
xnor U5004 (N_5004,N_2922,N_3075);
xnor U5005 (N_5005,N_3666,N_3658);
or U5006 (N_5006,N_3037,N_2510);
nor U5007 (N_5007,N_2229,N_2722);
nand U5008 (N_5008,N_3721,N_2341);
nand U5009 (N_5009,N_3406,N_2869);
nand U5010 (N_5010,N_3579,N_3967);
and U5011 (N_5011,N_2565,N_3759);
nand U5012 (N_5012,N_3473,N_2400);
nor U5013 (N_5013,N_3402,N_3672);
and U5014 (N_5014,N_3806,N_3055);
nor U5015 (N_5015,N_2761,N_3029);
or U5016 (N_5016,N_3346,N_3053);
xor U5017 (N_5017,N_3786,N_3245);
xor U5018 (N_5018,N_3053,N_2899);
nor U5019 (N_5019,N_3979,N_2488);
or U5020 (N_5020,N_3240,N_3091);
and U5021 (N_5021,N_2871,N_2299);
nand U5022 (N_5022,N_3978,N_2626);
or U5023 (N_5023,N_2910,N_3018);
nand U5024 (N_5024,N_3244,N_2220);
nor U5025 (N_5025,N_3314,N_3161);
xor U5026 (N_5026,N_3098,N_3990);
nand U5027 (N_5027,N_2742,N_3263);
xnor U5028 (N_5028,N_3172,N_2332);
nand U5029 (N_5029,N_3647,N_3198);
and U5030 (N_5030,N_2492,N_3103);
and U5031 (N_5031,N_3900,N_2156);
nor U5032 (N_5032,N_3746,N_2272);
nand U5033 (N_5033,N_3985,N_2657);
nand U5034 (N_5034,N_3941,N_2060);
or U5035 (N_5035,N_2792,N_2493);
and U5036 (N_5036,N_2190,N_2463);
or U5037 (N_5037,N_2259,N_2284);
and U5038 (N_5038,N_3840,N_3783);
xor U5039 (N_5039,N_2720,N_2302);
or U5040 (N_5040,N_3130,N_2183);
nor U5041 (N_5041,N_3426,N_3366);
nor U5042 (N_5042,N_3402,N_3606);
nor U5043 (N_5043,N_2492,N_2281);
nand U5044 (N_5044,N_3997,N_2330);
or U5045 (N_5045,N_3112,N_3804);
and U5046 (N_5046,N_3165,N_2473);
nor U5047 (N_5047,N_3146,N_2531);
nand U5048 (N_5048,N_2295,N_2192);
xnor U5049 (N_5049,N_2664,N_3650);
xnor U5050 (N_5050,N_2897,N_3297);
and U5051 (N_5051,N_3708,N_2948);
xor U5052 (N_5052,N_2751,N_2476);
nor U5053 (N_5053,N_2525,N_3891);
xor U5054 (N_5054,N_3181,N_3411);
or U5055 (N_5055,N_3404,N_2032);
xor U5056 (N_5056,N_3837,N_2953);
nor U5057 (N_5057,N_3711,N_3531);
nand U5058 (N_5058,N_2093,N_3212);
xnor U5059 (N_5059,N_3837,N_3659);
nand U5060 (N_5060,N_3310,N_2593);
xnor U5061 (N_5061,N_3419,N_2147);
nand U5062 (N_5062,N_3981,N_2886);
and U5063 (N_5063,N_3702,N_3538);
and U5064 (N_5064,N_2584,N_3481);
or U5065 (N_5065,N_2039,N_3176);
and U5066 (N_5066,N_2549,N_3232);
xor U5067 (N_5067,N_2679,N_3582);
or U5068 (N_5068,N_2337,N_3000);
nor U5069 (N_5069,N_2941,N_2624);
nor U5070 (N_5070,N_3901,N_3531);
nor U5071 (N_5071,N_2165,N_2133);
nand U5072 (N_5072,N_2740,N_2043);
xor U5073 (N_5073,N_3395,N_2097);
xnor U5074 (N_5074,N_2917,N_3298);
and U5075 (N_5075,N_2443,N_2139);
nand U5076 (N_5076,N_3546,N_2619);
or U5077 (N_5077,N_3890,N_2153);
nor U5078 (N_5078,N_3489,N_3663);
and U5079 (N_5079,N_2279,N_2561);
and U5080 (N_5080,N_3408,N_2076);
and U5081 (N_5081,N_2736,N_3400);
nor U5082 (N_5082,N_2477,N_3226);
nor U5083 (N_5083,N_2379,N_2945);
nand U5084 (N_5084,N_2472,N_2059);
xnor U5085 (N_5085,N_3925,N_2426);
nand U5086 (N_5086,N_3673,N_2668);
nand U5087 (N_5087,N_2777,N_2353);
and U5088 (N_5088,N_3251,N_2899);
and U5089 (N_5089,N_2904,N_2070);
or U5090 (N_5090,N_3786,N_3274);
or U5091 (N_5091,N_3158,N_3769);
nand U5092 (N_5092,N_2766,N_3807);
nand U5093 (N_5093,N_2895,N_2369);
nand U5094 (N_5094,N_2721,N_3943);
nor U5095 (N_5095,N_3469,N_2386);
and U5096 (N_5096,N_3715,N_2384);
or U5097 (N_5097,N_2368,N_2345);
nand U5098 (N_5098,N_2096,N_2238);
nand U5099 (N_5099,N_2630,N_2146);
nand U5100 (N_5100,N_3172,N_3142);
or U5101 (N_5101,N_3990,N_2958);
and U5102 (N_5102,N_2376,N_2353);
and U5103 (N_5103,N_2877,N_2252);
or U5104 (N_5104,N_3557,N_3641);
xor U5105 (N_5105,N_3038,N_3414);
nor U5106 (N_5106,N_2032,N_2922);
nand U5107 (N_5107,N_2825,N_3228);
xnor U5108 (N_5108,N_3532,N_3210);
and U5109 (N_5109,N_3235,N_3342);
and U5110 (N_5110,N_3521,N_2213);
xor U5111 (N_5111,N_3761,N_3094);
nand U5112 (N_5112,N_2963,N_3396);
nor U5113 (N_5113,N_2174,N_2084);
and U5114 (N_5114,N_3749,N_3237);
and U5115 (N_5115,N_2581,N_2267);
and U5116 (N_5116,N_2319,N_2739);
xnor U5117 (N_5117,N_2763,N_3813);
or U5118 (N_5118,N_2958,N_3914);
or U5119 (N_5119,N_2868,N_2197);
nand U5120 (N_5120,N_2634,N_2220);
nand U5121 (N_5121,N_3351,N_3239);
nor U5122 (N_5122,N_2646,N_3379);
nor U5123 (N_5123,N_3767,N_2003);
xor U5124 (N_5124,N_3474,N_3052);
nand U5125 (N_5125,N_2252,N_3011);
or U5126 (N_5126,N_2129,N_2987);
nor U5127 (N_5127,N_3452,N_3273);
or U5128 (N_5128,N_2730,N_2939);
nor U5129 (N_5129,N_2923,N_2188);
nand U5130 (N_5130,N_2390,N_2849);
or U5131 (N_5131,N_2330,N_2064);
and U5132 (N_5132,N_3852,N_2278);
nor U5133 (N_5133,N_3192,N_3865);
and U5134 (N_5134,N_2956,N_3456);
and U5135 (N_5135,N_3447,N_2729);
nand U5136 (N_5136,N_3881,N_3138);
and U5137 (N_5137,N_2955,N_2808);
and U5138 (N_5138,N_2719,N_3021);
nor U5139 (N_5139,N_3187,N_2671);
and U5140 (N_5140,N_2036,N_3255);
nor U5141 (N_5141,N_3747,N_3454);
or U5142 (N_5142,N_2253,N_3911);
xor U5143 (N_5143,N_2329,N_3148);
nor U5144 (N_5144,N_2026,N_2133);
nor U5145 (N_5145,N_2683,N_2069);
nor U5146 (N_5146,N_3556,N_2213);
nand U5147 (N_5147,N_2229,N_3958);
and U5148 (N_5148,N_3218,N_2560);
xnor U5149 (N_5149,N_3398,N_3217);
or U5150 (N_5150,N_2789,N_3054);
or U5151 (N_5151,N_3960,N_2533);
nand U5152 (N_5152,N_2963,N_3363);
xor U5153 (N_5153,N_2325,N_3055);
and U5154 (N_5154,N_3628,N_3088);
nor U5155 (N_5155,N_3402,N_3765);
nor U5156 (N_5156,N_2668,N_3935);
and U5157 (N_5157,N_2265,N_3403);
xor U5158 (N_5158,N_3692,N_2345);
nor U5159 (N_5159,N_2190,N_2763);
nor U5160 (N_5160,N_2944,N_2173);
xnor U5161 (N_5161,N_3375,N_2080);
nor U5162 (N_5162,N_3443,N_3703);
nor U5163 (N_5163,N_2493,N_3003);
nor U5164 (N_5164,N_2137,N_2709);
nor U5165 (N_5165,N_3349,N_2237);
nand U5166 (N_5166,N_3715,N_2004);
and U5167 (N_5167,N_2743,N_3363);
or U5168 (N_5168,N_3775,N_3593);
nand U5169 (N_5169,N_3020,N_3188);
nor U5170 (N_5170,N_2274,N_2229);
xnor U5171 (N_5171,N_2802,N_2420);
xor U5172 (N_5172,N_3729,N_2212);
nand U5173 (N_5173,N_2639,N_3414);
xor U5174 (N_5174,N_2646,N_3847);
nor U5175 (N_5175,N_2792,N_2410);
xor U5176 (N_5176,N_2791,N_3270);
or U5177 (N_5177,N_3013,N_2926);
xor U5178 (N_5178,N_3197,N_2787);
nor U5179 (N_5179,N_2294,N_3727);
or U5180 (N_5180,N_3945,N_3486);
nor U5181 (N_5181,N_3923,N_3764);
nand U5182 (N_5182,N_3425,N_2002);
or U5183 (N_5183,N_3997,N_2636);
xor U5184 (N_5184,N_2780,N_2329);
or U5185 (N_5185,N_3564,N_2096);
xnor U5186 (N_5186,N_2067,N_2346);
nand U5187 (N_5187,N_2102,N_2230);
nor U5188 (N_5188,N_3323,N_3883);
nand U5189 (N_5189,N_2675,N_3090);
nand U5190 (N_5190,N_2733,N_3654);
nor U5191 (N_5191,N_2108,N_3999);
and U5192 (N_5192,N_3075,N_3249);
and U5193 (N_5193,N_3466,N_3836);
xor U5194 (N_5194,N_3627,N_3232);
nor U5195 (N_5195,N_3994,N_3068);
xnor U5196 (N_5196,N_2113,N_2019);
and U5197 (N_5197,N_2436,N_2152);
xnor U5198 (N_5198,N_2431,N_3419);
nor U5199 (N_5199,N_2177,N_3587);
xor U5200 (N_5200,N_2969,N_2926);
nor U5201 (N_5201,N_3341,N_2022);
nor U5202 (N_5202,N_2665,N_3423);
nor U5203 (N_5203,N_3290,N_2653);
nand U5204 (N_5204,N_3079,N_3153);
and U5205 (N_5205,N_2728,N_2017);
nor U5206 (N_5206,N_2797,N_3131);
xor U5207 (N_5207,N_2945,N_3566);
xnor U5208 (N_5208,N_2836,N_3566);
nor U5209 (N_5209,N_2280,N_3339);
xnor U5210 (N_5210,N_3541,N_3970);
xor U5211 (N_5211,N_3846,N_3685);
or U5212 (N_5212,N_3121,N_2060);
or U5213 (N_5213,N_2855,N_3103);
or U5214 (N_5214,N_3907,N_3178);
nand U5215 (N_5215,N_3060,N_2091);
nand U5216 (N_5216,N_2558,N_3616);
nand U5217 (N_5217,N_2533,N_3842);
or U5218 (N_5218,N_2601,N_2489);
xnor U5219 (N_5219,N_2251,N_2936);
nand U5220 (N_5220,N_3547,N_3877);
and U5221 (N_5221,N_3012,N_2441);
nor U5222 (N_5222,N_3064,N_2443);
nor U5223 (N_5223,N_3656,N_3838);
or U5224 (N_5224,N_2582,N_3986);
xnor U5225 (N_5225,N_2512,N_2632);
or U5226 (N_5226,N_2303,N_2252);
nand U5227 (N_5227,N_2690,N_3696);
or U5228 (N_5228,N_2733,N_3215);
nor U5229 (N_5229,N_3393,N_2885);
nand U5230 (N_5230,N_2983,N_2471);
or U5231 (N_5231,N_3528,N_3915);
or U5232 (N_5232,N_3401,N_3869);
xnor U5233 (N_5233,N_3399,N_3729);
and U5234 (N_5234,N_2880,N_3251);
and U5235 (N_5235,N_3966,N_2513);
nor U5236 (N_5236,N_3251,N_2104);
xor U5237 (N_5237,N_2805,N_2136);
xnor U5238 (N_5238,N_2947,N_3390);
nor U5239 (N_5239,N_3885,N_3360);
and U5240 (N_5240,N_3287,N_2187);
and U5241 (N_5241,N_3955,N_2663);
or U5242 (N_5242,N_2677,N_2534);
or U5243 (N_5243,N_3748,N_3085);
and U5244 (N_5244,N_3458,N_3353);
nor U5245 (N_5245,N_3246,N_2796);
or U5246 (N_5246,N_3363,N_3350);
nand U5247 (N_5247,N_2549,N_2049);
nand U5248 (N_5248,N_2186,N_3292);
xor U5249 (N_5249,N_3971,N_2329);
nand U5250 (N_5250,N_3499,N_2415);
xnor U5251 (N_5251,N_3722,N_3144);
nor U5252 (N_5252,N_2724,N_2005);
or U5253 (N_5253,N_3337,N_3836);
and U5254 (N_5254,N_3323,N_2434);
or U5255 (N_5255,N_3584,N_3939);
nand U5256 (N_5256,N_2233,N_2758);
or U5257 (N_5257,N_2984,N_3312);
nor U5258 (N_5258,N_3159,N_2554);
nand U5259 (N_5259,N_2706,N_2558);
or U5260 (N_5260,N_3938,N_3700);
or U5261 (N_5261,N_2704,N_3303);
nor U5262 (N_5262,N_3301,N_3087);
nor U5263 (N_5263,N_3488,N_3915);
nor U5264 (N_5264,N_3225,N_3883);
nand U5265 (N_5265,N_3621,N_3672);
nor U5266 (N_5266,N_2205,N_3258);
nand U5267 (N_5267,N_3503,N_2664);
or U5268 (N_5268,N_3711,N_3779);
xnor U5269 (N_5269,N_3064,N_2696);
nand U5270 (N_5270,N_3022,N_2473);
and U5271 (N_5271,N_3105,N_2659);
xor U5272 (N_5272,N_3808,N_3431);
and U5273 (N_5273,N_2420,N_2161);
xor U5274 (N_5274,N_3503,N_3329);
nand U5275 (N_5275,N_2727,N_3950);
or U5276 (N_5276,N_3589,N_3955);
or U5277 (N_5277,N_2831,N_2274);
nor U5278 (N_5278,N_2224,N_2952);
nor U5279 (N_5279,N_2352,N_3065);
nand U5280 (N_5280,N_3310,N_2143);
and U5281 (N_5281,N_2036,N_3781);
and U5282 (N_5282,N_3537,N_2020);
xor U5283 (N_5283,N_2536,N_2463);
or U5284 (N_5284,N_3046,N_2372);
nand U5285 (N_5285,N_2768,N_2743);
nor U5286 (N_5286,N_2512,N_2950);
nor U5287 (N_5287,N_2922,N_3393);
nor U5288 (N_5288,N_3385,N_2359);
and U5289 (N_5289,N_2555,N_2449);
or U5290 (N_5290,N_3319,N_2855);
xnor U5291 (N_5291,N_3572,N_3223);
nor U5292 (N_5292,N_3425,N_2652);
or U5293 (N_5293,N_3623,N_3320);
and U5294 (N_5294,N_2252,N_3089);
or U5295 (N_5295,N_3738,N_2743);
xor U5296 (N_5296,N_2577,N_3164);
xnor U5297 (N_5297,N_2148,N_2538);
or U5298 (N_5298,N_3098,N_2907);
nand U5299 (N_5299,N_3385,N_3933);
nor U5300 (N_5300,N_3921,N_3945);
and U5301 (N_5301,N_3876,N_2223);
or U5302 (N_5302,N_3491,N_3231);
and U5303 (N_5303,N_3927,N_3899);
or U5304 (N_5304,N_3471,N_3903);
nand U5305 (N_5305,N_3570,N_2287);
and U5306 (N_5306,N_2544,N_3190);
xor U5307 (N_5307,N_3558,N_2945);
xnor U5308 (N_5308,N_2013,N_3751);
nand U5309 (N_5309,N_2501,N_2374);
and U5310 (N_5310,N_2730,N_2855);
nand U5311 (N_5311,N_2948,N_3251);
or U5312 (N_5312,N_2360,N_3330);
nor U5313 (N_5313,N_2909,N_3121);
or U5314 (N_5314,N_2204,N_3874);
nand U5315 (N_5315,N_2064,N_2817);
xor U5316 (N_5316,N_2159,N_2327);
xor U5317 (N_5317,N_3900,N_3012);
xor U5318 (N_5318,N_3890,N_3286);
or U5319 (N_5319,N_3783,N_2718);
and U5320 (N_5320,N_3610,N_2618);
nand U5321 (N_5321,N_2355,N_2043);
and U5322 (N_5322,N_2986,N_3022);
xor U5323 (N_5323,N_2546,N_3244);
nor U5324 (N_5324,N_3878,N_2206);
xor U5325 (N_5325,N_3529,N_3732);
or U5326 (N_5326,N_2810,N_2050);
or U5327 (N_5327,N_2246,N_2372);
nand U5328 (N_5328,N_3194,N_3606);
and U5329 (N_5329,N_3902,N_3653);
and U5330 (N_5330,N_2701,N_3408);
nand U5331 (N_5331,N_2478,N_2329);
nand U5332 (N_5332,N_3935,N_3795);
nand U5333 (N_5333,N_2762,N_2464);
nand U5334 (N_5334,N_3637,N_3706);
and U5335 (N_5335,N_3086,N_2566);
nor U5336 (N_5336,N_3326,N_3428);
xor U5337 (N_5337,N_3443,N_2210);
and U5338 (N_5338,N_2678,N_3415);
nand U5339 (N_5339,N_3865,N_2142);
and U5340 (N_5340,N_2762,N_3143);
nor U5341 (N_5341,N_3715,N_3798);
nor U5342 (N_5342,N_2465,N_2048);
and U5343 (N_5343,N_2779,N_3302);
and U5344 (N_5344,N_3318,N_2911);
nor U5345 (N_5345,N_3472,N_2155);
nand U5346 (N_5346,N_2562,N_3609);
nor U5347 (N_5347,N_2287,N_3607);
and U5348 (N_5348,N_2590,N_2448);
and U5349 (N_5349,N_2721,N_2689);
nor U5350 (N_5350,N_2755,N_2675);
xnor U5351 (N_5351,N_2720,N_3455);
xnor U5352 (N_5352,N_3862,N_3233);
and U5353 (N_5353,N_3657,N_3623);
nand U5354 (N_5354,N_3000,N_2612);
xnor U5355 (N_5355,N_3408,N_2208);
and U5356 (N_5356,N_2705,N_2961);
nor U5357 (N_5357,N_3014,N_2033);
nand U5358 (N_5358,N_3207,N_2344);
nor U5359 (N_5359,N_2446,N_2225);
nor U5360 (N_5360,N_3737,N_3488);
nand U5361 (N_5361,N_2491,N_3917);
or U5362 (N_5362,N_2049,N_2985);
nand U5363 (N_5363,N_2501,N_2012);
xor U5364 (N_5364,N_3329,N_2493);
and U5365 (N_5365,N_2884,N_3586);
and U5366 (N_5366,N_3227,N_3292);
xor U5367 (N_5367,N_2788,N_2179);
nor U5368 (N_5368,N_3192,N_2082);
nor U5369 (N_5369,N_3923,N_2283);
nand U5370 (N_5370,N_3968,N_2941);
nor U5371 (N_5371,N_2314,N_2039);
and U5372 (N_5372,N_2594,N_3710);
and U5373 (N_5373,N_3972,N_2760);
and U5374 (N_5374,N_3883,N_2117);
and U5375 (N_5375,N_3584,N_2899);
nand U5376 (N_5376,N_2220,N_3658);
and U5377 (N_5377,N_3514,N_3222);
and U5378 (N_5378,N_3278,N_2943);
xor U5379 (N_5379,N_2660,N_2940);
nand U5380 (N_5380,N_2468,N_3363);
or U5381 (N_5381,N_3333,N_2131);
and U5382 (N_5382,N_2871,N_3825);
nor U5383 (N_5383,N_2302,N_3252);
xnor U5384 (N_5384,N_2736,N_2581);
xor U5385 (N_5385,N_2956,N_2053);
xnor U5386 (N_5386,N_3524,N_3438);
nand U5387 (N_5387,N_3611,N_3273);
xnor U5388 (N_5388,N_3142,N_2959);
and U5389 (N_5389,N_2981,N_2311);
or U5390 (N_5390,N_3902,N_2583);
nor U5391 (N_5391,N_3579,N_3900);
nand U5392 (N_5392,N_2693,N_3998);
xnor U5393 (N_5393,N_3901,N_3639);
xnor U5394 (N_5394,N_2888,N_2465);
xnor U5395 (N_5395,N_2341,N_2816);
xnor U5396 (N_5396,N_2905,N_2792);
nand U5397 (N_5397,N_2824,N_2969);
and U5398 (N_5398,N_3425,N_3741);
xor U5399 (N_5399,N_2671,N_2760);
nor U5400 (N_5400,N_3617,N_3865);
xor U5401 (N_5401,N_3729,N_2986);
or U5402 (N_5402,N_2828,N_2534);
xnor U5403 (N_5403,N_2744,N_2039);
nor U5404 (N_5404,N_3781,N_3417);
nor U5405 (N_5405,N_3959,N_3484);
xnor U5406 (N_5406,N_2852,N_3788);
nand U5407 (N_5407,N_3131,N_2691);
or U5408 (N_5408,N_2150,N_2956);
and U5409 (N_5409,N_3065,N_3335);
nor U5410 (N_5410,N_2439,N_2928);
nor U5411 (N_5411,N_2377,N_2496);
or U5412 (N_5412,N_3755,N_3773);
xnor U5413 (N_5413,N_3713,N_3049);
and U5414 (N_5414,N_3661,N_2941);
nand U5415 (N_5415,N_2771,N_2164);
nor U5416 (N_5416,N_2548,N_2252);
nor U5417 (N_5417,N_2824,N_2025);
xnor U5418 (N_5418,N_3332,N_3068);
or U5419 (N_5419,N_3546,N_3519);
xor U5420 (N_5420,N_3772,N_2408);
and U5421 (N_5421,N_3913,N_2688);
xor U5422 (N_5422,N_2707,N_2202);
or U5423 (N_5423,N_3637,N_2345);
nor U5424 (N_5424,N_3668,N_2805);
nor U5425 (N_5425,N_2086,N_3968);
nand U5426 (N_5426,N_3898,N_2912);
and U5427 (N_5427,N_3619,N_3841);
nand U5428 (N_5428,N_3637,N_3634);
and U5429 (N_5429,N_3868,N_2199);
and U5430 (N_5430,N_2335,N_3063);
nor U5431 (N_5431,N_3102,N_2743);
nor U5432 (N_5432,N_3356,N_3463);
xnor U5433 (N_5433,N_2904,N_3110);
nor U5434 (N_5434,N_3369,N_3460);
nor U5435 (N_5435,N_2850,N_3080);
or U5436 (N_5436,N_3106,N_2494);
or U5437 (N_5437,N_2305,N_2340);
xor U5438 (N_5438,N_2946,N_2840);
nand U5439 (N_5439,N_2288,N_2557);
nand U5440 (N_5440,N_3464,N_3685);
and U5441 (N_5441,N_3667,N_2464);
nand U5442 (N_5442,N_2687,N_3606);
or U5443 (N_5443,N_3474,N_3348);
or U5444 (N_5444,N_3640,N_3539);
or U5445 (N_5445,N_3465,N_3295);
xor U5446 (N_5446,N_3070,N_3877);
or U5447 (N_5447,N_3883,N_2439);
and U5448 (N_5448,N_3838,N_2670);
xnor U5449 (N_5449,N_3758,N_3826);
or U5450 (N_5450,N_2532,N_2737);
xor U5451 (N_5451,N_3492,N_3791);
xnor U5452 (N_5452,N_3945,N_2177);
nand U5453 (N_5453,N_2532,N_3194);
nand U5454 (N_5454,N_2291,N_3558);
nand U5455 (N_5455,N_3356,N_2955);
or U5456 (N_5456,N_3365,N_2438);
nand U5457 (N_5457,N_2161,N_3547);
xnor U5458 (N_5458,N_2991,N_2545);
nor U5459 (N_5459,N_2595,N_3770);
nand U5460 (N_5460,N_2041,N_3625);
xor U5461 (N_5461,N_2720,N_2234);
xnor U5462 (N_5462,N_2367,N_2046);
or U5463 (N_5463,N_3617,N_3715);
or U5464 (N_5464,N_2618,N_3985);
nor U5465 (N_5465,N_3358,N_3291);
nor U5466 (N_5466,N_2164,N_3475);
or U5467 (N_5467,N_2506,N_3205);
and U5468 (N_5468,N_2647,N_2739);
and U5469 (N_5469,N_2404,N_2571);
and U5470 (N_5470,N_2067,N_2752);
xnor U5471 (N_5471,N_2538,N_2340);
nand U5472 (N_5472,N_2892,N_3816);
nor U5473 (N_5473,N_2869,N_2137);
nand U5474 (N_5474,N_3005,N_2423);
nor U5475 (N_5475,N_3519,N_3575);
xnor U5476 (N_5476,N_2837,N_3971);
nand U5477 (N_5477,N_3425,N_2183);
and U5478 (N_5478,N_2038,N_2355);
nand U5479 (N_5479,N_3680,N_3128);
nand U5480 (N_5480,N_3327,N_3465);
or U5481 (N_5481,N_3076,N_2835);
xnor U5482 (N_5482,N_2150,N_2426);
nand U5483 (N_5483,N_2700,N_3251);
nor U5484 (N_5484,N_2721,N_2908);
xnor U5485 (N_5485,N_3073,N_3278);
or U5486 (N_5486,N_3125,N_2848);
nor U5487 (N_5487,N_3128,N_2727);
or U5488 (N_5488,N_3988,N_3915);
nand U5489 (N_5489,N_3690,N_3769);
xor U5490 (N_5490,N_2744,N_2755);
or U5491 (N_5491,N_2529,N_3071);
nand U5492 (N_5492,N_2583,N_3660);
xor U5493 (N_5493,N_3254,N_3551);
and U5494 (N_5494,N_3096,N_2078);
nor U5495 (N_5495,N_2527,N_2332);
nand U5496 (N_5496,N_2072,N_2360);
xor U5497 (N_5497,N_3750,N_2415);
and U5498 (N_5498,N_3964,N_2566);
or U5499 (N_5499,N_2864,N_2726);
nand U5500 (N_5500,N_2540,N_2026);
nand U5501 (N_5501,N_3156,N_3007);
nand U5502 (N_5502,N_2178,N_3271);
or U5503 (N_5503,N_2684,N_3456);
xnor U5504 (N_5504,N_3614,N_2380);
or U5505 (N_5505,N_3640,N_3370);
and U5506 (N_5506,N_3531,N_2475);
or U5507 (N_5507,N_3329,N_3909);
nand U5508 (N_5508,N_2414,N_2412);
and U5509 (N_5509,N_2233,N_2868);
nor U5510 (N_5510,N_2694,N_2870);
xnor U5511 (N_5511,N_3328,N_3553);
nor U5512 (N_5512,N_3411,N_3452);
nor U5513 (N_5513,N_3222,N_2582);
and U5514 (N_5514,N_3525,N_3926);
xnor U5515 (N_5515,N_3342,N_3188);
or U5516 (N_5516,N_2929,N_2433);
and U5517 (N_5517,N_2880,N_2652);
nand U5518 (N_5518,N_3850,N_3728);
and U5519 (N_5519,N_3923,N_2038);
and U5520 (N_5520,N_2855,N_3743);
and U5521 (N_5521,N_3008,N_2005);
nand U5522 (N_5522,N_3365,N_2909);
xnor U5523 (N_5523,N_3920,N_2988);
or U5524 (N_5524,N_2890,N_2247);
nand U5525 (N_5525,N_2676,N_3725);
and U5526 (N_5526,N_2707,N_2863);
or U5527 (N_5527,N_2481,N_3065);
nor U5528 (N_5528,N_3495,N_2856);
or U5529 (N_5529,N_2145,N_2633);
or U5530 (N_5530,N_3292,N_2835);
nor U5531 (N_5531,N_2196,N_3942);
and U5532 (N_5532,N_2007,N_3635);
nand U5533 (N_5533,N_2864,N_3770);
and U5534 (N_5534,N_2961,N_3735);
and U5535 (N_5535,N_2357,N_2319);
nand U5536 (N_5536,N_3863,N_2239);
and U5537 (N_5537,N_3515,N_2052);
and U5538 (N_5538,N_3209,N_2860);
xor U5539 (N_5539,N_3230,N_3308);
and U5540 (N_5540,N_3745,N_2768);
and U5541 (N_5541,N_3660,N_2691);
xnor U5542 (N_5542,N_3663,N_3379);
or U5543 (N_5543,N_2474,N_2785);
nand U5544 (N_5544,N_3875,N_3261);
and U5545 (N_5545,N_3788,N_2626);
nand U5546 (N_5546,N_3166,N_2681);
xor U5547 (N_5547,N_2493,N_3246);
nand U5548 (N_5548,N_3756,N_2604);
xor U5549 (N_5549,N_2459,N_2858);
nor U5550 (N_5550,N_2686,N_3605);
nand U5551 (N_5551,N_3297,N_3425);
or U5552 (N_5552,N_2395,N_3181);
nand U5553 (N_5553,N_2175,N_3629);
nand U5554 (N_5554,N_3798,N_3291);
and U5555 (N_5555,N_3463,N_2307);
nand U5556 (N_5556,N_3516,N_2706);
and U5557 (N_5557,N_3842,N_3732);
xor U5558 (N_5558,N_2549,N_3886);
nor U5559 (N_5559,N_2706,N_2009);
xor U5560 (N_5560,N_2091,N_2718);
or U5561 (N_5561,N_3177,N_2141);
and U5562 (N_5562,N_2290,N_3129);
nor U5563 (N_5563,N_3432,N_2308);
xor U5564 (N_5564,N_2463,N_2124);
and U5565 (N_5565,N_2783,N_3963);
or U5566 (N_5566,N_3586,N_3835);
nor U5567 (N_5567,N_3619,N_2404);
or U5568 (N_5568,N_2246,N_3332);
xnor U5569 (N_5569,N_2889,N_3629);
xor U5570 (N_5570,N_2165,N_2377);
xnor U5571 (N_5571,N_2321,N_3455);
nor U5572 (N_5572,N_2141,N_2314);
or U5573 (N_5573,N_3226,N_3440);
nand U5574 (N_5574,N_2962,N_2748);
or U5575 (N_5575,N_3162,N_2249);
or U5576 (N_5576,N_3958,N_3591);
nand U5577 (N_5577,N_2370,N_3107);
nand U5578 (N_5578,N_3874,N_2510);
or U5579 (N_5579,N_2794,N_2106);
nor U5580 (N_5580,N_3011,N_3416);
xnor U5581 (N_5581,N_2790,N_3965);
nor U5582 (N_5582,N_2327,N_2825);
or U5583 (N_5583,N_2300,N_3004);
or U5584 (N_5584,N_3135,N_2726);
nor U5585 (N_5585,N_2625,N_2029);
and U5586 (N_5586,N_3164,N_2002);
or U5587 (N_5587,N_2274,N_2416);
nor U5588 (N_5588,N_2226,N_3135);
nor U5589 (N_5589,N_2436,N_3906);
nand U5590 (N_5590,N_3368,N_2924);
and U5591 (N_5591,N_2136,N_2457);
nand U5592 (N_5592,N_2395,N_2329);
and U5593 (N_5593,N_2919,N_3093);
xor U5594 (N_5594,N_3878,N_2078);
nand U5595 (N_5595,N_3595,N_2311);
nand U5596 (N_5596,N_2472,N_2581);
nor U5597 (N_5597,N_2001,N_3745);
or U5598 (N_5598,N_2979,N_3037);
and U5599 (N_5599,N_2069,N_3007);
xnor U5600 (N_5600,N_3861,N_3821);
nor U5601 (N_5601,N_2707,N_2213);
nand U5602 (N_5602,N_3192,N_2258);
or U5603 (N_5603,N_3490,N_2673);
or U5604 (N_5604,N_3458,N_3843);
nand U5605 (N_5605,N_2439,N_2297);
or U5606 (N_5606,N_3235,N_2676);
xnor U5607 (N_5607,N_2475,N_3378);
or U5608 (N_5608,N_2922,N_2889);
nand U5609 (N_5609,N_2616,N_3691);
nor U5610 (N_5610,N_2800,N_2929);
nand U5611 (N_5611,N_2824,N_3112);
nor U5612 (N_5612,N_2197,N_2045);
and U5613 (N_5613,N_3778,N_2744);
nor U5614 (N_5614,N_2964,N_2783);
or U5615 (N_5615,N_2966,N_2322);
nor U5616 (N_5616,N_2519,N_3495);
and U5617 (N_5617,N_2979,N_3156);
and U5618 (N_5618,N_3828,N_3814);
nor U5619 (N_5619,N_3763,N_2001);
or U5620 (N_5620,N_2994,N_3913);
nand U5621 (N_5621,N_2277,N_3098);
nor U5622 (N_5622,N_2962,N_2180);
nand U5623 (N_5623,N_3083,N_2689);
nor U5624 (N_5624,N_3135,N_3974);
or U5625 (N_5625,N_3164,N_2638);
or U5626 (N_5626,N_3301,N_2556);
nor U5627 (N_5627,N_3079,N_3673);
or U5628 (N_5628,N_2707,N_2110);
or U5629 (N_5629,N_3049,N_3320);
nand U5630 (N_5630,N_2268,N_3257);
nand U5631 (N_5631,N_2199,N_2273);
and U5632 (N_5632,N_3910,N_2083);
nand U5633 (N_5633,N_2118,N_2215);
xnor U5634 (N_5634,N_2982,N_3196);
or U5635 (N_5635,N_2983,N_3698);
nor U5636 (N_5636,N_2958,N_3750);
nor U5637 (N_5637,N_3632,N_3423);
and U5638 (N_5638,N_2527,N_2534);
and U5639 (N_5639,N_2884,N_3022);
nor U5640 (N_5640,N_2157,N_3752);
or U5641 (N_5641,N_2344,N_2623);
nor U5642 (N_5642,N_2148,N_3186);
and U5643 (N_5643,N_3562,N_3786);
or U5644 (N_5644,N_2100,N_2931);
or U5645 (N_5645,N_2193,N_2838);
or U5646 (N_5646,N_3377,N_2866);
and U5647 (N_5647,N_2628,N_3412);
nor U5648 (N_5648,N_3258,N_3523);
nor U5649 (N_5649,N_2652,N_2466);
nand U5650 (N_5650,N_2006,N_2076);
or U5651 (N_5651,N_3864,N_2189);
nor U5652 (N_5652,N_2087,N_2937);
nor U5653 (N_5653,N_2331,N_3988);
nand U5654 (N_5654,N_2789,N_3015);
nand U5655 (N_5655,N_2851,N_2108);
nor U5656 (N_5656,N_2985,N_3772);
nand U5657 (N_5657,N_3243,N_2846);
or U5658 (N_5658,N_2508,N_3930);
xnor U5659 (N_5659,N_3662,N_3032);
xnor U5660 (N_5660,N_2226,N_3941);
or U5661 (N_5661,N_2845,N_3912);
nand U5662 (N_5662,N_2542,N_2500);
nand U5663 (N_5663,N_3840,N_3612);
nor U5664 (N_5664,N_2440,N_2642);
xnor U5665 (N_5665,N_3397,N_2620);
xor U5666 (N_5666,N_3744,N_3388);
nand U5667 (N_5667,N_2236,N_2169);
xor U5668 (N_5668,N_3141,N_2201);
xor U5669 (N_5669,N_2800,N_2451);
nor U5670 (N_5670,N_3273,N_3430);
or U5671 (N_5671,N_3937,N_3976);
nand U5672 (N_5672,N_3555,N_2983);
nor U5673 (N_5673,N_3040,N_3944);
xor U5674 (N_5674,N_3809,N_2101);
or U5675 (N_5675,N_2494,N_2757);
and U5676 (N_5676,N_3810,N_3039);
or U5677 (N_5677,N_3731,N_2304);
xnor U5678 (N_5678,N_2566,N_2175);
nor U5679 (N_5679,N_2146,N_3939);
nor U5680 (N_5680,N_3086,N_2716);
or U5681 (N_5681,N_3467,N_3970);
or U5682 (N_5682,N_2028,N_3902);
nand U5683 (N_5683,N_3602,N_3777);
nor U5684 (N_5684,N_2845,N_2776);
and U5685 (N_5685,N_2224,N_2312);
nand U5686 (N_5686,N_2710,N_2834);
nand U5687 (N_5687,N_3550,N_2379);
xor U5688 (N_5688,N_3764,N_3597);
and U5689 (N_5689,N_2891,N_3954);
xor U5690 (N_5690,N_3471,N_3744);
or U5691 (N_5691,N_2227,N_3418);
or U5692 (N_5692,N_2228,N_3696);
xnor U5693 (N_5693,N_3038,N_2540);
nand U5694 (N_5694,N_3040,N_2378);
or U5695 (N_5695,N_3414,N_2470);
nand U5696 (N_5696,N_3188,N_3453);
nand U5697 (N_5697,N_2898,N_3523);
and U5698 (N_5698,N_2808,N_3724);
nand U5699 (N_5699,N_3424,N_3624);
or U5700 (N_5700,N_2258,N_2600);
xnor U5701 (N_5701,N_2204,N_3096);
nor U5702 (N_5702,N_2710,N_3229);
and U5703 (N_5703,N_2251,N_2198);
xnor U5704 (N_5704,N_3290,N_3177);
and U5705 (N_5705,N_2528,N_3873);
and U5706 (N_5706,N_3321,N_3276);
xnor U5707 (N_5707,N_2368,N_2582);
nand U5708 (N_5708,N_3050,N_2285);
nor U5709 (N_5709,N_2813,N_3130);
nand U5710 (N_5710,N_2706,N_2321);
xor U5711 (N_5711,N_2874,N_3882);
nand U5712 (N_5712,N_3781,N_3224);
and U5713 (N_5713,N_2354,N_3881);
xnor U5714 (N_5714,N_3895,N_3778);
nand U5715 (N_5715,N_2798,N_2084);
nand U5716 (N_5716,N_3200,N_2802);
nand U5717 (N_5717,N_2254,N_3978);
xor U5718 (N_5718,N_3986,N_2652);
nor U5719 (N_5719,N_3568,N_3106);
or U5720 (N_5720,N_3168,N_2672);
or U5721 (N_5721,N_3797,N_3288);
xor U5722 (N_5722,N_3997,N_3695);
nor U5723 (N_5723,N_2183,N_3842);
nand U5724 (N_5724,N_2631,N_3777);
nor U5725 (N_5725,N_3669,N_3089);
or U5726 (N_5726,N_3021,N_3458);
nand U5727 (N_5727,N_2259,N_2709);
nor U5728 (N_5728,N_2502,N_2530);
nand U5729 (N_5729,N_3029,N_2741);
nand U5730 (N_5730,N_2977,N_3311);
or U5731 (N_5731,N_2205,N_3986);
or U5732 (N_5732,N_3237,N_2015);
and U5733 (N_5733,N_2668,N_2758);
xnor U5734 (N_5734,N_2726,N_3840);
and U5735 (N_5735,N_3535,N_3877);
or U5736 (N_5736,N_3816,N_3730);
or U5737 (N_5737,N_3811,N_3650);
nand U5738 (N_5738,N_3042,N_3867);
or U5739 (N_5739,N_3572,N_3690);
and U5740 (N_5740,N_3929,N_3283);
xnor U5741 (N_5741,N_3270,N_3135);
or U5742 (N_5742,N_2755,N_2992);
nor U5743 (N_5743,N_3954,N_3600);
nand U5744 (N_5744,N_2644,N_2007);
and U5745 (N_5745,N_3740,N_3633);
xor U5746 (N_5746,N_2954,N_2031);
nor U5747 (N_5747,N_2828,N_2575);
nor U5748 (N_5748,N_3625,N_3121);
nand U5749 (N_5749,N_2462,N_2482);
xnor U5750 (N_5750,N_2440,N_3083);
nand U5751 (N_5751,N_3759,N_3927);
and U5752 (N_5752,N_2337,N_2959);
xnor U5753 (N_5753,N_2788,N_3664);
nor U5754 (N_5754,N_3326,N_2992);
or U5755 (N_5755,N_2401,N_3598);
nor U5756 (N_5756,N_2603,N_3036);
or U5757 (N_5757,N_2233,N_3590);
and U5758 (N_5758,N_3308,N_3634);
or U5759 (N_5759,N_2739,N_2783);
or U5760 (N_5760,N_2557,N_2193);
or U5761 (N_5761,N_2186,N_2165);
xor U5762 (N_5762,N_2120,N_2961);
xnor U5763 (N_5763,N_2068,N_2960);
and U5764 (N_5764,N_2630,N_3014);
nand U5765 (N_5765,N_2773,N_3384);
and U5766 (N_5766,N_2073,N_2845);
or U5767 (N_5767,N_3152,N_2149);
xor U5768 (N_5768,N_2408,N_2754);
and U5769 (N_5769,N_2079,N_3711);
xor U5770 (N_5770,N_2923,N_3297);
xor U5771 (N_5771,N_2757,N_2722);
xnor U5772 (N_5772,N_2381,N_3889);
and U5773 (N_5773,N_3997,N_3798);
and U5774 (N_5774,N_2815,N_2512);
nor U5775 (N_5775,N_3710,N_3276);
and U5776 (N_5776,N_3603,N_2228);
or U5777 (N_5777,N_2809,N_3050);
and U5778 (N_5778,N_2200,N_2971);
or U5779 (N_5779,N_2879,N_3959);
nor U5780 (N_5780,N_2869,N_3815);
xnor U5781 (N_5781,N_2150,N_2616);
nor U5782 (N_5782,N_3407,N_3930);
and U5783 (N_5783,N_2448,N_2035);
or U5784 (N_5784,N_3630,N_2725);
nand U5785 (N_5785,N_3436,N_3931);
xor U5786 (N_5786,N_2077,N_3049);
xor U5787 (N_5787,N_3996,N_3222);
xnor U5788 (N_5788,N_3734,N_3949);
nand U5789 (N_5789,N_3103,N_3711);
or U5790 (N_5790,N_3227,N_3651);
xor U5791 (N_5791,N_2014,N_2259);
or U5792 (N_5792,N_3703,N_3163);
xor U5793 (N_5793,N_3498,N_3522);
xnor U5794 (N_5794,N_3077,N_3701);
nor U5795 (N_5795,N_2535,N_3209);
or U5796 (N_5796,N_3046,N_2636);
or U5797 (N_5797,N_2026,N_3683);
and U5798 (N_5798,N_3016,N_2349);
or U5799 (N_5799,N_2044,N_3612);
nand U5800 (N_5800,N_3270,N_3115);
nand U5801 (N_5801,N_2721,N_2643);
and U5802 (N_5802,N_3635,N_3760);
nand U5803 (N_5803,N_2389,N_2100);
nand U5804 (N_5804,N_3504,N_3045);
or U5805 (N_5805,N_3977,N_3613);
nor U5806 (N_5806,N_3933,N_3166);
or U5807 (N_5807,N_2556,N_2363);
xnor U5808 (N_5808,N_2801,N_3776);
and U5809 (N_5809,N_3328,N_3047);
or U5810 (N_5810,N_3238,N_3626);
and U5811 (N_5811,N_2869,N_3522);
nand U5812 (N_5812,N_3332,N_2612);
or U5813 (N_5813,N_2572,N_3610);
nand U5814 (N_5814,N_3623,N_2182);
or U5815 (N_5815,N_3537,N_3991);
nor U5816 (N_5816,N_2530,N_3491);
and U5817 (N_5817,N_3741,N_3325);
nor U5818 (N_5818,N_3171,N_3874);
and U5819 (N_5819,N_2192,N_3425);
or U5820 (N_5820,N_3269,N_3975);
nand U5821 (N_5821,N_3227,N_2530);
nor U5822 (N_5822,N_3613,N_2104);
nand U5823 (N_5823,N_2626,N_2277);
and U5824 (N_5824,N_3061,N_3733);
nand U5825 (N_5825,N_2249,N_2164);
and U5826 (N_5826,N_2866,N_3920);
nand U5827 (N_5827,N_3976,N_2208);
and U5828 (N_5828,N_3290,N_3041);
nor U5829 (N_5829,N_2629,N_2007);
nor U5830 (N_5830,N_3752,N_2237);
or U5831 (N_5831,N_2577,N_2442);
nand U5832 (N_5832,N_3556,N_2896);
and U5833 (N_5833,N_3386,N_3703);
nor U5834 (N_5834,N_3048,N_2102);
and U5835 (N_5835,N_3885,N_2287);
xor U5836 (N_5836,N_2464,N_2808);
and U5837 (N_5837,N_2726,N_3065);
and U5838 (N_5838,N_3384,N_2460);
xor U5839 (N_5839,N_2894,N_3114);
and U5840 (N_5840,N_3456,N_3600);
nor U5841 (N_5841,N_3879,N_3757);
xor U5842 (N_5842,N_2759,N_2225);
or U5843 (N_5843,N_3488,N_2286);
nand U5844 (N_5844,N_2489,N_2824);
nand U5845 (N_5845,N_2458,N_3504);
nor U5846 (N_5846,N_3283,N_3215);
and U5847 (N_5847,N_2212,N_2308);
nand U5848 (N_5848,N_3865,N_2480);
nor U5849 (N_5849,N_3571,N_3416);
nand U5850 (N_5850,N_3923,N_3666);
nand U5851 (N_5851,N_3307,N_2581);
or U5852 (N_5852,N_2434,N_2339);
nor U5853 (N_5853,N_3689,N_2010);
nand U5854 (N_5854,N_3209,N_3349);
xor U5855 (N_5855,N_3732,N_2115);
or U5856 (N_5856,N_3087,N_3813);
nand U5857 (N_5857,N_3208,N_2601);
and U5858 (N_5858,N_2784,N_3377);
nand U5859 (N_5859,N_3547,N_3080);
nor U5860 (N_5860,N_2095,N_2002);
nand U5861 (N_5861,N_2930,N_2733);
nor U5862 (N_5862,N_3091,N_2504);
and U5863 (N_5863,N_3261,N_3673);
and U5864 (N_5864,N_3288,N_3392);
nand U5865 (N_5865,N_3970,N_2208);
and U5866 (N_5866,N_2468,N_3833);
xor U5867 (N_5867,N_3486,N_2278);
xnor U5868 (N_5868,N_2874,N_3009);
nand U5869 (N_5869,N_2047,N_2365);
nor U5870 (N_5870,N_3686,N_2494);
xor U5871 (N_5871,N_3554,N_3066);
nand U5872 (N_5872,N_3767,N_2509);
and U5873 (N_5873,N_2719,N_3028);
xor U5874 (N_5874,N_2928,N_3918);
nor U5875 (N_5875,N_2265,N_2986);
and U5876 (N_5876,N_2004,N_2269);
and U5877 (N_5877,N_3342,N_2549);
or U5878 (N_5878,N_2657,N_3837);
and U5879 (N_5879,N_2010,N_3096);
nand U5880 (N_5880,N_2514,N_3567);
xnor U5881 (N_5881,N_2273,N_2309);
and U5882 (N_5882,N_2828,N_3852);
and U5883 (N_5883,N_3185,N_2607);
and U5884 (N_5884,N_2166,N_2211);
or U5885 (N_5885,N_2198,N_2591);
or U5886 (N_5886,N_2767,N_2896);
nor U5887 (N_5887,N_2575,N_3515);
nor U5888 (N_5888,N_3734,N_3629);
or U5889 (N_5889,N_3447,N_2325);
nor U5890 (N_5890,N_3533,N_3391);
or U5891 (N_5891,N_2398,N_2758);
xor U5892 (N_5892,N_2207,N_3531);
nor U5893 (N_5893,N_3475,N_2377);
or U5894 (N_5894,N_2424,N_2285);
nor U5895 (N_5895,N_3045,N_3836);
or U5896 (N_5896,N_2914,N_2888);
nand U5897 (N_5897,N_2174,N_2680);
xor U5898 (N_5898,N_2916,N_3033);
xor U5899 (N_5899,N_3220,N_2073);
nor U5900 (N_5900,N_2944,N_3974);
nand U5901 (N_5901,N_3068,N_2849);
nand U5902 (N_5902,N_3443,N_3163);
or U5903 (N_5903,N_2894,N_2887);
nand U5904 (N_5904,N_3372,N_3759);
and U5905 (N_5905,N_2104,N_3135);
nor U5906 (N_5906,N_3177,N_2541);
xnor U5907 (N_5907,N_3506,N_2799);
or U5908 (N_5908,N_2608,N_3635);
nor U5909 (N_5909,N_2091,N_3505);
xnor U5910 (N_5910,N_3867,N_3361);
and U5911 (N_5911,N_2352,N_3223);
or U5912 (N_5912,N_2101,N_3690);
or U5913 (N_5913,N_3380,N_2350);
nand U5914 (N_5914,N_3331,N_2073);
nor U5915 (N_5915,N_3176,N_3159);
nor U5916 (N_5916,N_2908,N_2755);
or U5917 (N_5917,N_2518,N_3324);
or U5918 (N_5918,N_3659,N_3618);
xnor U5919 (N_5919,N_3641,N_3837);
or U5920 (N_5920,N_2794,N_3577);
nand U5921 (N_5921,N_2214,N_3450);
xnor U5922 (N_5922,N_3019,N_2511);
xor U5923 (N_5923,N_2428,N_2605);
and U5924 (N_5924,N_2561,N_3169);
or U5925 (N_5925,N_2380,N_2026);
nand U5926 (N_5926,N_3816,N_2006);
xor U5927 (N_5927,N_2697,N_3036);
nor U5928 (N_5928,N_3124,N_3639);
or U5929 (N_5929,N_3193,N_2866);
nand U5930 (N_5930,N_2853,N_3115);
nand U5931 (N_5931,N_2706,N_2772);
and U5932 (N_5932,N_2486,N_3988);
or U5933 (N_5933,N_3235,N_3911);
xnor U5934 (N_5934,N_3772,N_3617);
or U5935 (N_5935,N_3853,N_2909);
nand U5936 (N_5936,N_2321,N_3155);
xor U5937 (N_5937,N_3905,N_2699);
and U5938 (N_5938,N_2688,N_3077);
or U5939 (N_5939,N_2709,N_3288);
xor U5940 (N_5940,N_2479,N_2877);
xor U5941 (N_5941,N_3319,N_2782);
xor U5942 (N_5942,N_2939,N_3404);
nand U5943 (N_5943,N_2950,N_2452);
xor U5944 (N_5944,N_3462,N_3558);
nor U5945 (N_5945,N_3779,N_2409);
nor U5946 (N_5946,N_2453,N_2695);
and U5947 (N_5947,N_3019,N_2248);
nor U5948 (N_5948,N_2217,N_3291);
or U5949 (N_5949,N_3108,N_2626);
nor U5950 (N_5950,N_3598,N_2735);
or U5951 (N_5951,N_2082,N_2472);
and U5952 (N_5952,N_3274,N_2721);
and U5953 (N_5953,N_2377,N_3718);
or U5954 (N_5954,N_2424,N_3797);
and U5955 (N_5955,N_3453,N_2830);
xor U5956 (N_5956,N_3066,N_3308);
nor U5957 (N_5957,N_2994,N_3648);
and U5958 (N_5958,N_3227,N_2379);
or U5959 (N_5959,N_2398,N_2957);
xnor U5960 (N_5960,N_3713,N_3390);
xnor U5961 (N_5961,N_2295,N_2524);
xnor U5962 (N_5962,N_2131,N_2119);
nand U5963 (N_5963,N_3547,N_2128);
nand U5964 (N_5964,N_3302,N_3990);
and U5965 (N_5965,N_3035,N_2251);
nand U5966 (N_5966,N_2700,N_2727);
nand U5967 (N_5967,N_2095,N_2509);
nand U5968 (N_5968,N_2469,N_3426);
or U5969 (N_5969,N_2497,N_3621);
xnor U5970 (N_5970,N_2585,N_2793);
and U5971 (N_5971,N_2696,N_2684);
and U5972 (N_5972,N_3141,N_3508);
or U5973 (N_5973,N_3283,N_3450);
and U5974 (N_5974,N_3023,N_2156);
nand U5975 (N_5975,N_3928,N_2350);
xnor U5976 (N_5976,N_2409,N_3369);
nor U5977 (N_5977,N_3917,N_2057);
nand U5978 (N_5978,N_3862,N_2947);
nand U5979 (N_5979,N_3724,N_2648);
nor U5980 (N_5980,N_3857,N_2475);
xor U5981 (N_5981,N_2917,N_2363);
nand U5982 (N_5982,N_3027,N_2858);
xor U5983 (N_5983,N_2956,N_2557);
nor U5984 (N_5984,N_2606,N_2604);
or U5985 (N_5985,N_3015,N_2451);
and U5986 (N_5986,N_3880,N_3765);
and U5987 (N_5987,N_3344,N_3799);
nor U5988 (N_5988,N_3250,N_3787);
nand U5989 (N_5989,N_2797,N_3296);
or U5990 (N_5990,N_3549,N_2388);
xor U5991 (N_5991,N_3716,N_3060);
nor U5992 (N_5992,N_3190,N_2246);
and U5993 (N_5993,N_2212,N_3692);
nand U5994 (N_5994,N_3055,N_3589);
nand U5995 (N_5995,N_2460,N_2463);
nand U5996 (N_5996,N_2027,N_2200);
nand U5997 (N_5997,N_2930,N_2535);
xnor U5998 (N_5998,N_3320,N_3016);
or U5999 (N_5999,N_2277,N_3416);
nand U6000 (N_6000,N_4516,N_4777);
and U6001 (N_6001,N_5442,N_4255);
nor U6002 (N_6002,N_5695,N_5705);
xor U6003 (N_6003,N_4410,N_4452);
nor U6004 (N_6004,N_5875,N_4674);
xor U6005 (N_6005,N_4395,N_4078);
and U6006 (N_6006,N_4281,N_4604);
nor U6007 (N_6007,N_4213,N_4322);
xnor U6008 (N_6008,N_4787,N_5037);
and U6009 (N_6009,N_4494,N_5313);
xnor U6010 (N_6010,N_4485,N_5608);
nor U6011 (N_6011,N_5527,N_4127);
or U6012 (N_6012,N_5579,N_5847);
xor U6013 (N_6013,N_4178,N_4130);
nor U6014 (N_6014,N_4907,N_5147);
or U6015 (N_6015,N_5176,N_4039);
nor U6016 (N_6016,N_4967,N_5321);
nand U6017 (N_6017,N_5134,N_5757);
nor U6018 (N_6018,N_5363,N_5961);
nand U6019 (N_6019,N_5184,N_5574);
and U6020 (N_6020,N_4641,N_4229);
nand U6021 (N_6021,N_4900,N_5106);
xor U6022 (N_6022,N_5137,N_5666);
or U6023 (N_6023,N_4275,N_4580);
nor U6024 (N_6024,N_4404,N_4341);
nand U6025 (N_6025,N_4160,N_4131);
nand U6026 (N_6026,N_4665,N_4508);
nor U6027 (N_6027,N_5067,N_4473);
or U6028 (N_6028,N_5979,N_4757);
or U6029 (N_6029,N_4937,N_4203);
or U6030 (N_6030,N_4511,N_4881);
xnor U6031 (N_6031,N_5436,N_4501);
nand U6032 (N_6032,N_4152,N_5471);
nor U6033 (N_6033,N_4792,N_5131);
nand U6034 (N_6034,N_5936,N_5975);
nor U6035 (N_6035,N_4183,N_5978);
and U6036 (N_6036,N_4686,N_5098);
xnor U6037 (N_6037,N_5942,N_4558);
and U6038 (N_6038,N_4133,N_4345);
and U6039 (N_6039,N_5309,N_4679);
and U6040 (N_6040,N_5824,N_4601);
nor U6041 (N_6041,N_5553,N_4675);
and U6042 (N_6042,N_5329,N_5731);
and U6043 (N_6043,N_4128,N_4776);
nor U6044 (N_6044,N_4938,N_4918);
nand U6045 (N_6045,N_4902,N_5125);
nand U6046 (N_6046,N_4840,N_5908);
nor U6047 (N_6047,N_5514,N_5160);
nand U6048 (N_6048,N_4228,N_5153);
nor U6049 (N_6049,N_4234,N_5849);
xnor U6050 (N_6050,N_5177,N_4474);
xor U6051 (N_6051,N_5141,N_4442);
xor U6052 (N_6052,N_4236,N_5361);
or U6053 (N_6053,N_5499,N_4979);
xnor U6054 (N_6054,N_5158,N_5439);
nor U6055 (N_6055,N_5539,N_5909);
xor U6056 (N_6056,N_4858,N_5054);
nor U6057 (N_6057,N_4155,N_5333);
nand U6058 (N_6058,N_5733,N_4172);
and U6059 (N_6059,N_5492,N_5627);
nand U6060 (N_6060,N_5836,N_5586);
and U6061 (N_6061,N_4744,N_5216);
and U6062 (N_6062,N_5868,N_5116);
or U6063 (N_6063,N_4374,N_4481);
nand U6064 (N_6064,N_5244,N_5905);
and U6065 (N_6065,N_5466,N_5315);
or U6066 (N_6066,N_5193,N_4138);
nand U6067 (N_6067,N_5181,N_4600);
nor U6068 (N_6068,N_4871,N_4930);
xnor U6069 (N_6069,N_5569,N_5251);
nand U6070 (N_6070,N_5648,N_4908);
nor U6071 (N_6071,N_4661,N_5538);
xor U6072 (N_6072,N_5959,N_4096);
nand U6073 (N_6073,N_5250,N_5448);
nor U6074 (N_6074,N_4008,N_4310);
xnor U6075 (N_6075,N_5214,N_4115);
xnor U6076 (N_6076,N_4505,N_5982);
nand U6077 (N_6077,N_4239,N_4118);
or U6078 (N_6078,N_4567,N_4295);
nand U6079 (N_6079,N_5587,N_5521);
nor U6080 (N_6080,N_4610,N_4763);
nor U6081 (N_6081,N_4478,N_5071);
xor U6082 (N_6082,N_4707,N_4126);
xor U6083 (N_6083,N_4996,N_5736);
or U6084 (N_6084,N_4443,N_4260);
xnor U6085 (N_6085,N_4681,N_5743);
nor U6086 (N_6086,N_4687,N_5928);
xor U6087 (N_6087,N_4323,N_5678);
xnor U6088 (N_6088,N_4286,N_5612);
and U6089 (N_6089,N_4193,N_5740);
nand U6090 (N_6090,N_5676,N_4755);
nand U6091 (N_6091,N_4873,N_5179);
and U6092 (N_6092,N_4640,N_4406);
and U6093 (N_6093,N_4054,N_5080);
nand U6094 (N_6094,N_5613,N_4314);
and U6095 (N_6095,N_5159,N_4164);
nor U6096 (N_6096,N_4643,N_5667);
and U6097 (N_6097,N_4841,N_5960);
nor U6098 (N_6098,N_4882,N_4734);
nor U6099 (N_6099,N_4664,N_5324);
and U6100 (N_6100,N_4036,N_5095);
nor U6101 (N_6101,N_5291,N_5500);
or U6102 (N_6102,N_4090,N_4555);
nor U6103 (N_6103,N_5215,N_4232);
nand U6104 (N_6104,N_4968,N_4267);
nor U6105 (N_6105,N_5674,N_4951);
and U6106 (N_6106,N_4997,N_5078);
nand U6107 (N_6107,N_4257,N_5248);
and U6108 (N_6108,N_5772,N_5008);
and U6109 (N_6109,N_5649,N_5175);
nand U6110 (N_6110,N_4954,N_5461);
xnor U6111 (N_6111,N_4433,N_4527);
nor U6112 (N_6112,N_5422,N_5338);
nand U6113 (N_6113,N_4392,N_4446);
or U6114 (N_6114,N_4905,N_5884);
and U6115 (N_6115,N_4585,N_5317);
nand U6116 (N_6116,N_5891,N_4344);
or U6117 (N_6117,N_5292,N_5433);
or U6118 (N_6118,N_5644,N_4283);
nor U6119 (N_6119,N_4480,N_5014);
or U6120 (N_6120,N_4593,N_4955);
nand U6121 (N_6121,N_4885,N_4596);
xor U6122 (N_6122,N_4020,N_5617);
nor U6123 (N_6123,N_4572,N_4316);
or U6124 (N_6124,N_5033,N_5257);
xnor U6125 (N_6125,N_5459,N_4284);
xnor U6126 (N_6126,N_5778,N_4093);
nor U6127 (N_6127,N_5127,N_5092);
and U6128 (N_6128,N_5786,N_5922);
nor U6129 (N_6129,N_5630,N_5993);
and U6130 (N_6130,N_5104,N_5166);
or U6131 (N_6131,N_5918,N_4876);
nor U6132 (N_6132,N_5373,N_4301);
xnor U6133 (N_6133,N_4676,N_4758);
nand U6134 (N_6134,N_4923,N_4924);
nand U6135 (N_6135,N_4919,N_4754);
nand U6136 (N_6136,N_4101,N_5332);
nor U6137 (N_6137,N_5618,N_5969);
and U6138 (N_6138,N_4415,N_4067);
xnor U6139 (N_6139,N_5706,N_4429);
nor U6140 (N_6140,N_5407,N_4496);
and U6141 (N_6141,N_5105,N_4856);
and U6142 (N_6142,N_5227,N_4500);
nand U6143 (N_6143,N_5755,N_4512);
or U6144 (N_6144,N_5045,N_4804);
nor U6145 (N_6145,N_4028,N_5645);
xor U6146 (N_6146,N_5984,N_4079);
xnor U6147 (N_6147,N_4171,N_4177);
nor U6148 (N_6148,N_4689,N_5531);
and U6149 (N_6149,N_4261,N_4911);
and U6150 (N_6150,N_4723,N_5896);
and U6151 (N_6151,N_5821,N_4196);
and U6152 (N_6152,N_4844,N_4439);
or U6153 (N_6153,N_5737,N_4308);
xor U6154 (N_6154,N_5111,N_5224);
and U6155 (N_6155,N_4035,N_4716);
and U6156 (N_6156,N_5591,N_4351);
nand U6157 (N_6157,N_4386,N_5314);
xor U6158 (N_6158,N_5920,N_4578);
or U6159 (N_6159,N_4337,N_4595);
and U6160 (N_6160,N_4520,N_5869);
and U6161 (N_6161,N_5885,N_4484);
and U6162 (N_6162,N_5119,N_4735);
and U6163 (N_6163,N_4813,N_5677);
nand U6164 (N_6164,N_5915,N_4546);
or U6165 (N_6165,N_4801,N_5351);
and U6166 (N_6166,N_5528,N_4065);
nor U6167 (N_6167,N_4153,N_4498);
xnor U6168 (N_6168,N_4461,N_4909);
xor U6169 (N_6169,N_5290,N_5218);
nand U6170 (N_6170,N_4389,N_5983);
nand U6171 (N_6171,N_4615,N_5861);
and U6172 (N_6172,N_4960,N_5203);
xnor U6173 (N_6173,N_5780,N_4605);
nand U6174 (N_6174,N_5062,N_5398);
nand U6175 (N_6175,N_5404,N_5515);
or U6176 (N_6176,N_5495,N_4852);
nor U6177 (N_6177,N_5256,N_5540);
xnor U6178 (N_6178,N_4248,N_5082);
nor U6179 (N_6179,N_5242,N_5563);
and U6180 (N_6180,N_4680,N_5653);
nor U6181 (N_6181,N_5811,N_4708);
xnor U6182 (N_6182,N_4878,N_4764);
or U6183 (N_6183,N_5712,N_5164);
nor U6184 (N_6184,N_5491,N_5651);
nor U6185 (N_6185,N_4904,N_5451);
nor U6186 (N_6186,N_4659,N_4857);
nor U6187 (N_6187,N_4850,N_5118);
and U6188 (N_6188,N_4989,N_5659);
and U6189 (N_6189,N_5031,N_5526);
nor U6190 (N_6190,N_4948,N_5505);
nand U6191 (N_6191,N_4252,N_4538);
or U6192 (N_6192,N_4746,N_4145);
xnor U6193 (N_6193,N_5124,N_4751);
nand U6194 (N_6194,N_5409,N_5717);
or U6195 (N_6195,N_4618,N_4025);
and U6196 (N_6196,N_4574,N_4202);
nand U6197 (N_6197,N_5340,N_4427);
xor U6198 (N_6198,N_5243,N_4306);
and U6199 (N_6199,N_5862,N_5254);
and U6200 (N_6200,N_5679,N_4957);
or U6201 (N_6201,N_4720,N_5749);
xnor U6202 (N_6202,N_5196,N_4271);
nand U6203 (N_6203,N_4545,N_5343);
xnor U6204 (N_6204,N_5319,N_5155);
and U6205 (N_6205,N_4727,N_5728);
nand U6206 (N_6206,N_5482,N_5610);
nor U6207 (N_6207,N_4666,N_4941);
xnor U6208 (N_6208,N_5446,N_5415);
and U6209 (N_6209,N_4276,N_5994);
xnor U6210 (N_6210,N_5413,N_5932);
or U6211 (N_6211,N_5434,N_4944);
nor U6212 (N_6212,N_4129,N_4667);
nand U6213 (N_6213,N_5396,N_4015);
xor U6214 (N_6214,N_4430,N_5680);
nor U6215 (N_6215,N_5472,N_4011);
nor U6216 (N_6216,N_4471,N_5464);
and U6217 (N_6217,N_4087,N_5819);
or U6218 (N_6218,N_4220,N_5543);
xnor U6219 (N_6219,N_5814,N_5370);
nor U6220 (N_6220,N_5567,N_5596);
nor U6221 (N_6221,N_4952,N_5083);
or U6222 (N_6222,N_5665,N_4898);
xor U6223 (N_6223,N_4318,N_5637);
xnor U6224 (N_6224,N_4273,N_5304);
or U6225 (N_6225,N_5704,N_4633);
and U6226 (N_6226,N_4534,N_5641);
nand U6227 (N_6227,N_5399,N_4245);
nand U6228 (N_6228,N_4612,N_4401);
or U6229 (N_6229,N_4377,N_4802);
nand U6230 (N_6230,N_5890,N_5688);
or U6231 (N_6231,N_5592,N_5110);
or U6232 (N_6232,N_4737,N_5508);
xnor U6233 (N_6233,N_5601,N_5206);
nand U6234 (N_6234,N_5519,N_4431);
nor U6235 (N_6235,N_5072,N_4269);
and U6236 (N_6236,N_4851,N_4265);
xnor U6237 (N_6237,N_5352,N_4791);
xor U6238 (N_6238,N_4311,N_5209);
nand U6239 (N_6239,N_4730,N_4719);
or U6240 (N_6240,N_5079,N_4290);
or U6241 (N_6241,N_4515,N_4003);
xnor U6242 (N_6242,N_5555,N_4411);
xor U6243 (N_6243,N_5701,N_5981);
nand U6244 (N_6244,N_5086,N_4901);
nor U6245 (N_6245,N_4903,N_4820);
or U6246 (N_6246,N_4060,N_5792);
and U6247 (N_6247,N_4068,N_5170);
or U6248 (N_6248,N_5096,N_4992);
nor U6249 (N_6249,N_5832,N_4073);
or U6250 (N_6250,N_5943,N_5359);
xor U6251 (N_6251,N_5146,N_5270);
nand U6252 (N_6252,N_4910,N_4075);
nand U6253 (N_6253,N_4663,N_4187);
or U6254 (N_6254,N_5228,N_5020);
nor U6255 (N_6255,N_4379,N_4916);
xor U6256 (N_6256,N_5582,N_5202);
or U6257 (N_6257,N_5498,N_5428);
nor U6258 (N_6258,N_4999,N_5801);
or U6259 (N_6259,N_5190,N_5962);
and U6260 (N_6260,N_4143,N_5052);
xnor U6261 (N_6261,N_5523,N_5661);
nor U6262 (N_6262,N_5001,N_5235);
or U6263 (N_6263,N_5377,N_5600);
or U6264 (N_6264,N_5000,N_4365);
or U6265 (N_6265,N_5326,N_4636);
nor U6266 (N_6266,N_4782,N_4083);
or U6267 (N_6267,N_5197,N_5026);
xor U6268 (N_6268,N_5604,N_4483);
nand U6269 (N_6269,N_5093,N_5097);
xor U6270 (N_6270,N_4583,N_4420);
or U6271 (N_6271,N_5631,N_4082);
xnor U6272 (N_6272,N_4051,N_4625);
nand U6273 (N_6273,N_4049,N_5076);
nor U6274 (N_6274,N_5199,N_4147);
xnor U6275 (N_6275,N_5501,N_4210);
xor U6276 (N_6276,N_4581,N_4548);
nor U6277 (N_6277,N_4722,N_5522);
or U6278 (N_6278,N_5360,N_4590);
or U6279 (N_6279,N_5041,N_4437);
nor U6280 (N_6280,N_4380,N_4463);
or U6281 (N_6281,N_4653,N_5264);
nand U6282 (N_6282,N_4435,N_4588);
or U6283 (N_6283,N_4331,N_4259);
nor U6284 (N_6284,N_4603,N_5525);
or U6285 (N_6285,N_4778,N_5132);
and U6286 (N_6286,N_5576,N_4945);
xnor U6287 (N_6287,N_4211,N_5873);
xnor U6288 (N_6288,N_5504,N_4726);
and U6289 (N_6289,N_4022,N_4409);
nor U6290 (N_6290,N_4497,N_5350);
nand U6291 (N_6291,N_4414,N_4859);
or U6292 (N_6292,N_5136,N_5622);
xnor U6293 (N_6293,N_4825,N_4630);
nor U6294 (N_6294,N_5957,N_4785);
xnor U6295 (N_6295,N_5476,N_5513);
nor U6296 (N_6296,N_5729,N_4611);
nor U6297 (N_6297,N_5887,N_5584);
xor U6298 (N_6298,N_5298,N_4589);
nand U6299 (N_6299,N_5063,N_5019);
nand U6300 (N_6300,N_5931,N_4398);
or U6301 (N_6301,N_4030,N_4305);
and U6302 (N_6302,N_4510,N_4010);
nor U6303 (N_6303,N_4888,N_4956);
xnor U6304 (N_6304,N_5178,N_5796);
nand U6305 (N_6305,N_4094,N_4298);
xnor U6306 (N_6306,N_4334,N_4080);
nor U6307 (N_6307,N_5417,N_5198);
nand U6308 (N_6308,N_5296,N_5262);
nor U6309 (N_6309,N_5061,N_4350);
or U6310 (N_6310,N_5906,N_5099);
and U6311 (N_6311,N_5968,N_5839);
nor U6312 (N_6312,N_4346,N_4218);
nand U6313 (N_6313,N_4436,N_5646);
nand U6314 (N_6314,N_4691,N_4521);
nor U6315 (N_6315,N_4262,N_4912);
xnor U6316 (N_6316,N_5963,N_5907);
and U6317 (N_6317,N_4491,N_4274);
or U6318 (N_6318,N_5550,N_4642);
xnor U6319 (N_6319,N_4227,N_4826);
xor U6320 (N_6320,N_5595,N_4032);
nand U6321 (N_6321,N_5140,N_5858);
xnor U6322 (N_6322,N_4116,N_4326);
nand U6323 (N_6323,N_4037,N_5169);
and U6324 (N_6324,N_5381,N_4112);
nand U6325 (N_6325,N_5489,N_5779);
xnor U6326 (N_6326,N_5060,N_5878);
xor U6327 (N_6327,N_4045,N_5025);
xor U6328 (N_6328,N_4673,N_4703);
nand U6329 (N_6329,N_4906,N_4291);
nor U6330 (N_6330,N_5911,N_5813);
nand U6331 (N_6331,N_4747,N_4416);
and U6332 (N_6332,N_5782,N_4557);
or U6333 (N_6333,N_4529,N_5837);
and U6334 (N_6334,N_5308,N_4560);
nand U6335 (N_6335,N_4750,N_5967);
xnor U6336 (N_6336,N_5284,N_5267);
nor U6337 (N_6337,N_4695,N_4362);
and U6338 (N_6338,N_4829,N_5845);
xor U6339 (N_6339,N_4013,N_4076);
nand U6340 (N_6340,N_4895,N_5009);
or U6341 (N_6341,N_4303,N_4835);
and U6342 (N_6342,N_5174,N_5785);
xor U6343 (N_6343,N_4623,N_5217);
or U6344 (N_6344,N_5767,N_5115);
xor U6345 (N_6345,N_5259,N_5658);
xor U6346 (N_6346,N_5855,N_4978);
nor U6347 (N_6347,N_5864,N_5485);
nor U6348 (N_6348,N_4752,N_4833);
nor U6349 (N_6349,N_5794,N_4249);
and U6350 (N_6350,N_4169,N_4507);
and U6351 (N_6351,N_5053,N_4815);
and U6352 (N_6352,N_4634,N_5117);
nor U6353 (N_6353,N_4942,N_5479);
xnor U6354 (N_6354,N_5789,N_5854);
xor U6355 (N_6355,N_4215,N_4200);
or U6356 (N_6356,N_5827,N_4440);
nand U6357 (N_6357,N_5133,N_4405);
xor U6358 (N_6358,N_5694,N_5330);
and U6359 (N_6359,N_5161,N_5220);
or U6360 (N_6360,N_4897,N_4185);
and U6361 (N_6361,N_4671,N_5902);
xor U6362 (N_6362,N_5683,N_5764);
nand U6363 (N_6363,N_5403,N_5900);
nand U6364 (N_6364,N_4421,N_4104);
or U6365 (N_6365,N_4124,N_5379);
xnor U6366 (N_6366,N_4853,N_5278);
xor U6367 (N_6367,N_4523,N_5230);
nand U6368 (N_6368,N_4765,N_5225);
nand U6369 (N_6369,N_5725,N_5271);
and U6370 (N_6370,N_5709,N_5817);
and U6371 (N_6371,N_5964,N_5486);
and U6372 (N_6372,N_5893,N_5088);
and U6373 (N_6373,N_5572,N_5418);
xor U6374 (N_6374,N_5990,N_5213);
nor U6375 (N_6375,N_4041,N_5444);
nor U6376 (N_6376,N_4732,N_5210);
or U6377 (N_6377,N_5496,N_4816);
or U6378 (N_6378,N_4502,N_4475);
or U6379 (N_6379,N_5263,N_5369);
or U6380 (N_6380,N_4385,N_4970);
xnor U6381 (N_6381,N_4432,N_5735);
nand U6382 (N_6382,N_5713,N_4694);
nor U6383 (N_6383,N_5633,N_4874);
and U6384 (N_6384,N_4993,N_5283);
nor U6385 (N_6385,N_4683,N_4216);
and U6386 (N_6386,N_5310,N_4140);
nor U6387 (N_6387,N_5822,N_4517);
or U6388 (N_6388,N_5708,N_4980);
and U6389 (N_6389,N_4293,N_4479);
nand U6390 (N_6390,N_5970,N_4890);
xor U6391 (N_6391,N_5803,N_4455);
nand U6392 (N_6392,N_4532,N_4977);
nand U6393 (N_6393,N_4426,N_4845);
and U6394 (N_6394,N_4861,N_4438);
xor U6395 (N_6395,N_4288,N_5260);
nand U6396 (N_6396,N_4103,N_5745);
xor U6397 (N_6397,N_4340,N_4822);
nand U6398 (N_6398,N_5372,N_4591);
and U6399 (N_6399,N_5761,N_4119);
or U6400 (N_6400,N_5952,N_5195);
nor U6401 (N_6401,N_4760,N_4624);
and U6402 (N_6402,N_5848,N_4134);
and U6403 (N_6403,N_5039,N_4050);
xnor U6404 (N_6404,N_4847,N_4167);
or U6405 (N_6405,N_5081,N_5353);
or U6406 (N_6406,N_4713,N_4669);
nor U6407 (N_6407,N_5863,N_5976);
xor U6408 (N_6408,N_4328,N_5376);
nor U6409 (N_6409,N_5287,N_4191);
xnor U6410 (N_6410,N_5867,N_4132);
nand U6411 (N_6411,N_4509,N_4107);
nand U6412 (N_6412,N_5853,N_4806);
nand U6413 (N_6413,N_4343,N_5165);
nand U6414 (N_6414,N_4360,N_4846);
nand U6415 (N_6415,N_4525,N_5297);
xor U6416 (N_6416,N_5406,N_4289);
nor U6417 (N_6417,N_5306,N_4865);
nor U6418 (N_6418,N_5989,N_4608);
nand U6419 (N_6419,N_4577,N_4662);
nand U6420 (N_6420,N_4650,N_5130);
nor U6421 (N_6421,N_5686,N_4863);
xnor U6422 (N_6422,N_5397,N_5662);
nor U6423 (N_6423,N_4136,N_5689);
and U6424 (N_6424,N_4690,N_5383);
xnor U6425 (N_6425,N_5240,N_4117);
or U6426 (N_6426,N_5807,N_5393);
nand U6427 (N_6427,N_4598,N_5253);
xnor U6428 (N_6428,N_4984,N_5529);
xor U6429 (N_6429,N_5429,N_5589);
nand U6430 (N_6430,N_4969,N_5939);
nand U6431 (N_6431,N_5611,N_5746);
or U6432 (N_6432,N_4091,N_4870);
and U6433 (N_6433,N_4823,N_5722);
xnor U6434 (N_6434,N_4609,N_5938);
or U6435 (N_6435,N_4646,N_4297);
or U6436 (N_6436,N_4194,N_5307);
nor U6437 (N_6437,N_4917,N_4238);
xor U6438 (N_6438,N_5895,N_5050);
nand U6439 (N_6439,N_4710,N_4372);
or U6440 (N_6440,N_4849,N_4394);
and U6441 (N_6441,N_5438,N_4149);
xnor U6442 (N_6442,N_5234,N_5231);
nor U6443 (N_6443,N_5573,N_5289);
nand U6444 (N_6444,N_4613,N_5510);
xor U6445 (N_6445,N_4098,N_5995);
or U6446 (N_6446,N_4206,N_4862);
and U6447 (N_6447,N_5833,N_4472);
and U6448 (N_6448,N_4053,N_5354);
and U6449 (N_6449,N_5044,N_4170);
or U6450 (N_6450,N_4794,N_4564);
nand U6451 (N_6451,N_4146,N_5070);
or U6452 (N_6452,N_4729,N_5002);
or U6453 (N_6453,N_5342,N_4017);
or U6454 (N_6454,N_5899,N_4740);
nor U6455 (N_6455,N_5488,N_5549);
nand U6456 (N_6456,N_5507,N_5541);
nand U6457 (N_6457,N_4995,N_4469);
xor U6458 (N_6458,N_5835,N_4417);
nand U6459 (N_6459,N_5901,N_5503);
and U6460 (N_6460,N_4006,N_5634);
nand U6461 (N_6461,N_5856,N_4355);
and U6462 (N_6462,N_4280,N_5747);
xor U6463 (N_6463,N_5762,N_5998);
nor U6464 (N_6464,N_5800,N_5987);
or U6465 (N_6465,N_5018,N_4736);
and U6466 (N_6466,N_4795,N_5288);
and U6467 (N_6467,N_4922,N_4559);
xor U6468 (N_6468,N_5974,N_4990);
nor U6469 (N_6469,N_4031,N_4561);
xnor U6470 (N_6470,N_4958,N_4597);
nor U6471 (N_6471,N_4838,N_5844);
and U6472 (N_6472,N_5180,N_5593);
nor U6473 (N_6473,N_4120,N_4552);
and U6474 (N_6474,N_5512,N_4189);
nand U6475 (N_6475,N_5904,N_5015);
xor U6476 (N_6476,N_4382,N_4617);
nand U6477 (N_6477,N_4450,N_5414);
or U6478 (N_6478,N_5109,N_5742);
or U6479 (N_6479,N_4807,N_4963);
xnor U6480 (N_6480,N_5684,N_4180);
xor U6481 (N_6481,N_5065,N_5721);
and U6482 (N_6482,N_5598,N_4972);
nor U6483 (N_6483,N_5710,N_4587);
xnor U6484 (N_6484,N_4805,N_5578);
xor U6485 (N_6485,N_4453,N_4869);
xnor U6486 (N_6486,N_4855,N_5058);
or U6487 (N_6487,N_5337,N_4637);
nor U6488 (N_6488,N_4062,N_5973);
xor U6489 (N_6489,N_5723,N_5344);
xnor U6490 (N_6490,N_5866,N_4161);
nand U6491 (N_6491,N_5205,N_5465);
xor U6492 (N_6492,N_5423,N_5346);
or U6493 (N_6493,N_4444,N_5375);
nand U6494 (N_6494,N_4190,N_4569);
xor U6495 (N_6495,N_5650,N_4940);
and U6496 (N_6496,N_5171,N_5951);
nor U6497 (N_6497,N_5953,N_4179);
nand U6498 (N_6498,N_5450,N_5636);
nor U6499 (N_6499,N_5405,N_4487);
nor U6500 (N_6500,N_5440,N_4933);
or U6501 (N_6501,N_4626,N_5286);
or U6502 (N_6502,N_5185,N_5484);
xor U6503 (N_6503,N_5865,N_4766);
and U6504 (N_6504,N_4247,N_4012);
or U6505 (N_6505,N_5532,N_5506);
and U6506 (N_6506,N_4513,N_4700);
and U6507 (N_6507,N_5886,N_5966);
xnor U6508 (N_6508,N_4536,N_4607);
and U6509 (N_6509,N_5016,N_4629);
or U6510 (N_6510,N_4797,N_4761);
xnor U6511 (N_6511,N_5467,N_5364);
or U6512 (N_6512,N_4860,N_4867);
xor U6513 (N_6513,N_5138,N_4798);
and U6514 (N_6514,N_5711,N_5192);
or U6515 (N_6515,N_4834,N_5157);
or U6516 (N_6516,N_5268,N_5791);
or U6517 (N_6517,N_4019,N_4553);
nor U6518 (N_6518,N_5380,N_4779);
nand U6519 (N_6519,N_5797,N_5590);
xor U6520 (N_6520,N_5917,N_5300);
nor U6521 (N_6521,N_4742,N_5172);
xnor U6522 (N_6522,N_5387,N_5898);
nor U6523 (N_6523,N_5101,N_5236);
nor U6524 (N_6524,N_4085,N_4915);
and U6525 (N_6525,N_5580,N_5715);
and U6526 (N_6526,N_4089,N_4964);
and U6527 (N_6527,N_4880,N_5013);
nor U6528 (N_6528,N_5933,N_5734);
xor U6529 (N_6529,N_5923,N_4931);
or U6530 (N_6530,N_5524,N_4872);
nand U6531 (N_6531,N_4309,N_4712);
or U6532 (N_6532,N_4541,N_5102);
and U6533 (N_6533,N_5481,N_4056);
nand U6534 (N_6534,N_5458,N_4256);
and U6535 (N_6535,N_5435,N_5881);
and U6536 (N_6536,N_5077,N_4201);
xnor U6537 (N_6537,N_4105,N_5536);
xnor U6538 (N_6538,N_5302,N_4875);
nor U6539 (N_6539,N_4704,N_4009);
or U6540 (N_6540,N_5201,N_5470);
xnor U6541 (N_6541,N_5949,N_4396);
xnor U6542 (N_6542,N_4959,N_4198);
or U6543 (N_6543,N_5280,N_4125);
nand U6544 (N_6544,N_5556,N_4226);
nor U6545 (N_6545,N_4384,N_5846);
nand U6546 (N_6546,N_4176,N_5402);
and U6547 (N_6547,N_4222,N_5126);
nand U6548 (N_6548,N_4454,N_4205);
and U6549 (N_6549,N_5294,N_5520);
nand U6550 (N_6550,N_5872,N_5771);
nor U6551 (N_6551,N_4877,N_5888);
and U6552 (N_6552,N_5187,N_4457);
nand U6553 (N_6553,N_5823,N_5671);
nand U6554 (N_6554,N_5150,N_5643);
nand U6555 (N_6555,N_4935,N_4052);
and U6556 (N_6556,N_5698,N_5697);
xnor U6557 (N_6557,N_4866,N_5788);
nand U6558 (N_6558,N_4606,N_4886);
nand U6559 (N_6559,N_5620,N_4451);
nor U6560 (N_6560,N_5473,N_5301);
and U6561 (N_6561,N_4824,N_5699);
and U6562 (N_6562,N_5091,N_5335);
nor U6563 (N_6563,N_5090,N_5247);
nand U6564 (N_6564,N_4251,N_5258);
nor U6565 (N_6565,N_5410,N_4522);
and U6566 (N_6566,N_4099,N_5017);
and U6567 (N_6567,N_4352,N_4005);
nor U6568 (N_6568,N_4748,N_4893);
or U6569 (N_6569,N_4055,N_5239);
and U6570 (N_6570,N_4594,N_5903);
or U6571 (N_6571,N_5894,N_5535);
nor U6572 (N_6572,N_5769,N_5820);
or U6573 (N_6573,N_4582,N_4543);
nor U6574 (N_6574,N_5850,N_4021);
and U6575 (N_6575,N_4258,N_5879);
or U6576 (N_6576,N_4266,N_5112);
nor U6577 (N_6577,N_4057,N_4329);
xor U6578 (N_6578,N_5707,N_4086);
xnor U6579 (N_6579,N_5341,N_5431);
xnor U6580 (N_6580,N_5921,N_5685);
xnor U6581 (N_6581,N_5690,N_5274);
and U6582 (N_6582,N_4971,N_4034);
nand U6583 (N_6583,N_4635,N_4739);
and U6584 (N_6584,N_5838,N_5773);
and U6585 (N_6585,N_4084,N_5103);
and U6586 (N_6586,N_4027,N_5924);
nor U6587 (N_6587,N_5806,N_4499);
nor U6588 (N_6588,N_5607,N_4818);
or U6589 (N_6589,N_4468,N_4325);
nor U6590 (N_6590,N_5121,N_5047);
and U6591 (N_6591,N_5718,N_5143);
nand U6592 (N_6592,N_5732,N_4264);
nand U6593 (N_6593,N_4571,N_4749);
nor U6594 (N_6594,N_4425,N_5411);
and U6595 (N_6595,N_5985,N_5223);
and U6596 (N_6596,N_5537,N_4026);
xnor U6597 (N_6597,N_4447,N_5562);
xnor U6598 (N_6598,N_4836,N_5493);
nand U6599 (N_6599,N_4810,N_4839);
nor U6600 (N_6600,N_5812,N_4781);
or U6601 (N_6601,N_5055,N_5965);
nor U6602 (N_6602,N_4848,N_4706);
or U6603 (N_6603,N_4715,N_5443);
nand U6604 (N_6604,N_4771,N_5603);
xor U6605 (N_6605,N_4173,N_4418);
nor U6606 (N_6606,N_5564,N_5546);
xnor U6607 (N_6607,N_4400,N_5834);
xnor U6608 (N_6608,N_4786,N_4029);
nand U6609 (N_6609,N_5560,N_5934);
and U6610 (N_6610,N_4482,N_5222);
or U6611 (N_6611,N_5781,N_4312);
and U6612 (N_6612,N_5100,N_4358);
or U6613 (N_6613,N_5925,N_5490);
and U6614 (N_6614,N_5066,N_4648);
and U6615 (N_6615,N_4950,N_4000);
and U6616 (N_6616,N_4622,N_4974);
nand U6617 (N_6617,N_5432,N_5916);
xnor U6618 (N_6618,N_5480,N_4214);
and U6619 (N_6619,N_4693,N_5509);
and U6620 (N_6620,N_4390,N_5305);
or U6621 (N_6621,N_5775,N_4524);
or U6622 (N_6622,N_5219,N_5412);
xor U6623 (N_6623,N_4649,N_4619);
nand U6624 (N_6624,N_5669,N_4982);
and U6625 (N_6625,N_5084,N_4774);
nor U6626 (N_6626,N_5828,N_5716);
and U6627 (N_6627,N_4393,N_4991);
xor U6628 (N_6628,N_4889,N_4913);
nand U6629 (N_6629,N_4184,N_5770);
xor U6630 (N_6630,N_5605,N_5320);
and U6631 (N_6631,N_5281,N_4599);
nor U6632 (N_6632,N_5972,N_5692);
and U6633 (N_6633,N_4058,N_5419);
nor U6634 (N_6634,N_4016,N_5559);
and U6635 (N_6635,N_5420,N_5012);
or U6636 (N_6636,N_5548,N_5790);
nand U6637 (N_6637,N_4460,N_5581);
or U6638 (N_6638,N_4685,N_4059);
xnor U6639 (N_6639,N_5182,N_4678);
nand U6640 (N_6640,N_5874,N_5349);
or U6641 (N_6641,N_4651,N_5011);
nor U6642 (N_6642,N_4246,N_5358);
nand U6643 (N_6643,N_4985,N_5793);
or U6644 (N_6644,N_5497,N_4277);
nor U6645 (N_6645,N_5616,N_5910);
and U6646 (N_6646,N_5583,N_4368);
nand U6647 (N_6647,N_4883,N_5057);
or U6648 (N_6648,N_5628,N_5588);
or U6649 (N_6649,N_4002,N_4040);
nor U6650 (N_6650,N_5483,N_4620);
and U6651 (N_6651,N_4899,N_5599);
and U6652 (N_6652,N_4458,N_4230);
xor U6653 (N_6653,N_5421,N_4966);
nand U6654 (N_6654,N_5148,N_5469);
or U6655 (N_6655,N_5135,N_5424);
or U6656 (N_6656,N_4743,N_5738);
nor U6657 (N_6657,N_5763,N_4225);
nor U6658 (N_6658,N_4294,N_5113);
nor U6659 (N_6659,N_4504,N_5768);
xor U6660 (N_6660,N_4235,N_4562);
nor U6661 (N_6661,N_5038,N_4731);
nand U6662 (N_6662,N_4224,N_5075);
nand U6663 (N_6663,N_4388,N_5388);
or U6664 (N_6664,N_5787,N_5204);
or U6665 (N_6665,N_5107,N_4223);
or U6666 (N_6666,N_4614,N_4927);
nor U6667 (N_6667,N_4519,N_4925);
or U6668 (N_6668,N_4109,N_5005);
nand U6669 (N_6669,N_5255,N_4278);
xnor U6670 (N_6670,N_5362,N_4891);
nor U6671 (N_6671,N_5334,N_5365);
or U6672 (N_6672,N_4812,N_5566);
nor U6673 (N_6673,N_4403,N_5986);
nand U6674 (N_6674,N_5642,N_4645);
and U6675 (N_6675,N_5594,N_5368);
nor U6676 (N_6676,N_5655,N_5670);
and U6677 (N_6677,N_5272,N_4592);
nand U6678 (N_6678,N_5183,N_5453);
nand U6679 (N_6679,N_5394,N_5269);
and U6680 (N_6680,N_4638,N_5912);
or U6681 (N_6681,N_4533,N_5703);
and U6682 (N_6682,N_5328,N_4556);
or U6683 (N_6683,N_4539,N_5744);
nand U6684 (N_6684,N_4139,N_5945);
and U6685 (N_6685,N_5356,N_4983);
xnor U6686 (N_6686,N_5046,N_4654);
or U6687 (N_6687,N_5691,N_5241);
and U6688 (N_6688,N_5477,N_5825);
or U6689 (N_6689,N_5249,N_5144);
nor U6690 (N_6690,N_5547,N_5632);
or U6691 (N_6691,N_4711,N_4563);
nor U6692 (N_6692,N_5777,N_5006);
nor U6693 (N_6693,N_4165,N_4800);
xor U6694 (N_6694,N_4423,N_4784);
nor U6695 (N_6695,N_5545,N_5561);
or U6696 (N_6696,N_4492,N_4699);
nor U6697 (N_6697,N_4934,N_5427);
xor U6698 (N_6698,N_4462,N_4046);
xor U6699 (N_6699,N_4383,N_4181);
xor U6700 (N_6700,N_4682,N_4767);
nor U6701 (N_6701,N_4113,N_4338);
or U6702 (N_6702,N_4014,N_5391);
nand U6703 (N_6703,N_4321,N_4408);
nand U6704 (N_6704,N_5226,N_4315);
nand U6705 (N_6705,N_5366,N_4106);
or U6706 (N_6706,N_5714,N_4412);
nand U6707 (N_6707,N_4336,N_5245);
or U6708 (N_6708,N_5212,N_4066);
xor U6709 (N_6709,N_5675,N_5401);
nand U6710 (N_6710,N_4803,N_4495);
and U6711 (N_6711,N_4647,N_4413);
xor U6712 (N_6712,N_5852,N_5285);
xnor U6713 (N_6713,N_4854,N_4364);
and U6714 (N_6714,N_5233,N_5720);
and U6715 (N_6715,N_5445,N_4547);
nand U6716 (N_6716,N_4814,N_5609);
or U6717 (N_6717,N_4327,N_4357);
nor U6718 (N_6718,N_4048,N_4551);
and U6719 (N_6719,N_4962,N_4631);
and U6720 (N_6720,N_5007,N_4464);
and U6721 (N_6721,N_5577,N_5754);
nand U6722 (N_6722,N_5883,N_4530);
nor U6723 (N_6723,N_4655,N_5048);
nand U6724 (N_6724,N_5378,N_4570);
nand U6725 (N_6725,N_5815,N_4549);
nor U6726 (N_6726,N_5051,N_4168);
and U6727 (N_6727,N_4926,N_4044);
nor U6728 (N_6728,N_5322,N_4465);
and U6729 (N_6729,N_5914,N_5494);
nand U6730 (N_6730,N_4141,N_5988);
and U6731 (N_6731,N_4111,N_5068);
xor U6732 (N_6732,N_4166,N_5937);
and U6733 (N_6733,N_5727,N_4292);
nor U6734 (N_6734,N_5739,N_5724);
nand U6735 (N_6735,N_4158,N_4565);
xor U6736 (N_6736,N_4627,N_4375);
and U6737 (N_6737,N_4243,N_4879);
nor U6738 (N_6738,N_5336,N_4644);
or U6739 (N_6739,N_4672,N_5238);
nor U6740 (N_6740,N_5882,N_5656);
or U6741 (N_6741,N_5639,N_5279);
xor U6742 (N_6742,N_5700,N_4381);
or U6743 (N_6743,N_5384,N_4070);
nand U6744 (N_6744,N_5750,N_5129);
and U6745 (N_6745,N_4717,N_4043);
nor U6746 (N_6746,N_5357,N_5460);
nand U6747 (N_6747,N_4378,N_4137);
and U6748 (N_6748,N_5623,N_5252);
or U6749 (N_6749,N_4809,N_5400);
nor U6750 (N_6750,N_5452,N_4242);
nand U6751 (N_6751,N_4554,N_5892);
xor U6752 (N_6752,N_4579,N_4363);
xnor U6753 (N_6753,N_4489,N_4769);
xnor U6754 (N_6754,N_4307,N_5926);
and U6755 (N_6755,N_4796,N_4069);
nor U6756 (N_6756,N_4753,N_4821);
and U6757 (N_6757,N_5087,N_4354);
or U6758 (N_6758,N_4936,N_5652);
xnor U6759 (N_6759,N_5518,N_5282);
nand U6760 (N_6760,N_4939,N_4441);
nand U6761 (N_6761,N_5374,N_4688);
xnor U6762 (N_6762,N_5295,N_4998);
xnor U6763 (N_6763,N_5447,N_4095);
nand U6764 (N_6764,N_4745,N_4296);
xnor U6765 (N_6765,N_5189,N_5069);
and U6766 (N_6766,N_4568,N_5303);
and U6767 (N_6767,N_5802,N_4887);
nand U6768 (N_6768,N_5673,N_4466);
nor U6769 (N_6769,N_5897,N_4965);
and U6770 (N_6770,N_5751,N_4961);
and U6771 (N_6771,N_5311,N_4772);
xnor U6772 (N_6772,N_4947,N_5999);
and U6773 (N_6773,N_5425,N_5437);
xnor U6774 (N_6774,N_4503,N_5430);
or U6775 (N_6775,N_4914,N_5551);
or U6776 (N_6776,N_4300,N_4376);
or U6777 (N_6777,N_4584,N_4424);
or U6778 (N_6778,N_4738,N_5035);
nor U6779 (N_6779,N_5826,N_5681);
and U6780 (N_6780,N_4407,N_4221);
nor U6781 (N_6781,N_5876,N_5568);
xor U6782 (N_6782,N_5693,N_5570);
nor U6783 (N_6783,N_5029,N_5074);
nand U6784 (N_6784,N_5935,N_5647);
nand U6785 (N_6785,N_4071,N_5036);
and U6786 (N_6786,N_5913,N_4233);
nand U6787 (N_6787,N_5085,N_5347);
and U6788 (N_6788,N_4268,N_4456);
nor U6789 (N_6789,N_4728,N_5208);
xnor U6790 (N_6790,N_5843,N_5774);
nand U6791 (N_6791,N_5530,N_5167);
nor U6792 (N_6792,N_4151,N_5621);
or U6793 (N_6793,N_5312,N_4488);
or U6794 (N_6794,N_5759,N_4896);
xor U6795 (N_6795,N_4422,N_5663);
or U6796 (N_6796,N_5955,N_4828);
xnor U6797 (N_6797,N_5123,N_4330);
or U6798 (N_6798,N_4154,N_4892);
nand U6799 (N_6799,N_4576,N_4186);
nor U6800 (N_6800,N_4121,N_4790);
and U6801 (N_6801,N_4808,N_5149);
nor U6802 (N_6802,N_4001,N_5162);
nand U6803 (N_6803,N_4263,N_4632);
nor U6804 (N_6804,N_5186,N_4843);
nor U6805 (N_6805,N_4061,N_5457);
and U6806 (N_6806,N_4544,N_5299);
or U6807 (N_6807,N_5367,N_4253);
nor U6808 (N_6808,N_5571,N_5371);
or U6809 (N_6809,N_5151,N_4949);
and U6810 (N_6810,N_5954,N_4526);
nor U6811 (N_6811,N_5810,N_4347);
or U6812 (N_6812,N_5946,N_5606);
and U6813 (N_6813,N_4157,N_4486);
nand U6814 (N_6814,N_5753,N_4399);
nor U6815 (N_6815,N_4696,N_5191);
or U6816 (N_6816,N_4921,N_5765);
xnor U6817 (N_6817,N_4199,N_5385);
and U6818 (N_6818,N_4467,N_5108);
nand U6819 (N_6819,N_4528,N_5857);
and U6820 (N_6820,N_5534,N_5682);
nor U6821 (N_6821,N_4459,N_5640);
nor U6822 (N_6822,N_4319,N_5840);
xnor U6823 (N_6823,N_5089,N_5654);
nand U6824 (N_6824,N_4658,N_5672);
and U6825 (N_6825,N_4102,N_5168);
and U6826 (N_6826,N_5042,N_4490);
xnor U6827 (N_6827,N_4197,N_4370);
nor U6828 (N_6828,N_4832,N_4212);
nor U6829 (N_6829,N_4114,N_4279);
nor U6830 (N_6830,N_5635,N_5059);
and U6831 (N_6831,N_4373,N_4219);
xnor U6832 (N_6832,N_4988,N_5237);
and U6833 (N_6833,N_4692,N_4677);
or U6834 (N_6834,N_5805,N_5511);
xor U6835 (N_6835,N_4419,N_4007);
xnor U6836 (N_6836,N_4208,N_5958);
and U6837 (N_6837,N_5552,N_4387);
or U6838 (N_6838,N_4542,N_5956);
and U6839 (N_6839,N_5024,N_5056);
nor U6840 (N_6840,N_5851,N_4759);
and U6841 (N_6841,N_4811,N_4449);
nand U6842 (N_6842,N_5122,N_4304);
xor U6843 (N_6843,N_4042,N_5073);
nand U6844 (N_6844,N_5163,N_5638);
or U6845 (N_6845,N_5625,N_4773);
or U6846 (N_6846,N_5355,N_4793);
nor U6847 (N_6847,N_4929,N_4342);
or U6848 (N_6848,N_4953,N_4162);
nor U6849 (N_6849,N_4697,N_5558);
nor U6850 (N_6850,N_4270,N_5799);
or U6851 (N_6851,N_4110,N_4540);
nand U6852 (N_6852,N_5741,N_4209);
nand U6853 (N_6853,N_4788,N_4038);
or U6854 (N_6854,N_4077,N_4770);
nor U6855 (N_6855,N_5246,N_4150);
and U6856 (N_6856,N_5516,N_5474);
xor U6857 (N_6857,N_5877,N_4333);
and U6858 (N_6858,N_5207,N_4537);
nor U6859 (N_6859,N_4830,N_4317);
or U6860 (N_6860,N_4733,N_4448);
or U6861 (N_6861,N_4122,N_5094);
or U6862 (N_6862,N_5585,N_5416);
or U6863 (N_6863,N_5040,N_4339);
nor U6864 (N_6864,N_5475,N_5390);
nor U6865 (N_6865,N_4518,N_4709);
or U6866 (N_6866,N_5795,N_4100);
nor U6867 (N_6867,N_5668,N_5730);
nor U6868 (N_6868,N_5804,N_5454);
xor U6869 (N_6869,N_5831,N_5991);
and U6870 (N_6870,N_5980,N_4762);
nor U6871 (N_6871,N_4135,N_5977);
nor U6872 (N_6872,N_4335,N_5043);
and U6873 (N_6873,N_5028,N_5173);
nand U6874 (N_6874,N_4367,N_4244);
or U6875 (N_6875,N_4175,N_4660);
and U6876 (N_6876,N_4313,N_4024);
xor U6877 (N_6877,N_4349,N_5316);
xor U6878 (N_6878,N_4586,N_4573);
nand U6879 (N_6879,N_4092,N_5325);
or U6880 (N_6880,N_5997,N_5619);
or U6881 (N_6881,N_4097,N_5265);
xor U6882 (N_6882,N_4285,N_4639);
xor U6883 (N_6883,N_5478,N_5760);
nand U6884 (N_6884,N_5719,N_5232);
or U6885 (N_6885,N_5200,N_4698);
nor U6886 (N_6886,N_4831,N_5114);
nand U6887 (N_6887,N_5266,N_5657);
nand U6888 (N_6888,N_5152,N_4817);
xor U6889 (N_6889,N_4868,N_4240);
and U6890 (N_6890,N_5502,N_4023);
and U6891 (N_6891,N_5575,N_5660);
and U6892 (N_6892,N_4842,N_5142);
or U6893 (N_6893,N_5003,N_5348);
nand U6894 (N_6894,N_5293,N_4254);
or U6895 (N_6895,N_4535,N_5331);
nand U6896 (N_6896,N_4783,N_5766);
xnor U6897 (N_6897,N_5261,N_4302);
or U6898 (N_6898,N_4976,N_5614);
nor U6899 (N_6899,N_5211,N_5629);
nand U6900 (N_6900,N_5565,N_5455);
nor U6901 (N_6901,N_5758,N_5426);
or U6902 (N_6902,N_5188,N_4324);
nor U6903 (N_6903,N_5023,N_4628);
or U6904 (N_6904,N_4204,N_4207);
nor U6905 (N_6905,N_4195,N_4391);
or U6906 (N_6906,N_5010,N_4159);
and U6907 (N_6907,N_5992,N_4231);
xor U6908 (N_6908,N_5120,N_5808);
or U6909 (N_6909,N_4074,N_4081);
or U6910 (N_6910,N_5602,N_4356);
xor U6911 (N_6911,N_4656,N_4241);
and U6912 (N_6912,N_5798,N_4837);
nor U6913 (N_6913,N_5022,N_5809);
nand U6914 (N_6914,N_4670,N_5941);
and U6915 (N_6915,N_5463,N_4148);
and U6916 (N_6916,N_4575,N_4943);
nand U6917 (N_6917,N_5139,N_4768);
xor U6918 (N_6918,N_5395,N_4718);
nor U6919 (N_6919,N_4470,N_5462);
nand U6920 (N_6920,N_5034,N_5940);
nand U6921 (N_6921,N_4721,N_5533);
nand U6922 (N_6922,N_4602,N_5327);
nand U6923 (N_6923,N_5702,N_5392);
nor U6924 (N_6924,N_5783,N_4514);
and U6925 (N_6925,N_5664,N_5756);
xnor U6926 (N_6926,N_5032,N_4756);
or U6927 (N_6927,N_5318,N_4920);
nand U6928 (N_6928,N_4827,N_4884);
nand U6929 (N_6929,N_4724,N_4780);
nand U6930 (N_6930,N_4108,N_5927);
nand U6931 (N_6931,N_4684,N_4428);
xor U6932 (N_6932,N_5221,N_4142);
and U6933 (N_6933,N_4701,N_4144);
or U6934 (N_6934,N_4657,N_5544);
and U6935 (N_6935,N_5950,N_4353);
xnor U6936 (N_6936,N_4477,N_5860);
and U6937 (N_6937,N_5382,N_5748);
or U6938 (N_6938,N_5389,N_4434);
and U6939 (N_6939,N_5929,N_5154);
nand U6940 (N_6940,N_4894,N_5021);
and U6941 (N_6941,N_4348,N_4182);
xnor U6942 (N_6942,N_5128,N_5870);
nor U6943 (N_6943,N_4550,N_4986);
and U6944 (N_6944,N_5687,N_4004);
nor U6945 (N_6945,N_5449,N_5273);
nor U6946 (N_6946,N_5776,N_5859);
or U6947 (N_6947,N_5880,N_5784);
and U6948 (N_6948,N_4668,N_5841);
nand U6949 (N_6949,N_4725,N_5027);
xor U6950 (N_6950,N_4493,N_4088);
and U6951 (N_6951,N_5830,N_5408);
or U6952 (N_6952,N_4946,N_5944);
nor U6953 (N_6953,N_5004,N_4188);
nand U6954 (N_6954,N_5194,N_4819);
nor U6955 (N_6955,N_5948,N_4072);
or U6956 (N_6956,N_4192,N_4566);
nor U6957 (N_6957,N_4799,N_4237);
xor U6958 (N_6958,N_5842,N_5275);
and U6959 (N_6959,N_5752,N_5468);
and U6960 (N_6960,N_4445,N_5889);
or U6961 (N_6961,N_4994,N_4332);
nand U6962 (N_6962,N_5339,N_5229);
and U6963 (N_6963,N_4932,N_4174);
and U6964 (N_6964,N_5947,N_5696);
nand U6965 (N_6965,N_4402,N_4397);
or U6966 (N_6966,N_5276,N_5030);
xnor U6967 (N_6967,N_4714,N_4366);
or U6968 (N_6968,N_4047,N_4652);
nand U6969 (N_6969,N_4928,N_4299);
or U6970 (N_6970,N_4272,N_5557);
or U6971 (N_6971,N_5487,N_4282);
or U6972 (N_6972,N_4359,N_5554);
xnor U6973 (N_6973,N_4621,N_4789);
nand U6974 (N_6974,N_5626,N_4320);
nor U6975 (N_6975,N_5049,N_4369);
nand U6976 (N_6976,N_4371,N_5277);
nor U6977 (N_6977,N_4987,N_4018);
or U6978 (N_6978,N_4250,N_4033);
nand U6979 (N_6979,N_5818,N_4705);
xnor U6980 (N_6980,N_5871,N_5930);
nand U6981 (N_6981,N_5517,N_5456);
xnor U6982 (N_6982,N_5441,N_5323);
nand U6983 (N_6983,N_5919,N_4775);
nor U6984 (N_6984,N_4864,N_5156);
xor U6985 (N_6985,N_4616,N_5597);
or U6986 (N_6986,N_4361,N_5829);
or U6987 (N_6987,N_4156,N_5542);
nor U6988 (N_6988,N_4531,N_4476);
or U6989 (N_6989,N_4063,N_4973);
nor U6990 (N_6990,N_4123,N_5726);
and U6991 (N_6991,N_4741,N_5615);
and U6992 (N_6992,N_4163,N_4702);
xnor U6993 (N_6993,N_5624,N_5145);
and U6994 (N_6994,N_4506,N_5971);
nor U6995 (N_6995,N_4217,N_5816);
or U6996 (N_6996,N_5386,N_5064);
nor U6997 (N_6997,N_4287,N_4981);
or U6998 (N_6998,N_5345,N_5996);
or U6999 (N_6999,N_4064,N_4975);
nor U7000 (N_7000,N_4364,N_4020);
nor U7001 (N_7001,N_5368,N_4176);
xnor U7002 (N_7002,N_4575,N_4159);
and U7003 (N_7003,N_5662,N_5828);
or U7004 (N_7004,N_5283,N_5070);
nand U7005 (N_7005,N_4595,N_5869);
nand U7006 (N_7006,N_4571,N_4704);
nand U7007 (N_7007,N_4924,N_5933);
xnor U7008 (N_7008,N_4040,N_4156);
nand U7009 (N_7009,N_5749,N_5599);
or U7010 (N_7010,N_5784,N_5535);
nor U7011 (N_7011,N_4123,N_4454);
xnor U7012 (N_7012,N_4611,N_4972);
and U7013 (N_7013,N_5451,N_5598);
nor U7014 (N_7014,N_4619,N_4192);
or U7015 (N_7015,N_5813,N_4474);
or U7016 (N_7016,N_5333,N_5405);
xnor U7017 (N_7017,N_5026,N_5441);
or U7018 (N_7018,N_5192,N_4517);
xnor U7019 (N_7019,N_5883,N_5457);
xor U7020 (N_7020,N_4017,N_5739);
or U7021 (N_7021,N_4283,N_5424);
nor U7022 (N_7022,N_4817,N_5245);
and U7023 (N_7023,N_5982,N_4531);
nor U7024 (N_7024,N_5291,N_5778);
or U7025 (N_7025,N_5567,N_5962);
or U7026 (N_7026,N_5226,N_5671);
xor U7027 (N_7027,N_4463,N_5200);
xnor U7028 (N_7028,N_5358,N_5588);
or U7029 (N_7029,N_4994,N_4250);
nand U7030 (N_7030,N_5228,N_5040);
nand U7031 (N_7031,N_5410,N_5568);
or U7032 (N_7032,N_5307,N_4830);
xor U7033 (N_7033,N_4032,N_5012);
and U7034 (N_7034,N_5915,N_4508);
and U7035 (N_7035,N_5689,N_5216);
nor U7036 (N_7036,N_4435,N_5143);
or U7037 (N_7037,N_5360,N_4733);
nor U7038 (N_7038,N_4725,N_5295);
and U7039 (N_7039,N_4425,N_4488);
or U7040 (N_7040,N_5120,N_5896);
xor U7041 (N_7041,N_5468,N_5505);
and U7042 (N_7042,N_4826,N_5907);
nand U7043 (N_7043,N_4899,N_4995);
or U7044 (N_7044,N_5278,N_4096);
or U7045 (N_7045,N_5561,N_4474);
and U7046 (N_7046,N_5305,N_4033);
nor U7047 (N_7047,N_5443,N_5706);
nand U7048 (N_7048,N_5417,N_4986);
or U7049 (N_7049,N_5035,N_4480);
nand U7050 (N_7050,N_5562,N_4821);
and U7051 (N_7051,N_5532,N_4756);
xor U7052 (N_7052,N_5137,N_4729);
or U7053 (N_7053,N_4561,N_5033);
nand U7054 (N_7054,N_5268,N_4420);
or U7055 (N_7055,N_5850,N_5210);
nor U7056 (N_7056,N_5003,N_4686);
xor U7057 (N_7057,N_5081,N_5612);
and U7058 (N_7058,N_5751,N_4813);
and U7059 (N_7059,N_5134,N_5337);
nand U7060 (N_7060,N_5944,N_5977);
nor U7061 (N_7061,N_4327,N_5132);
or U7062 (N_7062,N_4845,N_4411);
nor U7063 (N_7063,N_5942,N_4464);
or U7064 (N_7064,N_5447,N_4394);
xor U7065 (N_7065,N_5591,N_4043);
nand U7066 (N_7066,N_4352,N_4337);
and U7067 (N_7067,N_4906,N_4275);
nand U7068 (N_7068,N_5074,N_4963);
nor U7069 (N_7069,N_5157,N_5610);
nand U7070 (N_7070,N_5306,N_5040);
or U7071 (N_7071,N_5804,N_5862);
nor U7072 (N_7072,N_5984,N_4858);
xnor U7073 (N_7073,N_5110,N_4224);
or U7074 (N_7074,N_5487,N_4573);
xnor U7075 (N_7075,N_5512,N_4663);
nor U7076 (N_7076,N_5855,N_5205);
and U7077 (N_7077,N_5515,N_4472);
nand U7078 (N_7078,N_4684,N_5130);
xor U7079 (N_7079,N_5809,N_5399);
nand U7080 (N_7080,N_5780,N_5771);
nor U7081 (N_7081,N_4588,N_5594);
nand U7082 (N_7082,N_5073,N_4822);
and U7083 (N_7083,N_4018,N_5302);
nand U7084 (N_7084,N_5010,N_5789);
or U7085 (N_7085,N_5518,N_4992);
nand U7086 (N_7086,N_5474,N_5624);
xor U7087 (N_7087,N_4049,N_4030);
and U7088 (N_7088,N_5546,N_4805);
nor U7089 (N_7089,N_5875,N_5533);
nor U7090 (N_7090,N_4590,N_5048);
and U7091 (N_7091,N_5177,N_4073);
or U7092 (N_7092,N_5401,N_5246);
nor U7093 (N_7093,N_4209,N_4690);
and U7094 (N_7094,N_4128,N_5187);
nand U7095 (N_7095,N_5483,N_5275);
nor U7096 (N_7096,N_4854,N_5940);
nor U7097 (N_7097,N_5935,N_5308);
and U7098 (N_7098,N_5565,N_4382);
or U7099 (N_7099,N_5239,N_4341);
nor U7100 (N_7100,N_5313,N_4637);
xor U7101 (N_7101,N_4959,N_4736);
nor U7102 (N_7102,N_4745,N_5396);
and U7103 (N_7103,N_4290,N_5963);
xor U7104 (N_7104,N_5609,N_4645);
nand U7105 (N_7105,N_4836,N_5566);
nand U7106 (N_7106,N_4762,N_5413);
nor U7107 (N_7107,N_4986,N_4431);
nand U7108 (N_7108,N_4727,N_5082);
nand U7109 (N_7109,N_4710,N_5923);
or U7110 (N_7110,N_5472,N_5265);
and U7111 (N_7111,N_4980,N_4303);
nor U7112 (N_7112,N_4132,N_4872);
nand U7113 (N_7113,N_5762,N_4328);
nand U7114 (N_7114,N_4696,N_5941);
and U7115 (N_7115,N_4411,N_5902);
nand U7116 (N_7116,N_5350,N_4896);
or U7117 (N_7117,N_4420,N_5260);
xor U7118 (N_7118,N_4009,N_4317);
nand U7119 (N_7119,N_5848,N_4679);
nand U7120 (N_7120,N_4873,N_5795);
and U7121 (N_7121,N_5856,N_5302);
nand U7122 (N_7122,N_4491,N_5854);
or U7123 (N_7123,N_5324,N_5409);
xor U7124 (N_7124,N_4159,N_5930);
nand U7125 (N_7125,N_5507,N_5783);
nor U7126 (N_7126,N_4067,N_5982);
or U7127 (N_7127,N_4889,N_4290);
and U7128 (N_7128,N_4623,N_4126);
or U7129 (N_7129,N_4920,N_5382);
or U7130 (N_7130,N_5615,N_4398);
nor U7131 (N_7131,N_5546,N_4703);
nand U7132 (N_7132,N_4998,N_5517);
xor U7133 (N_7133,N_5037,N_4157);
or U7134 (N_7134,N_4649,N_4334);
xor U7135 (N_7135,N_5240,N_4831);
and U7136 (N_7136,N_5439,N_4121);
or U7137 (N_7137,N_4284,N_4643);
xor U7138 (N_7138,N_4006,N_4961);
xnor U7139 (N_7139,N_5730,N_4580);
nor U7140 (N_7140,N_4086,N_5017);
or U7141 (N_7141,N_4880,N_5654);
or U7142 (N_7142,N_4750,N_4543);
nor U7143 (N_7143,N_5996,N_4158);
and U7144 (N_7144,N_4614,N_5101);
and U7145 (N_7145,N_5748,N_5809);
nand U7146 (N_7146,N_4190,N_5576);
nor U7147 (N_7147,N_5619,N_4855);
and U7148 (N_7148,N_4388,N_4551);
nand U7149 (N_7149,N_5055,N_5777);
or U7150 (N_7150,N_4066,N_5322);
xnor U7151 (N_7151,N_5613,N_5594);
xnor U7152 (N_7152,N_4408,N_5694);
and U7153 (N_7153,N_5330,N_5319);
or U7154 (N_7154,N_5796,N_5869);
nand U7155 (N_7155,N_4396,N_4020);
or U7156 (N_7156,N_5139,N_5014);
nor U7157 (N_7157,N_4004,N_4368);
nor U7158 (N_7158,N_4712,N_4243);
xor U7159 (N_7159,N_5790,N_4819);
nand U7160 (N_7160,N_4882,N_5560);
and U7161 (N_7161,N_4725,N_4677);
xnor U7162 (N_7162,N_5679,N_5736);
nand U7163 (N_7163,N_5591,N_4160);
or U7164 (N_7164,N_5663,N_5470);
and U7165 (N_7165,N_5324,N_5175);
or U7166 (N_7166,N_4766,N_5136);
nor U7167 (N_7167,N_4501,N_4423);
xnor U7168 (N_7168,N_4916,N_4444);
nand U7169 (N_7169,N_4708,N_5532);
nand U7170 (N_7170,N_5875,N_4948);
or U7171 (N_7171,N_4172,N_4471);
or U7172 (N_7172,N_5280,N_4616);
nand U7173 (N_7173,N_5403,N_4813);
or U7174 (N_7174,N_4240,N_4942);
xor U7175 (N_7175,N_4081,N_4810);
xnor U7176 (N_7176,N_5299,N_4525);
nor U7177 (N_7177,N_5818,N_4711);
nand U7178 (N_7178,N_5840,N_4857);
or U7179 (N_7179,N_5874,N_4620);
or U7180 (N_7180,N_5596,N_5927);
and U7181 (N_7181,N_5429,N_4341);
xnor U7182 (N_7182,N_4910,N_5354);
nand U7183 (N_7183,N_4120,N_4984);
nand U7184 (N_7184,N_4730,N_4466);
xnor U7185 (N_7185,N_4099,N_5093);
nor U7186 (N_7186,N_5756,N_5090);
nand U7187 (N_7187,N_5711,N_4828);
and U7188 (N_7188,N_5155,N_4161);
nand U7189 (N_7189,N_4370,N_5436);
nand U7190 (N_7190,N_5881,N_5010);
nor U7191 (N_7191,N_4634,N_5305);
and U7192 (N_7192,N_5703,N_4190);
or U7193 (N_7193,N_4486,N_5578);
nand U7194 (N_7194,N_5176,N_5081);
nor U7195 (N_7195,N_4267,N_5812);
nor U7196 (N_7196,N_5947,N_4392);
xor U7197 (N_7197,N_5125,N_5710);
or U7198 (N_7198,N_4471,N_5165);
nor U7199 (N_7199,N_4002,N_5323);
or U7200 (N_7200,N_5000,N_4742);
and U7201 (N_7201,N_4167,N_5194);
and U7202 (N_7202,N_5660,N_4930);
nand U7203 (N_7203,N_4807,N_4329);
nor U7204 (N_7204,N_4310,N_4278);
xnor U7205 (N_7205,N_5267,N_5824);
and U7206 (N_7206,N_4201,N_5760);
nor U7207 (N_7207,N_4286,N_4634);
or U7208 (N_7208,N_5764,N_4821);
xnor U7209 (N_7209,N_4346,N_5089);
or U7210 (N_7210,N_5707,N_5329);
nand U7211 (N_7211,N_4261,N_5779);
nand U7212 (N_7212,N_4575,N_5290);
or U7213 (N_7213,N_5412,N_5479);
or U7214 (N_7214,N_5544,N_5572);
and U7215 (N_7215,N_4770,N_4913);
or U7216 (N_7216,N_4644,N_5833);
nand U7217 (N_7217,N_5099,N_4007);
or U7218 (N_7218,N_5822,N_4246);
and U7219 (N_7219,N_5316,N_5119);
nand U7220 (N_7220,N_4758,N_5975);
or U7221 (N_7221,N_4669,N_4993);
nor U7222 (N_7222,N_5222,N_5271);
xnor U7223 (N_7223,N_5347,N_5847);
nand U7224 (N_7224,N_5494,N_5718);
nor U7225 (N_7225,N_5596,N_4821);
xnor U7226 (N_7226,N_4905,N_5902);
xnor U7227 (N_7227,N_4217,N_4658);
nand U7228 (N_7228,N_4263,N_5484);
nand U7229 (N_7229,N_4144,N_5339);
xor U7230 (N_7230,N_5051,N_4770);
nand U7231 (N_7231,N_5162,N_5192);
xnor U7232 (N_7232,N_4916,N_4380);
xor U7233 (N_7233,N_4285,N_4430);
nor U7234 (N_7234,N_5909,N_4685);
and U7235 (N_7235,N_5810,N_4846);
nor U7236 (N_7236,N_5731,N_4281);
nor U7237 (N_7237,N_4348,N_5574);
or U7238 (N_7238,N_5319,N_4985);
or U7239 (N_7239,N_5430,N_5359);
and U7240 (N_7240,N_4003,N_4159);
nor U7241 (N_7241,N_5301,N_4441);
nand U7242 (N_7242,N_5735,N_4921);
and U7243 (N_7243,N_5672,N_5779);
nand U7244 (N_7244,N_5049,N_4997);
and U7245 (N_7245,N_5965,N_4725);
nand U7246 (N_7246,N_5756,N_4423);
or U7247 (N_7247,N_4588,N_4952);
or U7248 (N_7248,N_5141,N_5043);
or U7249 (N_7249,N_5548,N_4701);
and U7250 (N_7250,N_4452,N_4046);
nor U7251 (N_7251,N_5377,N_4751);
or U7252 (N_7252,N_5202,N_4804);
or U7253 (N_7253,N_5332,N_4966);
and U7254 (N_7254,N_5365,N_5508);
and U7255 (N_7255,N_4584,N_4525);
nor U7256 (N_7256,N_5610,N_5105);
nand U7257 (N_7257,N_5173,N_5376);
or U7258 (N_7258,N_5634,N_4684);
and U7259 (N_7259,N_4693,N_5895);
nor U7260 (N_7260,N_4806,N_4114);
nor U7261 (N_7261,N_5804,N_4604);
nand U7262 (N_7262,N_4491,N_4745);
or U7263 (N_7263,N_4448,N_5262);
or U7264 (N_7264,N_4159,N_4483);
and U7265 (N_7265,N_4413,N_4681);
and U7266 (N_7266,N_5108,N_5241);
nor U7267 (N_7267,N_5382,N_5472);
nor U7268 (N_7268,N_4093,N_4985);
or U7269 (N_7269,N_5540,N_4833);
nor U7270 (N_7270,N_5252,N_4552);
or U7271 (N_7271,N_5488,N_5707);
and U7272 (N_7272,N_4975,N_4971);
nor U7273 (N_7273,N_5575,N_5728);
or U7274 (N_7274,N_5509,N_5291);
nand U7275 (N_7275,N_5947,N_4235);
and U7276 (N_7276,N_4514,N_4769);
nand U7277 (N_7277,N_5898,N_5069);
and U7278 (N_7278,N_4453,N_5069);
xor U7279 (N_7279,N_5600,N_5111);
nor U7280 (N_7280,N_5690,N_5942);
and U7281 (N_7281,N_5639,N_5748);
xor U7282 (N_7282,N_4508,N_4885);
xor U7283 (N_7283,N_5044,N_4960);
or U7284 (N_7284,N_5047,N_4695);
or U7285 (N_7285,N_5915,N_4862);
and U7286 (N_7286,N_4629,N_4617);
nor U7287 (N_7287,N_4986,N_4699);
nand U7288 (N_7288,N_5807,N_5971);
and U7289 (N_7289,N_5465,N_4362);
nor U7290 (N_7290,N_5795,N_4571);
nor U7291 (N_7291,N_4053,N_5509);
nor U7292 (N_7292,N_5841,N_4109);
or U7293 (N_7293,N_5026,N_4171);
and U7294 (N_7294,N_4908,N_4366);
xnor U7295 (N_7295,N_4486,N_5658);
and U7296 (N_7296,N_4204,N_5253);
xor U7297 (N_7297,N_5500,N_5552);
or U7298 (N_7298,N_5338,N_5075);
xor U7299 (N_7299,N_4542,N_5688);
xor U7300 (N_7300,N_4956,N_5419);
nand U7301 (N_7301,N_5667,N_4743);
or U7302 (N_7302,N_5018,N_4165);
and U7303 (N_7303,N_4854,N_4633);
and U7304 (N_7304,N_4636,N_4918);
or U7305 (N_7305,N_4607,N_5102);
xnor U7306 (N_7306,N_5016,N_5763);
and U7307 (N_7307,N_5036,N_4702);
or U7308 (N_7308,N_5988,N_5572);
nor U7309 (N_7309,N_4042,N_5542);
nor U7310 (N_7310,N_4195,N_5447);
xnor U7311 (N_7311,N_4781,N_4560);
or U7312 (N_7312,N_4735,N_4085);
nor U7313 (N_7313,N_4141,N_4439);
nand U7314 (N_7314,N_4985,N_4101);
nor U7315 (N_7315,N_5140,N_5082);
nand U7316 (N_7316,N_4611,N_4648);
and U7317 (N_7317,N_4959,N_5792);
or U7318 (N_7318,N_4010,N_4023);
or U7319 (N_7319,N_4922,N_4049);
or U7320 (N_7320,N_5656,N_4599);
nor U7321 (N_7321,N_5258,N_5145);
xnor U7322 (N_7322,N_4448,N_4962);
and U7323 (N_7323,N_4653,N_4104);
or U7324 (N_7324,N_4765,N_5781);
nor U7325 (N_7325,N_5399,N_4699);
xnor U7326 (N_7326,N_4791,N_4877);
nor U7327 (N_7327,N_5819,N_5206);
nor U7328 (N_7328,N_4356,N_5115);
or U7329 (N_7329,N_5479,N_5418);
and U7330 (N_7330,N_4675,N_4900);
or U7331 (N_7331,N_4836,N_4827);
or U7332 (N_7332,N_4171,N_4964);
and U7333 (N_7333,N_4741,N_5912);
nor U7334 (N_7334,N_4254,N_4657);
nand U7335 (N_7335,N_4804,N_5864);
or U7336 (N_7336,N_4600,N_5026);
nor U7337 (N_7337,N_5571,N_5556);
and U7338 (N_7338,N_4378,N_4678);
nor U7339 (N_7339,N_4424,N_5259);
nand U7340 (N_7340,N_5800,N_4775);
xnor U7341 (N_7341,N_4300,N_4698);
and U7342 (N_7342,N_5723,N_5580);
xnor U7343 (N_7343,N_5229,N_4705);
nor U7344 (N_7344,N_5834,N_4016);
xnor U7345 (N_7345,N_4188,N_5957);
and U7346 (N_7346,N_4838,N_5624);
xor U7347 (N_7347,N_4497,N_5451);
and U7348 (N_7348,N_4850,N_4333);
nand U7349 (N_7349,N_4234,N_4156);
nand U7350 (N_7350,N_5798,N_5805);
nor U7351 (N_7351,N_4816,N_5546);
or U7352 (N_7352,N_5325,N_4031);
or U7353 (N_7353,N_5370,N_5988);
nor U7354 (N_7354,N_4383,N_5413);
xor U7355 (N_7355,N_5541,N_5505);
xnor U7356 (N_7356,N_4100,N_4226);
and U7357 (N_7357,N_4802,N_4446);
and U7358 (N_7358,N_5261,N_5314);
nor U7359 (N_7359,N_4454,N_4559);
nor U7360 (N_7360,N_4216,N_5493);
and U7361 (N_7361,N_5014,N_5346);
nor U7362 (N_7362,N_5848,N_5210);
or U7363 (N_7363,N_5295,N_5678);
and U7364 (N_7364,N_5802,N_4020);
nor U7365 (N_7365,N_4316,N_4896);
nand U7366 (N_7366,N_5889,N_4208);
or U7367 (N_7367,N_5619,N_5833);
or U7368 (N_7368,N_5059,N_4019);
nor U7369 (N_7369,N_5844,N_5196);
nand U7370 (N_7370,N_5554,N_4725);
xnor U7371 (N_7371,N_5644,N_5939);
xor U7372 (N_7372,N_5565,N_5915);
nor U7373 (N_7373,N_4974,N_4832);
xor U7374 (N_7374,N_4162,N_5735);
nor U7375 (N_7375,N_4866,N_4605);
nand U7376 (N_7376,N_4350,N_5909);
nor U7377 (N_7377,N_5955,N_5249);
nand U7378 (N_7378,N_5774,N_5487);
and U7379 (N_7379,N_4304,N_5361);
and U7380 (N_7380,N_4694,N_4087);
or U7381 (N_7381,N_4864,N_5623);
and U7382 (N_7382,N_5997,N_4909);
and U7383 (N_7383,N_5784,N_4012);
nor U7384 (N_7384,N_5431,N_4814);
xor U7385 (N_7385,N_4119,N_4255);
xnor U7386 (N_7386,N_4564,N_4291);
and U7387 (N_7387,N_5259,N_5734);
nor U7388 (N_7388,N_5218,N_5704);
nor U7389 (N_7389,N_5194,N_4045);
or U7390 (N_7390,N_4391,N_5704);
xnor U7391 (N_7391,N_5789,N_5722);
nor U7392 (N_7392,N_4729,N_4345);
and U7393 (N_7393,N_4461,N_5944);
or U7394 (N_7394,N_4755,N_5649);
xor U7395 (N_7395,N_4659,N_4446);
or U7396 (N_7396,N_5322,N_4610);
nor U7397 (N_7397,N_4207,N_4008);
nor U7398 (N_7398,N_4940,N_4275);
xor U7399 (N_7399,N_5710,N_5807);
nor U7400 (N_7400,N_5184,N_5629);
xnor U7401 (N_7401,N_4880,N_4334);
nor U7402 (N_7402,N_5722,N_5452);
and U7403 (N_7403,N_5228,N_4377);
xnor U7404 (N_7404,N_4030,N_5535);
nand U7405 (N_7405,N_5712,N_5417);
xnor U7406 (N_7406,N_4034,N_4487);
nor U7407 (N_7407,N_5455,N_4663);
nor U7408 (N_7408,N_4319,N_5231);
and U7409 (N_7409,N_4198,N_5912);
nor U7410 (N_7410,N_5888,N_5970);
and U7411 (N_7411,N_5087,N_5237);
and U7412 (N_7412,N_5350,N_4925);
or U7413 (N_7413,N_4835,N_4026);
and U7414 (N_7414,N_5255,N_4155);
and U7415 (N_7415,N_5364,N_4318);
xnor U7416 (N_7416,N_4579,N_5878);
nand U7417 (N_7417,N_4691,N_4518);
nand U7418 (N_7418,N_5548,N_4229);
and U7419 (N_7419,N_5973,N_5693);
nor U7420 (N_7420,N_5828,N_5585);
nor U7421 (N_7421,N_4081,N_5377);
and U7422 (N_7422,N_5273,N_4278);
xnor U7423 (N_7423,N_4030,N_5185);
and U7424 (N_7424,N_5204,N_4291);
or U7425 (N_7425,N_4329,N_5614);
and U7426 (N_7426,N_4576,N_5891);
or U7427 (N_7427,N_4221,N_5899);
and U7428 (N_7428,N_5597,N_4485);
nand U7429 (N_7429,N_5919,N_4619);
and U7430 (N_7430,N_4780,N_5921);
nand U7431 (N_7431,N_4438,N_4933);
nand U7432 (N_7432,N_5868,N_5150);
xnor U7433 (N_7433,N_5992,N_4554);
nor U7434 (N_7434,N_4193,N_5675);
nor U7435 (N_7435,N_4183,N_5718);
nor U7436 (N_7436,N_4875,N_4656);
nor U7437 (N_7437,N_5622,N_5830);
nand U7438 (N_7438,N_4451,N_4482);
or U7439 (N_7439,N_4935,N_4640);
and U7440 (N_7440,N_4292,N_5716);
xor U7441 (N_7441,N_4350,N_5870);
nor U7442 (N_7442,N_4655,N_5310);
xor U7443 (N_7443,N_4537,N_4284);
nor U7444 (N_7444,N_5306,N_4815);
and U7445 (N_7445,N_4231,N_5696);
nand U7446 (N_7446,N_4154,N_4574);
xor U7447 (N_7447,N_4779,N_5456);
or U7448 (N_7448,N_4475,N_4425);
nor U7449 (N_7449,N_4280,N_5160);
or U7450 (N_7450,N_4980,N_5266);
or U7451 (N_7451,N_4573,N_4228);
and U7452 (N_7452,N_4314,N_4313);
nor U7453 (N_7453,N_4890,N_4682);
nor U7454 (N_7454,N_5471,N_4731);
xor U7455 (N_7455,N_4670,N_4768);
or U7456 (N_7456,N_5823,N_4316);
and U7457 (N_7457,N_5479,N_5719);
nand U7458 (N_7458,N_4822,N_5460);
nand U7459 (N_7459,N_5350,N_5689);
xor U7460 (N_7460,N_4029,N_4542);
and U7461 (N_7461,N_5204,N_4925);
and U7462 (N_7462,N_4382,N_4025);
nand U7463 (N_7463,N_4288,N_4151);
nand U7464 (N_7464,N_4473,N_5574);
and U7465 (N_7465,N_5042,N_5061);
and U7466 (N_7466,N_4982,N_5380);
xnor U7467 (N_7467,N_5620,N_5507);
and U7468 (N_7468,N_4894,N_4335);
nand U7469 (N_7469,N_4870,N_5671);
or U7470 (N_7470,N_4349,N_4578);
or U7471 (N_7471,N_4548,N_5748);
xnor U7472 (N_7472,N_4034,N_4726);
xor U7473 (N_7473,N_4924,N_5192);
and U7474 (N_7474,N_4941,N_5788);
or U7475 (N_7475,N_4917,N_4278);
xnor U7476 (N_7476,N_5888,N_4276);
or U7477 (N_7477,N_4808,N_4249);
nor U7478 (N_7478,N_4729,N_5890);
or U7479 (N_7479,N_5442,N_5395);
or U7480 (N_7480,N_4670,N_4883);
xor U7481 (N_7481,N_5745,N_4503);
nand U7482 (N_7482,N_4717,N_4979);
nor U7483 (N_7483,N_4238,N_5344);
or U7484 (N_7484,N_5960,N_5979);
and U7485 (N_7485,N_5625,N_4135);
or U7486 (N_7486,N_5534,N_4776);
nor U7487 (N_7487,N_5792,N_5103);
nand U7488 (N_7488,N_5077,N_5854);
or U7489 (N_7489,N_5565,N_4787);
or U7490 (N_7490,N_4096,N_5706);
nor U7491 (N_7491,N_4402,N_5250);
and U7492 (N_7492,N_5517,N_4726);
xor U7493 (N_7493,N_4122,N_5174);
and U7494 (N_7494,N_5651,N_4758);
nand U7495 (N_7495,N_4627,N_5560);
xor U7496 (N_7496,N_4581,N_4420);
and U7497 (N_7497,N_4822,N_5349);
nand U7498 (N_7498,N_4124,N_4598);
nor U7499 (N_7499,N_5823,N_4541);
nor U7500 (N_7500,N_4200,N_5547);
xor U7501 (N_7501,N_5500,N_4505);
or U7502 (N_7502,N_4216,N_5435);
or U7503 (N_7503,N_5051,N_5728);
xnor U7504 (N_7504,N_4359,N_4203);
xor U7505 (N_7505,N_4505,N_5456);
or U7506 (N_7506,N_5548,N_5375);
and U7507 (N_7507,N_4314,N_5044);
and U7508 (N_7508,N_5432,N_5443);
xnor U7509 (N_7509,N_4990,N_4228);
or U7510 (N_7510,N_5769,N_4876);
nor U7511 (N_7511,N_4300,N_5366);
nor U7512 (N_7512,N_4972,N_4112);
and U7513 (N_7513,N_5530,N_5578);
or U7514 (N_7514,N_4400,N_5444);
and U7515 (N_7515,N_4078,N_4960);
nor U7516 (N_7516,N_4628,N_4172);
and U7517 (N_7517,N_4876,N_4627);
nand U7518 (N_7518,N_4926,N_5856);
or U7519 (N_7519,N_4912,N_5800);
nand U7520 (N_7520,N_4971,N_5993);
xor U7521 (N_7521,N_5615,N_5624);
and U7522 (N_7522,N_4044,N_5857);
nand U7523 (N_7523,N_5704,N_5031);
nand U7524 (N_7524,N_5296,N_4117);
or U7525 (N_7525,N_5858,N_5460);
nor U7526 (N_7526,N_5789,N_5725);
nor U7527 (N_7527,N_5886,N_4374);
nor U7528 (N_7528,N_5218,N_4935);
nor U7529 (N_7529,N_4402,N_4930);
nand U7530 (N_7530,N_4935,N_4880);
xor U7531 (N_7531,N_4943,N_5266);
or U7532 (N_7532,N_5241,N_4281);
nor U7533 (N_7533,N_5568,N_5919);
nand U7534 (N_7534,N_5524,N_4065);
xnor U7535 (N_7535,N_4055,N_4033);
or U7536 (N_7536,N_4703,N_4619);
nand U7537 (N_7537,N_5130,N_4452);
and U7538 (N_7538,N_4895,N_5780);
or U7539 (N_7539,N_5505,N_4896);
and U7540 (N_7540,N_5364,N_4371);
nor U7541 (N_7541,N_5361,N_4760);
xnor U7542 (N_7542,N_5504,N_5291);
xnor U7543 (N_7543,N_4081,N_4171);
xnor U7544 (N_7544,N_5758,N_4279);
and U7545 (N_7545,N_5070,N_4612);
and U7546 (N_7546,N_4449,N_4471);
xor U7547 (N_7547,N_5321,N_4923);
or U7548 (N_7548,N_5897,N_4296);
nor U7549 (N_7549,N_4520,N_4268);
or U7550 (N_7550,N_5600,N_5753);
and U7551 (N_7551,N_5168,N_5741);
or U7552 (N_7552,N_4652,N_4575);
nor U7553 (N_7553,N_4400,N_5727);
and U7554 (N_7554,N_5612,N_4029);
nor U7555 (N_7555,N_4027,N_5217);
nand U7556 (N_7556,N_5821,N_5040);
nand U7557 (N_7557,N_4054,N_4152);
nand U7558 (N_7558,N_4297,N_5560);
and U7559 (N_7559,N_5601,N_5929);
xor U7560 (N_7560,N_4150,N_5102);
or U7561 (N_7561,N_4334,N_5786);
nor U7562 (N_7562,N_5427,N_4171);
or U7563 (N_7563,N_5414,N_5947);
xor U7564 (N_7564,N_4219,N_5281);
and U7565 (N_7565,N_5074,N_5653);
xor U7566 (N_7566,N_5275,N_5459);
and U7567 (N_7567,N_5840,N_4189);
nor U7568 (N_7568,N_4677,N_4498);
nor U7569 (N_7569,N_5326,N_5564);
and U7570 (N_7570,N_4209,N_4535);
nand U7571 (N_7571,N_4867,N_4843);
or U7572 (N_7572,N_4022,N_5224);
nand U7573 (N_7573,N_4460,N_4624);
xnor U7574 (N_7574,N_4027,N_4619);
nor U7575 (N_7575,N_5566,N_5181);
nor U7576 (N_7576,N_5241,N_4971);
xnor U7577 (N_7577,N_5507,N_4966);
xnor U7578 (N_7578,N_4166,N_4876);
and U7579 (N_7579,N_4605,N_5782);
or U7580 (N_7580,N_5101,N_4580);
nor U7581 (N_7581,N_4312,N_5897);
and U7582 (N_7582,N_4936,N_5777);
and U7583 (N_7583,N_4033,N_5134);
xnor U7584 (N_7584,N_4935,N_5524);
nand U7585 (N_7585,N_5875,N_4498);
or U7586 (N_7586,N_5096,N_5300);
nand U7587 (N_7587,N_5031,N_4470);
xnor U7588 (N_7588,N_5303,N_5675);
and U7589 (N_7589,N_5118,N_5424);
and U7590 (N_7590,N_5054,N_4885);
and U7591 (N_7591,N_4214,N_5654);
or U7592 (N_7592,N_4846,N_4168);
nor U7593 (N_7593,N_5371,N_5475);
and U7594 (N_7594,N_5852,N_4503);
nor U7595 (N_7595,N_4708,N_4339);
nand U7596 (N_7596,N_5301,N_5779);
nand U7597 (N_7597,N_4293,N_5656);
and U7598 (N_7598,N_4958,N_4901);
xnor U7599 (N_7599,N_4168,N_4357);
or U7600 (N_7600,N_4902,N_5620);
or U7601 (N_7601,N_4894,N_5645);
nor U7602 (N_7602,N_5100,N_5059);
or U7603 (N_7603,N_4396,N_5034);
nor U7604 (N_7604,N_4408,N_4363);
nand U7605 (N_7605,N_4477,N_5506);
nand U7606 (N_7606,N_5294,N_5382);
xnor U7607 (N_7607,N_4018,N_4035);
xnor U7608 (N_7608,N_4463,N_5899);
nor U7609 (N_7609,N_5370,N_5744);
or U7610 (N_7610,N_4692,N_5911);
nand U7611 (N_7611,N_5290,N_5383);
nor U7612 (N_7612,N_4678,N_4962);
or U7613 (N_7613,N_5433,N_5693);
or U7614 (N_7614,N_4888,N_4347);
or U7615 (N_7615,N_5197,N_4934);
or U7616 (N_7616,N_5926,N_5016);
and U7617 (N_7617,N_4864,N_5248);
nor U7618 (N_7618,N_4298,N_5950);
and U7619 (N_7619,N_4664,N_5372);
nand U7620 (N_7620,N_5935,N_4172);
and U7621 (N_7621,N_5450,N_5383);
and U7622 (N_7622,N_5912,N_5385);
and U7623 (N_7623,N_4549,N_4865);
or U7624 (N_7624,N_4080,N_5490);
xnor U7625 (N_7625,N_5526,N_5633);
nor U7626 (N_7626,N_5189,N_5435);
or U7627 (N_7627,N_5403,N_5544);
xnor U7628 (N_7628,N_4607,N_5413);
nand U7629 (N_7629,N_5229,N_4934);
or U7630 (N_7630,N_5795,N_4521);
nand U7631 (N_7631,N_5186,N_4211);
or U7632 (N_7632,N_4753,N_4465);
or U7633 (N_7633,N_5726,N_4370);
or U7634 (N_7634,N_5426,N_5059);
and U7635 (N_7635,N_4346,N_5542);
and U7636 (N_7636,N_4998,N_5580);
nor U7637 (N_7637,N_4411,N_5771);
or U7638 (N_7638,N_5998,N_4666);
nor U7639 (N_7639,N_5292,N_4898);
and U7640 (N_7640,N_4550,N_5747);
and U7641 (N_7641,N_4316,N_4584);
nand U7642 (N_7642,N_4174,N_5462);
nand U7643 (N_7643,N_5828,N_5343);
xor U7644 (N_7644,N_5985,N_5395);
nor U7645 (N_7645,N_4417,N_5243);
and U7646 (N_7646,N_4246,N_4295);
or U7647 (N_7647,N_5990,N_4624);
or U7648 (N_7648,N_5712,N_5515);
and U7649 (N_7649,N_5845,N_5241);
or U7650 (N_7650,N_4165,N_4943);
and U7651 (N_7651,N_5857,N_5747);
xor U7652 (N_7652,N_4749,N_5625);
and U7653 (N_7653,N_4366,N_4499);
and U7654 (N_7654,N_5478,N_5282);
nor U7655 (N_7655,N_4360,N_5769);
xor U7656 (N_7656,N_5523,N_4640);
nor U7657 (N_7657,N_4992,N_5938);
or U7658 (N_7658,N_4347,N_5956);
and U7659 (N_7659,N_4900,N_5013);
nand U7660 (N_7660,N_4474,N_5722);
or U7661 (N_7661,N_4952,N_4229);
and U7662 (N_7662,N_4119,N_4065);
and U7663 (N_7663,N_5698,N_4985);
xnor U7664 (N_7664,N_4596,N_4841);
nor U7665 (N_7665,N_5311,N_4204);
or U7666 (N_7666,N_4205,N_4965);
nor U7667 (N_7667,N_4487,N_4209);
xor U7668 (N_7668,N_5105,N_5451);
and U7669 (N_7669,N_5485,N_4779);
or U7670 (N_7670,N_4615,N_4733);
xnor U7671 (N_7671,N_5775,N_5889);
nand U7672 (N_7672,N_5417,N_4792);
nand U7673 (N_7673,N_5155,N_4690);
nand U7674 (N_7674,N_5238,N_4232);
and U7675 (N_7675,N_5555,N_4710);
nor U7676 (N_7676,N_5696,N_4911);
or U7677 (N_7677,N_4234,N_4184);
nor U7678 (N_7678,N_4058,N_5908);
xor U7679 (N_7679,N_5219,N_4508);
and U7680 (N_7680,N_5795,N_4768);
xnor U7681 (N_7681,N_5338,N_5285);
and U7682 (N_7682,N_5407,N_5045);
nand U7683 (N_7683,N_5788,N_4318);
nor U7684 (N_7684,N_5655,N_5350);
and U7685 (N_7685,N_5391,N_4883);
xor U7686 (N_7686,N_5260,N_5873);
and U7687 (N_7687,N_4572,N_4584);
nor U7688 (N_7688,N_4375,N_5072);
nand U7689 (N_7689,N_5538,N_4747);
nand U7690 (N_7690,N_4025,N_5892);
nor U7691 (N_7691,N_5557,N_4158);
or U7692 (N_7692,N_4386,N_5933);
nor U7693 (N_7693,N_4666,N_5922);
nand U7694 (N_7694,N_4672,N_5540);
nand U7695 (N_7695,N_4427,N_4673);
and U7696 (N_7696,N_4515,N_5254);
nand U7697 (N_7697,N_5460,N_4313);
nand U7698 (N_7698,N_5463,N_5692);
and U7699 (N_7699,N_4263,N_5545);
nor U7700 (N_7700,N_5303,N_5348);
or U7701 (N_7701,N_4783,N_4913);
xor U7702 (N_7702,N_4574,N_5528);
and U7703 (N_7703,N_5675,N_5264);
nor U7704 (N_7704,N_5937,N_4791);
or U7705 (N_7705,N_4382,N_5627);
nand U7706 (N_7706,N_4429,N_4305);
and U7707 (N_7707,N_4138,N_4263);
nor U7708 (N_7708,N_5313,N_5247);
xnor U7709 (N_7709,N_4767,N_5334);
nor U7710 (N_7710,N_5145,N_4899);
nand U7711 (N_7711,N_4608,N_4136);
or U7712 (N_7712,N_4610,N_4233);
nor U7713 (N_7713,N_4506,N_5506);
and U7714 (N_7714,N_5733,N_5527);
and U7715 (N_7715,N_4722,N_4217);
nor U7716 (N_7716,N_4342,N_4205);
nand U7717 (N_7717,N_4386,N_4438);
nand U7718 (N_7718,N_5538,N_5987);
nor U7719 (N_7719,N_4963,N_4892);
nand U7720 (N_7720,N_5976,N_5598);
and U7721 (N_7721,N_5291,N_5852);
nor U7722 (N_7722,N_5113,N_5105);
nor U7723 (N_7723,N_5538,N_4191);
nand U7724 (N_7724,N_4244,N_4522);
nor U7725 (N_7725,N_4334,N_4250);
or U7726 (N_7726,N_4290,N_5551);
and U7727 (N_7727,N_4353,N_4681);
and U7728 (N_7728,N_5000,N_5481);
nor U7729 (N_7729,N_4979,N_5922);
nand U7730 (N_7730,N_4435,N_5747);
xor U7731 (N_7731,N_4376,N_5614);
and U7732 (N_7732,N_5120,N_5622);
xnor U7733 (N_7733,N_5485,N_4581);
xnor U7734 (N_7734,N_5414,N_4145);
nand U7735 (N_7735,N_4255,N_4071);
nor U7736 (N_7736,N_5061,N_5052);
and U7737 (N_7737,N_4821,N_5303);
xnor U7738 (N_7738,N_4243,N_5407);
xor U7739 (N_7739,N_4538,N_5492);
nand U7740 (N_7740,N_4495,N_5065);
xor U7741 (N_7741,N_4413,N_5737);
or U7742 (N_7742,N_5243,N_5393);
nor U7743 (N_7743,N_5491,N_4162);
nor U7744 (N_7744,N_5278,N_5722);
nand U7745 (N_7745,N_5400,N_5245);
xor U7746 (N_7746,N_5068,N_5064);
nand U7747 (N_7747,N_5592,N_5466);
or U7748 (N_7748,N_5976,N_5702);
nor U7749 (N_7749,N_5374,N_5560);
nor U7750 (N_7750,N_5934,N_4825);
or U7751 (N_7751,N_5340,N_5914);
nor U7752 (N_7752,N_4117,N_4712);
or U7753 (N_7753,N_5305,N_4895);
and U7754 (N_7754,N_4147,N_5520);
nor U7755 (N_7755,N_4665,N_4459);
nor U7756 (N_7756,N_5087,N_4426);
and U7757 (N_7757,N_5473,N_5046);
nor U7758 (N_7758,N_4144,N_5728);
or U7759 (N_7759,N_4084,N_4915);
or U7760 (N_7760,N_4751,N_4336);
nor U7761 (N_7761,N_5036,N_4939);
xnor U7762 (N_7762,N_4304,N_5315);
nand U7763 (N_7763,N_5733,N_5397);
nand U7764 (N_7764,N_5583,N_5336);
and U7765 (N_7765,N_4544,N_5883);
nand U7766 (N_7766,N_4831,N_4039);
nor U7767 (N_7767,N_4304,N_5014);
or U7768 (N_7768,N_4632,N_5308);
or U7769 (N_7769,N_5796,N_5093);
nand U7770 (N_7770,N_4019,N_5381);
nand U7771 (N_7771,N_5979,N_4225);
or U7772 (N_7772,N_5021,N_4871);
nand U7773 (N_7773,N_5601,N_4596);
nor U7774 (N_7774,N_4137,N_5461);
nand U7775 (N_7775,N_5886,N_4878);
nor U7776 (N_7776,N_4612,N_5502);
nor U7777 (N_7777,N_4817,N_4163);
nand U7778 (N_7778,N_4990,N_4584);
or U7779 (N_7779,N_4946,N_5459);
xor U7780 (N_7780,N_5543,N_4309);
nor U7781 (N_7781,N_4302,N_4039);
xnor U7782 (N_7782,N_5989,N_4687);
and U7783 (N_7783,N_5796,N_4891);
nor U7784 (N_7784,N_5808,N_4868);
and U7785 (N_7785,N_5835,N_5154);
xnor U7786 (N_7786,N_4696,N_4347);
xnor U7787 (N_7787,N_4109,N_5041);
and U7788 (N_7788,N_5184,N_4275);
or U7789 (N_7789,N_4945,N_5373);
and U7790 (N_7790,N_5699,N_5561);
nor U7791 (N_7791,N_4262,N_4189);
xor U7792 (N_7792,N_5379,N_4761);
nor U7793 (N_7793,N_5125,N_5482);
nor U7794 (N_7794,N_4912,N_4538);
nand U7795 (N_7795,N_5404,N_5750);
nand U7796 (N_7796,N_5898,N_5053);
xor U7797 (N_7797,N_4383,N_4042);
nand U7798 (N_7798,N_4493,N_5135);
xnor U7799 (N_7799,N_5630,N_4543);
nor U7800 (N_7800,N_4496,N_4280);
or U7801 (N_7801,N_5684,N_4988);
and U7802 (N_7802,N_5647,N_4603);
nand U7803 (N_7803,N_5934,N_4228);
xor U7804 (N_7804,N_4794,N_5184);
nand U7805 (N_7805,N_4858,N_4027);
xor U7806 (N_7806,N_4560,N_4046);
nand U7807 (N_7807,N_5448,N_4819);
xnor U7808 (N_7808,N_5508,N_5862);
nand U7809 (N_7809,N_4819,N_5475);
nor U7810 (N_7810,N_4135,N_4917);
nand U7811 (N_7811,N_5545,N_4340);
or U7812 (N_7812,N_5236,N_4283);
nor U7813 (N_7813,N_5112,N_4991);
nand U7814 (N_7814,N_5151,N_5208);
xnor U7815 (N_7815,N_5400,N_4931);
nand U7816 (N_7816,N_4481,N_5173);
xnor U7817 (N_7817,N_5459,N_5592);
or U7818 (N_7818,N_4971,N_5202);
and U7819 (N_7819,N_5877,N_5146);
xnor U7820 (N_7820,N_5078,N_4395);
xor U7821 (N_7821,N_4175,N_4746);
and U7822 (N_7822,N_4842,N_5259);
nand U7823 (N_7823,N_5343,N_5283);
or U7824 (N_7824,N_5031,N_4822);
xor U7825 (N_7825,N_5705,N_5818);
or U7826 (N_7826,N_4138,N_5430);
nand U7827 (N_7827,N_4373,N_5716);
xor U7828 (N_7828,N_4904,N_5951);
nand U7829 (N_7829,N_5389,N_5193);
and U7830 (N_7830,N_4772,N_4754);
or U7831 (N_7831,N_5524,N_5274);
nand U7832 (N_7832,N_4693,N_5372);
xor U7833 (N_7833,N_4748,N_4770);
or U7834 (N_7834,N_5841,N_4116);
xnor U7835 (N_7835,N_5192,N_5327);
xnor U7836 (N_7836,N_4964,N_5107);
nand U7837 (N_7837,N_4685,N_4700);
and U7838 (N_7838,N_4422,N_4724);
nor U7839 (N_7839,N_5866,N_5167);
nand U7840 (N_7840,N_5718,N_5166);
nor U7841 (N_7841,N_5636,N_5226);
nand U7842 (N_7842,N_5170,N_4429);
nor U7843 (N_7843,N_4157,N_5856);
xnor U7844 (N_7844,N_4195,N_5477);
and U7845 (N_7845,N_4296,N_4294);
or U7846 (N_7846,N_4485,N_5856);
nor U7847 (N_7847,N_4631,N_4644);
nor U7848 (N_7848,N_4387,N_5049);
and U7849 (N_7849,N_5525,N_5135);
nor U7850 (N_7850,N_5319,N_4200);
xnor U7851 (N_7851,N_5999,N_4317);
xnor U7852 (N_7852,N_4400,N_5858);
and U7853 (N_7853,N_4907,N_5833);
xor U7854 (N_7854,N_4491,N_5433);
nand U7855 (N_7855,N_4009,N_4120);
and U7856 (N_7856,N_4775,N_5825);
nand U7857 (N_7857,N_4791,N_4131);
and U7858 (N_7858,N_5464,N_5904);
and U7859 (N_7859,N_4116,N_4398);
xnor U7860 (N_7860,N_5226,N_4190);
xnor U7861 (N_7861,N_4311,N_5656);
and U7862 (N_7862,N_4369,N_5982);
and U7863 (N_7863,N_4528,N_4848);
nand U7864 (N_7864,N_4841,N_5262);
nand U7865 (N_7865,N_5054,N_5523);
and U7866 (N_7866,N_5845,N_5163);
xor U7867 (N_7867,N_4583,N_4561);
nand U7868 (N_7868,N_5241,N_5248);
xor U7869 (N_7869,N_4198,N_5459);
xnor U7870 (N_7870,N_5234,N_4190);
or U7871 (N_7871,N_5968,N_4354);
and U7872 (N_7872,N_5020,N_4537);
nor U7873 (N_7873,N_4119,N_4740);
and U7874 (N_7874,N_5617,N_4179);
nand U7875 (N_7875,N_4817,N_4800);
xor U7876 (N_7876,N_5586,N_5025);
xnor U7877 (N_7877,N_5518,N_5019);
nor U7878 (N_7878,N_5613,N_4521);
and U7879 (N_7879,N_5820,N_4164);
or U7880 (N_7880,N_4759,N_4454);
or U7881 (N_7881,N_5408,N_4949);
or U7882 (N_7882,N_4238,N_4955);
and U7883 (N_7883,N_4854,N_4991);
or U7884 (N_7884,N_4282,N_5090);
nand U7885 (N_7885,N_5881,N_4414);
nand U7886 (N_7886,N_4134,N_5369);
nor U7887 (N_7887,N_4399,N_4091);
nand U7888 (N_7888,N_4963,N_5079);
and U7889 (N_7889,N_5270,N_5566);
and U7890 (N_7890,N_5976,N_5763);
or U7891 (N_7891,N_5183,N_4059);
nor U7892 (N_7892,N_5207,N_4831);
xor U7893 (N_7893,N_5975,N_4484);
nand U7894 (N_7894,N_4896,N_5924);
and U7895 (N_7895,N_5090,N_4353);
and U7896 (N_7896,N_5590,N_4049);
xnor U7897 (N_7897,N_4711,N_4741);
xor U7898 (N_7898,N_4926,N_4621);
nor U7899 (N_7899,N_4362,N_5220);
nor U7900 (N_7900,N_4438,N_4840);
and U7901 (N_7901,N_4465,N_5015);
xor U7902 (N_7902,N_4885,N_5796);
xnor U7903 (N_7903,N_5148,N_5780);
nand U7904 (N_7904,N_4874,N_5334);
or U7905 (N_7905,N_5617,N_4903);
or U7906 (N_7906,N_5263,N_5042);
nand U7907 (N_7907,N_4048,N_4011);
xor U7908 (N_7908,N_4310,N_5072);
xor U7909 (N_7909,N_4933,N_5165);
nand U7910 (N_7910,N_4800,N_4706);
nor U7911 (N_7911,N_4651,N_5956);
nand U7912 (N_7912,N_4698,N_5303);
and U7913 (N_7913,N_4332,N_4230);
or U7914 (N_7914,N_5685,N_5736);
and U7915 (N_7915,N_4571,N_5944);
xnor U7916 (N_7916,N_5177,N_4331);
and U7917 (N_7917,N_5021,N_4021);
xor U7918 (N_7918,N_4337,N_5277);
nand U7919 (N_7919,N_4757,N_4348);
nor U7920 (N_7920,N_4840,N_5185);
and U7921 (N_7921,N_5998,N_5160);
nand U7922 (N_7922,N_4868,N_5713);
and U7923 (N_7923,N_4492,N_5188);
nand U7924 (N_7924,N_5515,N_5408);
xor U7925 (N_7925,N_4208,N_5719);
or U7926 (N_7926,N_4779,N_4276);
nor U7927 (N_7927,N_5285,N_4265);
xor U7928 (N_7928,N_5241,N_5462);
xnor U7929 (N_7929,N_5247,N_5249);
or U7930 (N_7930,N_5115,N_5810);
xnor U7931 (N_7931,N_5231,N_4198);
nor U7932 (N_7932,N_4650,N_5010);
nand U7933 (N_7933,N_5598,N_4198);
and U7934 (N_7934,N_5048,N_4931);
or U7935 (N_7935,N_4672,N_5559);
nor U7936 (N_7936,N_5729,N_5857);
nand U7937 (N_7937,N_5051,N_4648);
nor U7938 (N_7938,N_4983,N_5832);
or U7939 (N_7939,N_5425,N_4239);
xor U7940 (N_7940,N_5763,N_4741);
xor U7941 (N_7941,N_4099,N_4837);
nand U7942 (N_7942,N_4890,N_5252);
nor U7943 (N_7943,N_5880,N_4535);
or U7944 (N_7944,N_4236,N_4080);
nor U7945 (N_7945,N_5883,N_4669);
and U7946 (N_7946,N_5726,N_5743);
nor U7947 (N_7947,N_5395,N_5609);
or U7948 (N_7948,N_4072,N_4646);
xnor U7949 (N_7949,N_5643,N_5164);
xnor U7950 (N_7950,N_4295,N_5566);
nand U7951 (N_7951,N_5224,N_5607);
or U7952 (N_7952,N_4577,N_4084);
and U7953 (N_7953,N_4040,N_4696);
xnor U7954 (N_7954,N_5440,N_4079);
nor U7955 (N_7955,N_4699,N_5605);
nand U7956 (N_7956,N_5760,N_5640);
xnor U7957 (N_7957,N_5327,N_4792);
xor U7958 (N_7958,N_4863,N_4039);
or U7959 (N_7959,N_4473,N_4211);
xnor U7960 (N_7960,N_5183,N_4981);
nand U7961 (N_7961,N_5601,N_5798);
nor U7962 (N_7962,N_4040,N_5478);
or U7963 (N_7963,N_5647,N_4517);
and U7964 (N_7964,N_5761,N_4296);
nand U7965 (N_7965,N_4853,N_4653);
xor U7966 (N_7966,N_5834,N_4395);
nor U7967 (N_7967,N_4625,N_5045);
xor U7968 (N_7968,N_5990,N_4514);
and U7969 (N_7969,N_5811,N_4578);
nand U7970 (N_7970,N_4332,N_5732);
nand U7971 (N_7971,N_5678,N_4513);
xnor U7972 (N_7972,N_4037,N_5375);
nor U7973 (N_7973,N_5668,N_4227);
or U7974 (N_7974,N_4526,N_5379);
xnor U7975 (N_7975,N_5575,N_4508);
or U7976 (N_7976,N_4912,N_4280);
xor U7977 (N_7977,N_4023,N_4479);
and U7978 (N_7978,N_4641,N_5382);
or U7979 (N_7979,N_5256,N_5416);
or U7980 (N_7980,N_5592,N_4854);
or U7981 (N_7981,N_5985,N_5764);
nand U7982 (N_7982,N_4652,N_4647);
or U7983 (N_7983,N_4302,N_5683);
xnor U7984 (N_7984,N_5083,N_5546);
xnor U7985 (N_7985,N_4063,N_5068);
and U7986 (N_7986,N_4736,N_4333);
xnor U7987 (N_7987,N_5179,N_5042);
nor U7988 (N_7988,N_4499,N_4275);
nand U7989 (N_7989,N_5918,N_5870);
and U7990 (N_7990,N_4129,N_5440);
and U7991 (N_7991,N_5058,N_5339);
xor U7992 (N_7992,N_4291,N_4279);
or U7993 (N_7993,N_5881,N_5708);
or U7994 (N_7994,N_5364,N_4277);
or U7995 (N_7995,N_4697,N_4328);
nand U7996 (N_7996,N_5433,N_5138);
nor U7997 (N_7997,N_4770,N_4662);
nand U7998 (N_7998,N_4842,N_5473);
nor U7999 (N_7999,N_5625,N_5066);
and U8000 (N_8000,N_7893,N_7798);
and U8001 (N_8001,N_6655,N_7775);
xnor U8002 (N_8002,N_6937,N_6789);
or U8003 (N_8003,N_7304,N_6008);
nand U8004 (N_8004,N_6256,N_7297);
xor U8005 (N_8005,N_7565,N_6597);
or U8006 (N_8006,N_7786,N_7275);
nand U8007 (N_8007,N_6067,N_7961);
nor U8008 (N_8008,N_6377,N_6833);
nor U8009 (N_8009,N_7865,N_7403);
nand U8010 (N_8010,N_7020,N_7815);
xor U8011 (N_8011,N_6681,N_7420);
nand U8012 (N_8012,N_6090,N_7144);
nand U8013 (N_8013,N_7399,N_7721);
or U8014 (N_8014,N_7274,N_6138);
xnor U8015 (N_8015,N_7787,N_7758);
or U8016 (N_8016,N_7492,N_7630);
or U8017 (N_8017,N_7282,N_7281);
and U8018 (N_8018,N_6285,N_6701);
nand U8019 (N_8019,N_7043,N_7021);
or U8020 (N_8020,N_6867,N_6944);
xor U8021 (N_8021,N_7889,N_7435);
xnor U8022 (N_8022,N_6425,N_7876);
or U8023 (N_8023,N_7372,N_7169);
and U8024 (N_8024,N_7107,N_6910);
nor U8025 (N_8025,N_6508,N_6325);
nor U8026 (N_8026,N_6875,N_7869);
xnor U8027 (N_8027,N_7591,N_6258);
nor U8028 (N_8028,N_7750,N_6428);
xor U8029 (N_8029,N_7520,N_6427);
nand U8030 (N_8030,N_6912,N_7386);
or U8031 (N_8031,N_7631,N_6190);
or U8032 (N_8032,N_7925,N_6403);
xor U8033 (N_8033,N_6466,N_7133);
nand U8034 (N_8034,N_6668,N_7514);
nor U8035 (N_8035,N_6879,N_6922);
nand U8036 (N_8036,N_7227,N_6758);
nor U8037 (N_8037,N_6218,N_7789);
nand U8038 (N_8038,N_7013,N_7956);
and U8039 (N_8039,N_7725,N_7592);
nand U8040 (N_8040,N_7508,N_7195);
nand U8041 (N_8041,N_6660,N_7734);
and U8042 (N_8042,N_6368,N_6808);
nand U8043 (N_8043,N_6532,N_7858);
nor U8044 (N_8044,N_7945,N_6111);
xnor U8045 (N_8045,N_7821,N_7458);
xnor U8046 (N_8046,N_7023,N_7543);
nor U8047 (N_8047,N_6757,N_6225);
nor U8048 (N_8048,N_6180,N_7946);
or U8049 (N_8049,N_7232,N_7664);
and U8050 (N_8050,N_6239,N_6296);
xnor U8051 (N_8051,N_7042,N_6905);
xor U8052 (N_8052,N_6421,N_6737);
nor U8053 (N_8053,N_7727,N_6783);
or U8054 (N_8054,N_6350,N_6749);
or U8055 (N_8055,N_7763,N_6921);
nor U8056 (N_8056,N_6547,N_6027);
and U8057 (N_8057,N_7368,N_7729);
nand U8058 (N_8058,N_7004,N_7875);
nor U8059 (N_8059,N_7507,N_6306);
nand U8060 (N_8060,N_7394,N_7467);
nor U8061 (N_8061,N_6459,N_6792);
and U8062 (N_8062,N_7566,N_6826);
nand U8063 (N_8063,N_7935,N_6370);
and U8064 (N_8064,N_7730,N_6173);
nor U8065 (N_8065,N_7357,N_6687);
and U8066 (N_8066,N_6301,N_6522);
nor U8067 (N_8067,N_7430,N_6990);
nand U8068 (N_8068,N_6860,N_7857);
nand U8069 (N_8069,N_6623,N_6451);
or U8070 (N_8070,N_7012,N_6162);
and U8071 (N_8071,N_6521,N_7928);
nand U8072 (N_8072,N_7864,N_6886);
nor U8073 (N_8073,N_6513,N_7202);
and U8074 (N_8074,N_7257,N_6223);
and U8075 (N_8075,N_7689,N_6065);
nor U8076 (N_8076,N_7996,N_7222);
xnor U8077 (N_8077,N_6777,N_7438);
nor U8078 (N_8078,N_6514,N_7123);
or U8079 (N_8079,N_6398,N_6518);
nand U8080 (N_8080,N_6346,N_6026);
and U8081 (N_8081,N_6807,N_7207);
or U8082 (N_8082,N_7301,N_7620);
nand U8083 (N_8083,N_6132,N_6135);
or U8084 (N_8084,N_6952,N_6520);
or U8085 (N_8085,N_6836,N_6106);
nor U8086 (N_8086,N_7658,N_6574);
and U8087 (N_8087,N_7999,N_7086);
and U8088 (N_8088,N_6120,N_6298);
or U8089 (N_8089,N_7544,N_7283);
nand U8090 (N_8090,N_6166,N_7124);
xor U8091 (N_8091,N_6692,N_6433);
nand U8092 (N_8092,N_6738,N_6224);
nand U8093 (N_8093,N_7575,N_7453);
xor U8094 (N_8094,N_6900,N_6969);
xor U8095 (N_8095,N_6746,N_6903);
nor U8096 (N_8096,N_7518,N_7509);
xor U8097 (N_8097,N_6482,N_6195);
nand U8098 (N_8098,N_6556,N_6152);
or U8099 (N_8099,N_7940,N_7213);
xnor U8100 (N_8100,N_6449,N_7772);
nor U8101 (N_8101,N_7423,N_6571);
nand U8102 (N_8102,N_7986,N_6811);
and U8103 (N_8103,N_6322,N_6664);
and U8104 (N_8104,N_6230,N_7974);
or U8105 (N_8105,N_6958,N_6842);
nor U8106 (N_8106,N_6240,N_7950);
nand U8107 (N_8107,N_7597,N_7849);
or U8108 (N_8108,N_7173,N_7094);
xnor U8109 (N_8109,N_6321,N_7817);
nor U8110 (N_8110,N_7331,N_6885);
or U8111 (N_8111,N_7995,N_7054);
nand U8112 (N_8112,N_7223,N_6215);
or U8113 (N_8113,N_7446,N_7264);
xor U8114 (N_8114,N_7596,N_6145);
nand U8115 (N_8115,N_6515,N_7644);
and U8116 (N_8116,N_6412,N_6528);
nand U8117 (N_8117,N_7670,N_7036);
nor U8118 (N_8118,N_6628,N_7090);
nor U8119 (N_8119,N_6801,N_7549);
xor U8120 (N_8120,N_6973,N_6440);
or U8121 (N_8121,N_6197,N_7773);
nor U8122 (N_8122,N_7007,N_6585);
nor U8123 (N_8123,N_7879,N_7402);
or U8124 (N_8124,N_7861,N_7745);
or U8125 (N_8125,N_6915,N_7662);
and U8126 (N_8126,N_7258,N_7496);
nand U8127 (N_8127,N_7776,N_7424);
nand U8128 (N_8128,N_6881,N_6609);
nor U8129 (N_8129,N_7663,N_7505);
nand U8130 (N_8130,N_7583,N_6951);
nor U8131 (N_8131,N_7442,N_6624);
nor U8132 (N_8132,N_7330,N_6634);
nor U8133 (N_8133,N_6208,N_7038);
nor U8134 (N_8134,N_7382,N_7343);
nor U8135 (N_8135,N_6025,N_6728);
and U8136 (N_8136,N_6485,N_6610);
or U8137 (N_8137,N_6684,N_6541);
nor U8138 (N_8138,N_6032,N_7434);
and U8139 (N_8139,N_6607,N_7142);
or U8140 (N_8140,N_7308,N_7551);
or U8141 (N_8141,N_6380,N_6534);
or U8142 (N_8142,N_6529,N_7968);
xor U8143 (N_8143,N_6612,N_7694);
or U8144 (N_8144,N_6302,N_6772);
nand U8145 (N_8145,N_7531,N_6114);
xnor U8146 (N_8146,N_7672,N_7163);
nand U8147 (N_8147,N_6775,N_6966);
nand U8148 (N_8148,N_7450,N_6342);
nand U8149 (N_8149,N_7942,N_6865);
nor U8150 (N_8150,N_7955,N_7437);
xor U8151 (N_8151,N_6354,N_7754);
nand U8152 (N_8152,N_7062,N_6901);
or U8153 (N_8153,N_6677,N_7949);
nand U8154 (N_8154,N_7731,N_7418);
or U8155 (N_8155,N_7770,N_7693);
xnor U8156 (N_8156,N_6565,N_7319);
xnor U8157 (N_8157,N_7119,N_7494);
nand U8158 (N_8158,N_7310,N_6938);
nor U8159 (N_8159,N_7610,N_6784);
xnor U8160 (N_8160,N_6095,N_7024);
nor U8161 (N_8161,N_6845,N_7624);
xnor U8162 (N_8162,N_6551,N_7116);
xnor U8163 (N_8163,N_6590,N_7171);
nand U8164 (N_8164,N_6330,N_7084);
nor U8165 (N_8165,N_6712,N_6576);
or U8166 (N_8166,N_7586,N_7973);
nor U8167 (N_8167,N_7681,N_6128);
and U8168 (N_8168,N_7466,N_6533);
nor U8169 (N_8169,N_6066,N_7769);
or U8170 (N_8170,N_6110,N_7860);
nand U8171 (N_8171,N_6748,N_7646);
nor U8172 (N_8172,N_7045,N_6564);
xnor U8173 (N_8173,N_6656,N_7525);
nor U8174 (N_8174,N_7542,N_6072);
nor U8175 (N_8175,N_7335,N_6092);
and U8176 (N_8176,N_6391,N_6467);
or U8177 (N_8177,N_6101,N_7573);
xor U8178 (N_8178,N_6150,N_6275);
xor U8179 (N_8179,N_6667,N_6780);
and U8180 (N_8180,N_7419,N_7130);
and U8181 (N_8181,N_6201,N_6318);
nor U8182 (N_8182,N_7778,N_6484);
and U8183 (N_8183,N_7605,N_7621);
nor U8184 (N_8184,N_7501,N_7848);
and U8185 (N_8185,N_7654,N_6392);
nand U8186 (N_8186,N_7738,N_6048);
and U8187 (N_8187,N_7698,N_7978);
and U8188 (N_8188,N_7276,N_7498);
or U8189 (N_8189,N_7181,N_6381);
nand U8190 (N_8190,N_6844,N_7713);
xor U8191 (N_8191,N_7441,N_6112);
nor U8192 (N_8192,N_7005,N_7221);
and U8193 (N_8193,N_7229,N_6028);
xnor U8194 (N_8194,N_6024,N_7040);
nand U8195 (N_8195,N_6584,N_7648);
nand U8196 (N_8196,N_6434,N_6954);
and U8197 (N_8197,N_6081,N_6091);
nand U8198 (N_8198,N_6539,N_7572);
and U8199 (N_8199,N_6137,N_6323);
and U8200 (N_8200,N_6975,N_7483);
nor U8201 (N_8201,N_6893,N_7568);
nand U8202 (N_8202,N_7922,N_7495);
xnor U8203 (N_8203,N_7818,N_7072);
or U8204 (N_8204,N_6304,N_6261);
or U8205 (N_8205,N_6962,N_6993);
xor U8206 (N_8206,N_7063,N_7188);
xor U8207 (N_8207,N_7360,N_6269);
xnor U8208 (N_8208,N_7647,N_7219);
nor U8209 (N_8209,N_7993,N_6974);
xnor U8210 (N_8210,N_7214,N_6943);
xor U8211 (N_8211,N_6198,N_6897);
xnor U8212 (N_8212,N_6144,N_6653);
nand U8213 (N_8213,N_6248,N_7588);
nand U8214 (N_8214,N_7702,N_7369);
and U8215 (N_8215,N_6579,N_6396);
xnor U8216 (N_8216,N_6499,N_6124);
xnor U8217 (N_8217,N_7975,N_7711);
xnor U8218 (N_8218,N_6160,N_6636);
and U8219 (N_8219,N_6407,N_6070);
and U8220 (N_8220,N_6119,N_7703);
and U8221 (N_8221,N_7203,N_6217);
nand U8222 (N_8222,N_7156,N_7558);
xnor U8223 (N_8223,N_6817,N_6037);
nand U8224 (N_8224,N_6043,N_7839);
and U8225 (N_8225,N_6569,N_7158);
nor U8226 (N_8226,N_7376,N_6439);
or U8227 (N_8227,N_7480,N_6926);
or U8228 (N_8228,N_6108,N_6184);
or U8229 (N_8229,N_7890,N_7010);
xor U8230 (N_8230,N_6593,N_6373);
xnor U8231 (N_8231,N_6383,N_7355);
xnor U8232 (N_8232,N_7895,N_6658);
nand U8233 (N_8233,N_7829,N_6343);
nand U8234 (N_8234,N_6154,N_6333);
xor U8235 (N_8235,N_6729,N_7218);
nand U8236 (N_8236,N_7987,N_6204);
xnor U8237 (N_8237,N_7953,N_7179);
and U8238 (N_8238,N_6464,N_6861);
nand U8239 (N_8239,N_6967,N_7078);
nand U8240 (N_8240,N_7436,N_7557);
xor U8241 (N_8241,N_7649,N_6411);
nand U8242 (N_8242,N_7854,N_7808);
nor U8243 (N_8243,N_6400,N_7510);
and U8244 (N_8244,N_6320,N_7318);
nor U8245 (N_8245,N_6986,N_6290);
nand U8246 (N_8246,N_6683,N_7154);
nand U8247 (N_8247,N_6882,N_7032);
nor U8248 (N_8248,N_7868,N_7425);
xnor U8249 (N_8249,N_7679,N_6442);
and U8250 (N_8250,N_6418,N_7872);
and U8251 (N_8251,N_7992,N_7294);
nand U8252 (N_8252,N_7739,N_7464);
xor U8253 (N_8253,N_7306,N_7245);
or U8254 (N_8254,N_7580,N_7200);
or U8255 (N_8255,N_7055,N_6703);
nor U8256 (N_8256,N_6231,N_7058);
nor U8257 (N_8257,N_6813,N_7115);
nor U8258 (N_8258,N_6776,N_6570);
nand U8259 (N_8259,N_7533,N_6883);
nor U8260 (N_8260,N_6480,N_7487);
nand U8261 (N_8261,N_6531,N_6075);
or U8262 (N_8262,N_6353,N_6468);
nor U8263 (N_8263,N_6644,N_7847);
nand U8264 (N_8264,N_6251,N_7743);
or U8265 (N_8265,N_6507,N_7690);
nor U8266 (N_8266,N_6673,N_7801);
and U8267 (N_8267,N_6390,N_6995);
nor U8268 (N_8268,N_6047,N_7105);
nand U8269 (N_8269,N_6519,N_7131);
and U8270 (N_8270,N_7678,N_6489);
or U8271 (N_8271,N_7779,N_6422);
nand U8272 (N_8272,N_6140,N_6554);
nand U8273 (N_8273,N_6415,N_6730);
or U8274 (N_8274,N_7209,N_6212);
nand U8275 (N_8275,N_7211,N_7337);
nor U8276 (N_8276,N_7065,N_6193);
xor U8277 (N_8277,N_7234,N_6537);
nand U8278 (N_8278,N_6059,N_7717);
xor U8279 (N_8279,N_7326,N_7629);
nor U8280 (N_8280,N_7550,N_6620);
and U8281 (N_8281,N_7046,N_6115);
xor U8282 (N_8282,N_6147,N_7688);
or U8283 (N_8283,N_6525,N_7958);
xor U8284 (N_8284,N_7563,N_6049);
or U8285 (N_8285,N_6006,N_6093);
and U8286 (N_8286,N_7175,N_7250);
and U8287 (N_8287,N_7008,N_6751);
and U8288 (N_8288,N_7609,N_6245);
and U8289 (N_8289,N_7692,N_6698);
nor U8290 (N_8290,N_6676,N_6206);
xor U8291 (N_8291,N_6852,N_7059);
nand U8292 (N_8292,N_6778,N_7351);
nor U8293 (N_8293,N_7205,N_6641);
and U8294 (N_8294,N_6062,N_7742);
and U8295 (N_8295,N_7737,N_6311);
nor U8296 (N_8296,N_6010,N_7251);
and U8297 (N_8297,N_6890,N_6894);
nor U8298 (N_8298,N_7651,N_6512);
nand U8299 (N_8299,N_7137,N_7598);
nand U8300 (N_8300,N_6884,N_6267);
xnor U8301 (N_8301,N_6362,N_7354);
xor U8302 (N_8302,N_6465,N_6854);
nor U8303 (N_8303,N_6021,N_7041);
or U8304 (N_8304,N_6004,N_6659);
xnor U8305 (N_8305,N_7802,N_6294);
xor U8306 (N_8306,N_7208,N_7346);
nand U8307 (N_8307,N_6942,N_6243);
or U8308 (N_8308,N_7206,N_6767);
xnor U8309 (N_8309,N_6082,N_6395);
or U8310 (N_8310,N_6638,N_6210);
and U8311 (N_8311,N_7792,N_7931);
and U8312 (N_8312,N_6017,N_6542);
or U8313 (N_8313,N_7930,N_7892);
nor U8314 (N_8314,N_7166,N_7101);
or U8315 (N_8315,N_7440,N_6987);
nand U8316 (N_8316,N_7969,N_6790);
nand U8317 (N_8317,N_6312,N_6806);
nor U8318 (N_8318,N_6526,N_7669);
nor U8319 (N_8319,N_6742,N_7416);
nor U8320 (N_8320,N_7067,N_7793);
or U8321 (N_8321,N_6560,N_7093);
nand U8322 (N_8322,N_7607,N_7342);
xor U8323 (N_8323,N_6672,N_7025);
xor U8324 (N_8324,N_7377,N_6211);
nand U8325 (N_8325,N_6992,N_7056);
or U8326 (N_8326,N_6196,N_6583);
xor U8327 (N_8327,N_7350,N_6031);
and U8328 (N_8328,N_7292,N_6016);
or U8329 (N_8329,N_6594,N_6341);
or U8330 (N_8330,N_6950,N_6674);
nor U8331 (N_8331,N_6804,N_7290);
xnor U8332 (N_8332,N_7001,N_7085);
or U8333 (N_8333,N_7850,N_6394);
and U8334 (N_8334,N_7488,N_6074);
nand U8335 (N_8335,N_6419,N_6107);
nand U8336 (N_8336,N_7286,N_7233);
and U8337 (N_8337,N_7356,N_6869);
and U8338 (N_8338,N_7180,N_7951);
or U8339 (N_8339,N_7295,N_6819);
and U8340 (N_8340,N_6219,N_7988);
or U8341 (N_8341,N_6443,N_6935);
nor U8342 (N_8342,N_6447,N_7659);
and U8343 (N_8343,N_7528,N_7236);
nand U8344 (N_8344,N_7548,N_6941);
or U8345 (N_8345,N_7113,N_6479);
xor U8346 (N_8346,N_6297,N_7867);
and U8347 (N_8347,N_6538,N_7117);
and U8348 (N_8348,N_7345,N_7655);
nor U8349 (N_8349,N_7366,N_6891);
and U8350 (N_8350,N_7489,N_6292);
and U8351 (N_8351,N_6168,N_6156);
xnor U8352 (N_8352,N_7537,N_7433);
or U8353 (N_8353,N_6731,N_6360);
xor U8354 (N_8354,N_6151,N_6142);
or U8355 (N_8355,N_7880,N_6176);
nand U8356 (N_8356,N_6889,N_6726);
and U8357 (N_8357,N_6498,N_6445);
nor U8358 (N_8358,N_6899,N_7810);
nand U8359 (N_8359,N_7613,N_7720);
and U8360 (N_8360,N_7881,N_7852);
xor U8361 (N_8361,N_7392,N_6469);
or U8362 (N_8362,N_7019,N_7615);
or U8363 (N_8363,N_6588,N_6994);
or U8364 (N_8364,N_7619,N_6616);
nor U8365 (N_8365,N_6118,N_6100);
nor U8366 (N_8366,N_7128,N_7162);
nand U8367 (N_8367,N_6782,N_6977);
nand U8368 (N_8368,N_7513,N_6446);
nor U8369 (N_8369,N_6870,N_6626);
xnor U8370 (N_8370,N_7783,N_7291);
xor U8371 (N_8371,N_6172,N_6606);
nand U8372 (N_8372,N_6050,N_6740);
nand U8373 (N_8373,N_7069,N_6492);
nand U8374 (N_8374,N_6877,N_7807);
nor U8375 (N_8375,N_6924,N_6798);
xnor U8376 (N_8376,N_7896,N_6083);
nor U8377 (N_8377,N_6930,N_7167);
and U8378 (N_8378,N_7919,N_6153);
and U8379 (N_8379,N_7135,N_6727);
and U8380 (N_8380,N_7553,N_6087);
xnor U8381 (N_8381,N_7096,N_7411);
nor U8382 (N_8382,N_6076,N_6134);
nor U8383 (N_8383,N_6452,N_7226);
or U8384 (N_8384,N_6980,N_6948);
and U8385 (N_8385,N_6247,N_6316);
nand U8386 (N_8386,N_6823,N_6797);
and U8387 (N_8387,N_6094,N_6345);
or U8388 (N_8388,N_7191,N_7500);
nor U8389 (N_8389,N_7159,N_6351);
nor U8390 (N_8390,N_7336,N_6029);
nand U8391 (N_8391,N_6327,N_6209);
xor U8392 (N_8392,N_7674,N_7344);
xnor U8393 (N_8393,N_6545,N_6287);
nand U8394 (N_8394,N_6608,N_6171);
xor U8395 (N_8395,N_7943,N_6042);
and U8396 (N_8396,N_7866,N_6192);
xor U8397 (N_8397,N_7475,N_6933);
nor U8398 (N_8398,N_6155,N_6985);
nor U8399 (N_8399,N_7751,N_7316);
and U8400 (N_8400,N_7788,N_7748);
xor U8401 (N_8401,N_6393,N_6690);
and U8402 (N_8402,N_7088,N_7774);
xor U8403 (N_8403,N_7585,N_7302);
and U8404 (N_8404,N_6490,N_6898);
nand U8405 (N_8405,N_6336,N_6241);
or U8406 (N_8406,N_7519,N_6573);
or U8407 (N_8407,N_6688,N_7391);
and U8408 (N_8408,N_7715,N_7835);
nor U8409 (N_8409,N_7584,N_7256);
and U8410 (N_8410,N_7724,N_6663);
and U8411 (N_8411,N_6073,N_6559);
and U8412 (N_8412,N_7053,N_7320);
nand U8413 (N_8413,N_6295,N_6259);
nand U8414 (N_8414,N_6461,N_7490);
xor U8415 (N_8415,N_7933,N_6163);
nand U8416 (N_8416,N_7602,N_7016);
xnor U8417 (N_8417,N_7271,N_7176);
xor U8418 (N_8418,N_7015,N_6580);
nor U8419 (N_8419,N_7333,N_7077);
and U8420 (N_8420,N_6505,N_6934);
nor U8421 (N_8421,N_7979,N_7100);
nor U8422 (N_8422,N_6996,N_7287);
or U8423 (N_8423,N_6130,N_6379);
and U8424 (N_8424,N_7653,N_7324);
and U8425 (N_8425,N_6274,N_7853);
and U8426 (N_8426,N_6165,N_6229);
or U8427 (N_8427,N_6265,N_7497);
nand U8428 (N_8428,N_6491,N_6796);
or U8429 (N_8429,N_6991,N_7027);
xor U8430 (N_8430,N_6838,N_7756);
xor U8431 (N_8431,N_7753,N_6769);
xor U8432 (N_8432,N_7691,N_7846);
and U8433 (N_8433,N_6558,N_6544);
and U8434 (N_8434,N_7099,N_6178);
nor U8435 (N_8435,N_6843,N_7851);
nand U8436 (N_8436,N_6376,N_7831);
or U8437 (N_8437,N_7383,N_6864);
xnor U8438 (N_8438,N_6289,N_6770);
xnor U8439 (N_8439,N_7569,N_6799);
and U8440 (N_8440,N_6802,N_6483);
or U8441 (N_8441,N_6277,N_6696);
xor U8442 (N_8442,N_6855,N_7472);
xnor U8443 (N_8443,N_6735,N_7239);
xnor U8444 (N_8444,N_6968,N_6825);
xor U8445 (N_8445,N_7825,N_6786);
or U8446 (N_8446,N_7459,N_7460);
and U8447 (N_8447,N_7534,N_6366);
and U8448 (N_8448,N_6242,N_6283);
or U8449 (N_8449,N_7899,N_6959);
xor U8450 (N_8450,N_7122,N_6699);
or U8451 (N_8451,N_7590,N_6927);
and U8452 (N_8452,N_7421,N_7529);
xnor U8453 (N_8453,N_7735,N_6014);
and U8454 (N_8454,N_7883,N_7474);
xor U8455 (N_8455,N_6754,N_7079);
xnor U8456 (N_8456,N_7948,N_6733);
nor U8457 (N_8457,N_7578,N_6019);
nor U8458 (N_8458,N_7177,N_6907);
xnor U8459 (N_8459,N_7339,N_7960);
or U8460 (N_8460,N_7947,N_7427);
xnor U8461 (N_8461,N_7790,N_6424);
xor U8462 (N_8462,N_6768,N_6779);
xnor U8463 (N_8463,N_7601,N_7741);
nor U8464 (N_8464,N_6553,N_6919);
nand U8465 (N_8465,N_6841,N_7364);
nand U8466 (N_8466,N_6957,N_6643);
nor U8467 (N_8467,N_7803,N_7622);
nor U8468 (N_8468,N_7070,N_6793);
nand U8469 (N_8469,N_6572,N_7120);
xnor U8470 (N_8470,N_6805,N_7305);
nand U8471 (N_8471,N_6857,N_7822);
nand U8472 (N_8472,N_7665,N_7608);
nor U8473 (N_8473,N_7026,N_6601);
or U8474 (N_8474,N_7707,N_7260);
nand U8475 (N_8475,N_7577,N_7449);
or U8476 (N_8476,N_7125,N_6272);
and U8477 (N_8477,N_6913,N_6709);
xnor U8478 (N_8478,N_7706,N_6456);
or U8479 (N_8479,N_6906,N_7512);
or U8480 (N_8480,N_6335,N_7348);
nor U8481 (N_8481,N_7760,N_6646);
nand U8482 (N_8482,N_7804,N_7401);
xor U8483 (N_8483,N_7249,N_7044);
xnor U8484 (N_8484,N_7606,N_6058);
nor U8485 (N_8485,N_7626,N_7722);
nor U8486 (N_8486,N_7224,N_7298);
nor U8487 (N_8487,N_7455,N_7856);
or U8488 (N_8488,N_7431,N_6504);
and U8489 (N_8489,N_7317,N_6308);
or U8490 (N_8490,N_7618,N_7547);
nand U8491 (N_8491,N_7030,N_7684);
or U8492 (N_8492,N_6567,N_7073);
nor U8493 (N_8493,N_7140,N_6762);
xnor U8494 (N_8494,N_6918,N_7970);
xor U8495 (N_8495,N_7595,N_7358);
xnor U8496 (N_8496,N_6410,N_7642);
and U8497 (N_8497,N_6022,N_6408);
xor U8498 (N_8498,N_7118,N_6680);
or U8499 (N_8499,N_7311,N_7000);
nor U8500 (N_8500,N_7641,N_6185);
nand U8501 (N_8501,N_6079,N_6603);
xnor U8502 (N_8502,N_6051,N_7980);
xnor U8503 (N_8503,N_7832,N_6271);
and U8504 (N_8504,N_7714,N_7511);
or U8505 (N_8505,N_6621,N_7262);
nand U8506 (N_8506,N_6876,N_7068);
or U8507 (N_8507,N_6693,N_6849);
nor U8508 (N_8508,N_7160,N_6795);
or U8509 (N_8509,N_7151,N_6691);
nand U8510 (N_8510,N_6057,N_6589);
xor U8511 (N_8511,N_6286,N_6310);
nor U8512 (N_8512,N_6633,N_6714);
or U8513 (N_8513,N_7749,N_7907);
and U8514 (N_8514,N_7736,N_6237);
or U8515 (N_8515,N_7397,N_7014);
nor U8516 (N_8516,N_7134,N_7152);
nor U8517 (N_8517,N_6164,N_6475);
or U8518 (N_8518,N_7461,N_6281);
nor U8519 (N_8519,N_6332,N_7182);
nand U8520 (N_8520,N_6818,N_7981);
nand U8521 (N_8521,N_7982,N_6654);
nor U8522 (N_8522,N_6471,N_6324);
nor U8523 (N_8523,N_7048,N_6071);
xor U8524 (N_8524,N_7676,N_7667);
or U8525 (N_8525,N_7523,N_6328);
or U8526 (N_8526,N_6760,N_7447);
nor U8527 (N_8527,N_7904,N_6997);
xnor U8528 (N_8528,N_6946,N_6161);
nor U8529 (N_8529,N_6543,N_6060);
or U8530 (N_8530,N_7562,N_7268);
and U8531 (N_8531,N_6916,N_7915);
nor U8532 (N_8532,N_6868,N_7834);
xor U8533 (N_8533,N_7673,N_7571);
nand U8534 (N_8534,N_7139,N_6374);
or U8535 (N_8535,N_6183,N_6694);
xnor U8536 (N_8536,N_7367,N_7840);
or U8537 (N_8537,N_7938,N_7238);
nand U8538 (N_8538,N_7050,N_6753);
or U8539 (N_8539,N_7363,N_6367);
nand U8540 (N_8540,N_7185,N_7912);
nor U8541 (N_8541,N_6866,N_6887);
or U8542 (N_8542,N_6174,N_6619);
and U8543 (N_8543,N_7457,N_7076);
nand U8544 (N_8544,N_6450,N_6548);
xnor U8545 (N_8545,N_6126,N_7353);
nor U8546 (N_8546,N_7964,N_7761);
and U8547 (N_8547,N_6384,N_7898);
nor U8548 (N_8548,N_7768,N_7917);
xnor U8549 (N_8549,N_6413,N_6999);
nor U8550 (N_8550,N_7503,N_6334);
nor U8551 (N_8551,N_7683,N_6697);
nand U8552 (N_8552,N_6568,N_6555);
xor U8553 (N_8553,N_6084,N_7957);
nand U8554 (N_8554,N_7150,N_7841);
nor U8555 (N_8555,N_6355,N_6207);
nand U8556 (N_8556,N_7632,N_7954);
xnor U8557 (N_8557,N_7296,N_6222);
xor U8558 (N_8558,N_7805,N_6369);
and U8559 (N_8559,N_7414,N_7241);
nand U8560 (N_8560,N_6309,N_7022);
xnor U8561 (N_8561,N_6622,N_6575);
nand U8562 (N_8562,N_6960,N_7280);
nor U8563 (N_8563,N_6435,N_7796);
or U8564 (N_8564,N_6488,N_6056);
nand U8565 (N_8565,N_6473,N_7109);
xor U8566 (N_8566,N_6679,N_6266);
xor U8567 (N_8567,N_6253,N_7398);
nand U8568 (N_8568,N_7092,N_7149);
xnor U8569 (N_8569,N_7235,N_7108);
and U8570 (N_8570,N_6794,N_6255);
and U8571 (N_8571,N_6858,N_7255);
or U8572 (N_8572,N_6523,N_7926);
and U8573 (N_8573,N_6406,N_6098);
nor U8574 (N_8574,N_7322,N_7340);
xnor U8575 (N_8575,N_6121,N_6116);
or U8576 (N_8576,N_6736,N_7066);
and U8577 (N_8577,N_7006,N_7699);
nor U8578 (N_8578,N_6426,N_7976);
nand U8579 (N_8579,N_7242,N_7972);
nand U8580 (N_8580,N_6472,N_7143);
or U8581 (N_8581,N_6284,N_6781);
or U8582 (N_8582,N_6743,N_6262);
nor U8583 (N_8583,N_7998,N_7473);
and U8584 (N_8584,N_7600,N_6517);
and U8585 (N_8585,N_7341,N_7556);
xnor U8586 (N_8586,N_7328,N_7625);
xnor U8587 (N_8587,N_7538,N_6348);
nor U8588 (N_8588,N_7932,N_7465);
nand U8589 (N_8589,N_6496,N_6839);
nor U8590 (N_8590,N_6947,N_7710);
xnor U8591 (N_8591,N_7894,N_7052);
or U8592 (N_8592,N_6068,N_7884);
nand U8593 (N_8593,N_6339,N_7806);
nand U8594 (N_8594,N_7797,N_7603);
xnor U8595 (N_8595,N_6278,N_6103);
nor U8596 (N_8596,N_6561,N_6766);
nand U8597 (N_8597,N_6214,N_6257);
nand U8598 (N_8598,N_6536,N_7643);
nand U8599 (N_8599,N_6280,N_7539);
or U8600 (N_8600,N_6244,N_7165);
or U8601 (N_8601,N_6650,N_6009);
or U8602 (N_8602,N_6631,N_7897);
nor U8603 (N_8603,N_6850,N_7874);
or U8604 (N_8604,N_7104,N_6812);
xnor U8605 (N_8605,N_6829,N_7429);
and U8606 (N_8606,N_7811,N_7660);
or U8607 (N_8607,N_6080,N_6649);
or U8608 (N_8608,N_6725,N_6552);
or U8609 (N_8609,N_7404,N_7791);
nor U8610 (N_8610,N_6096,N_7704);
or U8611 (N_8611,N_6592,N_6437);
and U8612 (N_8612,N_6707,N_6613);
nand U8613 (N_8613,N_7412,N_7541);
nand U8614 (N_8614,N_6704,N_7470);
nand U8615 (N_8615,N_6635,N_6493);
and U8616 (N_8616,N_6527,N_6365);
and U8617 (N_8617,N_7471,N_7220);
nand U8618 (N_8618,N_7499,N_6002);
nor U8619 (N_8619,N_7836,N_6288);
nand U8620 (N_8620,N_7408,N_6097);
nand U8621 (N_8621,N_6357,N_6220);
and U8622 (N_8622,N_7842,N_7900);
or U8623 (N_8623,N_6361,N_6053);
nand U8624 (N_8624,N_7552,N_7486);
and U8625 (N_8625,N_6510,N_7716);
and U8626 (N_8626,N_6063,N_7701);
xnor U8627 (N_8627,N_6578,N_6417);
and U8628 (N_8628,N_6928,N_6713);
nand U8629 (N_8629,N_6739,N_7002);
nand U8630 (N_8630,N_6034,N_7903);
and U8631 (N_8631,N_6431,N_7217);
and U8632 (N_8632,N_7187,N_7530);
and U8633 (N_8633,N_7081,N_6953);
nand U8634 (N_8634,N_7819,N_7627);
xor U8635 (N_8635,N_6319,N_7635);
nor U8636 (N_8636,N_6036,N_6363);
xor U8637 (N_8637,N_7270,N_6293);
nand U8638 (N_8638,N_7687,N_7155);
or U8639 (N_8639,N_7089,N_7444);
nand U8640 (N_8640,N_7161,N_7587);
xnor U8641 (N_8641,N_6205,N_7515);
nand U8642 (N_8642,N_6678,N_7886);
and U8643 (N_8643,N_7762,N_6359);
xor U8644 (N_8644,N_6356,N_6313);
nand U8645 (N_8645,N_7269,N_7983);
or U8646 (N_8646,N_7709,N_6495);
nand U8647 (N_8647,N_6939,N_7478);
or U8648 (N_8648,N_6652,N_7989);
nand U8649 (N_8649,N_6477,N_6186);
or U8650 (N_8650,N_7871,N_6416);
xnor U8651 (N_8651,N_7332,N_7259);
nor U8652 (N_8652,N_6454,N_6810);
nor U8653 (N_8653,N_7527,N_7493);
nor U8654 (N_8654,N_7682,N_7757);
or U8655 (N_8655,N_7733,N_7253);
and U8656 (N_8656,N_6689,N_7574);
or U8657 (N_8657,N_6895,N_7984);
xor U8658 (N_8658,N_6856,N_7189);
xor U8659 (N_8659,N_7920,N_6385);
and U8660 (N_8660,N_6216,N_7278);
and U8661 (N_8661,N_7240,N_6511);
xor U8662 (N_8662,N_6880,N_6352);
nor U8663 (N_8663,N_7755,N_6557);
and U8664 (N_8664,N_7833,N_7452);
nor U8665 (N_8665,N_6936,N_6448);
or U8666 (N_8666,N_7764,N_7929);
xnor U8667 (N_8667,N_7502,N_7671);
and U8668 (N_8668,N_7141,N_7747);
xor U8669 (N_8669,N_6719,N_6824);
and U8670 (N_8670,N_7445,N_6920);
and U8671 (N_8671,N_7172,N_6878);
nor U8672 (N_8672,N_7468,N_7375);
nor U8673 (N_8673,N_7506,N_7406);
or U8674 (N_8674,N_6371,N_7564);
or U8675 (N_8675,N_6840,N_7075);
xnor U8676 (N_8676,N_6187,N_7132);
nor U8677 (N_8677,N_7114,N_7567);
and U8678 (N_8678,N_6279,N_6591);
nor U8679 (N_8679,N_6705,N_7147);
nor U8680 (N_8680,N_7082,N_7400);
nor U8681 (N_8681,N_6614,N_7908);
xor U8682 (N_8682,N_6129,N_7617);
and U8683 (N_8683,N_6822,N_6965);
nand U8684 (N_8684,N_6078,N_6389);
nor U8685 (N_8685,N_7428,N_6260);
and U8686 (N_8686,N_7110,N_7321);
nand U8687 (N_8687,N_6148,N_7190);
xor U8688 (N_8688,N_7247,N_7902);
xor U8689 (N_8689,N_7201,N_6476);
or U8690 (N_8690,N_7843,N_6089);
nand U8691 (N_8691,N_6785,N_7723);
nor U8692 (N_8692,N_7634,N_6453);
xor U8693 (N_8693,N_6175,N_7112);
or U8694 (N_8694,N_7668,N_6979);
nand U8695 (N_8695,N_7863,N_6268);
xnor U8696 (N_8696,N_6501,N_6909);
xnor U8697 (N_8697,N_6349,N_6896);
nand U8698 (N_8698,N_7410,N_6651);
nand U8699 (N_8699,N_6146,N_7380);
and U8700 (N_8700,N_7031,N_7288);
xor U8701 (N_8701,N_6455,N_7732);
xor U8702 (N_8702,N_7873,N_7039);
xnor U8703 (N_8703,N_7164,N_6771);
nand U8704 (N_8704,N_6436,N_7910);
xnor U8705 (N_8705,N_6998,N_7359);
nand U8706 (N_8706,N_7314,N_7148);
xor U8707 (N_8707,N_7794,N_7049);
nand U8708 (N_8708,N_6815,N_6054);
nor U8709 (N_8709,N_6015,N_6710);
and U8710 (N_8710,N_6282,N_7859);
or U8711 (N_8711,N_6329,N_6637);
or U8712 (N_8712,N_6181,N_7153);
xor U8713 (N_8713,N_6788,N_7589);
nand U8714 (N_8714,N_7325,N_7485);
and U8715 (N_8715,N_6199,N_7186);
nand U8716 (N_8716,N_6249,N_7766);
nor U8717 (N_8717,N_7482,N_6404);
or U8718 (N_8718,N_6662,N_7481);
nor U8719 (N_8719,N_6364,N_6582);
and U8720 (N_8720,N_6157,N_7561);
xor U8721 (N_8721,N_7204,N_6671);
nor U8722 (N_8722,N_6099,N_7413);
nor U8723 (N_8723,N_6577,N_6566);
or U8724 (N_8724,N_7611,N_7307);
nand U8725 (N_8725,N_6828,N_6013);
nand U8726 (N_8726,N_7028,N_7570);
xor U8727 (N_8727,N_6432,N_6596);
xor U8728 (N_8728,N_7443,N_7554);
nand U8729 (N_8729,N_7265,N_7237);
xnor U8730 (N_8730,N_7371,N_6167);
nor U8731 (N_8731,N_6011,N_6046);
nand U8732 (N_8732,N_7640,N_7157);
nor U8733 (N_8733,N_6276,N_7532);
and U8734 (N_8734,N_7905,N_6238);
nor U8735 (N_8735,N_6862,N_7997);
or U8736 (N_8736,N_6003,N_6604);
nor U8737 (N_8737,N_7559,N_6695);
and U8738 (N_8738,N_6639,N_6402);
nor U8739 (N_8739,N_7248,N_7909);
xnor U8740 (N_8740,N_7263,N_7827);
nand U8741 (N_8741,N_7246,N_6045);
xor U8742 (N_8742,N_6388,N_7913);
and U8743 (N_8743,N_7594,N_6397);
nor U8744 (N_8744,N_7633,N_7639);
and U8745 (N_8745,N_7612,N_7432);
and U8746 (N_8746,N_6300,N_6535);
or U8747 (N_8747,N_7170,N_7771);
nor U8748 (N_8748,N_7261,N_7677);
nor U8749 (N_8749,N_6872,N_7726);
or U8750 (N_8750,N_6665,N_7780);
nand U8751 (N_8751,N_7309,N_6420);
nor U8752 (N_8752,N_6200,N_6685);
xnor U8753 (N_8753,N_7415,N_7934);
xor U8754 (N_8754,N_7451,N_6102);
xnor U8755 (N_8755,N_7967,N_6964);
or U8756 (N_8756,N_7409,N_7535);
nor U8757 (N_8757,N_7329,N_7193);
or U8758 (N_8758,N_7799,N_7491);
or U8759 (N_8759,N_7614,N_7405);
or U8760 (N_8760,N_6012,N_6133);
and U8761 (N_8761,N_7809,N_6202);
or U8762 (N_8762,N_6618,N_7448);
and U8763 (N_8763,N_6820,N_7824);
nand U8764 (N_8764,N_6888,N_6549);
or U8765 (N_8765,N_6143,N_6438);
nor U8766 (N_8766,N_7560,N_6718);
xor U8767 (N_8767,N_7267,N_7385);
xnor U8768 (N_8768,N_7645,N_7315);
or U8769 (N_8769,N_6170,N_7944);
and U8770 (N_8770,N_7719,N_7303);
or U8771 (N_8771,N_6562,N_6611);
nand U8772 (N_8772,N_7379,N_7087);
nor U8773 (N_8773,N_7034,N_7524);
nand U8774 (N_8774,N_7837,N_6500);
nand U8775 (N_8775,N_6487,N_6595);
and U8776 (N_8776,N_7705,N_6605);
nand U8777 (N_8777,N_6020,N_6627);
nand U8778 (N_8778,N_6834,N_6642);
nor U8779 (N_8779,N_7914,N_6931);
and U8780 (N_8780,N_6194,N_7599);
nor U8781 (N_8781,N_6832,N_7272);
nor U8782 (N_8782,N_6039,N_7035);
xor U8783 (N_8783,N_7362,N_6720);
or U8784 (N_8784,N_6773,N_7924);
xor U8785 (N_8785,N_6530,N_7784);
or U8786 (N_8786,N_7870,N_7718);
nor U8787 (N_8787,N_6816,N_6179);
xnor U8788 (N_8788,N_6666,N_6982);
nand U8789 (N_8789,N_6474,N_6989);
nand U8790 (N_8790,N_6423,N_7183);
nor U8791 (N_8791,N_7327,N_6972);
or U8792 (N_8792,N_6661,N_6141);
and U8793 (N_8793,N_6540,N_7127);
nand U8794 (N_8794,N_6005,N_6470);
nor U8795 (N_8795,N_7820,N_7198);
and U8796 (N_8796,N_6444,N_6405);
and U8797 (N_8797,N_7888,N_7814);
nor U8798 (N_8798,N_6189,N_6506);
nor U8799 (N_8799,N_6961,N_7666);
nor U8800 (N_8800,N_7700,N_7991);
nor U8801 (N_8801,N_6127,N_7370);
or U8802 (N_8802,N_7911,N_7365);
xnor U8803 (N_8803,N_6040,N_7126);
and U8804 (N_8804,N_7289,N_6136);
xor U8805 (N_8805,N_6038,N_7047);
nand U8806 (N_8806,N_7695,N_7579);
nor U8807 (N_8807,N_6717,N_7576);
nor U8808 (N_8808,N_6509,N_7252);
nor U8809 (N_8809,N_7844,N_6716);
nand U8810 (N_8810,N_7098,N_6481);
nor U8811 (N_8811,N_6847,N_7196);
xnor U8812 (N_8812,N_6904,N_6803);
and U8813 (N_8813,N_6955,N_7243);
xnor U8814 (N_8814,N_7728,N_7254);
xnor U8815 (N_8815,N_6759,N_7244);
or U8816 (N_8816,N_7009,N_7812);
nand U8817 (N_8817,N_6457,N_6494);
nand U8818 (N_8818,N_6983,N_7767);
xor U8819 (N_8819,N_6203,N_6932);
nor U8820 (N_8820,N_7216,N_6925);
nand U8821 (N_8821,N_7277,N_7977);
xnor U8822 (N_8822,N_7361,N_6546);
or U8823 (N_8823,N_7536,N_6326);
or U8824 (N_8824,N_7168,N_7877);
and U8825 (N_8825,N_7396,N_7285);
nand U8826 (N_8826,N_6235,N_6629);
nand U8827 (N_8827,N_6044,N_7816);
or U8828 (N_8828,N_6851,N_6052);
nor U8829 (N_8829,N_6227,N_7061);
nand U8830 (N_8830,N_7071,N_6809);
nor U8831 (N_8831,N_7299,N_7916);
nand U8832 (N_8832,N_7746,N_6956);
xnor U8833 (N_8833,N_7017,N_7378);
xnor U8834 (N_8834,N_6711,N_6625);
nor U8835 (N_8835,N_7628,N_6723);
nand U8836 (N_8836,N_6502,N_7095);
and U8837 (N_8837,N_6524,N_7145);
nand U8838 (N_8838,N_7279,N_6516);
and U8839 (N_8839,N_7965,N_7097);
or U8840 (N_8840,N_7136,N_6745);
nand U8841 (N_8841,N_7744,N_7901);
nand U8842 (N_8842,N_6859,N_7212);
or U8843 (N_8843,N_6503,N_6399);
or U8844 (N_8844,N_6337,N_6599);
nand U8845 (N_8845,N_6023,N_7941);
nor U8846 (N_8846,N_6252,N_7765);
xnor U8847 (N_8847,N_6478,N_7966);
xnor U8848 (N_8848,N_6949,N_6800);
nand U8849 (N_8849,N_6550,N_7349);
xor U8850 (N_8850,N_7823,N_6273);
nand U8851 (N_8851,N_7426,N_6007);
and U8852 (N_8852,N_6069,N_6863);
and U8853 (N_8853,N_6586,N_6747);
nor U8854 (N_8854,N_7862,N_7210);
nand U8855 (N_8855,N_6686,N_7680);
and U8856 (N_8856,N_6765,N_6835);
and U8857 (N_8857,N_6221,N_7300);
and U8858 (N_8858,N_6228,N_6682);
or U8859 (N_8859,N_7393,N_6978);
xor U8860 (N_8860,N_6462,N_6827);
and U8861 (N_8861,N_6375,N_6232);
nand U8862 (N_8862,N_7555,N_7033);
xnor U8863 (N_8863,N_7740,N_7313);
and U8864 (N_8864,N_6874,N_7581);
xnor U8865 (N_8865,N_6064,N_6314);
nor U8866 (N_8866,N_6923,N_7194);
xor U8867 (N_8867,N_6303,N_6401);
xor U8868 (N_8868,N_6409,N_7923);
nor U8869 (N_8869,N_7390,N_6984);
or U8870 (N_8870,N_6264,N_6908);
nand U8871 (N_8871,N_6191,N_7963);
or U8872 (N_8872,N_6441,N_6340);
nand U8873 (N_8873,N_7057,N_6158);
nor U8874 (N_8874,N_6131,N_6246);
xnor U8875 (N_8875,N_7939,N_6600);
xor U8876 (N_8876,N_6085,N_6233);
xnor U8877 (N_8877,N_7060,N_7546);
xor U8878 (N_8878,N_6830,N_6774);
nand U8879 (N_8879,N_6917,N_6741);
nand U8880 (N_8880,N_6981,N_6250);
nand U8881 (N_8881,N_6236,N_7462);
or U8882 (N_8882,N_7029,N_7111);
nor U8883 (N_8883,N_6831,N_6338);
xor U8884 (N_8884,N_6497,N_7708);
and U8885 (N_8885,N_7604,N_6647);
nor U8886 (N_8886,N_6970,N_6640);
and U8887 (N_8887,N_7656,N_7637);
or U8888 (N_8888,N_6317,N_7826);
xor U8889 (N_8889,N_7937,N_7885);
and U8890 (N_8890,N_6213,N_6299);
nor U8891 (N_8891,N_7003,N_7381);
xnor U8892 (N_8892,N_6035,N_7685);
xnor U8893 (N_8893,N_6117,N_6061);
xnor U8894 (N_8894,N_7781,N_6429);
nand U8895 (N_8895,N_6911,N_7293);
or U8896 (N_8896,N_6648,N_6563);
nand U8897 (N_8897,N_7422,N_6657);
and U8898 (N_8898,N_7696,N_7231);
nor U8899 (N_8899,N_6234,N_7657);
nand U8900 (N_8900,N_7878,N_7782);
nor U8901 (N_8901,N_6263,N_6088);
or U8902 (N_8902,N_7373,N_7439);
xor U8903 (N_8903,N_6700,N_7838);
nor U8904 (N_8904,N_7477,N_6000);
nor U8905 (N_8905,N_6732,N_6086);
nand U8906 (N_8906,N_7887,N_7990);
nor U8907 (N_8907,N_7129,N_7338);
xor U8908 (N_8908,N_6382,N_6669);
xor U8909 (N_8909,N_7891,N_6715);
nor U8910 (N_8910,N_6378,N_7388);
nor U8911 (N_8911,N_6945,N_6615);
and U8912 (N_8912,N_7197,N_7273);
nor U8913 (N_8913,N_7521,N_7225);
or U8914 (N_8914,N_6486,N_6430);
nand U8915 (N_8915,N_6291,N_6744);
nand U8916 (N_8916,N_6940,N_7083);
or U8917 (N_8917,N_6722,N_7323);
or U8918 (N_8918,N_7174,N_6460);
nor U8919 (N_8919,N_6001,N_7051);
nand U8920 (N_8920,N_7484,N_7623);
and U8921 (N_8921,N_7994,N_6104);
and U8922 (N_8922,N_7417,N_6976);
nor U8923 (N_8923,N_6764,N_7830);
nand U8924 (N_8924,N_6149,N_7582);
and U8925 (N_8925,N_6226,N_6873);
or U8926 (N_8926,N_7652,N_7192);
nor U8927 (N_8927,N_7374,N_7828);
and U8928 (N_8928,N_7636,N_6750);
xor U8929 (N_8929,N_7334,N_7985);
nand U8930 (N_8930,N_6902,N_7959);
or U8931 (N_8931,N_7215,N_7284);
nor U8932 (N_8932,N_7650,N_7813);
or U8933 (N_8933,N_6724,N_6617);
and U8934 (N_8934,N_7759,N_6708);
nand U8935 (N_8935,N_7228,N_7352);
nor U8936 (N_8936,N_7675,N_7479);
and U8937 (N_8937,N_6105,N_7074);
nor U8938 (N_8938,N_7184,N_7785);
xor U8939 (N_8939,N_6914,N_7593);
xor U8940 (N_8940,N_6358,N_7384);
xor U8941 (N_8941,N_7199,N_7106);
nor U8942 (N_8942,N_6414,N_6721);
nand U8943 (N_8943,N_6331,N_6791);
and U8944 (N_8944,N_6041,N_6387);
nand U8945 (N_8945,N_7522,N_6598);
nand U8946 (N_8946,N_6386,N_7516);
nor U8947 (N_8947,N_6458,N_7697);
nor U8948 (N_8948,N_7407,N_7752);
and U8949 (N_8949,N_6122,N_7102);
xor U8950 (N_8950,N_6853,N_7921);
nor U8951 (N_8951,N_7800,N_7476);
nand U8952 (N_8952,N_6344,N_7918);
nor U8953 (N_8953,N_6033,N_7540);
or U8954 (N_8954,N_6892,N_7018);
nand U8955 (N_8955,N_7146,N_6055);
nand U8956 (N_8956,N_6602,N_6761);
and U8957 (N_8957,N_6763,N_7504);
nor U8958 (N_8958,N_7138,N_7312);
and U8959 (N_8959,N_6307,N_7454);
nand U8960 (N_8960,N_6463,N_7037);
xnor U8961 (N_8961,N_6706,N_7080);
nor U8962 (N_8962,N_6188,N_6846);
nand U8963 (N_8963,N_7121,N_7456);
nand U8964 (N_8964,N_7347,N_6837);
or U8965 (N_8965,N_7795,N_6347);
nand U8966 (N_8966,N_7712,N_7686);
and U8967 (N_8967,N_6113,N_6988);
or U8968 (N_8968,N_6123,N_6963);
xor U8969 (N_8969,N_6125,N_6581);
nor U8970 (N_8970,N_6734,N_6169);
or U8971 (N_8971,N_7927,N_7616);
and U8972 (N_8972,N_7952,N_6254);
nor U8973 (N_8973,N_6630,N_6182);
and U8974 (N_8974,N_6139,N_6871);
nor U8975 (N_8975,N_6372,N_6787);
and U8976 (N_8976,N_6756,N_6929);
nor U8977 (N_8977,N_6159,N_7962);
xor U8978 (N_8978,N_7230,N_7387);
or U8979 (N_8979,N_7103,N_6177);
nor U8980 (N_8980,N_7845,N_6587);
or U8981 (N_8981,N_6670,N_6848);
nor U8982 (N_8982,N_6755,N_6821);
xor U8983 (N_8983,N_6971,N_7545);
nor U8984 (N_8984,N_6109,N_6305);
nand U8985 (N_8985,N_7178,N_6018);
xnor U8986 (N_8986,N_7517,N_7064);
nor U8987 (N_8987,N_7469,N_7661);
or U8988 (N_8988,N_7463,N_7011);
nor U8989 (N_8989,N_6702,N_7091);
and U8990 (N_8990,N_6675,N_6814);
nor U8991 (N_8991,N_7936,N_7906);
nor U8992 (N_8992,N_7526,N_7389);
nor U8993 (N_8993,N_6645,N_7266);
and U8994 (N_8994,N_6030,N_7638);
nor U8995 (N_8995,N_6632,N_7882);
or U8996 (N_8996,N_7777,N_6315);
xnor U8997 (N_8997,N_7395,N_7971);
or U8998 (N_8998,N_6270,N_6077);
nand U8999 (N_8999,N_7855,N_6752);
nor U9000 (N_9000,N_6725,N_7140);
nor U9001 (N_9001,N_7109,N_6026);
xnor U9002 (N_9002,N_7785,N_6060);
nor U9003 (N_9003,N_7811,N_6286);
and U9004 (N_9004,N_6166,N_6141);
and U9005 (N_9005,N_7167,N_6503);
xor U9006 (N_9006,N_7812,N_7780);
xor U9007 (N_9007,N_6912,N_6223);
and U9008 (N_9008,N_7061,N_6151);
and U9009 (N_9009,N_7198,N_6868);
xnor U9010 (N_9010,N_6368,N_6967);
nand U9011 (N_9011,N_7990,N_6315);
or U9012 (N_9012,N_6969,N_6470);
nand U9013 (N_9013,N_7589,N_6462);
xnor U9014 (N_9014,N_6286,N_7169);
nor U9015 (N_9015,N_7069,N_6150);
and U9016 (N_9016,N_7139,N_6267);
or U9017 (N_9017,N_6709,N_6556);
nand U9018 (N_9018,N_7520,N_6158);
nor U9019 (N_9019,N_6656,N_7763);
and U9020 (N_9020,N_7424,N_6639);
nor U9021 (N_9021,N_6960,N_6462);
nand U9022 (N_9022,N_6135,N_7888);
and U9023 (N_9023,N_6655,N_6845);
xnor U9024 (N_9024,N_7778,N_6615);
xnor U9025 (N_9025,N_7330,N_7357);
and U9026 (N_9026,N_6996,N_6481);
and U9027 (N_9027,N_7264,N_6807);
and U9028 (N_9028,N_7019,N_7486);
xor U9029 (N_9029,N_7568,N_7863);
xnor U9030 (N_9030,N_6564,N_6471);
or U9031 (N_9031,N_7425,N_7930);
nor U9032 (N_9032,N_6663,N_6574);
nand U9033 (N_9033,N_6327,N_7456);
xnor U9034 (N_9034,N_7538,N_7442);
and U9035 (N_9035,N_6025,N_7648);
xnor U9036 (N_9036,N_6850,N_7517);
and U9037 (N_9037,N_7292,N_7746);
nor U9038 (N_9038,N_6172,N_7918);
and U9039 (N_9039,N_6582,N_7345);
nand U9040 (N_9040,N_6190,N_7272);
nor U9041 (N_9041,N_6194,N_7359);
nand U9042 (N_9042,N_6608,N_7597);
nor U9043 (N_9043,N_7185,N_6651);
nor U9044 (N_9044,N_6071,N_6983);
and U9045 (N_9045,N_7772,N_6416);
xor U9046 (N_9046,N_7532,N_7412);
nand U9047 (N_9047,N_6525,N_6747);
nor U9048 (N_9048,N_7380,N_6478);
nor U9049 (N_9049,N_7617,N_7691);
or U9050 (N_9050,N_7575,N_7019);
nor U9051 (N_9051,N_7656,N_6613);
and U9052 (N_9052,N_7113,N_7770);
or U9053 (N_9053,N_6665,N_6233);
nor U9054 (N_9054,N_6599,N_7365);
nand U9055 (N_9055,N_6205,N_6862);
nand U9056 (N_9056,N_6252,N_7415);
and U9057 (N_9057,N_7075,N_6784);
and U9058 (N_9058,N_6836,N_7238);
or U9059 (N_9059,N_7038,N_6146);
and U9060 (N_9060,N_6456,N_6972);
or U9061 (N_9061,N_7046,N_7822);
or U9062 (N_9062,N_6472,N_6851);
nor U9063 (N_9063,N_6408,N_6866);
xor U9064 (N_9064,N_7278,N_6064);
nor U9065 (N_9065,N_7047,N_6669);
nand U9066 (N_9066,N_6298,N_7176);
or U9067 (N_9067,N_6656,N_7751);
or U9068 (N_9068,N_7585,N_6455);
nor U9069 (N_9069,N_7508,N_7256);
nor U9070 (N_9070,N_7604,N_7338);
nand U9071 (N_9071,N_6725,N_6665);
and U9072 (N_9072,N_7488,N_7994);
nand U9073 (N_9073,N_6853,N_7610);
or U9074 (N_9074,N_6275,N_6651);
and U9075 (N_9075,N_6693,N_6279);
nor U9076 (N_9076,N_6865,N_7873);
or U9077 (N_9077,N_6171,N_6744);
or U9078 (N_9078,N_7992,N_7798);
nand U9079 (N_9079,N_7308,N_7961);
nand U9080 (N_9080,N_6493,N_6670);
or U9081 (N_9081,N_6196,N_6939);
nand U9082 (N_9082,N_7637,N_7808);
nand U9083 (N_9083,N_7377,N_7285);
nor U9084 (N_9084,N_7331,N_6593);
nand U9085 (N_9085,N_6089,N_6867);
or U9086 (N_9086,N_7000,N_7201);
nor U9087 (N_9087,N_6984,N_6468);
xor U9088 (N_9088,N_6318,N_7275);
nand U9089 (N_9089,N_7300,N_6162);
or U9090 (N_9090,N_7623,N_7434);
or U9091 (N_9091,N_7828,N_6415);
nand U9092 (N_9092,N_7845,N_7204);
or U9093 (N_9093,N_7100,N_7688);
nor U9094 (N_9094,N_7492,N_6675);
nand U9095 (N_9095,N_6208,N_6397);
nand U9096 (N_9096,N_6220,N_6672);
nand U9097 (N_9097,N_6930,N_6391);
and U9098 (N_9098,N_6091,N_7310);
nand U9099 (N_9099,N_6894,N_6919);
or U9100 (N_9100,N_6113,N_7720);
and U9101 (N_9101,N_7252,N_6820);
or U9102 (N_9102,N_6188,N_6661);
and U9103 (N_9103,N_7916,N_6044);
and U9104 (N_9104,N_7938,N_7952);
and U9105 (N_9105,N_6661,N_6502);
and U9106 (N_9106,N_6383,N_7263);
and U9107 (N_9107,N_6900,N_6151);
xor U9108 (N_9108,N_6309,N_7364);
nor U9109 (N_9109,N_7271,N_7474);
xor U9110 (N_9110,N_7944,N_7196);
nor U9111 (N_9111,N_6584,N_7741);
nand U9112 (N_9112,N_7438,N_6892);
or U9113 (N_9113,N_6484,N_7192);
and U9114 (N_9114,N_7828,N_7876);
or U9115 (N_9115,N_7925,N_7191);
and U9116 (N_9116,N_7712,N_6252);
nand U9117 (N_9117,N_6198,N_7336);
nor U9118 (N_9118,N_7031,N_7482);
xor U9119 (N_9119,N_7628,N_7298);
and U9120 (N_9120,N_7923,N_6125);
nor U9121 (N_9121,N_6320,N_6253);
nor U9122 (N_9122,N_6999,N_6958);
or U9123 (N_9123,N_7934,N_6081);
nor U9124 (N_9124,N_7000,N_6615);
xnor U9125 (N_9125,N_7212,N_7174);
nor U9126 (N_9126,N_7237,N_6212);
and U9127 (N_9127,N_6010,N_7827);
xor U9128 (N_9128,N_6732,N_6838);
nor U9129 (N_9129,N_7327,N_7349);
or U9130 (N_9130,N_7459,N_7823);
and U9131 (N_9131,N_7224,N_7769);
nand U9132 (N_9132,N_7265,N_6817);
nand U9133 (N_9133,N_6358,N_6243);
or U9134 (N_9134,N_7651,N_7758);
nand U9135 (N_9135,N_7166,N_7555);
nand U9136 (N_9136,N_6332,N_7097);
or U9137 (N_9137,N_6037,N_7486);
nor U9138 (N_9138,N_7545,N_6022);
or U9139 (N_9139,N_6304,N_6033);
xor U9140 (N_9140,N_6643,N_6630);
xor U9141 (N_9141,N_7637,N_6492);
and U9142 (N_9142,N_6908,N_6145);
and U9143 (N_9143,N_6463,N_6038);
or U9144 (N_9144,N_7717,N_6601);
nand U9145 (N_9145,N_7242,N_6268);
and U9146 (N_9146,N_6879,N_6892);
xor U9147 (N_9147,N_7925,N_7293);
xnor U9148 (N_9148,N_7795,N_7798);
xnor U9149 (N_9149,N_6965,N_7457);
nand U9150 (N_9150,N_6366,N_7514);
xnor U9151 (N_9151,N_7054,N_6605);
nand U9152 (N_9152,N_7880,N_7188);
nand U9153 (N_9153,N_6714,N_6855);
nand U9154 (N_9154,N_6510,N_6551);
and U9155 (N_9155,N_7427,N_6835);
nor U9156 (N_9156,N_7985,N_6915);
xnor U9157 (N_9157,N_6543,N_6844);
nand U9158 (N_9158,N_7605,N_6795);
nand U9159 (N_9159,N_6760,N_6851);
and U9160 (N_9160,N_7515,N_7456);
xor U9161 (N_9161,N_6455,N_7246);
nand U9162 (N_9162,N_6754,N_6142);
and U9163 (N_9163,N_6280,N_6397);
xor U9164 (N_9164,N_7826,N_7006);
xor U9165 (N_9165,N_7987,N_6287);
nor U9166 (N_9166,N_6128,N_7858);
nand U9167 (N_9167,N_6952,N_7405);
xor U9168 (N_9168,N_6643,N_7198);
or U9169 (N_9169,N_6187,N_7026);
xnor U9170 (N_9170,N_6966,N_6130);
nand U9171 (N_9171,N_7826,N_7584);
nor U9172 (N_9172,N_6586,N_6931);
and U9173 (N_9173,N_6514,N_7242);
nor U9174 (N_9174,N_7221,N_7253);
and U9175 (N_9175,N_7531,N_7998);
nor U9176 (N_9176,N_6293,N_6590);
nor U9177 (N_9177,N_7463,N_6323);
nor U9178 (N_9178,N_6515,N_6767);
nor U9179 (N_9179,N_6323,N_6148);
and U9180 (N_9180,N_6807,N_7896);
or U9181 (N_9181,N_6371,N_6538);
xnor U9182 (N_9182,N_6795,N_7107);
or U9183 (N_9183,N_7780,N_6248);
or U9184 (N_9184,N_6241,N_6565);
nor U9185 (N_9185,N_6469,N_7188);
and U9186 (N_9186,N_7245,N_6923);
xnor U9187 (N_9187,N_6242,N_7868);
nor U9188 (N_9188,N_7362,N_6344);
nand U9189 (N_9189,N_6405,N_7786);
xnor U9190 (N_9190,N_6440,N_7477);
or U9191 (N_9191,N_7674,N_6928);
xnor U9192 (N_9192,N_7497,N_7349);
xor U9193 (N_9193,N_7713,N_6482);
and U9194 (N_9194,N_7671,N_7553);
nand U9195 (N_9195,N_6694,N_7297);
or U9196 (N_9196,N_7612,N_7842);
or U9197 (N_9197,N_6606,N_6660);
nor U9198 (N_9198,N_6188,N_6899);
or U9199 (N_9199,N_7306,N_7564);
xnor U9200 (N_9200,N_7308,N_6329);
xnor U9201 (N_9201,N_6383,N_6796);
nor U9202 (N_9202,N_7158,N_6525);
or U9203 (N_9203,N_6558,N_6228);
xor U9204 (N_9204,N_7146,N_7024);
nand U9205 (N_9205,N_7877,N_7441);
or U9206 (N_9206,N_7346,N_6405);
nor U9207 (N_9207,N_7215,N_7186);
nor U9208 (N_9208,N_6712,N_7454);
xor U9209 (N_9209,N_7603,N_6066);
xnor U9210 (N_9210,N_7964,N_6584);
nand U9211 (N_9211,N_7581,N_7882);
xor U9212 (N_9212,N_7042,N_6581);
or U9213 (N_9213,N_6115,N_7366);
nand U9214 (N_9214,N_6767,N_7067);
or U9215 (N_9215,N_7181,N_7417);
nand U9216 (N_9216,N_6427,N_6439);
or U9217 (N_9217,N_7482,N_7585);
xnor U9218 (N_9218,N_7719,N_6655);
nand U9219 (N_9219,N_6627,N_7226);
nor U9220 (N_9220,N_7253,N_7297);
xnor U9221 (N_9221,N_6658,N_7597);
nor U9222 (N_9222,N_7660,N_7382);
nand U9223 (N_9223,N_6221,N_6426);
or U9224 (N_9224,N_6959,N_6720);
nand U9225 (N_9225,N_6080,N_6928);
xnor U9226 (N_9226,N_6651,N_7551);
xor U9227 (N_9227,N_7973,N_7358);
or U9228 (N_9228,N_6813,N_7162);
nand U9229 (N_9229,N_7675,N_6616);
xnor U9230 (N_9230,N_6719,N_7041);
nand U9231 (N_9231,N_7285,N_6607);
nand U9232 (N_9232,N_6772,N_7943);
xnor U9233 (N_9233,N_7848,N_7864);
nand U9234 (N_9234,N_6369,N_6602);
xnor U9235 (N_9235,N_7983,N_7848);
nand U9236 (N_9236,N_6069,N_6116);
nand U9237 (N_9237,N_7082,N_6064);
nor U9238 (N_9238,N_6804,N_6729);
xor U9239 (N_9239,N_7167,N_6324);
nand U9240 (N_9240,N_6183,N_6498);
nand U9241 (N_9241,N_7237,N_6496);
or U9242 (N_9242,N_6600,N_7987);
or U9243 (N_9243,N_7996,N_6948);
nor U9244 (N_9244,N_7332,N_7468);
xor U9245 (N_9245,N_6753,N_6114);
and U9246 (N_9246,N_7444,N_6667);
or U9247 (N_9247,N_7001,N_6190);
or U9248 (N_9248,N_6742,N_7439);
nand U9249 (N_9249,N_6134,N_7759);
nand U9250 (N_9250,N_7296,N_7715);
and U9251 (N_9251,N_6145,N_6681);
or U9252 (N_9252,N_7020,N_6949);
xor U9253 (N_9253,N_6246,N_6289);
nor U9254 (N_9254,N_7967,N_7265);
and U9255 (N_9255,N_7520,N_7862);
nor U9256 (N_9256,N_6501,N_7186);
nand U9257 (N_9257,N_7041,N_7866);
or U9258 (N_9258,N_7041,N_6833);
and U9259 (N_9259,N_6634,N_7136);
nand U9260 (N_9260,N_6695,N_7205);
nand U9261 (N_9261,N_6607,N_7211);
or U9262 (N_9262,N_6016,N_6251);
xor U9263 (N_9263,N_7219,N_6484);
nor U9264 (N_9264,N_7883,N_7641);
nand U9265 (N_9265,N_6585,N_6202);
or U9266 (N_9266,N_7095,N_7908);
xor U9267 (N_9267,N_7296,N_6862);
or U9268 (N_9268,N_7363,N_7265);
xor U9269 (N_9269,N_7200,N_7142);
nor U9270 (N_9270,N_6924,N_6849);
xnor U9271 (N_9271,N_7511,N_6308);
xnor U9272 (N_9272,N_6364,N_6159);
nand U9273 (N_9273,N_7021,N_6281);
or U9274 (N_9274,N_7264,N_7545);
nand U9275 (N_9275,N_6844,N_7833);
xor U9276 (N_9276,N_6886,N_7533);
nand U9277 (N_9277,N_7821,N_6089);
nand U9278 (N_9278,N_7311,N_7356);
nor U9279 (N_9279,N_7598,N_6114);
and U9280 (N_9280,N_7033,N_6405);
or U9281 (N_9281,N_7778,N_6915);
or U9282 (N_9282,N_7450,N_7226);
and U9283 (N_9283,N_6031,N_7966);
and U9284 (N_9284,N_6612,N_7569);
nor U9285 (N_9285,N_7039,N_7562);
xnor U9286 (N_9286,N_7237,N_7503);
nand U9287 (N_9287,N_7859,N_7484);
or U9288 (N_9288,N_7730,N_6697);
nor U9289 (N_9289,N_7691,N_6092);
or U9290 (N_9290,N_6514,N_7924);
or U9291 (N_9291,N_6458,N_6687);
and U9292 (N_9292,N_7960,N_7223);
or U9293 (N_9293,N_7060,N_7176);
nor U9294 (N_9294,N_7863,N_6221);
nand U9295 (N_9295,N_7161,N_6625);
nor U9296 (N_9296,N_6079,N_7602);
xor U9297 (N_9297,N_7061,N_7493);
nand U9298 (N_9298,N_6494,N_6640);
xor U9299 (N_9299,N_7884,N_7869);
and U9300 (N_9300,N_6408,N_6242);
or U9301 (N_9301,N_6937,N_7597);
nor U9302 (N_9302,N_6394,N_7919);
nor U9303 (N_9303,N_7686,N_6331);
and U9304 (N_9304,N_6502,N_6775);
nor U9305 (N_9305,N_7495,N_6556);
xor U9306 (N_9306,N_6337,N_7264);
nor U9307 (N_9307,N_6611,N_6147);
or U9308 (N_9308,N_6182,N_6491);
and U9309 (N_9309,N_6443,N_7339);
nand U9310 (N_9310,N_7925,N_6076);
xor U9311 (N_9311,N_7722,N_7198);
nor U9312 (N_9312,N_7287,N_6103);
xnor U9313 (N_9313,N_6176,N_7077);
nor U9314 (N_9314,N_7636,N_7985);
xor U9315 (N_9315,N_6946,N_6225);
or U9316 (N_9316,N_7729,N_6335);
nor U9317 (N_9317,N_7230,N_7810);
xor U9318 (N_9318,N_6973,N_6805);
or U9319 (N_9319,N_7758,N_7996);
nor U9320 (N_9320,N_6701,N_7385);
and U9321 (N_9321,N_7019,N_6084);
or U9322 (N_9322,N_6645,N_7635);
or U9323 (N_9323,N_7120,N_6365);
or U9324 (N_9324,N_6878,N_6571);
and U9325 (N_9325,N_6055,N_6948);
xnor U9326 (N_9326,N_6304,N_7899);
xor U9327 (N_9327,N_7025,N_7155);
xor U9328 (N_9328,N_6209,N_6933);
and U9329 (N_9329,N_6823,N_6626);
and U9330 (N_9330,N_7464,N_7864);
and U9331 (N_9331,N_7437,N_7995);
nor U9332 (N_9332,N_7163,N_7443);
or U9333 (N_9333,N_6749,N_7672);
nand U9334 (N_9334,N_7505,N_6325);
and U9335 (N_9335,N_7224,N_7542);
and U9336 (N_9336,N_7896,N_7253);
or U9337 (N_9337,N_6805,N_7191);
and U9338 (N_9338,N_7625,N_7575);
xnor U9339 (N_9339,N_7406,N_7426);
nand U9340 (N_9340,N_7950,N_6167);
xor U9341 (N_9341,N_7685,N_6849);
xnor U9342 (N_9342,N_7498,N_6996);
or U9343 (N_9343,N_7130,N_6173);
xor U9344 (N_9344,N_7882,N_7772);
xnor U9345 (N_9345,N_6457,N_6737);
or U9346 (N_9346,N_7296,N_7965);
xor U9347 (N_9347,N_7804,N_6222);
nor U9348 (N_9348,N_6956,N_6492);
nor U9349 (N_9349,N_6704,N_7030);
and U9350 (N_9350,N_7930,N_7446);
or U9351 (N_9351,N_6972,N_6076);
or U9352 (N_9352,N_7252,N_7703);
and U9353 (N_9353,N_7414,N_6826);
nand U9354 (N_9354,N_7681,N_7308);
and U9355 (N_9355,N_7745,N_7594);
nand U9356 (N_9356,N_7316,N_7026);
or U9357 (N_9357,N_6078,N_7462);
xor U9358 (N_9358,N_7092,N_7762);
and U9359 (N_9359,N_7865,N_7117);
nand U9360 (N_9360,N_6028,N_7858);
nor U9361 (N_9361,N_6915,N_6606);
nor U9362 (N_9362,N_7896,N_7249);
and U9363 (N_9363,N_7008,N_7726);
or U9364 (N_9364,N_7096,N_7493);
or U9365 (N_9365,N_6336,N_7741);
nand U9366 (N_9366,N_7331,N_6987);
nor U9367 (N_9367,N_7087,N_7104);
xnor U9368 (N_9368,N_7397,N_6249);
nor U9369 (N_9369,N_6261,N_6708);
and U9370 (N_9370,N_6068,N_6647);
or U9371 (N_9371,N_6350,N_7825);
or U9372 (N_9372,N_6406,N_6730);
and U9373 (N_9373,N_7937,N_7318);
xnor U9374 (N_9374,N_7395,N_6816);
nor U9375 (N_9375,N_7811,N_7587);
xor U9376 (N_9376,N_7750,N_6011);
and U9377 (N_9377,N_6529,N_7047);
nor U9378 (N_9378,N_6213,N_7511);
nand U9379 (N_9379,N_7030,N_7704);
nor U9380 (N_9380,N_6282,N_6742);
xor U9381 (N_9381,N_6633,N_7628);
and U9382 (N_9382,N_6813,N_6167);
and U9383 (N_9383,N_7293,N_6372);
or U9384 (N_9384,N_6143,N_7944);
nand U9385 (N_9385,N_7548,N_6664);
or U9386 (N_9386,N_7170,N_7555);
nand U9387 (N_9387,N_6705,N_6106);
nor U9388 (N_9388,N_6016,N_7387);
xor U9389 (N_9389,N_6119,N_6172);
or U9390 (N_9390,N_6947,N_6522);
nand U9391 (N_9391,N_7187,N_6132);
xnor U9392 (N_9392,N_6313,N_6062);
nand U9393 (N_9393,N_7505,N_7109);
or U9394 (N_9394,N_6742,N_7985);
or U9395 (N_9395,N_6981,N_6489);
nand U9396 (N_9396,N_6113,N_6162);
nand U9397 (N_9397,N_7118,N_7253);
and U9398 (N_9398,N_6017,N_7590);
or U9399 (N_9399,N_6569,N_6470);
and U9400 (N_9400,N_6395,N_6227);
and U9401 (N_9401,N_7256,N_7546);
nor U9402 (N_9402,N_6994,N_7762);
xnor U9403 (N_9403,N_6549,N_7170);
nand U9404 (N_9404,N_6356,N_6969);
nor U9405 (N_9405,N_6907,N_7227);
and U9406 (N_9406,N_7992,N_7586);
nand U9407 (N_9407,N_7272,N_6141);
xor U9408 (N_9408,N_7738,N_7214);
and U9409 (N_9409,N_7798,N_7849);
nor U9410 (N_9410,N_7251,N_6828);
or U9411 (N_9411,N_6593,N_6131);
and U9412 (N_9412,N_7058,N_6058);
nand U9413 (N_9413,N_7794,N_7420);
xor U9414 (N_9414,N_6040,N_6022);
and U9415 (N_9415,N_6824,N_6984);
xnor U9416 (N_9416,N_6341,N_6126);
nor U9417 (N_9417,N_7038,N_6324);
or U9418 (N_9418,N_7197,N_6463);
and U9419 (N_9419,N_6107,N_6883);
or U9420 (N_9420,N_7132,N_7957);
xnor U9421 (N_9421,N_6295,N_6062);
and U9422 (N_9422,N_6321,N_7613);
or U9423 (N_9423,N_7077,N_7790);
nor U9424 (N_9424,N_6749,N_6278);
nand U9425 (N_9425,N_7099,N_7979);
and U9426 (N_9426,N_7831,N_7711);
xor U9427 (N_9427,N_7800,N_6596);
and U9428 (N_9428,N_6217,N_7413);
xnor U9429 (N_9429,N_7663,N_7412);
or U9430 (N_9430,N_6167,N_6893);
and U9431 (N_9431,N_6468,N_7514);
nand U9432 (N_9432,N_6967,N_7241);
or U9433 (N_9433,N_7876,N_7499);
or U9434 (N_9434,N_7969,N_6613);
xor U9435 (N_9435,N_7087,N_6181);
or U9436 (N_9436,N_7446,N_6443);
xor U9437 (N_9437,N_7916,N_7561);
or U9438 (N_9438,N_7196,N_7937);
xor U9439 (N_9439,N_6129,N_7859);
and U9440 (N_9440,N_6037,N_6690);
xor U9441 (N_9441,N_6130,N_7670);
nor U9442 (N_9442,N_7644,N_6707);
nor U9443 (N_9443,N_7432,N_7560);
nand U9444 (N_9444,N_6770,N_6191);
or U9445 (N_9445,N_7029,N_6887);
or U9446 (N_9446,N_7015,N_7500);
xor U9447 (N_9447,N_7747,N_6495);
or U9448 (N_9448,N_6642,N_7333);
nand U9449 (N_9449,N_7568,N_7525);
or U9450 (N_9450,N_7449,N_7337);
nor U9451 (N_9451,N_6207,N_6976);
xor U9452 (N_9452,N_7810,N_6313);
and U9453 (N_9453,N_7534,N_6517);
xor U9454 (N_9454,N_6681,N_6650);
and U9455 (N_9455,N_6388,N_6547);
xor U9456 (N_9456,N_6738,N_7486);
nor U9457 (N_9457,N_6843,N_6916);
and U9458 (N_9458,N_6155,N_7517);
nor U9459 (N_9459,N_6720,N_7444);
or U9460 (N_9460,N_6280,N_7275);
xnor U9461 (N_9461,N_6724,N_6390);
nor U9462 (N_9462,N_7522,N_6073);
nor U9463 (N_9463,N_6147,N_6481);
and U9464 (N_9464,N_7835,N_6989);
or U9465 (N_9465,N_6500,N_7935);
nor U9466 (N_9466,N_7861,N_6064);
or U9467 (N_9467,N_7973,N_7500);
and U9468 (N_9468,N_6778,N_7684);
nand U9469 (N_9469,N_7526,N_6182);
nand U9470 (N_9470,N_7519,N_6508);
nor U9471 (N_9471,N_7212,N_6232);
nand U9472 (N_9472,N_7404,N_6828);
and U9473 (N_9473,N_7252,N_7337);
nor U9474 (N_9474,N_6486,N_6759);
and U9475 (N_9475,N_6087,N_7903);
or U9476 (N_9476,N_7804,N_7707);
xnor U9477 (N_9477,N_7156,N_6040);
xor U9478 (N_9478,N_6560,N_7994);
xnor U9479 (N_9479,N_6259,N_6834);
and U9480 (N_9480,N_7327,N_6805);
or U9481 (N_9481,N_6223,N_6903);
xor U9482 (N_9482,N_7621,N_7812);
or U9483 (N_9483,N_7788,N_6096);
or U9484 (N_9484,N_6138,N_6461);
xor U9485 (N_9485,N_6498,N_6513);
xnor U9486 (N_9486,N_7544,N_6811);
nor U9487 (N_9487,N_6763,N_7670);
xnor U9488 (N_9488,N_6080,N_7889);
or U9489 (N_9489,N_6163,N_7242);
xnor U9490 (N_9490,N_6911,N_7948);
or U9491 (N_9491,N_6338,N_6855);
and U9492 (N_9492,N_7697,N_7634);
nand U9493 (N_9493,N_6640,N_7669);
nand U9494 (N_9494,N_7441,N_7039);
and U9495 (N_9495,N_6737,N_7559);
or U9496 (N_9496,N_6930,N_6898);
or U9497 (N_9497,N_7365,N_7330);
and U9498 (N_9498,N_6178,N_7984);
nor U9499 (N_9499,N_6245,N_7127);
xor U9500 (N_9500,N_6344,N_6422);
or U9501 (N_9501,N_6510,N_7055);
nand U9502 (N_9502,N_7004,N_6179);
nand U9503 (N_9503,N_6226,N_7101);
and U9504 (N_9504,N_6736,N_7082);
xnor U9505 (N_9505,N_6735,N_6641);
nand U9506 (N_9506,N_7340,N_7785);
nor U9507 (N_9507,N_6293,N_7487);
nor U9508 (N_9508,N_7624,N_7582);
and U9509 (N_9509,N_6038,N_6824);
xnor U9510 (N_9510,N_6434,N_6757);
nand U9511 (N_9511,N_7653,N_7463);
xor U9512 (N_9512,N_6661,N_6836);
nor U9513 (N_9513,N_6679,N_7484);
xor U9514 (N_9514,N_6603,N_6009);
and U9515 (N_9515,N_6324,N_6996);
nor U9516 (N_9516,N_7409,N_7961);
nand U9517 (N_9517,N_6891,N_6480);
or U9518 (N_9518,N_7092,N_7938);
xnor U9519 (N_9519,N_6513,N_6543);
nor U9520 (N_9520,N_7227,N_7980);
and U9521 (N_9521,N_6306,N_7528);
nand U9522 (N_9522,N_6653,N_7058);
nand U9523 (N_9523,N_7657,N_6465);
and U9524 (N_9524,N_7733,N_7768);
nor U9525 (N_9525,N_7521,N_7762);
and U9526 (N_9526,N_7655,N_7937);
and U9527 (N_9527,N_7728,N_7817);
or U9528 (N_9528,N_6547,N_7885);
nand U9529 (N_9529,N_7460,N_7457);
xnor U9530 (N_9530,N_6328,N_7543);
nand U9531 (N_9531,N_7419,N_6824);
nor U9532 (N_9532,N_7659,N_6249);
xor U9533 (N_9533,N_7488,N_6878);
xnor U9534 (N_9534,N_7726,N_6214);
or U9535 (N_9535,N_7668,N_6876);
nand U9536 (N_9536,N_6997,N_7162);
nand U9537 (N_9537,N_7378,N_7881);
xor U9538 (N_9538,N_7216,N_7239);
nor U9539 (N_9539,N_7325,N_6275);
xor U9540 (N_9540,N_6832,N_7054);
xor U9541 (N_9541,N_7042,N_6671);
nand U9542 (N_9542,N_7693,N_7299);
or U9543 (N_9543,N_7343,N_7511);
xnor U9544 (N_9544,N_7513,N_6449);
or U9545 (N_9545,N_7857,N_7934);
nand U9546 (N_9546,N_7828,N_7430);
nor U9547 (N_9547,N_6893,N_6503);
nand U9548 (N_9548,N_6753,N_6958);
nand U9549 (N_9549,N_7763,N_7779);
nor U9550 (N_9550,N_7565,N_6516);
xnor U9551 (N_9551,N_7611,N_6947);
and U9552 (N_9552,N_7438,N_6977);
nand U9553 (N_9553,N_6080,N_7826);
or U9554 (N_9554,N_6138,N_6984);
and U9555 (N_9555,N_7122,N_7435);
xor U9556 (N_9556,N_7321,N_6653);
nand U9557 (N_9557,N_6942,N_7269);
and U9558 (N_9558,N_6985,N_7216);
nand U9559 (N_9559,N_7105,N_6682);
or U9560 (N_9560,N_6620,N_6769);
and U9561 (N_9561,N_6705,N_6860);
xnor U9562 (N_9562,N_7209,N_6908);
or U9563 (N_9563,N_6062,N_6672);
nor U9564 (N_9564,N_6739,N_7974);
nand U9565 (N_9565,N_7182,N_7081);
xnor U9566 (N_9566,N_7895,N_7371);
xnor U9567 (N_9567,N_6589,N_7141);
nor U9568 (N_9568,N_7991,N_6157);
nand U9569 (N_9569,N_6814,N_6407);
or U9570 (N_9570,N_6572,N_6804);
nand U9571 (N_9571,N_6363,N_6273);
nor U9572 (N_9572,N_7068,N_6338);
nand U9573 (N_9573,N_6753,N_6285);
or U9574 (N_9574,N_7181,N_7447);
nand U9575 (N_9575,N_7281,N_6240);
nand U9576 (N_9576,N_6696,N_7845);
xnor U9577 (N_9577,N_6526,N_7923);
xnor U9578 (N_9578,N_7661,N_7833);
nor U9579 (N_9579,N_7179,N_7832);
nand U9580 (N_9580,N_6989,N_6747);
nand U9581 (N_9581,N_7788,N_6508);
nor U9582 (N_9582,N_6344,N_6637);
and U9583 (N_9583,N_6023,N_6102);
and U9584 (N_9584,N_6603,N_7553);
nor U9585 (N_9585,N_6885,N_7908);
nand U9586 (N_9586,N_7966,N_6137);
and U9587 (N_9587,N_6997,N_6419);
nor U9588 (N_9588,N_7769,N_7882);
xnor U9589 (N_9589,N_6801,N_7807);
or U9590 (N_9590,N_7370,N_7423);
nor U9591 (N_9591,N_6950,N_6304);
or U9592 (N_9592,N_7806,N_7581);
and U9593 (N_9593,N_7562,N_6653);
and U9594 (N_9594,N_6683,N_6240);
nand U9595 (N_9595,N_7052,N_6216);
and U9596 (N_9596,N_7550,N_7261);
or U9597 (N_9597,N_7193,N_6829);
or U9598 (N_9598,N_6541,N_6429);
nor U9599 (N_9599,N_6261,N_7687);
nor U9600 (N_9600,N_7702,N_7853);
xnor U9601 (N_9601,N_7194,N_7308);
xor U9602 (N_9602,N_6298,N_6106);
xor U9603 (N_9603,N_7982,N_6030);
or U9604 (N_9604,N_7573,N_7791);
nand U9605 (N_9605,N_6358,N_6353);
nor U9606 (N_9606,N_7173,N_6419);
or U9607 (N_9607,N_6575,N_6849);
nand U9608 (N_9608,N_7565,N_7487);
or U9609 (N_9609,N_6804,N_7716);
xnor U9610 (N_9610,N_7636,N_6484);
xnor U9611 (N_9611,N_7324,N_6759);
xnor U9612 (N_9612,N_7621,N_7316);
nand U9613 (N_9613,N_7322,N_7659);
nor U9614 (N_9614,N_6089,N_6600);
xnor U9615 (N_9615,N_6216,N_7776);
nor U9616 (N_9616,N_6105,N_7037);
xnor U9617 (N_9617,N_7000,N_7905);
xor U9618 (N_9618,N_6239,N_7621);
xnor U9619 (N_9619,N_6128,N_7430);
nand U9620 (N_9620,N_7271,N_6672);
or U9621 (N_9621,N_7635,N_6206);
and U9622 (N_9622,N_6877,N_6508);
nor U9623 (N_9623,N_6673,N_7922);
or U9624 (N_9624,N_7889,N_6567);
nor U9625 (N_9625,N_6200,N_7691);
and U9626 (N_9626,N_7903,N_6660);
nand U9627 (N_9627,N_6520,N_6063);
and U9628 (N_9628,N_6051,N_7832);
nor U9629 (N_9629,N_7687,N_7352);
nor U9630 (N_9630,N_7040,N_6655);
or U9631 (N_9631,N_6402,N_7682);
and U9632 (N_9632,N_7015,N_6904);
and U9633 (N_9633,N_7926,N_6452);
and U9634 (N_9634,N_6319,N_6337);
and U9635 (N_9635,N_6785,N_6317);
or U9636 (N_9636,N_7856,N_6871);
nor U9637 (N_9637,N_6227,N_7314);
nand U9638 (N_9638,N_7058,N_6071);
or U9639 (N_9639,N_6007,N_6689);
xor U9640 (N_9640,N_6723,N_6380);
nor U9641 (N_9641,N_7909,N_6013);
nand U9642 (N_9642,N_7902,N_7392);
and U9643 (N_9643,N_7435,N_7987);
nand U9644 (N_9644,N_7454,N_6385);
nand U9645 (N_9645,N_7430,N_7238);
nand U9646 (N_9646,N_6343,N_6533);
and U9647 (N_9647,N_6875,N_7321);
or U9648 (N_9648,N_6178,N_6796);
xor U9649 (N_9649,N_6992,N_6911);
or U9650 (N_9650,N_7761,N_6760);
nand U9651 (N_9651,N_7648,N_7547);
or U9652 (N_9652,N_6721,N_7834);
xor U9653 (N_9653,N_6623,N_7166);
and U9654 (N_9654,N_6104,N_6578);
or U9655 (N_9655,N_6815,N_7702);
nand U9656 (N_9656,N_6500,N_6146);
xnor U9657 (N_9657,N_7918,N_6356);
nand U9658 (N_9658,N_7635,N_7175);
xnor U9659 (N_9659,N_6058,N_7862);
nand U9660 (N_9660,N_6032,N_7265);
nor U9661 (N_9661,N_7030,N_7289);
nand U9662 (N_9662,N_6746,N_6179);
nand U9663 (N_9663,N_6681,N_7181);
nor U9664 (N_9664,N_7184,N_6841);
nand U9665 (N_9665,N_7714,N_7704);
nand U9666 (N_9666,N_7699,N_7657);
nor U9667 (N_9667,N_6388,N_6057);
and U9668 (N_9668,N_6978,N_7049);
and U9669 (N_9669,N_6612,N_7606);
and U9670 (N_9670,N_7599,N_7911);
nor U9671 (N_9671,N_7157,N_7295);
or U9672 (N_9672,N_6497,N_6065);
and U9673 (N_9673,N_6772,N_7681);
or U9674 (N_9674,N_7883,N_7998);
xnor U9675 (N_9675,N_6418,N_6039);
xor U9676 (N_9676,N_6035,N_7523);
xor U9677 (N_9677,N_7987,N_7932);
and U9678 (N_9678,N_7599,N_7130);
xor U9679 (N_9679,N_7077,N_6882);
or U9680 (N_9680,N_6346,N_6663);
and U9681 (N_9681,N_7925,N_7795);
and U9682 (N_9682,N_7073,N_7233);
nor U9683 (N_9683,N_6691,N_6323);
nor U9684 (N_9684,N_7420,N_7659);
nor U9685 (N_9685,N_7315,N_7407);
and U9686 (N_9686,N_7207,N_7464);
xor U9687 (N_9687,N_6873,N_7984);
nand U9688 (N_9688,N_7665,N_7334);
or U9689 (N_9689,N_7950,N_7843);
and U9690 (N_9690,N_6704,N_6275);
xnor U9691 (N_9691,N_6705,N_6579);
xnor U9692 (N_9692,N_7520,N_7874);
xnor U9693 (N_9693,N_7127,N_7468);
nand U9694 (N_9694,N_6994,N_7646);
nand U9695 (N_9695,N_7520,N_6941);
xnor U9696 (N_9696,N_6393,N_6623);
xnor U9697 (N_9697,N_6356,N_7406);
xor U9698 (N_9698,N_7643,N_6565);
nor U9699 (N_9699,N_7242,N_6031);
nand U9700 (N_9700,N_7301,N_7009);
xor U9701 (N_9701,N_6836,N_6704);
or U9702 (N_9702,N_6385,N_7474);
nor U9703 (N_9703,N_6297,N_6934);
xnor U9704 (N_9704,N_6506,N_7979);
xnor U9705 (N_9705,N_7284,N_7815);
or U9706 (N_9706,N_7101,N_6297);
nand U9707 (N_9707,N_6430,N_7887);
xnor U9708 (N_9708,N_6662,N_6509);
and U9709 (N_9709,N_6348,N_6976);
nor U9710 (N_9710,N_6815,N_7279);
nand U9711 (N_9711,N_7427,N_7059);
and U9712 (N_9712,N_6694,N_6727);
or U9713 (N_9713,N_6136,N_7534);
nor U9714 (N_9714,N_7122,N_6401);
nand U9715 (N_9715,N_7375,N_6990);
nor U9716 (N_9716,N_7524,N_6454);
and U9717 (N_9717,N_6873,N_6817);
nand U9718 (N_9718,N_7437,N_6720);
or U9719 (N_9719,N_7798,N_6839);
or U9720 (N_9720,N_6751,N_7877);
nor U9721 (N_9721,N_6511,N_6194);
nand U9722 (N_9722,N_7984,N_7444);
and U9723 (N_9723,N_6795,N_6753);
or U9724 (N_9724,N_6418,N_6898);
and U9725 (N_9725,N_7311,N_6274);
and U9726 (N_9726,N_7213,N_7183);
nand U9727 (N_9727,N_7013,N_7448);
nor U9728 (N_9728,N_6721,N_6716);
nor U9729 (N_9729,N_7191,N_7505);
and U9730 (N_9730,N_6009,N_6643);
nor U9731 (N_9731,N_7318,N_6173);
nand U9732 (N_9732,N_6868,N_6970);
xnor U9733 (N_9733,N_6173,N_6730);
xor U9734 (N_9734,N_6194,N_7335);
or U9735 (N_9735,N_7951,N_6003);
xor U9736 (N_9736,N_6320,N_7343);
xor U9737 (N_9737,N_7749,N_7012);
nor U9738 (N_9738,N_6614,N_7774);
nand U9739 (N_9739,N_7057,N_6892);
nand U9740 (N_9740,N_7458,N_7520);
or U9741 (N_9741,N_6496,N_7362);
and U9742 (N_9742,N_6465,N_7554);
nand U9743 (N_9743,N_7264,N_6059);
and U9744 (N_9744,N_6093,N_6271);
nor U9745 (N_9745,N_6703,N_6084);
nand U9746 (N_9746,N_6091,N_6123);
and U9747 (N_9747,N_7689,N_6911);
nand U9748 (N_9748,N_6336,N_6793);
nor U9749 (N_9749,N_6712,N_7082);
xor U9750 (N_9750,N_7667,N_6126);
or U9751 (N_9751,N_6789,N_6756);
nand U9752 (N_9752,N_6543,N_6510);
and U9753 (N_9753,N_7583,N_7017);
and U9754 (N_9754,N_7633,N_7748);
or U9755 (N_9755,N_7234,N_7638);
or U9756 (N_9756,N_7765,N_7737);
nor U9757 (N_9757,N_6814,N_6881);
xor U9758 (N_9758,N_7330,N_6140);
or U9759 (N_9759,N_6773,N_6817);
and U9760 (N_9760,N_7278,N_7888);
and U9761 (N_9761,N_6054,N_7651);
or U9762 (N_9762,N_6387,N_6249);
and U9763 (N_9763,N_7630,N_7514);
and U9764 (N_9764,N_7274,N_7636);
and U9765 (N_9765,N_6299,N_6410);
nand U9766 (N_9766,N_7269,N_7625);
and U9767 (N_9767,N_6745,N_7476);
nor U9768 (N_9768,N_7631,N_6196);
or U9769 (N_9769,N_7171,N_6527);
or U9770 (N_9770,N_6935,N_6823);
and U9771 (N_9771,N_7362,N_7421);
nor U9772 (N_9772,N_6814,N_7477);
or U9773 (N_9773,N_7631,N_7075);
xor U9774 (N_9774,N_7424,N_7441);
or U9775 (N_9775,N_7474,N_7845);
xor U9776 (N_9776,N_7633,N_6658);
and U9777 (N_9777,N_6429,N_6844);
or U9778 (N_9778,N_7048,N_6717);
xnor U9779 (N_9779,N_7829,N_6237);
nand U9780 (N_9780,N_6215,N_6476);
xor U9781 (N_9781,N_7010,N_6872);
or U9782 (N_9782,N_7264,N_7095);
nor U9783 (N_9783,N_6260,N_7317);
xnor U9784 (N_9784,N_6671,N_7588);
nand U9785 (N_9785,N_7217,N_6982);
nor U9786 (N_9786,N_7306,N_6299);
xor U9787 (N_9787,N_6032,N_7948);
xor U9788 (N_9788,N_7748,N_6053);
nor U9789 (N_9789,N_7390,N_7714);
xor U9790 (N_9790,N_6945,N_6775);
or U9791 (N_9791,N_7321,N_6052);
nand U9792 (N_9792,N_6660,N_6053);
nor U9793 (N_9793,N_6647,N_6055);
nand U9794 (N_9794,N_7579,N_6071);
xnor U9795 (N_9795,N_7868,N_7765);
and U9796 (N_9796,N_6594,N_6709);
and U9797 (N_9797,N_7247,N_7000);
and U9798 (N_9798,N_7563,N_7305);
or U9799 (N_9799,N_6243,N_6769);
or U9800 (N_9800,N_7326,N_6583);
nand U9801 (N_9801,N_6437,N_7083);
nor U9802 (N_9802,N_7769,N_7285);
or U9803 (N_9803,N_6857,N_6380);
nor U9804 (N_9804,N_7154,N_7084);
or U9805 (N_9805,N_6429,N_7856);
and U9806 (N_9806,N_6294,N_6904);
nor U9807 (N_9807,N_6584,N_6919);
and U9808 (N_9808,N_7507,N_7438);
xnor U9809 (N_9809,N_6338,N_6558);
xor U9810 (N_9810,N_7261,N_7064);
or U9811 (N_9811,N_7417,N_6443);
xor U9812 (N_9812,N_6730,N_7526);
nand U9813 (N_9813,N_7046,N_6062);
nor U9814 (N_9814,N_6945,N_7106);
xnor U9815 (N_9815,N_6548,N_7127);
xnor U9816 (N_9816,N_6228,N_6361);
nor U9817 (N_9817,N_7461,N_6406);
or U9818 (N_9818,N_6107,N_6586);
xor U9819 (N_9819,N_7672,N_6693);
nand U9820 (N_9820,N_6071,N_6949);
nor U9821 (N_9821,N_6921,N_6578);
and U9822 (N_9822,N_7649,N_6742);
xor U9823 (N_9823,N_7735,N_7458);
nand U9824 (N_9824,N_7828,N_6896);
nor U9825 (N_9825,N_7445,N_7870);
xor U9826 (N_9826,N_6158,N_6682);
xnor U9827 (N_9827,N_7623,N_6173);
or U9828 (N_9828,N_7721,N_7206);
or U9829 (N_9829,N_7441,N_7745);
or U9830 (N_9830,N_6003,N_7360);
nand U9831 (N_9831,N_6464,N_6110);
or U9832 (N_9832,N_7817,N_6143);
xor U9833 (N_9833,N_7299,N_7811);
or U9834 (N_9834,N_6632,N_6239);
and U9835 (N_9835,N_6616,N_6901);
xor U9836 (N_9836,N_7674,N_7853);
nor U9837 (N_9837,N_7188,N_7151);
and U9838 (N_9838,N_7124,N_7505);
xnor U9839 (N_9839,N_6319,N_6600);
xor U9840 (N_9840,N_6738,N_6564);
or U9841 (N_9841,N_6671,N_7786);
xor U9842 (N_9842,N_6293,N_6987);
nand U9843 (N_9843,N_7703,N_7341);
nor U9844 (N_9844,N_6805,N_6530);
or U9845 (N_9845,N_7292,N_7831);
nand U9846 (N_9846,N_6077,N_6222);
and U9847 (N_9847,N_6356,N_7156);
xor U9848 (N_9848,N_6935,N_6051);
or U9849 (N_9849,N_6375,N_6455);
or U9850 (N_9850,N_7669,N_6891);
xnor U9851 (N_9851,N_7049,N_7703);
nor U9852 (N_9852,N_6044,N_6907);
or U9853 (N_9853,N_6898,N_7876);
and U9854 (N_9854,N_6162,N_7765);
nor U9855 (N_9855,N_6417,N_6749);
or U9856 (N_9856,N_6301,N_7240);
nor U9857 (N_9857,N_7433,N_7183);
nand U9858 (N_9858,N_6668,N_6321);
or U9859 (N_9859,N_7520,N_6478);
xnor U9860 (N_9860,N_6597,N_6181);
nor U9861 (N_9861,N_6769,N_7893);
and U9862 (N_9862,N_6465,N_6063);
and U9863 (N_9863,N_6301,N_6789);
nor U9864 (N_9864,N_7184,N_6915);
xnor U9865 (N_9865,N_7575,N_7470);
and U9866 (N_9866,N_6969,N_6269);
and U9867 (N_9867,N_6488,N_7464);
nand U9868 (N_9868,N_7409,N_7807);
xor U9869 (N_9869,N_7717,N_6729);
xnor U9870 (N_9870,N_6566,N_6644);
or U9871 (N_9871,N_7587,N_6526);
nor U9872 (N_9872,N_7948,N_6547);
xor U9873 (N_9873,N_6023,N_6877);
nor U9874 (N_9874,N_7636,N_7501);
and U9875 (N_9875,N_6715,N_6857);
and U9876 (N_9876,N_7124,N_7330);
nand U9877 (N_9877,N_7118,N_6482);
or U9878 (N_9878,N_6330,N_7729);
nor U9879 (N_9879,N_6852,N_7447);
and U9880 (N_9880,N_7119,N_6452);
nand U9881 (N_9881,N_7636,N_7572);
xor U9882 (N_9882,N_7137,N_7811);
or U9883 (N_9883,N_6485,N_7081);
xnor U9884 (N_9884,N_7309,N_7989);
xor U9885 (N_9885,N_6291,N_6702);
xor U9886 (N_9886,N_6451,N_7770);
and U9887 (N_9887,N_7023,N_7643);
xor U9888 (N_9888,N_6724,N_7155);
nor U9889 (N_9889,N_7046,N_7950);
nor U9890 (N_9890,N_7384,N_7825);
or U9891 (N_9891,N_7792,N_7609);
nand U9892 (N_9892,N_7450,N_7816);
xor U9893 (N_9893,N_6936,N_7592);
nand U9894 (N_9894,N_7692,N_6692);
nor U9895 (N_9895,N_7964,N_7509);
nor U9896 (N_9896,N_6185,N_6108);
nand U9897 (N_9897,N_7830,N_6959);
nor U9898 (N_9898,N_6027,N_7141);
nand U9899 (N_9899,N_6511,N_6198);
and U9900 (N_9900,N_6053,N_6849);
nand U9901 (N_9901,N_6201,N_6812);
xnor U9902 (N_9902,N_7762,N_6326);
or U9903 (N_9903,N_6217,N_7432);
or U9904 (N_9904,N_7048,N_7657);
or U9905 (N_9905,N_6624,N_6796);
nor U9906 (N_9906,N_6404,N_7655);
nor U9907 (N_9907,N_7148,N_7904);
xor U9908 (N_9908,N_7452,N_6245);
nand U9909 (N_9909,N_6017,N_6678);
nand U9910 (N_9910,N_6480,N_6049);
xor U9911 (N_9911,N_7691,N_7844);
and U9912 (N_9912,N_7856,N_7916);
and U9913 (N_9913,N_6519,N_7587);
xnor U9914 (N_9914,N_7434,N_7365);
nand U9915 (N_9915,N_6173,N_7759);
xor U9916 (N_9916,N_6613,N_6095);
xor U9917 (N_9917,N_7409,N_6169);
nor U9918 (N_9918,N_7757,N_7828);
xnor U9919 (N_9919,N_6169,N_6805);
nor U9920 (N_9920,N_7381,N_7982);
xor U9921 (N_9921,N_7495,N_7970);
nor U9922 (N_9922,N_7575,N_6895);
and U9923 (N_9923,N_6851,N_7261);
nand U9924 (N_9924,N_7664,N_6555);
and U9925 (N_9925,N_7886,N_7599);
and U9926 (N_9926,N_6802,N_7649);
xor U9927 (N_9927,N_7965,N_7947);
xor U9928 (N_9928,N_6533,N_7484);
nand U9929 (N_9929,N_7243,N_7709);
nand U9930 (N_9930,N_6381,N_7606);
nor U9931 (N_9931,N_7673,N_7219);
nor U9932 (N_9932,N_7744,N_6142);
or U9933 (N_9933,N_7183,N_7933);
nor U9934 (N_9934,N_7065,N_6392);
or U9935 (N_9935,N_7115,N_6920);
nand U9936 (N_9936,N_6566,N_6311);
nor U9937 (N_9937,N_6514,N_7681);
xor U9938 (N_9938,N_6461,N_6941);
or U9939 (N_9939,N_7369,N_6559);
nor U9940 (N_9940,N_7211,N_7769);
nor U9941 (N_9941,N_6447,N_7294);
nand U9942 (N_9942,N_7933,N_7884);
xnor U9943 (N_9943,N_7909,N_7923);
nand U9944 (N_9944,N_7173,N_6922);
or U9945 (N_9945,N_7853,N_6776);
and U9946 (N_9946,N_7039,N_7507);
nand U9947 (N_9947,N_6386,N_7023);
xnor U9948 (N_9948,N_6351,N_7836);
nand U9949 (N_9949,N_7257,N_7224);
and U9950 (N_9950,N_7455,N_7394);
and U9951 (N_9951,N_7080,N_7647);
nor U9952 (N_9952,N_6013,N_7171);
and U9953 (N_9953,N_6195,N_6473);
nor U9954 (N_9954,N_6053,N_6021);
nor U9955 (N_9955,N_7438,N_6318);
nand U9956 (N_9956,N_6630,N_6156);
nand U9957 (N_9957,N_7595,N_7448);
or U9958 (N_9958,N_6472,N_7284);
nor U9959 (N_9959,N_6212,N_6581);
nand U9960 (N_9960,N_6693,N_6687);
nor U9961 (N_9961,N_6792,N_6347);
xnor U9962 (N_9962,N_6086,N_7523);
and U9963 (N_9963,N_7233,N_7816);
xor U9964 (N_9964,N_7159,N_7803);
and U9965 (N_9965,N_7634,N_7930);
and U9966 (N_9966,N_7974,N_7179);
and U9967 (N_9967,N_6995,N_6782);
nand U9968 (N_9968,N_7656,N_6518);
xnor U9969 (N_9969,N_6087,N_7174);
and U9970 (N_9970,N_6956,N_7070);
and U9971 (N_9971,N_7099,N_7708);
or U9972 (N_9972,N_6820,N_6319);
and U9973 (N_9973,N_6578,N_7121);
or U9974 (N_9974,N_7051,N_7733);
or U9975 (N_9975,N_7908,N_6251);
nand U9976 (N_9976,N_7143,N_6674);
nand U9977 (N_9977,N_6355,N_7446);
nand U9978 (N_9978,N_7516,N_6382);
or U9979 (N_9979,N_7677,N_6002);
or U9980 (N_9980,N_6349,N_7493);
or U9981 (N_9981,N_7276,N_7271);
and U9982 (N_9982,N_6933,N_6494);
nor U9983 (N_9983,N_6112,N_6300);
nor U9984 (N_9984,N_7451,N_7755);
nor U9985 (N_9985,N_7548,N_7810);
or U9986 (N_9986,N_6436,N_7635);
or U9987 (N_9987,N_7763,N_7813);
xnor U9988 (N_9988,N_6896,N_6729);
xnor U9989 (N_9989,N_6603,N_6011);
and U9990 (N_9990,N_7857,N_7952);
xor U9991 (N_9991,N_7963,N_6063);
or U9992 (N_9992,N_7314,N_7039);
nand U9993 (N_9993,N_7137,N_6980);
nor U9994 (N_9994,N_6047,N_7741);
nor U9995 (N_9995,N_6031,N_7035);
or U9996 (N_9996,N_6325,N_6227);
nand U9997 (N_9997,N_7495,N_7583);
and U9998 (N_9998,N_7179,N_7567);
and U9999 (N_9999,N_6600,N_6608);
xor UO_0 (O_0,N_9357,N_8324);
and UO_1 (O_1,N_8927,N_9434);
nor UO_2 (O_2,N_9541,N_9078);
xor UO_3 (O_3,N_9897,N_9909);
or UO_4 (O_4,N_9620,N_8827);
or UO_5 (O_5,N_8181,N_8501);
xnor UO_6 (O_6,N_8071,N_9458);
nand UO_7 (O_7,N_8303,N_8460);
or UO_8 (O_8,N_8268,N_8540);
xnor UO_9 (O_9,N_9067,N_8241);
nand UO_10 (O_10,N_9930,N_9091);
nand UO_11 (O_11,N_8760,N_9614);
nand UO_12 (O_12,N_9532,N_9638);
nand UO_13 (O_13,N_9422,N_8140);
nand UO_14 (O_14,N_9608,N_9831);
or UO_15 (O_15,N_9315,N_8750);
or UO_16 (O_16,N_9330,N_8444);
or UO_17 (O_17,N_9157,N_8811);
nor UO_18 (O_18,N_8189,N_9153);
or UO_19 (O_19,N_8023,N_8002);
nor UO_20 (O_20,N_8193,N_9943);
and UO_21 (O_21,N_8840,N_9632);
nand UO_22 (O_22,N_9810,N_9832);
and UO_23 (O_23,N_9347,N_8228);
xnor UO_24 (O_24,N_9631,N_9507);
xnor UO_25 (O_25,N_9471,N_9130);
nor UO_26 (O_26,N_9323,N_9158);
nand UO_27 (O_27,N_9010,N_9031);
or UO_28 (O_28,N_9421,N_9318);
xor UO_29 (O_29,N_8367,N_9990);
nand UO_30 (O_30,N_9363,N_8706);
xor UO_31 (O_31,N_9871,N_9705);
or UO_32 (O_32,N_8877,N_8828);
nor UO_33 (O_33,N_9436,N_8157);
nor UO_34 (O_34,N_8244,N_8031);
xor UO_35 (O_35,N_9531,N_8653);
xor UO_36 (O_36,N_9259,N_9023);
nor UO_37 (O_37,N_9284,N_9512);
nor UO_38 (O_38,N_9971,N_8350);
xnor UO_39 (O_39,N_9992,N_8547);
or UO_40 (O_40,N_8217,N_8930);
nand UO_41 (O_41,N_8083,N_9246);
xnor UO_42 (O_42,N_9178,N_8705);
and UO_43 (O_43,N_9090,N_8110);
xnor UO_44 (O_44,N_8732,N_9723);
or UO_45 (O_45,N_8542,N_9216);
or UO_46 (O_46,N_8022,N_9661);
nor UO_47 (O_47,N_8159,N_8512);
and UO_48 (O_48,N_9503,N_9406);
xor UO_49 (O_49,N_9752,N_8937);
or UO_50 (O_50,N_8068,N_8533);
or UO_51 (O_51,N_9081,N_8014);
nand UO_52 (O_52,N_8650,N_9762);
nor UO_53 (O_53,N_8139,N_8858);
xnor UO_54 (O_54,N_9309,N_9355);
nand UO_55 (O_55,N_8282,N_9188);
and UO_56 (O_56,N_9869,N_9559);
nor UO_57 (O_57,N_8514,N_9305);
and UO_58 (O_58,N_9163,N_8972);
and UO_59 (O_59,N_8506,N_8669);
or UO_60 (O_60,N_8882,N_9497);
nor UO_61 (O_61,N_9999,N_8919);
and UO_62 (O_62,N_9120,N_9449);
nor UO_63 (O_63,N_8346,N_9367);
xor UO_64 (O_64,N_8341,N_8856);
and UO_65 (O_65,N_9229,N_9402);
xnor UO_66 (O_66,N_8935,N_8605);
xnor UO_67 (O_67,N_8142,N_8690);
nand UO_68 (O_68,N_8988,N_8236);
nor UO_69 (O_69,N_8621,N_9485);
xor UO_70 (O_70,N_8318,N_8826);
nor UO_71 (O_71,N_8920,N_9852);
and UO_72 (O_72,N_9779,N_8450);
or UO_73 (O_73,N_9230,N_8312);
and UO_74 (O_74,N_9365,N_9272);
and UO_75 (O_75,N_8046,N_8242);
xor UO_76 (O_76,N_8073,N_8006);
and UO_77 (O_77,N_9283,N_9797);
xnor UO_78 (O_78,N_9165,N_9772);
and UO_79 (O_79,N_9009,N_8399);
nor UO_80 (O_80,N_9635,N_9933);
nand UO_81 (O_81,N_9949,N_8195);
nor UO_82 (O_82,N_8513,N_8360);
and UO_83 (O_83,N_8797,N_8757);
xor UO_84 (O_84,N_8825,N_8135);
or UO_85 (O_85,N_9711,N_8850);
xnor UO_86 (O_86,N_9533,N_9214);
nand UO_87 (O_87,N_8573,N_8932);
and UO_88 (O_88,N_8597,N_9170);
xnor UO_89 (O_89,N_8560,N_8429);
xor UO_90 (O_90,N_8394,N_8072);
or UO_91 (O_91,N_8986,N_9702);
xnor UO_92 (O_92,N_8577,N_9416);
nand UO_93 (O_93,N_9277,N_9006);
xor UO_94 (O_94,N_9961,N_8194);
nand UO_95 (O_95,N_9149,N_9645);
and UO_96 (O_96,N_9469,N_8043);
or UO_97 (O_97,N_8611,N_8373);
nor UO_98 (O_98,N_9053,N_9922);
xor UO_99 (O_99,N_9247,N_9407);
nor UO_100 (O_100,N_9144,N_9640);
and UO_101 (O_101,N_9328,N_9475);
nand UO_102 (O_102,N_8285,N_9110);
or UO_103 (O_103,N_9627,N_8051);
xor UO_104 (O_104,N_8531,N_9254);
and UO_105 (O_105,N_9058,N_9231);
or UO_106 (O_106,N_8326,N_9744);
xnor UO_107 (O_107,N_8032,N_8302);
and UO_108 (O_108,N_8205,N_9528);
xor UO_109 (O_109,N_8586,N_8117);
and UO_110 (O_110,N_8048,N_8267);
or UO_111 (O_111,N_9108,N_8275);
xor UO_112 (O_112,N_9420,N_8461);
xor UO_113 (O_113,N_8163,N_9213);
or UO_114 (O_114,N_9886,N_9984);
and UO_115 (O_115,N_9268,N_9221);
nor UO_116 (O_116,N_9515,N_9974);
or UO_117 (O_117,N_9798,N_9666);
or UO_118 (O_118,N_8146,N_9823);
xor UO_119 (O_119,N_9651,N_9036);
and UO_120 (O_120,N_9862,N_9065);
or UO_121 (O_121,N_8876,N_8299);
and UO_122 (O_122,N_9432,N_9607);
or UO_123 (O_123,N_9498,N_8094);
nor UO_124 (O_124,N_9524,N_9735);
nor UO_125 (O_125,N_8295,N_9673);
nor UO_126 (O_126,N_9424,N_8941);
or UO_127 (O_127,N_9579,N_9682);
xor UO_128 (O_128,N_8013,N_9615);
nor UO_129 (O_129,N_9311,N_9479);
nand UO_130 (O_130,N_9902,N_9000);
and UO_131 (O_131,N_8539,N_8996);
nand UO_132 (O_132,N_9914,N_9547);
or UO_133 (O_133,N_8761,N_9415);
or UO_134 (O_134,N_8216,N_9942);
or UO_135 (O_135,N_8891,N_9398);
nand UO_136 (O_136,N_9346,N_8132);
nand UO_137 (O_137,N_8630,N_9709);
and UO_138 (O_138,N_9513,N_8477);
nor UO_139 (O_139,N_8585,N_9546);
nand UO_140 (O_140,N_9394,N_8736);
or UO_141 (O_141,N_9098,N_8622);
nand UO_142 (O_142,N_8136,N_8917);
or UO_143 (O_143,N_8535,N_8390);
nand UO_144 (O_144,N_8247,N_9835);
and UO_145 (O_145,N_8728,N_8860);
xnor UO_146 (O_146,N_9390,N_9552);
or UO_147 (O_147,N_8028,N_8454);
and UO_148 (O_148,N_9655,N_9456);
and UO_149 (O_149,N_9099,N_8400);
or UO_150 (O_150,N_8847,N_9982);
xnor UO_151 (O_151,N_8519,N_8204);
or UO_152 (O_152,N_8016,N_9019);
nor UO_153 (O_153,N_9803,N_8198);
xor UO_154 (O_154,N_8832,N_8620);
and UO_155 (O_155,N_8614,N_9240);
or UO_156 (O_156,N_8026,N_9013);
nand UO_157 (O_157,N_8162,N_8809);
and UO_158 (O_158,N_9501,N_8306);
and UO_159 (O_159,N_9804,N_8122);
and UO_160 (O_160,N_8594,N_9731);
xnor UO_161 (O_161,N_8700,N_9795);
xnor UO_162 (O_162,N_9440,N_8387);
nor UO_163 (O_163,N_9257,N_9491);
nand UO_164 (O_164,N_9874,N_8018);
xnor UO_165 (O_165,N_8381,N_8419);
nand UO_166 (O_166,N_8829,N_9083);
nand UO_167 (O_167,N_9410,N_8721);
xnor UO_168 (O_168,N_9605,N_8724);
and UO_169 (O_169,N_8409,N_9298);
xnor UO_170 (O_170,N_8333,N_8246);
or UO_171 (O_171,N_9740,N_8225);
and UO_172 (O_172,N_9393,N_8378);
xnor UO_173 (O_173,N_9796,N_9629);
and UO_174 (O_174,N_8869,N_8354);
xnor UO_175 (O_175,N_9868,N_8226);
and UO_176 (O_176,N_8235,N_8323);
nor UO_177 (O_177,N_8056,N_8551);
nand UO_178 (O_178,N_8179,N_9292);
nor UO_179 (O_179,N_9612,N_8380);
nand UO_180 (O_180,N_8277,N_8695);
xnor UO_181 (O_181,N_8680,N_8480);
nor UO_182 (O_182,N_8288,N_8015);
or UO_183 (O_183,N_8012,N_8528);
nor UO_184 (O_184,N_9506,N_9888);
and UO_185 (O_185,N_9511,N_8095);
or UO_186 (O_186,N_8970,N_8138);
nor UO_187 (O_187,N_9502,N_8662);
and UO_188 (O_188,N_8590,N_9400);
or UO_189 (O_189,N_8973,N_8600);
and UO_190 (O_190,N_9817,N_8376);
and UO_191 (O_191,N_8173,N_9728);
and UO_192 (O_192,N_8633,N_8906);
nor UO_193 (O_193,N_8115,N_9807);
or UO_194 (O_194,N_8794,N_9181);
or UO_195 (O_195,N_9085,N_9116);
xor UO_196 (O_196,N_9299,N_9572);
nand UO_197 (O_197,N_9156,N_9706);
nand UO_198 (O_198,N_8744,N_8591);
nor UO_199 (O_199,N_8239,N_9453);
nand UO_200 (O_200,N_8961,N_8715);
xnor UO_201 (O_201,N_9996,N_8908);
and UO_202 (O_202,N_9557,N_8686);
nand UO_203 (O_203,N_8793,N_8702);
nor UO_204 (O_204,N_9736,N_9877);
and UO_205 (O_205,N_8783,N_9293);
nand UO_206 (O_206,N_8923,N_8664);
nand UO_207 (O_207,N_9487,N_9336);
nand UO_208 (O_208,N_8635,N_9162);
and UO_209 (O_209,N_9026,N_9088);
or UO_210 (O_210,N_8088,N_8274);
and UO_211 (O_211,N_8910,N_9414);
nand UO_212 (O_212,N_9204,N_8598);
xor UO_213 (O_213,N_8442,N_8045);
nand UO_214 (O_214,N_9142,N_9486);
xor UO_215 (O_215,N_9070,N_8966);
and UO_216 (O_216,N_8112,N_9238);
xor UO_217 (O_217,N_8294,N_9894);
xor UO_218 (O_218,N_8994,N_9174);
or UO_219 (O_219,N_9870,N_9077);
nand UO_220 (O_220,N_9074,N_8304);
nor UO_221 (O_221,N_8537,N_9191);
nor UO_222 (O_222,N_8888,N_8098);
nand UO_223 (O_223,N_9332,N_9027);
xnor UO_224 (O_224,N_8458,N_9701);
nand UO_225 (O_225,N_8903,N_9841);
and UO_226 (O_226,N_8165,N_9780);
xnor UO_227 (O_227,N_9684,N_8546);
or UO_228 (O_228,N_9068,N_8147);
nor UO_229 (O_229,N_9660,N_8854);
xnor UO_230 (O_230,N_9049,N_8907);
nand UO_231 (O_231,N_8953,N_9122);
nand UO_232 (O_232,N_8918,N_9461);
nor UO_233 (O_233,N_8358,N_9193);
nand UO_234 (O_234,N_8522,N_8145);
nand UO_235 (O_235,N_9048,N_9801);
or UO_236 (O_236,N_8768,N_8441);
or UO_237 (O_237,N_8316,N_8494);
nand UO_238 (O_238,N_8637,N_8368);
or UO_239 (O_239,N_9126,N_9087);
and UO_240 (O_240,N_9399,N_9334);
or UO_241 (O_241,N_8474,N_8260);
and UO_242 (O_242,N_8261,N_9202);
xnor UO_243 (O_243,N_8300,N_9634);
and UO_244 (O_244,N_9419,N_9225);
or UO_245 (O_245,N_9227,N_8152);
and UO_246 (O_246,N_8892,N_9525);
nor UO_247 (O_247,N_8722,N_9131);
nor UO_248 (O_248,N_8787,N_8886);
nand UO_249 (O_249,N_8796,N_9106);
nor UO_250 (O_250,N_9960,N_9725);
and UO_251 (O_251,N_8393,N_9973);
nand UO_252 (O_252,N_9593,N_9397);
or UO_253 (O_253,N_9335,N_9383);
and UO_254 (O_254,N_8345,N_8199);
xnor UO_255 (O_255,N_9302,N_8898);
and UO_256 (O_256,N_9681,N_9250);
and UO_257 (O_257,N_8626,N_8612);
nand UO_258 (O_258,N_8799,N_8987);
and UO_259 (O_259,N_8777,N_8417);
xor UO_260 (O_260,N_8938,N_8253);
and UO_261 (O_261,N_8714,N_8915);
xnor UO_262 (O_262,N_9109,N_8232);
nor UO_263 (O_263,N_8197,N_9128);
xor UO_264 (O_264,N_9704,N_8839);
nor UO_265 (O_265,N_9321,N_8849);
nand UO_266 (O_266,N_9164,N_8486);
nand UO_267 (O_267,N_9693,N_8307);
and UO_268 (O_268,N_9741,N_9342);
or UO_269 (O_269,N_8178,N_8320);
nor UO_270 (O_270,N_9339,N_8789);
xnor UO_271 (O_271,N_9903,N_8921);
or UO_272 (O_272,N_8631,N_8509);
xnor UO_273 (O_273,N_9584,N_8371);
or UO_274 (O_274,N_8881,N_9413);
nor UO_275 (O_275,N_9360,N_8564);
xor UO_276 (O_276,N_9270,N_8064);
nor UO_277 (O_277,N_8557,N_9028);
or UO_278 (O_278,N_9901,N_9401);
nor UO_279 (O_279,N_8488,N_9792);
nand UO_280 (O_280,N_8144,N_8308);
nor UO_281 (O_281,N_8476,N_8503);
xor UO_282 (O_282,N_9508,N_8156);
nand UO_283 (O_283,N_9097,N_9569);
and UO_284 (O_284,N_8118,N_9375);
nand UO_285 (O_285,N_8983,N_8786);
and UO_286 (O_286,N_9883,N_9939);
nand UO_287 (O_287,N_9039,N_9016);
and UO_288 (O_288,N_8698,N_8003);
nand UO_289 (O_289,N_9613,N_9904);
or UO_290 (O_290,N_9782,N_8672);
nand UO_291 (O_291,N_8743,N_8643);
nand UO_292 (O_292,N_9001,N_9956);
and UO_293 (O_293,N_8815,N_9929);
nand UO_294 (O_294,N_8770,N_8357);
xor UO_295 (O_295,N_9906,N_9760);
nor UO_296 (O_296,N_9173,N_8845);
or UO_297 (O_297,N_8889,N_8599);
nand UO_298 (O_298,N_9395,N_9935);
nand UO_299 (O_299,N_9443,N_8831);
xor UO_300 (O_300,N_8762,N_8291);
and UO_301 (O_301,N_9226,N_9260);
and UO_302 (O_302,N_8822,N_9545);
xnor UO_303 (O_303,N_9566,N_9970);
nor UO_304 (O_304,N_8337,N_9426);
and UO_305 (O_305,N_8500,N_8431);
and UO_306 (O_306,N_8334,N_8971);
xnor UO_307 (O_307,N_9585,N_8864);
nor UO_308 (O_308,N_8169,N_9758);
xor UO_309 (O_309,N_8758,N_8833);
and UO_310 (O_310,N_8674,N_8682);
xor UO_311 (O_311,N_9137,N_9884);
nand UO_312 (O_312,N_9024,N_9721);
nand UO_313 (O_313,N_9898,N_9527);
nor UO_314 (O_314,N_8331,N_9697);
xnor UO_315 (O_315,N_9370,N_8049);
and UO_316 (O_316,N_8418,N_9518);
or UO_317 (O_317,N_9916,N_8692);
nand UO_318 (O_318,N_8667,N_9815);
nor UO_319 (O_319,N_8126,N_9755);
or UO_320 (O_320,N_9151,N_8078);
and UO_321 (O_321,N_8818,N_8120);
nand UO_322 (O_322,N_9534,N_9451);
and UO_323 (O_323,N_9781,N_9172);
xnor UO_324 (O_324,N_9644,N_9757);
nor UO_325 (O_325,N_8391,N_8201);
and UO_326 (O_326,N_9376,N_8438);
nand UO_327 (O_327,N_8678,N_8472);
or UO_328 (O_328,N_9115,N_9699);
xor UO_329 (O_329,N_8171,N_9959);
nand UO_330 (O_330,N_9127,N_8188);
nor UO_331 (O_331,N_9769,N_9079);
or UO_332 (O_332,N_9712,N_9882);
xor UO_333 (O_333,N_8423,N_8894);
nand UO_334 (O_334,N_9663,N_8149);
xnor UO_335 (O_335,N_8775,N_8047);
nor UO_336 (O_336,N_9344,N_8718);
and UO_337 (O_337,N_8230,N_9437);
xnor UO_338 (O_338,N_8658,N_8592);
nor UO_339 (O_339,N_9391,N_9125);
xor UO_340 (O_340,N_9905,N_8437);
or UO_341 (O_341,N_9313,N_9952);
and UO_342 (O_342,N_9950,N_9450);
or UO_343 (O_343,N_8940,N_9520);
or UO_344 (O_344,N_9045,N_8617);
xnor UO_345 (O_345,N_8946,N_9073);
nor UO_346 (O_346,N_9958,N_9096);
nor UO_347 (O_347,N_9060,N_9764);
and UO_348 (O_348,N_8607,N_9953);
nor UO_349 (O_349,N_9733,N_9517);
and UO_350 (O_350,N_9842,N_9601);
and UO_351 (O_351,N_8523,N_8455);
nor UO_352 (O_352,N_9911,N_8266);
nand UO_353 (O_353,N_8278,N_8315);
and UO_354 (O_354,N_9827,N_9718);
nor UO_355 (O_355,N_8756,N_8264);
xnor UO_356 (O_356,N_8942,N_9556);
xor UO_357 (O_357,N_9766,N_9182);
nor UO_358 (O_358,N_8616,N_9899);
or UO_359 (O_359,N_9678,N_8141);
xnor UO_360 (O_360,N_9320,N_9387);
and UO_361 (O_361,N_9679,N_9878);
and UO_362 (O_362,N_9924,N_8703);
or UO_363 (O_363,N_8553,N_8675);
xor UO_364 (O_364,N_9848,N_9530);
nor UO_365 (O_365,N_8977,N_8992);
nand UO_366 (O_366,N_9044,N_8440);
and UO_367 (O_367,N_9431,N_9154);
nand UO_368 (O_368,N_9765,N_9977);
nand UO_369 (O_369,N_9537,N_9738);
or UO_370 (O_370,N_8065,N_8844);
nand UO_371 (O_371,N_9094,N_8639);
nand UO_372 (O_372,N_8810,N_9080);
nand UO_373 (O_373,N_9117,N_9671);
or UO_374 (O_374,N_9816,N_9307);
nor UO_375 (O_375,N_9988,N_8897);
nand UO_376 (O_376,N_8584,N_9843);
xnor UO_377 (O_377,N_8835,N_9124);
nand UO_378 (O_378,N_8314,N_9337);
nor UO_379 (O_379,N_8091,N_8769);
nor UO_380 (O_380,N_8449,N_8168);
nor UO_381 (O_381,N_8207,N_8990);
nor UO_382 (O_382,N_9177,N_9768);
nor UO_383 (O_383,N_9312,N_9480);
nor UO_384 (O_384,N_8511,N_9002);
nand UO_385 (O_385,N_8878,N_8401);
nor UO_386 (O_386,N_9194,N_9944);
nor UO_387 (O_387,N_9567,N_8432);
nand UO_388 (O_388,N_8305,N_8559);
or UO_389 (O_389,N_8569,N_9824);
nand UO_390 (O_390,N_9314,N_8862);
nor UO_391 (O_391,N_8857,N_9794);
nor UO_392 (O_392,N_8255,N_8552);
nand UO_393 (O_393,N_8279,N_8075);
nor UO_394 (O_394,N_8957,N_8991);
nand UO_395 (O_395,N_8211,N_8224);
and UO_396 (O_396,N_8934,N_9140);
or UO_397 (O_397,N_8166,N_9821);
nand UO_398 (O_398,N_9482,N_9329);
or UO_399 (O_399,N_9136,N_9427);
or UO_400 (O_400,N_8801,N_9799);
nand UO_401 (O_401,N_9887,N_8052);
xnor UO_402 (O_402,N_8067,N_9987);
xor UO_403 (O_403,N_9927,N_9576);
or UO_404 (O_404,N_9641,N_8446);
or UO_405 (O_405,N_9602,N_9111);
xor UO_406 (O_406,N_9264,N_9121);
nor UO_407 (O_407,N_8689,N_9300);
or UO_408 (O_408,N_8629,N_8459);
xnor UO_409 (O_409,N_9611,N_9331);
nand UO_410 (O_410,N_8451,N_9896);
nand UO_411 (O_411,N_9811,N_9778);
nand UO_412 (O_412,N_9015,N_9492);
or UO_413 (O_413,N_8883,N_9281);
nand UO_414 (O_414,N_8164,N_8792);
nand UO_415 (O_415,N_9713,N_8292);
and UO_416 (O_416,N_9717,N_9361);
nand UO_417 (O_417,N_9295,N_9197);
nor UO_418 (O_418,N_8676,N_8286);
nor UO_419 (O_419,N_9991,N_8984);
and UO_420 (O_420,N_8251,N_8836);
and UO_421 (O_421,N_9237,N_8250);
nand UO_422 (O_422,N_8238,N_9596);
nor UO_423 (O_423,N_9965,N_9428);
nor UO_424 (O_424,N_9565,N_9720);
xor UO_425 (O_425,N_8119,N_8924);
xor UO_426 (O_426,N_9621,N_9885);
and UO_427 (O_427,N_9253,N_9219);
xor UO_428 (O_428,N_8510,N_8330);
xnor UO_429 (O_429,N_9043,N_9269);
nand UO_430 (O_430,N_8403,N_9873);
nand UO_431 (O_431,N_9368,N_8838);
or UO_432 (O_432,N_8507,N_8059);
xor UO_433 (O_433,N_9266,N_8070);
xnor UO_434 (O_434,N_8384,N_9051);
and UO_435 (O_435,N_9470,N_9442);
xnor UO_436 (O_436,N_8086,N_9362);
xnor UO_437 (O_437,N_8021,N_9377);
nor UO_438 (O_438,N_8624,N_8753);
xor UO_439 (O_439,N_9203,N_9756);
nor UO_440 (O_440,N_8604,N_9834);
nor UO_441 (O_441,N_9095,N_9806);
or UO_442 (O_442,N_9021,N_9071);
xnor UO_443 (O_443,N_9966,N_8099);
xor UO_444 (O_444,N_9086,N_8968);
or UO_445 (O_445,N_8730,N_8725);
nand UO_446 (O_446,N_8949,N_8567);
and UO_447 (O_447,N_8814,N_9289);
or UO_448 (O_448,N_9890,N_9919);
nor UO_449 (O_449,N_9190,N_9448);
and UO_450 (O_450,N_9822,N_8107);
nand UO_451 (O_451,N_9550,N_8276);
xnor UO_452 (O_452,N_9409,N_8428);
and UO_453 (O_453,N_9388,N_8066);
and UO_454 (O_454,N_8491,N_8773);
xor UO_455 (O_455,N_8074,N_8955);
nor UO_456 (O_456,N_8038,N_9734);
or UO_457 (O_457,N_9891,N_8943);
nand UO_458 (O_458,N_8673,N_8213);
and UO_459 (O_459,N_8361,N_9774);
and UO_460 (O_460,N_9505,N_9228);
and UO_461 (O_461,N_9654,N_9220);
nand UO_462 (O_462,N_9102,N_9809);
nor UO_463 (O_463,N_9637,N_8130);
nor UO_464 (O_464,N_9476,N_9836);
nand UO_465 (O_465,N_9438,N_9784);
and UO_466 (O_466,N_9030,N_9864);
nor UO_467 (O_467,N_8129,N_9510);
or UO_468 (O_468,N_9747,N_8561);
and UO_469 (O_469,N_9493,N_8104);
xnor UO_470 (O_470,N_8939,N_9819);
or UO_471 (O_471,N_9997,N_9011);
and UO_472 (O_472,N_8041,N_9600);
xor UO_473 (O_473,N_9152,N_8402);
xnor UO_474 (O_474,N_8520,N_8338);
nand UO_475 (O_475,N_8817,N_8999);
xor UO_476 (O_476,N_9159,N_9521);
nor UO_477 (O_477,N_9255,N_9618);
and UO_478 (O_478,N_9773,N_9785);
or UO_479 (O_479,N_8663,N_8317);
nor UO_480 (O_480,N_8044,N_9932);
xnor UO_481 (O_481,N_8754,N_9879);
xnor UO_482 (O_482,N_8874,N_8985);
nand UO_483 (O_483,N_8336,N_9195);
xor UO_484 (O_484,N_9789,N_9969);
and UO_485 (O_485,N_8069,N_8463);
and UO_486 (O_486,N_9326,N_9201);
xor UO_487 (O_487,N_9542,N_8707);
nand UO_488 (O_488,N_9103,N_9038);
or UO_489 (O_489,N_8425,N_8548);
xor UO_490 (O_490,N_8603,N_8788);
or UO_491 (O_491,N_8057,N_8081);
nand UO_492 (O_492,N_9404,N_8234);
and UO_493 (O_493,N_9571,N_8259);
and UO_494 (O_494,N_8200,N_9786);
nand UO_495 (O_495,N_9509,N_9865);
or UO_496 (O_496,N_9316,N_8103);
and UO_497 (O_497,N_8035,N_9688);
and UO_498 (O_498,N_8398,N_9649);
nor UO_499 (O_499,N_9677,N_9069);
xnor UO_500 (O_500,N_8293,N_9910);
and UO_501 (O_501,N_8896,N_8566);
and UO_502 (O_502,N_8034,N_8063);
or UO_503 (O_503,N_8723,N_8875);
or UO_504 (O_504,N_8805,N_8386);
nand UO_505 (O_505,N_9359,N_9222);
or UO_506 (O_506,N_8273,N_9683);
xnor UO_507 (O_507,N_9241,N_9856);
nor UO_508 (O_508,N_9529,N_8790);
nor UO_509 (O_509,N_9296,N_8478);
and UO_510 (O_510,N_8711,N_8290);
xnor UO_511 (O_511,N_8610,N_8641);
xnor UO_512 (O_512,N_9630,N_8905);
nor UO_513 (O_513,N_8209,N_9052);
nor UO_514 (O_514,N_9946,N_9452);
or UO_515 (O_515,N_9742,N_9860);
or UO_516 (O_516,N_8448,N_9358);
nand UO_517 (O_517,N_9866,N_9653);
nand UO_518 (O_518,N_8978,N_8421);
and UO_519 (O_519,N_8319,N_9171);
xor UO_520 (O_520,N_9746,N_9770);
nor UO_521 (O_521,N_8697,N_8912);
nor UO_522 (O_522,N_8579,N_9790);
nor UO_523 (O_523,N_8019,N_8415);
xnor UO_524 (O_524,N_9833,N_9207);
nand UO_525 (O_525,N_8283,N_9995);
nand UO_526 (O_526,N_8998,N_9234);
nand UO_527 (O_527,N_9105,N_8694);
and UO_528 (O_528,N_8037,N_9350);
nor UO_529 (O_529,N_9783,N_8652);
nand UO_530 (O_530,N_8656,N_9372);
and UO_531 (O_531,N_8263,N_9196);
nor UO_532 (O_532,N_8379,N_8859);
and UO_533 (O_533,N_9212,N_8976);
and UO_534 (O_534,N_8529,N_9454);
or UO_535 (O_535,N_8240,N_9113);
xor UO_536 (O_536,N_9658,N_8089);
nor UO_537 (O_537,N_8177,N_8270);
xnor UO_538 (O_538,N_9349,N_8508);
xnor UO_539 (O_539,N_8550,N_8414);
xnor UO_540 (O_540,N_9129,N_8563);
nor UO_541 (O_541,N_8980,N_8496);
or UO_542 (O_542,N_8654,N_9430);
nand UO_543 (O_543,N_9826,N_8865);
nor UO_544 (O_544,N_9918,N_9138);
or UO_545 (O_545,N_9583,N_9389);
xor UO_546 (O_546,N_9353,N_9366);
nor UO_547 (O_547,N_8359,N_9468);
or UO_548 (O_548,N_8310,N_8007);
nor UO_549 (O_549,N_9575,N_8816);
xor UO_550 (O_550,N_9141,N_9662);
and UO_551 (O_551,N_8696,N_8413);
or UO_552 (O_552,N_8952,N_9648);
or UO_553 (O_553,N_9917,N_9055);
xnor UO_554 (O_554,N_8900,N_8175);
nand UO_555 (O_555,N_9133,N_9590);
nor UO_556 (O_556,N_8576,N_8804);
nor UO_557 (O_557,N_8516,N_8495);
nor UO_558 (O_558,N_9692,N_8807);
and UO_559 (O_559,N_8911,N_9345);
nor UO_560 (O_560,N_8490,N_9652);
and UO_561 (O_561,N_9354,N_8681);
xnor UO_562 (O_562,N_9076,N_9265);
nand UO_563 (O_563,N_8185,N_9775);
nand UO_564 (O_564,N_9751,N_9962);
nand UO_565 (O_565,N_9233,N_8893);
nor UO_566 (O_566,N_9582,N_8830);
nor UO_567 (O_567,N_9333,N_9863);
or UO_568 (O_568,N_9304,N_9107);
nor UO_569 (O_569,N_9185,N_8114);
nand UO_570 (O_570,N_9748,N_8846);
and UO_571 (O_571,N_9659,N_9867);
xnor UO_572 (O_572,N_8342,N_8568);
nor UO_573 (O_573,N_9519,N_9004);
nor UO_574 (O_574,N_8080,N_8369);
xor UO_575 (O_575,N_9290,N_9937);
or UO_576 (O_576,N_8870,N_8502);
nor UO_577 (O_577,N_9457,N_9522);
xor UO_578 (O_578,N_8589,N_8947);
or UO_579 (O_579,N_8471,N_9441);
nand UO_580 (O_580,N_9369,N_9032);
or UO_581 (O_581,N_8097,N_8427);
or UO_582 (O_582,N_8524,N_9280);
nand UO_583 (O_583,N_8571,N_8203);
nand UO_584 (O_584,N_9167,N_8671);
and UO_585 (O_585,N_8975,N_8027);
nand UO_586 (O_586,N_8751,N_9554);
or UO_587 (O_587,N_8887,N_9968);
nor UO_588 (O_588,N_9854,N_8085);
or UO_589 (O_589,N_8487,N_8623);
nor UO_590 (O_590,N_9948,N_9020);
nand UO_591 (O_591,N_8647,N_8541);
nor UO_592 (O_592,N_8473,N_9199);
nand UO_593 (O_593,N_9907,N_9808);
or UO_594 (O_594,N_9439,N_9687);
and UO_595 (O_595,N_9484,N_8462);
nand UO_596 (O_596,N_8127,N_8752);
and UO_597 (O_597,N_8229,N_9447);
nand UO_598 (O_598,N_8780,N_8190);
xor UO_599 (O_599,N_9496,N_8759);
xor UO_600 (O_600,N_8737,N_8134);
and UO_601 (O_601,N_8392,N_9563);
nand UO_602 (O_602,N_9592,N_8925);
or UO_603 (O_603,N_9558,N_8745);
nand UO_604 (O_604,N_9327,N_8964);
xor UO_605 (O_605,N_8741,N_8582);
or UO_606 (O_606,N_9408,N_9690);
nand UO_607 (O_607,N_9814,N_9716);
or UO_608 (O_608,N_8735,N_9235);
nand UO_609 (O_609,N_9034,N_9570);
and UO_610 (O_610,N_9695,N_9465);
or UO_611 (O_611,N_9417,N_8210);
or UO_612 (O_612,N_8465,N_9514);
nand UO_613 (O_613,N_8969,N_9893);
and UO_614 (O_614,N_9622,N_8183);
xor UO_615 (O_615,N_8020,N_9285);
or UO_616 (O_616,N_9239,N_8746);
nand UO_617 (O_617,N_8712,N_9633);
and UO_618 (O_618,N_9972,N_9249);
or UO_619 (O_619,N_8766,N_8340);
or UO_620 (O_620,N_8090,N_9364);
nor UO_621 (O_621,N_9975,N_9211);
xnor UO_622 (O_622,N_8902,N_9536);
or UO_623 (O_623,N_9892,N_9423);
xor UO_624 (O_624,N_8374,N_8030);
nand UO_625 (O_625,N_9035,N_9217);
and UO_626 (O_626,N_8872,N_9925);
nor UO_627 (O_627,N_8684,N_8806);
or UO_628 (O_628,N_9135,N_8457);
or UO_629 (O_629,N_9847,N_8332);
nand UO_630 (O_630,N_8691,N_8562);
and UO_631 (O_631,N_8954,N_8042);
nor UO_632 (O_632,N_9920,N_8824);
xnor UO_633 (O_633,N_8287,N_9729);
and UO_634 (O_634,N_8764,N_9338);
nand UO_635 (O_635,N_8245,N_8765);
and UO_636 (O_636,N_9947,N_9540);
xor UO_637 (O_637,N_9477,N_8111);
and UO_638 (O_638,N_8534,N_9727);
and UO_639 (O_639,N_9005,N_8951);
nor UO_640 (O_640,N_9722,N_8484);
or UO_641 (O_641,N_8366,N_8172);
or UO_642 (O_642,N_9564,N_8880);
nand UO_643 (O_643,N_8936,N_9754);
nor UO_644 (O_644,N_8959,N_8929);
nand UO_645 (O_645,N_8842,N_8913);
or UO_646 (O_646,N_9046,N_9017);
and UO_647 (O_647,N_8648,N_8101);
or UO_648 (O_648,N_9236,N_8556);
xor UO_649 (O_649,N_9745,N_8885);
nand UO_650 (O_650,N_9084,N_9606);
nor UO_651 (O_651,N_8530,N_9675);
or UO_652 (O_652,N_9278,N_8284);
and UO_653 (O_653,N_8646,N_8543);
nor UO_654 (O_654,N_8096,N_9964);
xnor UO_655 (O_655,N_8105,N_9411);
nand UO_656 (O_656,N_8174,N_9184);
or UO_657 (O_657,N_8965,N_8729);
and UO_658 (O_658,N_9646,N_8475);
or UO_659 (O_659,N_9691,N_8388);
or UO_660 (O_660,N_9625,N_9732);
nand UO_661 (O_661,N_8351,N_9589);
xnor UO_662 (O_662,N_8521,N_9526);
nor UO_663 (O_663,N_8884,N_8325);
nor UO_664 (O_664,N_9912,N_9580);
nand UO_665 (O_665,N_8219,N_8008);
and UO_666 (O_666,N_8688,N_9763);
nand UO_667 (O_667,N_8483,N_8154);
and UO_668 (O_668,N_9262,N_8489);
xor UO_669 (O_669,N_9846,N_9218);
nor UO_670 (O_670,N_8931,N_9610);
xor UO_671 (O_671,N_9037,N_9146);
xor UO_672 (O_672,N_9371,N_8661);
nor UO_673 (O_673,N_8795,N_9881);
nor UO_674 (O_674,N_9945,N_9696);
nand UO_675 (O_675,N_9104,N_8464);
and UO_676 (O_676,N_9813,N_9041);
xor UO_677 (O_677,N_8079,N_8798);
xnor UO_678 (O_678,N_8311,N_8679);
and UO_679 (O_679,N_9147,N_9274);
and UO_680 (O_680,N_9724,N_9636);
nand UO_681 (O_681,N_9271,N_8153);
xor UO_682 (O_682,N_8372,N_8587);
nor UO_683 (O_683,N_8375,N_9664);
or UO_684 (O_684,N_9872,N_8412);
xor UO_685 (O_685,N_8956,N_9405);
xnor UO_686 (O_686,N_9343,N_8328);
and UO_687 (O_687,N_8227,N_9018);
or UO_688 (O_688,N_9850,N_9179);
nor UO_689 (O_689,N_8109,N_8485);
nor UO_690 (O_690,N_9639,N_8092);
nor UO_691 (O_691,N_8385,N_9445);
or UO_692 (O_692,N_9776,N_8498);
and UO_693 (O_693,N_8659,N_8186);
xnor UO_694 (O_694,N_9676,N_9275);
and UO_695 (O_695,N_8608,N_8644);
nand UO_696 (O_696,N_9642,N_9750);
and UO_697 (O_697,N_9761,N_9980);
or UO_698 (O_698,N_8602,N_8271);
or UO_699 (O_699,N_9954,N_8660);
and UO_700 (O_700,N_9489,N_8055);
and UO_701 (O_701,N_8396,N_8170);
or UO_702 (O_702,N_8532,N_9539);
and UO_703 (O_703,N_9093,N_8733);
or UO_704 (O_704,N_8493,N_9993);
nor UO_705 (O_705,N_9698,N_9112);
and UO_706 (O_706,N_8355,N_9148);
xnor UO_707 (O_707,N_9829,N_9994);
xor UO_708 (O_708,N_8269,N_8687);
and UO_709 (O_709,N_9082,N_8583);
and UO_710 (O_710,N_8005,N_8191);
nand UO_711 (O_711,N_9464,N_9287);
or UO_712 (O_712,N_8017,N_9012);
nor UO_713 (O_713,N_8871,N_8363);
or UO_714 (O_714,N_8618,N_8916);
or UO_715 (O_715,N_8843,N_9976);
xnor UO_716 (O_716,N_9543,N_9499);
and UO_717 (O_717,N_8272,N_9187);
or UO_718 (O_718,N_8029,N_9340);
xor UO_719 (O_719,N_8812,N_9029);
or UO_720 (O_720,N_9626,N_8347);
and UO_721 (O_721,N_9101,N_8143);
xnor UO_722 (O_722,N_9198,N_9189);
and UO_723 (O_723,N_8024,N_9007);
nand UO_724 (O_724,N_9672,N_8280);
xor UO_725 (O_725,N_9915,N_8499);
nand UO_726 (O_726,N_9063,N_8879);
xor UO_727 (O_727,N_8439,N_8322);
or UO_728 (O_728,N_9478,N_8601);
or UO_729 (O_729,N_8150,N_9538);
xnor UO_730 (O_730,N_9297,N_9880);
nand UO_731 (O_731,N_9474,N_8452);
or UO_732 (O_732,N_8382,N_8453);
nand UO_733 (O_733,N_9715,N_8365);
and UO_734 (O_734,N_9139,N_9014);
nor UO_735 (O_735,N_9245,N_9481);
and UO_736 (O_736,N_8479,N_9500);
and UO_737 (O_737,N_8128,N_9805);
xor UO_738 (O_738,N_8082,N_9791);
nand UO_739 (O_739,N_9276,N_8774);
and UO_740 (O_740,N_8298,N_9261);
or UO_741 (O_741,N_9710,N_9433);
nor UO_742 (O_742,N_9483,N_9694);
xnor UO_743 (O_743,N_9674,N_8651);
nand UO_744 (O_744,N_8445,N_8851);
nand UO_745 (O_745,N_8084,N_8327);
nor UO_746 (O_746,N_8004,N_9588);
or UO_747 (O_747,N_8220,N_9771);
and UO_748 (O_748,N_9574,N_9812);
xor UO_749 (O_749,N_8781,N_9040);
xor UO_750 (O_750,N_8716,N_9380);
or UO_751 (O_751,N_9066,N_8785);
nand UO_752 (O_752,N_8593,N_8979);
nand UO_753 (O_753,N_8709,N_9403);
xnor UO_754 (O_754,N_9057,N_8221);
and UO_755 (O_755,N_9168,N_8206);
nor UO_756 (O_756,N_8467,N_8125);
and UO_757 (O_757,N_8549,N_9379);
nor UO_758 (O_758,N_8352,N_9166);
nor UO_759 (O_759,N_9726,N_8642);
or UO_760 (O_760,N_9382,N_9186);
and UO_761 (O_761,N_9800,N_8058);
nor UO_762 (O_762,N_8410,N_9876);
nor UO_763 (O_763,N_9488,N_9123);
nor UO_764 (O_764,N_9983,N_9455);
and UO_765 (O_765,N_8329,N_9665);
xnor UO_766 (O_766,N_8861,N_8009);
or UO_767 (O_767,N_8036,N_9616);
and UO_768 (O_768,N_9926,N_9114);
nand UO_769 (O_769,N_8062,N_8377);
nor UO_770 (O_770,N_8383,N_8158);
nand UO_771 (O_771,N_9176,N_8895);
xor UO_772 (O_772,N_9941,N_9119);
nor UO_773 (O_773,N_8570,N_8727);
or UO_774 (O_774,N_8819,N_8609);
or UO_775 (O_775,N_8113,N_8405);
and UO_776 (O_776,N_9373,N_8625);
and UO_777 (O_777,N_9351,N_9951);
xnor UO_778 (O_778,N_9444,N_9928);
nor UO_779 (O_779,N_8748,N_8666);
nand UO_780 (O_780,N_8436,N_8993);
and UO_781 (O_781,N_8525,N_8422);
nand UO_782 (O_782,N_9656,N_8778);
and UO_783 (O_783,N_9820,N_8636);
and UO_784 (O_784,N_8734,N_8670);
nor UO_785 (O_785,N_9861,N_9940);
and UO_786 (O_786,N_8944,N_8739);
xor UO_787 (O_787,N_8834,N_8640);
nand UO_788 (O_788,N_8772,N_9059);
and UO_789 (O_789,N_8634,N_8578);
and UO_790 (O_790,N_9802,N_8231);
nor UO_791 (O_791,N_8755,N_8108);
nand UO_792 (O_792,N_8747,N_8565);
nand UO_793 (O_793,N_8151,N_9767);
nand UO_794 (O_794,N_8989,N_8767);
nor UO_795 (O_795,N_9913,N_9668);
xnor UO_796 (O_796,N_9169,N_8087);
nand UO_797 (O_797,N_9669,N_8742);
and UO_798 (O_798,N_9923,N_9551);
nor UO_799 (O_799,N_9495,N_9418);
and UO_800 (O_800,N_9604,N_9308);
xnor UO_801 (O_801,N_9003,N_9291);
xnor UO_802 (O_802,N_8558,N_8710);
and UO_803 (O_803,N_9061,N_9022);
nand UO_804 (O_804,N_9042,N_8481);
nor UO_805 (O_805,N_9573,N_9288);
nand UO_806 (O_806,N_8685,N_8054);
or UO_807 (O_807,N_8505,N_8821);
nand UO_808 (O_808,N_9341,N_9900);
xnor UO_809 (O_809,N_8665,N_9145);
xnor UO_810 (O_810,N_9686,N_8784);
xor UO_811 (O_811,N_8581,N_8782);
and UO_812 (O_812,N_8704,N_9595);
nor UO_813 (O_813,N_9714,N_8699);
and UO_814 (O_814,N_9730,N_8873);
or UO_815 (O_815,N_8853,N_9549);
xnor UO_816 (O_816,N_8243,N_9934);
or UO_817 (O_817,N_9875,N_9279);
or UO_818 (O_818,N_9985,N_8196);
or UO_819 (O_819,N_8148,N_9374);
xor UO_820 (O_820,N_8606,N_8370);
xnor UO_821 (O_821,N_9619,N_9739);
and UO_822 (O_822,N_9175,N_8053);
nand UO_823 (O_823,N_9150,N_9303);
or UO_824 (O_824,N_8321,N_8281);
xnor UO_825 (O_825,N_8580,N_8349);
nor UO_826 (O_826,N_9719,N_8116);
xor UO_827 (O_827,N_9412,N_9516);
xnor UO_828 (O_828,N_8025,N_8933);
xor UO_829 (O_829,N_8960,N_8344);
xor UO_830 (O_830,N_8214,N_8837);
nor UO_831 (O_831,N_8202,N_8060);
nand UO_832 (O_832,N_8435,N_8588);
or UO_833 (O_833,N_8167,N_9273);
or UO_834 (O_834,N_9462,N_9979);
xnor UO_835 (O_835,N_9931,N_8619);
nor UO_836 (O_836,N_8544,N_8121);
nor UO_837 (O_837,N_8456,N_9348);
and UO_838 (O_838,N_9963,N_8389);
nor UO_839 (O_839,N_9703,N_9356);
and UO_840 (O_840,N_9050,N_8497);
nor UO_841 (O_841,N_8866,N_9957);
nand UO_842 (O_842,N_9643,N_8890);
xor UO_843 (O_843,N_9054,N_9209);
nor UO_844 (O_844,N_8904,N_8237);
nand UO_845 (O_845,N_8033,N_9205);
and UO_846 (O_846,N_8628,N_9317);
xnor UO_847 (O_847,N_9072,N_8249);
and UO_848 (O_848,N_9306,N_9591);
and UO_849 (O_849,N_8395,N_8106);
and UO_850 (O_850,N_8776,N_8575);
and UO_851 (O_851,N_9352,N_8708);
and UO_852 (O_852,N_8356,N_9180);
nand UO_853 (O_853,N_9594,N_8076);
nand UO_854 (O_854,N_8256,N_9788);
or UO_855 (O_855,N_9429,N_9689);
xnor UO_856 (O_856,N_9825,N_9210);
or UO_857 (O_857,N_9828,N_9062);
nand UO_858 (O_858,N_8192,N_9243);
xor UO_859 (O_859,N_8050,N_9859);
xnor UO_860 (O_860,N_8406,N_8482);
and UO_861 (O_861,N_9223,N_8974);
and UO_862 (O_862,N_9385,N_8967);
or UO_863 (O_863,N_9446,N_8997);
or UO_864 (O_864,N_8713,N_8301);
and UO_865 (O_865,N_8468,N_9586);
xnor UO_866 (O_866,N_8848,N_9793);
nand UO_867 (O_867,N_9889,N_9624);
and UO_868 (O_868,N_9561,N_8408);
and UO_869 (O_869,N_9100,N_8420);
xnor UO_870 (O_870,N_8855,N_8504);
nand UO_871 (O_871,N_8791,N_9936);
or UO_872 (O_872,N_8852,N_9425);
and UO_873 (O_873,N_9294,N_8254);
or UO_874 (O_874,N_8001,N_8124);
or UO_875 (O_875,N_8257,N_8645);
nand UO_876 (O_876,N_8813,N_8011);
nand UO_877 (O_877,N_8424,N_8763);
nor UO_878 (O_878,N_8962,N_9256);
xor UO_879 (O_879,N_8416,N_8000);
or UO_880 (O_880,N_8981,N_8928);
nand UO_881 (O_881,N_9560,N_9504);
nand UO_882 (O_882,N_8963,N_8447);
and UO_883 (O_883,N_8407,N_8215);
xnor UO_884 (O_884,N_8517,N_9599);
and UO_885 (O_885,N_9628,N_8155);
nor UO_886 (O_886,N_9324,N_9258);
nor UO_887 (O_887,N_9459,N_8536);
nor UO_888 (O_888,N_8343,N_9839);
and UO_889 (O_889,N_8948,N_8720);
xor UO_890 (O_890,N_8841,N_8469);
and UO_891 (O_891,N_8161,N_8868);
nor UO_892 (O_892,N_8638,N_8218);
nor UO_893 (O_893,N_8726,N_8717);
nand UO_894 (O_894,N_8518,N_9578);
xor UO_895 (O_895,N_9435,N_9064);
or UO_896 (O_896,N_9242,N_9160);
nand UO_897 (O_897,N_9818,N_8668);
or UO_898 (O_898,N_8364,N_9310);
nand UO_899 (O_899,N_9248,N_9251);
nor UO_900 (O_900,N_8187,N_8252);
or UO_901 (O_901,N_9381,N_8527);
nand UO_902 (O_902,N_8803,N_9472);
nand UO_903 (O_903,N_9089,N_9555);
nor UO_904 (O_904,N_9118,N_9267);
xor UO_905 (O_905,N_8223,N_9849);
or UO_906 (O_906,N_8433,N_8100);
nand UO_907 (O_907,N_8430,N_8061);
nand UO_908 (O_908,N_9553,N_9989);
xnor UO_909 (O_909,N_9938,N_9075);
or UO_910 (O_910,N_9787,N_8353);
nor UO_911 (O_911,N_8296,N_8515);
and UO_912 (O_912,N_8160,N_8596);
nand UO_913 (O_913,N_9008,N_9467);
or UO_914 (O_914,N_9753,N_9603);
nor UO_915 (O_915,N_8909,N_8208);
nor UO_916 (O_916,N_8863,N_9215);
or UO_917 (O_917,N_9244,N_9535);
and UO_918 (O_918,N_8426,N_9562);
or UO_919 (O_919,N_8265,N_8133);
nand UO_920 (O_920,N_9598,N_9647);
nor UO_921 (O_921,N_9263,N_8411);
xnor UO_922 (O_922,N_8800,N_9047);
or UO_923 (O_923,N_9845,N_9325);
nor UO_924 (O_924,N_9282,N_8649);
and UO_925 (O_925,N_9056,N_9837);
or UO_926 (O_926,N_8926,N_9025);
and UO_927 (O_927,N_9378,N_9161);
or UO_928 (O_928,N_8657,N_9921);
nor UO_929 (O_929,N_8683,N_9685);
or UO_930 (O_930,N_9844,N_9597);
nand UO_931 (O_931,N_9155,N_9206);
or UO_932 (O_932,N_8950,N_8982);
nor UO_933 (O_933,N_8470,N_8995);
or UO_934 (O_934,N_9568,N_8901);
and UO_935 (O_935,N_8077,N_8914);
and UO_936 (O_936,N_8434,N_8693);
xor UO_937 (O_937,N_8123,N_9548);
or UO_938 (O_938,N_8466,N_8899);
xnor UO_939 (O_939,N_8289,N_9749);
nand UO_940 (O_940,N_9853,N_8131);
and UO_941 (O_941,N_9224,N_9650);
or UO_942 (O_942,N_8554,N_9986);
xor UO_943 (O_943,N_9617,N_8040);
and UO_944 (O_944,N_8572,N_8749);
nor UO_945 (O_945,N_9998,N_9544);
or UO_946 (O_946,N_9322,N_8248);
and UO_947 (O_947,N_8719,N_8297);
nand UO_948 (O_948,N_8309,N_8655);
xnor UO_949 (O_949,N_9473,N_8771);
nand UO_950 (O_950,N_8233,N_9707);
nor UO_951 (O_951,N_9830,N_9908);
nor UO_952 (O_952,N_9777,N_9033);
xor UO_953 (O_953,N_9840,N_9384);
or UO_954 (O_954,N_9319,N_9143);
nand UO_955 (O_955,N_9609,N_8262);
and UO_956 (O_956,N_8102,N_9670);
or UO_957 (O_957,N_9396,N_8958);
nor UO_958 (O_958,N_9851,N_8212);
nor UO_959 (O_959,N_8595,N_8010);
nor UO_960 (O_960,N_8802,N_8677);
nand UO_961 (O_961,N_9581,N_8335);
nor UO_962 (O_962,N_9460,N_8731);
and UO_963 (O_963,N_9587,N_9623);
nand UO_964 (O_964,N_8443,N_9301);
nor UO_965 (O_965,N_8222,N_8258);
or UO_966 (O_966,N_9386,N_8574);
nand UO_967 (O_967,N_8627,N_8820);
and UO_968 (O_968,N_9208,N_8738);
and UO_969 (O_969,N_8701,N_8945);
and UO_970 (O_970,N_8039,N_8313);
or UO_971 (O_971,N_8922,N_9955);
and UO_972 (O_972,N_8779,N_9895);
or UO_973 (O_973,N_9967,N_9577);
nand UO_974 (O_974,N_9857,N_9232);
nand UO_975 (O_975,N_8555,N_9183);
and UO_976 (O_976,N_9981,N_9200);
nand UO_977 (O_977,N_8339,N_9192);
and UO_978 (O_978,N_9092,N_8404);
xnor UO_979 (O_979,N_8613,N_8492);
and UO_980 (O_980,N_8526,N_9252);
or UO_981 (O_981,N_8137,N_9855);
nor UO_982 (O_982,N_8632,N_9858);
or UO_983 (O_983,N_9523,N_9700);
or UO_984 (O_984,N_8615,N_8545);
nand UO_985 (O_985,N_9463,N_9286);
xnor UO_986 (O_986,N_8538,N_9743);
nand UO_987 (O_987,N_9667,N_9838);
and UO_988 (O_988,N_8180,N_8823);
nor UO_989 (O_989,N_9759,N_9134);
and UO_990 (O_990,N_9466,N_8348);
and UO_991 (O_991,N_8093,N_8740);
nor UO_992 (O_992,N_9490,N_9132);
nand UO_993 (O_993,N_8176,N_8867);
nand UO_994 (O_994,N_8397,N_8362);
nand UO_995 (O_995,N_9737,N_8182);
nor UO_996 (O_996,N_8808,N_9978);
nor UO_997 (O_997,N_9708,N_9680);
and UO_998 (O_998,N_9494,N_8184);
nand UO_999 (O_999,N_9657,N_9392);
and UO_1000 (O_1000,N_9151,N_9860);
or UO_1001 (O_1001,N_9774,N_9814);
nor UO_1002 (O_1002,N_8035,N_8974);
xnor UO_1003 (O_1003,N_8441,N_9753);
and UO_1004 (O_1004,N_9469,N_9518);
nand UO_1005 (O_1005,N_8994,N_8904);
xnor UO_1006 (O_1006,N_9691,N_8680);
nor UO_1007 (O_1007,N_8855,N_8010);
nand UO_1008 (O_1008,N_8542,N_9672);
nor UO_1009 (O_1009,N_8729,N_9798);
and UO_1010 (O_1010,N_9549,N_8172);
and UO_1011 (O_1011,N_8667,N_8719);
and UO_1012 (O_1012,N_9258,N_8134);
and UO_1013 (O_1013,N_9976,N_9948);
xor UO_1014 (O_1014,N_8070,N_9187);
or UO_1015 (O_1015,N_9320,N_8228);
nand UO_1016 (O_1016,N_9301,N_8775);
nor UO_1017 (O_1017,N_9328,N_8079);
nand UO_1018 (O_1018,N_8378,N_8897);
nor UO_1019 (O_1019,N_8950,N_9593);
or UO_1020 (O_1020,N_9632,N_8102);
nor UO_1021 (O_1021,N_8339,N_9368);
and UO_1022 (O_1022,N_9342,N_9156);
nor UO_1023 (O_1023,N_8864,N_8932);
and UO_1024 (O_1024,N_8305,N_9628);
nor UO_1025 (O_1025,N_9896,N_9198);
nor UO_1026 (O_1026,N_9443,N_9406);
nand UO_1027 (O_1027,N_8889,N_9166);
nand UO_1028 (O_1028,N_8451,N_9716);
nand UO_1029 (O_1029,N_9210,N_8468);
xnor UO_1030 (O_1030,N_8543,N_8156);
nor UO_1031 (O_1031,N_8344,N_9227);
xnor UO_1032 (O_1032,N_8708,N_9763);
nand UO_1033 (O_1033,N_8960,N_8296);
xor UO_1034 (O_1034,N_8502,N_8885);
nor UO_1035 (O_1035,N_8364,N_9840);
nor UO_1036 (O_1036,N_9542,N_8131);
nand UO_1037 (O_1037,N_8223,N_8145);
or UO_1038 (O_1038,N_9463,N_9106);
nor UO_1039 (O_1039,N_9063,N_9192);
xnor UO_1040 (O_1040,N_9389,N_9160);
and UO_1041 (O_1041,N_8589,N_8960);
and UO_1042 (O_1042,N_8566,N_8154);
and UO_1043 (O_1043,N_9606,N_9970);
nor UO_1044 (O_1044,N_9089,N_8179);
or UO_1045 (O_1045,N_9398,N_9996);
xnor UO_1046 (O_1046,N_9227,N_8326);
and UO_1047 (O_1047,N_9640,N_8650);
nor UO_1048 (O_1048,N_9587,N_9554);
nor UO_1049 (O_1049,N_8875,N_9218);
or UO_1050 (O_1050,N_9548,N_9371);
nor UO_1051 (O_1051,N_8461,N_8416);
and UO_1052 (O_1052,N_8470,N_8277);
or UO_1053 (O_1053,N_8090,N_9184);
and UO_1054 (O_1054,N_8011,N_9739);
or UO_1055 (O_1055,N_9722,N_8216);
nand UO_1056 (O_1056,N_8896,N_9751);
or UO_1057 (O_1057,N_9590,N_9621);
xnor UO_1058 (O_1058,N_8824,N_9390);
nand UO_1059 (O_1059,N_9513,N_8867);
nand UO_1060 (O_1060,N_8609,N_8814);
and UO_1061 (O_1061,N_9393,N_9085);
nand UO_1062 (O_1062,N_8703,N_9380);
and UO_1063 (O_1063,N_9343,N_9735);
nor UO_1064 (O_1064,N_8737,N_8466);
and UO_1065 (O_1065,N_9557,N_8084);
nand UO_1066 (O_1066,N_8478,N_9875);
and UO_1067 (O_1067,N_9200,N_8747);
or UO_1068 (O_1068,N_9796,N_9267);
nand UO_1069 (O_1069,N_9619,N_9921);
or UO_1070 (O_1070,N_8965,N_8767);
nor UO_1071 (O_1071,N_8567,N_9040);
xor UO_1072 (O_1072,N_9571,N_8081);
xnor UO_1073 (O_1073,N_9549,N_9129);
or UO_1074 (O_1074,N_8546,N_9909);
xor UO_1075 (O_1075,N_8393,N_8571);
nand UO_1076 (O_1076,N_9080,N_9698);
nand UO_1077 (O_1077,N_9748,N_8379);
nor UO_1078 (O_1078,N_8980,N_9868);
nor UO_1079 (O_1079,N_8028,N_9905);
nand UO_1080 (O_1080,N_8570,N_8065);
xnor UO_1081 (O_1081,N_8861,N_8073);
or UO_1082 (O_1082,N_8809,N_8369);
or UO_1083 (O_1083,N_8460,N_8352);
nor UO_1084 (O_1084,N_8559,N_9075);
or UO_1085 (O_1085,N_9731,N_8580);
xor UO_1086 (O_1086,N_9992,N_9895);
xnor UO_1087 (O_1087,N_8378,N_9836);
or UO_1088 (O_1088,N_8307,N_9953);
xor UO_1089 (O_1089,N_8103,N_8840);
nand UO_1090 (O_1090,N_8707,N_9872);
nand UO_1091 (O_1091,N_8231,N_8174);
or UO_1092 (O_1092,N_9217,N_9529);
and UO_1093 (O_1093,N_8590,N_8114);
nor UO_1094 (O_1094,N_8738,N_8565);
xor UO_1095 (O_1095,N_9326,N_9702);
and UO_1096 (O_1096,N_9126,N_9705);
or UO_1097 (O_1097,N_8566,N_9706);
nand UO_1098 (O_1098,N_8117,N_8932);
nand UO_1099 (O_1099,N_8053,N_8064);
and UO_1100 (O_1100,N_8501,N_8269);
nor UO_1101 (O_1101,N_8608,N_9181);
or UO_1102 (O_1102,N_9012,N_9432);
xnor UO_1103 (O_1103,N_9299,N_8529);
nor UO_1104 (O_1104,N_8168,N_8279);
and UO_1105 (O_1105,N_8817,N_9686);
nor UO_1106 (O_1106,N_8642,N_8990);
or UO_1107 (O_1107,N_8030,N_9339);
nand UO_1108 (O_1108,N_8469,N_8400);
xnor UO_1109 (O_1109,N_8476,N_8612);
and UO_1110 (O_1110,N_9241,N_9449);
and UO_1111 (O_1111,N_8986,N_8404);
xor UO_1112 (O_1112,N_9741,N_8795);
nand UO_1113 (O_1113,N_9913,N_9302);
and UO_1114 (O_1114,N_8423,N_9034);
or UO_1115 (O_1115,N_8411,N_8434);
xnor UO_1116 (O_1116,N_9412,N_9884);
xnor UO_1117 (O_1117,N_9407,N_9250);
nand UO_1118 (O_1118,N_9449,N_9606);
or UO_1119 (O_1119,N_8868,N_9567);
and UO_1120 (O_1120,N_9801,N_9701);
and UO_1121 (O_1121,N_8007,N_8615);
nor UO_1122 (O_1122,N_9660,N_8448);
xor UO_1123 (O_1123,N_9520,N_8321);
nor UO_1124 (O_1124,N_8393,N_8104);
nand UO_1125 (O_1125,N_9664,N_8580);
xor UO_1126 (O_1126,N_9086,N_9082);
xnor UO_1127 (O_1127,N_8967,N_9809);
xnor UO_1128 (O_1128,N_8894,N_8823);
nand UO_1129 (O_1129,N_8274,N_8032);
and UO_1130 (O_1130,N_9951,N_9642);
nor UO_1131 (O_1131,N_9703,N_8930);
and UO_1132 (O_1132,N_8648,N_8896);
nor UO_1133 (O_1133,N_8035,N_9822);
nand UO_1134 (O_1134,N_9796,N_9454);
or UO_1135 (O_1135,N_9981,N_9282);
nor UO_1136 (O_1136,N_9377,N_8394);
and UO_1137 (O_1137,N_9776,N_8251);
xor UO_1138 (O_1138,N_8385,N_8986);
or UO_1139 (O_1139,N_9690,N_9409);
xnor UO_1140 (O_1140,N_8951,N_9112);
or UO_1141 (O_1141,N_8107,N_8909);
or UO_1142 (O_1142,N_8898,N_9740);
nor UO_1143 (O_1143,N_8783,N_8819);
and UO_1144 (O_1144,N_9133,N_8971);
xor UO_1145 (O_1145,N_9860,N_9877);
xnor UO_1146 (O_1146,N_9244,N_9224);
nor UO_1147 (O_1147,N_9669,N_8343);
nand UO_1148 (O_1148,N_8892,N_9054);
nor UO_1149 (O_1149,N_8093,N_9516);
or UO_1150 (O_1150,N_9441,N_9484);
xor UO_1151 (O_1151,N_9041,N_8101);
and UO_1152 (O_1152,N_9269,N_8696);
and UO_1153 (O_1153,N_8219,N_9339);
xor UO_1154 (O_1154,N_9832,N_9619);
nand UO_1155 (O_1155,N_9448,N_8108);
nand UO_1156 (O_1156,N_9574,N_8018);
and UO_1157 (O_1157,N_8193,N_9998);
nor UO_1158 (O_1158,N_9969,N_9957);
or UO_1159 (O_1159,N_9245,N_9820);
nor UO_1160 (O_1160,N_8417,N_9374);
or UO_1161 (O_1161,N_8565,N_8294);
nand UO_1162 (O_1162,N_9699,N_8991);
nor UO_1163 (O_1163,N_8332,N_9707);
and UO_1164 (O_1164,N_8221,N_9988);
xnor UO_1165 (O_1165,N_9968,N_9484);
nor UO_1166 (O_1166,N_9348,N_9915);
or UO_1167 (O_1167,N_8045,N_9787);
or UO_1168 (O_1168,N_8161,N_8708);
and UO_1169 (O_1169,N_9937,N_8458);
xnor UO_1170 (O_1170,N_8882,N_8495);
xor UO_1171 (O_1171,N_8450,N_9506);
nand UO_1172 (O_1172,N_8172,N_9962);
nand UO_1173 (O_1173,N_9303,N_8726);
and UO_1174 (O_1174,N_9947,N_9845);
or UO_1175 (O_1175,N_9444,N_9476);
or UO_1176 (O_1176,N_9738,N_8638);
and UO_1177 (O_1177,N_9913,N_8488);
nand UO_1178 (O_1178,N_9555,N_8283);
xor UO_1179 (O_1179,N_8642,N_9049);
or UO_1180 (O_1180,N_8365,N_8293);
xnor UO_1181 (O_1181,N_8152,N_8284);
and UO_1182 (O_1182,N_8004,N_9458);
or UO_1183 (O_1183,N_8759,N_9444);
nand UO_1184 (O_1184,N_8020,N_8205);
nand UO_1185 (O_1185,N_8367,N_8900);
or UO_1186 (O_1186,N_9155,N_8290);
or UO_1187 (O_1187,N_8036,N_9377);
nor UO_1188 (O_1188,N_9218,N_8083);
or UO_1189 (O_1189,N_9748,N_9488);
and UO_1190 (O_1190,N_8131,N_9300);
and UO_1191 (O_1191,N_8262,N_9646);
and UO_1192 (O_1192,N_8929,N_8740);
nand UO_1193 (O_1193,N_8879,N_8638);
xor UO_1194 (O_1194,N_9260,N_8685);
nand UO_1195 (O_1195,N_8081,N_9938);
and UO_1196 (O_1196,N_9322,N_8228);
nand UO_1197 (O_1197,N_8892,N_8430);
and UO_1198 (O_1198,N_9959,N_9393);
or UO_1199 (O_1199,N_8876,N_9510);
xnor UO_1200 (O_1200,N_8922,N_9167);
nor UO_1201 (O_1201,N_8126,N_8651);
xnor UO_1202 (O_1202,N_9122,N_8065);
or UO_1203 (O_1203,N_8026,N_8071);
or UO_1204 (O_1204,N_9562,N_8651);
or UO_1205 (O_1205,N_8245,N_9220);
and UO_1206 (O_1206,N_9947,N_9149);
nand UO_1207 (O_1207,N_8749,N_9050);
or UO_1208 (O_1208,N_9957,N_9931);
nand UO_1209 (O_1209,N_8004,N_8044);
or UO_1210 (O_1210,N_9095,N_9170);
or UO_1211 (O_1211,N_9440,N_9045);
nor UO_1212 (O_1212,N_9067,N_8855);
nand UO_1213 (O_1213,N_9857,N_8728);
nand UO_1214 (O_1214,N_8797,N_8202);
xnor UO_1215 (O_1215,N_9235,N_9044);
and UO_1216 (O_1216,N_9647,N_8753);
nand UO_1217 (O_1217,N_9187,N_8786);
xor UO_1218 (O_1218,N_9249,N_8511);
or UO_1219 (O_1219,N_8230,N_9532);
and UO_1220 (O_1220,N_9211,N_8690);
nand UO_1221 (O_1221,N_8831,N_9152);
and UO_1222 (O_1222,N_9779,N_9812);
or UO_1223 (O_1223,N_9195,N_8212);
and UO_1224 (O_1224,N_8459,N_8619);
nand UO_1225 (O_1225,N_8000,N_9906);
and UO_1226 (O_1226,N_9824,N_9763);
or UO_1227 (O_1227,N_9848,N_9731);
or UO_1228 (O_1228,N_8383,N_9689);
nand UO_1229 (O_1229,N_8139,N_9993);
xnor UO_1230 (O_1230,N_9709,N_8971);
nor UO_1231 (O_1231,N_8278,N_8812);
nand UO_1232 (O_1232,N_8796,N_8510);
nor UO_1233 (O_1233,N_8253,N_8836);
or UO_1234 (O_1234,N_9849,N_8594);
and UO_1235 (O_1235,N_8539,N_9694);
nor UO_1236 (O_1236,N_9924,N_8919);
xnor UO_1237 (O_1237,N_8148,N_8703);
xnor UO_1238 (O_1238,N_9489,N_8947);
nor UO_1239 (O_1239,N_9125,N_9578);
and UO_1240 (O_1240,N_9652,N_9488);
and UO_1241 (O_1241,N_9439,N_9519);
and UO_1242 (O_1242,N_9482,N_8475);
and UO_1243 (O_1243,N_9628,N_8398);
and UO_1244 (O_1244,N_8395,N_8956);
nor UO_1245 (O_1245,N_8852,N_9887);
or UO_1246 (O_1246,N_8441,N_9399);
nand UO_1247 (O_1247,N_8469,N_8729);
nor UO_1248 (O_1248,N_8446,N_8256);
nand UO_1249 (O_1249,N_9862,N_9492);
and UO_1250 (O_1250,N_8611,N_9020);
and UO_1251 (O_1251,N_9108,N_8268);
or UO_1252 (O_1252,N_8072,N_9461);
nand UO_1253 (O_1253,N_9210,N_8778);
xnor UO_1254 (O_1254,N_9948,N_8225);
and UO_1255 (O_1255,N_8661,N_8570);
nor UO_1256 (O_1256,N_8257,N_9564);
nand UO_1257 (O_1257,N_9968,N_8575);
xor UO_1258 (O_1258,N_9300,N_9761);
xor UO_1259 (O_1259,N_9316,N_9971);
nor UO_1260 (O_1260,N_9218,N_8890);
nor UO_1261 (O_1261,N_8252,N_8353);
nand UO_1262 (O_1262,N_8110,N_8930);
or UO_1263 (O_1263,N_9674,N_8973);
nand UO_1264 (O_1264,N_9667,N_9768);
nand UO_1265 (O_1265,N_9106,N_9616);
nand UO_1266 (O_1266,N_9522,N_8877);
or UO_1267 (O_1267,N_9870,N_9667);
nand UO_1268 (O_1268,N_9508,N_8410);
nand UO_1269 (O_1269,N_9220,N_8309);
and UO_1270 (O_1270,N_9298,N_9492);
nor UO_1271 (O_1271,N_9486,N_8782);
xnor UO_1272 (O_1272,N_9453,N_9685);
nor UO_1273 (O_1273,N_9109,N_8151);
nand UO_1274 (O_1274,N_9623,N_8711);
and UO_1275 (O_1275,N_9481,N_9515);
or UO_1276 (O_1276,N_9648,N_8326);
and UO_1277 (O_1277,N_8463,N_9046);
xnor UO_1278 (O_1278,N_9201,N_8371);
or UO_1279 (O_1279,N_8339,N_8232);
nor UO_1280 (O_1280,N_9776,N_8918);
xnor UO_1281 (O_1281,N_8954,N_8588);
nor UO_1282 (O_1282,N_9226,N_8084);
and UO_1283 (O_1283,N_9675,N_9802);
or UO_1284 (O_1284,N_8485,N_8712);
or UO_1285 (O_1285,N_8852,N_8229);
xor UO_1286 (O_1286,N_9487,N_8501);
and UO_1287 (O_1287,N_8779,N_8247);
and UO_1288 (O_1288,N_9536,N_9153);
nand UO_1289 (O_1289,N_8468,N_8427);
nand UO_1290 (O_1290,N_8755,N_9392);
and UO_1291 (O_1291,N_9804,N_9699);
xor UO_1292 (O_1292,N_9881,N_8382);
xnor UO_1293 (O_1293,N_8482,N_9036);
and UO_1294 (O_1294,N_9144,N_8218);
nand UO_1295 (O_1295,N_8383,N_9007);
or UO_1296 (O_1296,N_8916,N_8249);
xor UO_1297 (O_1297,N_9109,N_8140);
xor UO_1298 (O_1298,N_9998,N_8671);
nor UO_1299 (O_1299,N_9197,N_8487);
nor UO_1300 (O_1300,N_8601,N_9104);
and UO_1301 (O_1301,N_8310,N_8991);
xnor UO_1302 (O_1302,N_8253,N_8507);
and UO_1303 (O_1303,N_9856,N_8582);
xnor UO_1304 (O_1304,N_9389,N_9271);
or UO_1305 (O_1305,N_8782,N_8515);
xor UO_1306 (O_1306,N_8874,N_8778);
and UO_1307 (O_1307,N_9390,N_9823);
or UO_1308 (O_1308,N_9342,N_8480);
and UO_1309 (O_1309,N_9746,N_8007);
nor UO_1310 (O_1310,N_8511,N_9661);
and UO_1311 (O_1311,N_9138,N_8907);
nor UO_1312 (O_1312,N_9233,N_8465);
xor UO_1313 (O_1313,N_9346,N_8321);
and UO_1314 (O_1314,N_8297,N_8890);
xor UO_1315 (O_1315,N_9460,N_8916);
xnor UO_1316 (O_1316,N_9969,N_8959);
nor UO_1317 (O_1317,N_9856,N_8250);
nor UO_1318 (O_1318,N_9250,N_9007);
and UO_1319 (O_1319,N_8692,N_9255);
and UO_1320 (O_1320,N_9545,N_8132);
nand UO_1321 (O_1321,N_8289,N_9363);
nand UO_1322 (O_1322,N_9511,N_8683);
nor UO_1323 (O_1323,N_9407,N_8636);
xor UO_1324 (O_1324,N_9875,N_8867);
or UO_1325 (O_1325,N_8957,N_9917);
and UO_1326 (O_1326,N_9684,N_8847);
xnor UO_1327 (O_1327,N_9406,N_8988);
and UO_1328 (O_1328,N_8291,N_9497);
nor UO_1329 (O_1329,N_9720,N_8141);
nand UO_1330 (O_1330,N_9639,N_9496);
nor UO_1331 (O_1331,N_8707,N_8540);
nand UO_1332 (O_1332,N_9274,N_8814);
nand UO_1333 (O_1333,N_8345,N_8904);
xor UO_1334 (O_1334,N_9675,N_9765);
xnor UO_1335 (O_1335,N_8412,N_9648);
nor UO_1336 (O_1336,N_9682,N_8351);
xnor UO_1337 (O_1337,N_9402,N_8599);
and UO_1338 (O_1338,N_9090,N_9932);
xor UO_1339 (O_1339,N_9064,N_9727);
and UO_1340 (O_1340,N_9659,N_9651);
nand UO_1341 (O_1341,N_8094,N_9309);
nor UO_1342 (O_1342,N_8432,N_8697);
or UO_1343 (O_1343,N_9099,N_9199);
nand UO_1344 (O_1344,N_9167,N_8281);
and UO_1345 (O_1345,N_9868,N_9926);
nand UO_1346 (O_1346,N_9584,N_8124);
or UO_1347 (O_1347,N_9607,N_8386);
xor UO_1348 (O_1348,N_9688,N_9624);
xnor UO_1349 (O_1349,N_8378,N_8389);
or UO_1350 (O_1350,N_8502,N_8428);
and UO_1351 (O_1351,N_9170,N_8804);
nand UO_1352 (O_1352,N_8776,N_8073);
or UO_1353 (O_1353,N_8025,N_9680);
or UO_1354 (O_1354,N_9861,N_8489);
or UO_1355 (O_1355,N_8187,N_8866);
nor UO_1356 (O_1356,N_8452,N_9581);
xnor UO_1357 (O_1357,N_9425,N_9567);
nor UO_1358 (O_1358,N_9457,N_9827);
and UO_1359 (O_1359,N_9417,N_8366);
nand UO_1360 (O_1360,N_9887,N_9952);
nor UO_1361 (O_1361,N_8089,N_9283);
and UO_1362 (O_1362,N_9320,N_8223);
xnor UO_1363 (O_1363,N_8971,N_9648);
or UO_1364 (O_1364,N_9853,N_9144);
nor UO_1365 (O_1365,N_8235,N_9958);
and UO_1366 (O_1366,N_9383,N_8686);
nand UO_1367 (O_1367,N_8541,N_8721);
or UO_1368 (O_1368,N_8668,N_8294);
xor UO_1369 (O_1369,N_9538,N_9890);
and UO_1370 (O_1370,N_9533,N_9446);
xnor UO_1371 (O_1371,N_8163,N_9201);
nand UO_1372 (O_1372,N_8323,N_9489);
xor UO_1373 (O_1373,N_9489,N_9851);
xnor UO_1374 (O_1374,N_8693,N_8095);
and UO_1375 (O_1375,N_8467,N_8247);
and UO_1376 (O_1376,N_8441,N_8993);
xnor UO_1377 (O_1377,N_9993,N_9633);
and UO_1378 (O_1378,N_8398,N_8308);
and UO_1379 (O_1379,N_8166,N_8921);
nor UO_1380 (O_1380,N_8414,N_9998);
nand UO_1381 (O_1381,N_9639,N_9579);
or UO_1382 (O_1382,N_8305,N_8406);
nand UO_1383 (O_1383,N_9984,N_9780);
and UO_1384 (O_1384,N_9898,N_8876);
or UO_1385 (O_1385,N_8815,N_9484);
and UO_1386 (O_1386,N_9279,N_9980);
xnor UO_1387 (O_1387,N_8358,N_9403);
or UO_1388 (O_1388,N_8078,N_9409);
nor UO_1389 (O_1389,N_8511,N_9485);
and UO_1390 (O_1390,N_9412,N_9363);
and UO_1391 (O_1391,N_9091,N_8348);
nor UO_1392 (O_1392,N_9790,N_9162);
nand UO_1393 (O_1393,N_9497,N_9766);
nand UO_1394 (O_1394,N_8215,N_8108);
and UO_1395 (O_1395,N_9734,N_9310);
xor UO_1396 (O_1396,N_9492,N_8130);
nor UO_1397 (O_1397,N_8102,N_8183);
nor UO_1398 (O_1398,N_8226,N_9901);
or UO_1399 (O_1399,N_8290,N_9321);
and UO_1400 (O_1400,N_9538,N_8547);
and UO_1401 (O_1401,N_9201,N_9608);
xor UO_1402 (O_1402,N_8322,N_9822);
and UO_1403 (O_1403,N_8370,N_9853);
or UO_1404 (O_1404,N_8045,N_8680);
xnor UO_1405 (O_1405,N_9443,N_9866);
or UO_1406 (O_1406,N_9356,N_9869);
or UO_1407 (O_1407,N_9535,N_8379);
nor UO_1408 (O_1408,N_9148,N_8584);
or UO_1409 (O_1409,N_9002,N_9325);
nor UO_1410 (O_1410,N_8435,N_9925);
or UO_1411 (O_1411,N_9186,N_8455);
nor UO_1412 (O_1412,N_9788,N_9995);
xnor UO_1413 (O_1413,N_9108,N_8465);
nand UO_1414 (O_1414,N_8366,N_8400);
xnor UO_1415 (O_1415,N_8583,N_8864);
nor UO_1416 (O_1416,N_8016,N_8413);
and UO_1417 (O_1417,N_8918,N_9379);
nand UO_1418 (O_1418,N_9669,N_9198);
and UO_1419 (O_1419,N_9528,N_8678);
and UO_1420 (O_1420,N_8096,N_8474);
nor UO_1421 (O_1421,N_9753,N_8136);
nand UO_1422 (O_1422,N_8800,N_8415);
nor UO_1423 (O_1423,N_8520,N_8859);
nor UO_1424 (O_1424,N_8975,N_9554);
xor UO_1425 (O_1425,N_8640,N_9833);
nand UO_1426 (O_1426,N_9453,N_8559);
nor UO_1427 (O_1427,N_8939,N_8517);
nor UO_1428 (O_1428,N_8915,N_8839);
or UO_1429 (O_1429,N_9169,N_9382);
and UO_1430 (O_1430,N_9782,N_9268);
nor UO_1431 (O_1431,N_8388,N_9504);
nor UO_1432 (O_1432,N_8654,N_9619);
nor UO_1433 (O_1433,N_8821,N_8960);
nand UO_1434 (O_1434,N_9676,N_8094);
nand UO_1435 (O_1435,N_9005,N_9280);
or UO_1436 (O_1436,N_8513,N_8183);
or UO_1437 (O_1437,N_8746,N_8648);
or UO_1438 (O_1438,N_8414,N_8556);
xor UO_1439 (O_1439,N_8334,N_9806);
nor UO_1440 (O_1440,N_8712,N_9469);
nand UO_1441 (O_1441,N_8461,N_8762);
nand UO_1442 (O_1442,N_9753,N_8284);
nand UO_1443 (O_1443,N_8165,N_9864);
or UO_1444 (O_1444,N_8310,N_8136);
nand UO_1445 (O_1445,N_9933,N_9466);
or UO_1446 (O_1446,N_9230,N_8979);
xor UO_1447 (O_1447,N_9296,N_9839);
nor UO_1448 (O_1448,N_9828,N_8425);
nor UO_1449 (O_1449,N_8833,N_9676);
and UO_1450 (O_1450,N_8336,N_9895);
nor UO_1451 (O_1451,N_9823,N_8904);
or UO_1452 (O_1452,N_8476,N_9312);
xnor UO_1453 (O_1453,N_9507,N_8110);
xor UO_1454 (O_1454,N_8309,N_9606);
nor UO_1455 (O_1455,N_9897,N_9179);
and UO_1456 (O_1456,N_9636,N_8254);
or UO_1457 (O_1457,N_9558,N_8531);
xor UO_1458 (O_1458,N_8146,N_9133);
nor UO_1459 (O_1459,N_9682,N_9491);
nor UO_1460 (O_1460,N_9497,N_8982);
or UO_1461 (O_1461,N_9827,N_9380);
nand UO_1462 (O_1462,N_9943,N_8067);
or UO_1463 (O_1463,N_8332,N_9142);
nor UO_1464 (O_1464,N_8078,N_9341);
and UO_1465 (O_1465,N_9625,N_8938);
nor UO_1466 (O_1466,N_9942,N_8333);
and UO_1467 (O_1467,N_8283,N_9256);
xnor UO_1468 (O_1468,N_8799,N_8974);
or UO_1469 (O_1469,N_8353,N_9569);
nand UO_1470 (O_1470,N_8667,N_8345);
or UO_1471 (O_1471,N_8483,N_9618);
xor UO_1472 (O_1472,N_8032,N_9111);
xnor UO_1473 (O_1473,N_9510,N_8064);
nand UO_1474 (O_1474,N_9437,N_8756);
or UO_1475 (O_1475,N_9581,N_8619);
or UO_1476 (O_1476,N_8290,N_8061);
nor UO_1477 (O_1477,N_9609,N_9708);
nor UO_1478 (O_1478,N_8389,N_9626);
nand UO_1479 (O_1479,N_8755,N_9715);
nand UO_1480 (O_1480,N_8919,N_9090);
and UO_1481 (O_1481,N_8901,N_9714);
xnor UO_1482 (O_1482,N_8361,N_8124);
or UO_1483 (O_1483,N_9164,N_9641);
nand UO_1484 (O_1484,N_9429,N_9687);
and UO_1485 (O_1485,N_8498,N_8815);
nand UO_1486 (O_1486,N_9256,N_8335);
nor UO_1487 (O_1487,N_8910,N_9980);
nor UO_1488 (O_1488,N_8652,N_9084);
nor UO_1489 (O_1489,N_9274,N_8916);
nand UO_1490 (O_1490,N_8058,N_9592);
xnor UO_1491 (O_1491,N_9993,N_9641);
or UO_1492 (O_1492,N_8889,N_8977);
nor UO_1493 (O_1493,N_8265,N_9414);
nor UO_1494 (O_1494,N_8222,N_9535);
xor UO_1495 (O_1495,N_9820,N_8123);
xnor UO_1496 (O_1496,N_8460,N_9334);
nor UO_1497 (O_1497,N_9919,N_8115);
and UO_1498 (O_1498,N_8376,N_8805);
nor UO_1499 (O_1499,N_9567,N_9038);
endmodule