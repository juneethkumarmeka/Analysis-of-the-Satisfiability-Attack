module basic_500_3000_500_6_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_68,In_25);
nand U1 (N_1,In_433,In_199);
or U2 (N_2,In_97,In_447);
or U3 (N_3,In_232,In_268);
or U4 (N_4,In_55,In_23);
nor U5 (N_5,In_468,In_435);
or U6 (N_6,In_17,In_34);
and U7 (N_7,In_77,In_186);
and U8 (N_8,In_273,In_93);
nand U9 (N_9,In_260,In_166);
and U10 (N_10,In_480,In_12);
and U11 (N_11,In_109,In_177);
and U12 (N_12,In_382,In_277);
and U13 (N_13,In_400,In_123);
nand U14 (N_14,In_308,In_137);
nor U15 (N_15,In_42,In_88);
nand U16 (N_16,In_191,In_290);
and U17 (N_17,In_224,In_271);
and U18 (N_18,In_487,In_147);
or U19 (N_19,In_262,In_154);
and U20 (N_20,In_194,In_252);
nand U21 (N_21,In_402,In_14);
nand U22 (N_22,In_218,In_391);
nand U23 (N_23,In_448,In_48);
xnor U24 (N_24,In_427,In_420);
and U25 (N_25,In_225,In_295);
xnor U26 (N_26,In_496,In_170);
nor U27 (N_27,In_43,In_160);
and U28 (N_28,In_326,In_19);
or U29 (N_29,In_263,In_60);
nor U30 (N_30,In_78,In_356);
and U31 (N_31,In_318,In_426);
or U32 (N_32,In_393,In_234);
and U33 (N_33,In_296,In_338);
or U34 (N_34,In_139,In_297);
nand U35 (N_35,In_182,In_413);
nand U36 (N_36,In_67,In_334);
or U37 (N_37,In_464,In_302);
or U38 (N_38,In_482,In_134);
nand U39 (N_39,In_370,In_229);
nand U40 (N_40,In_203,In_398);
or U41 (N_41,In_327,In_264);
nor U42 (N_42,In_21,In_220);
nor U43 (N_43,In_465,In_140);
or U44 (N_44,In_153,In_332);
nand U45 (N_45,In_399,In_462);
nand U46 (N_46,In_15,In_415);
or U47 (N_47,In_226,In_345);
or U48 (N_48,In_243,In_138);
and U49 (N_49,In_281,In_24);
nor U50 (N_50,In_176,In_411);
nor U51 (N_51,In_171,In_418);
nand U52 (N_52,In_275,In_286);
and U53 (N_53,In_364,In_16);
or U54 (N_54,In_127,In_189);
or U55 (N_55,In_294,In_28);
nand U56 (N_56,In_86,In_394);
nor U57 (N_57,In_269,In_217);
nand U58 (N_58,In_158,In_52);
nor U59 (N_59,In_27,In_183);
nor U60 (N_60,In_279,In_4);
or U61 (N_61,In_13,In_471);
and U62 (N_62,In_278,In_51);
or U63 (N_63,In_472,In_256);
nor U64 (N_64,In_227,In_467);
or U65 (N_65,In_397,In_131);
xor U66 (N_66,In_358,In_436);
nor U67 (N_67,In_246,In_307);
nand U68 (N_68,In_247,In_304);
or U69 (N_69,In_211,In_144);
or U70 (N_70,In_421,In_301);
or U71 (N_71,In_309,In_417);
xnor U72 (N_72,In_22,In_253);
nand U73 (N_73,In_54,In_280);
nand U74 (N_74,In_444,In_317);
nand U75 (N_75,In_344,In_352);
nand U76 (N_76,In_493,In_282);
and U77 (N_77,In_135,In_126);
or U78 (N_78,In_483,In_141);
and U79 (N_79,In_221,In_156);
nand U80 (N_80,In_75,In_384);
and U81 (N_81,In_452,In_456);
nand U82 (N_82,In_132,In_405);
nor U83 (N_83,In_474,In_486);
or U84 (N_84,In_213,In_347);
nand U85 (N_85,In_133,In_437);
nand U86 (N_86,In_209,In_178);
or U87 (N_87,In_212,In_38);
nand U88 (N_88,In_89,In_155);
nand U89 (N_89,In_136,In_162);
nand U90 (N_90,In_195,In_336);
and U91 (N_91,In_443,In_115);
nor U92 (N_92,In_216,In_241);
nand U93 (N_93,In_390,In_414);
xor U94 (N_94,In_129,In_254);
nor U95 (N_95,In_198,In_303);
nor U96 (N_96,In_335,In_44);
nand U97 (N_97,In_128,In_32);
or U98 (N_98,In_149,In_258);
and U99 (N_99,In_355,In_222);
nand U100 (N_100,In_320,In_428);
nand U101 (N_101,In_407,In_276);
nor U102 (N_102,In_284,In_492);
and U103 (N_103,In_380,In_120);
or U104 (N_104,In_261,In_200);
nor U105 (N_105,In_378,In_267);
and U106 (N_106,In_70,In_197);
and U107 (N_107,In_112,In_94);
or U108 (N_108,In_210,In_328);
nand U109 (N_109,In_499,In_432);
or U110 (N_110,In_342,In_466);
nor U111 (N_111,In_442,In_72);
or U112 (N_112,In_40,In_419);
or U113 (N_113,In_103,In_354);
or U114 (N_114,In_375,In_481);
and U115 (N_115,In_11,In_59);
nand U116 (N_116,In_497,In_409);
nor U117 (N_117,In_161,In_130);
xor U118 (N_118,In_396,In_385);
nand U119 (N_119,In_461,In_62);
nand U120 (N_120,In_376,In_325);
and U121 (N_121,In_498,In_239);
nor U122 (N_122,In_469,In_35);
or U123 (N_123,In_477,In_116);
and U124 (N_124,In_406,In_163);
and U125 (N_125,In_313,In_323);
or U126 (N_126,In_248,In_5);
or U127 (N_127,In_47,In_315);
and U128 (N_128,In_41,In_124);
or U129 (N_129,In_7,In_272);
xnor U130 (N_130,In_157,In_306);
or U131 (N_131,In_20,In_83);
or U132 (N_132,In_202,In_455);
nand U133 (N_133,In_244,In_374);
or U134 (N_134,In_228,In_33);
or U135 (N_135,In_37,In_236);
or U136 (N_136,In_441,In_90);
nand U137 (N_137,In_412,In_117);
nand U138 (N_138,In_285,In_288);
or U139 (N_139,In_172,In_167);
nor U140 (N_140,In_484,In_363);
nand U141 (N_141,In_460,In_395);
or U142 (N_142,In_489,In_53);
nor U143 (N_143,In_353,In_99);
and U144 (N_144,In_289,In_9);
or U145 (N_145,In_274,In_491);
and U146 (N_146,In_312,In_322);
nand U147 (N_147,In_381,In_410);
or U148 (N_148,In_449,In_488);
or U149 (N_149,In_39,In_180);
and U150 (N_150,In_235,In_367);
nand U151 (N_151,In_259,In_425);
or U152 (N_152,In_291,In_187);
nand U153 (N_153,In_207,In_388);
nor U154 (N_154,In_168,In_142);
or U155 (N_155,In_190,In_416);
or U156 (N_156,In_429,In_185);
or U157 (N_157,In_80,In_192);
nor U158 (N_158,In_230,In_362);
nor U159 (N_159,In_79,In_446);
and U160 (N_160,In_100,In_65);
or U161 (N_161,In_6,In_205);
or U162 (N_162,In_386,In_404);
nand U163 (N_163,In_283,In_26);
nor U164 (N_164,In_340,In_74);
and U165 (N_165,In_169,In_184);
nand U166 (N_166,In_101,In_82);
nand U167 (N_167,In_341,In_423);
nand U168 (N_168,In_445,In_403);
or U169 (N_169,In_18,In_463);
nand U170 (N_170,In_470,In_76);
nand U171 (N_171,In_331,In_359);
and U172 (N_172,In_125,In_3);
and U173 (N_173,In_453,In_343);
or U174 (N_174,In_434,In_196);
or U175 (N_175,In_0,In_150);
nand U176 (N_176,In_193,In_392);
nor U177 (N_177,In_95,In_494);
or U178 (N_178,In_475,In_250);
nor U179 (N_179,In_206,In_57);
nand U180 (N_180,In_201,In_321);
nand U181 (N_181,In_151,In_238);
nand U182 (N_182,In_91,In_245);
or U183 (N_183,In_270,In_36);
nand U184 (N_184,In_73,In_173);
nor U185 (N_185,In_377,In_164);
xor U186 (N_186,In_350,In_121);
nor U187 (N_187,In_108,In_451);
or U188 (N_188,In_237,In_365);
nand U189 (N_189,In_310,In_31);
or U190 (N_190,In_348,In_383);
nand U191 (N_191,In_122,In_119);
or U192 (N_192,In_64,In_58);
nor U193 (N_193,In_152,In_188);
and U194 (N_194,In_66,In_145);
or U195 (N_195,In_458,In_159);
or U196 (N_196,In_476,In_351);
nor U197 (N_197,In_118,In_85);
and U198 (N_198,In_104,In_242);
and U199 (N_199,In_479,In_287);
and U200 (N_200,In_495,In_56);
nand U201 (N_201,In_450,In_179);
nor U202 (N_202,In_454,In_69);
nand U203 (N_203,In_255,In_324);
nor U204 (N_204,In_2,In_249);
nor U205 (N_205,In_457,In_369);
nor U206 (N_206,In_231,In_81);
nand U207 (N_207,In_368,In_175);
nor U208 (N_208,In_379,In_146);
or U209 (N_209,In_63,In_424);
nand U210 (N_210,In_114,In_387);
nor U211 (N_211,In_329,In_438);
nand U212 (N_212,In_357,In_143);
nor U213 (N_213,In_110,In_339);
and U214 (N_214,In_430,In_107);
or U215 (N_215,In_490,In_371);
or U216 (N_216,In_305,In_148);
and U217 (N_217,In_111,In_113);
nand U218 (N_218,In_314,In_174);
and U219 (N_219,In_298,In_46);
and U220 (N_220,In_106,In_214);
and U221 (N_221,In_408,In_8);
and U222 (N_222,In_373,In_29);
or U223 (N_223,In_440,In_366);
nor U224 (N_224,In_372,In_257);
and U225 (N_225,In_319,In_215);
nand U226 (N_226,In_299,In_10);
nand U227 (N_227,In_181,In_422);
nor U228 (N_228,In_300,In_96);
and U229 (N_229,In_485,In_360);
or U230 (N_230,In_219,In_333);
nand U231 (N_231,In_204,In_346);
nor U232 (N_232,In_233,In_316);
or U233 (N_233,In_98,In_478);
nor U234 (N_234,In_105,In_102);
and U235 (N_235,In_349,In_30);
nand U236 (N_236,In_266,In_330);
nand U237 (N_237,In_361,In_45);
and U238 (N_238,In_389,In_84);
or U239 (N_239,In_311,In_165);
and U240 (N_240,In_401,In_473);
nor U241 (N_241,In_459,In_71);
and U242 (N_242,In_439,In_431);
nand U243 (N_243,In_208,In_49);
nor U244 (N_244,In_87,In_251);
or U245 (N_245,In_293,In_61);
nor U246 (N_246,In_92,In_292);
and U247 (N_247,In_337,In_223);
nand U248 (N_248,In_50,In_1);
nor U249 (N_249,In_240,In_265);
or U250 (N_250,In_114,In_149);
xnor U251 (N_251,In_209,In_155);
nand U252 (N_252,In_95,In_146);
and U253 (N_253,In_205,In_278);
nand U254 (N_254,In_345,In_182);
or U255 (N_255,In_410,In_203);
or U256 (N_256,In_432,In_454);
or U257 (N_257,In_359,In_89);
nand U258 (N_258,In_180,In_489);
or U259 (N_259,In_200,In_499);
and U260 (N_260,In_227,In_92);
or U261 (N_261,In_423,In_337);
nand U262 (N_262,In_166,In_91);
nand U263 (N_263,In_408,In_273);
xnor U264 (N_264,In_31,In_47);
and U265 (N_265,In_299,In_116);
nor U266 (N_266,In_333,In_336);
nand U267 (N_267,In_468,In_426);
or U268 (N_268,In_183,In_293);
nand U269 (N_269,In_410,In_77);
nand U270 (N_270,In_410,In_25);
or U271 (N_271,In_170,In_238);
or U272 (N_272,In_305,In_368);
nand U273 (N_273,In_498,In_150);
and U274 (N_274,In_192,In_245);
nor U275 (N_275,In_369,In_367);
nor U276 (N_276,In_132,In_262);
or U277 (N_277,In_42,In_315);
or U278 (N_278,In_180,In_257);
nor U279 (N_279,In_426,In_158);
and U280 (N_280,In_8,In_21);
or U281 (N_281,In_44,In_104);
or U282 (N_282,In_0,In_326);
or U283 (N_283,In_21,In_200);
or U284 (N_284,In_165,In_332);
nor U285 (N_285,In_22,In_260);
or U286 (N_286,In_107,In_367);
nand U287 (N_287,In_60,In_326);
or U288 (N_288,In_147,In_1);
nand U289 (N_289,In_387,In_127);
nand U290 (N_290,In_52,In_364);
nand U291 (N_291,In_16,In_413);
nand U292 (N_292,In_254,In_210);
and U293 (N_293,In_34,In_114);
nor U294 (N_294,In_199,In_79);
nor U295 (N_295,In_295,In_333);
nor U296 (N_296,In_141,In_77);
or U297 (N_297,In_218,In_62);
and U298 (N_298,In_27,In_128);
nand U299 (N_299,In_148,In_493);
nor U300 (N_300,In_250,In_201);
or U301 (N_301,In_471,In_3);
nand U302 (N_302,In_98,In_372);
nand U303 (N_303,In_317,In_156);
or U304 (N_304,In_385,In_485);
or U305 (N_305,In_461,In_16);
nor U306 (N_306,In_248,In_356);
and U307 (N_307,In_12,In_451);
nand U308 (N_308,In_234,In_134);
nand U309 (N_309,In_387,In_126);
or U310 (N_310,In_408,In_14);
and U311 (N_311,In_98,In_369);
and U312 (N_312,In_43,In_306);
or U313 (N_313,In_169,In_235);
or U314 (N_314,In_36,In_320);
nor U315 (N_315,In_78,In_406);
and U316 (N_316,In_358,In_382);
or U317 (N_317,In_226,In_282);
or U318 (N_318,In_57,In_483);
or U319 (N_319,In_458,In_5);
xnor U320 (N_320,In_470,In_211);
nor U321 (N_321,In_153,In_13);
or U322 (N_322,In_243,In_446);
or U323 (N_323,In_274,In_221);
nand U324 (N_324,In_78,In_95);
or U325 (N_325,In_436,In_300);
and U326 (N_326,In_258,In_106);
or U327 (N_327,In_407,In_275);
nor U328 (N_328,In_6,In_126);
nand U329 (N_329,In_119,In_473);
or U330 (N_330,In_107,In_33);
xnor U331 (N_331,In_190,In_211);
nand U332 (N_332,In_471,In_431);
nand U333 (N_333,In_56,In_258);
nand U334 (N_334,In_195,In_68);
nor U335 (N_335,In_347,In_362);
nor U336 (N_336,In_93,In_297);
and U337 (N_337,In_189,In_338);
and U338 (N_338,In_117,In_34);
nor U339 (N_339,In_283,In_221);
or U340 (N_340,In_452,In_312);
or U341 (N_341,In_465,In_156);
nor U342 (N_342,In_52,In_31);
and U343 (N_343,In_298,In_257);
nor U344 (N_344,In_336,In_21);
or U345 (N_345,In_437,In_364);
and U346 (N_346,In_347,In_140);
nand U347 (N_347,In_401,In_51);
or U348 (N_348,In_435,In_269);
or U349 (N_349,In_16,In_123);
nand U350 (N_350,In_248,In_184);
nand U351 (N_351,In_82,In_485);
or U352 (N_352,In_133,In_481);
or U353 (N_353,In_158,In_435);
nand U354 (N_354,In_342,In_169);
nand U355 (N_355,In_324,In_28);
or U356 (N_356,In_128,In_58);
nor U357 (N_357,In_227,In_115);
nor U358 (N_358,In_120,In_199);
nand U359 (N_359,In_435,In_241);
nand U360 (N_360,In_82,In_139);
nor U361 (N_361,In_64,In_301);
or U362 (N_362,In_481,In_403);
and U363 (N_363,In_21,In_313);
xor U364 (N_364,In_389,In_87);
or U365 (N_365,In_475,In_348);
nor U366 (N_366,In_343,In_497);
and U367 (N_367,In_197,In_116);
nand U368 (N_368,In_418,In_211);
and U369 (N_369,In_13,In_496);
nand U370 (N_370,In_431,In_490);
and U371 (N_371,In_300,In_146);
nand U372 (N_372,In_223,In_284);
and U373 (N_373,In_127,In_308);
and U374 (N_374,In_398,In_453);
nor U375 (N_375,In_391,In_389);
nor U376 (N_376,In_471,In_442);
nor U377 (N_377,In_111,In_150);
nand U378 (N_378,In_407,In_321);
and U379 (N_379,In_8,In_431);
nand U380 (N_380,In_336,In_45);
and U381 (N_381,In_251,In_181);
and U382 (N_382,In_163,In_250);
nand U383 (N_383,In_67,In_192);
and U384 (N_384,In_88,In_253);
or U385 (N_385,In_344,In_167);
nand U386 (N_386,In_217,In_400);
nor U387 (N_387,In_140,In_365);
or U388 (N_388,In_123,In_316);
or U389 (N_389,In_308,In_225);
and U390 (N_390,In_200,In_449);
nor U391 (N_391,In_404,In_26);
nand U392 (N_392,In_451,In_203);
or U393 (N_393,In_262,In_77);
nand U394 (N_394,In_205,In_415);
nor U395 (N_395,In_18,In_369);
and U396 (N_396,In_129,In_240);
or U397 (N_397,In_398,In_490);
and U398 (N_398,In_364,In_192);
xnor U399 (N_399,In_359,In_75);
nor U400 (N_400,In_363,In_227);
nor U401 (N_401,In_29,In_19);
or U402 (N_402,In_462,In_158);
nand U403 (N_403,In_245,In_173);
xnor U404 (N_404,In_230,In_396);
xnor U405 (N_405,In_188,In_104);
nor U406 (N_406,In_354,In_158);
nor U407 (N_407,In_299,In_407);
or U408 (N_408,In_431,In_153);
nor U409 (N_409,In_0,In_394);
nand U410 (N_410,In_212,In_80);
and U411 (N_411,In_414,In_103);
xnor U412 (N_412,In_95,In_491);
and U413 (N_413,In_200,In_394);
and U414 (N_414,In_256,In_206);
and U415 (N_415,In_0,In_355);
or U416 (N_416,In_276,In_192);
nor U417 (N_417,In_320,In_418);
nand U418 (N_418,In_494,In_62);
or U419 (N_419,In_225,In_467);
or U420 (N_420,In_380,In_274);
nor U421 (N_421,In_166,In_269);
and U422 (N_422,In_31,In_452);
and U423 (N_423,In_223,In_425);
or U424 (N_424,In_55,In_112);
nor U425 (N_425,In_14,In_293);
and U426 (N_426,In_218,In_125);
nand U427 (N_427,In_71,In_259);
nand U428 (N_428,In_88,In_58);
or U429 (N_429,In_471,In_245);
and U430 (N_430,In_329,In_19);
or U431 (N_431,In_272,In_111);
or U432 (N_432,In_383,In_81);
xnor U433 (N_433,In_457,In_0);
nor U434 (N_434,In_158,In_115);
nand U435 (N_435,In_282,In_235);
or U436 (N_436,In_256,In_5);
xnor U437 (N_437,In_398,In_220);
nor U438 (N_438,In_217,In_193);
nor U439 (N_439,In_457,In_165);
or U440 (N_440,In_162,In_440);
nor U441 (N_441,In_405,In_339);
nor U442 (N_442,In_218,In_163);
or U443 (N_443,In_393,In_372);
and U444 (N_444,In_374,In_272);
or U445 (N_445,In_333,In_476);
and U446 (N_446,In_390,In_228);
nand U447 (N_447,In_367,In_420);
xnor U448 (N_448,In_154,In_307);
nand U449 (N_449,In_464,In_244);
and U450 (N_450,In_399,In_38);
or U451 (N_451,In_227,In_471);
nor U452 (N_452,In_209,In_88);
nor U453 (N_453,In_376,In_317);
or U454 (N_454,In_122,In_54);
nor U455 (N_455,In_248,In_51);
or U456 (N_456,In_227,In_6);
and U457 (N_457,In_499,In_478);
nand U458 (N_458,In_379,In_283);
nand U459 (N_459,In_221,In_417);
or U460 (N_460,In_174,In_331);
nand U461 (N_461,In_51,In_471);
or U462 (N_462,In_46,In_91);
and U463 (N_463,In_69,In_164);
nor U464 (N_464,In_168,In_328);
nand U465 (N_465,In_376,In_414);
nor U466 (N_466,In_170,In_77);
and U467 (N_467,In_22,In_358);
or U468 (N_468,In_174,In_156);
nor U469 (N_469,In_91,In_210);
and U470 (N_470,In_136,In_473);
and U471 (N_471,In_392,In_461);
or U472 (N_472,In_283,In_168);
and U473 (N_473,In_265,In_446);
nand U474 (N_474,In_188,In_452);
nand U475 (N_475,In_393,In_21);
and U476 (N_476,In_68,In_228);
or U477 (N_477,In_336,In_184);
or U478 (N_478,In_423,In_172);
nor U479 (N_479,In_280,In_496);
or U480 (N_480,In_280,In_389);
or U481 (N_481,In_0,In_193);
or U482 (N_482,In_319,In_179);
nor U483 (N_483,In_496,In_105);
and U484 (N_484,In_72,In_194);
nand U485 (N_485,In_77,In_112);
nor U486 (N_486,In_282,In_5);
and U487 (N_487,In_427,In_380);
nor U488 (N_488,In_219,In_278);
or U489 (N_489,In_76,In_129);
or U490 (N_490,In_445,In_2);
and U491 (N_491,In_54,In_453);
nor U492 (N_492,In_385,In_164);
nand U493 (N_493,In_325,In_145);
nand U494 (N_494,In_3,In_193);
nand U495 (N_495,In_25,In_271);
xor U496 (N_496,In_487,In_444);
and U497 (N_497,In_313,In_113);
and U498 (N_498,In_399,In_143);
and U499 (N_499,In_459,In_55);
and U500 (N_500,N_231,N_135);
or U501 (N_501,N_441,N_218);
nand U502 (N_502,N_212,N_484);
nand U503 (N_503,N_423,N_146);
or U504 (N_504,N_442,N_387);
nand U505 (N_505,N_289,N_15);
nand U506 (N_506,N_48,N_41);
and U507 (N_507,N_127,N_297);
nor U508 (N_508,N_9,N_125);
nand U509 (N_509,N_106,N_397);
xnor U510 (N_510,N_456,N_294);
nand U511 (N_511,N_195,N_254);
nand U512 (N_512,N_103,N_247);
xor U513 (N_513,N_96,N_64);
and U514 (N_514,N_188,N_5);
nor U515 (N_515,N_38,N_226);
or U516 (N_516,N_178,N_269);
or U517 (N_517,N_401,N_265);
and U518 (N_518,N_222,N_486);
or U519 (N_519,N_235,N_392);
nor U520 (N_520,N_354,N_24);
nor U521 (N_521,N_40,N_182);
nand U522 (N_522,N_83,N_145);
and U523 (N_523,N_396,N_57);
nor U524 (N_524,N_60,N_94);
nor U525 (N_525,N_312,N_262);
and U526 (N_526,N_136,N_364);
nor U527 (N_527,N_452,N_453);
or U528 (N_528,N_264,N_8);
and U529 (N_529,N_325,N_149);
and U530 (N_530,N_58,N_37);
or U531 (N_531,N_191,N_316);
and U532 (N_532,N_51,N_147);
nor U533 (N_533,N_437,N_461);
nand U534 (N_534,N_98,N_102);
or U535 (N_535,N_322,N_55);
nor U536 (N_536,N_258,N_187);
nor U537 (N_537,N_223,N_408);
and U538 (N_538,N_221,N_66);
nor U539 (N_539,N_411,N_141);
and U540 (N_540,N_126,N_151);
nor U541 (N_541,N_478,N_311);
or U542 (N_542,N_35,N_403);
and U543 (N_543,N_365,N_215);
and U544 (N_544,N_199,N_14);
or U545 (N_545,N_53,N_450);
or U546 (N_546,N_313,N_20);
nor U547 (N_547,N_467,N_382);
and U548 (N_548,N_162,N_173);
nand U549 (N_549,N_74,N_131);
or U550 (N_550,N_39,N_70);
or U551 (N_551,N_248,N_308);
nand U552 (N_552,N_498,N_216);
nand U553 (N_553,N_306,N_388);
nor U554 (N_554,N_72,N_193);
nor U555 (N_555,N_255,N_204);
or U556 (N_556,N_232,N_110);
or U557 (N_557,N_389,N_261);
or U558 (N_558,N_302,N_319);
nand U559 (N_559,N_307,N_285);
nor U560 (N_560,N_253,N_448);
or U561 (N_561,N_263,N_495);
or U562 (N_562,N_288,N_295);
nand U563 (N_563,N_436,N_157);
or U564 (N_564,N_45,N_293);
and U565 (N_565,N_260,N_433);
and U566 (N_566,N_324,N_97);
and U567 (N_567,N_230,N_240);
nor U568 (N_568,N_59,N_0);
nand U569 (N_569,N_154,N_114);
and U570 (N_570,N_21,N_372);
nor U571 (N_571,N_205,N_400);
nand U572 (N_572,N_395,N_92);
and U573 (N_573,N_421,N_305);
nand U574 (N_574,N_337,N_394);
and U575 (N_575,N_79,N_170);
nor U576 (N_576,N_416,N_138);
and U577 (N_577,N_479,N_251);
nor U578 (N_578,N_237,N_329);
nor U579 (N_579,N_373,N_19);
or U580 (N_580,N_133,N_326);
nor U581 (N_581,N_327,N_213);
or U582 (N_582,N_426,N_161);
and U583 (N_583,N_12,N_298);
nand U584 (N_584,N_160,N_443);
xor U585 (N_585,N_300,N_301);
and U586 (N_586,N_225,N_415);
or U587 (N_587,N_129,N_243);
and U588 (N_588,N_291,N_259);
nor U589 (N_589,N_474,N_431);
nor U590 (N_590,N_367,N_470);
nand U591 (N_591,N_296,N_132);
xnor U592 (N_592,N_3,N_47);
nand U593 (N_593,N_444,N_22);
nor U594 (N_594,N_377,N_124);
nand U595 (N_595,N_116,N_328);
nand U596 (N_596,N_290,N_277);
nand U597 (N_597,N_424,N_158);
or U598 (N_598,N_32,N_391);
nor U599 (N_599,N_88,N_250);
and U600 (N_600,N_239,N_95);
and U601 (N_601,N_219,N_252);
nor U602 (N_602,N_379,N_180);
or U603 (N_603,N_359,N_87);
nor U604 (N_604,N_487,N_30);
and U605 (N_605,N_344,N_150);
xor U606 (N_606,N_466,N_440);
or U607 (N_607,N_460,N_343);
or U608 (N_608,N_435,N_349);
or U609 (N_609,N_50,N_197);
nor U610 (N_610,N_257,N_245);
and U611 (N_611,N_68,N_481);
and U612 (N_612,N_144,N_482);
nand U613 (N_613,N_29,N_211);
nor U614 (N_614,N_476,N_109);
and U615 (N_615,N_380,N_447);
nand U616 (N_616,N_27,N_156);
nand U617 (N_617,N_181,N_99);
and U618 (N_618,N_65,N_338);
or U619 (N_619,N_363,N_341);
and U620 (N_620,N_413,N_140);
or U621 (N_621,N_80,N_267);
nand U622 (N_622,N_34,N_249);
nor U623 (N_623,N_119,N_422);
nand U624 (N_624,N_176,N_280);
nand U625 (N_625,N_292,N_458);
or U626 (N_626,N_228,N_405);
nor U627 (N_627,N_4,N_407);
and U628 (N_628,N_26,N_206);
and U629 (N_629,N_353,N_346);
or U630 (N_630,N_355,N_104);
and U631 (N_631,N_321,N_445);
nand U632 (N_632,N_271,N_128);
and U633 (N_633,N_483,N_78);
nand U634 (N_634,N_77,N_340);
and U635 (N_635,N_121,N_56);
or U636 (N_636,N_153,N_69);
and U637 (N_637,N_381,N_2);
and U638 (N_638,N_275,N_220);
or U639 (N_639,N_494,N_432);
and U640 (N_640,N_44,N_282);
nand U641 (N_641,N_164,N_49);
or U642 (N_642,N_371,N_246);
and U643 (N_643,N_427,N_71);
nor U644 (N_644,N_33,N_1);
nor U645 (N_645,N_320,N_166);
nand U646 (N_646,N_412,N_75);
nand U647 (N_647,N_477,N_455);
nor U648 (N_648,N_142,N_475);
nor U649 (N_649,N_332,N_6);
or U650 (N_650,N_430,N_463);
nor U651 (N_651,N_434,N_208);
nor U652 (N_652,N_386,N_314);
or U653 (N_653,N_376,N_342);
nand U654 (N_654,N_179,N_283);
and U655 (N_655,N_310,N_315);
and U656 (N_656,N_334,N_214);
nand U657 (N_657,N_274,N_42);
and U658 (N_658,N_118,N_152);
and U659 (N_659,N_425,N_428);
nand U660 (N_660,N_471,N_406);
nand U661 (N_661,N_276,N_200);
or U662 (N_662,N_233,N_174);
nand U663 (N_663,N_167,N_10);
or U664 (N_664,N_304,N_61);
or U665 (N_665,N_446,N_414);
nor U666 (N_666,N_496,N_266);
nand U667 (N_667,N_375,N_360);
nor U668 (N_668,N_137,N_89);
or U669 (N_669,N_168,N_201);
nor U670 (N_670,N_336,N_36);
or U671 (N_671,N_62,N_492);
and U672 (N_672,N_279,N_350);
or U673 (N_673,N_177,N_112);
nand U674 (N_674,N_169,N_352);
nor U675 (N_675,N_497,N_438);
or U676 (N_676,N_82,N_244);
and U677 (N_677,N_370,N_419);
nor U678 (N_678,N_93,N_399);
or U679 (N_679,N_361,N_469);
nand U680 (N_680,N_374,N_7);
nand U681 (N_681,N_449,N_123);
nand U682 (N_682,N_194,N_238);
nand U683 (N_683,N_13,N_417);
nand U684 (N_684,N_429,N_272);
nand U685 (N_685,N_287,N_84);
or U686 (N_686,N_184,N_23);
and U687 (N_687,N_54,N_464);
nor U688 (N_688,N_499,N_462);
and U689 (N_689,N_159,N_91);
and U690 (N_690,N_409,N_86);
or U691 (N_691,N_76,N_345);
nand U692 (N_692,N_31,N_351);
nor U693 (N_693,N_333,N_286);
nand U694 (N_694,N_67,N_90);
nor U695 (N_695,N_190,N_242);
nand U696 (N_696,N_270,N_134);
nand U697 (N_697,N_491,N_369);
nor U698 (N_698,N_139,N_485);
nor U699 (N_699,N_348,N_331);
nand U700 (N_700,N_390,N_171);
nor U701 (N_701,N_148,N_209);
nand U702 (N_702,N_339,N_273);
nand U703 (N_703,N_468,N_490);
or U704 (N_704,N_451,N_317);
and U705 (N_705,N_101,N_473);
and U706 (N_706,N_234,N_163);
nand U707 (N_707,N_358,N_454);
or U708 (N_708,N_362,N_439);
or U709 (N_709,N_196,N_398);
and U710 (N_710,N_241,N_175);
nor U711 (N_711,N_393,N_107);
and U712 (N_712,N_335,N_299);
or U713 (N_713,N_227,N_493);
nor U714 (N_714,N_366,N_318);
or U715 (N_715,N_25,N_122);
or U716 (N_716,N_347,N_385);
nor U717 (N_717,N_198,N_410);
and U718 (N_718,N_309,N_420);
nand U719 (N_719,N_85,N_203);
nand U720 (N_720,N_189,N_192);
or U721 (N_721,N_185,N_143);
nand U722 (N_722,N_100,N_130);
nor U723 (N_723,N_73,N_281);
nand U724 (N_724,N_172,N_323);
or U725 (N_725,N_472,N_11);
or U726 (N_726,N_16,N_384);
nand U727 (N_727,N_202,N_480);
nor U728 (N_728,N_256,N_236);
and U729 (N_729,N_63,N_330);
or U730 (N_730,N_43,N_383);
nand U731 (N_731,N_28,N_165);
nand U732 (N_732,N_105,N_81);
nor U733 (N_733,N_229,N_357);
and U734 (N_734,N_113,N_489);
nand U735 (N_735,N_207,N_457);
nor U736 (N_736,N_111,N_224);
or U737 (N_737,N_52,N_284);
nand U738 (N_738,N_183,N_155);
nor U739 (N_739,N_356,N_465);
nand U740 (N_740,N_186,N_18);
and U741 (N_741,N_278,N_404);
xor U742 (N_742,N_210,N_120);
or U743 (N_743,N_368,N_378);
or U744 (N_744,N_108,N_402);
nor U745 (N_745,N_488,N_459);
nand U746 (N_746,N_46,N_268);
nor U747 (N_747,N_17,N_418);
nor U748 (N_748,N_115,N_303);
and U749 (N_749,N_117,N_217);
nand U750 (N_750,N_178,N_387);
nand U751 (N_751,N_58,N_251);
and U752 (N_752,N_72,N_257);
nand U753 (N_753,N_90,N_123);
and U754 (N_754,N_393,N_77);
nand U755 (N_755,N_226,N_451);
or U756 (N_756,N_464,N_98);
nand U757 (N_757,N_160,N_265);
nor U758 (N_758,N_237,N_153);
or U759 (N_759,N_54,N_258);
nand U760 (N_760,N_195,N_347);
or U761 (N_761,N_452,N_94);
or U762 (N_762,N_257,N_492);
nand U763 (N_763,N_205,N_286);
nor U764 (N_764,N_289,N_86);
nor U765 (N_765,N_250,N_269);
and U766 (N_766,N_96,N_30);
nor U767 (N_767,N_486,N_68);
and U768 (N_768,N_367,N_144);
nand U769 (N_769,N_272,N_137);
or U770 (N_770,N_219,N_64);
and U771 (N_771,N_117,N_168);
nand U772 (N_772,N_349,N_38);
nand U773 (N_773,N_63,N_452);
and U774 (N_774,N_105,N_308);
nor U775 (N_775,N_166,N_202);
or U776 (N_776,N_310,N_345);
and U777 (N_777,N_431,N_189);
nor U778 (N_778,N_258,N_373);
xnor U779 (N_779,N_196,N_66);
and U780 (N_780,N_261,N_496);
nand U781 (N_781,N_104,N_248);
nand U782 (N_782,N_371,N_486);
and U783 (N_783,N_307,N_456);
and U784 (N_784,N_320,N_363);
nor U785 (N_785,N_262,N_446);
or U786 (N_786,N_95,N_304);
or U787 (N_787,N_424,N_153);
nor U788 (N_788,N_317,N_263);
nor U789 (N_789,N_14,N_213);
and U790 (N_790,N_437,N_186);
nor U791 (N_791,N_41,N_425);
nor U792 (N_792,N_258,N_136);
nor U793 (N_793,N_322,N_184);
and U794 (N_794,N_471,N_290);
nand U795 (N_795,N_278,N_399);
nand U796 (N_796,N_27,N_471);
and U797 (N_797,N_173,N_255);
or U798 (N_798,N_81,N_179);
nor U799 (N_799,N_329,N_255);
nand U800 (N_800,N_310,N_1);
nand U801 (N_801,N_89,N_81);
nand U802 (N_802,N_254,N_112);
and U803 (N_803,N_182,N_455);
and U804 (N_804,N_183,N_162);
and U805 (N_805,N_243,N_469);
and U806 (N_806,N_470,N_446);
xnor U807 (N_807,N_146,N_141);
nor U808 (N_808,N_366,N_423);
and U809 (N_809,N_465,N_85);
nand U810 (N_810,N_39,N_100);
nand U811 (N_811,N_108,N_489);
or U812 (N_812,N_125,N_162);
nand U813 (N_813,N_40,N_27);
nor U814 (N_814,N_22,N_438);
and U815 (N_815,N_44,N_312);
or U816 (N_816,N_409,N_75);
nand U817 (N_817,N_262,N_46);
and U818 (N_818,N_422,N_374);
or U819 (N_819,N_81,N_489);
or U820 (N_820,N_156,N_183);
or U821 (N_821,N_299,N_455);
and U822 (N_822,N_91,N_212);
or U823 (N_823,N_12,N_90);
nor U824 (N_824,N_239,N_44);
and U825 (N_825,N_453,N_65);
or U826 (N_826,N_29,N_266);
nor U827 (N_827,N_454,N_452);
and U828 (N_828,N_234,N_145);
or U829 (N_829,N_412,N_306);
and U830 (N_830,N_418,N_364);
nand U831 (N_831,N_385,N_354);
nand U832 (N_832,N_163,N_70);
nor U833 (N_833,N_218,N_429);
nand U834 (N_834,N_33,N_173);
nand U835 (N_835,N_175,N_212);
and U836 (N_836,N_340,N_124);
and U837 (N_837,N_255,N_374);
and U838 (N_838,N_209,N_117);
or U839 (N_839,N_309,N_452);
xor U840 (N_840,N_161,N_360);
or U841 (N_841,N_318,N_160);
or U842 (N_842,N_349,N_241);
nand U843 (N_843,N_295,N_199);
nand U844 (N_844,N_377,N_320);
and U845 (N_845,N_261,N_337);
and U846 (N_846,N_492,N_18);
and U847 (N_847,N_296,N_227);
nor U848 (N_848,N_397,N_133);
nand U849 (N_849,N_428,N_293);
and U850 (N_850,N_457,N_64);
and U851 (N_851,N_20,N_152);
nor U852 (N_852,N_279,N_444);
nor U853 (N_853,N_13,N_395);
nor U854 (N_854,N_20,N_361);
nor U855 (N_855,N_286,N_219);
nor U856 (N_856,N_114,N_462);
nand U857 (N_857,N_46,N_118);
nor U858 (N_858,N_295,N_367);
nor U859 (N_859,N_191,N_446);
or U860 (N_860,N_48,N_208);
or U861 (N_861,N_358,N_478);
nor U862 (N_862,N_432,N_405);
nand U863 (N_863,N_166,N_440);
and U864 (N_864,N_474,N_378);
or U865 (N_865,N_182,N_7);
or U866 (N_866,N_488,N_460);
and U867 (N_867,N_321,N_139);
nand U868 (N_868,N_160,N_174);
nand U869 (N_869,N_182,N_410);
nand U870 (N_870,N_149,N_55);
or U871 (N_871,N_468,N_28);
and U872 (N_872,N_22,N_411);
nand U873 (N_873,N_298,N_373);
xor U874 (N_874,N_488,N_110);
or U875 (N_875,N_370,N_286);
nand U876 (N_876,N_86,N_440);
and U877 (N_877,N_88,N_330);
nor U878 (N_878,N_486,N_431);
and U879 (N_879,N_364,N_256);
or U880 (N_880,N_437,N_0);
nand U881 (N_881,N_419,N_235);
nand U882 (N_882,N_313,N_349);
and U883 (N_883,N_200,N_157);
nand U884 (N_884,N_437,N_466);
nand U885 (N_885,N_49,N_131);
and U886 (N_886,N_149,N_392);
and U887 (N_887,N_6,N_222);
nand U888 (N_888,N_37,N_76);
nand U889 (N_889,N_367,N_407);
nor U890 (N_890,N_73,N_150);
and U891 (N_891,N_28,N_475);
and U892 (N_892,N_4,N_335);
nor U893 (N_893,N_319,N_147);
nand U894 (N_894,N_211,N_338);
and U895 (N_895,N_230,N_30);
nand U896 (N_896,N_174,N_325);
nor U897 (N_897,N_196,N_172);
or U898 (N_898,N_96,N_378);
and U899 (N_899,N_302,N_30);
and U900 (N_900,N_236,N_325);
nor U901 (N_901,N_45,N_77);
or U902 (N_902,N_69,N_446);
or U903 (N_903,N_458,N_126);
or U904 (N_904,N_336,N_440);
and U905 (N_905,N_104,N_83);
nor U906 (N_906,N_6,N_204);
and U907 (N_907,N_482,N_207);
or U908 (N_908,N_396,N_265);
nor U909 (N_909,N_321,N_325);
nor U910 (N_910,N_195,N_10);
and U911 (N_911,N_139,N_46);
or U912 (N_912,N_109,N_81);
and U913 (N_913,N_135,N_487);
and U914 (N_914,N_140,N_361);
and U915 (N_915,N_26,N_473);
and U916 (N_916,N_379,N_83);
or U917 (N_917,N_255,N_224);
nor U918 (N_918,N_36,N_158);
or U919 (N_919,N_322,N_278);
or U920 (N_920,N_225,N_432);
and U921 (N_921,N_18,N_232);
or U922 (N_922,N_480,N_120);
nand U923 (N_923,N_213,N_114);
or U924 (N_924,N_206,N_176);
or U925 (N_925,N_435,N_258);
or U926 (N_926,N_470,N_33);
and U927 (N_927,N_361,N_104);
and U928 (N_928,N_207,N_234);
or U929 (N_929,N_162,N_324);
xor U930 (N_930,N_15,N_175);
and U931 (N_931,N_40,N_80);
nand U932 (N_932,N_156,N_206);
xor U933 (N_933,N_129,N_342);
nor U934 (N_934,N_265,N_210);
nand U935 (N_935,N_156,N_324);
nand U936 (N_936,N_25,N_211);
or U937 (N_937,N_108,N_77);
nor U938 (N_938,N_18,N_157);
nand U939 (N_939,N_489,N_478);
nand U940 (N_940,N_179,N_186);
or U941 (N_941,N_333,N_213);
and U942 (N_942,N_405,N_265);
or U943 (N_943,N_39,N_424);
and U944 (N_944,N_370,N_451);
nor U945 (N_945,N_127,N_336);
nor U946 (N_946,N_463,N_331);
or U947 (N_947,N_3,N_354);
nor U948 (N_948,N_200,N_439);
nor U949 (N_949,N_246,N_6);
and U950 (N_950,N_459,N_380);
and U951 (N_951,N_373,N_226);
and U952 (N_952,N_282,N_311);
nor U953 (N_953,N_207,N_432);
nor U954 (N_954,N_340,N_148);
nand U955 (N_955,N_65,N_5);
and U956 (N_956,N_213,N_78);
or U957 (N_957,N_88,N_75);
nor U958 (N_958,N_474,N_21);
nor U959 (N_959,N_412,N_368);
and U960 (N_960,N_92,N_320);
nand U961 (N_961,N_12,N_151);
nor U962 (N_962,N_149,N_25);
and U963 (N_963,N_268,N_391);
nand U964 (N_964,N_401,N_480);
or U965 (N_965,N_436,N_322);
and U966 (N_966,N_109,N_207);
nand U967 (N_967,N_437,N_419);
or U968 (N_968,N_202,N_161);
and U969 (N_969,N_422,N_273);
and U970 (N_970,N_328,N_306);
nand U971 (N_971,N_23,N_387);
or U972 (N_972,N_265,N_245);
or U973 (N_973,N_320,N_468);
and U974 (N_974,N_1,N_79);
nor U975 (N_975,N_473,N_199);
and U976 (N_976,N_418,N_110);
or U977 (N_977,N_356,N_109);
nor U978 (N_978,N_174,N_15);
and U979 (N_979,N_386,N_70);
nand U980 (N_980,N_472,N_363);
nor U981 (N_981,N_17,N_47);
or U982 (N_982,N_173,N_481);
nor U983 (N_983,N_13,N_99);
and U984 (N_984,N_101,N_310);
nor U985 (N_985,N_315,N_40);
nand U986 (N_986,N_40,N_231);
or U987 (N_987,N_413,N_407);
and U988 (N_988,N_30,N_440);
nand U989 (N_989,N_381,N_156);
nor U990 (N_990,N_362,N_80);
or U991 (N_991,N_311,N_81);
or U992 (N_992,N_184,N_56);
nand U993 (N_993,N_462,N_349);
or U994 (N_994,N_435,N_449);
and U995 (N_995,N_304,N_198);
or U996 (N_996,N_62,N_220);
or U997 (N_997,N_239,N_380);
and U998 (N_998,N_469,N_299);
or U999 (N_999,N_137,N_20);
nand U1000 (N_1000,N_866,N_949);
and U1001 (N_1001,N_661,N_794);
nor U1002 (N_1002,N_785,N_565);
and U1003 (N_1003,N_987,N_518);
nand U1004 (N_1004,N_626,N_554);
and U1005 (N_1005,N_510,N_665);
nand U1006 (N_1006,N_913,N_655);
nand U1007 (N_1007,N_622,N_985);
or U1008 (N_1008,N_810,N_783);
xor U1009 (N_1009,N_504,N_855);
nor U1010 (N_1010,N_743,N_780);
nand U1011 (N_1011,N_962,N_784);
or U1012 (N_1012,N_521,N_546);
nand U1013 (N_1013,N_627,N_539);
and U1014 (N_1014,N_587,N_628);
nand U1015 (N_1015,N_758,N_944);
and U1016 (N_1016,N_578,N_672);
nand U1017 (N_1017,N_909,N_968);
nand U1018 (N_1018,N_556,N_673);
or U1019 (N_1019,N_958,N_973);
nor U1020 (N_1020,N_845,N_983);
nor U1021 (N_1021,N_532,N_812);
or U1022 (N_1022,N_571,N_818);
or U1023 (N_1023,N_891,N_955);
nand U1024 (N_1024,N_905,N_572);
xor U1025 (N_1025,N_975,N_756);
nor U1026 (N_1026,N_735,N_937);
nand U1027 (N_1027,N_841,N_514);
nand U1028 (N_1028,N_809,N_746);
nand U1029 (N_1029,N_523,N_739);
nand U1030 (N_1030,N_912,N_524);
or U1031 (N_1031,N_718,N_522);
and U1032 (N_1032,N_804,N_954);
and U1033 (N_1033,N_779,N_641);
or U1034 (N_1034,N_789,N_834);
nor U1035 (N_1035,N_564,N_802);
or U1036 (N_1036,N_507,N_907);
nand U1037 (N_1037,N_536,N_515);
nand U1038 (N_1038,N_617,N_824);
nor U1039 (N_1039,N_755,N_823);
and U1040 (N_1040,N_753,N_679);
nand U1041 (N_1041,N_737,N_611);
nor U1042 (N_1042,N_871,N_730);
nand U1043 (N_1043,N_829,N_977);
and U1044 (N_1044,N_768,N_956);
and U1045 (N_1045,N_693,N_945);
nor U1046 (N_1046,N_652,N_960);
nor U1047 (N_1047,N_636,N_734);
nor U1048 (N_1048,N_867,N_659);
or U1049 (N_1049,N_586,N_632);
or U1050 (N_1050,N_569,N_864);
and U1051 (N_1051,N_748,N_860);
nand U1052 (N_1052,N_742,N_904);
nor U1053 (N_1053,N_926,N_512);
or U1054 (N_1054,N_674,N_639);
nor U1055 (N_1055,N_844,N_588);
nor U1056 (N_1056,N_579,N_581);
or U1057 (N_1057,N_508,N_813);
and U1058 (N_1058,N_751,N_885);
or U1059 (N_1059,N_869,N_682);
and U1060 (N_1060,N_921,N_553);
nor U1061 (N_1061,N_625,N_555);
and U1062 (N_1062,N_593,N_634);
nand U1063 (N_1063,N_965,N_807);
nand U1064 (N_1064,N_772,N_710);
and U1065 (N_1065,N_832,N_961);
nor U1066 (N_1066,N_910,N_600);
and U1067 (N_1067,N_999,N_876);
or U1068 (N_1068,N_924,N_967);
nor U1069 (N_1069,N_919,N_517);
nand U1070 (N_1070,N_687,N_724);
nand U1071 (N_1071,N_964,N_951);
or U1072 (N_1072,N_981,N_570);
and U1073 (N_1073,N_950,N_857);
nand U1074 (N_1074,N_915,N_574);
and U1075 (N_1075,N_979,N_914);
nand U1076 (N_1076,N_997,N_713);
nor U1077 (N_1077,N_584,N_879);
nor U1078 (N_1078,N_615,N_573);
or U1079 (N_1079,N_744,N_712);
nand U1080 (N_1080,N_596,N_676);
and U1081 (N_1081,N_604,N_660);
nand U1082 (N_1082,N_842,N_880);
or U1083 (N_1083,N_666,N_650);
nor U1084 (N_1084,N_959,N_566);
or U1085 (N_1085,N_653,N_745);
and U1086 (N_1086,N_668,N_662);
or U1087 (N_1087,N_685,N_643);
nand U1088 (N_1088,N_736,N_803);
and U1089 (N_1089,N_616,N_614);
or U1090 (N_1090,N_502,N_731);
nor U1091 (N_1091,N_692,N_870);
nor U1092 (N_1092,N_953,N_932);
nor U1093 (N_1093,N_843,N_778);
nand U1094 (N_1094,N_796,N_723);
nand U1095 (N_1095,N_763,N_852);
xnor U1096 (N_1096,N_911,N_873);
nand U1097 (N_1097,N_620,N_878);
and U1098 (N_1098,N_500,N_542);
nor U1099 (N_1099,N_769,N_791);
and U1100 (N_1100,N_766,N_854);
nor U1101 (N_1101,N_837,N_648);
nand U1102 (N_1102,N_929,N_846);
nand U1103 (N_1103,N_605,N_897);
or U1104 (N_1104,N_621,N_908);
nand U1105 (N_1105,N_757,N_941);
or U1106 (N_1106,N_696,N_705);
or U1107 (N_1107,N_557,N_896);
nor U1108 (N_1108,N_995,N_732);
nand U1109 (N_1109,N_820,N_899);
nand U1110 (N_1110,N_645,N_618);
nand U1111 (N_1111,N_826,N_856);
and U1112 (N_1112,N_669,N_568);
nand U1113 (N_1113,N_901,N_816);
nor U1114 (N_1114,N_825,N_702);
or U1115 (N_1115,N_725,N_946);
and U1116 (N_1116,N_551,N_830);
nor U1117 (N_1117,N_699,N_831);
nand U1118 (N_1118,N_863,N_940);
xor U1119 (N_1119,N_704,N_935);
nor U1120 (N_1120,N_683,N_801);
and U1121 (N_1121,N_637,N_582);
nand U1122 (N_1122,N_609,N_827);
or U1123 (N_1123,N_729,N_635);
xor U1124 (N_1124,N_861,N_630);
nor U1125 (N_1125,N_612,N_976);
and U1126 (N_1126,N_503,N_590);
nor U1127 (N_1127,N_752,N_550);
and U1128 (N_1128,N_681,N_580);
and U1129 (N_1129,N_540,N_547);
nor U1130 (N_1130,N_698,N_817);
and U1131 (N_1131,N_606,N_963);
and U1132 (N_1132,N_898,N_654);
and U1133 (N_1133,N_992,N_534);
or U1134 (N_1134,N_675,N_850);
xnor U1135 (N_1135,N_853,N_623);
nand U1136 (N_1136,N_649,N_776);
nand U1137 (N_1137,N_906,N_529);
or U1138 (N_1138,N_799,N_516);
nand U1139 (N_1139,N_717,N_691);
nor U1140 (N_1140,N_567,N_970);
nor U1141 (N_1141,N_619,N_598);
or U1142 (N_1142,N_722,N_957);
xor U1143 (N_1143,N_750,N_942);
or U1144 (N_1144,N_740,N_525);
or U1145 (N_1145,N_986,N_741);
nor U1146 (N_1146,N_893,N_978);
nand U1147 (N_1147,N_998,N_640);
and U1148 (N_1148,N_773,N_931);
nand U1149 (N_1149,N_642,N_782);
and U1150 (N_1150,N_974,N_689);
nor U1151 (N_1151,N_775,N_838);
and U1152 (N_1152,N_545,N_835);
and U1153 (N_1153,N_697,N_815);
nand U1154 (N_1154,N_948,N_651);
and U1155 (N_1155,N_526,N_786);
and U1156 (N_1156,N_916,N_790);
or U1157 (N_1157,N_805,N_996);
and U1158 (N_1158,N_886,N_501);
or U1159 (N_1159,N_530,N_667);
nand U1160 (N_1160,N_747,N_603);
or U1161 (N_1161,N_980,N_519);
and U1162 (N_1162,N_511,N_583);
nand U1163 (N_1163,N_848,N_943);
nand U1164 (N_1164,N_862,N_688);
nand U1165 (N_1165,N_930,N_684);
or U1166 (N_1166,N_882,N_828);
nor U1167 (N_1167,N_658,N_972);
nor U1168 (N_1168,N_520,N_918);
nor U1169 (N_1169,N_865,N_754);
nor U1170 (N_1170,N_677,N_680);
and U1171 (N_1171,N_938,N_700);
nor U1172 (N_1172,N_990,N_900);
nor U1173 (N_1173,N_721,N_624);
nor U1174 (N_1174,N_629,N_589);
or U1175 (N_1175,N_610,N_822);
and U1176 (N_1176,N_984,N_594);
and U1177 (N_1177,N_777,N_585);
nor U1178 (N_1178,N_638,N_788);
or U1179 (N_1179,N_560,N_719);
nand U1180 (N_1180,N_559,N_726);
or U1181 (N_1181,N_894,N_613);
and U1182 (N_1182,N_933,N_969);
or U1183 (N_1183,N_552,N_795);
or U1184 (N_1184,N_607,N_738);
or U1185 (N_1185,N_808,N_608);
nor U1186 (N_1186,N_708,N_877);
or U1187 (N_1187,N_670,N_599);
nand U1188 (N_1188,N_716,N_770);
and U1189 (N_1189,N_715,N_800);
nor U1190 (N_1190,N_849,N_819);
and U1191 (N_1191,N_814,N_994);
nor U1192 (N_1192,N_558,N_883);
nand U1193 (N_1193,N_947,N_934);
or U1194 (N_1194,N_709,N_592);
nor U1195 (N_1195,N_535,N_859);
nor U1196 (N_1196,N_601,N_836);
nand U1197 (N_1197,N_631,N_922);
or U1198 (N_1198,N_760,N_647);
and U1199 (N_1199,N_533,N_821);
and U1200 (N_1200,N_764,N_727);
nand U1201 (N_1201,N_531,N_591);
nand U1202 (N_1202,N_656,N_549);
or U1203 (N_1203,N_695,N_858);
or U1204 (N_1204,N_548,N_527);
and U1205 (N_1205,N_728,N_991);
nor U1206 (N_1206,N_646,N_561);
nor U1207 (N_1207,N_774,N_694);
nand U1208 (N_1208,N_884,N_762);
nand U1209 (N_1209,N_966,N_798);
or U1210 (N_1210,N_644,N_686);
nand U1211 (N_1211,N_633,N_707);
nand U1212 (N_1212,N_887,N_888);
nor U1213 (N_1213,N_847,N_806);
nor U1214 (N_1214,N_671,N_936);
or U1215 (N_1215,N_663,N_917);
nor U1216 (N_1216,N_923,N_982);
nor U1217 (N_1217,N_563,N_509);
and U1218 (N_1218,N_890,N_811);
nor U1219 (N_1219,N_706,N_597);
and U1220 (N_1220,N_749,N_839);
and U1221 (N_1221,N_840,N_927);
xor U1222 (N_1222,N_971,N_577);
nor U1223 (N_1223,N_720,N_664);
nor U1224 (N_1224,N_711,N_562);
nand U1225 (N_1225,N_690,N_781);
or U1226 (N_1226,N_792,N_513);
and U1227 (N_1227,N_889,N_505);
and U1228 (N_1228,N_902,N_928);
and U1229 (N_1229,N_988,N_602);
nand U1230 (N_1230,N_895,N_543);
xnor U1231 (N_1231,N_993,N_733);
and U1232 (N_1232,N_851,N_872);
or U1233 (N_1233,N_833,N_528);
and U1234 (N_1234,N_868,N_506);
nand U1235 (N_1235,N_881,N_892);
or U1236 (N_1236,N_701,N_989);
nand U1237 (N_1237,N_903,N_761);
nor U1238 (N_1238,N_703,N_925);
nand U1239 (N_1239,N_952,N_759);
nor U1240 (N_1240,N_538,N_874);
and U1241 (N_1241,N_771,N_657);
and U1242 (N_1242,N_678,N_595);
and U1243 (N_1243,N_920,N_575);
nor U1244 (N_1244,N_875,N_767);
and U1245 (N_1245,N_787,N_714);
nand U1246 (N_1246,N_793,N_797);
nand U1247 (N_1247,N_537,N_544);
or U1248 (N_1248,N_765,N_939);
nand U1249 (N_1249,N_576,N_541);
nand U1250 (N_1250,N_686,N_784);
nand U1251 (N_1251,N_969,N_862);
and U1252 (N_1252,N_654,N_681);
and U1253 (N_1253,N_545,N_761);
and U1254 (N_1254,N_715,N_891);
nor U1255 (N_1255,N_808,N_859);
nor U1256 (N_1256,N_791,N_703);
and U1257 (N_1257,N_645,N_934);
nand U1258 (N_1258,N_635,N_823);
nand U1259 (N_1259,N_841,N_778);
nor U1260 (N_1260,N_945,N_780);
or U1261 (N_1261,N_998,N_670);
and U1262 (N_1262,N_877,N_546);
nand U1263 (N_1263,N_936,N_818);
nor U1264 (N_1264,N_639,N_974);
and U1265 (N_1265,N_891,N_509);
nand U1266 (N_1266,N_731,N_670);
and U1267 (N_1267,N_904,N_686);
or U1268 (N_1268,N_648,N_647);
or U1269 (N_1269,N_701,N_744);
or U1270 (N_1270,N_818,N_839);
nand U1271 (N_1271,N_949,N_712);
nand U1272 (N_1272,N_700,N_576);
and U1273 (N_1273,N_564,N_842);
nand U1274 (N_1274,N_890,N_981);
nand U1275 (N_1275,N_533,N_616);
nand U1276 (N_1276,N_695,N_924);
or U1277 (N_1277,N_956,N_979);
nor U1278 (N_1278,N_905,N_734);
nand U1279 (N_1279,N_850,N_721);
and U1280 (N_1280,N_786,N_693);
nand U1281 (N_1281,N_586,N_504);
and U1282 (N_1282,N_912,N_601);
and U1283 (N_1283,N_662,N_681);
or U1284 (N_1284,N_544,N_605);
and U1285 (N_1285,N_821,N_914);
nor U1286 (N_1286,N_908,N_724);
nand U1287 (N_1287,N_668,N_641);
or U1288 (N_1288,N_575,N_931);
nor U1289 (N_1289,N_970,N_664);
nor U1290 (N_1290,N_973,N_795);
nand U1291 (N_1291,N_887,N_940);
and U1292 (N_1292,N_947,N_860);
and U1293 (N_1293,N_978,N_879);
nand U1294 (N_1294,N_524,N_677);
nand U1295 (N_1295,N_968,N_845);
nand U1296 (N_1296,N_520,N_956);
and U1297 (N_1297,N_997,N_879);
or U1298 (N_1298,N_825,N_996);
or U1299 (N_1299,N_862,N_507);
nor U1300 (N_1300,N_697,N_999);
nor U1301 (N_1301,N_890,N_950);
or U1302 (N_1302,N_611,N_932);
nor U1303 (N_1303,N_615,N_545);
nor U1304 (N_1304,N_728,N_961);
nand U1305 (N_1305,N_929,N_925);
and U1306 (N_1306,N_516,N_976);
xnor U1307 (N_1307,N_653,N_840);
or U1308 (N_1308,N_688,N_769);
nor U1309 (N_1309,N_696,N_539);
or U1310 (N_1310,N_511,N_903);
nor U1311 (N_1311,N_741,N_805);
and U1312 (N_1312,N_797,N_858);
nor U1313 (N_1313,N_829,N_504);
nor U1314 (N_1314,N_592,N_938);
nand U1315 (N_1315,N_633,N_911);
xor U1316 (N_1316,N_622,N_858);
nand U1317 (N_1317,N_882,N_696);
and U1318 (N_1318,N_749,N_657);
nor U1319 (N_1319,N_797,N_905);
and U1320 (N_1320,N_875,N_811);
or U1321 (N_1321,N_915,N_898);
nand U1322 (N_1322,N_968,N_599);
nor U1323 (N_1323,N_536,N_862);
nand U1324 (N_1324,N_557,N_797);
nor U1325 (N_1325,N_862,N_876);
nor U1326 (N_1326,N_680,N_853);
nor U1327 (N_1327,N_814,N_787);
nor U1328 (N_1328,N_824,N_557);
and U1329 (N_1329,N_861,N_939);
or U1330 (N_1330,N_992,N_640);
or U1331 (N_1331,N_508,N_659);
and U1332 (N_1332,N_537,N_753);
nand U1333 (N_1333,N_815,N_662);
and U1334 (N_1334,N_574,N_513);
and U1335 (N_1335,N_692,N_959);
nor U1336 (N_1336,N_720,N_825);
nand U1337 (N_1337,N_851,N_585);
and U1338 (N_1338,N_518,N_810);
or U1339 (N_1339,N_654,N_976);
nor U1340 (N_1340,N_919,N_868);
nor U1341 (N_1341,N_812,N_669);
and U1342 (N_1342,N_538,N_911);
and U1343 (N_1343,N_870,N_964);
nor U1344 (N_1344,N_531,N_654);
or U1345 (N_1345,N_992,N_610);
xnor U1346 (N_1346,N_524,N_639);
or U1347 (N_1347,N_979,N_988);
or U1348 (N_1348,N_600,N_665);
and U1349 (N_1349,N_593,N_878);
or U1350 (N_1350,N_538,N_765);
nor U1351 (N_1351,N_767,N_822);
or U1352 (N_1352,N_533,N_846);
nand U1353 (N_1353,N_983,N_851);
nand U1354 (N_1354,N_982,N_764);
nand U1355 (N_1355,N_530,N_632);
nand U1356 (N_1356,N_827,N_682);
and U1357 (N_1357,N_777,N_960);
nand U1358 (N_1358,N_610,N_737);
or U1359 (N_1359,N_874,N_750);
and U1360 (N_1360,N_669,N_838);
or U1361 (N_1361,N_848,N_526);
or U1362 (N_1362,N_998,N_972);
nand U1363 (N_1363,N_641,N_541);
nand U1364 (N_1364,N_861,N_587);
and U1365 (N_1365,N_827,N_551);
nand U1366 (N_1366,N_950,N_989);
nand U1367 (N_1367,N_732,N_849);
and U1368 (N_1368,N_540,N_800);
nand U1369 (N_1369,N_926,N_622);
and U1370 (N_1370,N_650,N_604);
or U1371 (N_1371,N_693,N_940);
or U1372 (N_1372,N_679,N_892);
or U1373 (N_1373,N_812,N_717);
or U1374 (N_1374,N_875,N_850);
or U1375 (N_1375,N_516,N_519);
nor U1376 (N_1376,N_634,N_954);
and U1377 (N_1377,N_816,N_797);
nand U1378 (N_1378,N_740,N_778);
and U1379 (N_1379,N_948,N_652);
nand U1380 (N_1380,N_785,N_855);
or U1381 (N_1381,N_795,N_856);
and U1382 (N_1382,N_979,N_503);
nor U1383 (N_1383,N_783,N_866);
or U1384 (N_1384,N_806,N_804);
or U1385 (N_1385,N_713,N_529);
nand U1386 (N_1386,N_979,N_933);
nor U1387 (N_1387,N_783,N_791);
nor U1388 (N_1388,N_828,N_878);
and U1389 (N_1389,N_552,N_593);
or U1390 (N_1390,N_893,N_977);
and U1391 (N_1391,N_769,N_929);
nand U1392 (N_1392,N_612,N_868);
nand U1393 (N_1393,N_733,N_723);
and U1394 (N_1394,N_743,N_575);
and U1395 (N_1395,N_761,N_962);
and U1396 (N_1396,N_973,N_612);
nor U1397 (N_1397,N_779,N_856);
or U1398 (N_1398,N_722,N_527);
nand U1399 (N_1399,N_640,N_755);
nand U1400 (N_1400,N_668,N_643);
nor U1401 (N_1401,N_955,N_686);
nor U1402 (N_1402,N_785,N_737);
and U1403 (N_1403,N_809,N_740);
or U1404 (N_1404,N_546,N_857);
nand U1405 (N_1405,N_544,N_500);
nand U1406 (N_1406,N_632,N_995);
nor U1407 (N_1407,N_953,N_669);
and U1408 (N_1408,N_705,N_868);
nor U1409 (N_1409,N_782,N_676);
nand U1410 (N_1410,N_693,N_670);
and U1411 (N_1411,N_743,N_729);
xnor U1412 (N_1412,N_539,N_709);
and U1413 (N_1413,N_784,N_715);
or U1414 (N_1414,N_839,N_978);
and U1415 (N_1415,N_985,N_686);
nor U1416 (N_1416,N_905,N_643);
or U1417 (N_1417,N_811,N_796);
nand U1418 (N_1418,N_949,N_736);
and U1419 (N_1419,N_530,N_935);
or U1420 (N_1420,N_711,N_623);
nor U1421 (N_1421,N_562,N_702);
nand U1422 (N_1422,N_948,N_591);
nand U1423 (N_1423,N_764,N_530);
nor U1424 (N_1424,N_829,N_605);
and U1425 (N_1425,N_508,N_791);
and U1426 (N_1426,N_837,N_649);
and U1427 (N_1427,N_823,N_627);
nand U1428 (N_1428,N_979,N_972);
nor U1429 (N_1429,N_968,N_591);
and U1430 (N_1430,N_990,N_547);
nand U1431 (N_1431,N_870,N_803);
and U1432 (N_1432,N_678,N_518);
nand U1433 (N_1433,N_886,N_644);
nor U1434 (N_1434,N_861,N_829);
nand U1435 (N_1435,N_938,N_559);
nor U1436 (N_1436,N_606,N_924);
nor U1437 (N_1437,N_982,N_797);
nor U1438 (N_1438,N_616,N_915);
or U1439 (N_1439,N_995,N_547);
xnor U1440 (N_1440,N_508,N_752);
and U1441 (N_1441,N_620,N_917);
nor U1442 (N_1442,N_919,N_999);
or U1443 (N_1443,N_683,N_995);
nor U1444 (N_1444,N_931,N_776);
nand U1445 (N_1445,N_888,N_966);
and U1446 (N_1446,N_694,N_726);
and U1447 (N_1447,N_808,N_556);
nand U1448 (N_1448,N_593,N_528);
or U1449 (N_1449,N_534,N_549);
or U1450 (N_1450,N_700,N_744);
or U1451 (N_1451,N_877,N_645);
and U1452 (N_1452,N_706,N_910);
and U1453 (N_1453,N_508,N_622);
or U1454 (N_1454,N_837,N_748);
or U1455 (N_1455,N_874,N_577);
nand U1456 (N_1456,N_639,N_867);
or U1457 (N_1457,N_691,N_863);
or U1458 (N_1458,N_982,N_581);
nor U1459 (N_1459,N_993,N_681);
or U1460 (N_1460,N_938,N_652);
nand U1461 (N_1461,N_913,N_528);
nand U1462 (N_1462,N_912,N_572);
nor U1463 (N_1463,N_517,N_959);
and U1464 (N_1464,N_790,N_697);
and U1465 (N_1465,N_852,N_955);
and U1466 (N_1466,N_727,N_883);
or U1467 (N_1467,N_671,N_757);
or U1468 (N_1468,N_531,N_637);
nor U1469 (N_1469,N_592,N_743);
and U1470 (N_1470,N_781,N_803);
and U1471 (N_1471,N_923,N_555);
or U1472 (N_1472,N_661,N_554);
nand U1473 (N_1473,N_684,N_766);
xnor U1474 (N_1474,N_943,N_685);
nand U1475 (N_1475,N_558,N_596);
nand U1476 (N_1476,N_771,N_680);
nand U1477 (N_1477,N_715,N_580);
or U1478 (N_1478,N_860,N_725);
xnor U1479 (N_1479,N_792,N_834);
nor U1480 (N_1480,N_905,N_891);
nand U1481 (N_1481,N_827,N_886);
or U1482 (N_1482,N_546,N_964);
nor U1483 (N_1483,N_974,N_622);
nor U1484 (N_1484,N_929,N_767);
xor U1485 (N_1485,N_559,N_557);
nor U1486 (N_1486,N_921,N_616);
or U1487 (N_1487,N_824,N_508);
and U1488 (N_1488,N_955,N_788);
nor U1489 (N_1489,N_799,N_684);
or U1490 (N_1490,N_600,N_662);
nand U1491 (N_1491,N_542,N_681);
or U1492 (N_1492,N_735,N_726);
xnor U1493 (N_1493,N_642,N_608);
nor U1494 (N_1494,N_931,N_661);
and U1495 (N_1495,N_600,N_979);
nor U1496 (N_1496,N_645,N_518);
nor U1497 (N_1497,N_875,N_652);
and U1498 (N_1498,N_800,N_947);
nand U1499 (N_1499,N_951,N_563);
and U1500 (N_1500,N_1426,N_1489);
and U1501 (N_1501,N_1384,N_1457);
and U1502 (N_1502,N_1174,N_1068);
and U1503 (N_1503,N_1157,N_1230);
nand U1504 (N_1504,N_1317,N_1051);
nor U1505 (N_1505,N_1013,N_1178);
or U1506 (N_1506,N_1477,N_1413);
nor U1507 (N_1507,N_1282,N_1213);
nand U1508 (N_1508,N_1333,N_1259);
nor U1509 (N_1509,N_1168,N_1304);
nand U1510 (N_1510,N_1476,N_1309);
or U1511 (N_1511,N_1375,N_1197);
nor U1512 (N_1512,N_1224,N_1034);
or U1513 (N_1513,N_1411,N_1049);
and U1514 (N_1514,N_1179,N_1371);
nand U1515 (N_1515,N_1402,N_1467);
or U1516 (N_1516,N_1439,N_1172);
and U1517 (N_1517,N_1189,N_1126);
or U1518 (N_1518,N_1058,N_1221);
and U1519 (N_1519,N_1407,N_1163);
nor U1520 (N_1520,N_1326,N_1130);
and U1521 (N_1521,N_1369,N_1095);
or U1522 (N_1522,N_1039,N_1316);
xnor U1523 (N_1523,N_1430,N_1212);
and U1524 (N_1524,N_1387,N_1208);
or U1525 (N_1525,N_1123,N_1142);
or U1526 (N_1526,N_1194,N_1285);
and U1527 (N_1527,N_1358,N_1061);
nor U1528 (N_1528,N_1480,N_1493);
nand U1529 (N_1529,N_1398,N_1075);
nand U1530 (N_1530,N_1349,N_1004);
or U1531 (N_1531,N_1283,N_1040);
and U1532 (N_1532,N_1138,N_1287);
nor U1533 (N_1533,N_1483,N_1492);
nand U1534 (N_1534,N_1159,N_1237);
nand U1535 (N_1535,N_1217,N_1320);
and U1536 (N_1536,N_1300,N_1268);
and U1537 (N_1537,N_1451,N_1105);
xnor U1538 (N_1538,N_1408,N_1462);
or U1539 (N_1539,N_1487,N_1052);
and U1540 (N_1540,N_1472,N_1114);
nor U1541 (N_1541,N_1288,N_1404);
and U1542 (N_1542,N_1137,N_1222);
nor U1543 (N_1543,N_1148,N_1295);
and U1544 (N_1544,N_1290,N_1002);
and U1545 (N_1545,N_1279,N_1323);
nand U1546 (N_1546,N_1044,N_1458);
nand U1547 (N_1547,N_1030,N_1464);
nand U1548 (N_1548,N_1352,N_1147);
and U1549 (N_1549,N_1399,N_1080);
or U1550 (N_1550,N_1264,N_1141);
nor U1551 (N_1551,N_1233,N_1028);
nor U1552 (N_1552,N_1247,N_1165);
and U1553 (N_1553,N_1225,N_1019);
or U1554 (N_1554,N_1433,N_1261);
nand U1555 (N_1555,N_1188,N_1447);
or U1556 (N_1556,N_1468,N_1424);
or U1557 (N_1557,N_1365,N_1348);
nand U1558 (N_1558,N_1175,N_1059);
xnor U1559 (N_1559,N_1111,N_1435);
and U1560 (N_1560,N_1297,N_1110);
nor U1561 (N_1561,N_1298,N_1332);
nand U1562 (N_1562,N_1379,N_1104);
or U1563 (N_1563,N_1215,N_1236);
nand U1564 (N_1564,N_1354,N_1335);
nor U1565 (N_1565,N_1334,N_1460);
or U1566 (N_1566,N_1419,N_1270);
nand U1567 (N_1567,N_1183,N_1299);
nor U1568 (N_1568,N_1312,N_1228);
or U1569 (N_1569,N_1377,N_1339);
or U1570 (N_1570,N_1146,N_1275);
or U1571 (N_1571,N_1362,N_1205);
and U1572 (N_1572,N_1015,N_1229);
and U1573 (N_1573,N_1461,N_1310);
nand U1574 (N_1574,N_1380,N_1429);
and U1575 (N_1575,N_1181,N_1344);
nor U1576 (N_1576,N_1294,N_1246);
or U1577 (N_1577,N_1200,N_1001);
nand U1578 (N_1578,N_1448,N_1242);
and U1579 (N_1579,N_1106,N_1390);
or U1580 (N_1580,N_1265,N_1441);
and U1581 (N_1581,N_1227,N_1238);
and U1582 (N_1582,N_1470,N_1177);
xnor U1583 (N_1583,N_1330,N_1289);
and U1584 (N_1584,N_1158,N_1026);
or U1585 (N_1585,N_1145,N_1386);
and U1586 (N_1586,N_1496,N_1083);
or U1587 (N_1587,N_1118,N_1047);
and U1588 (N_1588,N_1108,N_1251);
and U1589 (N_1589,N_1066,N_1060);
nor U1590 (N_1590,N_1240,N_1274);
nor U1591 (N_1591,N_1396,N_1056);
and U1592 (N_1592,N_1409,N_1069);
or U1593 (N_1593,N_1166,N_1219);
nand U1594 (N_1594,N_1389,N_1042);
nand U1595 (N_1595,N_1169,N_1154);
and U1596 (N_1596,N_1113,N_1440);
or U1597 (N_1597,N_1452,N_1363);
nand U1598 (N_1598,N_1436,N_1206);
nand U1599 (N_1599,N_1167,N_1432);
nand U1600 (N_1600,N_1007,N_1134);
nor U1601 (N_1601,N_1370,N_1100);
or U1602 (N_1602,N_1173,N_1164);
nor U1603 (N_1603,N_1491,N_1347);
nor U1604 (N_1604,N_1361,N_1416);
or U1605 (N_1605,N_1373,N_1437);
nor U1606 (N_1606,N_1277,N_1161);
or U1607 (N_1607,N_1280,N_1003);
nand U1608 (N_1608,N_1293,N_1239);
nand U1609 (N_1609,N_1121,N_1021);
nand U1610 (N_1610,N_1022,N_1186);
nor U1611 (N_1611,N_1490,N_1223);
nand U1612 (N_1612,N_1431,N_1421);
nor U1613 (N_1613,N_1356,N_1382);
nor U1614 (N_1614,N_1043,N_1091);
nand U1615 (N_1615,N_1392,N_1292);
nand U1616 (N_1616,N_1434,N_1391);
and U1617 (N_1617,N_1184,N_1325);
nand U1618 (N_1618,N_1263,N_1176);
nand U1619 (N_1619,N_1036,N_1202);
nand U1620 (N_1620,N_1449,N_1406);
or U1621 (N_1621,N_1256,N_1281);
nand U1622 (N_1622,N_1235,N_1395);
nor U1623 (N_1623,N_1008,N_1269);
and U1624 (N_1624,N_1364,N_1135);
xor U1625 (N_1625,N_1378,N_1357);
nor U1626 (N_1626,N_1079,N_1014);
or U1627 (N_1627,N_1445,N_1185);
or U1628 (N_1628,N_1000,N_1057);
nor U1629 (N_1629,N_1403,N_1331);
and U1630 (N_1630,N_1025,N_1053);
and U1631 (N_1631,N_1074,N_1423);
nand U1632 (N_1632,N_1063,N_1248);
nor U1633 (N_1633,N_1016,N_1474);
or U1634 (N_1634,N_1397,N_1345);
nand U1635 (N_1635,N_1143,N_1249);
xnor U1636 (N_1636,N_1351,N_1427);
and U1637 (N_1637,N_1045,N_1258);
and U1638 (N_1638,N_1254,N_1005);
xor U1639 (N_1639,N_1307,N_1267);
nor U1640 (N_1640,N_1355,N_1243);
and U1641 (N_1641,N_1198,N_1338);
nand U1642 (N_1642,N_1149,N_1082);
and U1643 (N_1643,N_1071,N_1131);
nor U1644 (N_1644,N_1006,N_1302);
nand U1645 (N_1645,N_1191,N_1284);
and U1646 (N_1646,N_1400,N_1327);
and U1647 (N_1647,N_1203,N_1276);
xnor U1648 (N_1648,N_1350,N_1089);
and U1649 (N_1649,N_1035,N_1466);
or U1650 (N_1650,N_1128,N_1315);
and U1651 (N_1651,N_1401,N_1313);
or U1652 (N_1652,N_1086,N_1046);
nand U1653 (N_1653,N_1182,N_1278);
nor U1654 (N_1654,N_1011,N_1455);
or U1655 (N_1655,N_1368,N_1346);
nand U1656 (N_1656,N_1475,N_1125);
or U1657 (N_1657,N_1062,N_1340);
nor U1658 (N_1658,N_1226,N_1443);
nor U1659 (N_1659,N_1498,N_1214);
nor U1660 (N_1660,N_1210,N_1442);
xnor U1661 (N_1661,N_1107,N_1101);
nand U1662 (N_1662,N_1065,N_1418);
and U1663 (N_1663,N_1207,N_1160);
nand U1664 (N_1664,N_1324,N_1497);
nor U1665 (N_1665,N_1253,N_1054);
or U1666 (N_1666,N_1076,N_1092);
nand U1667 (N_1667,N_1412,N_1456);
nand U1668 (N_1668,N_1372,N_1087);
xnor U1669 (N_1669,N_1038,N_1020);
and U1670 (N_1670,N_1446,N_1425);
xnor U1671 (N_1671,N_1311,N_1393);
and U1672 (N_1672,N_1232,N_1381);
or U1673 (N_1673,N_1192,N_1009);
nand U1674 (N_1674,N_1438,N_1454);
or U1675 (N_1675,N_1322,N_1070);
nand U1676 (N_1676,N_1231,N_1018);
nand U1677 (N_1677,N_1360,N_1140);
and U1678 (N_1678,N_1041,N_1394);
or U1679 (N_1679,N_1081,N_1099);
or U1680 (N_1680,N_1195,N_1252);
or U1681 (N_1681,N_1272,N_1048);
or U1682 (N_1682,N_1271,N_1144);
nand U1683 (N_1683,N_1090,N_1343);
and U1684 (N_1684,N_1193,N_1450);
and U1685 (N_1685,N_1266,N_1305);
nand U1686 (N_1686,N_1033,N_1120);
xor U1687 (N_1687,N_1481,N_1417);
and U1688 (N_1688,N_1170,N_1273);
or U1689 (N_1689,N_1129,N_1257);
or U1690 (N_1690,N_1024,N_1245);
nor U1691 (N_1691,N_1414,N_1353);
nand U1692 (N_1692,N_1415,N_1112);
or U1693 (N_1693,N_1337,N_1136);
nor U1694 (N_1694,N_1196,N_1156);
nor U1695 (N_1695,N_1064,N_1255);
nor U1696 (N_1696,N_1469,N_1211);
and U1697 (N_1697,N_1096,N_1201);
nor U1698 (N_1698,N_1488,N_1209);
or U1699 (N_1699,N_1204,N_1301);
nand U1700 (N_1700,N_1132,N_1055);
nand U1701 (N_1701,N_1341,N_1485);
or U1702 (N_1702,N_1139,N_1484);
nor U1703 (N_1703,N_1218,N_1102);
or U1704 (N_1704,N_1422,N_1097);
and U1705 (N_1705,N_1084,N_1029);
nand U1706 (N_1706,N_1494,N_1151);
and U1707 (N_1707,N_1199,N_1094);
or U1708 (N_1708,N_1319,N_1077);
and U1709 (N_1709,N_1085,N_1336);
or U1710 (N_1710,N_1495,N_1329);
nand U1711 (N_1711,N_1383,N_1190);
or U1712 (N_1712,N_1473,N_1321);
nor U1713 (N_1713,N_1410,N_1152);
and U1714 (N_1714,N_1465,N_1119);
nor U1715 (N_1715,N_1367,N_1187);
nor U1716 (N_1716,N_1482,N_1155);
nor U1717 (N_1717,N_1250,N_1328);
nand U1718 (N_1718,N_1098,N_1303);
and U1719 (N_1719,N_1359,N_1260);
nor U1720 (N_1720,N_1216,N_1117);
or U1721 (N_1721,N_1023,N_1318);
and U1722 (N_1722,N_1220,N_1162);
nor U1723 (N_1723,N_1241,N_1479);
nor U1724 (N_1724,N_1286,N_1116);
nor U1725 (N_1725,N_1133,N_1153);
or U1726 (N_1726,N_1122,N_1073);
and U1727 (N_1727,N_1027,N_1499);
nand U1728 (N_1728,N_1374,N_1031);
and U1729 (N_1729,N_1067,N_1308);
nand U1730 (N_1730,N_1420,N_1037);
nor U1731 (N_1731,N_1314,N_1017);
or U1732 (N_1732,N_1471,N_1050);
nand U1733 (N_1733,N_1388,N_1078);
and U1734 (N_1734,N_1124,N_1459);
or U1735 (N_1735,N_1180,N_1103);
nor U1736 (N_1736,N_1150,N_1453);
nand U1737 (N_1737,N_1486,N_1342);
and U1738 (N_1738,N_1010,N_1428);
nor U1739 (N_1739,N_1115,N_1262);
nand U1740 (N_1740,N_1244,N_1012);
nand U1741 (N_1741,N_1171,N_1093);
and U1742 (N_1742,N_1032,N_1366);
xor U1743 (N_1743,N_1088,N_1072);
nor U1744 (N_1744,N_1478,N_1234);
and U1745 (N_1745,N_1306,N_1127);
and U1746 (N_1746,N_1463,N_1109);
or U1747 (N_1747,N_1291,N_1385);
and U1748 (N_1748,N_1444,N_1405);
or U1749 (N_1749,N_1296,N_1376);
nand U1750 (N_1750,N_1348,N_1473);
nand U1751 (N_1751,N_1483,N_1362);
nand U1752 (N_1752,N_1171,N_1278);
nor U1753 (N_1753,N_1499,N_1258);
nand U1754 (N_1754,N_1255,N_1099);
or U1755 (N_1755,N_1123,N_1445);
and U1756 (N_1756,N_1342,N_1480);
nand U1757 (N_1757,N_1282,N_1359);
or U1758 (N_1758,N_1291,N_1142);
nand U1759 (N_1759,N_1039,N_1334);
nand U1760 (N_1760,N_1189,N_1014);
nand U1761 (N_1761,N_1033,N_1126);
or U1762 (N_1762,N_1049,N_1368);
or U1763 (N_1763,N_1332,N_1342);
or U1764 (N_1764,N_1030,N_1027);
or U1765 (N_1765,N_1223,N_1374);
nand U1766 (N_1766,N_1050,N_1375);
or U1767 (N_1767,N_1074,N_1270);
and U1768 (N_1768,N_1207,N_1428);
or U1769 (N_1769,N_1483,N_1323);
or U1770 (N_1770,N_1228,N_1293);
and U1771 (N_1771,N_1320,N_1372);
and U1772 (N_1772,N_1393,N_1096);
or U1773 (N_1773,N_1290,N_1148);
and U1774 (N_1774,N_1499,N_1289);
and U1775 (N_1775,N_1106,N_1314);
nand U1776 (N_1776,N_1281,N_1345);
nor U1777 (N_1777,N_1250,N_1396);
or U1778 (N_1778,N_1490,N_1241);
or U1779 (N_1779,N_1229,N_1230);
nand U1780 (N_1780,N_1130,N_1304);
and U1781 (N_1781,N_1130,N_1270);
or U1782 (N_1782,N_1177,N_1208);
and U1783 (N_1783,N_1382,N_1067);
and U1784 (N_1784,N_1195,N_1415);
nor U1785 (N_1785,N_1311,N_1392);
and U1786 (N_1786,N_1318,N_1410);
or U1787 (N_1787,N_1089,N_1372);
or U1788 (N_1788,N_1480,N_1436);
nor U1789 (N_1789,N_1297,N_1176);
and U1790 (N_1790,N_1358,N_1196);
nor U1791 (N_1791,N_1100,N_1163);
and U1792 (N_1792,N_1062,N_1129);
nor U1793 (N_1793,N_1409,N_1036);
and U1794 (N_1794,N_1315,N_1068);
nand U1795 (N_1795,N_1416,N_1237);
nor U1796 (N_1796,N_1238,N_1092);
xor U1797 (N_1797,N_1193,N_1290);
nor U1798 (N_1798,N_1173,N_1149);
nand U1799 (N_1799,N_1179,N_1497);
nor U1800 (N_1800,N_1425,N_1131);
and U1801 (N_1801,N_1028,N_1224);
nand U1802 (N_1802,N_1030,N_1374);
or U1803 (N_1803,N_1217,N_1103);
or U1804 (N_1804,N_1122,N_1305);
nand U1805 (N_1805,N_1292,N_1012);
nor U1806 (N_1806,N_1432,N_1300);
nand U1807 (N_1807,N_1168,N_1197);
and U1808 (N_1808,N_1028,N_1240);
and U1809 (N_1809,N_1059,N_1371);
or U1810 (N_1810,N_1021,N_1135);
xnor U1811 (N_1811,N_1451,N_1103);
nand U1812 (N_1812,N_1402,N_1479);
nand U1813 (N_1813,N_1298,N_1020);
or U1814 (N_1814,N_1232,N_1324);
nand U1815 (N_1815,N_1240,N_1166);
nand U1816 (N_1816,N_1179,N_1105);
or U1817 (N_1817,N_1048,N_1416);
nor U1818 (N_1818,N_1198,N_1219);
nor U1819 (N_1819,N_1217,N_1167);
and U1820 (N_1820,N_1356,N_1010);
xnor U1821 (N_1821,N_1224,N_1111);
or U1822 (N_1822,N_1407,N_1289);
or U1823 (N_1823,N_1187,N_1236);
nor U1824 (N_1824,N_1375,N_1043);
nor U1825 (N_1825,N_1344,N_1247);
nand U1826 (N_1826,N_1264,N_1473);
or U1827 (N_1827,N_1097,N_1155);
nand U1828 (N_1828,N_1401,N_1365);
nand U1829 (N_1829,N_1135,N_1262);
nor U1830 (N_1830,N_1206,N_1089);
nand U1831 (N_1831,N_1005,N_1364);
and U1832 (N_1832,N_1105,N_1284);
nand U1833 (N_1833,N_1163,N_1210);
and U1834 (N_1834,N_1336,N_1304);
and U1835 (N_1835,N_1052,N_1455);
nor U1836 (N_1836,N_1251,N_1293);
or U1837 (N_1837,N_1427,N_1266);
or U1838 (N_1838,N_1426,N_1187);
nand U1839 (N_1839,N_1486,N_1019);
and U1840 (N_1840,N_1137,N_1327);
nand U1841 (N_1841,N_1453,N_1003);
or U1842 (N_1842,N_1334,N_1187);
xor U1843 (N_1843,N_1205,N_1443);
nand U1844 (N_1844,N_1410,N_1086);
nand U1845 (N_1845,N_1436,N_1074);
nand U1846 (N_1846,N_1004,N_1353);
nor U1847 (N_1847,N_1310,N_1223);
or U1848 (N_1848,N_1229,N_1214);
and U1849 (N_1849,N_1402,N_1302);
or U1850 (N_1850,N_1169,N_1407);
and U1851 (N_1851,N_1376,N_1337);
nor U1852 (N_1852,N_1203,N_1342);
nand U1853 (N_1853,N_1019,N_1099);
or U1854 (N_1854,N_1084,N_1461);
and U1855 (N_1855,N_1371,N_1082);
or U1856 (N_1856,N_1322,N_1369);
nand U1857 (N_1857,N_1032,N_1372);
or U1858 (N_1858,N_1012,N_1067);
and U1859 (N_1859,N_1268,N_1153);
and U1860 (N_1860,N_1379,N_1393);
nand U1861 (N_1861,N_1035,N_1359);
nor U1862 (N_1862,N_1117,N_1185);
nand U1863 (N_1863,N_1225,N_1490);
and U1864 (N_1864,N_1149,N_1268);
nor U1865 (N_1865,N_1359,N_1425);
nor U1866 (N_1866,N_1428,N_1445);
and U1867 (N_1867,N_1439,N_1428);
or U1868 (N_1868,N_1280,N_1169);
nor U1869 (N_1869,N_1428,N_1212);
and U1870 (N_1870,N_1414,N_1261);
and U1871 (N_1871,N_1180,N_1184);
or U1872 (N_1872,N_1323,N_1086);
nor U1873 (N_1873,N_1073,N_1166);
nor U1874 (N_1874,N_1422,N_1024);
and U1875 (N_1875,N_1423,N_1063);
xor U1876 (N_1876,N_1005,N_1183);
nand U1877 (N_1877,N_1349,N_1289);
or U1878 (N_1878,N_1209,N_1087);
and U1879 (N_1879,N_1085,N_1322);
nand U1880 (N_1880,N_1407,N_1193);
and U1881 (N_1881,N_1491,N_1120);
nor U1882 (N_1882,N_1491,N_1485);
or U1883 (N_1883,N_1133,N_1408);
or U1884 (N_1884,N_1313,N_1193);
nor U1885 (N_1885,N_1444,N_1200);
and U1886 (N_1886,N_1448,N_1354);
or U1887 (N_1887,N_1213,N_1155);
or U1888 (N_1888,N_1190,N_1307);
xor U1889 (N_1889,N_1388,N_1387);
nand U1890 (N_1890,N_1480,N_1010);
or U1891 (N_1891,N_1499,N_1297);
nand U1892 (N_1892,N_1204,N_1167);
or U1893 (N_1893,N_1241,N_1085);
nand U1894 (N_1894,N_1423,N_1320);
or U1895 (N_1895,N_1227,N_1218);
nor U1896 (N_1896,N_1123,N_1443);
nor U1897 (N_1897,N_1476,N_1351);
and U1898 (N_1898,N_1136,N_1365);
and U1899 (N_1899,N_1299,N_1305);
nand U1900 (N_1900,N_1493,N_1460);
xnor U1901 (N_1901,N_1355,N_1329);
nand U1902 (N_1902,N_1109,N_1491);
nand U1903 (N_1903,N_1472,N_1381);
nor U1904 (N_1904,N_1060,N_1296);
nand U1905 (N_1905,N_1204,N_1006);
and U1906 (N_1906,N_1433,N_1290);
xor U1907 (N_1907,N_1461,N_1169);
nand U1908 (N_1908,N_1140,N_1379);
nor U1909 (N_1909,N_1012,N_1372);
nand U1910 (N_1910,N_1161,N_1385);
nand U1911 (N_1911,N_1364,N_1341);
and U1912 (N_1912,N_1238,N_1483);
and U1913 (N_1913,N_1012,N_1157);
and U1914 (N_1914,N_1002,N_1044);
nor U1915 (N_1915,N_1239,N_1209);
nor U1916 (N_1916,N_1041,N_1290);
nand U1917 (N_1917,N_1249,N_1273);
or U1918 (N_1918,N_1292,N_1255);
and U1919 (N_1919,N_1364,N_1179);
or U1920 (N_1920,N_1031,N_1118);
nor U1921 (N_1921,N_1014,N_1240);
nor U1922 (N_1922,N_1327,N_1223);
and U1923 (N_1923,N_1307,N_1247);
or U1924 (N_1924,N_1462,N_1219);
xor U1925 (N_1925,N_1476,N_1277);
and U1926 (N_1926,N_1301,N_1260);
or U1927 (N_1927,N_1392,N_1145);
nand U1928 (N_1928,N_1027,N_1473);
nor U1929 (N_1929,N_1463,N_1340);
and U1930 (N_1930,N_1007,N_1255);
or U1931 (N_1931,N_1067,N_1086);
nor U1932 (N_1932,N_1483,N_1040);
and U1933 (N_1933,N_1061,N_1187);
and U1934 (N_1934,N_1298,N_1462);
nor U1935 (N_1935,N_1084,N_1435);
xnor U1936 (N_1936,N_1456,N_1131);
and U1937 (N_1937,N_1468,N_1209);
and U1938 (N_1938,N_1376,N_1125);
and U1939 (N_1939,N_1348,N_1075);
or U1940 (N_1940,N_1234,N_1193);
and U1941 (N_1941,N_1456,N_1344);
nor U1942 (N_1942,N_1261,N_1143);
and U1943 (N_1943,N_1013,N_1396);
and U1944 (N_1944,N_1241,N_1129);
nand U1945 (N_1945,N_1072,N_1353);
nor U1946 (N_1946,N_1152,N_1219);
nor U1947 (N_1947,N_1399,N_1417);
and U1948 (N_1948,N_1014,N_1325);
nor U1949 (N_1949,N_1096,N_1385);
and U1950 (N_1950,N_1185,N_1372);
nor U1951 (N_1951,N_1356,N_1292);
or U1952 (N_1952,N_1362,N_1039);
nor U1953 (N_1953,N_1089,N_1143);
nor U1954 (N_1954,N_1439,N_1227);
nand U1955 (N_1955,N_1360,N_1011);
nor U1956 (N_1956,N_1263,N_1273);
nand U1957 (N_1957,N_1416,N_1391);
xor U1958 (N_1958,N_1463,N_1265);
nor U1959 (N_1959,N_1298,N_1264);
and U1960 (N_1960,N_1019,N_1375);
nor U1961 (N_1961,N_1284,N_1323);
and U1962 (N_1962,N_1223,N_1496);
nand U1963 (N_1963,N_1470,N_1445);
or U1964 (N_1964,N_1119,N_1396);
and U1965 (N_1965,N_1422,N_1041);
nand U1966 (N_1966,N_1004,N_1173);
nand U1967 (N_1967,N_1315,N_1293);
nand U1968 (N_1968,N_1443,N_1363);
nand U1969 (N_1969,N_1169,N_1054);
nor U1970 (N_1970,N_1169,N_1124);
or U1971 (N_1971,N_1135,N_1465);
or U1972 (N_1972,N_1125,N_1386);
nor U1973 (N_1973,N_1302,N_1409);
nor U1974 (N_1974,N_1154,N_1408);
and U1975 (N_1975,N_1240,N_1007);
nor U1976 (N_1976,N_1198,N_1177);
and U1977 (N_1977,N_1084,N_1069);
and U1978 (N_1978,N_1342,N_1083);
or U1979 (N_1979,N_1024,N_1075);
nor U1980 (N_1980,N_1106,N_1443);
or U1981 (N_1981,N_1471,N_1416);
or U1982 (N_1982,N_1475,N_1168);
and U1983 (N_1983,N_1108,N_1061);
or U1984 (N_1984,N_1128,N_1111);
or U1985 (N_1985,N_1246,N_1296);
or U1986 (N_1986,N_1066,N_1323);
or U1987 (N_1987,N_1231,N_1364);
and U1988 (N_1988,N_1329,N_1375);
and U1989 (N_1989,N_1066,N_1446);
and U1990 (N_1990,N_1425,N_1405);
or U1991 (N_1991,N_1387,N_1120);
nor U1992 (N_1992,N_1059,N_1165);
and U1993 (N_1993,N_1449,N_1149);
or U1994 (N_1994,N_1168,N_1370);
and U1995 (N_1995,N_1187,N_1342);
nor U1996 (N_1996,N_1400,N_1373);
or U1997 (N_1997,N_1226,N_1120);
and U1998 (N_1998,N_1072,N_1425);
nor U1999 (N_1999,N_1049,N_1459);
or U2000 (N_2000,N_1942,N_1655);
nor U2001 (N_2001,N_1637,N_1927);
or U2002 (N_2002,N_1576,N_1989);
nand U2003 (N_2003,N_1725,N_1509);
nand U2004 (N_2004,N_1963,N_1613);
nor U2005 (N_2005,N_1746,N_1717);
nor U2006 (N_2006,N_1667,N_1961);
and U2007 (N_2007,N_1917,N_1599);
nand U2008 (N_2008,N_1805,N_1618);
nand U2009 (N_2009,N_1515,N_1868);
nand U2010 (N_2010,N_1600,N_1561);
xor U2011 (N_2011,N_1593,N_1823);
and U2012 (N_2012,N_1825,N_1871);
nand U2013 (N_2013,N_1731,N_1960);
nand U2014 (N_2014,N_1700,N_1807);
nor U2015 (N_2015,N_1907,N_1730);
and U2016 (N_2016,N_1646,N_1545);
nor U2017 (N_2017,N_1943,N_1589);
or U2018 (N_2018,N_1970,N_1556);
nand U2019 (N_2019,N_1993,N_1761);
and U2020 (N_2020,N_1672,N_1581);
or U2021 (N_2021,N_1521,N_1912);
nand U2022 (N_2022,N_1678,N_1659);
nand U2023 (N_2023,N_1718,N_1842);
and U2024 (N_2024,N_1552,N_1564);
nor U2025 (N_2025,N_1844,N_1573);
xor U2026 (N_2026,N_1981,N_1565);
and U2027 (N_2027,N_1918,N_1703);
and U2028 (N_2028,N_1772,N_1794);
nand U2029 (N_2029,N_1550,N_1950);
nor U2030 (N_2030,N_1741,N_1877);
or U2031 (N_2031,N_1768,N_1585);
nand U2032 (N_2032,N_1607,N_1806);
or U2033 (N_2033,N_1959,N_1568);
or U2034 (N_2034,N_1929,N_1894);
and U2035 (N_2035,N_1559,N_1691);
and U2036 (N_2036,N_1699,N_1873);
and U2037 (N_2037,N_1834,N_1598);
nand U2038 (N_2038,N_1850,N_1945);
nand U2039 (N_2039,N_1533,N_1606);
and U2040 (N_2040,N_1546,N_1715);
or U2041 (N_2041,N_1903,N_1542);
nand U2042 (N_2042,N_1722,N_1865);
and U2043 (N_2043,N_1940,N_1838);
or U2044 (N_2044,N_1821,N_1944);
or U2045 (N_2045,N_1875,N_1810);
and U2046 (N_2046,N_1681,N_1666);
nand U2047 (N_2047,N_1892,N_1733);
and U2048 (N_2048,N_1904,N_1629);
nor U2049 (N_2049,N_1974,N_1849);
and U2050 (N_2050,N_1841,N_1994);
nand U2051 (N_2051,N_1740,N_1986);
nand U2052 (N_2052,N_1701,N_1869);
nand U2053 (N_2053,N_1935,N_1665);
nor U2054 (N_2054,N_1636,N_1967);
or U2055 (N_2055,N_1610,N_1764);
and U2056 (N_2056,N_1888,N_1955);
and U2057 (N_2057,N_1640,N_1962);
nor U2058 (N_2058,N_1574,N_1743);
nor U2059 (N_2059,N_1978,N_1669);
nor U2060 (N_2060,N_1774,N_1985);
and U2061 (N_2061,N_1558,N_1537);
nand U2062 (N_2062,N_1933,N_1815);
or U2063 (N_2063,N_1786,N_1541);
nand U2064 (N_2064,N_1532,N_1987);
nor U2065 (N_2065,N_1922,N_1548);
nor U2066 (N_2066,N_1938,N_1951);
nor U2067 (N_2067,N_1857,N_1853);
xnor U2068 (N_2068,N_1793,N_1964);
nand U2069 (N_2069,N_1779,N_1582);
nor U2070 (N_2070,N_1505,N_1982);
and U2071 (N_2071,N_1555,N_1801);
nand U2072 (N_2072,N_1587,N_1720);
nand U2073 (N_2073,N_1826,N_1642);
and U2074 (N_2074,N_1689,N_1579);
nand U2075 (N_2075,N_1872,N_1980);
and U2076 (N_2076,N_1519,N_1767);
nand U2077 (N_2077,N_1694,N_1921);
or U2078 (N_2078,N_1895,N_1736);
xnor U2079 (N_2079,N_1973,N_1705);
or U2080 (N_2080,N_1780,N_1650);
and U2081 (N_2081,N_1627,N_1712);
nor U2082 (N_2082,N_1831,N_1577);
nor U2083 (N_2083,N_1808,N_1652);
nand U2084 (N_2084,N_1709,N_1508);
nand U2085 (N_2085,N_1608,N_1603);
and U2086 (N_2086,N_1803,N_1939);
or U2087 (N_2087,N_1769,N_1995);
or U2088 (N_2088,N_1797,N_1941);
nor U2089 (N_2089,N_1957,N_1863);
nand U2090 (N_2090,N_1862,N_1504);
or U2091 (N_2091,N_1597,N_1996);
and U2092 (N_2092,N_1855,N_1527);
nand U2093 (N_2093,N_1811,N_1649);
or U2094 (N_2094,N_1592,N_1615);
and U2095 (N_2095,N_1643,N_1664);
nand U2096 (N_2096,N_1612,N_1870);
nor U2097 (N_2097,N_1910,N_1784);
nor U2098 (N_2098,N_1926,N_1824);
and U2099 (N_2099,N_1601,N_1915);
nand U2100 (N_2100,N_1626,N_1817);
nand U2101 (N_2101,N_1557,N_1762);
and U2102 (N_2102,N_1704,N_1638);
nor U2103 (N_2103,N_1832,N_1795);
or U2104 (N_2104,N_1724,N_1583);
nand U2105 (N_2105,N_1711,N_1525);
nand U2106 (N_2106,N_1688,N_1732);
nor U2107 (N_2107,N_1544,N_1859);
and U2108 (N_2108,N_1901,N_1596);
or U2109 (N_2109,N_1748,N_1848);
or U2110 (N_2110,N_1856,N_1734);
nor U2111 (N_2111,N_1773,N_1997);
nand U2112 (N_2112,N_1706,N_1887);
nand U2113 (N_2113,N_1674,N_1516);
nand U2114 (N_2114,N_1983,N_1625);
nor U2115 (N_2115,N_1896,N_1882);
nand U2116 (N_2116,N_1931,N_1551);
or U2117 (N_2117,N_1658,N_1909);
or U2118 (N_2118,N_1991,N_1648);
nor U2119 (N_2119,N_1713,N_1830);
and U2120 (N_2120,N_1539,N_1676);
nor U2121 (N_2121,N_1879,N_1507);
nand U2122 (N_2122,N_1816,N_1549);
nor U2123 (N_2123,N_1881,N_1790);
nor U2124 (N_2124,N_1946,N_1952);
nand U2125 (N_2125,N_1569,N_1632);
or U2126 (N_2126,N_1766,N_1710);
nor U2127 (N_2127,N_1819,N_1670);
nand U2128 (N_2128,N_1682,N_1977);
nand U2129 (N_2129,N_1614,N_1716);
and U2130 (N_2130,N_1889,N_1571);
nor U2131 (N_2131,N_1503,N_1645);
or U2132 (N_2132,N_1822,N_1534);
and U2133 (N_2133,N_1899,N_1885);
or U2134 (N_2134,N_1783,N_1858);
nand U2135 (N_2135,N_1923,N_1671);
nand U2136 (N_2136,N_1753,N_1580);
nor U2137 (N_2137,N_1623,N_1512);
and U2138 (N_2138,N_1570,N_1763);
nand U2139 (N_2139,N_1902,N_1804);
or U2140 (N_2140,N_1647,N_1538);
xnor U2141 (N_2141,N_1540,N_1609);
nor U2142 (N_2142,N_1520,N_1884);
nor U2143 (N_2143,N_1916,N_1644);
and U2144 (N_2144,N_1729,N_1752);
nand U2145 (N_2145,N_1886,N_1880);
or U2146 (N_2146,N_1714,N_1789);
and U2147 (N_2147,N_1616,N_1905);
nand U2148 (N_2148,N_1965,N_1936);
or U2149 (N_2149,N_1953,N_1727);
and U2150 (N_2150,N_1535,N_1878);
and U2151 (N_2151,N_1928,N_1900);
and U2152 (N_2152,N_1777,N_1523);
nor U2153 (N_2153,N_1634,N_1605);
and U2154 (N_2154,N_1782,N_1692);
and U2155 (N_2155,N_1584,N_1968);
nor U2156 (N_2156,N_1814,N_1662);
and U2157 (N_2157,N_1501,N_1698);
nand U2158 (N_2158,N_1990,N_1854);
nand U2159 (N_2159,N_1617,N_1776);
nand U2160 (N_2160,N_1765,N_1791);
or U2161 (N_2161,N_1737,N_1563);
nand U2162 (N_2162,N_1876,N_1781);
nor U2163 (N_2163,N_1526,N_1845);
and U2164 (N_2164,N_1920,N_1680);
or U2165 (N_2165,N_1992,N_1949);
and U2166 (N_2166,N_1620,N_1785);
nor U2167 (N_2167,N_1890,N_1745);
nor U2168 (N_2168,N_1677,N_1972);
or U2169 (N_2169,N_1639,N_1827);
nand U2170 (N_2170,N_1771,N_1751);
or U2171 (N_2171,N_1934,N_1575);
nor U2172 (N_2172,N_1792,N_1820);
and U2173 (N_2173,N_1622,N_1837);
nor U2174 (N_2174,N_1719,N_1663);
nand U2175 (N_2175,N_1693,N_1543);
nor U2176 (N_2176,N_1602,N_1653);
nand U2177 (N_2177,N_1702,N_1852);
nand U2178 (N_2178,N_1624,N_1708);
nor U2179 (N_2179,N_1802,N_1514);
nand U2180 (N_2180,N_1913,N_1760);
or U2181 (N_2181,N_1809,N_1969);
nor U2182 (N_2182,N_1843,N_1511);
nor U2183 (N_2183,N_1954,N_1510);
or U2184 (N_2184,N_1757,N_1518);
nand U2185 (N_2185,N_1937,N_1633);
nand U2186 (N_2186,N_1897,N_1536);
nor U2187 (N_2187,N_1818,N_1586);
nor U2188 (N_2188,N_1898,N_1787);
or U2189 (N_2189,N_1956,N_1828);
and U2190 (N_2190,N_1621,N_1628);
nor U2191 (N_2191,N_1891,N_1813);
xor U2192 (N_2192,N_1998,N_1864);
nand U2193 (N_2193,N_1778,N_1687);
nand U2194 (N_2194,N_1835,N_1911);
nor U2195 (N_2195,N_1775,N_1867);
nor U2196 (N_2196,N_1562,N_1924);
nor U2197 (N_2197,N_1966,N_1707);
nor U2198 (N_2198,N_1798,N_1932);
nor U2199 (N_2199,N_1930,N_1594);
nor U2200 (N_2200,N_1975,N_1979);
and U2201 (N_2201,N_1851,N_1925);
nand U2202 (N_2202,N_1756,N_1742);
nand U2203 (N_2203,N_1661,N_1759);
nand U2204 (N_2204,N_1919,N_1524);
or U2205 (N_2205,N_1947,N_1893);
and U2206 (N_2206,N_1553,N_1630);
nand U2207 (N_2207,N_1723,N_1726);
and U2208 (N_2208,N_1906,N_1800);
and U2209 (N_2209,N_1619,N_1588);
nand U2210 (N_2210,N_1685,N_1560);
nand U2211 (N_2211,N_1590,N_1747);
nor U2212 (N_2212,N_1531,N_1673);
nor U2213 (N_2213,N_1999,N_1744);
nor U2214 (N_2214,N_1988,N_1654);
and U2215 (N_2215,N_1611,N_1529);
or U2216 (N_2216,N_1735,N_1739);
nand U2217 (N_2217,N_1749,N_1738);
and U2218 (N_2218,N_1578,N_1517);
nor U2219 (N_2219,N_1958,N_1506);
nand U2220 (N_2220,N_1971,N_1675);
and U2221 (N_2221,N_1668,N_1839);
or U2222 (N_2222,N_1684,N_1513);
and U2223 (N_2223,N_1572,N_1528);
nand U2224 (N_2224,N_1641,N_1840);
nor U2225 (N_2225,N_1686,N_1522);
or U2226 (N_2226,N_1604,N_1721);
and U2227 (N_2227,N_1554,N_1883);
nor U2228 (N_2228,N_1755,N_1833);
and U2229 (N_2229,N_1812,N_1728);
nor U2230 (N_2230,N_1770,N_1799);
and U2231 (N_2231,N_1591,N_1595);
and U2232 (N_2232,N_1754,N_1860);
nor U2233 (N_2233,N_1696,N_1984);
nor U2234 (N_2234,N_1530,N_1547);
or U2235 (N_2235,N_1847,N_1502);
or U2236 (N_2236,N_1683,N_1690);
nand U2237 (N_2237,N_1976,N_1697);
or U2238 (N_2238,N_1656,N_1500);
or U2239 (N_2239,N_1861,N_1660);
nand U2240 (N_2240,N_1846,N_1914);
and U2241 (N_2241,N_1631,N_1836);
nand U2242 (N_2242,N_1788,N_1651);
nand U2243 (N_2243,N_1948,N_1750);
and U2244 (N_2244,N_1695,N_1866);
or U2245 (N_2245,N_1874,N_1567);
and U2246 (N_2246,N_1908,N_1796);
nor U2247 (N_2247,N_1657,N_1829);
or U2248 (N_2248,N_1758,N_1566);
xnor U2249 (N_2249,N_1679,N_1635);
or U2250 (N_2250,N_1537,N_1918);
nand U2251 (N_2251,N_1638,N_1814);
and U2252 (N_2252,N_1847,N_1710);
or U2253 (N_2253,N_1826,N_1783);
or U2254 (N_2254,N_1989,N_1958);
or U2255 (N_2255,N_1507,N_1618);
nor U2256 (N_2256,N_1582,N_1683);
and U2257 (N_2257,N_1711,N_1503);
and U2258 (N_2258,N_1769,N_1942);
nand U2259 (N_2259,N_1636,N_1929);
nand U2260 (N_2260,N_1818,N_1932);
or U2261 (N_2261,N_1713,N_1782);
xor U2262 (N_2262,N_1575,N_1937);
and U2263 (N_2263,N_1582,N_1610);
and U2264 (N_2264,N_1596,N_1847);
or U2265 (N_2265,N_1891,N_1641);
and U2266 (N_2266,N_1685,N_1576);
nand U2267 (N_2267,N_1810,N_1572);
nor U2268 (N_2268,N_1566,N_1559);
and U2269 (N_2269,N_1570,N_1510);
nor U2270 (N_2270,N_1508,N_1939);
nand U2271 (N_2271,N_1647,N_1569);
and U2272 (N_2272,N_1906,N_1595);
and U2273 (N_2273,N_1677,N_1727);
nor U2274 (N_2274,N_1834,N_1564);
nand U2275 (N_2275,N_1594,N_1792);
and U2276 (N_2276,N_1673,N_1842);
and U2277 (N_2277,N_1856,N_1912);
nor U2278 (N_2278,N_1840,N_1578);
nand U2279 (N_2279,N_1560,N_1853);
or U2280 (N_2280,N_1850,N_1581);
nand U2281 (N_2281,N_1735,N_1798);
or U2282 (N_2282,N_1686,N_1999);
and U2283 (N_2283,N_1782,N_1510);
nor U2284 (N_2284,N_1658,N_1557);
nor U2285 (N_2285,N_1736,N_1808);
and U2286 (N_2286,N_1802,N_1763);
and U2287 (N_2287,N_1649,N_1731);
or U2288 (N_2288,N_1505,N_1752);
nand U2289 (N_2289,N_1545,N_1831);
or U2290 (N_2290,N_1735,N_1835);
nand U2291 (N_2291,N_1505,N_1679);
nand U2292 (N_2292,N_1811,N_1792);
nand U2293 (N_2293,N_1663,N_1607);
or U2294 (N_2294,N_1856,N_1549);
xnor U2295 (N_2295,N_1980,N_1942);
or U2296 (N_2296,N_1826,N_1844);
nor U2297 (N_2297,N_1656,N_1952);
or U2298 (N_2298,N_1583,N_1711);
and U2299 (N_2299,N_1503,N_1525);
and U2300 (N_2300,N_1983,N_1570);
nor U2301 (N_2301,N_1899,N_1728);
nor U2302 (N_2302,N_1732,N_1830);
or U2303 (N_2303,N_1823,N_1828);
nand U2304 (N_2304,N_1713,N_1660);
nand U2305 (N_2305,N_1708,N_1897);
nor U2306 (N_2306,N_1796,N_1575);
nor U2307 (N_2307,N_1912,N_1997);
nand U2308 (N_2308,N_1854,N_1679);
and U2309 (N_2309,N_1978,N_1705);
nor U2310 (N_2310,N_1796,N_1691);
and U2311 (N_2311,N_1560,N_1551);
or U2312 (N_2312,N_1540,N_1890);
nor U2313 (N_2313,N_1578,N_1773);
nor U2314 (N_2314,N_1908,N_1547);
or U2315 (N_2315,N_1569,N_1874);
and U2316 (N_2316,N_1627,N_1699);
nor U2317 (N_2317,N_1814,N_1733);
or U2318 (N_2318,N_1931,N_1779);
and U2319 (N_2319,N_1695,N_1742);
nand U2320 (N_2320,N_1548,N_1742);
nor U2321 (N_2321,N_1519,N_1545);
nor U2322 (N_2322,N_1690,N_1877);
nor U2323 (N_2323,N_1883,N_1525);
nand U2324 (N_2324,N_1918,N_1958);
and U2325 (N_2325,N_1621,N_1547);
nor U2326 (N_2326,N_1779,N_1966);
nor U2327 (N_2327,N_1825,N_1632);
and U2328 (N_2328,N_1787,N_1925);
and U2329 (N_2329,N_1897,N_1857);
or U2330 (N_2330,N_1799,N_1830);
nor U2331 (N_2331,N_1851,N_1828);
nor U2332 (N_2332,N_1533,N_1953);
nor U2333 (N_2333,N_1501,N_1624);
nand U2334 (N_2334,N_1598,N_1588);
nand U2335 (N_2335,N_1626,N_1614);
and U2336 (N_2336,N_1617,N_1753);
or U2337 (N_2337,N_1833,N_1955);
and U2338 (N_2338,N_1548,N_1800);
or U2339 (N_2339,N_1764,N_1523);
nor U2340 (N_2340,N_1721,N_1743);
or U2341 (N_2341,N_1691,N_1849);
or U2342 (N_2342,N_1617,N_1787);
and U2343 (N_2343,N_1628,N_1939);
nand U2344 (N_2344,N_1934,N_1949);
nand U2345 (N_2345,N_1904,N_1721);
nand U2346 (N_2346,N_1948,N_1859);
or U2347 (N_2347,N_1792,N_1731);
and U2348 (N_2348,N_1674,N_1730);
nand U2349 (N_2349,N_1593,N_1503);
nor U2350 (N_2350,N_1970,N_1588);
or U2351 (N_2351,N_1733,N_1522);
and U2352 (N_2352,N_1719,N_1939);
nand U2353 (N_2353,N_1996,N_1961);
nand U2354 (N_2354,N_1801,N_1644);
and U2355 (N_2355,N_1993,N_1511);
nand U2356 (N_2356,N_1817,N_1943);
or U2357 (N_2357,N_1915,N_1856);
or U2358 (N_2358,N_1946,N_1509);
and U2359 (N_2359,N_1620,N_1664);
nor U2360 (N_2360,N_1936,N_1534);
or U2361 (N_2361,N_1640,N_1928);
nand U2362 (N_2362,N_1984,N_1963);
nor U2363 (N_2363,N_1611,N_1829);
nand U2364 (N_2364,N_1933,N_1974);
nor U2365 (N_2365,N_1760,N_1782);
nand U2366 (N_2366,N_1853,N_1697);
nand U2367 (N_2367,N_1522,N_1985);
or U2368 (N_2368,N_1752,N_1987);
or U2369 (N_2369,N_1663,N_1686);
and U2370 (N_2370,N_1900,N_1870);
nand U2371 (N_2371,N_1964,N_1525);
or U2372 (N_2372,N_1699,N_1816);
or U2373 (N_2373,N_1693,N_1876);
nand U2374 (N_2374,N_1504,N_1767);
or U2375 (N_2375,N_1817,N_1522);
nand U2376 (N_2376,N_1873,N_1761);
or U2377 (N_2377,N_1949,N_1571);
or U2378 (N_2378,N_1867,N_1581);
nor U2379 (N_2379,N_1649,N_1884);
nor U2380 (N_2380,N_1887,N_1769);
nand U2381 (N_2381,N_1910,N_1752);
nand U2382 (N_2382,N_1768,N_1545);
nor U2383 (N_2383,N_1815,N_1616);
or U2384 (N_2384,N_1829,N_1729);
or U2385 (N_2385,N_1969,N_1782);
and U2386 (N_2386,N_1873,N_1502);
nand U2387 (N_2387,N_1967,N_1514);
nand U2388 (N_2388,N_1740,N_1651);
nand U2389 (N_2389,N_1772,N_1586);
nor U2390 (N_2390,N_1677,N_1844);
and U2391 (N_2391,N_1788,N_1767);
or U2392 (N_2392,N_1976,N_1749);
or U2393 (N_2393,N_1833,N_1535);
nor U2394 (N_2394,N_1958,N_1984);
nor U2395 (N_2395,N_1965,N_1847);
and U2396 (N_2396,N_1706,N_1909);
or U2397 (N_2397,N_1878,N_1719);
or U2398 (N_2398,N_1768,N_1748);
or U2399 (N_2399,N_1766,N_1566);
nor U2400 (N_2400,N_1539,N_1945);
and U2401 (N_2401,N_1945,N_1867);
nor U2402 (N_2402,N_1513,N_1720);
or U2403 (N_2403,N_1591,N_1618);
nand U2404 (N_2404,N_1839,N_1650);
or U2405 (N_2405,N_1519,N_1574);
nor U2406 (N_2406,N_1571,N_1899);
nand U2407 (N_2407,N_1508,N_1736);
or U2408 (N_2408,N_1729,N_1570);
nor U2409 (N_2409,N_1823,N_1785);
nor U2410 (N_2410,N_1651,N_1820);
xnor U2411 (N_2411,N_1522,N_1910);
nand U2412 (N_2412,N_1909,N_1791);
and U2413 (N_2413,N_1989,N_1618);
nor U2414 (N_2414,N_1976,N_1858);
or U2415 (N_2415,N_1616,N_1549);
or U2416 (N_2416,N_1833,N_1771);
and U2417 (N_2417,N_1515,N_1569);
and U2418 (N_2418,N_1713,N_1530);
and U2419 (N_2419,N_1603,N_1648);
nand U2420 (N_2420,N_1834,N_1974);
nand U2421 (N_2421,N_1939,N_1613);
nor U2422 (N_2422,N_1735,N_1585);
and U2423 (N_2423,N_1872,N_1987);
or U2424 (N_2424,N_1801,N_1609);
or U2425 (N_2425,N_1815,N_1915);
nor U2426 (N_2426,N_1901,N_1913);
nor U2427 (N_2427,N_1844,N_1615);
nand U2428 (N_2428,N_1536,N_1849);
or U2429 (N_2429,N_1514,N_1632);
nor U2430 (N_2430,N_1765,N_1803);
or U2431 (N_2431,N_1919,N_1856);
nand U2432 (N_2432,N_1505,N_1527);
nand U2433 (N_2433,N_1608,N_1631);
or U2434 (N_2434,N_1942,N_1564);
or U2435 (N_2435,N_1930,N_1864);
or U2436 (N_2436,N_1536,N_1719);
or U2437 (N_2437,N_1676,N_1544);
nor U2438 (N_2438,N_1979,N_1898);
nor U2439 (N_2439,N_1711,N_1853);
nand U2440 (N_2440,N_1838,N_1745);
xnor U2441 (N_2441,N_1583,N_1922);
and U2442 (N_2442,N_1911,N_1653);
nand U2443 (N_2443,N_1936,N_1943);
nor U2444 (N_2444,N_1635,N_1742);
and U2445 (N_2445,N_1524,N_1918);
or U2446 (N_2446,N_1927,N_1616);
xor U2447 (N_2447,N_1583,N_1570);
nand U2448 (N_2448,N_1873,N_1541);
or U2449 (N_2449,N_1696,N_1554);
or U2450 (N_2450,N_1776,N_1517);
nor U2451 (N_2451,N_1877,N_1526);
nand U2452 (N_2452,N_1697,N_1521);
and U2453 (N_2453,N_1706,N_1621);
nor U2454 (N_2454,N_1905,N_1524);
and U2455 (N_2455,N_1760,N_1995);
nand U2456 (N_2456,N_1702,N_1537);
nand U2457 (N_2457,N_1666,N_1723);
xnor U2458 (N_2458,N_1670,N_1838);
nand U2459 (N_2459,N_1896,N_1751);
and U2460 (N_2460,N_1670,N_1663);
nor U2461 (N_2461,N_1896,N_1981);
or U2462 (N_2462,N_1679,N_1839);
nor U2463 (N_2463,N_1609,N_1796);
nand U2464 (N_2464,N_1832,N_1651);
or U2465 (N_2465,N_1604,N_1667);
nor U2466 (N_2466,N_1769,N_1676);
nor U2467 (N_2467,N_1532,N_1990);
xor U2468 (N_2468,N_1996,N_1518);
nor U2469 (N_2469,N_1711,N_1768);
and U2470 (N_2470,N_1995,N_1634);
and U2471 (N_2471,N_1896,N_1683);
nand U2472 (N_2472,N_1538,N_1887);
or U2473 (N_2473,N_1524,N_1687);
and U2474 (N_2474,N_1864,N_1963);
nor U2475 (N_2475,N_1801,N_1674);
or U2476 (N_2476,N_1779,N_1707);
nand U2477 (N_2477,N_1719,N_1628);
nand U2478 (N_2478,N_1716,N_1896);
nor U2479 (N_2479,N_1907,N_1739);
and U2480 (N_2480,N_1548,N_1618);
or U2481 (N_2481,N_1729,N_1559);
nor U2482 (N_2482,N_1989,N_1852);
nor U2483 (N_2483,N_1566,N_1633);
or U2484 (N_2484,N_1638,N_1870);
nor U2485 (N_2485,N_1660,N_1612);
or U2486 (N_2486,N_1518,N_1675);
or U2487 (N_2487,N_1648,N_1935);
and U2488 (N_2488,N_1532,N_1550);
and U2489 (N_2489,N_1958,N_1812);
or U2490 (N_2490,N_1504,N_1634);
nor U2491 (N_2491,N_1896,N_1642);
nor U2492 (N_2492,N_1614,N_1711);
nor U2493 (N_2493,N_1662,N_1546);
nand U2494 (N_2494,N_1506,N_1564);
and U2495 (N_2495,N_1985,N_1816);
or U2496 (N_2496,N_1747,N_1817);
or U2497 (N_2497,N_1887,N_1635);
and U2498 (N_2498,N_1610,N_1765);
nand U2499 (N_2499,N_1810,N_1656);
xnor U2500 (N_2500,N_2188,N_2049);
nand U2501 (N_2501,N_2157,N_2177);
nor U2502 (N_2502,N_2370,N_2489);
nand U2503 (N_2503,N_2119,N_2462);
nor U2504 (N_2504,N_2397,N_2291);
or U2505 (N_2505,N_2338,N_2217);
nor U2506 (N_2506,N_2421,N_2176);
or U2507 (N_2507,N_2463,N_2496);
and U2508 (N_2508,N_2237,N_2240);
and U2509 (N_2509,N_2303,N_2024);
or U2510 (N_2510,N_2021,N_2061);
nand U2511 (N_2511,N_2484,N_2435);
nand U2512 (N_2512,N_2043,N_2464);
or U2513 (N_2513,N_2292,N_2116);
or U2514 (N_2514,N_2098,N_2352);
nand U2515 (N_2515,N_2138,N_2159);
or U2516 (N_2516,N_2124,N_2359);
nor U2517 (N_2517,N_2473,N_2185);
nand U2518 (N_2518,N_2284,N_2209);
and U2519 (N_2519,N_2218,N_2206);
or U2520 (N_2520,N_2114,N_2332);
or U2521 (N_2521,N_2244,N_2305);
and U2522 (N_2522,N_2314,N_2055);
nand U2523 (N_2523,N_2497,N_2082);
or U2524 (N_2524,N_2113,N_2310);
nand U2525 (N_2525,N_2155,N_2200);
nor U2526 (N_2526,N_2219,N_2014);
nand U2527 (N_2527,N_2450,N_2094);
or U2528 (N_2528,N_2101,N_2153);
or U2529 (N_2529,N_2488,N_2449);
and U2530 (N_2530,N_2319,N_2042);
or U2531 (N_2531,N_2266,N_2053);
nor U2532 (N_2532,N_2459,N_2100);
nor U2533 (N_2533,N_2143,N_2228);
and U2534 (N_2534,N_2365,N_2036);
or U2535 (N_2535,N_2327,N_2348);
nand U2536 (N_2536,N_2045,N_2372);
and U2537 (N_2537,N_2181,N_2440);
or U2538 (N_2538,N_2039,N_2429);
xor U2539 (N_2539,N_2447,N_2382);
and U2540 (N_2540,N_2309,N_2202);
nor U2541 (N_2541,N_2121,N_2445);
and U2542 (N_2542,N_2135,N_2412);
nor U2543 (N_2543,N_2477,N_2080);
and U2544 (N_2544,N_2416,N_2354);
nor U2545 (N_2545,N_2057,N_2164);
nor U2546 (N_2546,N_2264,N_2499);
or U2547 (N_2547,N_2278,N_2259);
nor U2548 (N_2548,N_2443,N_2187);
nor U2549 (N_2549,N_2004,N_2019);
nand U2550 (N_2550,N_2353,N_2168);
nor U2551 (N_2551,N_2142,N_2469);
or U2552 (N_2552,N_2406,N_2417);
or U2553 (N_2553,N_2481,N_2494);
nor U2554 (N_2554,N_2232,N_2199);
or U2555 (N_2555,N_2350,N_2368);
or U2556 (N_2556,N_2363,N_2051);
nor U2557 (N_2557,N_2169,N_2016);
and U2558 (N_2558,N_2204,N_2261);
nand U2559 (N_2559,N_2180,N_2029);
or U2560 (N_2560,N_2070,N_2038);
and U2561 (N_2561,N_2380,N_2152);
and U2562 (N_2562,N_2133,N_2022);
nand U2563 (N_2563,N_2331,N_2106);
nor U2564 (N_2564,N_2139,N_2110);
or U2565 (N_2565,N_2233,N_2063);
nand U2566 (N_2566,N_2174,N_2461);
or U2567 (N_2567,N_2282,N_2486);
and U2568 (N_2568,N_2025,N_2230);
nor U2569 (N_2569,N_2222,N_2144);
or U2570 (N_2570,N_2103,N_2326);
and U2571 (N_2571,N_2383,N_2156);
or U2572 (N_2572,N_2125,N_2020);
and U2573 (N_2573,N_2446,N_2394);
nand U2574 (N_2574,N_2179,N_2288);
nand U2575 (N_2575,N_2092,N_2026);
nand U2576 (N_2576,N_2392,N_2492);
or U2577 (N_2577,N_2079,N_2283);
and U2578 (N_2578,N_2250,N_2148);
or U2579 (N_2579,N_2102,N_2298);
nor U2580 (N_2580,N_2387,N_2192);
and U2581 (N_2581,N_2431,N_2369);
xor U2582 (N_2582,N_2472,N_2050);
or U2583 (N_2583,N_2328,N_2318);
nand U2584 (N_2584,N_2090,N_2377);
or U2585 (N_2585,N_2393,N_2415);
or U2586 (N_2586,N_2389,N_2322);
or U2587 (N_2587,N_2189,N_2274);
nor U2588 (N_2588,N_2088,N_2078);
or U2589 (N_2589,N_2273,N_2210);
nand U2590 (N_2590,N_2207,N_2031);
and U2591 (N_2591,N_2149,N_2136);
and U2592 (N_2592,N_2493,N_2035);
nor U2593 (N_2593,N_2410,N_2251);
nand U2594 (N_2594,N_2003,N_2112);
or U2595 (N_2595,N_2087,N_2236);
nand U2596 (N_2596,N_2052,N_2089);
and U2597 (N_2597,N_2211,N_2467);
nand U2598 (N_2598,N_2011,N_2028);
nor U2599 (N_2599,N_2468,N_2123);
and U2600 (N_2600,N_2085,N_2256);
nand U2601 (N_2601,N_2096,N_2279);
nand U2602 (N_2602,N_2300,N_2041);
and U2603 (N_2603,N_2194,N_2296);
and U2604 (N_2604,N_2427,N_2390);
and U2605 (N_2605,N_2321,N_2018);
or U2606 (N_2606,N_2109,N_2171);
nand U2607 (N_2607,N_2460,N_2301);
or U2608 (N_2608,N_2441,N_2404);
nand U2609 (N_2609,N_2229,N_2347);
and U2610 (N_2610,N_2295,N_2485);
or U2611 (N_2611,N_2379,N_2285);
nor U2612 (N_2612,N_2411,N_2442);
nor U2613 (N_2613,N_2341,N_2430);
or U2614 (N_2614,N_2023,N_2239);
or U2615 (N_2615,N_2474,N_2129);
nor U2616 (N_2616,N_2386,N_2358);
nor U2617 (N_2617,N_2084,N_2315);
nand U2618 (N_2618,N_2466,N_2452);
nand U2619 (N_2619,N_2190,N_2306);
and U2620 (N_2620,N_2356,N_2099);
nand U2621 (N_2621,N_2420,N_2059);
and U2622 (N_2622,N_2402,N_2267);
and U2623 (N_2623,N_2032,N_2175);
nand U2624 (N_2624,N_2215,N_2374);
nor U2625 (N_2625,N_2037,N_2077);
nor U2626 (N_2626,N_2165,N_2064);
or U2627 (N_2627,N_2196,N_2373);
nand U2628 (N_2628,N_2396,N_2198);
nand U2629 (N_2629,N_2208,N_2060);
and U2630 (N_2630,N_2360,N_2095);
nand U2631 (N_2631,N_2405,N_2453);
and U2632 (N_2632,N_2010,N_2172);
or U2633 (N_2633,N_2317,N_2034);
and U2634 (N_2634,N_2375,N_2069);
and U2635 (N_2635,N_2105,N_2223);
nand U2636 (N_2636,N_2128,N_2395);
nor U2637 (N_2637,N_2361,N_2161);
and U2638 (N_2638,N_2436,N_2480);
and U2639 (N_2639,N_2150,N_2293);
nor U2640 (N_2640,N_2276,N_2400);
and U2641 (N_2641,N_2241,N_2399);
and U2642 (N_2642,N_2357,N_2335);
nor U2643 (N_2643,N_2257,N_2071);
or U2644 (N_2644,N_2245,N_2238);
nand U2645 (N_2645,N_2478,N_2479);
nand U2646 (N_2646,N_2433,N_2140);
or U2647 (N_2647,N_2158,N_2065);
nor U2648 (N_2648,N_2195,N_2385);
and U2649 (N_2649,N_2281,N_2455);
nand U2650 (N_2650,N_2253,N_2068);
and U2651 (N_2651,N_2255,N_2490);
nor U2652 (N_2652,N_2235,N_2265);
or U2653 (N_2653,N_2173,N_2339);
and U2654 (N_2654,N_2307,N_2482);
and U2655 (N_2655,N_2002,N_2491);
nor U2656 (N_2656,N_2424,N_2132);
or U2657 (N_2657,N_2419,N_2277);
or U2658 (N_2658,N_2407,N_2366);
nand U2659 (N_2659,N_2438,N_2439);
and U2660 (N_2660,N_2127,N_2378);
and U2661 (N_2661,N_2312,N_2117);
nand U2662 (N_2662,N_2345,N_2403);
nand U2663 (N_2663,N_2231,N_2476);
nor U2664 (N_2664,N_2330,N_2226);
nor U2665 (N_2665,N_2213,N_2391);
or U2666 (N_2666,N_2289,N_2325);
nor U2667 (N_2667,N_2304,N_2349);
and U2668 (N_2668,N_2268,N_2000);
nand U2669 (N_2669,N_2294,N_2048);
or U2670 (N_2670,N_2444,N_2362);
nor U2671 (N_2671,N_2252,N_2437);
nand U2672 (N_2672,N_2111,N_2495);
or U2673 (N_2673,N_2083,N_2457);
nand U2674 (N_2674,N_2333,N_2220);
nand U2675 (N_2675,N_2007,N_2093);
or U2676 (N_2676,N_2316,N_2081);
nand U2677 (N_2677,N_2141,N_2227);
xor U2678 (N_2678,N_2160,N_2418);
nand U2679 (N_2679,N_2147,N_2414);
nor U2680 (N_2680,N_2320,N_2201);
nand U2681 (N_2681,N_2425,N_2115);
nor U2682 (N_2682,N_2324,N_2342);
and U2683 (N_2683,N_2146,N_2280);
and U2684 (N_2684,N_2337,N_2299);
or U2685 (N_2685,N_2498,N_2334);
nand U2686 (N_2686,N_2166,N_2254);
nand U2687 (N_2687,N_2047,N_2302);
and U2688 (N_2688,N_2475,N_2262);
nor U2689 (N_2689,N_2074,N_2044);
nand U2690 (N_2690,N_2458,N_2184);
nor U2691 (N_2691,N_2263,N_2163);
or U2692 (N_2692,N_2046,N_2062);
nor U2693 (N_2693,N_2008,N_2423);
nor U2694 (N_2694,N_2009,N_2154);
or U2695 (N_2695,N_2308,N_2367);
or U2696 (N_2696,N_2027,N_2336);
and U2697 (N_2697,N_2162,N_2182);
nor U2698 (N_2698,N_2428,N_2167);
nand U2699 (N_2699,N_2072,N_2371);
nor U2700 (N_2700,N_2448,N_2130);
nor U2701 (N_2701,N_2040,N_2247);
nand U2702 (N_2702,N_2340,N_2323);
nor U2703 (N_2703,N_2270,N_2183);
xnor U2704 (N_2704,N_2122,N_2216);
nand U2705 (N_2705,N_2178,N_2422);
or U2706 (N_2706,N_2091,N_2454);
nand U2707 (N_2707,N_2271,N_2408);
and U2708 (N_2708,N_2013,N_2001);
nor U2709 (N_2709,N_2234,N_2398);
nor U2710 (N_2710,N_2145,N_2248);
and U2711 (N_2711,N_2134,N_2269);
or U2712 (N_2712,N_2203,N_2005);
or U2713 (N_2713,N_2104,N_2033);
and U2714 (N_2714,N_2272,N_2388);
nand U2715 (N_2715,N_2243,N_2214);
and U2716 (N_2716,N_2191,N_2355);
or U2717 (N_2717,N_2108,N_2413);
nor U2718 (N_2718,N_2170,N_2225);
nand U2719 (N_2719,N_2351,N_2017);
nand U2720 (N_2720,N_2076,N_2205);
or U2721 (N_2721,N_2287,N_2451);
or U2722 (N_2722,N_2275,N_2401);
or U2723 (N_2723,N_2120,N_2483);
nand U2724 (N_2724,N_2426,N_2197);
nand U2725 (N_2725,N_2456,N_2151);
nand U2726 (N_2726,N_2073,N_2487);
nor U2727 (N_2727,N_2056,N_2137);
or U2728 (N_2728,N_2432,N_2364);
nand U2729 (N_2729,N_2344,N_2118);
and U2730 (N_2730,N_2471,N_2376);
nand U2731 (N_2731,N_2311,N_2381);
and U2732 (N_2732,N_2258,N_2260);
and U2733 (N_2733,N_2058,N_2054);
or U2734 (N_2734,N_2107,N_2346);
nor U2735 (N_2735,N_2470,N_2030);
nand U2736 (N_2736,N_2186,N_2246);
xor U2737 (N_2737,N_2313,N_2224);
nor U2738 (N_2738,N_2075,N_2242);
or U2739 (N_2739,N_2015,N_2297);
nand U2740 (N_2740,N_2434,N_2290);
nor U2741 (N_2741,N_2329,N_2286);
nor U2742 (N_2742,N_2097,N_2066);
and U2743 (N_2743,N_2006,N_2067);
nor U2744 (N_2744,N_2212,N_2221);
or U2745 (N_2745,N_2465,N_2193);
or U2746 (N_2746,N_2343,N_2249);
nand U2747 (N_2747,N_2126,N_2384);
nand U2748 (N_2748,N_2131,N_2409);
nor U2749 (N_2749,N_2012,N_2086);
nor U2750 (N_2750,N_2455,N_2339);
or U2751 (N_2751,N_2121,N_2133);
nand U2752 (N_2752,N_2012,N_2210);
nor U2753 (N_2753,N_2133,N_2141);
nor U2754 (N_2754,N_2468,N_2461);
nor U2755 (N_2755,N_2498,N_2456);
and U2756 (N_2756,N_2210,N_2054);
or U2757 (N_2757,N_2227,N_2335);
or U2758 (N_2758,N_2248,N_2082);
or U2759 (N_2759,N_2197,N_2250);
nor U2760 (N_2760,N_2455,N_2356);
and U2761 (N_2761,N_2333,N_2289);
and U2762 (N_2762,N_2317,N_2103);
and U2763 (N_2763,N_2402,N_2380);
nor U2764 (N_2764,N_2048,N_2395);
nand U2765 (N_2765,N_2105,N_2186);
nand U2766 (N_2766,N_2097,N_2187);
nand U2767 (N_2767,N_2346,N_2104);
nor U2768 (N_2768,N_2450,N_2194);
nand U2769 (N_2769,N_2131,N_2092);
nor U2770 (N_2770,N_2463,N_2403);
or U2771 (N_2771,N_2008,N_2209);
nand U2772 (N_2772,N_2357,N_2448);
and U2773 (N_2773,N_2463,N_2297);
nor U2774 (N_2774,N_2008,N_2244);
and U2775 (N_2775,N_2277,N_2275);
or U2776 (N_2776,N_2380,N_2379);
and U2777 (N_2777,N_2161,N_2009);
and U2778 (N_2778,N_2448,N_2008);
or U2779 (N_2779,N_2247,N_2395);
and U2780 (N_2780,N_2031,N_2339);
and U2781 (N_2781,N_2446,N_2377);
and U2782 (N_2782,N_2227,N_2276);
or U2783 (N_2783,N_2029,N_2044);
nand U2784 (N_2784,N_2334,N_2030);
and U2785 (N_2785,N_2379,N_2304);
nor U2786 (N_2786,N_2330,N_2319);
or U2787 (N_2787,N_2040,N_2400);
nand U2788 (N_2788,N_2463,N_2013);
or U2789 (N_2789,N_2048,N_2266);
xnor U2790 (N_2790,N_2351,N_2293);
or U2791 (N_2791,N_2047,N_2007);
and U2792 (N_2792,N_2308,N_2190);
nor U2793 (N_2793,N_2186,N_2472);
nor U2794 (N_2794,N_2202,N_2070);
nor U2795 (N_2795,N_2117,N_2116);
nand U2796 (N_2796,N_2185,N_2059);
nor U2797 (N_2797,N_2146,N_2134);
or U2798 (N_2798,N_2025,N_2425);
or U2799 (N_2799,N_2170,N_2238);
or U2800 (N_2800,N_2009,N_2038);
nand U2801 (N_2801,N_2077,N_2117);
or U2802 (N_2802,N_2159,N_2316);
nand U2803 (N_2803,N_2499,N_2261);
and U2804 (N_2804,N_2078,N_2213);
and U2805 (N_2805,N_2474,N_2301);
nor U2806 (N_2806,N_2237,N_2085);
or U2807 (N_2807,N_2293,N_2162);
or U2808 (N_2808,N_2484,N_2285);
and U2809 (N_2809,N_2383,N_2030);
and U2810 (N_2810,N_2292,N_2234);
and U2811 (N_2811,N_2437,N_2237);
and U2812 (N_2812,N_2386,N_2136);
and U2813 (N_2813,N_2093,N_2282);
nand U2814 (N_2814,N_2407,N_2497);
nor U2815 (N_2815,N_2072,N_2373);
xor U2816 (N_2816,N_2371,N_2218);
and U2817 (N_2817,N_2288,N_2494);
xor U2818 (N_2818,N_2335,N_2103);
or U2819 (N_2819,N_2212,N_2158);
or U2820 (N_2820,N_2089,N_2378);
and U2821 (N_2821,N_2333,N_2394);
nand U2822 (N_2822,N_2040,N_2074);
and U2823 (N_2823,N_2413,N_2332);
and U2824 (N_2824,N_2408,N_2145);
or U2825 (N_2825,N_2125,N_2196);
and U2826 (N_2826,N_2417,N_2258);
nand U2827 (N_2827,N_2102,N_2079);
and U2828 (N_2828,N_2323,N_2479);
nand U2829 (N_2829,N_2220,N_2441);
nor U2830 (N_2830,N_2034,N_2283);
or U2831 (N_2831,N_2089,N_2007);
nand U2832 (N_2832,N_2467,N_2178);
nor U2833 (N_2833,N_2280,N_2170);
and U2834 (N_2834,N_2200,N_2134);
nand U2835 (N_2835,N_2122,N_2402);
nor U2836 (N_2836,N_2257,N_2269);
nor U2837 (N_2837,N_2496,N_2011);
nand U2838 (N_2838,N_2316,N_2170);
nor U2839 (N_2839,N_2168,N_2325);
nand U2840 (N_2840,N_2466,N_2486);
nand U2841 (N_2841,N_2443,N_2264);
or U2842 (N_2842,N_2231,N_2162);
nor U2843 (N_2843,N_2295,N_2035);
nor U2844 (N_2844,N_2180,N_2281);
nand U2845 (N_2845,N_2218,N_2042);
nor U2846 (N_2846,N_2184,N_2239);
or U2847 (N_2847,N_2136,N_2279);
or U2848 (N_2848,N_2133,N_2054);
and U2849 (N_2849,N_2369,N_2247);
and U2850 (N_2850,N_2406,N_2433);
and U2851 (N_2851,N_2093,N_2150);
nor U2852 (N_2852,N_2399,N_2087);
or U2853 (N_2853,N_2338,N_2250);
nand U2854 (N_2854,N_2155,N_2218);
nand U2855 (N_2855,N_2031,N_2377);
nand U2856 (N_2856,N_2472,N_2494);
and U2857 (N_2857,N_2246,N_2386);
or U2858 (N_2858,N_2104,N_2152);
xnor U2859 (N_2859,N_2317,N_2016);
nor U2860 (N_2860,N_2261,N_2327);
nor U2861 (N_2861,N_2433,N_2020);
nor U2862 (N_2862,N_2186,N_2074);
and U2863 (N_2863,N_2272,N_2371);
nand U2864 (N_2864,N_2361,N_2006);
nor U2865 (N_2865,N_2253,N_2056);
nand U2866 (N_2866,N_2332,N_2377);
and U2867 (N_2867,N_2198,N_2269);
nor U2868 (N_2868,N_2296,N_2270);
or U2869 (N_2869,N_2360,N_2252);
and U2870 (N_2870,N_2118,N_2040);
and U2871 (N_2871,N_2386,N_2093);
nor U2872 (N_2872,N_2059,N_2323);
nand U2873 (N_2873,N_2342,N_2456);
nand U2874 (N_2874,N_2121,N_2078);
nor U2875 (N_2875,N_2301,N_2366);
and U2876 (N_2876,N_2450,N_2034);
and U2877 (N_2877,N_2055,N_2287);
and U2878 (N_2878,N_2319,N_2055);
nand U2879 (N_2879,N_2069,N_2025);
nor U2880 (N_2880,N_2174,N_2044);
nand U2881 (N_2881,N_2471,N_2250);
or U2882 (N_2882,N_2411,N_2196);
nor U2883 (N_2883,N_2089,N_2313);
or U2884 (N_2884,N_2201,N_2455);
nand U2885 (N_2885,N_2231,N_2297);
or U2886 (N_2886,N_2036,N_2152);
or U2887 (N_2887,N_2106,N_2090);
nor U2888 (N_2888,N_2234,N_2020);
or U2889 (N_2889,N_2401,N_2084);
nor U2890 (N_2890,N_2486,N_2007);
nand U2891 (N_2891,N_2225,N_2133);
and U2892 (N_2892,N_2427,N_2074);
xor U2893 (N_2893,N_2168,N_2496);
nor U2894 (N_2894,N_2017,N_2310);
or U2895 (N_2895,N_2391,N_2242);
nor U2896 (N_2896,N_2436,N_2424);
nor U2897 (N_2897,N_2351,N_2150);
and U2898 (N_2898,N_2383,N_2351);
nand U2899 (N_2899,N_2145,N_2376);
xor U2900 (N_2900,N_2240,N_2103);
and U2901 (N_2901,N_2217,N_2443);
nor U2902 (N_2902,N_2100,N_2270);
nor U2903 (N_2903,N_2020,N_2149);
nor U2904 (N_2904,N_2353,N_2446);
or U2905 (N_2905,N_2403,N_2273);
nor U2906 (N_2906,N_2093,N_2448);
nand U2907 (N_2907,N_2044,N_2159);
and U2908 (N_2908,N_2346,N_2384);
nand U2909 (N_2909,N_2177,N_2110);
nand U2910 (N_2910,N_2443,N_2078);
and U2911 (N_2911,N_2183,N_2247);
nand U2912 (N_2912,N_2310,N_2225);
and U2913 (N_2913,N_2410,N_2401);
nor U2914 (N_2914,N_2251,N_2186);
nor U2915 (N_2915,N_2039,N_2472);
or U2916 (N_2916,N_2336,N_2047);
nand U2917 (N_2917,N_2475,N_2088);
nand U2918 (N_2918,N_2091,N_2380);
and U2919 (N_2919,N_2185,N_2127);
or U2920 (N_2920,N_2069,N_2390);
and U2921 (N_2921,N_2315,N_2098);
or U2922 (N_2922,N_2275,N_2257);
or U2923 (N_2923,N_2443,N_2490);
nand U2924 (N_2924,N_2021,N_2463);
nand U2925 (N_2925,N_2299,N_2253);
nand U2926 (N_2926,N_2174,N_2422);
or U2927 (N_2927,N_2396,N_2068);
and U2928 (N_2928,N_2393,N_2242);
or U2929 (N_2929,N_2319,N_2307);
and U2930 (N_2930,N_2149,N_2473);
nand U2931 (N_2931,N_2008,N_2077);
or U2932 (N_2932,N_2423,N_2252);
nor U2933 (N_2933,N_2486,N_2311);
nand U2934 (N_2934,N_2137,N_2022);
and U2935 (N_2935,N_2390,N_2225);
nand U2936 (N_2936,N_2439,N_2013);
xor U2937 (N_2937,N_2145,N_2388);
and U2938 (N_2938,N_2265,N_2156);
nor U2939 (N_2939,N_2462,N_2031);
or U2940 (N_2940,N_2346,N_2185);
nand U2941 (N_2941,N_2005,N_2110);
nor U2942 (N_2942,N_2192,N_2212);
nor U2943 (N_2943,N_2023,N_2229);
nand U2944 (N_2944,N_2120,N_2218);
nor U2945 (N_2945,N_2328,N_2305);
or U2946 (N_2946,N_2248,N_2171);
nor U2947 (N_2947,N_2097,N_2406);
or U2948 (N_2948,N_2267,N_2104);
nand U2949 (N_2949,N_2257,N_2402);
xor U2950 (N_2950,N_2414,N_2487);
xor U2951 (N_2951,N_2340,N_2473);
or U2952 (N_2952,N_2462,N_2448);
or U2953 (N_2953,N_2472,N_2167);
and U2954 (N_2954,N_2277,N_2165);
nand U2955 (N_2955,N_2337,N_2229);
or U2956 (N_2956,N_2012,N_2048);
nand U2957 (N_2957,N_2229,N_2308);
and U2958 (N_2958,N_2416,N_2483);
nand U2959 (N_2959,N_2474,N_2457);
or U2960 (N_2960,N_2204,N_2459);
nor U2961 (N_2961,N_2100,N_2408);
nand U2962 (N_2962,N_2122,N_2219);
nand U2963 (N_2963,N_2425,N_2444);
or U2964 (N_2964,N_2342,N_2401);
nand U2965 (N_2965,N_2339,N_2482);
nand U2966 (N_2966,N_2330,N_2311);
or U2967 (N_2967,N_2329,N_2149);
nand U2968 (N_2968,N_2266,N_2208);
and U2969 (N_2969,N_2219,N_2036);
and U2970 (N_2970,N_2095,N_2371);
nor U2971 (N_2971,N_2480,N_2044);
or U2972 (N_2972,N_2339,N_2459);
nand U2973 (N_2973,N_2499,N_2363);
nor U2974 (N_2974,N_2312,N_2428);
and U2975 (N_2975,N_2284,N_2092);
nand U2976 (N_2976,N_2208,N_2460);
nand U2977 (N_2977,N_2301,N_2445);
nor U2978 (N_2978,N_2261,N_2162);
and U2979 (N_2979,N_2482,N_2002);
or U2980 (N_2980,N_2184,N_2313);
nor U2981 (N_2981,N_2249,N_2366);
and U2982 (N_2982,N_2464,N_2449);
or U2983 (N_2983,N_2102,N_2262);
nand U2984 (N_2984,N_2358,N_2239);
and U2985 (N_2985,N_2153,N_2238);
nand U2986 (N_2986,N_2348,N_2128);
or U2987 (N_2987,N_2464,N_2481);
nor U2988 (N_2988,N_2390,N_2030);
nor U2989 (N_2989,N_2119,N_2010);
nor U2990 (N_2990,N_2494,N_2053);
nand U2991 (N_2991,N_2081,N_2384);
nor U2992 (N_2992,N_2427,N_2343);
and U2993 (N_2993,N_2479,N_2115);
nand U2994 (N_2994,N_2210,N_2044);
nand U2995 (N_2995,N_2309,N_2157);
nand U2996 (N_2996,N_2064,N_2453);
nor U2997 (N_2997,N_2414,N_2313);
nor U2998 (N_2998,N_2395,N_2466);
and U2999 (N_2999,N_2111,N_2077);
nor UO_0 (O_0,N_2547,N_2732);
and UO_1 (O_1,N_2845,N_2926);
and UO_2 (O_2,N_2885,N_2994);
nor UO_3 (O_3,N_2898,N_2544);
or UO_4 (O_4,N_2525,N_2857);
nand UO_5 (O_5,N_2522,N_2868);
or UO_6 (O_6,N_2801,N_2741);
nand UO_7 (O_7,N_2592,N_2643);
and UO_8 (O_8,N_2508,N_2862);
nor UO_9 (O_9,N_2852,N_2814);
nand UO_10 (O_10,N_2581,N_2844);
or UO_11 (O_11,N_2934,N_2823);
nand UO_12 (O_12,N_2891,N_2999);
or UO_13 (O_13,N_2510,N_2572);
nor UO_14 (O_14,N_2886,N_2747);
nor UO_15 (O_15,N_2746,N_2545);
nand UO_16 (O_16,N_2662,N_2507);
and UO_17 (O_17,N_2627,N_2760);
nand UO_18 (O_18,N_2523,N_2651);
or UO_19 (O_19,N_2663,N_2719);
xor UO_20 (O_20,N_2693,N_2708);
nor UO_21 (O_21,N_2610,N_2743);
nor UO_22 (O_22,N_2762,N_2751);
nand UO_23 (O_23,N_2820,N_2904);
and UO_24 (O_24,N_2952,N_2988);
nor UO_25 (O_25,N_2511,N_2772);
nand UO_26 (O_26,N_2642,N_2825);
and UO_27 (O_27,N_2556,N_2652);
nand UO_28 (O_28,N_2726,N_2764);
and UO_29 (O_29,N_2593,N_2660);
nor UO_30 (O_30,N_2724,N_2878);
nand UO_31 (O_31,N_2604,N_2661);
xor UO_32 (O_32,N_2799,N_2997);
or UO_33 (O_33,N_2910,N_2615);
and UO_34 (O_34,N_2899,N_2601);
and UO_35 (O_35,N_2786,N_2504);
nand UO_36 (O_36,N_2754,N_2518);
and UO_37 (O_37,N_2935,N_2633);
nor UO_38 (O_38,N_2552,N_2872);
and UO_39 (O_39,N_2861,N_2728);
and UO_40 (O_40,N_2710,N_2815);
nor UO_41 (O_41,N_2846,N_2509);
or UO_42 (O_42,N_2834,N_2722);
and UO_43 (O_43,N_2500,N_2829);
nand UO_44 (O_44,N_2656,N_2706);
nand UO_45 (O_45,N_2520,N_2915);
and UO_46 (O_46,N_2916,N_2526);
or UO_47 (O_47,N_2625,N_2616);
nor UO_48 (O_48,N_2953,N_2789);
or UO_49 (O_49,N_2513,N_2807);
nor UO_50 (O_50,N_2776,N_2648);
or UO_51 (O_51,N_2958,N_2721);
or UO_52 (O_52,N_2533,N_2683);
and UO_53 (O_53,N_2578,N_2870);
and UO_54 (O_54,N_2516,N_2809);
nor UO_55 (O_55,N_2599,N_2536);
and UO_56 (O_56,N_2647,N_2869);
nand UO_57 (O_57,N_2657,N_2691);
and UO_58 (O_58,N_2745,N_2841);
or UO_59 (O_59,N_2550,N_2827);
nor UO_60 (O_60,N_2680,N_2977);
nand UO_61 (O_61,N_2854,N_2538);
or UO_62 (O_62,N_2811,N_2860);
or UO_63 (O_63,N_2608,N_2636);
and UO_64 (O_64,N_2540,N_2613);
or UO_65 (O_65,N_2539,N_2794);
and UO_66 (O_66,N_2957,N_2569);
nor UO_67 (O_67,N_2871,N_2562);
or UO_68 (O_68,N_2546,N_2781);
and UO_69 (O_69,N_2612,N_2976);
nand UO_70 (O_70,N_2583,N_2750);
or UO_71 (O_71,N_2514,N_2987);
or UO_72 (O_72,N_2541,N_2557);
nor UO_73 (O_73,N_2923,N_2595);
or UO_74 (O_74,N_2911,N_2699);
or UO_75 (O_75,N_2564,N_2646);
nor UO_76 (O_76,N_2694,N_2664);
and UO_77 (O_77,N_2634,N_2905);
and UO_78 (O_78,N_2596,N_2573);
nor UO_79 (O_79,N_2527,N_2998);
and UO_80 (O_80,N_2936,N_2674);
nor UO_81 (O_81,N_2822,N_2549);
nor UO_82 (O_82,N_2949,N_2720);
nor UO_83 (O_83,N_2686,N_2713);
nor UO_84 (O_84,N_2880,N_2836);
nand UO_85 (O_85,N_2990,N_2669);
and UO_86 (O_86,N_2991,N_2687);
nand UO_87 (O_87,N_2995,N_2628);
and UO_88 (O_88,N_2912,N_2902);
nor UO_89 (O_89,N_2787,N_2512);
nor UO_90 (O_90,N_2665,N_2842);
nand UO_91 (O_91,N_2575,N_2524);
or UO_92 (O_92,N_2805,N_2849);
and UO_93 (O_93,N_2968,N_2590);
or UO_94 (O_94,N_2755,N_2875);
nand UO_95 (O_95,N_2874,N_2882);
nor UO_96 (O_96,N_2780,N_2688);
nand UO_97 (O_97,N_2671,N_2808);
nand UO_98 (O_98,N_2890,N_2618);
or UO_99 (O_99,N_2931,N_2913);
and UO_100 (O_100,N_2704,N_2975);
and UO_101 (O_101,N_2919,N_2566);
xor UO_102 (O_102,N_2795,N_2943);
nor UO_103 (O_103,N_2889,N_2587);
and UO_104 (O_104,N_2866,N_2729);
nor UO_105 (O_105,N_2692,N_2503);
and UO_106 (O_106,N_2909,N_2768);
or UO_107 (O_107,N_2757,N_2655);
and UO_108 (O_108,N_2922,N_2756);
nand UO_109 (O_109,N_2532,N_2903);
xor UO_110 (O_110,N_2530,N_2973);
nor UO_111 (O_111,N_2717,N_2939);
xnor UO_112 (O_112,N_2617,N_2961);
nand UO_113 (O_113,N_2812,N_2838);
or UO_114 (O_114,N_2966,N_2576);
or UO_115 (O_115,N_2594,N_2658);
or UO_116 (O_116,N_2983,N_2607);
and UO_117 (O_117,N_2908,N_2588);
and UO_118 (O_118,N_2964,N_2702);
nor UO_119 (O_119,N_2626,N_2734);
nor UO_120 (O_120,N_2597,N_2978);
or UO_121 (O_121,N_2894,N_2676);
and UO_122 (O_122,N_2985,N_2833);
or UO_123 (O_123,N_2640,N_2771);
or UO_124 (O_124,N_2716,N_2748);
or UO_125 (O_125,N_2907,N_2791);
nand UO_126 (O_126,N_2965,N_2816);
or UO_127 (O_127,N_2954,N_2619);
or UO_128 (O_128,N_2956,N_2864);
nand UO_129 (O_129,N_2879,N_2570);
nor UO_130 (O_130,N_2622,N_2621);
nand UO_131 (O_131,N_2979,N_2623);
or UO_132 (O_132,N_2785,N_2817);
nor UO_133 (O_133,N_2832,N_2519);
nand UO_134 (O_134,N_2715,N_2606);
or UO_135 (O_135,N_2737,N_2992);
or UO_136 (O_136,N_2932,N_2560);
and UO_137 (O_137,N_2993,N_2501);
or UO_138 (O_138,N_2804,N_2733);
and UO_139 (O_139,N_2797,N_2897);
xor UO_140 (O_140,N_2609,N_2837);
nand UO_141 (O_141,N_2506,N_2568);
nor UO_142 (O_142,N_2712,N_2782);
nor UO_143 (O_143,N_2537,N_2681);
or UO_144 (O_144,N_2896,N_2502);
or UO_145 (O_145,N_2584,N_2529);
or UO_146 (O_146,N_2873,N_2517);
nor UO_147 (O_147,N_2920,N_2790);
nor UO_148 (O_148,N_2653,N_2802);
or UO_149 (O_149,N_2641,N_2675);
nand UO_150 (O_150,N_2798,N_2843);
nor UO_151 (O_151,N_2586,N_2679);
nor UO_152 (O_152,N_2937,N_2645);
and UO_153 (O_153,N_2918,N_2947);
nand UO_154 (O_154,N_2685,N_2542);
nand UO_155 (O_155,N_2850,N_2725);
nor UO_156 (O_156,N_2826,N_2917);
nor UO_157 (O_157,N_2740,N_2974);
nand UO_158 (O_158,N_2951,N_2638);
and UO_159 (O_159,N_2528,N_2980);
or UO_160 (O_160,N_2859,N_2924);
nand UO_161 (O_161,N_2701,N_2614);
or UO_162 (O_162,N_2515,N_2824);
nand UO_163 (O_163,N_2810,N_2698);
nand UO_164 (O_164,N_2865,N_2773);
nand UO_165 (O_165,N_2666,N_2730);
nor UO_166 (O_166,N_2887,N_2962);
nand UO_167 (O_167,N_2996,N_2742);
and UO_168 (O_168,N_2941,N_2696);
nand UO_169 (O_169,N_2649,N_2598);
nor UO_170 (O_170,N_2883,N_2986);
nor UO_171 (O_171,N_2940,N_2700);
nand UO_172 (O_172,N_2984,N_2690);
or UO_173 (O_173,N_2813,N_2942);
nor UO_174 (O_174,N_2650,N_2806);
and UO_175 (O_175,N_2709,N_2981);
and UO_176 (O_176,N_2603,N_2707);
nand UO_177 (O_177,N_2759,N_2624);
nand UO_178 (O_178,N_2835,N_2777);
or UO_179 (O_179,N_2925,N_2585);
nand UO_180 (O_180,N_2677,N_2858);
and UO_181 (O_181,N_2605,N_2950);
or UO_182 (O_182,N_2901,N_2521);
nand UO_183 (O_183,N_2761,N_2579);
xnor UO_184 (O_184,N_2914,N_2856);
and UO_185 (O_185,N_2689,N_2654);
and UO_186 (O_186,N_2783,N_2774);
nor UO_187 (O_187,N_2863,N_2900);
nand UO_188 (O_188,N_2758,N_2895);
nand UO_189 (O_189,N_2543,N_2629);
and UO_190 (O_190,N_2739,N_2731);
nor UO_191 (O_191,N_2763,N_2946);
nor UO_192 (O_192,N_2611,N_2928);
or UO_193 (O_193,N_2884,N_2793);
and UO_194 (O_194,N_2989,N_2930);
nand UO_195 (O_195,N_2558,N_2705);
nand UO_196 (O_196,N_2784,N_2893);
xor UO_197 (O_197,N_2867,N_2944);
and UO_198 (O_198,N_2554,N_2819);
nand UO_199 (O_199,N_2561,N_2972);
or UO_200 (O_200,N_2788,N_2960);
and UO_201 (O_201,N_2667,N_2531);
and UO_202 (O_202,N_2766,N_2971);
nor UO_203 (O_203,N_2535,N_2955);
nand UO_204 (O_204,N_2567,N_2632);
and UO_205 (O_205,N_2770,N_2959);
nand UO_206 (O_206,N_2600,N_2718);
nand UO_207 (O_207,N_2830,N_2684);
xor UO_208 (O_208,N_2695,N_2591);
and UO_209 (O_209,N_2892,N_2945);
and UO_210 (O_210,N_2853,N_2589);
and UO_211 (O_211,N_2767,N_2505);
and UO_212 (O_212,N_2769,N_2851);
or UO_213 (O_213,N_2792,N_2921);
or UO_214 (O_214,N_2803,N_2775);
nand UO_215 (O_215,N_2565,N_2682);
or UO_216 (O_216,N_2672,N_2723);
or UO_217 (O_217,N_2620,N_2580);
nand UO_218 (O_218,N_2848,N_2635);
nor UO_219 (O_219,N_2796,N_2659);
and UO_220 (O_220,N_2778,N_2582);
nor UO_221 (O_221,N_2828,N_2881);
and UO_222 (O_222,N_2967,N_2563);
nor UO_223 (O_223,N_2602,N_2840);
or UO_224 (O_224,N_2821,N_2779);
nor UO_225 (O_225,N_2673,N_2548);
and UO_226 (O_226,N_2697,N_2982);
nor UO_227 (O_227,N_2736,N_2938);
and UO_228 (O_228,N_2637,N_2752);
nor UO_229 (O_229,N_2847,N_2855);
and UO_230 (O_230,N_2577,N_2551);
or UO_231 (O_231,N_2630,N_2555);
and UO_232 (O_232,N_2571,N_2735);
xor UO_233 (O_233,N_2668,N_2678);
nor UO_234 (O_234,N_2963,N_2639);
nand UO_235 (O_235,N_2644,N_2906);
nor UO_236 (O_236,N_2876,N_2948);
and UO_237 (O_237,N_2559,N_2831);
nand UO_238 (O_238,N_2800,N_2749);
nor UO_239 (O_239,N_2744,N_2927);
nand UO_240 (O_240,N_2969,N_2711);
nor UO_241 (O_241,N_2753,N_2553);
nor UO_242 (O_242,N_2888,N_2534);
or UO_243 (O_243,N_2703,N_2933);
and UO_244 (O_244,N_2929,N_2631);
nor UO_245 (O_245,N_2574,N_2727);
and UO_246 (O_246,N_2877,N_2765);
nand UO_247 (O_247,N_2970,N_2839);
nor UO_248 (O_248,N_2670,N_2738);
nor UO_249 (O_249,N_2818,N_2714);
and UO_250 (O_250,N_2777,N_2714);
nor UO_251 (O_251,N_2845,N_2996);
nand UO_252 (O_252,N_2653,N_2548);
nor UO_253 (O_253,N_2571,N_2965);
nand UO_254 (O_254,N_2554,N_2719);
or UO_255 (O_255,N_2773,N_2506);
nand UO_256 (O_256,N_2783,N_2877);
nor UO_257 (O_257,N_2854,N_2525);
nor UO_258 (O_258,N_2607,N_2990);
and UO_259 (O_259,N_2917,N_2915);
nor UO_260 (O_260,N_2829,N_2872);
or UO_261 (O_261,N_2927,N_2616);
nand UO_262 (O_262,N_2727,N_2521);
and UO_263 (O_263,N_2643,N_2571);
or UO_264 (O_264,N_2694,N_2781);
or UO_265 (O_265,N_2879,N_2506);
nand UO_266 (O_266,N_2801,N_2731);
and UO_267 (O_267,N_2862,N_2642);
nor UO_268 (O_268,N_2515,N_2658);
nand UO_269 (O_269,N_2948,N_2954);
and UO_270 (O_270,N_2796,N_2913);
xnor UO_271 (O_271,N_2599,N_2888);
and UO_272 (O_272,N_2603,N_2778);
nand UO_273 (O_273,N_2761,N_2912);
nor UO_274 (O_274,N_2654,N_2660);
nand UO_275 (O_275,N_2888,N_2812);
nor UO_276 (O_276,N_2539,N_2966);
or UO_277 (O_277,N_2849,N_2998);
nand UO_278 (O_278,N_2565,N_2927);
and UO_279 (O_279,N_2527,N_2938);
or UO_280 (O_280,N_2964,N_2808);
nor UO_281 (O_281,N_2953,N_2798);
nor UO_282 (O_282,N_2716,N_2704);
nor UO_283 (O_283,N_2977,N_2874);
nor UO_284 (O_284,N_2865,N_2982);
and UO_285 (O_285,N_2826,N_2685);
nor UO_286 (O_286,N_2863,N_2725);
and UO_287 (O_287,N_2596,N_2542);
nor UO_288 (O_288,N_2798,N_2872);
or UO_289 (O_289,N_2815,N_2738);
or UO_290 (O_290,N_2837,N_2633);
or UO_291 (O_291,N_2894,N_2741);
or UO_292 (O_292,N_2822,N_2987);
or UO_293 (O_293,N_2519,N_2922);
nand UO_294 (O_294,N_2637,N_2529);
and UO_295 (O_295,N_2554,N_2789);
nor UO_296 (O_296,N_2726,N_2619);
or UO_297 (O_297,N_2755,N_2779);
and UO_298 (O_298,N_2976,N_2515);
or UO_299 (O_299,N_2903,N_2799);
or UO_300 (O_300,N_2931,N_2547);
nor UO_301 (O_301,N_2883,N_2672);
and UO_302 (O_302,N_2949,N_2544);
or UO_303 (O_303,N_2655,N_2774);
nand UO_304 (O_304,N_2792,N_2834);
nand UO_305 (O_305,N_2761,N_2888);
xor UO_306 (O_306,N_2742,N_2915);
or UO_307 (O_307,N_2521,N_2640);
nand UO_308 (O_308,N_2721,N_2657);
or UO_309 (O_309,N_2914,N_2888);
nand UO_310 (O_310,N_2534,N_2519);
nand UO_311 (O_311,N_2518,N_2937);
and UO_312 (O_312,N_2856,N_2799);
or UO_313 (O_313,N_2783,N_2786);
and UO_314 (O_314,N_2561,N_2849);
nor UO_315 (O_315,N_2660,N_2936);
or UO_316 (O_316,N_2690,N_2687);
nor UO_317 (O_317,N_2642,N_2570);
nor UO_318 (O_318,N_2783,N_2831);
nor UO_319 (O_319,N_2699,N_2781);
or UO_320 (O_320,N_2958,N_2806);
nand UO_321 (O_321,N_2874,N_2518);
nand UO_322 (O_322,N_2943,N_2615);
or UO_323 (O_323,N_2968,N_2604);
and UO_324 (O_324,N_2861,N_2545);
and UO_325 (O_325,N_2701,N_2697);
nand UO_326 (O_326,N_2929,N_2722);
or UO_327 (O_327,N_2816,N_2804);
xnor UO_328 (O_328,N_2987,N_2949);
nand UO_329 (O_329,N_2997,N_2719);
and UO_330 (O_330,N_2715,N_2613);
nand UO_331 (O_331,N_2815,N_2999);
or UO_332 (O_332,N_2942,N_2555);
nand UO_333 (O_333,N_2635,N_2991);
nand UO_334 (O_334,N_2927,N_2824);
and UO_335 (O_335,N_2560,N_2871);
nand UO_336 (O_336,N_2670,N_2799);
or UO_337 (O_337,N_2926,N_2745);
nor UO_338 (O_338,N_2966,N_2684);
nand UO_339 (O_339,N_2703,N_2679);
nor UO_340 (O_340,N_2560,N_2611);
or UO_341 (O_341,N_2967,N_2778);
or UO_342 (O_342,N_2977,N_2889);
or UO_343 (O_343,N_2873,N_2796);
nand UO_344 (O_344,N_2596,N_2938);
nand UO_345 (O_345,N_2595,N_2642);
or UO_346 (O_346,N_2951,N_2889);
nor UO_347 (O_347,N_2805,N_2753);
nand UO_348 (O_348,N_2792,N_2681);
and UO_349 (O_349,N_2738,N_2872);
and UO_350 (O_350,N_2944,N_2736);
or UO_351 (O_351,N_2817,N_2824);
and UO_352 (O_352,N_2957,N_2517);
or UO_353 (O_353,N_2657,N_2715);
and UO_354 (O_354,N_2518,N_2917);
nor UO_355 (O_355,N_2836,N_2677);
nor UO_356 (O_356,N_2890,N_2814);
nand UO_357 (O_357,N_2766,N_2984);
nand UO_358 (O_358,N_2972,N_2993);
and UO_359 (O_359,N_2717,N_2988);
or UO_360 (O_360,N_2658,N_2653);
or UO_361 (O_361,N_2952,N_2783);
and UO_362 (O_362,N_2991,N_2751);
nand UO_363 (O_363,N_2956,N_2618);
and UO_364 (O_364,N_2522,N_2708);
or UO_365 (O_365,N_2927,N_2928);
or UO_366 (O_366,N_2715,N_2719);
or UO_367 (O_367,N_2721,N_2703);
nor UO_368 (O_368,N_2596,N_2504);
and UO_369 (O_369,N_2620,N_2873);
or UO_370 (O_370,N_2616,N_2578);
or UO_371 (O_371,N_2534,N_2875);
and UO_372 (O_372,N_2960,N_2596);
and UO_373 (O_373,N_2676,N_2956);
nor UO_374 (O_374,N_2503,N_2850);
and UO_375 (O_375,N_2524,N_2517);
or UO_376 (O_376,N_2630,N_2959);
nand UO_377 (O_377,N_2657,N_2777);
and UO_378 (O_378,N_2504,N_2555);
nand UO_379 (O_379,N_2664,N_2956);
nor UO_380 (O_380,N_2788,N_2618);
nand UO_381 (O_381,N_2991,N_2885);
nand UO_382 (O_382,N_2879,N_2650);
and UO_383 (O_383,N_2967,N_2665);
nor UO_384 (O_384,N_2677,N_2601);
or UO_385 (O_385,N_2922,N_2766);
nand UO_386 (O_386,N_2681,N_2764);
and UO_387 (O_387,N_2676,N_2773);
nor UO_388 (O_388,N_2608,N_2628);
nor UO_389 (O_389,N_2939,N_2550);
or UO_390 (O_390,N_2977,N_2751);
nor UO_391 (O_391,N_2814,N_2816);
nand UO_392 (O_392,N_2656,N_2892);
nand UO_393 (O_393,N_2784,N_2931);
nand UO_394 (O_394,N_2627,N_2842);
nor UO_395 (O_395,N_2909,N_2604);
and UO_396 (O_396,N_2834,N_2538);
nand UO_397 (O_397,N_2512,N_2629);
nor UO_398 (O_398,N_2710,N_2854);
nand UO_399 (O_399,N_2986,N_2941);
nor UO_400 (O_400,N_2765,N_2978);
or UO_401 (O_401,N_2852,N_2799);
or UO_402 (O_402,N_2963,N_2804);
nor UO_403 (O_403,N_2550,N_2791);
nand UO_404 (O_404,N_2544,N_2888);
and UO_405 (O_405,N_2966,N_2798);
and UO_406 (O_406,N_2752,N_2591);
or UO_407 (O_407,N_2749,N_2897);
nand UO_408 (O_408,N_2718,N_2551);
nor UO_409 (O_409,N_2702,N_2691);
nor UO_410 (O_410,N_2657,N_2635);
or UO_411 (O_411,N_2710,N_2632);
nand UO_412 (O_412,N_2543,N_2934);
or UO_413 (O_413,N_2637,N_2617);
and UO_414 (O_414,N_2828,N_2589);
or UO_415 (O_415,N_2771,N_2687);
xnor UO_416 (O_416,N_2687,N_2801);
nand UO_417 (O_417,N_2882,N_2780);
nor UO_418 (O_418,N_2771,N_2524);
nand UO_419 (O_419,N_2766,N_2883);
or UO_420 (O_420,N_2949,N_2914);
or UO_421 (O_421,N_2789,N_2990);
and UO_422 (O_422,N_2916,N_2705);
and UO_423 (O_423,N_2864,N_2658);
or UO_424 (O_424,N_2996,N_2817);
or UO_425 (O_425,N_2899,N_2666);
nand UO_426 (O_426,N_2577,N_2564);
or UO_427 (O_427,N_2858,N_2602);
and UO_428 (O_428,N_2773,N_2800);
and UO_429 (O_429,N_2518,N_2769);
nor UO_430 (O_430,N_2744,N_2892);
nor UO_431 (O_431,N_2823,N_2927);
nor UO_432 (O_432,N_2734,N_2858);
nand UO_433 (O_433,N_2892,N_2787);
and UO_434 (O_434,N_2532,N_2517);
and UO_435 (O_435,N_2754,N_2986);
nor UO_436 (O_436,N_2894,N_2559);
xnor UO_437 (O_437,N_2580,N_2618);
or UO_438 (O_438,N_2960,N_2932);
nor UO_439 (O_439,N_2571,N_2604);
nand UO_440 (O_440,N_2774,N_2941);
and UO_441 (O_441,N_2557,N_2579);
or UO_442 (O_442,N_2840,N_2817);
nor UO_443 (O_443,N_2604,N_2558);
nand UO_444 (O_444,N_2626,N_2524);
nand UO_445 (O_445,N_2527,N_2971);
nor UO_446 (O_446,N_2900,N_2611);
nand UO_447 (O_447,N_2538,N_2802);
or UO_448 (O_448,N_2962,N_2576);
or UO_449 (O_449,N_2711,N_2756);
nand UO_450 (O_450,N_2662,N_2572);
and UO_451 (O_451,N_2558,N_2718);
and UO_452 (O_452,N_2592,N_2742);
nand UO_453 (O_453,N_2710,N_2692);
and UO_454 (O_454,N_2509,N_2771);
and UO_455 (O_455,N_2519,N_2674);
nand UO_456 (O_456,N_2995,N_2930);
and UO_457 (O_457,N_2548,N_2681);
or UO_458 (O_458,N_2577,N_2664);
or UO_459 (O_459,N_2945,N_2888);
nor UO_460 (O_460,N_2785,N_2890);
nand UO_461 (O_461,N_2547,N_2724);
or UO_462 (O_462,N_2548,N_2712);
or UO_463 (O_463,N_2777,N_2779);
and UO_464 (O_464,N_2667,N_2747);
nand UO_465 (O_465,N_2595,N_2891);
nand UO_466 (O_466,N_2516,N_2708);
nor UO_467 (O_467,N_2647,N_2614);
xor UO_468 (O_468,N_2521,N_2752);
nand UO_469 (O_469,N_2952,N_2639);
nor UO_470 (O_470,N_2846,N_2834);
nor UO_471 (O_471,N_2791,N_2801);
nand UO_472 (O_472,N_2597,N_2857);
or UO_473 (O_473,N_2838,N_2963);
or UO_474 (O_474,N_2508,N_2836);
nand UO_475 (O_475,N_2793,N_2874);
and UO_476 (O_476,N_2738,N_2791);
nor UO_477 (O_477,N_2697,N_2684);
and UO_478 (O_478,N_2747,N_2791);
or UO_479 (O_479,N_2933,N_2919);
and UO_480 (O_480,N_2551,N_2568);
or UO_481 (O_481,N_2698,N_2842);
and UO_482 (O_482,N_2702,N_2672);
nor UO_483 (O_483,N_2697,N_2803);
nand UO_484 (O_484,N_2516,N_2801);
and UO_485 (O_485,N_2787,N_2504);
or UO_486 (O_486,N_2998,N_2851);
nand UO_487 (O_487,N_2588,N_2801);
nand UO_488 (O_488,N_2764,N_2593);
and UO_489 (O_489,N_2878,N_2802);
or UO_490 (O_490,N_2893,N_2628);
and UO_491 (O_491,N_2720,N_2761);
or UO_492 (O_492,N_2528,N_2745);
nand UO_493 (O_493,N_2551,N_2960);
nor UO_494 (O_494,N_2832,N_2872);
and UO_495 (O_495,N_2795,N_2886);
or UO_496 (O_496,N_2858,N_2574);
or UO_497 (O_497,N_2859,N_2811);
nor UO_498 (O_498,N_2568,N_2797);
nand UO_499 (O_499,N_2802,N_2746);
endmodule