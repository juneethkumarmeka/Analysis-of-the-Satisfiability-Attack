module basic_3000_30000_3500_25_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_2332,In_116);
or U1 (N_1,In_2974,In_739);
and U2 (N_2,In_1051,In_1435);
xor U3 (N_3,In_1926,In_618);
or U4 (N_4,In_1913,In_2496);
and U5 (N_5,In_370,In_2866);
and U6 (N_6,In_1995,In_1019);
nand U7 (N_7,In_2409,In_406);
xnor U8 (N_8,In_2497,In_1424);
xor U9 (N_9,In_2170,In_340);
nor U10 (N_10,In_863,In_827);
xor U11 (N_11,In_390,In_1123);
nor U12 (N_12,In_2269,In_236);
or U13 (N_13,In_1155,In_2614);
nand U14 (N_14,In_1638,In_1193);
nor U15 (N_15,In_2052,In_2350);
and U16 (N_16,In_2569,In_1356);
nor U17 (N_17,In_1074,In_478);
nand U18 (N_18,In_498,In_2049);
and U19 (N_19,In_612,In_1573);
nand U20 (N_20,In_1788,In_1446);
and U21 (N_21,In_79,In_1731);
and U22 (N_22,In_1598,In_1277);
nand U23 (N_23,In_1951,In_2187);
nand U24 (N_24,In_165,In_287);
xnor U25 (N_25,In_712,In_1223);
nand U26 (N_26,In_1620,In_690);
nand U27 (N_27,In_1642,In_2778);
and U28 (N_28,In_1159,In_1189);
nor U29 (N_29,In_1191,In_708);
xor U30 (N_30,In_846,In_553);
xor U31 (N_31,In_1279,In_417);
nor U32 (N_32,In_2585,In_1048);
and U33 (N_33,In_1254,In_1986);
and U34 (N_34,In_1666,In_2197);
or U35 (N_35,In_1643,In_2067);
nand U36 (N_36,In_2361,In_2270);
nand U37 (N_37,In_2916,In_660);
xnor U38 (N_38,In_2061,In_215);
or U39 (N_39,In_2669,In_1338);
xor U40 (N_40,In_759,In_2991);
or U41 (N_41,In_309,In_344);
nand U42 (N_42,In_798,In_436);
nand U43 (N_43,In_1082,In_2711);
xnor U44 (N_44,In_2157,In_126);
xnor U45 (N_45,In_71,In_350);
nor U46 (N_46,In_1372,In_516);
nor U47 (N_47,In_354,In_844);
nand U48 (N_48,In_1104,In_1410);
nand U49 (N_49,In_1095,In_401);
xor U50 (N_50,In_1534,In_675);
nor U51 (N_51,In_2150,In_1655);
and U52 (N_52,In_962,In_968);
and U53 (N_53,In_931,In_1963);
xnor U54 (N_54,In_1320,In_241);
and U55 (N_55,In_1201,In_2677);
nor U56 (N_56,In_599,In_2486);
or U57 (N_57,In_1807,In_826);
nor U58 (N_58,In_1284,In_565);
nor U59 (N_59,In_369,In_2079);
xor U60 (N_60,In_1991,In_1892);
and U61 (N_61,In_610,In_2848);
xor U62 (N_62,In_2764,In_2248);
or U63 (N_63,In_1239,In_682);
nand U64 (N_64,In_981,In_1618);
nand U65 (N_65,In_2971,In_960);
xnor U66 (N_66,In_2952,In_2356);
xnor U67 (N_67,In_696,In_2667);
and U68 (N_68,In_2771,In_2278);
nand U69 (N_69,In_2675,In_2177);
xnor U70 (N_70,In_2860,In_2640);
xnor U71 (N_71,In_2008,In_2096);
xnor U72 (N_72,In_943,In_509);
xor U73 (N_73,In_490,In_31);
nor U74 (N_74,In_2510,In_520);
xor U75 (N_75,In_328,In_2262);
and U76 (N_76,In_2135,In_469);
or U77 (N_77,In_2584,In_1656);
nand U78 (N_78,In_626,In_159);
and U79 (N_79,In_2163,In_281);
or U80 (N_80,In_1783,In_1779);
xor U81 (N_81,In_1661,In_607);
xor U82 (N_82,In_2593,In_2637);
xor U83 (N_83,In_2845,In_2118);
nor U84 (N_84,In_339,In_2898);
xnor U85 (N_85,In_2399,In_2040);
or U86 (N_86,In_1753,In_1972);
and U87 (N_87,In_1519,In_2457);
nor U88 (N_88,In_249,In_1378);
and U89 (N_89,In_2925,In_2542);
and U90 (N_90,In_997,In_644);
nand U91 (N_91,In_1084,In_2685);
and U92 (N_92,In_546,In_2573);
nand U93 (N_93,In_1557,In_764);
nand U94 (N_94,In_122,In_2029);
nor U95 (N_95,In_2762,In_2671);
nor U96 (N_96,In_464,In_665);
xor U97 (N_97,In_797,In_2415);
xnor U98 (N_98,In_1353,In_1129);
and U99 (N_99,In_754,In_2114);
or U100 (N_100,In_292,In_1778);
and U101 (N_101,In_2220,In_2330);
or U102 (N_102,In_508,In_2038);
and U103 (N_103,In_1025,In_622);
nand U104 (N_104,In_905,In_815);
xnor U105 (N_105,In_1984,In_2224);
nor U106 (N_106,In_1580,In_2741);
or U107 (N_107,In_204,In_902);
nand U108 (N_108,In_2219,In_2620);
and U109 (N_109,In_2055,In_2024);
xor U110 (N_110,In_1358,In_552);
or U111 (N_111,In_1309,In_152);
nand U112 (N_112,In_1131,In_55);
nand U113 (N_113,In_738,In_1158);
nand U114 (N_114,In_1018,In_2865);
or U115 (N_115,In_2093,In_443);
xor U116 (N_116,In_2473,In_1115);
nand U117 (N_117,In_1895,In_955);
or U118 (N_118,In_2401,In_2053);
nor U119 (N_119,In_1975,In_2251);
or U120 (N_120,In_1267,In_1881);
or U121 (N_121,In_744,In_1723);
nor U122 (N_122,In_2723,In_264);
or U123 (N_123,In_2239,In_2698);
nor U124 (N_124,In_1754,In_1287);
xnor U125 (N_125,In_94,In_2470);
nand U126 (N_126,In_2231,In_2390);
nor U127 (N_127,In_2835,In_330);
or U128 (N_128,In_1594,In_314);
xor U129 (N_129,In_101,In_1422);
or U130 (N_130,In_1415,In_2563);
or U131 (N_131,In_310,In_2081);
xor U132 (N_132,In_2891,In_1293);
xor U133 (N_133,In_1872,In_322);
nor U134 (N_134,In_683,In_2126);
and U135 (N_135,In_619,In_468);
or U136 (N_136,In_898,In_2789);
nor U137 (N_137,In_1840,In_2986);
xnor U138 (N_138,In_693,In_1292);
nand U139 (N_139,In_2946,In_1616);
and U140 (N_140,In_25,In_2425);
nand U141 (N_141,In_359,In_1489);
and U142 (N_142,In_1759,In_41);
and U143 (N_143,In_2166,In_1154);
xor U144 (N_144,In_2198,In_2010);
or U145 (N_145,In_2125,In_1015);
nor U146 (N_146,In_1905,In_518);
and U147 (N_147,In_2227,In_2892);
nor U148 (N_148,In_503,In_1752);
nand U149 (N_149,In_1069,In_517);
xnor U150 (N_150,In_2794,In_2805);
nand U151 (N_151,In_111,In_347);
or U152 (N_152,In_2641,In_562);
nand U153 (N_153,In_2403,In_1286);
nand U154 (N_154,In_1175,In_2381);
xnor U155 (N_155,In_691,In_747);
xor U156 (N_156,In_1767,In_1747);
and U157 (N_157,In_991,In_1071);
or U158 (N_158,In_2767,In_2196);
or U159 (N_159,In_1987,In_1760);
nor U160 (N_160,In_2016,In_425);
or U161 (N_161,In_870,In_2749);
xor U162 (N_162,In_641,In_226);
and U163 (N_163,In_2378,In_2562);
or U164 (N_164,In_2026,In_259);
nand U165 (N_165,In_2665,In_1343);
or U166 (N_166,In_2240,In_280);
xnor U167 (N_167,In_1464,In_2992);
nor U168 (N_168,In_2846,In_2368);
and U169 (N_169,In_1829,In_937);
nand U170 (N_170,In_1768,In_1670);
nor U171 (N_171,In_1417,In_2581);
and U172 (N_172,In_2012,In_289);
nor U173 (N_173,In_2937,In_2495);
or U174 (N_174,In_2629,In_2229);
nand U175 (N_175,In_2041,In_2062);
or U176 (N_176,In_1419,In_2632);
nand U177 (N_177,In_629,In_158);
nand U178 (N_178,In_1226,In_2627);
nor U179 (N_179,In_2277,In_1106);
and U180 (N_180,In_1512,In_2357);
nand U181 (N_181,In_1607,In_1225);
xnor U182 (N_182,In_1028,In_1800);
or U183 (N_183,In_2021,In_1936);
nand U184 (N_184,In_2463,In_1550);
nor U185 (N_185,In_647,In_1858);
and U186 (N_186,In_2518,In_2630);
nand U187 (N_187,In_2408,In_582);
or U188 (N_188,In_2327,In_1042);
and U189 (N_189,In_2088,In_849);
nand U190 (N_190,In_1736,In_2070);
and U191 (N_191,In_2343,In_32);
and U192 (N_192,In_2689,In_2142);
nor U193 (N_193,In_623,In_1339);
or U194 (N_194,In_1439,In_709);
nand U195 (N_195,In_2000,In_290);
xnor U196 (N_196,In_2193,In_790);
xor U197 (N_197,In_2259,In_2247);
xnor U198 (N_198,In_242,In_2424);
or U199 (N_199,In_65,In_1562);
or U200 (N_200,In_1163,In_1539);
xor U201 (N_201,In_42,In_632);
and U202 (N_202,In_884,In_631);
xor U203 (N_203,In_185,In_2595);
or U204 (N_204,In_853,In_378);
nor U205 (N_205,In_2571,In_2708);
and U206 (N_206,In_2984,In_1348);
and U207 (N_207,In_2321,In_1669);
nor U208 (N_208,In_49,In_2832);
nand U209 (N_209,In_1693,In_305);
nand U210 (N_210,In_2435,In_2107);
or U211 (N_211,In_2349,In_537);
xor U212 (N_212,In_115,In_365);
or U213 (N_213,In_1344,In_1482);
xnor U214 (N_214,In_2750,In_2017);
nand U215 (N_215,In_2284,In_1849);
xnor U216 (N_216,In_260,In_2333);
nor U217 (N_217,In_2215,In_2046);
or U218 (N_218,In_890,In_166);
and U219 (N_219,In_645,In_1035);
and U220 (N_220,In_2953,In_1382);
or U221 (N_221,In_2793,In_1471);
nand U222 (N_222,In_2309,In_2909);
nor U223 (N_223,In_805,In_2684);
nor U224 (N_224,In_2988,In_557);
nor U225 (N_225,In_1111,In_1043);
and U226 (N_226,In_2483,In_2138);
or U227 (N_227,In_276,In_1234);
nor U228 (N_228,In_2546,In_1192);
nand U229 (N_229,In_1125,In_2606);
or U230 (N_230,In_1981,In_715);
and U231 (N_231,In_1613,In_2951);
or U232 (N_232,In_832,In_2687);
nor U233 (N_233,In_1507,In_878);
nand U234 (N_234,In_345,In_541);
or U235 (N_235,In_1064,In_2642);
and U236 (N_236,In_2738,In_692);
nand U237 (N_237,In_1503,In_1114);
and U238 (N_238,In_2165,In_2590);
nor U239 (N_239,In_2109,In_306);
or U240 (N_240,In_1079,In_1836);
or U241 (N_241,In_1634,In_2926);
xnor U242 (N_242,In_2755,In_59);
nand U243 (N_243,In_1629,In_2252);
xnor U244 (N_244,In_523,In_664);
nand U245 (N_245,In_2131,In_2018);
or U246 (N_246,In_2236,In_448);
xor U247 (N_247,In_1864,In_1671);
or U248 (N_248,In_899,In_2422);
and U249 (N_249,In_2618,In_2790);
and U250 (N_250,In_1817,In_725);
nor U251 (N_251,In_2132,In_2928);
and U252 (N_252,In_2014,In_275);
and U253 (N_253,In_2212,In_942);
or U254 (N_254,In_1894,In_1165);
xor U255 (N_255,In_170,In_2872);
nand U256 (N_256,In_1774,In_1076);
or U257 (N_257,In_203,In_894);
xnor U258 (N_258,In_1238,In_2477);
xor U259 (N_259,In_2548,In_2316);
and U260 (N_260,In_335,In_2837);
xnor U261 (N_261,In_911,In_178);
nor U262 (N_262,In_452,In_1825);
and U263 (N_263,In_1057,In_950);
nand U264 (N_264,In_871,In_2727);
and U265 (N_265,In_1063,In_1097);
nor U266 (N_266,In_1432,In_1797);
xor U267 (N_267,In_1952,In_755);
nor U268 (N_268,In_1928,In_110);
xor U269 (N_269,In_1586,In_1041);
nand U270 (N_270,In_1360,In_1595);
nand U271 (N_271,In_580,In_1566);
nand U272 (N_272,In_296,In_2578);
nor U273 (N_273,In_1861,In_221);
or U274 (N_274,In_829,In_2146);
xnor U275 (N_275,In_394,In_2209);
nand U276 (N_276,In_2940,In_487);
and U277 (N_277,In_2533,In_2244);
nand U278 (N_278,In_1368,In_1182);
and U279 (N_279,In_633,In_2783);
nand U280 (N_280,In_82,In_2842);
or U281 (N_281,In_1515,In_934);
nor U282 (N_282,In_442,In_2869);
and U283 (N_283,In_1449,In_451);
nor U284 (N_284,In_1741,In_820);
and U285 (N_285,In_39,In_160);
and U286 (N_286,In_1603,In_1326);
and U287 (N_287,In_433,In_2704);
nor U288 (N_288,In_1141,In_2376);
nand U289 (N_289,In_661,In_689);
nand U290 (N_290,In_1483,In_2834);
and U291 (N_291,In_2173,In_216);
or U292 (N_292,In_1990,In_2861);
and U293 (N_293,In_76,In_672);
and U294 (N_294,In_3,In_2300);
or U295 (N_295,In_706,In_2084);
and U296 (N_296,In_23,In_1266);
or U297 (N_297,In_2337,In_1870);
and U298 (N_298,In_128,In_893);
nor U299 (N_299,In_1932,In_600);
xor U300 (N_300,In_219,In_1215);
and U301 (N_301,In_1050,In_209);
and U302 (N_302,In_796,In_323);
or U303 (N_303,In_2263,In_1833);
or U304 (N_304,In_1006,In_2976);
nor U305 (N_305,In_2101,In_333);
xnor U306 (N_306,In_1228,In_597);
and U307 (N_307,In_426,In_577);
or U308 (N_308,In_136,In_199);
xnor U309 (N_309,In_956,In_17);
or U310 (N_310,In_717,In_519);
nor U311 (N_311,In_620,In_1649);
or U312 (N_312,In_1506,In_87);
or U313 (N_313,In_234,In_1107);
xor U314 (N_314,In_2127,In_2168);
nand U315 (N_315,In_2206,In_2256);
nand U316 (N_316,In_1709,In_1855);
nand U317 (N_317,In_2526,In_2650);
nand U318 (N_318,In_1472,In_2128);
nor U319 (N_319,In_2394,In_2797);
nor U320 (N_320,In_1322,In_782);
and U321 (N_321,In_2466,In_528);
xnor U322 (N_322,In_2175,In_1965);
nand U323 (N_323,In_1915,In_86);
xnor U324 (N_324,In_367,In_2681);
nor U325 (N_325,In_422,In_247);
nand U326 (N_326,In_2763,In_1688);
xor U327 (N_327,In_1755,In_2739);
nand U328 (N_328,In_2781,In_2815);
nor U329 (N_329,In_2856,In_2480);
and U330 (N_330,In_1806,In_1939);
nor U331 (N_331,In_459,In_1136);
or U332 (N_332,In_1469,In_757);
xnor U333 (N_333,In_285,In_636);
and U334 (N_334,In_804,In_1574);
nor U335 (N_335,In_2897,In_2902);
nand U336 (N_336,In_2078,In_2775);
nand U337 (N_337,In_2977,In_467);
nand U338 (N_338,In_2180,In_402);
and U339 (N_339,In_9,In_1098);
nand U340 (N_340,In_2290,In_1721);
and U341 (N_341,In_527,In_1493);
xnor U342 (N_342,In_977,In_1854);
xnor U343 (N_343,In_2100,In_1186);
and U344 (N_344,In_2002,In_1319);
and U345 (N_345,In_428,In_2978);
xnor U346 (N_346,In_2760,In_2194);
nor U347 (N_347,In_2719,In_2817);
xor U348 (N_348,In_1216,In_1900);
nor U349 (N_349,In_1570,In_2025);
nand U350 (N_350,In_745,In_835);
xor U351 (N_351,In_1707,In_107);
nand U352 (N_352,In_2371,In_726);
nor U353 (N_353,In_2232,In_569);
nand U354 (N_354,In_540,In_2216);
xnor U355 (N_355,In_2450,In_1460);
or U356 (N_356,In_806,In_372);
or U357 (N_357,In_1862,In_2462);
or U358 (N_358,In_512,In_2961);
or U359 (N_359,In_1705,In_2154);
xor U360 (N_360,In_1416,In_2512);
nand U361 (N_361,In_392,In_81);
nand U362 (N_362,In_308,In_1758);
or U363 (N_363,In_767,In_1209);
nor U364 (N_364,In_2785,In_1887);
and U365 (N_365,In_1591,In_84);
nor U366 (N_366,In_2652,In_291);
nor U367 (N_367,In_2963,In_14);
xor U368 (N_368,In_830,In_2700);
xor U369 (N_369,In_793,In_1333);
and U370 (N_370,In_941,In_1860);
nor U371 (N_371,In_1204,In_1834);
or U372 (N_372,In_1185,In_1218);
and U373 (N_373,In_2275,In_180);
or U374 (N_374,In_2970,In_1466);
nand U375 (N_375,In_1233,In_24);
xnor U376 (N_376,In_2134,In_1835);
or U377 (N_377,In_999,In_141);
nand U378 (N_378,In_869,In_2028);
or U379 (N_379,In_2875,In_492);
xnor U380 (N_380,In_2520,In_172);
nor U381 (N_381,In_2661,In_687);
xor U382 (N_382,In_2519,In_1355);
xnor U383 (N_383,In_2812,In_2729);
nor U384 (N_384,In_1997,In_269);
nor U385 (N_385,In_1183,In_2281);
nor U386 (N_386,In_1579,In_1346);
nor U387 (N_387,In_2478,In_1306);
nor U388 (N_388,In_1663,In_1475);
or U389 (N_389,In_2530,In_313);
nor U390 (N_390,In_2124,In_1842);
xnor U391 (N_391,In_2306,In_2319);
or U392 (N_392,In_1636,In_2210);
nand U393 (N_393,In_1176,In_1038);
nand U394 (N_394,In_465,In_2123);
xnor U395 (N_395,In_1946,In_2416);
nand U396 (N_396,In_1062,In_773);
or U397 (N_397,In_1749,In_2862);
or U398 (N_398,In_11,In_2914);
and U399 (N_399,In_1792,In_1756);
nor U400 (N_400,In_720,In_2517);
nand U401 (N_401,In_2452,In_2340);
nor U402 (N_402,In_1942,In_1841);
xor U403 (N_403,In_1011,In_1625);
nor U404 (N_404,In_1032,In_2186);
or U405 (N_405,In_639,In_1787);
xor U406 (N_406,In_2811,In_1815);
and U407 (N_407,In_1605,In_1885);
nand U408 (N_408,In_918,In_1738);
or U409 (N_409,In_375,In_1102);
nor U410 (N_410,In_1013,In_2494);
nand U411 (N_411,In_1884,In_1660);
nand U412 (N_412,In_1350,In_1962);
nand U413 (N_413,In_97,In_2623);
nor U414 (N_414,In_1914,In_892);
nor U415 (N_415,In_1973,In_207);
nand U416 (N_416,In_1197,In_544);
nor U417 (N_417,In_1824,In_1589);
and U418 (N_418,In_2149,In_2857);
nand U419 (N_419,In_1677,In_312);
nand U420 (N_420,In_984,In_674);
xnor U421 (N_421,In_1325,In_2710);
nand U422 (N_422,In_379,In_2130);
or U423 (N_423,In_262,In_381);
or U424 (N_424,In_2151,In_975);
or U425 (N_425,In_2853,In_522);
nor U426 (N_426,In_188,In_535);
or U427 (N_427,In_2703,In_231);
or U428 (N_428,In_2304,In_95);
xnor U429 (N_429,In_928,In_2427);
nand U430 (N_430,In_1392,In_326);
or U431 (N_431,In_2858,In_1804);
and U432 (N_432,In_2476,In_1811);
nor U433 (N_433,In_1664,In_2728);
or U434 (N_434,In_2254,In_1704);
or U435 (N_435,In_51,In_2172);
nor U436 (N_436,In_2679,In_1614);
nand U437 (N_437,In_1575,In_2437);
and U438 (N_438,In_271,In_653);
and U439 (N_439,In_1526,In_1133);
nor U440 (N_440,In_817,In_47);
and U441 (N_441,In_1017,In_1784);
and U442 (N_442,In_455,In_377);
and U443 (N_443,In_676,In_1146);
xnor U444 (N_444,In_64,In_2358);
nand U445 (N_445,In_707,In_1940);
nor U446 (N_446,In_104,In_91);
nand U447 (N_447,In_2391,In_2688);
or U448 (N_448,In_2575,In_2923);
xor U449 (N_449,In_1441,In_1144);
and U450 (N_450,In_48,In_2459);
xnor U451 (N_451,In_2752,In_2110);
and U452 (N_452,In_1801,In_2499);
nand U453 (N_453,In_1726,In_635);
nor U454 (N_454,In_1822,In_385);
xnor U455 (N_455,In_54,In_195);
nand U456 (N_456,In_430,In_1554);
nand U457 (N_457,In_761,In_825);
or U458 (N_458,In_2449,In_2481);
xor U459 (N_459,In_1376,In_1092);
xor U460 (N_460,In_510,In_1949);
nand U461 (N_461,In_1879,In_1604);
or U462 (N_462,In_137,In_945);
nor U463 (N_463,In_60,In_879);
and U464 (N_464,In_901,In_753);
nor U465 (N_465,In_2874,In_954);
or U466 (N_466,In_2178,In_476);
and U467 (N_467,In_2344,In_98);
or U468 (N_468,In_1463,In_658);
xor U469 (N_469,In_189,In_334);
and U470 (N_470,In_1269,In_548);
and U471 (N_471,In_1413,In_662);
xnor U472 (N_472,In_2726,In_1790);
xor U473 (N_473,In_1899,In_1798);
or U474 (N_474,In_1733,In_2912);
or U475 (N_475,In_1901,In_2663);
nand U476 (N_476,In_1569,In_1610);
xnor U477 (N_477,In_1401,In_2831);
nand U478 (N_478,In_1737,In_970);
nand U479 (N_479,In_2328,In_1213);
nand U480 (N_480,In_2448,In_1331);
nand U481 (N_481,In_2164,In_1148);
and U482 (N_482,In_1166,In_1317);
nor U483 (N_483,In_818,In_1716);
nand U484 (N_484,In_2622,In_1179);
xor U485 (N_485,In_1672,In_1933);
and U486 (N_486,In_52,In_2608);
or U487 (N_487,In_716,In_2314);
or U488 (N_488,In_2324,In_888);
nor U489 (N_489,In_1626,In_2199);
xor U490 (N_490,In_1096,In_2160);
nor U491 (N_491,In_1559,In_109);
or U492 (N_492,In_831,In_2336);
nand U493 (N_493,In_803,In_2516);
nand U494 (N_494,In_337,In_1505);
nor U495 (N_495,In_1072,In_2543);
nor U496 (N_496,In_810,In_1044);
xor U497 (N_497,In_2202,In_811);
nand U498 (N_498,In_1711,In_2174);
nor U499 (N_499,In_1762,In_1674);
xnor U500 (N_500,In_1206,In_2718);
and U501 (N_501,In_549,In_923);
and U502 (N_502,In_602,In_2631);
nand U503 (N_503,In_50,In_2768);
and U504 (N_504,In_1468,In_2673);
or U505 (N_505,In_1808,In_646);
and U506 (N_506,In_2936,In_1087);
nand U507 (N_507,In_2929,In_383);
nor U508 (N_508,In_1911,In_1961);
xor U509 (N_509,In_925,In_842);
and U510 (N_510,In_1809,In_2934);
nor U511 (N_511,In_384,In_361);
nor U512 (N_512,In_475,In_2643);
nor U513 (N_513,In_996,In_1130);
nor U514 (N_514,In_2105,In_1746);
or U515 (N_515,In_2318,In_2967);
or U516 (N_516,In_1447,In_1692);
or U517 (N_517,In_1418,In_1280);
nor U518 (N_518,In_438,In_776);
and U519 (N_519,In_61,In_1303);
xnor U520 (N_520,In_1242,In_2464);
nand U521 (N_521,In_123,In_2443);
xor U522 (N_522,In_2057,In_1140);
or U523 (N_523,In_515,In_1295);
nand U524 (N_524,In_2267,In_1727);
nor U525 (N_525,In_824,In_2919);
or U526 (N_526,In_480,In_2558);
or U527 (N_527,In_1897,In_319);
xnor U528 (N_528,In_2887,In_2407);
nand U529 (N_529,In_2830,In_2159);
or U530 (N_530,In_2836,In_307);
xnor U531 (N_531,In_1243,In_2293);
nand U532 (N_532,In_193,In_2504);
xnor U533 (N_533,In_2468,In_457);
or U534 (N_534,In_880,In_261);
nand U535 (N_535,In_2249,In_293);
xor U536 (N_536,In_1918,In_1387);
and U537 (N_537,In_2436,In_2576);
xnor U538 (N_538,In_1135,In_56);
and U539 (N_539,In_415,In_2908);
xor U540 (N_540,In_2871,In_2171);
xnor U541 (N_541,In_2311,In_2523);
xor U542 (N_542,In_1066,In_868);
and U543 (N_543,In_456,In_1437);
nand U544 (N_544,In_1527,In_2555);
xor U545 (N_545,In_2279,In_2471);
xor U546 (N_546,In_867,In_2779);
nand U547 (N_547,In_1706,In_1630);
nand U548 (N_548,In_2522,In_1268);
nor U549 (N_549,In_1099,In_1635);
nor U550 (N_550,In_1820,In_1773);
or U551 (N_551,In_785,In_257);
and U552 (N_552,In_1908,In_2426);
xnor U553 (N_553,In_2372,In_2373);
nor U554 (N_554,In_1,In_1826);
xnor U555 (N_555,In_149,In_2291);
and U556 (N_556,In_601,In_2506);
and U557 (N_557,In_2092,In_2696);
or U558 (N_558,In_2889,In_1001);
and U559 (N_559,In_1480,In_1061);
nand U560 (N_560,In_673,In_765);
xnor U561 (N_561,In_35,In_2648);
nand U562 (N_562,In_2803,In_2037);
nand U563 (N_563,In_446,In_2932);
nand U564 (N_564,In_2264,In_727);
xor U565 (N_565,In_2359,In_325);
nand U566 (N_566,In_2377,In_1196);
nand U567 (N_567,In_801,In_1966);
nor U568 (N_568,In_1113,In_1147);
nor U569 (N_569,In_1717,In_171);
and U570 (N_570,In_2966,In_1985);
nand U571 (N_571,In_2713,In_1304);
xor U572 (N_572,In_729,In_1540);
xnor U573 (N_573,In_1745,In_2852);
nand U574 (N_574,In_238,In_2737);
xor U575 (N_575,In_2716,In_2042);
and U576 (N_576,In_802,In_1349);
xor U577 (N_577,In_883,In_1828);
or U578 (N_578,In_1054,In_2877);
nor U579 (N_579,In_396,In_1298);
nand U580 (N_580,In_2011,In_142);
xnor U581 (N_581,In_988,In_10);
and U582 (N_582,In_2702,In_1763);
xor U583 (N_583,In_1330,In_1149);
nor U584 (N_584,In_591,In_1379);
or U585 (N_585,In_2345,In_2983);
nand U586 (N_586,In_83,In_441);
nand U587 (N_587,In_881,In_714);
nand U588 (N_588,In_1587,In_2500);
and U589 (N_589,In_1549,In_2766);
nand U590 (N_590,In_447,In_2960);
and U591 (N_591,In_2190,In_2947);
or U592 (N_592,In_1518,In_481);
xor U593 (N_593,In_2392,In_651);
nand U594 (N_594,In_2451,In_1544);
and U595 (N_595,In_959,In_1199);
xor U596 (N_596,In_1335,In_2044);
and U597 (N_597,In_1487,In_670);
and U598 (N_598,In_1865,In_2985);
xor U599 (N_599,In_177,In_1290);
nand U600 (N_600,In_1305,In_2964);
nand U601 (N_601,In_1712,In_212);
and U602 (N_602,In_2120,In_1859);
nor U603 (N_603,In_364,In_795);
or U604 (N_604,In_2701,In_1511);
or U605 (N_605,In_294,In_2638);
or U606 (N_606,In_279,In_1262);
xor U607 (N_607,In_2694,In_1168);
nor U608 (N_608,In_2453,In_2907);
nor U609 (N_609,In_2136,In_1725);
or U610 (N_610,In_1137,In_799);
nand U611 (N_611,In_1632,In_1576);
and U612 (N_612,In_2829,In_812);
nor U613 (N_613,In_2060,In_2382);
and U614 (N_614,In_2939,In_2746);
or U615 (N_615,In_1599,In_1582);
nor U616 (N_616,In_1970,In_255);
or U617 (N_617,In_1026,In_2364);
and U618 (N_618,In_1195,In_1395);
nor U619 (N_619,In_1780,In_21);
xor U620 (N_620,In_780,In_1359);
or U621 (N_621,In_889,In_2514);
nand U622 (N_622,In_567,In_2440);
xnor U623 (N_623,In_486,In_1782);
and U624 (N_624,In_2111,In_427);
nor U625 (N_625,In_1454,In_2736);
and U626 (N_626,In_1375,In_1551);
and U627 (N_627,In_2354,In_2063);
nor U628 (N_628,In_2289,In_320);
nand U629 (N_629,In_1764,In_1361);
xor U630 (N_630,In_2621,In_477);
and U631 (N_631,In_1535,In_1474);
or U632 (N_632,In_1956,In_1005);
and U633 (N_633,In_2823,In_2137);
nor U634 (N_634,In_200,In_2802);
or U635 (N_635,In_327,In_1045);
nand U636 (N_636,In_1198,In_1299);
nor U637 (N_637,In_948,In_539);
xor U638 (N_638,In_1440,In_2885);
xnor U639 (N_639,In_963,In_668);
xnor U640 (N_640,In_413,In_1090);
nand U641 (N_641,In_961,In_1434);
and U642 (N_642,In_957,In_332);
xor U643 (N_643,In_538,In_2540);
nor U644 (N_644,In_2601,In_1430);
xor U645 (N_645,In_2863,In_69);
or U646 (N_646,In_239,In_1903);
nor U647 (N_647,In_2255,In_366);
and U648 (N_648,In_1485,In_2956);
nand U649 (N_649,In_2724,In_2626);
xnor U650 (N_650,In_671,In_787);
nand U651 (N_651,In_1283,In_821);
and U652 (N_652,In_2557,In_208);
or U653 (N_653,In_688,In_781);
xor U654 (N_654,In_1710,In_1012);
or U655 (N_655,In_667,In_2753);
and U656 (N_656,In_2266,In_1473);
nor U657 (N_657,In_2564,In_1886);
and U658 (N_658,In_1805,In_28);
and U659 (N_659,In_2505,In_560);
and U660 (N_660,In_2577,In_2086);
nor U661 (N_661,In_1093,In_2479);
and U662 (N_662,In_1769,In_1365);
xnor U663 (N_663,In_2876,In_1976);
and U664 (N_664,In_966,In_2844);
nor U665 (N_665,In_472,In_2276);
and U666 (N_666,In_1742,In_1033);
or U667 (N_667,In_1751,In_2366);
and U668 (N_668,In_838,In_229);
xor U669 (N_669,In_1016,In_1498);
and U670 (N_670,In_1960,In_710);
nor U671 (N_671,In_1311,In_561);
nor U672 (N_672,In_2998,In_613);
nand U673 (N_673,In_1999,In_217);
or U674 (N_674,In_432,In_27);
xnor U675 (N_675,In_1053,In_1813);
nand U676 (N_676,In_775,In_1786);
or U677 (N_677,In_2161,In_2094);
or U678 (N_678,In_2045,In_1930);
or U679 (N_679,In_2221,In_2954);
nand U680 (N_680,In_1907,In_2434);
nand U681 (N_681,In_2553,In_2103);
nor U682 (N_682,In_743,In_1328);
xnor U683 (N_683,In_1814,In_1214);
nor U684 (N_684,In_2666,In_584);
xnor U685 (N_685,In_1265,In_2776);
or U686 (N_686,In_316,In_1847);
or U687 (N_687,In_1927,In_926);
xor U688 (N_688,In_2204,In_1796);
and U689 (N_689,In_1488,In_1288);
or U690 (N_690,In_919,In_2561);
or U691 (N_691,In_2393,In_1509);
xor U692 (N_692,In_423,In_1252);
xor U693 (N_693,In_183,In_235);
nor U694 (N_694,In_282,In_2315);
nor U695 (N_695,In_2567,In_2987);
xor U696 (N_696,In_2234,In_1037);
nor U697 (N_697,In_2153,In_2313);
nor U698 (N_698,In_2551,In_2362);
or U699 (N_699,In_351,In_2133);
nand U700 (N_700,In_1420,In_2155);
nor U701 (N_701,In_62,In_1021);
xnor U702 (N_702,In_2810,In_2242);
nor U703 (N_703,In_603,In_877);
xnor U704 (N_704,In_1851,In_329);
and U705 (N_705,In_2879,In_295);
and U706 (N_706,In_2822,In_940);
or U707 (N_707,In_1954,In_408);
nor U708 (N_708,In_735,In_768);
and U709 (N_709,In_68,In_700);
nand U710 (N_710,In_2591,In_1386);
nand U711 (N_711,In_1408,In_2604);
xor U712 (N_712,In_2597,In_1910);
nor U713 (N_713,In_2417,In_2346);
or U714 (N_714,In_1470,In_434);
nor U715 (N_715,In_458,In_1715);
nor U716 (N_716,In_1389,In_1924);
nor U717 (N_717,In_263,In_75);
and U718 (N_718,In_2260,In_502);
and U719 (N_719,In_935,In_1263);
or U720 (N_720,In_1396,In_501);
nor U721 (N_721,In_833,In_823);
xnor U722 (N_722,In_2461,In_1402);
xor U723 (N_723,In_2899,In_2188);
nand U724 (N_724,In_1743,In_1167);
nand U725 (N_725,In_2302,In_2900);
nand U726 (N_726,In_450,In_2524);
or U727 (N_727,In_2388,In_1650);
or U728 (N_728,In_46,In_944);
nor U729 (N_729,In_232,In_1484);
nand U730 (N_730,In_694,In_2310);
and U731 (N_731,In_1948,In_1761);
and U732 (N_732,In_998,In_1555);
and U733 (N_733,In_283,In_1929);
or U734 (N_734,In_896,In_2959);
and U735 (N_735,In_1571,In_979);
and U736 (N_736,In_2341,In_1953);
or U737 (N_737,In_2709,In_2438);
xor U738 (N_738,In_1120,In_2493);
nor U739 (N_739,In_1893,In_2979);
xnor U740 (N_740,In_1058,In_1510);
nor U741 (N_741,In_1126,In_2509);
nor U742 (N_742,In_1945,In_57);
nor U743 (N_743,In_1882,In_1235);
or U744 (N_744,In_2535,In_1685);
and U745 (N_745,In_852,In_2348);
nand U746 (N_746,In_2600,In_1452);
nand U747 (N_747,In_1556,In_2731);
xor U748 (N_748,In_2184,In_1162);
nand U749 (N_749,In_2788,In_2054);
or U750 (N_750,In_779,In_1983);
nand U751 (N_751,In_1249,In_1091);
and U752 (N_752,In_2056,In_648);
or U753 (N_753,In_1878,In_1177);
nor U754 (N_754,In_2993,In_1221);
nor U755 (N_755,In_2467,In_1070);
nand U756 (N_756,In_1785,In_2331);
and U757 (N_757,In_99,In_1217);
nor U758 (N_758,In_2655,In_1294);
nor U759 (N_759,In_1332,In_2189);
nor U760 (N_760,In_711,In_752);
or U761 (N_761,In_299,In_2962);
nor U762 (N_762,In_2431,In_368);
nand U763 (N_763,In_2945,In_2469);
or U764 (N_764,In_2169,In_2430);
and U765 (N_765,In_2243,In_702);
xor U766 (N_766,In_938,In_2931);
or U767 (N_767,In_405,In_1810);
xor U768 (N_768,In_491,In_2207);
xnor U769 (N_769,In_70,In_1950);
or U770 (N_770,In_1081,In_1504);
nand U771 (N_771,In_1321,In_1445);
nor U772 (N_772,In_2784,In_627);
and U773 (N_773,In_2747,In_403);
nand U774 (N_774,In_2868,In_252);
or U775 (N_775,In_695,In_105);
nor U776 (N_776,In_2740,In_874);
nand U777 (N_777,In_497,In_1352);
and U778 (N_778,In_583,In_2756);
nand U779 (N_779,In_445,In_2446);
nand U780 (N_780,In_1465,In_1282);
xor U781 (N_781,In_2824,In_2213);
or U782 (N_782,In_414,In_214);
or U783 (N_783,In_2645,In_1730);
nor U784 (N_784,In_499,In_2757);
xnor U785 (N_785,In_1232,In_1560);
or U786 (N_786,In_2941,In_1203);
or U787 (N_787,In_2888,In_698);
and U788 (N_788,In_1367,In_1658);
or U789 (N_789,In_2413,In_2847);
xnor U790 (N_790,In_36,In_407);
and U791 (N_791,In_2818,In_444);
xnor U792 (N_792,In_1514,In_697);
nor U793 (N_793,In_1425,In_983);
xor U794 (N_794,In_2075,In_630);
nand U795 (N_795,In_2913,In_1490);
nand U796 (N_796,In_34,In_2930);
nor U797 (N_797,In_1307,In_2828);
nand U798 (N_798,In_1596,In_2880);
nor U799 (N_799,In_92,In_2441);
nand U800 (N_800,In_121,In_1852);
nor U801 (N_801,In_2228,In_164);
xnor U802 (N_802,In_1925,In_2678);
and U803 (N_803,In_809,In_595);
and U804 (N_804,In_1659,In_897);
and U805 (N_805,In_596,In_1651);
or U806 (N_806,In_1525,In_2754);
and U807 (N_807,In_1776,In_2218);
and U808 (N_808,In_1486,In_1673);
xnor U809 (N_809,In_1336,In_794);
or U810 (N_810,In_1547,In_2442);
xor U811 (N_811,In_202,In_834);
xnor U812 (N_812,In_1491,In_2676);
and U813 (N_813,In_573,In_547);
nor U814 (N_814,In_1967,In_643);
nor U815 (N_815,In_2725,In_733);
nor U816 (N_816,In_100,In_2566);
nand U817 (N_817,In_2065,In_1567);
or U818 (N_818,In_2734,In_1992);
or U819 (N_819,In_1548,In_2380);
nand U820 (N_820,In_1848,In_1429);
xor U821 (N_821,In_1968,In_1024);
nand U822 (N_822,In_1174,In_1912);
xnor U823 (N_823,In_1583,In_1543);
and U824 (N_824,In_1296,In_1552);
nor U825 (N_825,In_2774,In_2649);
xor U826 (N_826,In_127,In_1406);
nor U827 (N_827,In_228,In_1250);
nand U828 (N_828,In_1869,In_187);
or U829 (N_829,In_932,In_590);
nand U830 (N_830,In_1623,In_640);
and U831 (N_831,In_1362,In_1502);
nor U832 (N_832,In_22,In_1781);
nor U833 (N_833,In_1497,In_493);
and U834 (N_834,In_2273,In_2454);
or U835 (N_835,In_2465,In_1978);
or U836 (N_836,In_2820,In_1772);
and U837 (N_837,In_1285,In_2307);
nor U838 (N_838,In_958,In_680);
nor U839 (N_839,In_1433,In_2246);
nor U840 (N_840,In_2782,In_2644);
and U841 (N_841,In_642,In_352);
nor U842 (N_842,In_1492,In_2308);
or U843 (N_843,In_400,In_524);
nor U844 (N_844,In_162,In_1802);
nand U845 (N_845,In_2791,In_2955);
nor U846 (N_846,In_1724,In_2297);
or U847 (N_847,In_1236,In_2003);
nor U848 (N_848,In_2031,In_2200);
xor U849 (N_849,In_2288,In_2374);
or U850 (N_850,In_718,In_1403);
nor U851 (N_851,In_922,In_686);
nor U852 (N_852,In_1684,In_353);
xnor U853 (N_853,In_473,In_2099);
and U854 (N_854,In_1770,In_2968);
and U855 (N_855,In_585,In_734);
nand U856 (N_856,In_2780,In_1699);
and U857 (N_857,In_1046,In_1188);
nand U858 (N_858,In_2864,In_581);
or U859 (N_859,In_66,In_1411);
and U860 (N_860,In_2854,In_302);
or U861 (N_861,In_1397,In_2098);
nand U862 (N_862,In_967,In_300);
xnor U863 (N_863,In_1647,In_1993);
and U864 (N_864,In_2257,In_1691);
nand U865 (N_865,In_1390,In_223);
or U866 (N_866,In_453,In_192);
xnor U867 (N_867,In_2625,In_88);
and U868 (N_868,In_1029,In_274);
and U869 (N_869,In_2886,In_916);
or U870 (N_870,In_1371,In_1606);
nand U871 (N_871,In_749,In_1245);
or U872 (N_872,In_1347,In_2751);
nand U873 (N_873,In_1128,In_2657);
and U874 (N_874,In_424,In_398);
or U875 (N_875,In_33,In_2116);
nor U876 (N_876,In_534,In_2167);
and U877 (N_877,In_466,In_2020);
nor U878 (N_878,In_2195,In_1400);
nor U879 (N_879,In_650,In_1219);
and U880 (N_880,In_1047,In_2547);
or U881 (N_881,In_2541,In_2004);
or U882 (N_882,In_2398,In_2833);
and U883 (N_883,In_2492,In_995);
xnor U884 (N_884,In_336,In_1211);
or U885 (N_885,In_2117,In_243);
nor U886 (N_886,In_437,In_1979);
nand U887 (N_887,In_2855,In_2074);
xnor U888 (N_888,In_2490,In_854);
nor U889 (N_889,In_2660,In_246);
or U890 (N_890,In_637,In_862);
xnor U891 (N_891,In_2258,In_220);
nand U892 (N_892,In_701,In_256);
xnor U893 (N_893,In_531,In_1077);
xnor U894 (N_894,In_554,In_2647);
nand U895 (N_895,In_2122,In_1479);
and U896 (N_896,In_840,In_1085);
nand U897 (N_897,In_2141,In_2777);
and U898 (N_898,In_1541,In_856);
or U899 (N_899,In_2342,In_2176);
and U900 (N_900,In_1719,In_837);
nand U901 (N_901,In_1205,In_318);
xnor U902 (N_902,In_973,In_1904);
nand U903 (N_903,In_2683,In_1641);
xnor U904 (N_904,In_2949,In_904);
nand U905 (N_905,In_576,In_1405);
xor U906 (N_906,In_1315,In_1568);
nor U907 (N_907,In_1259,In_2634);
and U908 (N_908,In_2112,In_559);
nand U909 (N_909,In_2589,In_1530);
xnor U910 (N_910,In_2156,In_2896);
xor U911 (N_911,In_393,In_2211);
nor U912 (N_912,In_504,In_2744);
xor U913 (N_913,In_2922,In_1600);
or U914 (N_914,In_912,In_1178);
xor U915 (N_915,In_37,In_270);
nand U916 (N_916,In_2271,In_1334);
xor U917 (N_917,In_1722,In_1921);
or U918 (N_918,In_2580,In_1627);
nand U919 (N_919,In_617,In_1597);
or U920 (N_920,In_1224,In_699);
or U921 (N_921,In_872,In_1039);
xor U922 (N_922,In_1034,In_435);
nand U923 (N_923,In_628,In_2272);
or U924 (N_924,In_1301,In_1789);
xor U925 (N_925,In_2938,In_1545);
and U926 (N_926,In_1832,In_474);
nand U927 (N_927,In_1398,In_1698);
nor U928 (N_928,In_2851,In_2095);
nor U929 (N_929,In_1451,In_1522);
xnor U930 (N_930,In_2881,In_2106);
nor U931 (N_931,In_2973,In_1156);
nand U932 (N_932,In_2646,In_1837);
or U933 (N_933,In_858,In_1247);
nand U934 (N_934,In_1327,In_543);
nor U935 (N_935,In_740,In_1022);
xnor U936 (N_936,In_2556,In_1989);
and U937 (N_937,In_1577,In_1537);
or U938 (N_938,In_2867,In_2036);
xnor U939 (N_939,In_376,In_2813);
nor U940 (N_940,In_2745,In_1652);
nor U941 (N_941,In_5,In_288);
xor U942 (N_942,In_113,In_766);
nand U943 (N_943,In_190,In_1258);
nand U944 (N_944,In_608,In_240);
xnor U945 (N_945,In_677,In_1496);
or U946 (N_946,In_2568,In_106);
or U947 (N_947,In_2385,In_1380);
nand U948 (N_948,In_1208,In_855);
nand U949 (N_949,In_349,In_1152);
nor U950 (N_950,In_532,In_2712);
nor U951 (N_951,In_1257,In_1888);
nand U952 (N_952,In_866,In_2030);
nor U953 (N_953,In_2786,In_741);
xnor U954 (N_954,In_1867,In_355);
and U955 (N_955,In_1720,In_1703);
or U956 (N_956,In_416,In_1364);
xor U957 (N_957,In_2612,In_213);
xor U958 (N_958,In_2838,In_953);
nand U959 (N_959,In_1412,In_380);
or U960 (N_960,In_2748,In_1108);
and U961 (N_961,In_103,In_730);
and U962 (N_962,In_173,In_593);
and U963 (N_963,In_1794,In_2895);
nor U964 (N_964,In_1220,In_1920);
xor U965 (N_965,In_2082,In_784);
nor U966 (N_966,In_2806,In_903);
and U967 (N_967,In_1777,In_594);
or U968 (N_968,In_1383,In_120);
nand U969 (N_969,In_564,In_324);
nand U970 (N_970,In_1139,In_1889);
or U971 (N_971,In_1686,In_851);
xnor U972 (N_972,In_119,In_2335);
or U973 (N_973,In_2059,In_133);
xnor U974 (N_974,In_2261,In_598);
or U975 (N_975,In_1210,In_1399);
nor U976 (N_976,In_1996,In_1682);
nand U977 (N_977,In_30,In_222);
xnor U978 (N_978,In_460,In_1342);
or U979 (N_979,In_505,In_828);
or U980 (N_980,In_2699,In_2722);
nor U981 (N_981,In_989,In_1744);
xor U982 (N_982,In_1988,In_1590);
xor U983 (N_983,In_1003,In_1922);
and U984 (N_984,In_2411,In_2019);
and U985 (N_985,In_1812,In_1409);
nand U986 (N_986,In_822,In_1073);
xor U987 (N_987,In_2071,In_1883);
xnor U988 (N_988,In_861,In_2539);
nand U989 (N_989,In_1314,In_1612);
nand U990 (N_990,In_2607,In_1478);
and U991 (N_991,In_2073,In_429);
nand U992 (N_992,In_1680,In_550);
or U993 (N_993,In_2402,In_1819);
nor U994 (N_994,In_1083,In_1481);
nand U995 (N_995,In_1702,In_461);
or U996 (N_996,In_1040,In_704);
and U997 (N_997,In_1943,In_663);
nor U998 (N_998,In_885,In_154);
nor U999 (N_999,In_2691,In_2682);
xor U1000 (N_1000,In_412,In_1150);
and U1001 (N_1001,In_1495,In_2795);
xor U1002 (N_1002,In_800,In_1513);
nand U1003 (N_1003,In_1601,In_114);
nor U1004 (N_1004,In_572,In_363);
nor U1005 (N_1005,In_2594,In_1302);
and U1006 (N_1006,In_1151,In_2531);
nor U1007 (N_1007,In_2654,In_2148);
or U1008 (N_1008,In_936,In_1818);
xor U1009 (N_1009,In_2,In_2077);
nand U1010 (N_1010,In_927,In_2921);
nand U1011 (N_1011,In_2129,In_58);
and U1012 (N_1012,In_1110,In_2732);
nor U1013 (N_1013,In_900,In_2299);
and U1014 (N_1014,In_1275,In_125);
nor U1015 (N_1015,In_1443,In_1172);
and U1016 (N_1016,In_2347,In_254);
or U1017 (N_1017,In_2421,In_2384);
and U1018 (N_1018,In_1896,In_816);
nand U1019 (N_1019,In_507,In_1253);
and U1020 (N_1020,In_2670,In_1276);
nor U1021 (N_1021,In_135,In_2217);
nand U1022 (N_1022,In_186,In_2317);
nand U1023 (N_1023,In_2484,In_495);
xor U1024 (N_1024,In_1866,In_2807);
and U1025 (N_1025,In_2147,In_2383);
xor U1026 (N_1026,In_0,In_990);
nand U1027 (N_1027,In_1388,In_1687);
and U1028 (N_1028,In_2903,In_2989);
or U1029 (N_1029,In_2047,In_1639);
and U1030 (N_1030,In_2233,In_1791);
and U1031 (N_1031,In_638,In_1354);
or U1032 (N_1032,In_1718,In_2994);
or U1033 (N_1033,In_179,In_462);
nor U1034 (N_1034,In_2651,In_545);
and U1035 (N_1035,In_479,In_847);
or U1036 (N_1036,In_2808,In_1385);
xor U1037 (N_1037,In_939,In_304);
xor U1038 (N_1038,In_210,In_2162);
and U1039 (N_1039,In_994,In_2915);
nand U1040 (N_1040,In_974,In_789);
xnor U1041 (N_1041,In_1101,In_2274);
nand U1042 (N_1042,In_2033,In_67);
xor U1043 (N_1043,In_1407,In_2485);
nand U1044 (N_1044,In_758,In_1701);
nor U1045 (N_1045,In_669,In_514);
or U1046 (N_1046,In_1180,In_2456);
nor U1047 (N_1047,In_2668,In_130);
nor U1048 (N_1048,In_2102,In_681);
or U1049 (N_1049,In_1119,In_1494);
and U1050 (N_1050,In_1078,In_2367);
nor U1051 (N_1051,In_1971,In_1816);
xnor U1052 (N_1052,In_2982,In_388);
nor U1053 (N_1053,In_40,In_914);
nand U1054 (N_1054,In_2814,In_2662);
nand U1055 (N_1055,In_2066,In_1227);
nand U1056 (N_1056,In_1049,In_19);
nor U1057 (N_1057,In_2068,In_161);
xor U1058 (N_1058,In_201,In_891);
or U1059 (N_1059,In_2536,In_2433);
nor U1060 (N_1060,In_678,In_886);
or U1061 (N_1061,In_2873,In_850);
or U1062 (N_1062,In_1803,In_1020);
and U1063 (N_1063,In_1823,In_63);
nand U1064 (N_1064,In_1231,In_1771);
xor U1065 (N_1065,In_1947,In_2223);
nor U1066 (N_1066,In_2230,In_2305);
nor U1067 (N_1067,In_2113,In_2439);
xnor U1068 (N_1068,In_1345,In_563);
or U1069 (N_1069,In_530,In_331);
and U1070 (N_1070,In_420,In_2574);
nor U1071 (N_1071,In_2619,In_2287);
nor U1072 (N_1072,In_1300,In_1442);
nor U1073 (N_1073,In_2080,In_819);
and U1074 (N_1074,In_1427,In_1563);
nand U1075 (N_1075,In_788,In_317);
nor U1076 (N_1076,In_286,In_2995);
nand U1077 (N_1077,In_1909,In_2559);
and U1078 (N_1078,In_985,In_2883);
nor U1079 (N_1079,In_895,In_2592);
and U1080 (N_1080,In_2901,In_155);
and U1081 (N_1081,In_1007,In_2761);
xnor U1082 (N_1082,In_1341,In_2690);
xor U1083 (N_1083,In_2201,In_2532);
and U1084 (N_1084,In_2475,In_1075);
and U1085 (N_1085,In_1458,In_1516);
nand U1086 (N_1086,In_1637,In_1455);
xor U1087 (N_1087,In_542,In_1959);
and U1088 (N_1088,In_26,In_2529);
nor U1089 (N_1089,In_930,In_2043);
nor U1090 (N_1090,In_656,In_278);
xnor U1091 (N_1091,In_227,In_2119);
or U1092 (N_1092,In_358,In_1068);
nor U1093 (N_1093,In_1014,In_2226);
and U1094 (N_1094,In_1351,In_489);
xnor U1095 (N_1095,In_2695,In_2884);
xor U1096 (N_1096,In_933,In_1369);
xor U1097 (N_1097,In_2444,In_605);
or U1098 (N_1098,In_2432,In_2400);
nor U1099 (N_1099,In_1340,In_2292);
xnor U1100 (N_1100,In_529,In_315);
nand U1101 (N_1101,In_1467,In_174);
or U1102 (N_1102,In_1853,In_1241);
xnor U1103 (N_1103,In_1877,In_1461);
xor U1104 (N_1104,In_150,In_2538);
nand U1105 (N_1105,In_987,In_2714);
xor U1106 (N_1106,In_2550,In_1117);
xnor U1107 (N_1107,In_1845,In_2491);
xor U1108 (N_1108,In_485,In_1426);
nor U1109 (N_1109,In_1735,In_90);
nand U1110 (N_1110,In_1621,In_348);
and U1111 (N_1111,In_1890,In_719);
or U1112 (N_1112,In_182,In_2680);
nand U1113 (N_1113,In_2488,In_606);
and U1114 (N_1114,In_864,In_2827);
nor U1115 (N_1115,In_1871,In_1230);
nor U1116 (N_1116,In_2235,In_1421);
nand U1117 (N_1117,In_1457,In_1714);
and U1118 (N_1118,In_1103,In_2743);
nand U1119 (N_1119,In_386,In_1273);
or U1120 (N_1120,In_7,In_1324);
or U1121 (N_1121,In_1919,In_992);
or U1122 (N_1122,In_575,In_2503);
or U1123 (N_1123,In_1456,In_2352);
and U1124 (N_1124,In_1270,In_2799);
nor U1125 (N_1125,In_685,In_1157);
nand U1126 (N_1126,In_1700,In_2773);
xor U1127 (N_1127,In_1462,In_411);
nor U1128 (N_1128,In_814,In_131);
and U1129 (N_1129,In_2720,In_1765);
nand U1130 (N_1130,In_1648,In_1194);
nor U1131 (N_1131,In_604,In_1713);
nand U1132 (N_1132,In_1105,In_1088);
and U1133 (N_1133,In_2058,In_980);
nand U1134 (N_1134,In_728,In_2280);
nor U1135 (N_1135,In_2143,In_373);
nand U1136 (N_1136,In_124,In_1935);
or U1137 (N_1137,In_859,In_1622);
or U1138 (N_1138,In_1533,In_2537);
or U1139 (N_1139,In_118,In_1523);
or U1140 (N_1140,In_2253,In_1873);
or U1141 (N_1141,In_1384,In_2418);
nor U1142 (N_1142,In_1374,In_2617);
or U1143 (N_1143,In_2933,In_2849);
or U1144 (N_1144,In_1628,In_1528);
or U1145 (N_1145,In_1588,In_2801);
and U1146 (N_1146,In_2363,In_621);
nand U1147 (N_1147,In_2387,In_421);
xnor U1148 (N_1148,In_1381,In_148);
nor U1149 (N_1149,In_2588,In_978);
xor U1150 (N_1150,In_1145,In_2076);
nand U1151 (N_1151,In_2355,In_659);
xor U1152 (N_1152,In_2338,In_1009);
nor U1153 (N_1153,In_836,In_2323);
xnor U1154 (N_1154,In_151,In_568);
nand U1155 (N_1155,In_1450,In_2007);
or U1156 (N_1156,In_488,In_760);
nor U1157 (N_1157,In_1916,In_78);
or U1158 (N_1158,In_756,In_578);
xor U1159 (N_1159,In_157,In_2735);
and U1160 (N_1160,In_1581,In_494);
or U1161 (N_1161,In_2920,In_551);
or U1162 (N_1162,In_876,In_2423);
and U1163 (N_1163,In_2560,In_2369);
nor U1164 (N_1164,In_1200,In_1121);
xor U1165 (N_1165,In_483,In_2250);
nand U1166 (N_1166,In_2192,In_1318);
nand U1167 (N_1167,In_2090,In_722);
and U1168 (N_1168,In_2191,In_1558);
nand U1169 (N_1169,In_6,In_1874);
nor U1170 (N_1170,In_129,In_1289);
nor U1171 (N_1171,In_1880,In_1122);
nand U1172 (N_1172,In_1645,In_80);
xnor U1173 (N_1173,In_2513,In_649);
nor U1174 (N_1174,In_43,In_1982);
nor U1175 (N_1175,In_654,In_2905);
nand U1176 (N_1176,In_1831,In_2894);
or U1177 (N_1177,In_2798,In_2659);
nand U1178 (N_1178,In_1668,In_982);
or U1179 (N_1179,In_1584,In_29);
nor U1180 (N_1180,In_175,In_1729);
or U1181 (N_1181,In_1448,In_2145);
xor U1182 (N_1182,In_2286,In_225);
xnor U1183 (N_1183,In_1531,In_679);
and U1184 (N_1184,In_586,In_2521);
xor U1185 (N_1185,In_2545,In_1856);
xor U1186 (N_1186,In_146,In_1357);
nor U1187 (N_1187,In_2800,In_2511);
nand U1188 (N_1188,In_533,In_8);
and U1189 (N_1189,In_882,In_1414);
nand U1190 (N_1190,In_2351,In_860);
or U1191 (N_1191,In_2840,In_45);
nand U1192 (N_1192,In_1323,In_53);
xnor U1193 (N_1193,In_284,In_1060);
or U1194 (N_1194,In_2809,In_482);
nand U1195 (N_1195,In_1272,In_1917);
and U1196 (N_1196,In_1529,In_2770);
or U1197 (N_1197,In_2582,In_1585);
and U1198 (N_1198,In_2693,In_857);
nand U1199 (N_1199,In_73,In_1377);
xor U1200 (N_1200,N_252,N_755);
xnor U1201 (N_1201,In_1538,In_1373);
and U1202 (N_1202,In_774,N_345);
xor U1203 (N_1203,N_277,N_1084);
or U1204 (N_1204,In_2552,In_2674);
or U1205 (N_1205,N_552,N_975);
nand U1206 (N_1206,N_0,N_511);
nand U1207 (N_1207,In_1056,In_614);
or U1208 (N_1208,N_1195,N_709);
and U1209 (N_1209,N_713,N_1087);
nand U1210 (N_1210,In_1694,N_522);
xor U1211 (N_1211,N_65,In_1281);
xor U1212 (N_1212,In_2565,N_166);
xor U1213 (N_1213,N_331,N_309);
or U1214 (N_1214,N_390,N_1096);
or U1215 (N_1215,In_140,In_439);
xnor U1216 (N_1216,N_574,N_1061);
or U1217 (N_1217,In_588,N_292);
and U1218 (N_1218,In_972,N_834);
nor U1219 (N_1219,N_199,In_2804);
nand U1220 (N_1220,N_391,In_321);
nor U1221 (N_1221,In_634,N_447);
xor U1222 (N_1222,N_1022,In_404);
nor U1223 (N_1223,N_1005,N_669);
nor U1224 (N_1224,N_649,In_1766);
nor U1225 (N_1225,In_2329,N_61);
nor U1226 (N_1226,In_748,N_978);
and U1227 (N_1227,N_236,N_386);
nand U1228 (N_1228,N_139,In_579);
or U1229 (N_1229,N_1138,N_628);
xnor U1230 (N_1230,In_2414,In_356);
xnor U1231 (N_1231,N_16,N_733);
and U1232 (N_1232,In_2334,In_2023);
nand U1233 (N_1233,N_756,In_1844);
xnor U1234 (N_1234,N_561,N_357);
and U1235 (N_1235,In_1080,N_637);
or U1236 (N_1236,In_1229,In_449);
and U1237 (N_1237,In_2605,N_7);
nor U1238 (N_1238,In_2544,N_488);
nand U1239 (N_1239,N_544,N_182);
and U1240 (N_1240,In_2610,N_1183);
nand U1241 (N_1241,N_141,In_2322);
nand U1242 (N_1242,N_39,N_1120);
xor U1243 (N_1243,N_428,N_845);
and U1244 (N_1244,N_494,N_170);
xnor U1245 (N_1245,In_15,In_993);
and U1246 (N_1246,In_2006,N_722);
and U1247 (N_1247,N_749,N_346);
and U1248 (N_1248,N_71,N_738);
xnor U1249 (N_1249,N_777,N_186);
or U1250 (N_1250,N_1107,N_928);
nand U1251 (N_1251,N_870,In_419);
and U1252 (N_1252,In_2282,N_576);
or U1253 (N_1253,N_250,N_740);
or U1254 (N_1254,N_1086,In_1222);
and U1255 (N_1255,N_1071,N_360);
or U1256 (N_1256,In_2980,In_1517);
or U1257 (N_1257,In_625,In_1740);
xnor U1258 (N_1258,N_44,N_772);
nand U1259 (N_1259,N_272,In_2579);
xor U1260 (N_1260,N_460,In_2997);
or U1261 (N_1261,In_112,N_130);
or U1262 (N_1262,N_314,N_138);
xor U1263 (N_1263,N_1033,N_508);
or U1264 (N_1264,In_1052,In_277);
nor U1265 (N_1265,N_418,N_680);
xnor U1266 (N_1266,N_609,N_339);
or U1267 (N_1267,In_1500,N_22);
nor U1268 (N_1268,N_643,N_438);
or U1269 (N_1269,N_481,N_618);
xnor U1270 (N_1270,N_1032,N_446);
xor U1271 (N_1271,N_773,In_2115);
and U1272 (N_1272,N_1035,N_6);
nand U1273 (N_1273,In_1030,In_168);
nor U1274 (N_1274,N_249,In_609);
nand U1275 (N_1275,N_90,N_49);
nand U1276 (N_1276,N_915,N_316);
nand U1277 (N_1277,N_783,N_932);
or U1278 (N_1278,In_1728,N_686);
nor U1279 (N_1279,N_1063,In_2639);
or U1280 (N_1280,In_1690,N_864);
and U1281 (N_1281,N_736,In_2035);
xnor U1282 (N_1282,N_1129,N_203);
or U1283 (N_1283,N_1025,N_681);
and U1284 (N_1284,N_568,N_1147);
and U1285 (N_1285,N_626,N_290);
nand U1286 (N_1286,N_601,N_958);
nor U1287 (N_1287,In_1134,In_138);
nand U1288 (N_1288,N_999,In_268);
xor U1289 (N_1289,In_1004,N_1165);
nand U1290 (N_1290,N_638,In_924);
and U1291 (N_1291,In_2034,In_616);
and U1292 (N_1292,In_1561,N_468);
or U1293 (N_1293,In_2759,In_1875);
or U1294 (N_1294,N_879,In_1255);
and U1295 (N_1295,N_82,N_1046);
and U1296 (N_1296,N_383,In_471);
nand U1297 (N_1297,In_2906,N_429);
or U1298 (N_1298,N_745,N_885);
xor U1299 (N_1299,In_2370,N_1090);
nor U1300 (N_1300,N_746,In_2447);
nor U1301 (N_1301,N_704,N_1113);
nor U1302 (N_1302,N_714,N_1122);
or U1303 (N_1303,In_1313,In_1732);
and U1304 (N_1304,In_1181,N_35);
or U1305 (N_1305,In_2375,In_713);
nand U1306 (N_1306,N_367,N_225);
and U1307 (N_1307,N_105,In_1980);
and U1308 (N_1308,N_324,N_930);
nor U1309 (N_1309,N_925,N_1148);
nor U1310 (N_1310,N_92,N_695);
xor U1311 (N_1311,N_153,N_821);
nor U1312 (N_1312,In_410,In_1675);
nor U1313 (N_1313,In_2121,N_959);
xnor U1314 (N_1314,N_943,N_903);
nand U1315 (N_1315,In_2395,N_1196);
or U1316 (N_1316,In_1246,In_1898);
xor U1317 (N_1317,N_434,N_102);
or U1318 (N_1318,N_707,In_143);
and U1319 (N_1319,N_155,In_526);
nor U1320 (N_1320,N_780,N_115);
or U1321 (N_1321,N_439,In_792);
or U1322 (N_1322,N_1187,N_758);
and U1323 (N_1323,N_883,In_906);
xor U1324 (N_1324,N_1164,In_2633);
or U1325 (N_1325,N_227,N_216);
nand U1326 (N_1326,N_1002,In_1264);
xor U1327 (N_1327,N_207,N_335);
or U1328 (N_1328,In_2501,In_589);
nor U1329 (N_1329,N_392,In_2602);
or U1330 (N_1330,N_644,N_763);
or U1331 (N_1331,N_828,In_570);
xnor U1332 (N_1332,N_156,N_567);
and U1333 (N_1333,In_1955,In_1476);
xnor U1334 (N_1334,N_135,In_156);
and U1335 (N_1335,In_1363,In_2405);
and U1336 (N_1336,In_1271,In_2707);
xnor U1337 (N_1337,N_600,N_238);
nor U1338 (N_1338,In_74,N_317);
nor U1339 (N_1339,N_310,N_769);
or U1340 (N_1340,In_1838,N_807);
or U1341 (N_1341,N_245,N_363);
and U1342 (N_1342,In_2596,N_1112);
or U1343 (N_1343,N_161,In_1572);
nor U1344 (N_1344,N_848,N_151);
and U1345 (N_1345,In_96,N_829);
or U1346 (N_1346,N_913,In_145);
xnor U1347 (N_1347,In_1431,N_856);
nand U1348 (N_1348,N_952,N_1082);
or U1349 (N_1349,N_858,In_2911);
or U1350 (N_1350,In_338,In_244);
nor U1351 (N_1351,N_779,N_716);
nand U1352 (N_1352,In_2410,N_122);
nor U1353 (N_1353,N_241,N_584);
or U1354 (N_1354,In_2996,N_406);
nor U1355 (N_1355,N_825,N_1034);
nor U1356 (N_1356,N_657,In_2999);
and U1357 (N_1357,N_688,In_703);
xor U1358 (N_1358,N_334,N_1198);
nand U1359 (N_1359,N_661,N_1054);
nand U1360 (N_1360,N_876,In_1678);
and U1361 (N_1361,In_463,In_1739);
nor U1362 (N_1362,In_2050,N_771);
xor U1363 (N_1363,N_374,N_1101);
and U1364 (N_1364,In_2958,N_352);
xnor U1365 (N_1365,In_1261,N_937);
or U1366 (N_1366,N_405,In_2360);
or U1367 (N_1367,N_815,In_1173);
nand U1368 (N_1368,N_486,N_631);
nand U1369 (N_1369,In_2181,N_178);
nor U1370 (N_1370,N_776,N_853);
and U1371 (N_1371,N_1114,N_942);
nand U1372 (N_1372,N_653,In_1065);
or U1373 (N_1373,N_1173,N_1030);
nor U1374 (N_1374,N_860,N_775);
nand U1375 (N_1375,N_372,N_427);
or U1376 (N_1376,N_899,N_977);
xor U1377 (N_1377,In_1002,N_1099);
and U1378 (N_1378,N_946,N_315);
xnor U1379 (N_1379,N_974,N_531);
or U1380 (N_1380,In_2787,In_887);
and U1381 (N_1381,In_762,N_817);
and U1382 (N_1382,N_844,N_359);
nand U1383 (N_1383,N_366,N_1186);
xor U1384 (N_1384,N_530,In_1023);
nor U1385 (N_1385,N_757,N_254);
or U1386 (N_1386,N_45,In_38);
xnor U1387 (N_1387,N_332,N_307);
and U1388 (N_1388,N_800,N_1003);
and U1389 (N_1389,In_1969,In_592);
nand U1390 (N_1390,In_341,In_267);
nand U1391 (N_1391,N_1057,N_691);
xor U1392 (N_1392,N_191,N_291);
nand U1393 (N_1393,In_915,N_927);
xor U1394 (N_1394,N_752,In_1564);
nand U1395 (N_1395,In_2839,N_251);
or U1396 (N_1396,N_1007,N_1125);
nor U1397 (N_1397,N_276,N_298);
and U1398 (N_1398,In_976,N_514);
and U1399 (N_1399,N_562,N_452);
xnor U1400 (N_1400,N_991,N_791);
nor U1401 (N_1401,N_774,N_751);
nand U1402 (N_1402,N_673,N_666);
or U1403 (N_1403,N_179,N_420);
or U1404 (N_1404,N_503,N_833);
nor U1405 (N_1405,N_902,N_55);
xor U1406 (N_1406,N_53,In_845);
xnor U1407 (N_1407,N_444,N_1080);
nand U1408 (N_1408,N_350,In_1653);
or U1409 (N_1409,In_311,In_1546);
nand U1410 (N_1410,N_424,In_230);
or U1411 (N_1411,N_694,N_58);
nor U1412 (N_1412,N_555,In_2981);
nand U1413 (N_1413,In_1619,In_2320);
nand U1414 (N_1414,In_2283,In_454);
nor U1415 (N_1415,In_521,In_1404);
and U1416 (N_1416,N_811,N_563);
and U1417 (N_1417,In_265,In_2325);
and U1418 (N_1418,In_1256,In_2758);
nor U1419 (N_1419,In_1010,N_13);
nand U1420 (N_1420,N_1006,In_2139);
or U1421 (N_1421,In_176,In_2072);
xor U1422 (N_1422,In_2733,N_954);
and U1423 (N_1423,In_2944,In_2214);
and U1424 (N_1424,In_2572,In_2303);
nor U1425 (N_1425,N_767,N_1036);
or U1426 (N_1426,In_1142,In_1308);
nand U1427 (N_1427,In_2048,N_608);
nor U1428 (N_1428,In_1633,N_957);
and U1429 (N_1429,N_641,In_2489);
nand U1430 (N_1430,N_95,N_702);
and U1431 (N_1431,N_548,In_1423);
nand U1432 (N_1432,N_177,N_900);
xnor U1433 (N_1433,In_566,N_893);
and U1434 (N_1434,N_1169,N_847);
or U1435 (N_1435,N_96,In_2445);
nand U1436 (N_1436,N_24,N_449);
and U1437 (N_1437,N_577,N_1176);
or U1438 (N_1438,In_511,N_229);
or U1439 (N_1439,N_586,N_857);
nor U1440 (N_1440,N_539,N_454);
nor U1441 (N_1441,In_1202,N_998);
nor U1442 (N_1442,N_659,In_1278);
or U1443 (N_1443,N_518,N_152);
xnor U1444 (N_1444,In_536,N_1104);
and U1445 (N_1445,N_613,In_965);
nor U1446 (N_1446,N_86,N_1041);
or U1447 (N_1447,In_2301,N_1060);
nand U1448 (N_1448,N_253,In_1132);
nand U1449 (N_1449,N_29,N_540);
nor U1450 (N_1450,N_483,N_676);
or U1451 (N_1451,N_1143,In_2268);
xor U1452 (N_1452,N_21,In_2015);
xor U1453 (N_1453,In_2525,In_1608);
nand U1454 (N_1454,In_2927,N_570);
xor U1455 (N_1455,N_737,In_2935);
and U1456 (N_1456,In_2285,N_950);
nor U1457 (N_1457,N_840,N_934);
or U1458 (N_1458,N_81,N_408);
and U1459 (N_1459,N_1188,N_689);
and U1460 (N_1460,N_1159,N_510);
nand U1461 (N_1461,In_1696,N_73);
xor U1462 (N_1462,In_732,N_1121);
nor U1463 (N_1463,N_700,In_1444);
xnor U1464 (N_1464,N_128,N_57);
xnor U1465 (N_1465,N_851,In_2179);
nand U1466 (N_1466,N_967,N_917);
xnor U1467 (N_1467,In_2792,N_108);
xnor U1468 (N_1468,In_2658,N_545);
nand U1469 (N_1469,In_77,N_687);
and U1470 (N_1470,In_2412,In_772);
or U1471 (N_1471,N_287,In_1974);
or U1472 (N_1472,In_2389,In_2878);
nand U1473 (N_1473,N_515,N_134);
nand U1474 (N_1474,In_813,In_1187);
nand U1475 (N_1475,N_892,N_764);
and U1476 (N_1476,In_1938,In_1153);
or U1477 (N_1477,N_476,N_1156);
or U1478 (N_1478,N_1042,N_46);
nand U1479 (N_1479,In_807,In_1689);
nor U1480 (N_1480,In_946,N_489);
and U1481 (N_1481,In_153,N_595);
or U1482 (N_1482,N_364,In_2706);
or U1483 (N_1483,N_1052,In_921);
nor U1484 (N_1484,N_770,In_2312);
or U1485 (N_1485,N_672,In_2611);
xnor U1486 (N_1486,N_1167,N_538);
nand U1487 (N_1487,In_971,In_2406);
nor U1488 (N_1488,N_635,In_1795);
and U1489 (N_1489,In_2549,N_417);
or U1490 (N_1490,N_517,N_1043);
nand U1491 (N_1491,In_1891,In_1337);
or U1492 (N_1492,In_2064,In_848);
and U1493 (N_1493,N_131,In_751);
xnor U1494 (N_1494,In_2265,In_791);
nand U1495 (N_1495,N_744,In_986);
nor U1496 (N_1496,N_465,N_1181);
and U1497 (N_1497,N_349,N_875);
nor U1498 (N_1498,N_910,In_2825);
xnor U1499 (N_1499,N_665,In_1644);
or U1500 (N_1500,N_206,In_218);
xnor U1501 (N_1501,N_159,In_555);
nor U1502 (N_1502,In_1578,In_1708);
and U1503 (N_1503,N_243,In_1681);
nor U1504 (N_1504,N_432,N_690);
nor U1505 (N_1505,N_50,N_228);
or U1506 (N_1506,N_217,In_1657);
xnor U1507 (N_1507,In_2587,N_924);
and U1508 (N_1508,In_2089,N_861);
or U1509 (N_1509,N_968,In_2730);
nand U1510 (N_1510,N_34,In_1923);
nor U1511 (N_1511,N_981,In_2904);
nand U1512 (N_1512,N_1023,N_1047);
nor U1513 (N_1513,N_36,N_490);
nor U1514 (N_1514,N_1026,N_378);
xnor U1515 (N_1515,N_1027,N_841);
xnor U1516 (N_1516,N_1185,N_569);
nor U1517 (N_1517,N_533,N_306);
and U1518 (N_1518,N_933,N_72);
nor U1519 (N_1519,In_1665,N_461);
nor U1520 (N_1520,N_822,N_1108);
or U1521 (N_1521,N_97,N_380);
or U1522 (N_1522,N_940,N_1175);
and U1523 (N_1523,N_327,In_2051);
nor U1524 (N_1524,N_622,In_2460);
xor U1525 (N_1525,In_1902,In_910);
nor U1526 (N_1526,N_121,N_1139);
and U1527 (N_1527,N_127,N_99);
and U1528 (N_1528,N_919,N_886);
xnor U1529 (N_1529,N_308,N_399);
xor U1530 (N_1530,In_198,N_341);
nand U1531 (N_1531,N_1127,N_321);
nor U1532 (N_1532,N_565,N_914);
or U1533 (N_1533,N_835,In_18);
and U1534 (N_1534,In_1438,N_1008);
nor U1535 (N_1535,In_1089,N_1123);
nand U1536 (N_1536,In_657,N_765);
nand U1537 (N_1537,N_759,N_69);
nor U1538 (N_1538,N_467,N_302);
nor U1539 (N_1539,N_469,N_869);
or U1540 (N_1540,N_430,In_865);
or U1541 (N_1541,In_917,In_395);
nor U1542 (N_1542,N_1110,N_278);
or U1543 (N_1543,N_788,N_1150);
or U1544 (N_1544,In_587,N_581);
and U1545 (N_1545,N_9,N_20);
nor U1546 (N_1546,In_163,In_2972);
xor U1547 (N_1547,N_31,N_1095);
nor U1548 (N_1548,In_1977,N_411);
nand U1549 (N_1549,In_2027,N_660);
nand U1550 (N_1550,N_648,In_2487);
and U1551 (N_1551,N_630,In_2950);
nand U1552 (N_1552,N_168,In_1994);
and U1553 (N_1553,N_263,N_557);
nand U1554 (N_1554,In_2943,In_2158);
xnor U1555 (N_1555,N_148,N_623);
or U1556 (N_1556,N_655,In_1251);
or U1557 (N_1557,N_1031,In_2507);
nor U1558 (N_1558,In_1998,In_2924);
or U1559 (N_1559,N_333,N_1157);
or U1560 (N_1560,In_1109,N_247);
nor U1561 (N_1561,N_423,N_931);
nand U1562 (N_1562,N_84,N_664);
or U1563 (N_1563,In_1750,In_611);
nor U1564 (N_1564,N_393,In_2482);
xor U1565 (N_1565,N_342,In_1370);
nand U1566 (N_1566,N_652,In_908);
or U1567 (N_1567,N_1166,In_1931);
xnor U1568 (N_1568,N_389,N_564);
nand U1569 (N_1569,In_1393,N_1055);
xor U1570 (N_1570,In_2717,N_859);
xnor U1571 (N_1571,N_492,N_246);
and U1572 (N_1572,In_1850,N_204);
nand U1573 (N_1573,In_1662,In_205);
or U1574 (N_1574,In_949,In_2969);
and U1575 (N_1575,N_442,N_1013);
nor U1576 (N_1576,In_1958,In_16);
and U1577 (N_1577,N_270,In_1565);
xnor U1578 (N_1578,N_507,In_1757);
nor U1579 (N_1579,N_224,N_962);
nor U1580 (N_1580,N_210,In_1617);
and U1581 (N_1581,N_541,In_391);
nand U1582 (N_1582,N_375,In_873);
nor U1583 (N_1583,N_180,In_2515);
xor U1584 (N_1584,N_656,N_677);
and U1585 (N_1585,N_602,In_2420);
or U1586 (N_1586,N_1168,In_2298);
nand U1587 (N_1587,N_258,In_2686);
and U1588 (N_1588,N_909,In_771);
nor U1589 (N_1589,In_181,N_257);
nand U1590 (N_1590,N_760,N_1197);
nand U1591 (N_1591,N_698,In_169);
nor U1592 (N_1592,N_136,In_1171);
xnor U1593 (N_1593,In_343,In_2009);
and U1594 (N_1594,N_794,N_710);
xor U1595 (N_1595,N_582,N_878);
nand U1596 (N_1596,N_318,N_1155);
xnor U1597 (N_1597,N_929,In_1501);
nor U1598 (N_1598,N_304,In_397);
nand U1599 (N_1599,N_175,In_1748);
and U1600 (N_1600,In_1240,N_521);
nand U1601 (N_1601,N_158,N_262);
or U1602 (N_1602,N_674,N_201);
or U1603 (N_1603,N_734,N_273);
and U1604 (N_1604,N_523,In_2365);
xor U1605 (N_1605,N_213,N_1044);
or U1606 (N_1606,N_1058,In_2554);
xnor U1607 (N_1607,N_185,N_1049);
xor U1608 (N_1608,N_188,N_947);
or U1609 (N_1609,In_2850,N_256);
or U1610 (N_1610,In_2586,In_737);
nor U1611 (N_1611,N_233,N_329);
nor U1612 (N_1612,N_596,In_1524);
nor U1613 (N_1613,N_197,N_884);
nand U1614 (N_1614,In_1843,In_2583);
nand U1615 (N_1615,N_632,N_1191);
nand U1616 (N_1616,N_491,N_824);
xnor U1617 (N_1617,N_936,In_108);
and U1618 (N_1618,In_1316,In_1184);
or U1619 (N_1619,N_1136,N_150);
nand U1620 (N_1620,In_2656,N_819);
xnor U1621 (N_1621,N_1105,In_750);
and U1622 (N_1622,N_337,N_200);
and U1623 (N_1623,N_474,N_11);
xnor U1624 (N_1624,In_525,N_921);
nand U1625 (N_1625,N_519,N_477);
and U1626 (N_1626,N_987,In_1827);
or U1627 (N_1627,N_1018,N_955);
nand U1628 (N_1628,N_336,N_850);
nor U1629 (N_1629,N_855,N_1132);
xor U1630 (N_1630,N_259,N_14);
or U1631 (N_1631,N_571,In_389);
nand U1632 (N_1632,N_215,N_117);
and U1633 (N_1633,In_513,N_1070);
nor U1634 (N_1634,N_455,N_711);
xnor U1635 (N_1635,N_670,N_610);
nand U1636 (N_1636,In_770,N_365);
and U1637 (N_1637,N_74,N_94);
xor U1638 (N_1638,N_10,N_23);
nor U1639 (N_1639,N_802,N_590);
xor U1640 (N_1640,N_371,N_768);
and U1641 (N_1641,N_283,N_611);
and U1642 (N_1642,N_1004,In_196);
nor U1643 (N_1643,In_2826,N_167);
xor U1644 (N_1644,N_412,N_43);
nand U1645 (N_1645,N_814,N_647);
or U1646 (N_1646,N_994,In_2697);
or U1647 (N_1647,N_827,In_2458);
nand U1648 (N_1648,N_165,N_1137);
nand U1649 (N_1649,N_966,N_920);
nor U1650 (N_1650,N_312,N_1162);
and U1651 (N_1651,N_51,In_2140);
nor U1652 (N_1652,In_1520,N_1158);
xnor U1653 (N_1653,N_916,N_4);
nand U1654 (N_1654,In_272,N_813);
nand U1655 (N_1655,N_559,N_1000);
nand U1656 (N_1656,In_2948,N_338);
xnor U1657 (N_1657,In_1100,In_1944);
nand U1658 (N_1658,In_1536,N_340);
nand U1659 (N_1659,N_1152,In_2472);
or U1660 (N_1660,N_597,N_326);
xor U1661 (N_1661,N_471,N_1189);
nand U1662 (N_1662,N_897,In_951);
nor U1663 (N_1663,N_583,N_509);
nor U1664 (N_1664,In_357,N_496);
nor U1665 (N_1665,N_3,N_663);
and U1666 (N_1666,In_144,N_104);
nor U1667 (N_1667,In_248,N_1128);
and U1668 (N_1668,N_63,N_145);
xor U1669 (N_1669,N_526,N_705);
xnor U1670 (N_1670,N_30,N_796);
or U1671 (N_1671,N_1160,In_2225);
nor U1672 (N_1672,In_1138,N_747);
nor U1673 (N_1673,N_1078,N_485);
nand U1674 (N_1674,N_1075,N_404);
and U1675 (N_1675,N_502,N_1177);
xor U1676 (N_1676,In_731,N_741);
and U1677 (N_1677,N_1,N_558);
xor U1678 (N_1678,N_466,In_2653);
nor U1679 (N_1679,N_154,N_394);
and U1680 (N_1680,N_766,N_573);
or U1681 (N_1681,In_2721,N_603);
and U1682 (N_1682,N_173,N_580);
nor U1683 (N_1683,N_880,N_1182);
and U1684 (N_1684,In_500,N_831);
and U1685 (N_1685,N_1179,N_280);
nor U1686 (N_1686,N_500,In_2715);
nor U1687 (N_1687,N_535,N_28);
nand U1688 (N_1688,In_496,N_566);
nand U1689 (N_1689,N_877,In_2428);
nor U1690 (N_1690,N_60,In_2910);
nand U1691 (N_1691,N_1153,N_89);
nand U1692 (N_1692,N_192,N_351);
or U1693 (N_1693,N_214,N_701);
xor U1694 (N_1694,N_133,N_662);
or U1695 (N_1695,N_248,In_197);
or U1696 (N_1696,N_450,N_47);
nor U1697 (N_1697,N_546,N_101);
xnor U1698 (N_1698,N_862,In_1863);
and U1699 (N_1699,N_325,In_2527);
nor U1700 (N_1700,N_1174,N_1015);
nand U1701 (N_1701,N_66,In_1008);
xnor U1702 (N_1702,N_639,N_12);
and U1703 (N_1703,In_1436,In_409);
xnor U1704 (N_1704,N_18,N_328);
nor U1705 (N_1705,N_144,N_17);
and U1706 (N_1706,N_579,In_251);
and U1707 (N_1707,In_93,N_462);
or U1708 (N_1708,N_537,N_146);
nor U1709 (N_1709,N_1192,N_1012);
and U1710 (N_1710,N_872,N_556);
and U1711 (N_1711,N_112,N_640);
nor U1712 (N_1712,N_684,N_38);
and U1713 (N_1713,N_941,N_1009);
and U1714 (N_1714,N_264,N_787);
nand U1715 (N_1715,N_1069,N_753);
or U1716 (N_1716,In_2296,N_935);
and U1717 (N_1717,In_387,N_459);
or U1718 (N_1718,N_645,N_1074);
and U1719 (N_1719,N_832,N_697);
or U1720 (N_1720,N_1118,In_2182);
nand U1721 (N_1721,N_826,N_143);
nor U1722 (N_1722,N_88,N_232);
and U1723 (N_1723,N_296,N_724);
and U1724 (N_1724,N_984,N_896);
xnor U1725 (N_1725,N_1038,In_615);
and U1726 (N_1726,N_1098,N_113);
nand U1727 (N_1727,N_750,N_1029);
nand U1728 (N_1728,N_479,N_524);
or U1729 (N_1729,N_149,In_1821);
and U1730 (N_1730,N_493,N_1001);
or U1731 (N_1731,In_2379,N_1106);
xor U1732 (N_1732,In_1124,In_1067);
nor U1733 (N_1733,N_27,In_2295);
or U1734 (N_1734,N_1117,N_795);
and U1735 (N_1735,N_1144,N_1039);
nor U1736 (N_1736,N_1091,In_297);
xor U1737 (N_1737,N_904,N_1020);
and U1738 (N_1738,In_1868,In_211);
nor U1739 (N_1739,N_472,N_284);
xnor U1740 (N_1740,N_881,In_1127);
xor U1741 (N_1741,In_13,N_1149);
xnor U1742 (N_1742,N_116,In_2429);
nand U1743 (N_1743,In_132,N_693);
or U1744 (N_1744,N_98,N_497);
nor U1745 (N_1745,N_1051,In_1453);
nand U1746 (N_1746,N_549,N_554);
nor U1747 (N_1747,In_2616,N_983);
and U1748 (N_1748,In_303,In_2870);
nand U1749 (N_1749,In_2570,In_2032);
xnor U1750 (N_1750,In_2893,N_852);
xor U1751 (N_1751,N_416,In_1676);
xor U1752 (N_1752,N_355,N_456);
xnor U1753 (N_1753,N_593,N_654);
nand U1754 (N_1754,N_313,N_995);
nor U1755 (N_1755,In_2816,N_398);
nand U1756 (N_1756,In_1508,N_77);
and U1757 (N_1757,N_871,N_874);
or U1758 (N_1758,N_260,In_655);
nor U1759 (N_1759,N_732,N_482);
nor U1760 (N_1760,In_684,N_397);
or U1761 (N_1761,In_139,In_2672);
nor U1762 (N_1762,N_988,N_553);
or U1763 (N_1763,In_2615,N_985);
nand U1764 (N_1764,N_699,N_1163);
or U1765 (N_1765,N_422,N_119);
or U1766 (N_1766,N_912,N_1146);
or U1767 (N_1767,N_59,N_70);
nand U1768 (N_1768,N_542,N_606);
or U1769 (N_1769,In_2404,N_195);
xor U1770 (N_1770,N_873,N_803);
xnor U1771 (N_1771,N_498,N_895);
or U1772 (N_1772,In_2942,N_520);
nor U1773 (N_1773,N_100,N_965);
nand U1774 (N_1774,N_836,N_748);
and U1775 (N_1775,N_536,N_712);
or U1776 (N_1776,N_938,N_512);
or U1777 (N_1777,In_1248,N_504);
nor U1778 (N_1778,N_682,In_1615);
or U1779 (N_1779,N_1154,N_996);
xor U1780 (N_1780,N_810,N_319);
xor U1781 (N_1781,N_1133,In_736);
nor U1782 (N_1782,N_487,N_839);
and U1783 (N_1783,In_2069,In_258);
and U1784 (N_1784,N_762,N_809);
and U1785 (N_1785,N_37,In_1631);
or U1786 (N_1786,In_2692,N_911);
nor U1787 (N_1787,N_717,In_1934);
nand U1788 (N_1788,N_407,N_969);
nand U1789 (N_1789,N_785,N_592);
nand U1790 (N_1790,N_356,N_484);
xor U1791 (N_1791,In_1027,N_1170);
nor U1792 (N_1792,N_634,N_818);
and U1793 (N_1793,N_196,In_2237);
nand U1794 (N_1794,In_1116,N_1019);
and U1795 (N_1795,N_379,N_729);
or U1796 (N_1796,N_629,N_692);
and U1797 (N_1797,N_721,In_1170);
xor U1798 (N_1798,In_2386,N_52);
nand U1799 (N_1799,N_218,N_589);
and U1800 (N_1800,In_418,N_866);
nor U1801 (N_1801,N_230,N_587);
xnor U1802 (N_1802,N_1092,N_409);
or U1803 (N_1803,N_868,In_2534);
xor U1804 (N_1804,N_400,N_993);
or U1805 (N_1805,In_301,N_706);
or U1806 (N_1806,N_240,N_849);
and U1807 (N_1807,N_953,N_205);
nand U1808 (N_1808,N_1119,N_221);
and U1809 (N_1809,N_1151,N_157);
or U1810 (N_1810,N_370,In_506);
or U1811 (N_1811,N_384,N_147);
or U1812 (N_1812,N_621,In_382);
nor U1813 (N_1813,N_1056,N_651);
nand U1814 (N_1814,N_786,N_906);
and U1815 (N_1815,N_1140,In_2528);
xor U1816 (N_1816,In_2841,In_1957);
nor U1817 (N_1817,N_202,N_176);
nor U1818 (N_1818,N_986,In_2241);
or U1819 (N_1819,N_475,N_1172);
or U1820 (N_1820,N_617,In_839);
and U1821 (N_1821,N_960,N_343);
nand U1822 (N_1822,N_402,In_875);
or U1823 (N_1823,In_206,N_668);
and U1824 (N_1824,N_239,N_801);
nor U1825 (N_1825,N_901,N_1065);
nand U1826 (N_1826,N_132,N_730);
and U1827 (N_1827,N_183,In_2843);
or U1828 (N_1828,In_1207,In_723);
nand U1829 (N_1829,N_174,In_250);
or U1830 (N_1830,N_226,N_543);
nand U1831 (N_1831,In_2397,N_1037);
nand U1832 (N_1832,In_342,N_414);
nand U1833 (N_1833,N_1145,N_501);
and U1834 (N_1834,In_4,N_683);
nand U1835 (N_1835,N_211,In_2890);
xnor U1836 (N_1836,In_253,In_266);
nand U1837 (N_1837,N_41,N_505);
and U1838 (N_1838,N_54,In_2396);
nand U1839 (N_1839,N_281,N_193);
or U1840 (N_1840,In_2238,N_75);
nand U1841 (N_1841,In_147,N_671);
and U1842 (N_1842,N_1180,In_2957);
or U1843 (N_1843,N_171,In_1609);
nor U1844 (N_1844,In_1697,In_952);
nor U1845 (N_1845,In_947,N_1194);
nand U1846 (N_1846,In_1297,In_374);
nand U1847 (N_1847,In_167,N_2);
and U1848 (N_1848,N_125,In_224);
or U1849 (N_1849,In_742,N_48);
nand U1850 (N_1850,In_346,In_1310);
and U1851 (N_1851,N_1199,N_980);
and U1852 (N_1852,N_1130,In_431);
xor U1853 (N_1853,In_2765,N_735);
and U1854 (N_1854,In_2087,N_311);
or U1855 (N_1855,N_297,In_1086);
and U1856 (N_1856,N_322,N_137);
or U1857 (N_1857,N_169,In_12);
nor U1858 (N_1858,N_805,N_421);
and U1859 (N_1859,In_1244,In_1160);
nand U1860 (N_1860,N_437,N_598);
and U1861 (N_1861,N_792,In_1521);
or U1862 (N_1862,In_907,N_1076);
or U1863 (N_1863,N_387,N_368);
xor U1864 (N_1864,In_1459,N_347);
nor U1865 (N_1865,In_484,N_560);
xnor U1866 (N_1866,N_282,N_244);
or U1867 (N_1867,In_843,N_761);
nor U1868 (N_1868,In_2455,N_1077);
and U1869 (N_1869,In_2628,N_1073);
xor U1870 (N_1870,In_1428,In_89);
nand U1871 (N_1871,N_348,N_1184);
and U1872 (N_1872,N_945,In_783);
or U1873 (N_1873,N_410,N_267);
nand U1874 (N_1874,N_435,In_371);
xnor U1875 (N_1875,N_463,In_909);
nand U1876 (N_1876,N_797,N_812);
nand U1877 (N_1877,In_1602,N_898);
and U1878 (N_1878,In_2294,N_782);
or U1879 (N_1879,N_8,N_547);
nor U1880 (N_1880,In_1477,N_361);
and U1881 (N_1881,In_134,In_1274);
and U1882 (N_1882,N_1115,N_594);
nor U1883 (N_1883,N_118,N_742);
nor U1884 (N_1884,N_551,N_80);
nand U1885 (N_1885,In_1000,N_667);
xor U1886 (N_1886,N_1085,N_237);
nand U1887 (N_1887,N_110,In_1118);
nand U1888 (N_1888,N_78,In_2609);
nor U1889 (N_1889,N_894,In_2599);
or U1890 (N_1890,N_1066,N_140);
nand U1891 (N_1891,N_285,N_194);
and U1892 (N_1892,N_1103,N_939);
or U1893 (N_1893,N_473,N_1100);
or U1894 (N_1894,N_979,N_529);
and U1895 (N_1895,N_209,In_2664);
xor U1896 (N_1896,N_344,In_2859);
xnor U1897 (N_1897,N_728,In_2598);
xnor U1898 (N_1898,In_273,In_1291);
or U1899 (N_1899,N_164,N_91);
xnor U1900 (N_1900,N_1017,N_126);
or U1901 (N_1901,In_769,N_470);
and U1902 (N_1902,N_295,In_2624);
nor U1903 (N_1903,In_298,In_1143);
nor U1904 (N_1904,N_726,In_2474);
or U1905 (N_1905,In_2635,N_436);
and U1906 (N_1906,N_723,N_320);
or U1907 (N_1907,N_972,In_624);
and U1908 (N_1908,N_457,In_2353);
nand U1909 (N_1909,N_572,N_739);
or U1910 (N_1910,N_1024,N_1124);
nand U1911 (N_1911,In_85,In_1532);
and U1912 (N_1912,In_1169,In_191);
xnor U1913 (N_1913,N_123,N_396);
xor U1914 (N_1914,In_1646,N_516);
xor U1915 (N_1915,In_2185,N_358);
or U1916 (N_1916,N_495,N_25);
and U1917 (N_1917,N_142,In_1830);
and U1918 (N_1918,N_612,In_1237);
and U1919 (N_1919,N_323,In_470);
or U1920 (N_1920,In_1695,In_2705);
or U1921 (N_1921,N_266,N_1079);
xnor U1922 (N_1922,N_719,N_111);
or U1923 (N_1923,N_1190,N_114);
nor U1924 (N_1924,N_703,N_184);
nand U1925 (N_1925,N_172,N_231);
nor U1926 (N_1926,In_1654,N_303);
xnor U1927 (N_1927,N_846,N_76);
nand U1928 (N_1928,N_458,N_781);
nand U1929 (N_1929,N_650,In_2772);
and U1930 (N_1930,N_778,N_162);
xnor U1931 (N_1931,N_1028,N_26);
and U1932 (N_1932,N_923,In_2918);
and U1933 (N_1933,In_1793,N_806);
xor U1934 (N_1934,In_1031,N_982);
nor U1935 (N_1935,N_964,N_499);
and U1936 (N_1936,In_724,N_1102);
or U1937 (N_1937,In_2326,N_718);
or U1938 (N_1938,In_1161,In_1799);
xor U1939 (N_1939,N_804,In_746);
nand U1940 (N_1940,N_575,N_624);
xnor U1941 (N_1941,N_578,N_1171);
nor U1942 (N_1942,N_198,In_1394);
nor U1943 (N_1943,In_571,In_2001);
and U1944 (N_1944,In_913,In_1857);
nor U1945 (N_1945,N_1161,N_891);
or U1946 (N_1946,N_33,In_440);
or U1947 (N_1947,N_944,N_190);
nor U1948 (N_1948,N_990,N_743);
nor U1949 (N_1949,N_1062,In_1391);
nand U1950 (N_1950,N_1050,N_1178);
xnor U1951 (N_1951,N_642,N_1109);
xor U1952 (N_1952,N_513,N_1126);
or U1953 (N_1953,N_269,N_353);
nand U1954 (N_1954,In_245,In_556);
nand U1955 (N_1955,In_1839,N_1135);
and U1956 (N_1956,N_949,In_1164);
nand U1957 (N_1957,In_184,In_1542);
or U1958 (N_1958,N_636,N_300);
nand U1959 (N_1959,N_376,In_2091);
nand U1960 (N_1960,N_106,In_964);
xor U1961 (N_1961,N_882,N_678);
and U1962 (N_1962,N_604,In_1906);
nand U1963 (N_1963,N_685,N_93);
nand U1964 (N_1964,In_1366,In_1190);
nor U1965 (N_1965,N_448,N_956);
and U1966 (N_1966,N_443,In_2819);
or U1967 (N_1967,N_289,N_926);
nor U1968 (N_1968,N_288,N_109);
and U1969 (N_1969,N_1011,N_279);
xnor U1970 (N_1970,N_403,N_1089);
nor U1971 (N_1971,N_369,In_777);
nor U1972 (N_1972,In_2603,N_445);
xor U1973 (N_1973,In_117,In_841);
xnor U1974 (N_1974,In_2882,N_354);
or U1975 (N_1975,N_907,In_72);
nor U1976 (N_1976,In_721,N_299);
nand U1977 (N_1977,N_431,In_2104);
and U1978 (N_1978,In_2083,In_1059);
or U1979 (N_1979,N_948,N_189);
or U1980 (N_1980,N_658,N_441);
nand U1981 (N_1981,N_223,N_87);
and U1982 (N_1982,In_1593,N_255);
nand U1983 (N_1983,N_908,N_1093);
nor U1984 (N_1984,N_696,N_293);
nand U1985 (N_1985,In_778,N_989);
nand U1986 (N_1986,In_2085,N_330);
or U1987 (N_1987,N_887,N_890);
nand U1988 (N_1988,N_160,N_478);
nand U1989 (N_1989,N_528,In_2152);
nand U1990 (N_1990,N_830,In_2005);
xnor U1991 (N_1991,N_793,N_1021);
or U1992 (N_1992,N_419,In_1640);
nor U1993 (N_1993,N_56,N_1067);
nand U1994 (N_1994,N_32,In_1553);
xor U1995 (N_1995,N_725,In_2208);
nor U1996 (N_1996,In_1775,N_301);
or U1997 (N_1997,In_2742,N_1111);
xor U1998 (N_1998,N_918,In_1683);
and U1999 (N_1999,N_1068,N_922);
xor U2000 (N_2000,N_963,N_40);
or U2001 (N_2001,In_102,In_1667);
or U2002 (N_2002,N_274,N_837);
xnor U2003 (N_2003,N_971,N_863);
nor U2004 (N_2004,N_1059,N_888);
nand U2005 (N_2005,N_464,In_763);
or U2006 (N_2006,In_2508,In_1036);
or U2007 (N_2007,N_1081,N_532);
nand U2008 (N_2008,N_1193,In_2339);
xnor U2009 (N_2009,N_675,N_727);
nor U2010 (N_2010,N_715,N_679);
and U2011 (N_2011,N_401,N_525);
and U2012 (N_2012,N_5,N_1083);
or U2013 (N_2013,N_64,N_67);
or U2014 (N_2014,N_377,N_415);
or U2015 (N_2015,In_1876,In_1499);
nor U2016 (N_2016,N_163,In_2245);
xnor U2017 (N_2017,In_666,N_1088);
nand U2018 (N_2018,N_625,N_614);
and U2019 (N_2019,In_360,N_790);
xor U2020 (N_2020,N_271,N_286);
xnor U2021 (N_2021,N_85,N_129);
and U2022 (N_2022,N_585,In_1329);
nor U2023 (N_2023,N_620,N_708);
nand U2024 (N_2024,N_373,N_268);
xor U2025 (N_2025,N_1064,N_615);
or U2026 (N_2026,N_798,In_2796);
nor U2027 (N_2027,N_808,N_823);
and U2028 (N_2028,N_480,N_784);
nand U2029 (N_2029,N_426,N_838);
nand U2030 (N_2030,In_2108,In_2613);
or U2031 (N_2031,N_961,In_2097);
and U2032 (N_2032,N_976,In_1212);
xnor U2033 (N_2033,In_20,N_816);
or U2034 (N_2034,N_599,In_1611);
nand U2035 (N_2035,In_1941,N_534);
and U2036 (N_2036,N_19,N_1131);
xor U2037 (N_2037,N_395,In_2975);
nand U2038 (N_2038,N_1014,N_305);
or U2039 (N_2039,N_1016,N_605);
or U2040 (N_2040,In_1592,N_388);
xnor U2041 (N_2041,N_208,N_381);
and U2042 (N_2042,N_854,N_820);
and U2043 (N_2043,N_550,N_1072);
nand U2044 (N_2044,In_2965,N_1048);
or U2045 (N_2045,In_786,N_1045);
or U2046 (N_2046,N_951,N_62);
xor U2047 (N_2047,In_574,N_799);
and U2048 (N_2048,N_79,N_588);
or U2049 (N_2049,In_2013,N_261);
xor U2050 (N_2050,N_633,In_2039);
and U2051 (N_2051,N_1116,In_2144);
or U2052 (N_2052,N_1142,In_1679);
nand U2053 (N_2053,N_68,N_413);
and U2054 (N_2054,N_591,N_294);
and U2055 (N_2055,In_969,N_842);
nand U2056 (N_2056,N_607,N_382);
nand U2057 (N_2057,N_42,In_652);
xor U2058 (N_2058,In_1260,In_399);
xnor U2059 (N_2059,N_425,N_1053);
or U2060 (N_2060,N_1010,In_1734);
or U2061 (N_2061,In_1094,N_1094);
nor U2062 (N_2062,In_705,N_275);
nand U2063 (N_2063,N_506,N_219);
nand U2064 (N_2064,N_843,N_453);
nand U2065 (N_2065,N_235,In_2990);
xor U2066 (N_2066,N_889,N_362);
or U2067 (N_2067,In_2502,N_616);
or U2068 (N_2068,In_2205,N_120);
and U2069 (N_2069,N_865,N_220);
or U2070 (N_2070,In_2636,N_1134);
xor U2071 (N_2071,N_619,In_237);
and U2072 (N_2072,N_1040,N_124);
nor U2073 (N_2073,N_646,N_867);
and U2074 (N_2074,N_181,N_527);
nand U2075 (N_2075,N_265,N_905);
nand U2076 (N_2076,N_754,In_1055);
or U2077 (N_2077,N_720,In_233);
or U2078 (N_2078,In_2419,N_385);
or U2079 (N_2079,In_1112,In_1846);
xnor U2080 (N_2080,In_558,In_2183);
nor U2081 (N_2081,In_2498,N_1141);
nor U2082 (N_2082,N_83,In_2203);
or U2083 (N_2083,In_2222,N_973);
or U2084 (N_2084,N_992,In_929);
or U2085 (N_2085,N_627,In_1964);
or U2086 (N_2086,In_2917,N_234);
nor U2087 (N_2087,N_187,N_222);
and U2088 (N_2088,N_731,In_2022);
or U2089 (N_2089,N_433,N_997);
and U2090 (N_2090,N_970,In_362);
or U2091 (N_2091,N_242,In_808);
xor U2092 (N_2092,In_194,In_1937);
nand U2093 (N_2093,In_2769,N_15);
and U2094 (N_2094,N_451,In_1312);
xnor U2095 (N_2095,N_107,In_44);
or U2096 (N_2096,N_103,N_440);
nand U2097 (N_2097,N_789,N_212);
and U2098 (N_2098,In_2821,N_1097);
nand U2099 (N_2099,In_1624,In_920);
or U2100 (N_2100,N_389,N_570);
nand U2101 (N_2101,In_1902,N_575);
nor U2102 (N_2102,N_642,N_38);
nor U2103 (N_2103,In_2104,In_2182);
or U2104 (N_2104,In_2705,In_1255);
and U2105 (N_2105,N_54,N_117);
and U2106 (N_2106,In_2715,N_1161);
xnor U2107 (N_2107,N_329,N_1056);
and U2108 (N_2108,In_89,N_864);
nand U2109 (N_2109,N_1016,In_2395);
xnor U2110 (N_2110,N_582,N_412);
and U2111 (N_2111,N_64,In_431);
and U2112 (N_2112,In_357,N_806);
nor U2113 (N_2113,In_2069,N_199);
or U2114 (N_2114,N_666,N_663);
and U2115 (N_2115,N_148,In_2990);
nand U2116 (N_2116,N_657,In_1310);
xor U2117 (N_2117,N_1179,In_371);
xnor U2118 (N_2118,N_332,N_705);
and U2119 (N_2119,N_701,In_2706);
xnor U2120 (N_2120,In_513,N_627);
or U2121 (N_2121,N_177,In_2527);
xor U2122 (N_2122,N_916,In_196);
nor U2123 (N_2123,In_2013,In_947);
or U2124 (N_2124,In_1969,N_675);
xnor U2125 (N_2125,N_339,In_2935);
xor U2126 (N_2126,In_2605,N_842);
and U2127 (N_2127,N_423,N_7);
nand U2128 (N_2128,N_657,N_759);
nand U2129 (N_2129,N_77,In_915);
and U2130 (N_2130,N_870,N_1142);
nor U2131 (N_2131,N_5,In_920);
and U2132 (N_2132,In_1631,N_211);
and U2133 (N_2133,In_145,In_72);
and U2134 (N_2134,N_447,N_4);
nor U2135 (N_2135,N_1043,N_81);
xnor U2136 (N_2136,In_1056,N_209);
or U2137 (N_2137,N_855,N_1135);
and U2138 (N_2138,N_184,N_231);
xnor U2139 (N_2139,N_981,N_728);
nor U2140 (N_2140,In_1994,N_810);
or U2141 (N_2141,N_195,In_2301);
and U2142 (N_2142,N_914,N_169);
and U2143 (N_2143,N_105,In_153);
xnor U2144 (N_2144,N_362,In_2674);
or U2145 (N_2145,N_214,In_2225);
xor U2146 (N_2146,In_2238,N_9);
or U2147 (N_2147,N_849,N_693);
xor U2148 (N_2148,N_575,In_1678);
or U2149 (N_2149,N_1111,N_802);
and U2150 (N_2150,N_767,N_1047);
nand U2151 (N_2151,In_2893,N_618);
xor U2152 (N_2152,N_683,N_679);
xnor U2153 (N_2153,N_250,N_622);
or U2154 (N_2154,N_160,N_103);
and U2155 (N_2155,In_2035,N_597);
xor U2156 (N_2156,In_1561,In_2969);
or U2157 (N_2157,N_594,In_2935);
nor U2158 (N_2158,In_250,N_514);
nor U2159 (N_2159,In_267,N_1151);
and U2160 (N_2160,N_547,N_16);
nor U2161 (N_2161,N_367,N_342);
nor U2162 (N_2162,N_103,N_979);
and U2163 (N_2163,In_2458,N_271);
nor U2164 (N_2164,In_792,N_343);
nand U2165 (N_2165,N_430,N_450);
or U2166 (N_2166,N_1051,N_903);
nor U2167 (N_2167,N_196,N_47);
xor U2168 (N_2168,N_90,In_777);
nor U2169 (N_2169,N_1136,N_152);
nand U2170 (N_2170,N_154,In_1654);
and U2171 (N_2171,In_1750,In_2554);
and U2172 (N_2172,N_986,N_163);
nand U2173 (N_2173,N_257,In_1109);
xor U2174 (N_2174,N_772,In_1212);
or U2175 (N_2175,N_1047,N_172);
xnor U2176 (N_2176,In_1030,In_723);
xnor U2177 (N_2177,N_509,N_121);
and U2178 (N_2178,In_2633,In_356);
nand U2179 (N_2179,In_297,N_784);
or U2180 (N_2180,N_512,N_802);
nand U2181 (N_2181,In_909,In_2605);
or U2182 (N_2182,N_552,N_847);
xor U2183 (N_2183,N_557,N_500);
nor U2184 (N_2184,N_815,N_599);
and U2185 (N_2185,N_110,In_2596);
nor U2186 (N_2186,N_1194,N_353);
nor U2187 (N_2187,N_168,N_10);
and U2188 (N_2188,N_45,N_776);
and U2189 (N_2189,N_875,N_1072);
or U2190 (N_2190,In_2958,N_132);
and U2191 (N_2191,N_448,N_18);
nand U2192 (N_2192,In_2296,N_410);
nor U2193 (N_2193,In_1615,N_656);
and U2194 (N_2194,N_394,N_987);
and U2195 (N_2195,N_988,N_1028);
or U2196 (N_2196,N_160,In_724);
nor U2197 (N_2197,N_215,N_467);
nor U2198 (N_2198,In_2950,N_1152);
xnor U2199 (N_2199,N_547,In_2957);
nand U2200 (N_2200,N_847,N_38);
and U2201 (N_2201,In_2528,N_263);
nand U2202 (N_2202,N_810,N_734);
nand U2203 (N_2203,In_132,In_1757);
nand U2204 (N_2204,N_673,N_1034);
nand U2205 (N_2205,N_1029,In_2334);
nand U2206 (N_2206,In_1164,N_358);
nand U2207 (N_2207,In_382,N_462);
nor U2208 (N_2208,In_2410,N_1135);
nor U2209 (N_2209,N_966,N_917);
nand U2210 (N_2210,N_155,N_100);
and U2211 (N_2211,N_253,N_894);
nor U2212 (N_2212,N_136,N_1100);
or U2213 (N_2213,In_2294,N_445);
nand U2214 (N_2214,N_195,N_1148);
nand U2215 (N_2215,N_303,In_1160);
nor U2216 (N_2216,N_256,N_1185);
nor U2217 (N_2217,N_394,N_726);
nor U2218 (N_2218,In_2579,In_244);
xor U2219 (N_2219,N_1119,N_1019);
nand U2220 (N_2220,N_625,In_929);
nor U2221 (N_2221,N_382,In_1775);
or U2222 (N_2222,In_2792,N_328);
or U2223 (N_2223,In_1694,In_1667);
nor U2224 (N_2224,N_184,N_173);
nand U2225 (N_2225,In_145,In_2507);
nor U2226 (N_2226,N_498,In_1222);
xnor U2227 (N_2227,N_1024,In_2298);
or U2228 (N_2228,N_236,N_702);
nand U2229 (N_2229,N_421,In_176);
xnor U2230 (N_2230,N_1145,N_779);
nor U2231 (N_2231,In_1244,In_2804);
nand U2232 (N_2232,N_972,N_890);
xor U2233 (N_2233,In_908,In_145);
and U2234 (N_2234,In_2893,In_147);
xnor U2235 (N_2235,In_2489,N_649);
or U2236 (N_2236,N_1077,N_953);
xor U2237 (N_2237,N_232,In_2508);
and U2238 (N_2238,N_549,In_1453);
nand U2239 (N_2239,In_1059,N_511);
and U2240 (N_2240,N_714,N_501);
and U2241 (N_2241,In_2489,In_2048);
or U2242 (N_2242,N_879,N_259);
or U2243 (N_2243,N_353,In_1564);
nor U2244 (N_2244,N_1182,In_769);
xnor U2245 (N_2245,N_525,In_1313);
nand U2246 (N_2246,N_599,N_359);
xor U2247 (N_2247,N_845,N_627);
nand U2248 (N_2248,In_2958,In_2353);
nor U2249 (N_2249,N_469,N_275);
xnor U2250 (N_2250,N_7,In_297);
nand U2251 (N_2251,N_848,N_133);
nand U2252 (N_2252,N_739,N_327);
xor U2253 (N_2253,N_183,In_2664);
and U2254 (N_2254,In_736,In_2965);
and U2255 (N_2255,N_925,N_716);
and U2256 (N_2256,N_42,N_723);
and U2257 (N_2257,N_674,N_19);
nand U2258 (N_2258,N_921,N_538);
and U2259 (N_2259,N_981,N_364);
or U2260 (N_2260,In_139,In_77);
and U2261 (N_2261,N_429,N_230);
nor U2262 (N_2262,N_500,N_1030);
nand U2263 (N_2263,N_447,In_2121);
xnor U2264 (N_2264,N_1122,In_1906);
nor U2265 (N_2265,N_322,In_1654);
xor U2266 (N_2266,In_2428,N_1018);
xor U2267 (N_2267,N_1124,N_655);
and U2268 (N_2268,In_410,In_431);
nand U2269 (N_2269,In_2183,N_432);
xnor U2270 (N_2270,N_762,In_1202);
and U2271 (N_2271,N_1136,N_756);
or U2272 (N_2272,N_931,N_65);
and U2273 (N_2273,N_1137,N_1084);
xnor U2274 (N_2274,In_2616,N_328);
or U2275 (N_2275,N_799,N_1107);
and U2276 (N_2276,N_883,N_392);
or U2277 (N_2277,N_96,N_566);
nand U2278 (N_2278,In_251,In_910);
and U2279 (N_2279,In_1994,In_211);
and U2280 (N_2280,In_952,N_441);
xnor U2281 (N_2281,N_871,In_1944);
nor U2282 (N_2282,N_111,N_760);
or U2283 (N_2283,N_1161,N_1001);
nand U2284 (N_2284,N_934,N_8);
and U2285 (N_2285,In_1657,N_1049);
nand U2286 (N_2286,N_231,In_2507);
or U2287 (N_2287,N_197,In_906);
nand U2288 (N_2288,N_1009,In_1404);
and U2289 (N_2289,N_965,N_1114);
nor U2290 (N_2290,In_387,N_372);
nand U2291 (N_2291,In_1477,N_965);
nor U2292 (N_2292,N_303,N_213);
nor U2293 (N_2293,In_245,In_1459);
nor U2294 (N_2294,In_2990,N_168);
and U2295 (N_2295,N_631,N_671);
nand U2296 (N_2296,N_983,In_184);
or U2297 (N_2297,In_1274,N_624);
nor U2298 (N_2298,N_330,In_705);
xnor U2299 (N_2299,In_1329,N_730);
nor U2300 (N_2300,N_809,N_1131);
nand U2301 (N_2301,In_611,N_552);
nor U2302 (N_2302,In_2957,In_2334);
xnor U2303 (N_2303,N_693,N_130);
xor U2304 (N_2304,In_2507,N_822);
or U2305 (N_2305,N_435,N_632);
xnor U2306 (N_2306,N_507,In_1617);
xor U2307 (N_2307,N_966,N_62);
or U2308 (N_2308,N_503,N_1077);
and U2309 (N_2309,N_661,N_97);
nand U2310 (N_2310,In_1244,In_2396);
nand U2311 (N_2311,In_2375,In_1863);
and U2312 (N_2312,N_773,N_893);
nand U2313 (N_2313,N_451,N_464);
nor U2314 (N_2314,In_813,N_1147);
xor U2315 (N_2315,N_425,N_158);
xnor U2316 (N_2316,N_197,N_313);
nor U2317 (N_2317,N_81,N_548);
nand U2318 (N_2318,In_2904,N_1073);
or U2319 (N_2319,N_753,N_431);
nor U2320 (N_2320,N_856,N_655);
or U2321 (N_2321,N_739,In_2839);
nand U2322 (N_2322,In_2579,In_1264);
xnor U2323 (N_2323,N_1,N_883);
and U2324 (N_2324,N_779,N_34);
or U2325 (N_2325,N_224,N_565);
nor U2326 (N_2326,In_1732,N_730);
and U2327 (N_2327,In_2552,N_407);
xnor U2328 (N_2328,N_1127,In_2730);
xor U2329 (N_2329,N_144,N_359);
or U2330 (N_2330,N_109,N_557);
nand U2331 (N_2331,N_1148,N_966);
or U2332 (N_2332,N_102,N_460);
nor U2333 (N_2333,N_500,N_717);
nand U2334 (N_2334,In_2121,In_20);
and U2335 (N_2335,In_2282,N_78);
nor U2336 (N_2336,N_1045,N_331);
nor U2337 (N_2337,N_282,N_1102);
and U2338 (N_2338,In_513,N_561);
and U2339 (N_2339,In_1564,N_301);
and U2340 (N_2340,N_734,In_1237);
xnor U2341 (N_2341,N_998,In_1428);
nand U2342 (N_2342,In_500,N_719);
or U2343 (N_2343,N_278,N_300);
nor U2344 (N_2344,N_195,N_739);
or U2345 (N_2345,In_1977,In_2707);
or U2346 (N_2346,N_1117,In_134);
or U2347 (N_2347,N_1060,N_329);
nor U2348 (N_2348,N_807,N_359);
xnor U2349 (N_2349,In_971,N_709);
nor U2350 (N_2350,N_205,N_1004);
xor U2351 (N_2351,N_626,N_110);
xor U2352 (N_2352,N_450,In_357);
xnor U2353 (N_2353,In_145,N_730);
nor U2354 (N_2354,N_1069,N_233);
xnor U2355 (N_2355,N_434,N_1011);
or U2356 (N_2356,N_576,N_435);
and U2357 (N_2357,N_876,N_54);
nor U2358 (N_2358,N_1185,N_829);
or U2359 (N_2359,N_645,In_624);
or U2360 (N_2360,N_479,N_824);
and U2361 (N_2361,N_211,N_746);
or U2362 (N_2362,N_38,In_1431);
and U2363 (N_2363,N_821,N_720);
and U2364 (N_2364,N_919,N_665);
or U2365 (N_2365,N_161,In_1052);
or U2366 (N_2366,N_783,N_825);
xor U2367 (N_2367,N_315,N_66);
and U2368 (N_2368,N_887,N_857);
xor U2369 (N_2369,N_897,N_688);
nand U2370 (N_2370,In_713,N_340);
nor U2371 (N_2371,N_39,In_1561);
and U2372 (N_2372,N_881,N_436);
or U2373 (N_2373,N_134,N_1108);
nor U2374 (N_2374,N_986,N_242);
nand U2375 (N_2375,In_389,N_614);
nor U2376 (N_2376,In_2917,N_1182);
and U2377 (N_2377,In_2674,In_233);
or U2378 (N_2378,In_705,N_507);
nand U2379 (N_2379,In_2183,N_967);
nand U2380 (N_2380,In_792,In_1964);
or U2381 (N_2381,N_502,In_2498);
and U2382 (N_2382,N_379,In_742);
nor U2383 (N_2383,In_2870,N_660);
nor U2384 (N_2384,In_791,In_1602);
and U2385 (N_2385,N_289,N_798);
nand U2386 (N_2386,N_128,In_2032);
xor U2387 (N_2387,N_697,In_1274);
nand U2388 (N_2388,N_1066,N_749);
nor U2389 (N_2389,In_1615,N_662);
or U2390 (N_2390,N_555,N_431);
or U2391 (N_2391,N_278,In_1274);
or U2392 (N_2392,In_1438,N_836);
nor U2393 (N_2393,N_933,In_2152);
xnor U2394 (N_2394,N_144,N_464);
nand U2395 (N_2395,N_171,In_2792);
or U2396 (N_2396,N_816,N_351);
nand U2397 (N_2397,In_1190,N_561);
xor U2398 (N_2398,N_115,N_853);
nand U2399 (N_2399,N_628,N_24);
xnor U2400 (N_2400,N_1801,N_1583);
xnor U2401 (N_2401,N_1218,N_1958);
or U2402 (N_2402,N_1393,N_2138);
nand U2403 (N_2403,N_1841,N_1299);
xor U2404 (N_2404,N_1296,N_2069);
nor U2405 (N_2405,N_1365,N_2083);
nand U2406 (N_2406,N_1873,N_2166);
or U2407 (N_2407,N_2393,N_1919);
or U2408 (N_2408,N_1656,N_1658);
or U2409 (N_2409,N_1771,N_2171);
or U2410 (N_2410,N_2297,N_1434);
and U2411 (N_2411,N_2137,N_1861);
and U2412 (N_2412,N_2139,N_1741);
nor U2413 (N_2413,N_2046,N_1837);
xnor U2414 (N_2414,N_1854,N_1551);
and U2415 (N_2415,N_2263,N_2006);
and U2416 (N_2416,N_1680,N_1473);
and U2417 (N_2417,N_1904,N_1376);
or U2418 (N_2418,N_1884,N_1791);
nand U2419 (N_2419,N_1682,N_1731);
xnor U2420 (N_2420,N_1864,N_1310);
xor U2421 (N_2421,N_2024,N_1881);
or U2422 (N_2422,N_2042,N_1575);
and U2423 (N_2423,N_2034,N_2243);
or U2424 (N_2424,N_1664,N_1942);
or U2425 (N_2425,N_2193,N_1219);
xnor U2426 (N_2426,N_1311,N_2076);
nor U2427 (N_2427,N_2224,N_2308);
and U2428 (N_2428,N_2296,N_1670);
or U2429 (N_2429,N_1825,N_1866);
or U2430 (N_2430,N_1389,N_2347);
nand U2431 (N_2431,N_1996,N_1776);
nand U2432 (N_2432,N_1792,N_2064);
nand U2433 (N_2433,N_2339,N_1752);
nor U2434 (N_2434,N_1449,N_1208);
nor U2435 (N_2435,N_1924,N_1785);
nor U2436 (N_2436,N_1464,N_1348);
and U2437 (N_2437,N_2159,N_2092);
xor U2438 (N_2438,N_1950,N_2055);
and U2439 (N_2439,N_1725,N_2309);
xnor U2440 (N_2440,N_2188,N_1428);
nand U2441 (N_2441,N_1654,N_1323);
xnor U2442 (N_2442,N_1250,N_1306);
nor U2443 (N_2443,N_1522,N_1346);
or U2444 (N_2444,N_1511,N_1369);
or U2445 (N_2445,N_1615,N_2161);
xnor U2446 (N_2446,N_1391,N_2189);
nor U2447 (N_2447,N_1759,N_2081);
xor U2448 (N_2448,N_2218,N_2269);
or U2449 (N_2449,N_1778,N_1253);
nor U2450 (N_2450,N_1733,N_2094);
nand U2451 (N_2451,N_2180,N_1216);
or U2452 (N_2452,N_2281,N_1377);
xor U2453 (N_2453,N_1698,N_1274);
or U2454 (N_2454,N_2089,N_1380);
xnor U2455 (N_2455,N_2254,N_2082);
or U2456 (N_2456,N_2031,N_2118);
xnor U2457 (N_2457,N_1364,N_2372);
nand U2458 (N_2458,N_1634,N_2172);
and U2459 (N_2459,N_2348,N_2387);
nor U2460 (N_2460,N_1852,N_1651);
or U2461 (N_2461,N_1246,N_2066);
nor U2462 (N_2462,N_2268,N_1401);
nand U2463 (N_2463,N_1489,N_2025);
and U2464 (N_2464,N_1640,N_2345);
nor U2465 (N_2465,N_1315,N_1435);
and U2466 (N_2466,N_1977,N_2020);
xor U2467 (N_2467,N_1684,N_1674);
xor U2468 (N_2468,N_1840,N_1321);
nand U2469 (N_2469,N_1912,N_1993);
or U2470 (N_2470,N_1662,N_1363);
nand U2471 (N_2471,N_1200,N_2340);
and U2472 (N_2472,N_1520,N_1989);
or U2473 (N_2473,N_1598,N_2298);
and U2474 (N_2474,N_1477,N_1342);
nand U2475 (N_2475,N_1782,N_2100);
xor U2476 (N_2476,N_1202,N_2014);
xor U2477 (N_2477,N_1987,N_2003);
and U2478 (N_2478,N_1659,N_2107);
xor U2479 (N_2479,N_2067,N_1982);
and U2480 (N_2480,N_1984,N_1638);
xor U2481 (N_2481,N_1563,N_2214);
nand U2482 (N_2482,N_1675,N_1382);
xor U2483 (N_2483,N_1749,N_2292);
xnor U2484 (N_2484,N_1480,N_1609);
xnor U2485 (N_2485,N_1244,N_2049);
nand U2486 (N_2486,N_1230,N_2145);
nand U2487 (N_2487,N_1234,N_2197);
or U2488 (N_2488,N_1605,N_2096);
xnor U2489 (N_2489,N_2132,N_2093);
xor U2490 (N_2490,N_1264,N_2070);
or U2491 (N_2491,N_1702,N_1407);
xor U2492 (N_2492,N_1343,N_1751);
and U2493 (N_2493,N_2277,N_1220);
xor U2494 (N_2494,N_1655,N_1732);
and U2495 (N_2495,N_1813,N_1880);
or U2496 (N_2496,N_2129,N_2141);
xnor U2497 (N_2497,N_1829,N_1593);
or U2498 (N_2498,N_2349,N_1330);
xor U2499 (N_2499,N_1454,N_1579);
nor U2500 (N_2500,N_1737,N_1341);
or U2501 (N_2501,N_2110,N_2160);
nor U2502 (N_2502,N_2383,N_1436);
or U2503 (N_2503,N_1663,N_2265);
or U2504 (N_2504,N_2379,N_2163);
xnor U2505 (N_2505,N_1602,N_1902);
nand U2506 (N_2506,N_1440,N_2285);
xnor U2507 (N_2507,N_1843,N_1922);
xnor U2508 (N_2508,N_2019,N_2208);
xor U2509 (N_2509,N_1328,N_1576);
xnor U2510 (N_2510,N_1953,N_2264);
nand U2511 (N_2511,N_2305,N_1398);
or U2512 (N_2512,N_2078,N_1236);
and U2513 (N_2513,N_2018,N_1552);
or U2514 (N_2514,N_1985,N_1340);
or U2515 (N_2515,N_2050,N_2358);
or U2516 (N_2516,N_1920,N_2356);
nor U2517 (N_2517,N_1603,N_1915);
or U2518 (N_2518,N_1974,N_1907);
and U2519 (N_2519,N_1859,N_1764);
and U2520 (N_2520,N_1925,N_1461);
and U2521 (N_2521,N_1860,N_2306);
nand U2522 (N_2522,N_1894,N_1476);
xor U2523 (N_2523,N_1292,N_1877);
and U2524 (N_2524,N_1952,N_2182);
nand U2525 (N_2525,N_1734,N_2157);
xor U2526 (N_2526,N_1758,N_1333);
nor U2527 (N_2527,N_1217,N_2337);
nand U2528 (N_2528,N_1972,N_1788);
xor U2529 (N_2529,N_2017,N_2116);
or U2530 (N_2530,N_1694,N_1370);
nor U2531 (N_2531,N_2114,N_1558);
nand U2532 (N_2532,N_2127,N_1688);
nand U2533 (N_2533,N_1503,N_1505);
and U2534 (N_2534,N_1297,N_1997);
xnor U2535 (N_2535,N_2242,N_1275);
xor U2536 (N_2536,N_2183,N_1222);
nand U2537 (N_2537,N_1258,N_1312);
nor U2538 (N_2538,N_2205,N_1381);
nand U2539 (N_2539,N_2385,N_1903);
or U2540 (N_2540,N_2131,N_1777);
or U2541 (N_2541,N_2290,N_1945);
nor U2542 (N_2542,N_2375,N_1644);
nor U2543 (N_2543,N_1452,N_1283);
and U2544 (N_2544,N_1307,N_1775);
xnor U2545 (N_2545,N_1999,N_1351);
nand U2546 (N_2546,N_2152,N_1541);
nor U2547 (N_2547,N_1613,N_1232);
nand U2548 (N_2548,N_2270,N_2267);
and U2549 (N_2549,N_1677,N_1951);
xnor U2550 (N_2550,N_1665,N_2261);
nor U2551 (N_2551,N_1429,N_2235);
nor U2552 (N_2552,N_1905,N_2158);
or U2553 (N_2553,N_2097,N_2051);
or U2554 (N_2554,N_1286,N_1544);
nand U2555 (N_2555,N_2148,N_1700);
or U2556 (N_2556,N_1445,N_2090);
nor U2557 (N_2557,N_1448,N_2095);
nor U2558 (N_2558,N_1358,N_1291);
nor U2559 (N_2559,N_1462,N_1366);
and U2560 (N_2560,N_2319,N_1507);
nand U2561 (N_2561,N_1490,N_1709);
and U2562 (N_2562,N_1846,N_2043);
or U2563 (N_2563,N_1225,N_1529);
nor U2564 (N_2564,N_1303,N_1305);
nand U2565 (N_2565,N_1413,N_1475);
and U2566 (N_2566,N_1320,N_1392);
or U2567 (N_2567,N_1833,N_1616);
xor U2568 (N_2568,N_1517,N_1645);
nor U2569 (N_2569,N_1523,N_1271);
nand U2570 (N_2570,N_1223,N_1772);
or U2571 (N_2571,N_2362,N_2212);
nand U2572 (N_2572,N_1302,N_2217);
nor U2573 (N_2573,N_2185,N_2350);
nor U2574 (N_2574,N_1963,N_1712);
nor U2575 (N_2575,N_1612,N_1756);
or U2576 (N_2576,N_1988,N_2035);
or U2577 (N_2577,N_2237,N_2251);
nor U2578 (N_2578,N_1339,N_1930);
or U2579 (N_2579,N_1637,N_1409);
or U2580 (N_2580,N_2143,N_2029);
and U2581 (N_2581,N_1269,N_1789);
nand U2582 (N_2582,N_1543,N_1584);
nor U2583 (N_2583,N_2311,N_1898);
or U2584 (N_2584,N_1360,N_1278);
xor U2585 (N_2585,N_1309,N_2213);
and U2586 (N_2586,N_1273,N_2088);
nand U2587 (N_2587,N_2073,N_1243);
and U2588 (N_2588,N_2147,N_1395);
nand U2589 (N_2589,N_1750,N_1578);
and U2590 (N_2590,N_1815,N_1760);
nor U2591 (N_2591,N_1384,N_1743);
and U2592 (N_2592,N_1808,N_1876);
and U2593 (N_2593,N_2388,N_1372);
xnor U2594 (N_2594,N_1798,N_2004);
nor U2595 (N_2595,N_1221,N_1574);
or U2596 (N_2596,N_1538,N_2109);
and U2597 (N_2597,N_2239,N_1835);
and U2598 (N_2598,N_1405,N_1590);
and U2599 (N_2599,N_2300,N_2316);
nand U2600 (N_2600,N_1617,N_1493);
nand U2601 (N_2601,N_1308,N_1806);
or U2602 (N_2602,N_2156,N_1765);
xor U2603 (N_2603,N_1948,N_2274);
nor U2604 (N_2604,N_1444,N_1937);
nor U2605 (N_2605,N_1495,N_2091);
nand U2606 (N_2606,N_1685,N_1931);
xor U2607 (N_2607,N_2133,N_1716);
nor U2608 (N_2608,N_1539,N_1497);
and U2609 (N_2609,N_2048,N_1823);
and U2610 (N_2610,N_1726,N_2085);
nand U2611 (N_2611,N_1766,N_2325);
xnor U2612 (N_2612,N_2200,N_1371);
xor U2613 (N_2613,N_1783,N_2226);
xor U2614 (N_2614,N_1414,N_2369);
nand U2615 (N_2615,N_1272,N_2164);
or U2616 (N_2616,N_2009,N_1865);
or U2617 (N_2617,N_1532,N_2355);
and U2618 (N_2618,N_1588,N_1839);
nand U2619 (N_2619,N_1828,N_1779);
and U2620 (N_2620,N_1387,N_1367);
xor U2621 (N_2621,N_2351,N_1239);
and U2622 (N_2622,N_1738,N_2357);
and U2623 (N_2623,N_2253,N_1285);
nor U2624 (N_2624,N_1241,N_1991);
nand U2625 (N_2625,N_1453,N_1643);
xor U2626 (N_2626,N_2317,N_1567);
nand U2627 (N_2627,N_2244,N_1883);
xnor U2628 (N_2628,N_2016,N_1862);
and U2629 (N_2629,N_2045,N_1425);
or U2630 (N_2630,N_1550,N_1418);
and U2631 (N_2631,N_1796,N_2262);
nand U2632 (N_2632,N_1513,N_2390);
or U2633 (N_2633,N_1857,N_2255);
nand U2634 (N_2634,N_1383,N_2104);
or U2635 (N_2635,N_1284,N_1251);
or U2636 (N_2636,N_1368,N_2230);
and U2637 (N_2637,N_1402,N_1975);
and U2638 (N_2638,N_2001,N_1838);
xnor U2639 (N_2639,N_2123,N_2209);
or U2640 (N_2640,N_1591,N_1926);
and U2641 (N_2641,N_1349,N_2284);
nand U2642 (N_2642,N_1748,N_1800);
xnor U2643 (N_2643,N_1938,N_2301);
nor U2644 (N_2644,N_2323,N_1396);
or U2645 (N_2645,N_2010,N_1882);
xnor U2646 (N_2646,N_1636,N_1795);
xnor U2647 (N_2647,N_2063,N_2169);
nand U2648 (N_2648,N_1652,N_1728);
nor U2649 (N_2649,N_1889,N_1548);
and U2650 (N_2650,N_2338,N_1786);
or U2651 (N_2651,N_2008,N_1207);
xnor U2652 (N_2652,N_1667,N_2059);
or U2653 (N_2653,N_1531,N_1842);
and U2654 (N_2654,N_1754,N_1630);
xor U2655 (N_2655,N_1356,N_1720);
and U2656 (N_2656,N_2115,N_1502);
nor U2657 (N_2657,N_1727,N_2130);
xnor U2658 (N_2658,N_1515,N_1679);
xnor U2659 (N_2659,N_1212,N_1488);
or U2660 (N_2660,N_1594,N_1460);
and U2661 (N_2661,N_1281,N_1474);
nor U2662 (N_2662,N_2223,N_1962);
or U2663 (N_2663,N_1411,N_1378);
or U2664 (N_2664,N_1535,N_1561);
nand U2665 (N_2665,N_1932,N_1954);
or U2666 (N_2666,N_1500,N_2135);
xnor U2667 (N_2667,N_2366,N_2330);
xnor U2668 (N_2668,N_1885,N_1908);
or U2669 (N_2669,N_1794,N_1501);
xor U2670 (N_2670,N_1465,N_1471);
nor U2671 (N_2671,N_1277,N_1830);
nor U2672 (N_2672,N_1441,N_1247);
nand U2673 (N_2673,N_2077,N_2038);
nor U2674 (N_2674,N_1821,N_2221);
nor U2675 (N_2675,N_1438,N_1761);
nand U2676 (N_2676,N_1781,N_2275);
xor U2677 (N_2677,N_1432,N_1479);
nand U2678 (N_2678,N_1293,N_2322);
and U2679 (N_2679,N_1468,N_1201);
nand U2680 (N_2680,N_1611,N_2178);
and U2681 (N_2681,N_2032,N_1762);
xnor U2682 (N_2682,N_2273,N_2304);
or U2683 (N_2683,N_1929,N_2030);
xnor U2684 (N_2684,N_2344,N_1856);
and U2685 (N_2685,N_1868,N_1506);
nor U2686 (N_2686,N_1521,N_2392);
and U2687 (N_2687,N_1601,N_1362);
and U2688 (N_2688,N_2398,N_1899);
nand U2689 (N_2689,N_1450,N_2288);
nor U2690 (N_2690,N_2062,N_1256);
xor U2691 (N_2691,N_2376,N_1580);
nor U2692 (N_2692,N_2382,N_1624);
and U2693 (N_2693,N_1276,N_2365);
and U2694 (N_2694,N_1487,N_2187);
and U2695 (N_2695,N_2236,N_1946);
nor U2696 (N_2696,N_1910,N_2037);
xor U2697 (N_2697,N_1970,N_1562);
xor U2698 (N_2698,N_1990,N_2011);
and U2699 (N_2699,N_2053,N_1206);
nor U2700 (N_2700,N_1397,N_1417);
nor U2701 (N_2701,N_1683,N_1755);
nor U2702 (N_2702,N_1824,N_1867);
nor U2703 (N_2703,N_1242,N_1848);
nand U2704 (N_2704,N_1690,N_2151);
or U2705 (N_2705,N_1357,N_2314);
nor U2706 (N_2706,N_2012,N_1324);
nand U2707 (N_2707,N_1971,N_1676);
or U2708 (N_2708,N_1622,N_1470);
xor U2709 (N_2709,N_1210,N_1510);
xor U2710 (N_2710,N_1701,N_1485);
and U2711 (N_2711,N_1718,N_2033);
and U2712 (N_2712,N_1836,N_2216);
xor U2713 (N_2713,N_1729,N_2287);
nand U2714 (N_2714,N_2179,N_1966);
or U2715 (N_2715,N_1648,N_2399);
and U2716 (N_2716,N_1205,N_2334);
and U2717 (N_2717,N_1623,N_1629);
nand U2718 (N_2718,N_1774,N_1433);
nor U2719 (N_2719,N_1812,N_1322);
xnor U2720 (N_2720,N_1332,N_1335);
or U2721 (N_2721,N_1304,N_2154);
xor U2722 (N_2722,N_2155,N_1282);
xor U2723 (N_2723,N_2234,N_2289);
and U2724 (N_2724,N_1509,N_2136);
and U2725 (N_2725,N_1592,N_1831);
and U2726 (N_2726,N_2260,N_1618);
or U2727 (N_2727,N_1534,N_1900);
xor U2728 (N_2728,N_1625,N_1939);
and U2729 (N_2729,N_1666,N_1537);
xnor U2730 (N_2730,N_1847,N_1635);
and U2731 (N_2731,N_2039,N_1375);
xnor U2732 (N_2732,N_1496,N_2283);
nand U2733 (N_2733,N_1810,N_1514);
and U2734 (N_2734,N_1607,N_1295);
and U2735 (N_2735,N_2346,N_1226);
and U2736 (N_2736,N_1359,N_2302);
xor U2737 (N_2737,N_1944,N_2201);
or U2738 (N_2738,N_1257,N_1653);
and U2739 (N_2739,N_1909,N_1901);
nor U2740 (N_2740,N_1849,N_2353);
xor U2741 (N_2741,N_1650,N_2219);
nand U2742 (N_2742,N_2103,N_2240);
and U2743 (N_2743,N_1459,N_2360);
nor U2744 (N_2744,N_1252,N_1995);
nand U2745 (N_2745,N_2199,N_1316);
xnor U2746 (N_2746,N_1446,N_1294);
xnor U2747 (N_2747,N_2086,N_1784);
xnor U2748 (N_2748,N_1317,N_1259);
nor U2749 (N_2749,N_2047,N_1681);
xnor U2750 (N_2750,N_2105,N_1628);
nor U2751 (N_2751,N_1710,N_1355);
nand U2752 (N_2752,N_1326,N_1227);
nor U2753 (N_2753,N_2162,N_2056);
xor U2754 (N_2754,N_1739,N_1527);
nand U2755 (N_2755,N_1268,N_1672);
xor U2756 (N_2756,N_2370,N_2052);
xnor U2757 (N_2757,N_1668,N_1211);
xnor U2758 (N_2758,N_1818,N_2175);
nand U2759 (N_2759,N_1519,N_1770);
xor U2760 (N_2760,N_2331,N_2238);
nor U2761 (N_2761,N_1373,N_1641);
nor U2762 (N_2762,N_1319,N_1879);
nand U2763 (N_2763,N_1458,N_1832);
xor U2764 (N_2764,N_1735,N_1482);
nand U2765 (N_2765,N_1853,N_2198);
and U2766 (N_2766,N_1714,N_1385);
xor U2767 (N_2767,N_1965,N_1255);
nand U2768 (N_2768,N_2380,N_1516);
nand U2769 (N_2769,N_1705,N_1826);
or U2770 (N_2770,N_2326,N_1466);
xor U2771 (N_2771,N_1267,N_2386);
or U2772 (N_2772,N_2315,N_2303);
and U2773 (N_2773,N_1298,N_2168);
xnor U2774 (N_2774,N_1213,N_1911);
nor U2775 (N_2775,N_1757,N_1960);
nor U2776 (N_2776,N_1621,N_1586);
nand U2777 (N_2777,N_2057,N_2395);
nor U2778 (N_2778,N_1695,N_1707);
nand U2779 (N_2779,N_1708,N_1642);
and U2780 (N_2780,N_1888,N_1745);
or U2781 (N_2781,N_1992,N_1973);
or U2782 (N_2782,N_2246,N_2332);
or U2783 (N_2783,N_2027,N_2101);
or U2784 (N_2784,N_1631,N_1768);
xor U2785 (N_2785,N_1740,N_2391);
and U2786 (N_2786,N_1261,N_1978);
or U2787 (N_2787,N_2146,N_2000);
xor U2788 (N_2788,N_2333,N_2191);
and U2789 (N_2789,N_2065,N_1290);
and U2790 (N_2790,N_2310,N_1265);
xor U2791 (N_2791,N_1235,N_1518);
or U2792 (N_2792,N_1270,N_1964);
xor U2793 (N_2793,N_1231,N_1439);
or U2794 (N_2794,N_1671,N_1412);
nand U2795 (N_2795,N_1935,N_2227);
or U2796 (N_2796,N_1215,N_1240);
or U2797 (N_2797,N_1814,N_2225);
and U2798 (N_2798,N_1981,N_1715);
or U2799 (N_2799,N_1921,N_2228);
nand U2800 (N_2800,N_2271,N_1742);
xor U2801 (N_2801,N_1689,N_1704);
or U2802 (N_2802,N_2007,N_2134);
or U2803 (N_2803,N_2215,N_1870);
or U2804 (N_2804,N_1325,N_2194);
or U2805 (N_2805,N_1570,N_1390);
xor U2806 (N_2806,N_1336,N_1481);
xor U2807 (N_2807,N_1416,N_1906);
nor U2808 (N_2808,N_2026,N_1546);
nor U2809 (N_2809,N_1573,N_1933);
nor U2810 (N_2810,N_2282,N_1969);
nor U2811 (N_2811,N_1260,N_2327);
xor U2812 (N_2812,N_1338,N_1895);
nor U2813 (N_2813,N_1940,N_2318);
nor U2814 (N_2814,N_1404,N_1891);
nand U2815 (N_2815,N_1803,N_2378);
or U2816 (N_2816,N_2108,N_1976);
or U2817 (N_2817,N_1540,N_1352);
and U2818 (N_2818,N_1887,N_1620);
or U2819 (N_2819,N_1724,N_1787);
or U2820 (N_2820,N_1746,N_1632);
nand U2821 (N_2821,N_1331,N_1673);
or U2822 (N_2822,N_1424,N_1566);
nor U2823 (N_2823,N_2125,N_1400);
and U2824 (N_2824,N_1512,N_1804);
or U2825 (N_2825,N_1499,N_2071);
nand U2826 (N_2826,N_1585,N_1530);
nand U2827 (N_2827,N_1819,N_1203);
and U2828 (N_2828,N_1721,N_2374);
and U2829 (N_2829,N_1722,N_1427);
xor U2830 (N_2830,N_1442,N_1279);
and U2831 (N_2831,N_1869,N_1457);
and U2832 (N_2832,N_1560,N_2196);
nor U2833 (N_2833,N_2248,N_1802);
xnor U2834 (N_2834,N_1587,N_1536);
nand U2835 (N_2835,N_1229,N_1245);
nor U2836 (N_2836,N_1415,N_1896);
and U2837 (N_2837,N_1918,N_1492);
and U2838 (N_2838,N_1811,N_2329);
and U2839 (N_2839,N_1564,N_2257);
nand U2840 (N_2840,N_1855,N_1957);
xnor U2841 (N_2841,N_1559,N_2258);
nand U2842 (N_2842,N_2256,N_1753);
nand U2843 (N_2843,N_1713,N_1554);
or U2844 (N_2844,N_1955,N_2394);
and U2845 (N_2845,N_1334,N_2294);
and U2846 (N_2846,N_2079,N_1287);
or U2847 (N_2847,N_2022,N_1483);
and U2848 (N_2848,N_1890,N_1508);
or U2849 (N_2849,N_1809,N_1524);
xor U2850 (N_2850,N_1968,N_1967);
xnor U2851 (N_2851,N_1249,N_1805);
nand U2852 (N_2852,N_2099,N_1769);
nand U2853 (N_2853,N_1678,N_2174);
nand U2854 (N_2854,N_1597,N_2074);
or U2855 (N_2855,N_2211,N_2259);
or U2856 (N_2856,N_1610,N_1467);
nor U2857 (N_2857,N_1379,N_2142);
or U2858 (N_2858,N_2222,N_1844);
or U2859 (N_2859,N_1350,N_1525);
xor U2860 (N_2860,N_1595,N_1542);
and U2861 (N_2861,N_1872,N_1913);
or U2862 (N_2862,N_1820,N_1431);
or U2863 (N_2863,N_2015,N_1947);
or U2864 (N_2864,N_1699,N_1943);
xor U2865 (N_2865,N_1314,N_1248);
nand U2866 (N_2866,N_1914,N_1301);
and U2867 (N_2867,N_1565,N_2286);
nand U2868 (N_2868,N_1851,N_1289);
and U2869 (N_2869,N_1797,N_1263);
xor U2870 (N_2870,N_1410,N_2140);
and U2871 (N_2871,N_2352,N_2021);
and U2872 (N_2872,N_2150,N_1555);
xnor U2873 (N_2873,N_1353,N_2312);
xnor U2874 (N_2874,N_1577,N_1419);
and U2875 (N_2875,N_1730,N_1723);
and U2876 (N_2876,N_1691,N_1692);
nand U2877 (N_2877,N_2328,N_1545);
nand U2878 (N_2878,N_2124,N_1443);
xor U2879 (N_2879,N_2266,N_1661);
nor U2880 (N_2880,N_1706,N_1646);
nor U2881 (N_2881,N_1669,N_2186);
nor U2882 (N_2882,N_1486,N_1994);
nor U2883 (N_2883,N_1214,N_2291);
and U2884 (N_2884,N_2364,N_1568);
xor U2885 (N_2885,N_1850,N_1209);
xor U2886 (N_2886,N_2206,N_2190);
xnor U2887 (N_2887,N_2084,N_1347);
xnor U2888 (N_2888,N_1233,N_1822);
or U2889 (N_2889,N_2232,N_1858);
nor U2890 (N_2890,N_1547,N_1799);
and U2891 (N_2891,N_1936,N_2343);
or U2892 (N_2892,N_2192,N_2195);
nand U2893 (N_2893,N_1557,N_2181);
or U2894 (N_2894,N_1686,N_1927);
and U2895 (N_2895,N_1817,N_2220);
nand U2896 (N_2896,N_1361,N_1875);
nand U2897 (N_2897,N_1288,N_1604);
nand U2898 (N_2898,N_1633,N_2245);
nand U2899 (N_2899,N_2361,N_2167);
xnor U2900 (N_2900,N_2111,N_2013);
xor U2901 (N_2901,N_2359,N_1581);
nand U2902 (N_2902,N_1569,N_2247);
xor U2903 (N_2903,N_2335,N_1934);
nor U2904 (N_2904,N_2117,N_1923);
nand U2905 (N_2905,N_1478,N_1834);
xnor U2906 (N_2906,N_2170,N_1816);
or U2907 (N_2907,N_2307,N_1998);
and U2908 (N_2908,N_2144,N_2272);
nor U2909 (N_2909,N_1874,N_2023);
and U2910 (N_2910,N_1455,N_2068);
nand U2911 (N_2911,N_1979,N_1437);
xor U2912 (N_2912,N_1430,N_1793);
and U2913 (N_2913,N_1949,N_2377);
and U2914 (N_2914,N_1456,N_1980);
and U2915 (N_2915,N_1807,N_2396);
nor U2916 (N_2916,N_2250,N_1344);
nor U2917 (N_2917,N_1916,N_1484);
nand U2918 (N_2918,N_1494,N_2373);
and U2919 (N_2919,N_1491,N_1703);
nor U2920 (N_2920,N_1845,N_1498);
xor U2921 (N_2921,N_2354,N_1388);
or U2922 (N_2922,N_2389,N_2295);
xnor U2923 (N_2923,N_1983,N_2153);
nand U2924 (N_2924,N_1329,N_2061);
or U2925 (N_2925,N_2336,N_1599);
and U2926 (N_2926,N_2293,N_1941);
xor U2927 (N_2927,N_1719,N_1556);
nand U2928 (N_2928,N_1451,N_1571);
nand U2929 (N_2929,N_1928,N_2002);
nor U2930 (N_2930,N_2204,N_1408);
or U2931 (N_2931,N_2075,N_2102);
or U2932 (N_2932,N_1959,N_1300);
nor U2933 (N_2933,N_1626,N_2368);
and U2934 (N_2934,N_1986,N_2060);
or U2935 (N_2935,N_2276,N_1827);
or U2936 (N_2936,N_1463,N_2210);
nor U2937 (N_2937,N_1886,N_1687);
nand U2938 (N_2938,N_1717,N_2041);
or U2939 (N_2939,N_2249,N_2233);
nand U2940 (N_2940,N_1572,N_1606);
xnor U2941 (N_2941,N_2313,N_2367);
nand U2942 (N_2942,N_1878,N_1374);
or U2943 (N_2943,N_1711,N_1619);
and U2944 (N_2944,N_1649,N_2005);
nand U2945 (N_2945,N_2342,N_1394);
xnor U2946 (N_2946,N_1354,N_1744);
nand U2947 (N_2947,N_1736,N_2371);
and U2948 (N_2948,N_1627,N_2112);
nand U2949 (N_2949,N_2184,N_2119);
or U2950 (N_2950,N_1266,N_1447);
nand U2951 (N_2951,N_1747,N_1254);
and U2952 (N_2952,N_1533,N_1526);
xor U2953 (N_2953,N_2054,N_2241);
or U2954 (N_2954,N_1917,N_1614);
nand U2955 (N_2955,N_2397,N_1956);
nand U2956 (N_2956,N_2252,N_1780);
nand U2957 (N_2957,N_1596,N_2177);
nand U2958 (N_2958,N_2106,N_1696);
nand U2959 (N_2959,N_1237,N_2229);
or U2960 (N_2960,N_1660,N_2058);
xnor U2961 (N_2961,N_1280,N_1386);
nor U2962 (N_2962,N_1469,N_1763);
or U2963 (N_2963,N_1582,N_1697);
or U2964 (N_2964,N_1224,N_2128);
nand U2965 (N_2965,N_2384,N_2080);
nand U2966 (N_2966,N_2324,N_1420);
or U2967 (N_2967,N_2176,N_2072);
nand U2968 (N_2968,N_2122,N_1647);
or U2969 (N_2969,N_1897,N_2113);
xnor U2970 (N_2970,N_1406,N_1773);
and U2971 (N_2971,N_2363,N_2087);
and U2972 (N_2972,N_1600,N_1549);
or U2973 (N_2973,N_2203,N_1228);
or U2974 (N_2974,N_1553,N_2040);
nand U2975 (N_2975,N_1403,N_1345);
or U2976 (N_2976,N_1693,N_1422);
nand U2977 (N_2977,N_2036,N_1337);
or U2978 (N_2978,N_1893,N_2202);
or U2979 (N_2979,N_1426,N_1318);
nor U2980 (N_2980,N_2278,N_1767);
or U2981 (N_2981,N_1327,N_1421);
xor U2982 (N_2982,N_1204,N_2280);
nor U2983 (N_2983,N_1639,N_2173);
nor U2984 (N_2984,N_1589,N_1528);
nand U2985 (N_2985,N_2279,N_2028);
or U2986 (N_2986,N_1262,N_2165);
nor U2987 (N_2987,N_1871,N_1423);
and U2988 (N_2988,N_2321,N_1863);
or U2989 (N_2989,N_1472,N_2120);
and U2990 (N_2990,N_2044,N_1238);
nor U2991 (N_2991,N_2207,N_2231);
nor U2992 (N_2992,N_1657,N_1504);
or U2993 (N_2993,N_1399,N_1608);
nor U2994 (N_2994,N_1892,N_2320);
xor U2995 (N_2995,N_2299,N_2126);
and U2996 (N_2996,N_2381,N_2341);
or U2997 (N_2997,N_1961,N_1313);
xnor U2998 (N_2998,N_1790,N_2098);
nand U2999 (N_2999,N_2149,N_2121);
xor U3000 (N_3000,N_1532,N_1565);
and U3001 (N_3001,N_1734,N_2061);
xor U3002 (N_3002,N_2392,N_1433);
or U3003 (N_3003,N_2251,N_1843);
nor U3004 (N_3004,N_2387,N_1338);
xor U3005 (N_3005,N_2075,N_2088);
and U3006 (N_3006,N_2292,N_1565);
and U3007 (N_3007,N_1543,N_1489);
nor U3008 (N_3008,N_2088,N_1369);
xnor U3009 (N_3009,N_1948,N_1380);
or U3010 (N_3010,N_1641,N_2027);
nor U3011 (N_3011,N_1755,N_2039);
and U3012 (N_3012,N_1614,N_2392);
and U3013 (N_3013,N_1250,N_1294);
and U3014 (N_3014,N_2041,N_1850);
nor U3015 (N_3015,N_1627,N_1986);
nand U3016 (N_3016,N_1521,N_2056);
nand U3017 (N_3017,N_1275,N_1571);
or U3018 (N_3018,N_2307,N_1514);
or U3019 (N_3019,N_2324,N_1733);
nand U3020 (N_3020,N_1919,N_2200);
nand U3021 (N_3021,N_1262,N_1368);
nand U3022 (N_3022,N_1878,N_1589);
xor U3023 (N_3023,N_2130,N_1838);
or U3024 (N_3024,N_1866,N_1943);
or U3025 (N_3025,N_2068,N_2331);
nand U3026 (N_3026,N_1868,N_1728);
and U3027 (N_3027,N_1351,N_2019);
xor U3028 (N_3028,N_2059,N_1973);
xor U3029 (N_3029,N_2099,N_1885);
nand U3030 (N_3030,N_1530,N_1716);
nand U3031 (N_3031,N_1323,N_1578);
xor U3032 (N_3032,N_1563,N_2222);
and U3033 (N_3033,N_1200,N_1587);
nor U3034 (N_3034,N_1439,N_1330);
nor U3035 (N_3035,N_2052,N_1921);
nor U3036 (N_3036,N_1810,N_1493);
and U3037 (N_3037,N_2102,N_1386);
and U3038 (N_3038,N_2306,N_1723);
nand U3039 (N_3039,N_1966,N_1480);
and U3040 (N_3040,N_1337,N_1622);
xor U3041 (N_3041,N_1709,N_2329);
nand U3042 (N_3042,N_1308,N_1496);
nor U3043 (N_3043,N_2041,N_1347);
nor U3044 (N_3044,N_2292,N_2339);
nor U3045 (N_3045,N_1533,N_2228);
nand U3046 (N_3046,N_1826,N_1563);
nor U3047 (N_3047,N_2006,N_1325);
and U3048 (N_3048,N_2127,N_2334);
and U3049 (N_3049,N_1223,N_1631);
nand U3050 (N_3050,N_2351,N_1287);
or U3051 (N_3051,N_1679,N_1311);
and U3052 (N_3052,N_2219,N_1589);
xnor U3053 (N_3053,N_2121,N_2285);
xnor U3054 (N_3054,N_1661,N_2293);
nor U3055 (N_3055,N_2093,N_2269);
and U3056 (N_3056,N_1213,N_1278);
xor U3057 (N_3057,N_1261,N_1783);
nand U3058 (N_3058,N_1802,N_2359);
nand U3059 (N_3059,N_1410,N_1503);
nor U3060 (N_3060,N_2298,N_1559);
xor U3061 (N_3061,N_1461,N_1618);
and U3062 (N_3062,N_1615,N_1571);
or U3063 (N_3063,N_2185,N_1939);
nor U3064 (N_3064,N_1756,N_1367);
nor U3065 (N_3065,N_1608,N_1937);
nand U3066 (N_3066,N_1680,N_1712);
xnor U3067 (N_3067,N_2267,N_1997);
and U3068 (N_3068,N_2111,N_2038);
nor U3069 (N_3069,N_2103,N_1355);
or U3070 (N_3070,N_2354,N_1977);
and U3071 (N_3071,N_2206,N_2294);
nand U3072 (N_3072,N_1308,N_1801);
or U3073 (N_3073,N_1305,N_2367);
and U3074 (N_3074,N_1243,N_2375);
xor U3075 (N_3075,N_2270,N_1217);
and U3076 (N_3076,N_1895,N_1533);
or U3077 (N_3077,N_1623,N_1959);
and U3078 (N_3078,N_1500,N_2382);
and U3079 (N_3079,N_1820,N_1764);
and U3080 (N_3080,N_1419,N_1433);
or U3081 (N_3081,N_2053,N_1409);
nor U3082 (N_3082,N_1585,N_1413);
and U3083 (N_3083,N_1781,N_1780);
nor U3084 (N_3084,N_1359,N_2034);
and U3085 (N_3085,N_2096,N_2289);
or U3086 (N_3086,N_2277,N_2221);
nor U3087 (N_3087,N_1562,N_2008);
and U3088 (N_3088,N_2366,N_1354);
nor U3089 (N_3089,N_2194,N_1392);
or U3090 (N_3090,N_1435,N_2297);
nand U3091 (N_3091,N_2298,N_2365);
nand U3092 (N_3092,N_1744,N_1965);
or U3093 (N_3093,N_1859,N_2141);
xnor U3094 (N_3094,N_2316,N_2299);
and U3095 (N_3095,N_1985,N_2174);
nand U3096 (N_3096,N_1707,N_2026);
and U3097 (N_3097,N_1285,N_1886);
nor U3098 (N_3098,N_2193,N_2362);
and U3099 (N_3099,N_1203,N_1842);
or U3100 (N_3100,N_1255,N_2093);
and U3101 (N_3101,N_1322,N_1776);
or U3102 (N_3102,N_2006,N_1432);
or U3103 (N_3103,N_1697,N_1542);
xor U3104 (N_3104,N_1626,N_1484);
and U3105 (N_3105,N_1478,N_1709);
xor U3106 (N_3106,N_1381,N_1368);
or U3107 (N_3107,N_2183,N_1683);
nand U3108 (N_3108,N_1217,N_1455);
or U3109 (N_3109,N_1899,N_1679);
or U3110 (N_3110,N_1931,N_2066);
xnor U3111 (N_3111,N_2398,N_2314);
nand U3112 (N_3112,N_1611,N_2299);
nor U3113 (N_3113,N_1273,N_1933);
nor U3114 (N_3114,N_1769,N_1687);
xnor U3115 (N_3115,N_1773,N_2287);
nor U3116 (N_3116,N_1883,N_1213);
nor U3117 (N_3117,N_2199,N_1461);
xnor U3118 (N_3118,N_1655,N_1800);
or U3119 (N_3119,N_2279,N_1383);
nor U3120 (N_3120,N_1745,N_1697);
and U3121 (N_3121,N_1900,N_2178);
nor U3122 (N_3122,N_1954,N_2022);
and U3123 (N_3123,N_1227,N_1909);
or U3124 (N_3124,N_1528,N_2103);
nor U3125 (N_3125,N_1783,N_2159);
and U3126 (N_3126,N_1781,N_2007);
nand U3127 (N_3127,N_1674,N_1503);
and U3128 (N_3128,N_1767,N_2333);
or U3129 (N_3129,N_2051,N_1714);
and U3130 (N_3130,N_1289,N_1841);
xnor U3131 (N_3131,N_1719,N_2014);
nor U3132 (N_3132,N_1585,N_1643);
xor U3133 (N_3133,N_1858,N_2315);
nand U3134 (N_3134,N_2393,N_1476);
and U3135 (N_3135,N_1607,N_1279);
or U3136 (N_3136,N_1291,N_1212);
nand U3137 (N_3137,N_1924,N_1540);
nor U3138 (N_3138,N_1915,N_2363);
and U3139 (N_3139,N_1367,N_1694);
and U3140 (N_3140,N_1228,N_1378);
or U3141 (N_3141,N_1419,N_2184);
xnor U3142 (N_3142,N_1907,N_1998);
nand U3143 (N_3143,N_1913,N_1332);
xor U3144 (N_3144,N_1531,N_1833);
nor U3145 (N_3145,N_1672,N_1520);
and U3146 (N_3146,N_2323,N_1478);
and U3147 (N_3147,N_1224,N_1217);
or U3148 (N_3148,N_2128,N_2348);
nor U3149 (N_3149,N_1380,N_1781);
nor U3150 (N_3150,N_1649,N_1955);
nand U3151 (N_3151,N_2123,N_1648);
xnor U3152 (N_3152,N_2101,N_2127);
nor U3153 (N_3153,N_1690,N_1798);
or U3154 (N_3154,N_2272,N_1916);
nand U3155 (N_3155,N_2210,N_1505);
or U3156 (N_3156,N_1808,N_2328);
and U3157 (N_3157,N_1310,N_1419);
nand U3158 (N_3158,N_2050,N_1749);
xor U3159 (N_3159,N_1625,N_1924);
and U3160 (N_3160,N_1593,N_2208);
and U3161 (N_3161,N_1645,N_1504);
and U3162 (N_3162,N_1783,N_1445);
or U3163 (N_3163,N_1206,N_2125);
or U3164 (N_3164,N_2208,N_2365);
nor U3165 (N_3165,N_1415,N_2396);
or U3166 (N_3166,N_1304,N_1213);
and U3167 (N_3167,N_2143,N_2121);
or U3168 (N_3168,N_1661,N_2111);
or U3169 (N_3169,N_1549,N_2072);
and U3170 (N_3170,N_1208,N_1989);
nor U3171 (N_3171,N_1496,N_2333);
nand U3172 (N_3172,N_2362,N_2017);
and U3173 (N_3173,N_2145,N_1951);
xor U3174 (N_3174,N_2255,N_1778);
nand U3175 (N_3175,N_1407,N_1793);
xnor U3176 (N_3176,N_2083,N_1678);
and U3177 (N_3177,N_1924,N_1970);
or U3178 (N_3178,N_1384,N_1658);
xor U3179 (N_3179,N_2381,N_2084);
xor U3180 (N_3180,N_2374,N_1893);
nor U3181 (N_3181,N_2101,N_1300);
and U3182 (N_3182,N_2211,N_2133);
and U3183 (N_3183,N_1502,N_1929);
xor U3184 (N_3184,N_1309,N_1997);
xor U3185 (N_3185,N_1878,N_1791);
nor U3186 (N_3186,N_1455,N_1450);
nor U3187 (N_3187,N_1416,N_2331);
nor U3188 (N_3188,N_1721,N_1573);
nand U3189 (N_3189,N_2126,N_2178);
or U3190 (N_3190,N_2119,N_1451);
or U3191 (N_3191,N_2215,N_2279);
nand U3192 (N_3192,N_1952,N_1495);
or U3193 (N_3193,N_2032,N_1931);
nand U3194 (N_3194,N_1646,N_2186);
or U3195 (N_3195,N_1351,N_1698);
and U3196 (N_3196,N_1862,N_1470);
nand U3197 (N_3197,N_2336,N_2013);
xnor U3198 (N_3198,N_1626,N_1342);
xnor U3199 (N_3199,N_1578,N_1444);
xnor U3200 (N_3200,N_1578,N_1870);
nor U3201 (N_3201,N_1599,N_1712);
xor U3202 (N_3202,N_1222,N_1859);
nor U3203 (N_3203,N_1399,N_1413);
nor U3204 (N_3204,N_2355,N_1861);
nand U3205 (N_3205,N_1288,N_1874);
xor U3206 (N_3206,N_1334,N_2201);
nand U3207 (N_3207,N_1840,N_1806);
nand U3208 (N_3208,N_1836,N_1679);
or U3209 (N_3209,N_1976,N_2109);
xor U3210 (N_3210,N_1925,N_1536);
and U3211 (N_3211,N_1930,N_1802);
or U3212 (N_3212,N_1888,N_1728);
and U3213 (N_3213,N_2181,N_2279);
xor U3214 (N_3214,N_1911,N_1920);
or U3215 (N_3215,N_2082,N_1256);
and U3216 (N_3216,N_1594,N_2359);
or U3217 (N_3217,N_1440,N_2363);
nand U3218 (N_3218,N_2231,N_1385);
xor U3219 (N_3219,N_1325,N_1595);
or U3220 (N_3220,N_1636,N_1296);
or U3221 (N_3221,N_1995,N_1929);
and U3222 (N_3222,N_1984,N_1822);
or U3223 (N_3223,N_2144,N_1878);
and U3224 (N_3224,N_1803,N_2295);
xnor U3225 (N_3225,N_1960,N_1408);
nand U3226 (N_3226,N_1972,N_2375);
nor U3227 (N_3227,N_1533,N_1386);
and U3228 (N_3228,N_1839,N_2206);
nand U3229 (N_3229,N_1463,N_2258);
or U3230 (N_3230,N_1304,N_1796);
nor U3231 (N_3231,N_1620,N_2282);
nor U3232 (N_3232,N_1217,N_2089);
or U3233 (N_3233,N_2288,N_2150);
xor U3234 (N_3234,N_1218,N_1648);
xnor U3235 (N_3235,N_1411,N_1999);
nor U3236 (N_3236,N_1506,N_1675);
nor U3237 (N_3237,N_1727,N_1726);
and U3238 (N_3238,N_2058,N_2197);
xor U3239 (N_3239,N_1542,N_1622);
and U3240 (N_3240,N_1234,N_1519);
nand U3241 (N_3241,N_1907,N_2165);
nor U3242 (N_3242,N_1678,N_2158);
nand U3243 (N_3243,N_2128,N_2052);
and U3244 (N_3244,N_2296,N_1419);
and U3245 (N_3245,N_1588,N_2305);
or U3246 (N_3246,N_2077,N_1394);
and U3247 (N_3247,N_2082,N_1892);
xnor U3248 (N_3248,N_1623,N_1604);
nor U3249 (N_3249,N_2269,N_1280);
or U3250 (N_3250,N_1563,N_1642);
xnor U3251 (N_3251,N_2269,N_1599);
or U3252 (N_3252,N_1973,N_2253);
nand U3253 (N_3253,N_2297,N_2349);
xnor U3254 (N_3254,N_1841,N_2318);
and U3255 (N_3255,N_1385,N_2122);
or U3256 (N_3256,N_2333,N_1537);
or U3257 (N_3257,N_1532,N_2072);
xnor U3258 (N_3258,N_1203,N_1328);
nand U3259 (N_3259,N_1863,N_2112);
nor U3260 (N_3260,N_1743,N_1332);
nand U3261 (N_3261,N_1701,N_1644);
nand U3262 (N_3262,N_1232,N_2324);
nor U3263 (N_3263,N_1294,N_1526);
and U3264 (N_3264,N_1232,N_1376);
and U3265 (N_3265,N_2305,N_1753);
and U3266 (N_3266,N_1261,N_1692);
nand U3267 (N_3267,N_2091,N_1932);
and U3268 (N_3268,N_1404,N_1385);
xor U3269 (N_3269,N_2039,N_1628);
xor U3270 (N_3270,N_1920,N_1251);
xor U3271 (N_3271,N_1771,N_1342);
xnor U3272 (N_3272,N_1756,N_2147);
or U3273 (N_3273,N_2125,N_2167);
nor U3274 (N_3274,N_2309,N_2215);
or U3275 (N_3275,N_1619,N_1772);
nor U3276 (N_3276,N_2116,N_1874);
or U3277 (N_3277,N_2035,N_2057);
and U3278 (N_3278,N_2170,N_1586);
xor U3279 (N_3279,N_1226,N_2045);
or U3280 (N_3280,N_2027,N_1404);
nand U3281 (N_3281,N_2234,N_1627);
xor U3282 (N_3282,N_1966,N_2211);
xnor U3283 (N_3283,N_2388,N_1620);
nand U3284 (N_3284,N_1932,N_1646);
nand U3285 (N_3285,N_1764,N_1749);
nor U3286 (N_3286,N_1641,N_2158);
and U3287 (N_3287,N_1620,N_1281);
and U3288 (N_3288,N_1502,N_1467);
and U3289 (N_3289,N_1405,N_1208);
or U3290 (N_3290,N_1582,N_1542);
xnor U3291 (N_3291,N_2164,N_1789);
or U3292 (N_3292,N_2167,N_2251);
nor U3293 (N_3293,N_2232,N_1290);
nor U3294 (N_3294,N_1264,N_2232);
xnor U3295 (N_3295,N_1301,N_1337);
and U3296 (N_3296,N_1717,N_1928);
or U3297 (N_3297,N_1887,N_1497);
nor U3298 (N_3298,N_1999,N_1630);
and U3299 (N_3299,N_1943,N_1603);
or U3300 (N_3300,N_2129,N_2089);
nand U3301 (N_3301,N_1943,N_1888);
xor U3302 (N_3302,N_2067,N_2159);
nand U3303 (N_3303,N_1396,N_1572);
and U3304 (N_3304,N_1849,N_1543);
and U3305 (N_3305,N_2068,N_1821);
nand U3306 (N_3306,N_1319,N_1330);
nor U3307 (N_3307,N_2125,N_1281);
nor U3308 (N_3308,N_2171,N_1459);
nor U3309 (N_3309,N_1982,N_1923);
or U3310 (N_3310,N_2361,N_2113);
nand U3311 (N_3311,N_1356,N_1251);
xor U3312 (N_3312,N_2087,N_2349);
nor U3313 (N_3313,N_1878,N_1289);
nand U3314 (N_3314,N_2228,N_1823);
nand U3315 (N_3315,N_2273,N_2275);
nor U3316 (N_3316,N_1420,N_1380);
or U3317 (N_3317,N_1692,N_1759);
nor U3318 (N_3318,N_1288,N_1483);
or U3319 (N_3319,N_1836,N_2326);
and U3320 (N_3320,N_2049,N_1548);
and U3321 (N_3321,N_1220,N_1425);
xnor U3322 (N_3322,N_1995,N_1345);
and U3323 (N_3323,N_2100,N_2117);
nand U3324 (N_3324,N_1428,N_1377);
xnor U3325 (N_3325,N_1745,N_1969);
nand U3326 (N_3326,N_1600,N_1250);
nand U3327 (N_3327,N_2174,N_2022);
xnor U3328 (N_3328,N_2059,N_1461);
xnor U3329 (N_3329,N_1271,N_2303);
xnor U3330 (N_3330,N_2128,N_1960);
nor U3331 (N_3331,N_1459,N_1820);
nand U3332 (N_3332,N_1754,N_2308);
or U3333 (N_3333,N_2296,N_1754);
nor U3334 (N_3334,N_1350,N_2027);
nand U3335 (N_3335,N_1959,N_2386);
and U3336 (N_3336,N_2371,N_1318);
or U3337 (N_3337,N_2281,N_1691);
nor U3338 (N_3338,N_2233,N_1757);
nor U3339 (N_3339,N_1887,N_1805);
or U3340 (N_3340,N_1616,N_1816);
nand U3341 (N_3341,N_2113,N_1279);
and U3342 (N_3342,N_1455,N_2260);
xnor U3343 (N_3343,N_2367,N_1844);
nand U3344 (N_3344,N_1505,N_1420);
xnor U3345 (N_3345,N_1681,N_1846);
and U3346 (N_3346,N_1573,N_1941);
and U3347 (N_3347,N_2317,N_2135);
xnor U3348 (N_3348,N_1390,N_1938);
nand U3349 (N_3349,N_2162,N_2156);
nor U3350 (N_3350,N_2123,N_2215);
and U3351 (N_3351,N_1711,N_2297);
and U3352 (N_3352,N_2255,N_1364);
and U3353 (N_3353,N_2133,N_1536);
nand U3354 (N_3354,N_1745,N_2379);
and U3355 (N_3355,N_1641,N_1572);
or U3356 (N_3356,N_1281,N_1537);
nand U3357 (N_3357,N_1641,N_1212);
xor U3358 (N_3358,N_1923,N_1325);
and U3359 (N_3359,N_1697,N_2393);
or U3360 (N_3360,N_1472,N_1697);
or U3361 (N_3361,N_1636,N_1280);
nand U3362 (N_3362,N_2132,N_1780);
nor U3363 (N_3363,N_1229,N_1541);
nand U3364 (N_3364,N_2068,N_1977);
nand U3365 (N_3365,N_1384,N_2178);
nor U3366 (N_3366,N_2390,N_1314);
xor U3367 (N_3367,N_1590,N_2309);
nor U3368 (N_3368,N_1613,N_1722);
xor U3369 (N_3369,N_2238,N_1382);
nand U3370 (N_3370,N_1341,N_1617);
nand U3371 (N_3371,N_2086,N_1755);
nand U3372 (N_3372,N_1942,N_1286);
nand U3373 (N_3373,N_1301,N_1824);
or U3374 (N_3374,N_2110,N_2198);
or U3375 (N_3375,N_2265,N_1383);
nor U3376 (N_3376,N_2227,N_2246);
and U3377 (N_3377,N_1719,N_2062);
or U3378 (N_3378,N_1223,N_1983);
or U3379 (N_3379,N_1969,N_1624);
xor U3380 (N_3380,N_1585,N_1934);
or U3381 (N_3381,N_2122,N_2394);
and U3382 (N_3382,N_1710,N_2314);
nand U3383 (N_3383,N_1848,N_2207);
nand U3384 (N_3384,N_1910,N_2041);
nand U3385 (N_3385,N_2132,N_1380);
nand U3386 (N_3386,N_1593,N_1273);
or U3387 (N_3387,N_2375,N_2151);
or U3388 (N_3388,N_2081,N_1362);
nor U3389 (N_3389,N_1538,N_1331);
nand U3390 (N_3390,N_1332,N_1469);
nor U3391 (N_3391,N_1486,N_1481);
nand U3392 (N_3392,N_1914,N_1942);
or U3393 (N_3393,N_1939,N_1701);
or U3394 (N_3394,N_2215,N_1240);
nor U3395 (N_3395,N_1900,N_2397);
xnor U3396 (N_3396,N_1367,N_1681);
nand U3397 (N_3397,N_2091,N_2384);
and U3398 (N_3398,N_1280,N_1949);
nand U3399 (N_3399,N_1489,N_1796);
xnor U3400 (N_3400,N_1598,N_1836);
xor U3401 (N_3401,N_1361,N_1312);
xnor U3402 (N_3402,N_1459,N_1519);
nand U3403 (N_3403,N_2179,N_2161);
or U3404 (N_3404,N_2123,N_2316);
or U3405 (N_3405,N_1911,N_2139);
xnor U3406 (N_3406,N_1804,N_1949);
nand U3407 (N_3407,N_1769,N_1538);
nor U3408 (N_3408,N_1904,N_2032);
nand U3409 (N_3409,N_2004,N_2182);
nand U3410 (N_3410,N_2391,N_2352);
or U3411 (N_3411,N_2257,N_2088);
and U3412 (N_3412,N_1572,N_1578);
or U3413 (N_3413,N_1240,N_1493);
xor U3414 (N_3414,N_2222,N_1676);
or U3415 (N_3415,N_2222,N_2202);
and U3416 (N_3416,N_2009,N_1539);
xor U3417 (N_3417,N_2323,N_1522);
and U3418 (N_3418,N_1607,N_1473);
and U3419 (N_3419,N_1352,N_2140);
xnor U3420 (N_3420,N_2399,N_1342);
or U3421 (N_3421,N_2387,N_2114);
xor U3422 (N_3422,N_2383,N_1803);
or U3423 (N_3423,N_1946,N_2190);
nor U3424 (N_3424,N_2124,N_1886);
and U3425 (N_3425,N_2255,N_1739);
or U3426 (N_3426,N_1759,N_2302);
and U3427 (N_3427,N_1970,N_2184);
nand U3428 (N_3428,N_2221,N_1921);
xnor U3429 (N_3429,N_1503,N_2397);
nor U3430 (N_3430,N_1454,N_2275);
nor U3431 (N_3431,N_2309,N_1312);
nand U3432 (N_3432,N_1772,N_1633);
xor U3433 (N_3433,N_2390,N_2074);
or U3434 (N_3434,N_1525,N_1724);
or U3435 (N_3435,N_2274,N_1521);
nor U3436 (N_3436,N_1384,N_1784);
or U3437 (N_3437,N_2343,N_1694);
nand U3438 (N_3438,N_1854,N_2298);
nor U3439 (N_3439,N_2368,N_2285);
and U3440 (N_3440,N_1489,N_1810);
or U3441 (N_3441,N_1413,N_2160);
nand U3442 (N_3442,N_2296,N_1261);
nor U3443 (N_3443,N_2323,N_1525);
and U3444 (N_3444,N_1801,N_1872);
nor U3445 (N_3445,N_2338,N_1981);
and U3446 (N_3446,N_2345,N_1369);
nor U3447 (N_3447,N_2312,N_2040);
xor U3448 (N_3448,N_1828,N_1862);
and U3449 (N_3449,N_2260,N_1996);
nand U3450 (N_3450,N_1774,N_1972);
nor U3451 (N_3451,N_1920,N_1221);
nand U3452 (N_3452,N_1355,N_1677);
or U3453 (N_3453,N_2190,N_2171);
and U3454 (N_3454,N_1793,N_1294);
nor U3455 (N_3455,N_2054,N_2101);
or U3456 (N_3456,N_2062,N_2126);
xor U3457 (N_3457,N_1718,N_1739);
xnor U3458 (N_3458,N_2376,N_1687);
and U3459 (N_3459,N_2351,N_1811);
or U3460 (N_3460,N_1576,N_1215);
and U3461 (N_3461,N_2382,N_2052);
xor U3462 (N_3462,N_1354,N_2377);
xor U3463 (N_3463,N_1868,N_1443);
nand U3464 (N_3464,N_1482,N_1234);
nand U3465 (N_3465,N_1224,N_2107);
xnor U3466 (N_3466,N_2169,N_2082);
nor U3467 (N_3467,N_1891,N_1625);
nor U3468 (N_3468,N_1606,N_1331);
nor U3469 (N_3469,N_1558,N_1490);
xor U3470 (N_3470,N_2110,N_1316);
xor U3471 (N_3471,N_1200,N_2242);
nor U3472 (N_3472,N_2231,N_1511);
nor U3473 (N_3473,N_1719,N_2319);
nand U3474 (N_3474,N_1902,N_1226);
or U3475 (N_3475,N_2068,N_1215);
nand U3476 (N_3476,N_1863,N_2366);
or U3477 (N_3477,N_1719,N_1588);
nor U3478 (N_3478,N_1865,N_2253);
or U3479 (N_3479,N_1877,N_1368);
nand U3480 (N_3480,N_1316,N_1393);
xnor U3481 (N_3481,N_1704,N_2229);
nor U3482 (N_3482,N_1663,N_1348);
nand U3483 (N_3483,N_1415,N_1341);
or U3484 (N_3484,N_1451,N_2345);
xor U3485 (N_3485,N_1252,N_1455);
or U3486 (N_3486,N_1219,N_1684);
nand U3487 (N_3487,N_1608,N_2094);
nand U3488 (N_3488,N_2043,N_2249);
and U3489 (N_3489,N_1315,N_2167);
or U3490 (N_3490,N_1833,N_1850);
nor U3491 (N_3491,N_1500,N_1996);
xor U3492 (N_3492,N_1445,N_1678);
xnor U3493 (N_3493,N_1516,N_2228);
nand U3494 (N_3494,N_1723,N_1512);
nor U3495 (N_3495,N_1778,N_1642);
or U3496 (N_3496,N_1729,N_2230);
nand U3497 (N_3497,N_2145,N_2124);
xor U3498 (N_3498,N_2149,N_1712);
xor U3499 (N_3499,N_1634,N_1210);
and U3500 (N_3500,N_2132,N_1761);
nor U3501 (N_3501,N_1398,N_1520);
and U3502 (N_3502,N_1446,N_1271);
xor U3503 (N_3503,N_2259,N_1423);
and U3504 (N_3504,N_1404,N_1559);
and U3505 (N_3505,N_1859,N_1958);
and U3506 (N_3506,N_2235,N_1484);
or U3507 (N_3507,N_1383,N_2083);
and U3508 (N_3508,N_2011,N_1204);
and U3509 (N_3509,N_2324,N_1579);
and U3510 (N_3510,N_1747,N_2114);
or U3511 (N_3511,N_1697,N_1903);
or U3512 (N_3512,N_1713,N_1467);
nor U3513 (N_3513,N_1658,N_2394);
and U3514 (N_3514,N_1375,N_1527);
nand U3515 (N_3515,N_1238,N_2132);
or U3516 (N_3516,N_1643,N_2285);
or U3517 (N_3517,N_1635,N_1588);
and U3518 (N_3518,N_1201,N_1816);
and U3519 (N_3519,N_1270,N_2358);
and U3520 (N_3520,N_2390,N_2020);
and U3521 (N_3521,N_1413,N_1843);
nor U3522 (N_3522,N_2250,N_1366);
xor U3523 (N_3523,N_2158,N_1707);
and U3524 (N_3524,N_2207,N_2160);
and U3525 (N_3525,N_2276,N_1808);
or U3526 (N_3526,N_1765,N_1743);
and U3527 (N_3527,N_2389,N_2219);
or U3528 (N_3528,N_1590,N_1396);
nand U3529 (N_3529,N_1555,N_2345);
or U3530 (N_3530,N_2347,N_2274);
or U3531 (N_3531,N_2372,N_1653);
nor U3532 (N_3532,N_1467,N_1798);
xnor U3533 (N_3533,N_1698,N_1799);
nand U3534 (N_3534,N_1884,N_1456);
xnor U3535 (N_3535,N_1465,N_1575);
nor U3536 (N_3536,N_1287,N_1690);
nand U3537 (N_3537,N_1864,N_1265);
xnor U3538 (N_3538,N_2274,N_1567);
or U3539 (N_3539,N_1578,N_1319);
or U3540 (N_3540,N_1412,N_2056);
and U3541 (N_3541,N_2313,N_1867);
xnor U3542 (N_3542,N_2160,N_1650);
nor U3543 (N_3543,N_1532,N_1296);
nor U3544 (N_3544,N_1495,N_2045);
and U3545 (N_3545,N_2098,N_1475);
xor U3546 (N_3546,N_1541,N_1572);
xnor U3547 (N_3547,N_2309,N_2281);
nand U3548 (N_3548,N_2181,N_2052);
xnor U3549 (N_3549,N_1444,N_1692);
xor U3550 (N_3550,N_2111,N_1231);
nand U3551 (N_3551,N_1593,N_1698);
or U3552 (N_3552,N_2348,N_2079);
xnor U3553 (N_3553,N_2205,N_1896);
nand U3554 (N_3554,N_2355,N_1895);
xnor U3555 (N_3555,N_1781,N_1750);
xnor U3556 (N_3556,N_1301,N_2054);
nor U3557 (N_3557,N_1378,N_1816);
and U3558 (N_3558,N_1486,N_1970);
xnor U3559 (N_3559,N_2237,N_1679);
or U3560 (N_3560,N_1295,N_1237);
xor U3561 (N_3561,N_1722,N_1840);
nand U3562 (N_3562,N_2062,N_2174);
or U3563 (N_3563,N_2310,N_1338);
nand U3564 (N_3564,N_1542,N_1715);
and U3565 (N_3565,N_1368,N_2141);
nor U3566 (N_3566,N_1997,N_2265);
and U3567 (N_3567,N_2198,N_2243);
xnor U3568 (N_3568,N_2179,N_2125);
and U3569 (N_3569,N_1399,N_2252);
nand U3570 (N_3570,N_1893,N_1694);
xnor U3571 (N_3571,N_1875,N_2191);
xnor U3572 (N_3572,N_1836,N_1426);
nor U3573 (N_3573,N_1595,N_2326);
nor U3574 (N_3574,N_1215,N_2192);
or U3575 (N_3575,N_1391,N_1766);
or U3576 (N_3576,N_1495,N_1338);
nand U3577 (N_3577,N_1391,N_2082);
xnor U3578 (N_3578,N_1631,N_1333);
nor U3579 (N_3579,N_2036,N_1343);
and U3580 (N_3580,N_2186,N_1652);
and U3581 (N_3581,N_2028,N_1735);
nor U3582 (N_3582,N_2195,N_2365);
nand U3583 (N_3583,N_1746,N_1943);
nor U3584 (N_3584,N_1491,N_1387);
and U3585 (N_3585,N_1484,N_2369);
and U3586 (N_3586,N_1520,N_1609);
xnor U3587 (N_3587,N_1611,N_1208);
xnor U3588 (N_3588,N_1429,N_1446);
xor U3589 (N_3589,N_1439,N_1597);
and U3590 (N_3590,N_1552,N_1235);
or U3591 (N_3591,N_1903,N_2115);
xnor U3592 (N_3592,N_1508,N_1487);
nand U3593 (N_3593,N_2028,N_2385);
or U3594 (N_3594,N_1570,N_1329);
or U3595 (N_3595,N_2045,N_1362);
nand U3596 (N_3596,N_1387,N_1563);
and U3597 (N_3597,N_1736,N_1565);
and U3598 (N_3598,N_1439,N_1998);
nand U3599 (N_3599,N_1936,N_2372);
nand U3600 (N_3600,N_2587,N_3565);
nor U3601 (N_3601,N_3347,N_2921);
nand U3602 (N_3602,N_2554,N_3065);
or U3603 (N_3603,N_2864,N_2481);
and U3604 (N_3604,N_3342,N_3529);
and U3605 (N_3605,N_3358,N_3404);
or U3606 (N_3606,N_2793,N_3010);
or U3607 (N_3607,N_3353,N_3526);
or U3608 (N_3608,N_2953,N_2958);
nor U3609 (N_3609,N_2704,N_2705);
or U3610 (N_3610,N_3287,N_2829);
nor U3611 (N_3611,N_2780,N_3471);
nand U3612 (N_3612,N_3475,N_2421);
nor U3613 (N_3613,N_3171,N_3382);
nand U3614 (N_3614,N_2440,N_3024);
and U3615 (N_3615,N_2878,N_2612);
or U3616 (N_3616,N_3399,N_2451);
or U3617 (N_3617,N_3088,N_3491);
nor U3618 (N_3618,N_2960,N_2867);
nor U3619 (N_3619,N_3325,N_3551);
or U3620 (N_3620,N_2431,N_2491);
nand U3621 (N_3621,N_2962,N_2606);
nand U3622 (N_3622,N_2846,N_3022);
xnor U3623 (N_3623,N_3313,N_3137);
and U3624 (N_3624,N_3219,N_3444);
nand U3625 (N_3625,N_2795,N_3032);
or U3626 (N_3626,N_3135,N_2540);
or U3627 (N_3627,N_2418,N_2403);
and U3628 (N_3628,N_3069,N_3510);
xor U3629 (N_3629,N_3552,N_3216);
xor U3630 (N_3630,N_3285,N_3322);
or U3631 (N_3631,N_2954,N_3321);
nor U3632 (N_3632,N_2879,N_2836);
nand U3633 (N_3633,N_3450,N_2724);
or U3634 (N_3634,N_3006,N_3407);
nand U3635 (N_3635,N_2433,N_3258);
and U3636 (N_3636,N_3060,N_2690);
nand U3637 (N_3637,N_2955,N_3581);
nand U3638 (N_3638,N_2735,N_3376);
or U3639 (N_3639,N_3091,N_3563);
nand U3640 (N_3640,N_2872,N_2676);
xor U3641 (N_3641,N_3078,N_3122);
and U3642 (N_3642,N_3441,N_2607);
and U3643 (N_3643,N_2579,N_2956);
xor U3644 (N_3644,N_2972,N_2966);
or U3645 (N_3645,N_3294,N_3072);
xnor U3646 (N_3646,N_2450,N_3596);
or U3647 (N_3647,N_3261,N_2664);
xnor U3648 (N_3648,N_3493,N_3089);
nand U3649 (N_3649,N_2764,N_3394);
nand U3650 (N_3650,N_3405,N_3220);
nand U3651 (N_3651,N_2539,N_2455);
nor U3652 (N_3652,N_2681,N_3369);
xor U3653 (N_3653,N_3474,N_2636);
or U3654 (N_3654,N_3046,N_3571);
and U3655 (N_3655,N_3501,N_3239);
nand U3656 (N_3656,N_2558,N_3438);
xnor U3657 (N_3657,N_2977,N_3517);
and U3658 (N_3658,N_2760,N_2738);
nand U3659 (N_3659,N_2801,N_2550);
nand U3660 (N_3660,N_3011,N_2987);
or U3661 (N_3661,N_3243,N_2856);
or U3662 (N_3662,N_3201,N_2474);
nand U3663 (N_3663,N_2400,N_2447);
and U3664 (N_3664,N_3139,N_3590);
nor U3665 (N_3665,N_3092,N_3016);
and U3666 (N_3666,N_3275,N_2901);
nor U3667 (N_3667,N_3598,N_2434);
xnor U3668 (N_3668,N_2976,N_2970);
nand U3669 (N_3669,N_3231,N_3109);
or U3670 (N_3670,N_2556,N_2682);
or U3671 (N_3671,N_2832,N_3013);
xor U3672 (N_3672,N_3211,N_3225);
nor U3673 (N_3673,N_2952,N_3550);
and U3674 (N_3674,N_3415,N_2610);
or U3675 (N_3675,N_2797,N_3164);
or U3676 (N_3676,N_3026,N_3064);
and U3677 (N_3677,N_2565,N_2930);
or U3678 (N_3678,N_3177,N_3393);
xor U3679 (N_3679,N_2898,N_3311);
and U3680 (N_3680,N_2806,N_2686);
nand U3681 (N_3681,N_3421,N_3543);
nand U3682 (N_3682,N_2635,N_3435);
xnor U3683 (N_3683,N_2571,N_3279);
xnor U3684 (N_3684,N_2799,N_2895);
xor U3685 (N_3685,N_3038,N_2880);
nor U3686 (N_3686,N_2726,N_3318);
and U3687 (N_3687,N_2849,N_2733);
or U3688 (N_3688,N_2412,N_2893);
or U3689 (N_3689,N_2638,N_3198);
and U3690 (N_3690,N_2417,N_3351);
and U3691 (N_3691,N_2986,N_3063);
or U3692 (N_3692,N_2788,N_2499);
or U3693 (N_3693,N_3387,N_2715);
and U3694 (N_3694,N_3015,N_3367);
nor U3695 (N_3695,N_2751,N_2416);
xor U3696 (N_3696,N_2741,N_3497);
xor U3697 (N_3697,N_3297,N_2415);
nand U3698 (N_3698,N_3210,N_3136);
nand U3699 (N_3699,N_3385,N_3056);
nor U3700 (N_3700,N_2743,N_3386);
nor U3701 (N_3701,N_2967,N_2406);
nand U3702 (N_3702,N_3107,N_3185);
or U3703 (N_3703,N_3520,N_3406);
and U3704 (N_3704,N_2575,N_2653);
nand U3705 (N_3705,N_3541,N_2845);
nor U3706 (N_3706,N_3338,N_2831);
xnor U3707 (N_3707,N_2548,N_3308);
xor U3708 (N_3708,N_3319,N_3593);
xor U3709 (N_3709,N_2525,N_2659);
xor U3710 (N_3710,N_3317,N_3383);
nand U3711 (N_3711,N_2768,N_2993);
xor U3712 (N_3712,N_2527,N_2975);
and U3713 (N_3713,N_2584,N_3200);
and U3714 (N_3714,N_3036,N_3058);
nand U3715 (N_3715,N_3434,N_3138);
xor U3716 (N_3716,N_3106,N_3237);
nand U3717 (N_3717,N_2428,N_2851);
nor U3718 (N_3718,N_2407,N_2461);
and U3719 (N_3719,N_2553,N_3576);
nand U3720 (N_3720,N_2826,N_2561);
nand U3721 (N_3721,N_2919,N_3331);
xnor U3722 (N_3722,N_3222,N_2410);
or U3723 (N_3723,N_2591,N_2853);
xor U3724 (N_3724,N_3217,N_3554);
nand U3725 (N_3725,N_3470,N_3265);
or U3726 (N_3726,N_2702,N_3044);
or U3727 (N_3727,N_2475,N_3365);
or U3728 (N_3728,N_2448,N_3524);
nand U3729 (N_3729,N_3445,N_3228);
nand U3730 (N_3730,N_2580,N_3586);
and U3731 (N_3731,N_3448,N_2621);
and U3732 (N_3732,N_3084,N_3489);
xor U3733 (N_3733,N_2489,N_3316);
or U3734 (N_3734,N_3537,N_3150);
or U3735 (N_3735,N_2503,N_3085);
nor U3736 (N_3736,N_2514,N_2711);
nand U3737 (N_3737,N_2625,N_3167);
or U3738 (N_3738,N_3504,N_2520);
nor U3739 (N_3739,N_3148,N_3569);
xnor U3740 (N_3740,N_3492,N_2902);
xor U3741 (N_3741,N_2445,N_3431);
xnor U3742 (N_3742,N_2913,N_2763);
nand U3743 (N_3743,N_3412,N_3246);
and U3744 (N_3744,N_2603,N_2983);
xor U3745 (N_3745,N_3472,N_2529);
nor U3746 (N_3746,N_3362,N_2516);
nand U3747 (N_3747,N_3395,N_2929);
or U3748 (N_3748,N_3221,N_3253);
nand U3749 (N_3749,N_3051,N_2923);
and U3750 (N_3750,N_2509,N_2742);
or U3751 (N_3751,N_3086,N_3267);
nor U3752 (N_3752,N_3156,N_2865);
nor U3753 (N_3753,N_2528,N_3396);
nand U3754 (N_3754,N_2816,N_3131);
nor U3755 (N_3755,N_2655,N_2854);
nor U3756 (N_3756,N_3354,N_2559);
xnor U3757 (N_3757,N_3499,N_3436);
and U3758 (N_3758,N_3323,N_3498);
xnor U3759 (N_3759,N_2914,N_2555);
xnor U3760 (N_3760,N_3288,N_3256);
or U3761 (N_3761,N_2629,N_2734);
nand U3762 (N_3762,N_3055,N_3241);
or U3763 (N_3763,N_3248,N_2656);
and U3764 (N_3764,N_3154,N_3556);
nor U3765 (N_3765,N_3273,N_2942);
xnor U3766 (N_3766,N_2643,N_3527);
or U3767 (N_3767,N_2492,N_2598);
nor U3768 (N_3768,N_3260,N_3513);
nand U3769 (N_3769,N_3230,N_3487);
nor U3770 (N_3770,N_3417,N_2678);
and U3771 (N_3771,N_2994,N_3227);
nand U3772 (N_3772,N_3269,N_3123);
and U3773 (N_3773,N_2602,N_2912);
or U3774 (N_3774,N_2688,N_2671);
nor U3775 (N_3775,N_2568,N_2524);
xor U3776 (N_3776,N_2841,N_2971);
nand U3777 (N_3777,N_2683,N_3213);
or U3778 (N_3778,N_2870,N_3119);
xor U3779 (N_3779,N_3511,N_2718);
and U3780 (N_3780,N_3207,N_2778);
xnor U3781 (N_3781,N_2782,N_3140);
or U3782 (N_3782,N_3070,N_2753);
or U3783 (N_3783,N_2999,N_3430);
nor U3784 (N_3784,N_3447,N_3202);
nand U3785 (N_3785,N_2820,N_3484);
or U3786 (N_3786,N_2478,N_2409);
xnor U3787 (N_3787,N_2574,N_2968);
nand U3788 (N_3788,N_2615,N_3264);
nand U3789 (N_3789,N_2490,N_3208);
xor U3790 (N_3790,N_3329,N_3559);
nor U3791 (N_3791,N_2585,N_3449);
xor U3792 (N_3792,N_3465,N_2985);
xnor U3793 (N_3793,N_2748,N_2807);
nor U3794 (N_3794,N_2484,N_3163);
and U3795 (N_3795,N_3364,N_2595);
and U3796 (N_3796,N_3312,N_2507);
and U3797 (N_3797,N_3049,N_2422);
and U3798 (N_3798,N_2660,N_2712);
nand U3799 (N_3799,N_3205,N_2632);
and U3800 (N_3800,N_2680,N_2819);
and U3801 (N_3801,N_2511,N_2570);
nand U3802 (N_3802,N_2984,N_3336);
or U3803 (N_3803,N_3439,N_3532);
nand U3804 (N_3804,N_3274,N_3182);
xor U3805 (N_3805,N_3224,N_2419);
and U3806 (N_3806,N_2486,N_2505);
nand U3807 (N_3807,N_3223,N_3054);
or U3808 (N_3808,N_2663,N_2988);
or U3809 (N_3809,N_2679,N_2843);
nor U3810 (N_3810,N_2508,N_3134);
or U3811 (N_3811,N_3374,N_3542);
xnor U3812 (N_3812,N_2978,N_2519);
nand U3813 (N_3813,N_3538,N_3309);
xnor U3814 (N_3814,N_2943,N_3120);
and U3815 (N_3815,N_3488,N_2446);
or U3816 (N_3816,N_3390,N_2631);
and U3817 (N_3817,N_2533,N_2411);
or U3818 (N_3818,N_3410,N_2973);
or U3819 (N_3819,N_3061,N_3127);
and U3820 (N_3820,N_2670,N_3068);
nor U3821 (N_3821,N_2771,N_2874);
nor U3822 (N_3822,N_3034,N_3306);
xor U3823 (N_3823,N_3584,N_3141);
nor U3824 (N_3824,N_2560,N_2847);
nand U3825 (N_3825,N_3192,N_2582);
or U3826 (N_3826,N_2927,N_3464);
and U3827 (N_3827,N_3149,N_2463);
nor U3828 (N_3828,N_3573,N_3519);
nand U3829 (N_3829,N_3583,N_3007);
nor U3830 (N_3830,N_2749,N_3515);
nand U3831 (N_3831,N_3144,N_3268);
nor U3832 (N_3832,N_3428,N_2767);
or U3833 (N_3833,N_2979,N_2714);
nand U3834 (N_3834,N_3400,N_3426);
xor U3835 (N_3835,N_3454,N_2777);
xor U3836 (N_3836,N_2932,N_3112);
and U3837 (N_3837,N_2639,N_2926);
or U3838 (N_3838,N_2803,N_3203);
and U3839 (N_3839,N_3392,N_3480);
nand U3840 (N_3840,N_3116,N_3043);
or U3841 (N_3841,N_2909,N_3234);
or U3842 (N_3842,N_2696,N_2905);
nor U3843 (N_3843,N_2472,N_3066);
xor U3844 (N_3844,N_3263,N_3195);
nor U3845 (N_3845,N_3009,N_2640);
and U3846 (N_3846,N_2961,N_3486);
nor U3847 (N_3847,N_2811,N_3408);
nand U3848 (N_3848,N_2989,N_3566);
nor U3849 (N_3849,N_2637,N_3057);
or U3850 (N_3850,N_3293,N_3516);
and U3851 (N_3851,N_3276,N_2813);
and U3852 (N_3852,N_3166,N_2617);
and U3853 (N_3853,N_2838,N_3025);
nand U3854 (N_3854,N_3012,N_2906);
xnor U3855 (N_3855,N_3372,N_2850);
xnor U3856 (N_3856,N_3359,N_2562);
nand U3857 (N_3857,N_2882,N_3553);
nor U3858 (N_3858,N_3528,N_3337);
xor U3859 (N_3859,N_2697,N_3425);
nand U3860 (N_3860,N_2589,N_3352);
nand U3861 (N_3861,N_2649,N_3184);
or U3862 (N_3862,N_3255,N_3468);
or U3863 (N_3863,N_2896,N_3340);
and U3864 (N_3864,N_3547,N_3496);
xor U3865 (N_3865,N_2464,N_2883);
or U3866 (N_3866,N_3523,N_3191);
nand U3867 (N_3867,N_3429,N_2835);
nor U3868 (N_3868,N_2668,N_2439);
xor U3869 (N_3869,N_3277,N_3121);
nor U3870 (N_3870,N_3076,N_2420);
or U3871 (N_3871,N_2452,N_2442);
nand U3872 (N_3872,N_3291,N_3204);
nor U3873 (N_3873,N_2996,N_3262);
and U3874 (N_3874,N_2936,N_2497);
or U3875 (N_3875,N_3310,N_2673);
and U3876 (N_3876,N_3162,N_2859);
or U3877 (N_3877,N_2583,N_3355);
or U3878 (N_3878,N_3422,N_3172);
or U3879 (N_3879,N_3567,N_3170);
nor U3880 (N_3880,N_3099,N_3245);
nor U3881 (N_3881,N_2834,N_2934);
or U3882 (N_3882,N_3419,N_2911);
or U3883 (N_3883,N_2844,N_3380);
nand U3884 (N_3884,N_2868,N_3502);
xnor U3885 (N_3885,N_2592,N_3442);
nor U3886 (N_3886,N_2667,N_3190);
or U3887 (N_3887,N_3008,N_2922);
xor U3888 (N_3888,N_3104,N_3577);
nand U3889 (N_3889,N_3373,N_3580);
xnor U3890 (N_3890,N_2737,N_2732);
and U3891 (N_3891,N_2567,N_3161);
nor U3892 (N_3892,N_3165,N_2674);
nor U3893 (N_3893,N_2885,N_2687);
nor U3894 (N_3894,N_3521,N_3437);
and U3895 (N_3895,N_3345,N_2980);
or U3896 (N_3896,N_3495,N_3023);
and U3897 (N_3897,N_3476,N_3549);
nand U3898 (N_3898,N_3282,N_3168);
and U3899 (N_3899,N_3173,N_3096);
xor U3900 (N_3900,N_2616,N_2487);
or U3901 (N_3901,N_2564,N_3074);
xnor U3902 (N_3902,N_2627,N_3053);
xnor U3903 (N_3903,N_2488,N_3244);
and U3904 (N_3904,N_3522,N_3111);
xnor U3905 (N_3905,N_2761,N_3401);
and U3906 (N_3906,N_3503,N_2910);
xnor U3907 (N_3907,N_3266,N_3302);
nor U3908 (N_3908,N_2708,N_3478);
or U3909 (N_3909,N_3414,N_3443);
nand U3910 (N_3910,N_2689,N_2758);
nand U3911 (N_3911,N_2920,N_2833);
and U3912 (N_3912,N_2775,N_3283);
xor U3913 (N_3913,N_3423,N_2646);
and U3914 (N_3914,N_3377,N_3562);
and U3915 (N_3915,N_3000,N_3506);
or U3916 (N_3916,N_3242,N_3589);
xnor U3917 (N_3917,N_2941,N_2776);
nand U3918 (N_3918,N_3531,N_3229);
nand U3919 (N_3919,N_3592,N_3591);
nor U3920 (N_3920,N_3176,N_2739);
xnor U3921 (N_3921,N_3514,N_2691);
xnor U3922 (N_3922,N_2766,N_2677);
or U3923 (N_3923,N_3193,N_2541);
or U3924 (N_3924,N_2916,N_3505);
xor U3925 (N_3925,N_2703,N_2873);
and U3926 (N_3926,N_3042,N_2745);
and U3927 (N_3927,N_2802,N_3579);
xor U3928 (N_3928,N_2815,N_3546);
nor U3929 (N_3929,N_3232,N_2495);
nor U3930 (N_3930,N_3100,N_2658);
nor U3931 (N_3931,N_3178,N_2787);
xor U3932 (N_3932,N_2402,N_2522);
nor U3933 (N_3933,N_3574,N_2950);
or U3934 (N_3934,N_3530,N_3098);
xor U3935 (N_3935,N_2469,N_3278);
and U3936 (N_3936,N_3328,N_3284);
and U3937 (N_3937,N_3048,N_3544);
or U3938 (N_3938,N_3469,N_2494);
nand U3939 (N_3939,N_3067,N_2804);
and U3940 (N_3940,N_2611,N_3102);
nand U3941 (N_3941,N_2538,N_2863);
xnor U3942 (N_3942,N_2423,N_3597);
or U3943 (N_3943,N_2752,N_2662);
nor U3944 (N_3944,N_2963,N_3363);
and U3945 (N_3945,N_2675,N_2684);
and U3946 (N_3946,N_2907,N_3017);
nor U3947 (N_3947,N_2889,N_3295);
and U3948 (N_3948,N_2812,N_3560);
xnor U3949 (N_3949,N_2785,N_2644);
and U3950 (N_3950,N_2552,N_2500);
xor U3951 (N_3951,N_3050,N_3536);
and U3952 (N_3952,N_2783,N_2931);
and U3953 (N_3953,N_3021,N_3002);
nor U3954 (N_3954,N_2827,N_3071);
or U3955 (N_3955,N_2483,N_3087);
nand U3956 (N_3956,N_2665,N_3424);
or U3957 (N_3957,N_3461,N_3535);
or U3958 (N_3958,N_2669,N_3314);
nand U3959 (N_3959,N_2817,N_2609);
xnor U3960 (N_3960,N_3339,N_3341);
nor U3961 (N_3961,N_2948,N_3272);
nor U3962 (N_3962,N_2736,N_2651);
and U3963 (N_3963,N_3077,N_2551);
nand U3964 (N_3964,N_2619,N_2457);
nor U3965 (N_3965,N_3458,N_2730);
or U3966 (N_3966,N_2731,N_3389);
xnor U3967 (N_3967,N_2501,N_3349);
or U3968 (N_3968,N_3575,N_3147);
nand U3969 (N_3969,N_2654,N_2545);
and U3970 (N_3970,N_2779,N_3233);
nand U3971 (N_3971,N_2861,N_2805);
and U3972 (N_3972,N_2740,N_3108);
xnor U3973 (N_3973,N_3360,N_2641);
nor U3974 (N_3974,N_3247,N_2425);
and U3975 (N_3975,N_2789,N_3196);
xor U3976 (N_3976,N_2717,N_2477);
nor U3977 (N_3977,N_2762,N_2842);
nor U3978 (N_3978,N_2900,N_2502);
xnor U3979 (N_3979,N_2685,N_2642);
xnor U3980 (N_3980,N_2496,N_2858);
nor U3981 (N_3981,N_2781,N_3081);
nand U3982 (N_3982,N_2476,N_2769);
nand U3983 (N_3983,N_3332,N_2454);
and U3984 (N_3984,N_2546,N_3459);
xor U3985 (N_3985,N_2435,N_2535);
or U3986 (N_3986,N_3518,N_3254);
and U3987 (N_3987,N_3304,N_2468);
or U3988 (N_3988,N_2809,N_2918);
nand U3989 (N_3989,N_2459,N_2626);
and U3990 (N_3990,N_3045,N_2523);
nor U3991 (N_3991,N_2765,N_3418);
and U3992 (N_3992,N_2808,N_3427);
and U3993 (N_3993,N_2701,N_2650);
xnor U3994 (N_3994,N_2605,N_3333);
nand U3995 (N_3995,N_3080,N_3482);
or U3996 (N_3996,N_2513,N_2600);
nand U3997 (N_3997,N_3001,N_2596);
xnor U3998 (N_3998,N_2810,N_3142);
nand U3999 (N_3999,N_2757,N_2634);
xor U4000 (N_4000,N_3296,N_3420);
and U4001 (N_4001,N_2924,N_3183);
nor U4002 (N_4002,N_3483,N_2657);
nor U4003 (N_4003,N_2964,N_2935);
xor U4004 (N_4004,N_3271,N_3500);
and U4005 (N_4005,N_2756,N_2536);
or U4006 (N_4006,N_3212,N_2672);
nor U4007 (N_4007,N_3181,N_3578);
nand U4008 (N_4008,N_2818,N_3507);
xor U4009 (N_4009,N_3381,N_3020);
xnor U4010 (N_4010,N_3151,N_2728);
nor U4011 (N_4011,N_2581,N_2908);
or U4012 (N_4012,N_3027,N_2998);
nor U4013 (N_4013,N_3075,N_2729);
nor U4014 (N_4014,N_2465,N_3124);
and U4015 (N_4015,N_3197,N_2543);
xor U4016 (N_4016,N_3327,N_3416);
xnor U4017 (N_4017,N_2622,N_2414);
nor U4018 (N_4018,N_2852,N_3152);
and U4019 (N_4019,N_2517,N_2594);
and U4020 (N_4020,N_3290,N_3433);
nor U4021 (N_4021,N_2821,N_2563);
and U4022 (N_4022,N_3175,N_2597);
and U4023 (N_4023,N_3031,N_3095);
nand U4024 (N_4024,N_2959,N_2997);
nand U4025 (N_4025,N_2430,N_2974);
and U4026 (N_4026,N_3326,N_3252);
or U4027 (N_4027,N_3093,N_2720);
nand U4028 (N_4028,N_3270,N_3079);
and U4029 (N_4029,N_2706,N_3169);
nand U4030 (N_4030,N_3101,N_2991);
nand U4031 (N_4031,N_3361,N_3019);
nand U4032 (N_4032,N_2413,N_3409);
and U4033 (N_4033,N_3343,N_2937);
or U4034 (N_4034,N_3324,N_3462);
or U4035 (N_4035,N_2772,N_3249);
nor U4036 (N_4036,N_2443,N_3062);
or U4037 (N_4037,N_3280,N_3187);
and U4038 (N_4038,N_3402,N_2613);
and U4039 (N_4039,N_2530,N_2569);
and U4040 (N_4040,N_2759,N_2512);
and U4041 (N_4041,N_2648,N_2946);
nor U4042 (N_4042,N_3158,N_2630);
nand U4043 (N_4043,N_2957,N_3555);
xor U4044 (N_4044,N_2981,N_2645);
or U4045 (N_4045,N_3029,N_2429);
and U4046 (N_4046,N_2888,N_2939);
and U4047 (N_4047,N_3357,N_3334);
nor U4048 (N_4048,N_3125,N_3315);
nand U4049 (N_4049,N_3375,N_2770);
xnor U4050 (N_4050,N_2549,N_2408);
or U4051 (N_4051,N_3411,N_2624);
nor U4052 (N_4052,N_3041,N_3238);
xnor U4053 (N_4053,N_2857,N_2709);
and U4054 (N_4054,N_3378,N_3194);
and U4055 (N_4055,N_3494,N_3368);
nand U4056 (N_4056,N_2693,N_3466);
xnor U4057 (N_4057,N_2652,N_2573);
or U4058 (N_4058,N_2578,N_2604);
or U4059 (N_4059,N_3186,N_3179);
and U4060 (N_4060,N_2723,N_2666);
xor U4061 (N_4061,N_3525,N_2586);
and U4062 (N_4062,N_2557,N_2449);
or U4063 (N_4063,N_3572,N_3281);
nor U4064 (N_4064,N_2426,N_3350);
or U4065 (N_4065,N_2746,N_3113);
or U4066 (N_4066,N_2990,N_2661);
and U4067 (N_4067,N_3477,N_2894);
xor U4068 (N_4068,N_2504,N_2456);
and U4069 (N_4069,N_2839,N_3218);
or U4070 (N_4070,N_3118,N_2506);
nand U4071 (N_4071,N_3115,N_2436);
or U4072 (N_4072,N_3508,N_2904);
xor U4073 (N_4073,N_2725,N_2462);
nor U4074 (N_4074,N_2969,N_2887);
nor U4075 (N_4075,N_3240,N_2515);
xor U4076 (N_4076,N_2510,N_3540);
nor U4077 (N_4077,N_3129,N_3083);
and U4078 (N_4078,N_3545,N_2790);
nand U4079 (N_4079,N_2944,N_2695);
nand U4080 (N_4080,N_3371,N_2860);
and U4081 (N_4081,N_3481,N_2940);
and U4082 (N_4082,N_3509,N_2800);
nand U4083 (N_4083,N_3206,N_3174);
nand U4084 (N_4084,N_3047,N_2432);
or U4085 (N_4085,N_3456,N_2796);
nand U4086 (N_4086,N_3126,N_2791);
or U4087 (N_4087,N_2698,N_3132);
xnor U4088 (N_4088,N_3300,N_3463);
and U4089 (N_4089,N_3014,N_2722);
nor U4090 (N_4090,N_2837,N_2521);
nand U4091 (N_4091,N_3344,N_2572);
or U4092 (N_4092,N_2577,N_2877);
nor U4093 (N_4093,N_3485,N_2493);
nor U4094 (N_4094,N_2938,N_3005);
or U4095 (N_4095,N_2534,N_2618);
nand U4096 (N_4096,N_2750,N_3286);
and U4097 (N_4097,N_2825,N_2719);
xnor U4098 (N_4098,N_3533,N_2897);
or U4099 (N_4099,N_3446,N_2544);
nand U4100 (N_4100,N_2855,N_2405);
xor U4101 (N_4101,N_3391,N_3040);
and U4102 (N_4102,N_3539,N_2965);
nand U4103 (N_4103,N_2547,N_2862);
or U4104 (N_4104,N_2875,N_3453);
nor U4105 (N_4105,N_3035,N_3455);
nand U4106 (N_4106,N_2482,N_3292);
or U4107 (N_4107,N_3117,N_3534);
nor U4108 (N_4108,N_3153,N_2792);
xor U4109 (N_4109,N_2438,N_3298);
nor U4110 (N_4110,N_3114,N_2647);
nor U4111 (N_4111,N_2424,N_3214);
xor U4112 (N_4112,N_3479,N_2822);
nand U4113 (N_4113,N_2982,N_2427);
xnor U4114 (N_4114,N_2480,N_3452);
or U4115 (N_4115,N_3250,N_2992);
nand U4116 (N_4116,N_3215,N_2566);
or U4117 (N_4117,N_3346,N_2576);
xor U4118 (N_4118,N_2891,N_2537);
nor U4119 (N_4119,N_2532,N_2814);
or U4120 (N_4120,N_3413,N_3398);
and U4121 (N_4121,N_3180,N_2744);
nor U4122 (N_4122,N_3133,N_2892);
and U4123 (N_4123,N_2928,N_3570);
nor U4124 (N_4124,N_3128,N_2755);
nand U4125 (N_4125,N_3003,N_3143);
nand U4126 (N_4126,N_2869,N_2526);
or U4127 (N_4127,N_3039,N_2866);
and U4128 (N_4128,N_2949,N_3105);
nand U4129 (N_4129,N_3094,N_2466);
or U4130 (N_4130,N_2707,N_2518);
or U4131 (N_4131,N_3037,N_2794);
and U4132 (N_4132,N_3564,N_3594);
xor U4133 (N_4133,N_2633,N_3582);
xor U4134 (N_4134,N_2774,N_2444);
nand U4135 (N_4135,N_3236,N_3397);
nor U4136 (N_4136,N_3356,N_3490);
or U4137 (N_4137,N_2620,N_2608);
and U4138 (N_4138,N_2823,N_2915);
nand U4139 (N_4139,N_2599,N_2890);
nor U4140 (N_4140,N_3259,N_2453);
or U4141 (N_4141,N_3366,N_3082);
nand U4142 (N_4142,N_2754,N_3384);
or U4143 (N_4143,N_2798,N_3251);
or U4144 (N_4144,N_3157,N_3299);
nand U4145 (N_4145,N_3561,N_2470);
nand U4146 (N_4146,N_3097,N_2404);
and U4147 (N_4147,N_3568,N_2840);
nand U4148 (N_4148,N_3209,N_2458);
nor U4149 (N_4149,N_3403,N_3033);
xnor U4150 (N_4150,N_3018,N_3460);
and U4151 (N_4151,N_2460,N_3130);
nand U4152 (N_4152,N_3585,N_2716);
nor U4153 (N_4153,N_3103,N_2694);
or U4154 (N_4154,N_2542,N_3145);
nand U4155 (N_4155,N_3370,N_2588);
or U4156 (N_4156,N_3588,N_2786);
xor U4157 (N_4157,N_2471,N_2899);
nand U4158 (N_4158,N_2692,N_2614);
xnor U4159 (N_4159,N_3558,N_3599);
and U4160 (N_4160,N_3320,N_2945);
nor U4161 (N_4161,N_2713,N_2601);
nor U4162 (N_4162,N_3595,N_3307);
xor U4163 (N_4163,N_3440,N_2947);
or U4164 (N_4164,N_3059,N_2747);
xor U4165 (N_4165,N_2773,N_3110);
nand U4166 (N_4166,N_3335,N_2623);
or U4167 (N_4167,N_3467,N_3188);
or U4168 (N_4168,N_2479,N_3388);
and U4169 (N_4169,N_3587,N_2933);
and U4170 (N_4170,N_2884,N_3330);
nor U4171 (N_4171,N_2590,N_2593);
xor U4172 (N_4172,N_3457,N_2828);
xnor U4173 (N_4173,N_2531,N_3289);
xor U4174 (N_4174,N_3301,N_2721);
xnor U4175 (N_4175,N_2903,N_2498);
nand U4176 (N_4176,N_2925,N_3432);
and U4177 (N_4177,N_2886,N_3160);
or U4178 (N_4178,N_3379,N_2700);
xor U4179 (N_4179,N_3226,N_3348);
nand U4180 (N_4180,N_2441,N_2710);
nand U4181 (N_4181,N_3473,N_2876);
xnor U4182 (N_4182,N_2871,N_2727);
xnor U4183 (N_4183,N_3090,N_3451);
or U4184 (N_4184,N_3189,N_2995);
and U4185 (N_4185,N_3199,N_2628);
xor U4186 (N_4186,N_2401,N_2467);
or U4187 (N_4187,N_3052,N_2784);
xnor U4188 (N_4188,N_3004,N_2951);
xor U4189 (N_4189,N_2824,N_3235);
and U4190 (N_4190,N_3548,N_3146);
xor U4191 (N_4191,N_2917,N_3303);
and U4192 (N_4192,N_2485,N_3028);
xor U4193 (N_4193,N_2848,N_2699);
nand U4194 (N_4194,N_2437,N_3512);
and U4195 (N_4195,N_2473,N_2881);
nor U4196 (N_4196,N_3159,N_3155);
xor U4197 (N_4197,N_2830,N_3557);
nor U4198 (N_4198,N_3305,N_3257);
xor U4199 (N_4199,N_3073,N_3030);
nor U4200 (N_4200,N_3538,N_3317);
and U4201 (N_4201,N_3047,N_3378);
or U4202 (N_4202,N_2938,N_2927);
xor U4203 (N_4203,N_3069,N_3025);
nand U4204 (N_4204,N_2565,N_2639);
and U4205 (N_4205,N_3124,N_2823);
nand U4206 (N_4206,N_2877,N_2690);
xnor U4207 (N_4207,N_3490,N_3257);
xnor U4208 (N_4208,N_2760,N_2590);
xor U4209 (N_4209,N_2848,N_2559);
nand U4210 (N_4210,N_3282,N_3323);
or U4211 (N_4211,N_3447,N_2679);
and U4212 (N_4212,N_2628,N_3076);
or U4213 (N_4213,N_2507,N_3479);
xor U4214 (N_4214,N_3425,N_2779);
nand U4215 (N_4215,N_3582,N_3506);
nor U4216 (N_4216,N_2557,N_2636);
xnor U4217 (N_4217,N_3374,N_3388);
and U4218 (N_4218,N_3281,N_3210);
and U4219 (N_4219,N_2915,N_2725);
or U4220 (N_4220,N_2417,N_3557);
xor U4221 (N_4221,N_3286,N_3588);
and U4222 (N_4222,N_2884,N_3414);
or U4223 (N_4223,N_3036,N_3455);
xnor U4224 (N_4224,N_3590,N_2913);
nor U4225 (N_4225,N_3562,N_2801);
and U4226 (N_4226,N_2999,N_3521);
xor U4227 (N_4227,N_3145,N_2787);
nor U4228 (N_4228,N_3379,N_3141);
nand U4229 (N_4229,N_3206,N_2988);
or U4230 (N_4230,N_2520,N_2628);
nand U4231 (N_4231,N_3053,N_2521);
or U4232 (N_4232,N_2711,N_3102);
or U4233 (N_4233,N_3124,N_2793);
nor U4234 (N_4234,N_2874,N_2542);
nor U4235 (N_4235,N_2829,N_3064);
xnor U4236 (N_4236,N_2412,N_2934);
nand U4237 (N_4237,N_3357,N_2451);
xnor U4238 (N_4238,N_2518,N_2560);
xor U4239 (N_4239,N_3355,N_3287);
nor U4240 (N_4240,N_3408,N_2799);
nor U4241 (N_4241,N_2796,N_2461);
and U4242 (N_4242,N_3492,N_3166);
and U4243 (N_4243,N_2556,N_2496);
or U4244 (N_4244,N_3540,N_3370);
and U4245 (N_4245,N_3440,N_3568);
or U4246 (N_4246,N_3219,N_3217);
nor U4247 (N_4247,N_2751,N_2537);
nand U4248 (N_4248,N_2796,N_2691);
nand U4249 (N_4249,N_2981,N_2475);
xor U4250 (N_4250,N_2432,N_2562);
xnor U4251 (N_4251,N_2805,N_3058);
nor U4252 (N_4252,N_2681,N_2530);
or U4253 (N_4253,N_2742,N_2655);
nor U4254 (N_4254,N_3336,N_2804);
nor U4255 (N_4255,N_3155,N_2731);
or U4256 (N_4256,N_3334,N_3038);
or U4257 (N_4257,N_3009,N_2615);
and U4258 (N_4258,N_2908,N_2703);
and U4259 (N_4259,N_3053,N_2578);
nand U4260 (N_4260,N_2479,N_2500);
and U4261 (N_4261,N_3391,N_3464);
or U4262 (N_4262,N_3356,N_2643);
or U4263 (N_4263,N_3469,N_2439);
nand U4264 (N_4264,N_2922,N_2782);
nand U4265 (N_4265,N_2733,N_2511);
and U4266 (N_4266,N_2965,N_2610);
or U4267 (N_4267,N_3359,N_2598);
nor U4268 (N_4268,N_2602,N_3551);
xor U4269 (N_4269,N_3140,N_2779);
and U4270 (N_4270,N_3233,N_3324);
or U4271 (N_4271,N_3008,N_3388);
xnor U4272 (N_4272,N_2722,N_2604);
xnor U4273 (N_4273,N_3278,N_3216);
or U4274 (N_4274,N_3122,N_2654);
xnor U4275 (N_4275,N_3287,N_2736);
or U4276 (N_4276,N_3377,N_3077);
and U4277 (N_4277,N_2616,N_3226);
nor U4278 (N_4278,N_2792,N_2502);
xor U4279 (N_4279,N_2954,N_3285);
nand U4280 (N_4280,N_2438,N_3294);
and U4281 (N_4281,N_2492,N_3085);
and U4282 (N_4282,N_3453,N_3171);
and U4283 (N_4283,N_2653,N_2998);
nand U4284 (N_4284,N_3283,N_2472);
nand U4285 (N_4285,N_3257,N_2601);
or U4286 (N_4286,N_3426,N_2887);
nor U4287 (N_4287,N_3137,N_3371);
or U4288 (N_4288,N_2985,N_3186);
or U4289 (N_4289,N_3237,N_2418);
nor U4290 (N_4290,N_3286,N_2581);
nor U4291 (N_4291,N_2986,N_2968);
xor U4292 (N_4292,N_3572,N_2605);
nor U4293 (N_4293,N_2684,N_2530);
xnor U4294 (N_4294,N_3402,N_3049);
or U4295 (N_4295,N_2628,N_2792);
and U4296 (N_4296,N_2566,N_2461);
or U4297 (N_4297,N_2700,N_3238);
or U4298 (N_4298,N_2934,N_3403);
and U4299 (N_4299,N_3551,N_2738);
xor U4300 (N_4300,N_2647,N_3576);
xor U4301 (N_4301,N_2555,N_2610);
or U4302 (N_4302,N_3568,N_2946);
xor U4303 (N_4303,N_2475,N_2577);
and U4304 (N_4304,N_3437,N_2424);
and U4305 (N_4305,N_3015,N_3121);
xnor U4306 (N_4306,N_2562,N_3147);
and U4307 (N_4307,N_3355,N_2419);
nand U4308 (N_4308,N_2523,N_2961);
nor U4309 (N_4309,N_2474,N_2946);
or U4310 (N_4310,N_2613,N_2909);
nand U4311 (N_4311,N_3449,N_2576);
and U4312 (N_4312,N_2642,N_2960);
nor U4313 (N_4313,N_2670,N_2763);
nand U4314 (N_4314,N_2809,N_2671);
xnor U4315 (N_4315,N_2928,N_2813);
xor U4316 (N_4316,N_2676,N_2576);
or U4317 (N_4317,N_3533,N_2664);
nor U4318 (N_4318,N_3095,N_3355);
or U4319 (N_4319,N_3473,N_2911);
xnor U4320 (N_4320,N_3048,N_2740);
xor U4321 (N_4321,N_3510,N_2939);
xor U4322 (N_4322,N_2673,N_3193);
nor U4323 (N_4323,N_2401,N_2893);
and U4324 (N_4324,N_3497,N_2556);
nand U4325 (N_4325,N_2443,N_2697);
or U4326 (N_4326,N_3346,N_3457);
nand U4327 (N_4327,N_3224,N_3397);
xnor U4328 (N_4328,N_2830,N_3359);
or U4329 (N_4329,N_2846,N_3196);
xor U4330 (N_4330,N_3399,N_2833);
or U4331 (N_4331,N_2766,N_2512);
xnor U4332 (N_4332,N_2654,N_3434);
and U4333 (N_4333,N_2951,N_2643);
nor U4334 (N_4334,N_2499,N_3288);
xor U4335 (N_4335,N_3051,N_3101);
and U4336 (N_4336,N_2411,N_3360);
nor U4337 (N_4337,N_2782,N_2584);
or U4338 (N_4338,N_2631,N_2480);
or U4339 (N_4339,N_2469,N_3437);
or U4340 (N_4340,N_2665,N_3092);
nor U4341 (N_4341,N_3589,N_3530);
or U4342 (N_4342,N_2498,N_3178);
or U4343 (N_4343,N_2433,N_3532);
nand U4344 (N_4344,N_2949,N_2700);
nand U4345 (N_4345,N_2882,N_3239);
nand U4346 (N_4346,N_2898,N_3383);
xor U4347 (N_4347,N_3030,N_2901);
xnor U4348 (N_4348,N_3073,N_3279);
or U4349 (N_4349,N_3030,N_2915);
xnor U4350 (N_4350,N_2870,N_2761);
or U4351 (N_4351,N_3252,N_2778);
nand U4352 (N_4352,N_2465,N_2767);
nor U4353 (N_4353,N_3543,N_2407);
nand U4354 (N_4354,N_3156,N_3128);
or U4355 (N_4355,N_3106,N_2839);
nand U4356 (N_4356,N_2838,N_2534);
nor U4357 (N_4357,N_2978,N_2403);
or U4358 (N_4358,N_3048,N_2659);
and U4359 (N_4359,N_3183,N_2533);
nor U4360 (N_4360,N_2822,N_3093);
or U4361 (N_4361,N_3556,N_3514);
or U4362 (N_4362,N_2960,N_2701);
or U4363 (N_4363,N_2577,N_3201);
or U4364 (N_4364,N_2553,N_2950);
and U4365 (N_4365,N_2730,N_2521);
and U4366 (N_4366,N_2651,N_2635);
nand U4367 (N_4367,N_2553,N_2752);
and U4368 (N_4368,N_2887,N_2654);
xnor U4369 (N_4369,N_2565,N_2486);
nor U4370 (N_4370,N_3158,N_3370);
or U4371 (N_4371,N_3181,N_3532);
nand U4372 (N_4372,N_2848,N_3586);
and U4373 (N_4373,N_2951,N_3241);
and U4374 (N_4374,N_2597,N_3441);
nand U4375 (N_4375,N_3200,N_3507);
nor U4376 (N_4376,N_3574,N_2629);
nor U4377 (N_4377,N_3128,N_2573);
or U4378 (N_4378,N_2929,N_3580);
nor U4379 (N_4379,N_2442,N_2932);
or U4380 (N_4380,N_3455,N_2625);
xor U4381 (N_4381,N_2946,N_2737);
nand U4382 (N_4382,N_2601,N_2677);
nor U4383 (N_4383,N_2881,N_2860);
and U4384 (N_4384,N_2442,N_3424);
xor U4385 (N_4385,N_3329,N_2643);
nand U4386 (N_4386,N_2540,N_2517);
xor U4387 (N_4387,N_2459,N_2516);
and U4388 (N_4388,N_2679,N_3107);
nor U4389 (N_4389,N_3553,N_2517);
xor U4390 (N_4390,N_3595,N_3403);
nand U4391 (N_4391,N_3439,N_3487);
or U4392 (N_4392,N_3295,N_2645);
nand U4393 (N_4393,N_2426,N_3578);
nand U4394 (N_4394,N_3249,N_3419);
nor U4395 (N_4395,N_2565,N_3092);
nor U4396 (N_4396,N_2955,N_3445);
nand U4397 (N_4397,N_3577,N_3528);
xor U4398 (N_4398,N_2414,N_2406);
nand U4399 (N_4399,N_3590,N_2851);
xor U4400 (N_4400,N_2871,N_2901);
or U4401 (N_4401,N_3229,N_2908);
xnor U4402 (N_4402,N_3413,N_3084);
nand U4403 (N_4403,N_3171,N_3457);
nand U4404 (N_4404,N_3425,N_3125);
nand U4405 (N_4405,N_3308,N_3536);
nor U4406 (N_4406,N_2520,N_3211);
nor U4407 (N_4407,N_2667,N_3083);
xnor U4408 (N_4408,N_3097,N_3181);
nand U4409 (N_4409,N_3315,N_2404);
nand U4410 (N_4410,N_3425,N_2850);
nor U4411 (N_4411,N_3004,N_3241);
or U4412 (N_4412,N_2586,N_2543);
nor U4413 (N_4413,N_2452,N_2550);
or U4414 (N_4414,N_2782,N_3076);
or U4415 (N_4415,N_2667,N_2762);
xor U4416 (N_4416,N_3456,N_3026);
or U4417 (N_4417,N_2690,N_2530);
or U4418 (N_4418,N_3311,N_2642);
nor U4419 (N_4419,N_2507,N_3574);
nor U4420 (N_4420,N_3348,N_3524);
or U4421 (N_4421,N_2557,N_3490);
nor U4422 (N_4422,N_3556,N_3270);
or U4423 (N_4423,N_2848,N_2931);
nor U4424 (N_4424,N_2735,N_3354);
or U4425 (N_4425,N_2799,N_3488);
nor U4426 (N_4426,N_3081,N_2761);
xnor U4427 (N_4427,N_3315,N_2481);
or U4428 (N_4428,N_3293,N_2798);
and U4429 (N_4429,N_3358,N_2485);
and U4430 (N_4430,N_2925,N_2910);
and U4431 (N_4431,N_2433,N_2911);
nand U4432 (N_4432,N_2574,N_3364);
and U4433 (N_4433,N_3479,N_3195);
xor U4434 (N_4434,N_3021,N_2587);
nand U4435 (N_4435,N_2956,N_3434);
and U4436 (N_4436,N_3102,N_2605);
and U4437 (N_4437,N_2859,N_2955);
and U4438 (N_4438,N_2506,N_2563);
nor U4439 (N_4439,N_3589,N_2956);
and U4440 (N_4440,N_3389,N_2699);
or U4441 (N_4441,N_3104,N_3238);
nand U4442 (N_4442,N_2984,N_2597);
or U4443 (N_4443,N_2661,N_2791);
nand U4444 (N_4444,N_2832,N_3284);
nand U4445 (N_4445,N_3553,N_2693);
nand U4446 (N_4446,N_3432,N_2527);
xor U4447 (N_4447,N_2652,N_2530);
or U4448 (N_4448,N_2933,N_2503);
or U4449 (N_4449,N_2623,N_2540);
nor U4450 (N_4450,N_3397,N_3057);
nor U4451 (N_4451,N_2625,N_2513);
and U4452 (N_4452,N_2597,N_3316);
xor U4453 (N_4453,N_2960,N_3569);
and U4454 (N_4454,N_2716,N_2766);
nor U4455 (N_4455,N_3535,N_3030);
nand U4456 (N_4456,N_3191,N_2571);
xnor U4457 (N_4457,N_3053,N_2785);
and U4458 (N_4458,N_3412,N_2859);
nor U4459 (N_4459,N_2903,N_2856);
nand U4460 (N_4460,N_3521,N_3097);
nor U4461 (N_4461,N_3130,N_2606);
nand U4462 (N_4462,N_3342,N_3466);
nor U4463 (N_4463,N_2949,N_2419);
xor U4464 (N_4464,N_2716,N_2710);
xor U4465 (N_4465,N_2849,N_2593);
or U4466 (N_4466,N_2517,N_3210);
and U4467 (N_4467,N_2976,N_2663);
or U4468 (N_4468,N_3400,N_3051);
xnor U4469 (N_4469,N_2895,N_3160);
nand U4470 (N_4470,N_3349,N_2693);
xnor U4471 (N_4471,N_2420,N_3465);
nand U4472 (N_4472,N_3226,N_3527);
or U4473 (N_4473,N_2580,N_2941);
xor U4474 (N_4474,N_3439,N_3078);
nor U4475 (N_4475,N_2578,N_3271);
nand U4476 (N_4476,N_2609,N_2645);
nand U4477 (N_4477,N_3202,N_2868);
and U4478 (N_4478,N_3346,N_2444);
nor U4479 (N_4479,N_2818,N_3444);
or U4480 (N_4480,N_2574,N_3392);
nor U4481 (N_4481,N_2492,N_3402);
xnor U4482 (N_4482,N_2449,N_3332);
nor U4483 (N_4483,N_2754,N_3494);
and U4484 (N_4484,N_2890,N_3385);
or U4485 (N_4485,N_3198,N_3022);
or U4486 (N_4486,N_2446,N_3517);
and U4487 (N_4487,N_3026,N_3059);
or U4488 (N_4488,N_3148,N_3505);
nand U4489 (N_4489,N_3375,N_3367);
nor U4490 (N_4490,N_3041,N_3223);
or U4491 (N_4491,N_3428,N_2792);
nor U4492 (N_4492,N_3457,N_2869);
nor U4493 (N_4493,N_2970,N_3259);
nor U4494 (N_4494,N_3400,N_2509);
nor U4495 (N_4495,N_3090,N_3194);
nor U4496 (N_4496,N_2432,N_2553);
and U4497 (N_4497,N_2855,N_2778);
nor U4498 (N_4498,N_2409,N_2879);
nand U4499 (N_4499,N_2659,N_3030);
or U4500 (N_4500,N_2753,N_2948);
xnor U4501 (N_4501,N_3447,N_3394);
xnor U4502 (N_4502,N_3495,N_3425);
and U4503 (N_4503,N_3486,N_3513);
and U4504 (N_4504,N_3113,N_3052);
or U4505 (N_4505,N_2836,N_3032);
nand U4506 (N_4506,N_2576,N_2642);
nand U4507 (N_4507,N_3534,N_2993);
nand U4508 (N_4508,N_2895,N_3415);
and U4509 (N_4509,N_2621,N_2912);
nand U4510 (N_4510,N_2908,N_2440);
nand U4511 (N_4511,N_2460,N_3193);
nand U4512 (N_4512,N_3213,N_2556);
nor U4513 (N_4513,N_3563,N_2668);
nand U4514 (N_4514,N_3590,N_3562);
and U4515 (N_4515,N_3567,N_3516);
or U4516 (N_4516,N_2617,N_3348);
nand U4517 (N_4517,N_3359,N_2893);
or U4518 (N_4518,N_3132,N_2659);
nand U4519 (N_4519,N_3371,N_2815);
and U4520 (N_4520,N_3129,N_3274);
nand U4521 (N_4521,N_3098,N_3542);
nor U4522 (N_4522,N_3555,N_2824);
nand U4523 (N_4523,N_2479,N_3040);
nor U4524 (N_4524,N_3599,N_3491);
xor U4525 (N_4525,N_2878,N_3341);
nor U4526 (N_4526,N_3486,N_2817);
nand U4527 (N_4527,N_3337,N_2990);
nor U4528 (N_4528,N_3015,N_2646);
nand U4529 (N_4529,N_3040,N_2422);
nor U4530 (N_4530,N_2656,N_3512);
xor U4531 (N_4531,N_3586,N_3390);
nand U4532 (N_4532,N_2879,N_3265);
xor U4533 (N_4533,N_3011,N_2659);
nor U4534 (N_4534,N_2764,N_3467);
or U4535 (N_4535,N_2861,N_3407);
and U4536 (N_4536,N_2704,N_2418);
and U4537 (N_4537,N_3091,N_2573);
nor U4538 (N_4538,N_2523,N_3006);
xor U4539 (N_4539,N_3172,N_2730);
nand U4540 (N_4540,N_3323,N_2765);
nand U4541 (N_4541,N_2917,N_2490);
nand U4542 (N_4542,N_2595,N_3249);
or U4543 (N_4543,N_3340,N_3555);
xor U4544 (N_4544,N_2481,N_3114);
and U4545 (N_4545,N_3034,N_2865);
and U4546 (N_4546,N_3178,N_3095);
nand U4547 (N_4547,N_2594,N_2706);
nand U4548 (N_4548,N_2698,N_3331);
nand U4549 (N_4549,N_2874,N_3024);
nor U4550 (N_4550,N_3230,N_2756);
nand U4551 (N_4551,N_3451,N_2521);
or U4552 (N_4552,N_2695,N_2939);
nor U4553 (N_4553,N_2908,N_2849);
or U4554 (N_4554,N_3126,N_2953);
nor U4555 (N_4555,N_2869,N_2639);
and U4556 (N_4556,N_3066,N_2903);
and U4557 (N_4557,N_3231,N_2579);
or U4558 (N_4558,N_2525,N_2637);
nand U4559 (N_4559,N_2932,N_3473);
nor U4560 (N_4560,N_3086,N_2678);
xnor U4561 (N_4561,N_2508,N_2487);
nand U4562 (N_4562,N_3171,N_3537);
xnor U4563 (N_4563,N_2954,N_2932);
xnor U4564 (N_4564,N_3235,N_3529);
xor U4565 (N_4565,N_2506,N_2457);
or U4566 (N_4566,N_2572,N_2789);
nand U4567 (N_4567,N_2557,N_3078);
or U4568 (N_4568,N_3232,N_2738);
nor U4569 (N_4569,N_3127,N_2402);
nand U4570 (N_4570,N_3440,N_2452);
or U4571 (N_4571,N_3555,N_2664);
nand U4572 (N_4572,N_3545,N_3230);
and U4573 (N_4573,N_3334,N_2506);
nand U4574 (N_4574,N_3269,N_3178);
nand U4575 (N_4575,N_2446,N_2665);
or U4576 (N_4576,N_2490,N_3458);
and U4577 (N_4577,N_2899,N_3173);
and U4578 (N_4578,N_3571,N_2556);
and U4579 (N_4579,N_2458,N_3444);
or U4580 (N_4580,N_3597,N_3434);
and U4581 (N_4581,N_2955,N_3161);
nor U4582 (N_4582,N_3514,N_2748);
and U4583 (N_4583,N_2898,N_3070);
nand U4584 (N_4584,N_3592,N_3170);
xor U4585 (N_4585,N_2590,N_2569);
nand U4586 (N_4586,N_2584,N_3306);
xnor U4587 (N_4587,N_2581,N_2859);
nand U4588 (N_4588,N_3443,N_2454);
and U4589 (N_4589,N_3138,N_3062);
nand U4590 (N_4590,N_2813,N_2982);
and U4591 (N_4591,N_3549,N_2644);
xnor U4592 (N_4592,N_2468,N_2805);
and U4593 (N_4593,N_2527,N_3470);
nand U4594 (N_4594,N_2534,N_3187);
and U4595 (N_4595,N_3290,N_3051);
or U4596 (N_4596,N_2532,N_2732);
nand U4597 (N_4597,N_2633,N_3327);
and U4598 (N_4598,N_2464,N_2738);
nor U4599 (N_4599,N_3001,N_3239);
or U4600 (N_4600,N_2945,N_2585);
nand U4601 (N_4601,N_3243,N_3044);
nand U4602 (N_4602,N_3364,N_2441);
and U4603 (N_4603,N_2569,N_3414);
nor U4604 (N_4604,N_3054,N_2980);
and U4605 (N_4605,N_2608,N_3215);
nor U4606 (N_4606,N_3539,N_2496);
or U4607 (N_4607,N_2490,N_3067);
or U4608 (N_4608,N_3298,N_2780);
nand U4609 (N_4609,N_2517,N_2704);
nor U4610 (N_4610,N_3279,N_2837);
nor U4611 (N_4611,N_3429,N_3046);
nand U4612 (N_4612,N_2549,N_2847);
xnor U4613 (N_4613,N_2516,N_2729);
xor U4614 (N_4614,N_3008,N_3108);
or U4615 (N_4615,N_2879,N_3440);
xnor U4616 (N_4616,N_3542,N_2684);
nor U4617 (N_4617,N_3220,N_3379);
or U4618 (N_4618,N_3093,N_2787);
nand U4619 (N_4619,N_3177,N_3374);
xor U4620 (N_4620,N_3171,N_3598);
and U4621 (N_4621,N_3185,N_2901);
nor U4622 (N_4622,N_2502,N_2716);
and U4623 (N_4623,N_3319,N_2493);
or U4624 (N_4624,N_3007,N_2449);
nor U4625 (N_4625,N_2715,N_2660);
nor U4626 (N_4626,N_3367,N_2686);
nor U4627 (N_4627,N_3471,N_2789);
nor U4628 (N_4628,N_2478,N_3310);
nand U4629 (N_4629,N_2570,N_3427);
nand U4630 (N_4630,N_3091,N_3075);
nor U4631 (N_4631,N_2852,N_3576);
xnor U4632 (N_4632,N_2495,N_2768);
or U4633 (N_4633,N_3011,N_2928);
xor U4634 (N_4634,N_3101,N_2779);
or U4635 (N_4635,N_3310,N_2539);
nand U4636 (N_4636,N_3389,N_2941);
nand U4637 (N_4637,N_3422,N_2460);
and U4638 (N_4638,N_3307,N_3592);
or U4639 (N_4639,N_3291,N_3325);
nor U4640 (N_4640,N_3418,N_2485);
nor U4641 (N_4641,N_3236,N_3418);
nor U4642 (N_4642,N_2499,N_2898);
and U4643 (N_4643,N_3053,N_3384);
and U4644 (N_4644,N_3169,N_2579);
nor U4645 (N_4645,N_3166,N_3512);
nand U4646 (N_4646,N_2530,N_2450);
nand U4647 (N_4647,N_2931,N_2524);
xnor U4648 (N_4648,N_3011,N_2409);
nor U4649 (N_4649,N_3121,N_3403);
nor U4650 (N_4650,N_2601,N_3070);
and U4651 (N_4651,N_3028,N_3135);
and U4652 (N_4652,N_2735,N_3170);
or U4653 (N_4653,N_3191,N_2969);
nor U4654 (N_4654,N_3099,N_2649);
nor U4655 (N_4655,N_3257,N_2860);
and U4656 (N_4656,N_3310,N_3085);
nor U4657 (N_4657,N_3076,N_3110);
nor U4658 (N_4658,N_3359,N_3549);
nor U4659 (N_4659,N_3187,N_2528);
nor U4660 (N_4660,N_3396,N_2970);
and U4661 (N_4661,N_2595,N_3234);
or U4662 (N_4662,N_3066,N_2747);
nand U4663 (N_4663,N_2688,N_3235);
nand U4664 (N_4664,N_3068,N_3387);
and U4665 (N_4665,N_2871,N_2660);
nand U4666 (N_4666,N_2436,N_3352);
xnor U4667 (N_4667,N_3386,N_3458);
xnor U4668 (N_4668,N_3128,N_3370);
xor U4669 (N_4669,N_3591,N_2675);
and U4670 (N_4670,N_2919,N_2738);
nor U4671 (N_4671,N_2990,N_2795);
xnor U4672 (N_4672,N_3406,N_3118);
xor U4673 (N_4673,N_3434,N_2853);
nor U4674 (N_4674,N_3308,N_2845);
nand U4675 (N_4675,N_2429,N_3148);
nor U4676 (N_4676,N_2550,N_2800);
nor U4677 (N_4677,N_2646,N_2749);
nor U4678 (N_4678,N_3408,N_2838);
xnor U4679 (N_4679,N_2918,N_3226);
nand U4680 (N_4680,N_2792,N_3259);
nor U4681 (N_4681,N_3174,N_2531);
and U4682 (N_4682,N_2927,N_3107);
xnor U4683 (N_4683,N_2524,N_3371);
xor U4684 (N_4684,N_3087,N_3441);
and U4685 (N_4685,N_2431,N_3308);
xnor U4686 (N_4686,N_2925,N_3131);
xnor U4687 (N_4687,N_2583,N_2477);
xor U4688 (N_4688,N_2851,N_2754);
xor U4689 (N_4689,N_3469,N_3091);
nand U4690 (N_4690,N_3521,N_2932);
nor U4691 (N_4691,N_2978,N_3076);
and U4692 (N_4692,N_2611,N_2607);
and U4693 (N_4693,N_3503,N_2899);
or U4694 (N_4694,N_2454,N_2912);
xor U4695 (N_4695,N_2883,N_3448);
or U4696 (N_4696,N_2686,N_2874);
or U4697 (N_4697,N_3154,N_2970);
xnor U4698 (N_4698,N_3516,N_3351);
nor U4699 (N_4699,N_3312,N_2907);
nand U4700 (N_4700,N_3242,N_3596);
nand U4701 (N_4701,N_3069,N_2516);
nor U4702 (N_4702,N_2489,N_3353);
and U4703 (N_4703,N_2576,N_3559);
and U4704 (N_4704,N_3491,N_3018);
nand U4705 (N_4705,N_2452,N_2553);
nor U4706 (N_4706,N_2653,N_2918);
nor U4707 (N_4707,N_2569,N_2937);
nor U4708 (N_4708,N_2842,N_2607);
nand U4709 (N_4709,N_3325,N_3461);
nor U4710 (N_4710,N_3043,N_2954);
nand U4711 (N_4711,N_3238,N_2795);
nor U4712 (N_4712,N_2857,N_2557);
nor U4713 (N_4713,N_3075,N_3014);
nand U4714 (N_4714,N_3106,N_2713);
xnor U4715 (N_4715,N_2744,N_2431);
nor U4716 (N_4716,N_3001,N_3000);
nor U4717 (N_4717,N_3029,N_2860);
nor U4718 (N_4718,N_2927,N_2839);
and U4719 (N_4719,N_3485,N_2838);
nor U4720 (N_4720,N_2613,N_3355);
or U4721 (N_4721,N_3096,N_2915);
and U4722 (N_4722,N_2850,N_3193);
nand U4723 (N_4723,N_2935,N_3000);
and U4724 (N_4724,N_2451,N_2813);
nand U4725 (N_4725,N_3286,N_2607);
nor U4726 (N_4726,N_2529,N_2522);
and U4727 (N_4727,N_2782,N_2846);
nand U4728 (N_4728,N_2613,N_2904);
nor U4729 (N_4729,N_3500,N_2464);
nand U4730 (N_4730,N_2437,N_2840);
nor U4731 (N_4731,N_3023,N_3126);
nor U4732 (N_4732,N_2625,N_3436);
nor U4733 (N_4733,N_2532,N_3097);
xnor U4734 (N_4734,N_3566,N_2763);
xnor U4735 (N_4735,N_2541,N_3107);
and U4736 (N_4736,N_2698,N_3408);
or U4737 (N_4737,N_3331,N_2568);
and U4738 (N_4738,N_2589,N_2880);
and U4739 (N_4739,N_2527,N_3218);
nand U4740 (N_4740,N_2916,N_2876);
or U4741 (N_4741,N_3116,N_3354);
nand U4742 (N_4742,N_3379,N_3158);
xnor U4743 (N_4743,N_3080,N_3246);
and U4744 (N_4744,N_2615,N_3141);
nand U4745 (N_4745,N_2878,N_2953);
nor U4746 (N_4746,N_3093,N_3252);
or U4747 (N_4747,N_2766,N_3327);
or U4748 (N_4748,N_2590,N_3159);
nor U4749 (N_4749,N_2736,N_3219);
or U4750 (N_4750,N_2984,N_2602);
and U4751 (N_4751,N_3418,N_3458);
nor U4752 (N_4752,N_2482,N_3283);
or U4753 (N_4753,N_2645,N_2654);
or U4754 (N_4754,N_2735,N_2720);
nand U4755 (N_4755,N_3562,N_3021);
and U4756 (N_4756,N_3569,N_3405);
xnor U4757 (N_4757,N_2709,N_3296);
nor U4758 (N_4758,N_2749,N_2881);
and U4759 (N_4759,N_2548,N_2695);
nor U4760 (N_4760,N_3154,N_3292);
nor U4761 (N_4761,N_3512,N_3535);
or U4762 (N_4762,N_3155,N_2578);
nor U4763 (N_4763,N_2473,N_2862);
and U4764 (N_4764,N_3074,N_3554);
xor U4765 (N_4765,N_3036,N_3055);
nor U4766 (N_4766,N_2471,N_2949);
nand U4767 (N_4767,N_3055,N_2782);
nor U4768 (N_4768,N_3229,N_3320);
xnor U4769 (N_4769,N_3333,N_3231);
nor U4770 (N_4770,N_2566,N_2449);
or U4771 (N_4771,N_3051,N_3538);
xnor U4772 (N_4772,N_3085,N_3211);
nor U4773 (N_4773,N_2692,N_2671);
nor U4774 (N_4774,N_3571,N_2908);
nor U4775 (N_4775,N_2774,N_3162);
or U4776 (N_4776,N_2920,N_3172);
nand U4777 (N_4777,N_2549,N_2938);
nand U4778 (N_4778,N_3437,N_2428);
or U4779 (N_4779,N_2668,N_2495);
or U4780 (N_4780,N_2410,N_3001);
nor U4781 (N_4781,N_2794,N_3082);
xor U4782 (N_4782,N_3370,N_3228);
nand U4783 (N_4783,N_3186,N_2825);
and U4784 (N_4784,N_3320,N_2452);
or U4785 (N_4785,N_3049,N_2569);
and U4786 (N_4786,N_2907,N_3092);
or U4787 (N_4787,N_3275,N_3284);
and U4788 (N_4788,N_2990,N_2744);
nand U4789 (N_4789,N_3165,N_3256);
or U4790 (N_4790,N_2966,N_2555);
xor U4791 (N_4791,N_3080,N_2672);
xor U4792 (N_4792,N_3402,N_2786);
and U4793 (N_4793,N_3450,N_3005);
or U4794 (N_4794,N_3277,N_2813);
and U4795 (N_4795,N_3524,N_3139);
nor U4796 (N_4796,N_3589,N_2574);
nor U4797 (N_4797,N_3029,N_3190);
xnor U4798 (N_4798,N_3443,N_2685);
and U4799 (N_4799,N_3510,N_2476);
nand U4800 (N_4800,N_4255,N_3964);
nand U4801 (N_4801,N_4219,N_3673);
or U4802 (N_4802,N_3952,N_4642);
xor U4803 (N_4803,N_4032,N_4726);
nor U4804 (N_4804,N_4061,N_4363);
nand U4805 (N_4805,N_4762,N_3674);
nor U4806 (N_4806,N_4586,N_4253);
or U4807 (N_4807,N_4756,N_4095);
nand U4808 (N_4808,N_4536,N_4393);
nand U4809 (N_4809,N_3903,N_4161);
and U4810 (N_4810,N_4239,N_4070);
xnor U4811 (N_4811,N_3758,N_3751);
and U4812 (N_4812,N_4582,N_4330);
and U4813 (N_4813,N_4394,N_4606);
or U4814 (N_4814,N_4758,N_4538);
nand U4815 (N_4815,N_4662,N_4052);
nor U4816 (N_4816,N_4595,N_4531);
or U4817 (N_4817,N_4130,N_4735);
or U4818 (N_4818,N_3830,N_4764);
or U4819 (N_4819,N_3995,N_4710);
xnor U4820 (N_4820,N_4521,N_4366);
and U4821 (N_4821,N_3852,N_3868);
or U4822 (N_4822,N_4146,N_3948);
and U4823 (N_4823,N_3794,N_3780);
nand U4824 (N_4824,N_4262,N_4285);
and U4825 (N_4825,N_4499,N_4315);
and U4826 (N_4826,N_3963,N_3657);
nor U4827 (N_4827,N_4411,N_3768);
nor U4828 (N_4828,N_3601,N_4769);
nand U4829 (N_4829,N_4122,N_4541);
and U4830 (N_4830,N_3842,N_4429);
nor U4831 (N_4831,N_3623,N_3775);
nor U4832 (N_4832,N_4016,N_4216);
and U4833 (N_4833,N_3772,N_4208);
xor U4834 (N_4834,N_4400,N_3992);
and U4835 (N_4835,N_3881,N_4086);
nand U4836 (N_4836,N_3695,N_4263);
xor U4837 (N_4837,N_3813,N_3985);
xnor U4838 (N_4838,N_4082,N_3606);
or U4839 (N_4839,N_4724,N_4204);
nor U4840 (N_4840,N_4229,N_3764);
nor U4841 (N_4841,N_4583,N_4490);
or U4842 (N_4842,N_3987,N_4527);
nand U4843 (N_4843,N_4092,N_4381);
nor U4844 (N_4844,N_4534,N_4029);
nand U4845 (N_4845,N_3997,N_3901);
xnor U4846 (N_4846,N_4269,N_4175);
or U4847 (N_4847,N_4057,N_4702);
or U4848 (N_4848,N_4231,N_4437);
nor U4849 (N_4849,N_4080,N_4442);
or U4850 (N_4850,N_4607,N_3787);
and U4851 (N_4851,N_3883,N_4312);
xor U4852 (N_4852,N_4410,N_4633);
xor U4853 (N_4853,N_3640,N_3954);
xor U4854 (N_4854,N_4605,N_4386);
xnor U4855 (N_4855,N_4010,N_3940);
or U4856 (N_4856,N_4151,N_3799);
nand U4857 (N_4857,N_4436,N_4578);
xor U4858 (N_4858,N_4213,N_4604);
nor U4859 (N_4859,N_4439,N_4569);
nand U4860 (N_4860,N_4611,N_4709);
xor U4861 (N_4861,N_4500,N_4037);
and U4862 (N_4862,N_4600,N_4031);
nand U4863 (N_4863,N_4640,N_4347);
or U4864 (N_4864,N_3730,N_4301);
nand U4865 (N_4865,N_3839,N_4528);
nor U4866 (N_4866,N_3976,N_3982);
and U4867 (N_4867,N_4722,N_4162);
nor U4868 (N_4868,N_3689,N_3624);
nor U4869 (N_4869,N_4355,N_4030);
nor U4870 (N_4870,N_4336,N_4214);
nand U4871 (N_4871,N_4547,N_4223);
nor U4872 (N_4872,N_4416,N_3728);
nor U4873 (N_4873,N_3862,N_4668);
nand U4874 (N_4874,N_4178,N_4518);
nand U4875 (N_4875,N_4243,N_4091);
xnor U4876 (N_4876,N_4725,N_3650);
or U4877 (N_4877,N_4079,N_4050);
or U4878 (N_4878,N_4241,N_4324);
xnor U4879 (N_4879,N_3704,N_4711);
and U4880 (N_4880,N_4357,N_3972);
or U4881 (N_4881,N_4172,N_4261);
or U4882 (N_4882,N_3899,N_3653);
nor U4883 (N_4883,N_4690,N_4124);
and U4884 (N_4884,N_4636,N_3757);
xor U4885 (N_4885,N_4560,N_3652);
and U4886 (N_4886,N_4034,N_3840);
and U4887 (N_4887,N_3691,N_4071);
nor U4888 (N_4888,N_4542,N_4483);
nor U4889 (N_4889,N_4723,N_4486);
nor U4890 (N_4890,N_4383,N_4040);
xor U4891 (N_4891,N_3721,N_3988);
xor U4892 (N_4892,N_3861,N_3918);
nor U4893 (N_4893,N_4740,N_3743);
nand U4894 (N_4894,N_4217,N_4680);
or U4895 (N_4895,N_4593,N_4712);
nand U4896 (N_4896,N_4648,N_4478);
and U4897 (N_4897,N_4549,N_4054);
xor U4898 (N_4898,N_3661,N_4280);
nand U4899 (N_4899,N_4247,N_3894);
and U4900 (N_4900,N_4323,N_4691);
xor U4901 (N_4901,N_3878,N_4007);
or U4902 (N_4902,N_4718,N_3677);
or U4903 (N_4903,N_4211,N_3701);
xnor U4904 (N_4904,N_3639,N_3891);
and U4905 (N_4905,N_4579,N_4373);
nor U4906 (N_4906,N_4188,N_3684);
and U4907 (N_4907,N_3938,N_3675);
or U4908 (N_4908,N_4065,N_3970);
xor U4909 (N_4909,N_4069,N_3798);
and U4910 (N_4910,N_4548,N_3932);
nand U4911 (N_4911,N_4568,N_3801);
xor U4912 (N_4912,N_3824,N_4265);
or U4913 (N_4913,N_3714,N_3655);
xor U4914 (N_4914,N_3867,N_3649);
nand U4915 (N_4915,N_4097,N_4566);
xor U4916 (N_4916,N_3685,N_4327);
nor U4917 (N_4917,N_4795,N_3943);
xor U4918 (N_4918,N_4658,N_4730);
nand U4919 (N_4919,N_3810,N_4205);
or U4920 (N_4920,N_4591,N_3958);
or U4921 (N_4921,N_4321,N_3729);
or U4922 (N_4922,N_4099,N_3771);
and U4923 (N_4923,N_3734,N_4655);
nand U4924 (N_4924,N_3807,N_3666);
or U4925 (N_4925,N_3828,N_4290);
nor U4926 (N_4926,N_4523,N_4625);
or U4927 (N_4927,N_4046,N_4440);
and U4928 (N_4928,N_3866,N_3694);
nor U4929 (N_4929,N_4176,N_4457);
and U4930 (N_4930,N_3908,N_4182);
nand U4931 (N_4931,N_4294,N_4344);
or U4932 (N_4932,N_4173,N_4484);
and U4933 (N_4933,N_4152,N_3740);
and U4934 (N_4934,N_4398,N_3825);
nand U4935 (N_4935,N_4314,N_4624);
and U4936 (N_4936,N_3919,N_4326);
nor U4937 (N_4937,N_4369,N_4288);
nor U4938 (N_4938,N_3617,N_4281);
and U4939 (N_4939,N_3863,N_4520);
or U4940 (N_4940,N_3804,N_4035);
xor U4941 (N_4941,N_3817,N_4708);
or U4942 (N_4942,N_3800,N_4529);
nor U4943 (N_4943,N_4663,N_4317);
and U4944 (N_4944,N_4438,N_3784);
nand U4945 (N_4945,N_4649,N_3603);
and U4946 (N_4946,N_4351,N_4653);
nand U4947 (N_4947,N_4445,N_3697);
nor U4948 (N_4948,N_4698,N_4617);
nor U4949 (N_4949,N_3924,N_4696);
nand U4950 (N_4950,N_4657,N_3776);
nand U4951 (N_4951,N_3897,N_4169);
nand U4952 (N_4952,N_4333,N_4179);
and U4953 (N_4953,N_4135,N_4372);
xnor U4954 (N_4954,N_4537,N_4378);
or U4955 (N_4955,N_4230,N_3662);
nor U4956 (N_4956,N_4044,N_4361);
nand U4957 (N_4957,N_4707,N_4405);
xnor U4958 (N_4958,N_3769,N_4557);
nor U4959 (N_4959,N_3746,N_3898);
or U4960 (N_4960,N_4206,N_3980);
and U4961 (N_4961,N_4268,N_3609);
xnor U4962 (N_4962,N_4299,N_4632);
xnor U4963 (N_4963,N_3869,N_3837);
nand U4964 (N_4964,N_3951,N_4003);
and U4965 (N_4965,N_4187,N_3942);
and U4966 (N_4966,N_3686,N_4433);
nand U4967 (N_4967,N_3838,N_4119);
or U4968 (N_4968,N_3887,N_3632);
and U4969 (N_4969,N_4417,N_4127);
xnor U4970 (N_4970,N_4687,N_3966);
nand U4971 (N_4971,N_4626,N_4209);
and U4972 (N_4972,N_4013,N_4258);
or U4973 (N_4973,N_3950,N_4788);
nand U4974 (N_4974,N_4441,N_4492);
and U4975 (N_4975,N_3687,N_4038);
and U4976 (N_4976,N_3809,N_3871);
nand U4977 (N_4977,N_3880,N_3930);
and U4978 (N_4978,N_4513,N_4570);
nand U4979 (N_4979,N_4062,N_3710);
nand U4980 (N_4980,N_4706,N_4123);
nor U4981 (N_4981,N_3703,N_4248);
xnor U4982 (N_4982,N_4613,N_4011);
xor U4983 (N_4983,N_4664,N_4621);
or U4984 (N_4984,N_4546,N_4510);
nor U4985 (N_4985,N_4670,N_4249);
nand U4986 (N_4986,N_4755,N_4390);
or U4987 (N_4987,N_3795,N_3907);
nor U4988 (N_4988,N_4310,N_3879);
and U4989 (N_4989,N_3818,N_3731);
nand U4990 (N_4990,N_4550,N_4641);
nand U4991 (N_4991,N_4462,N_3886);
and U4992 (N_4992,N_4777,N_4671);
or U4993 (N_4993,N_4020,N_3763);
xnor U4994 (N_4994,N_4564,N_4472);
xnor U4995 (N_4995,N_4444,N_4218);
nand U4996 (N_4996,N_4328,N_4341);
xnor U4997 (N_4997,N_4374,N_4667);
nor U4998 (N_4998,N_3600,N_3767);
nor U4999 (N_4999,N_3984,N_4332);
nand U5000 (N_5000,N_4058,N_4283);
nor U5001 (N_5001,N_4073,N_3668);
or U5002 (N_5002,N_4496,N_4602);
xor U5003 (N_5003,N_4553,N_4552);
xnor U5004 (N_5004,N_4264,N_4337);
nand U5005 (N_5005,N_4747,N_4753);
nand U5006 (N_5006,N_4587,N_4556);
nor U5007 (N_5007,N_3916,N_3974);
nor U5008 (N_5008,N_4107,N_4460);
nor U5009 (N_5009,N_4620,N_3900);
nor U5010 (N_5010,N_3853,N_3856);
xor U5011 (N_5011,N_3658,N_4103);
or U5012 (N_5012,N_4459,N_4661);
or U5013 (N_5013,N_3616,N_4503);
or U5014 (N_5014,N_4126,N_3742);
and U5015 (N_5015,N_4155,N_4746);
nor U5016 (N_5016,N_4609,N_3688);
and U5017 (N_5017,N_3773,N_4000);
nand U5018 (N_5018,N_3629,N_3875);
or U5019 (N_5019,N_3766,N_4488);
nor U5020 (N_5020,N_4192,N_4237);
nor U5021 (N_5021,N_4631,N_4259);
nand U5022 (N_5022,N_4701,N_4049);
xnor U5023 (N_5023,N_4509,N_3857);
or U5024 (N_5024,N_4053,N_3739);
nand U5025 (N_5025,N_4036,N_3744);
nor U5026 (N_5026,N_4105,N_3915);
and U5027 (N_5027,N_4200,N_3611);
or U5028 (N_5028,N_3877,N_4193);
or U5029 (N_5029,N_3789,N_4647);
nor U5030 (N_5030,N_4791,N_4102);
and U5031 (N_5031,N_4563,N_4171);
xnor U5032 (N_5032,N_4512,N_4311);
or U5033 (N_5033,N_3962,N_4308);
and U5034 (N_5034,N_4027,N_3882);
nor U5035 (N_5035,N_4212,N_4271);
or U5036 (N_5036,N_4743,N_3820);
or U5037 (N_5037,N_4651,N_3893);
nor U5038 (N_5038,N_4425,N_4463);
xnor U5039 (N_5039,N_4286,N_4683);
nor U5040 (N_5040,N_4257,N_4768);
or U5041 (N_5041,N_4754,N_3865);
or U5042 (N_5042,N_4493,N_4619);
and U5043 (N_5043,N_3874,N_4678);
nand U5044 (N_5044,N_4409,N_3725);
or U5045 (N_5045,N_4284,N_4396);
and U5046 (N_5046,N_4422,N_3910);
and U5047 (N_5047,N_3849,N_3859);
nand U5048 (N_5048,N_3864,N_4432);
xnor U5049 (N_5049,N_4201,N_3612);
or U5050 (N_5050,N_4018,N_4427);
nor U5051 (N_5051,N_4395,N_4138);
and U5052 (N_5052,N_4561,N_4502);
or U5053 (N_5053,N_4158,N_4544);
or U5054 (N_5054,N_3917,N_4190);
and U5055 (N_5055,N_4266,N_4598);
nand U5056 (N_5056,N_3831,N_4506);
and U5057 (N_5057,N_3802,N_4716);
xnor U5058 (N_5058,N_4421,N_4392);
and U5059 (N_5059,N_3636,N_4234);
or U5060 (N_5060,N_4423,N_4728);
or U5061 (N_5061,N_4732,N_4183);
xor U5062 (N_5062,N_4644,N_3797);
and U5063 (N_5063,N_3929,N_4166);
and U5064 (N_5064,N_4603,N_4116);
nand U5065 (N_5065,N_4379,N_3613);
nor U5066 (N_5066,N_4084,N_4799);
xnor U5067 (N_5067,N_4741,N_4491);
or U5068 (N_5068,N_4345,N_4385);
nand U5069 (N_5069,N_4026,N_4665);
nor U5070 (N_5070,N_3975,N_3656);
xnor U5071 (N_5071,N_3783,N_3778);
nand U5072 (N_5072,N_3659,N_4713);
nor U5073 (N_5073,N_4362,N_4589);
xor U5074 (N_5074,N_4376,N_4770);
and U5075 (N_5075,N_4794,N_3884);
nor U5076 (N_5076,N_3607,N_4154);
xor U5077 (N_5077,N_3667,N_4309);
or U5078 (N_5078,N_4227,N_4674);
nand U5079 (N_5079,N_4339,N_4380);
or U5080 (N_5080,N_4128,N_3850);
and U5081 (N_5081,N_3727,N_4739);
and U5082 (N_5082,N_4516,N_3812);
nor U5083 (N_5083,N_4094,N_3716);
nand U5084 (N_5084,N_4751,N_3705);
nand U5085 (N_5085,N_3712,N_4508);
and U5086 (N_5086,N_3835,N_4535);
nand U5087 (N_5087,N_4786,N_4573);
or U5088 (N_5088,N_3790,N_3937);
and U5089 (N_5089,N_4594,N_4562);
or U5090 (N_5090,N_3990,N_4643);
or U5091 (N_5091,N_4614,N_3643);
nor U5092 (N_5092,N_4303,N_4414);
nand U5093 (N_5093,N_4420,N_4015);
nor U5094 (N_5094,N_4377,N_4108);
xnor U5095 (N_5095,N_4199,N_4325);
nand U5096 (N_5096,N_4615,N_4164);
xnor U5097 (N_5097,N_4470,N_3633);
and U5098 (N_5098,N_4693,N_3814);
nor U5099 (N_5099,N_4412,N_3692);
nand U5100 (N_5100,N_4540,N_4195);
and U5101 (N_5101,N_4101,N_4068);
and U5102 (N_5102,N_4571,N_3717);
xor U5103 (N_5103,N_3793,N_4464);
xnor U5104 (N_5104,N_3827,N_4646);
nor U5105 (N_5105,N_4300,N_3637);
nor U5106 (N_5106,N_4497,N_4250);
and U5107 (N_5107,N_3872,N_3774);
nand U5108 (N_5108,N_3702,N_3620);
xor U5109 (N_5109,N_4186,N_4783);
or U5110 (N_5110,N_4004,N_4485);
or U5111 (N_5111,N_4120,N_4349);
nand U5112 (N_5112,N_4767,N_3671);
nor U5113 (N_5113,N_4222,N_4699);
and U5114 (N_5114,N_4451,N_4404);
and U5115 (N_5115,N_4477,N_4215);
nor U5116 (N_5116,N_4334,N_4514);
nor U5117 (N_5117,N_3682,N_4532);
xnor U5118 (N_5118,N_3890,N_3978);
nor U5119 (N_5119,N_4745,N_3833);
or U5120 (N_5120,N_4163,N_4495);
or U5121 (N_5121,N_4525,N_4399);
nand U5122 (N_5122,N_4370,N_3902);
xor U5123 (N_5123,N_4139,N_4639);
or U5124 (N_5124,N_4584,N_4041);
nand U5125 (N_5125,N_3888,N_3645);
nor U5126 (N_5126,N_4543,N_4466);
nand U5127 (N_5127,N_3933,N_4313);
nor U5128 (N_5128,N_3770,N_4220);
and U5129 (N_5129,N_4356,N_4511);
xnor U5130 (N_5130,N_4279,N_4715);
nor U5131 (N_5131,N_4059,N_4577);
nor U5132 (N_5132,N_3967,N_4637);
nand U5133 (N_5133,N_3870,N_4047);
and U5134 (N_5134,N_3718,N_3843);
and U5135 (N_5135,N_4289,N_4689);
and U5136 (N_5136,N_3991,N_4447);
nor U5137 (N_5137,N_4067,N_4159);
xnor U5138 (N_5138,N_3905,N_4630);
and U5139 (N_5139,N_4100,N_4426);
or U5140 (N_5140,N_3847,N_4153);
or U5141 (N_5141,N_4242,N_3854);
and U5142 (N_5142,N_4150,N_4367);
or U5143 (N_5143,N_4719,N_4467);
nor U5144 (N_5144,N_4505,N_4350);
xnor U5145 (N_5145,N_4305,N_3885);
nand U5146 (N_5146,N_4793,N_3841);
and U5147 (N_5147,N_4471,N_3604);
and U5148 (N_5148,N_4225,N_4145);
xnor U5149 (N_5149,N_4522,N_4087);
nand U5150 (N_5150,N_3680,N_4567);
nor U5151 (N_5151,N_4185,N_4254);
xnor U5152 (N_5152,N_3858,N_4686);
nand U5153 (N_5153,N_4494,N_3977);
xnor U5154 (N_5154,N_4077,N_4453);
and U5155 (N_5155,N_4202,N_3996);
nor U5156 (N_5156,N_4074,N_4006);
nand U5157 (N_5157,N_4781,N_4652);
nor U5158 (N_5158,N_3786,N_4267);
or U5159 (N_5159,N_4700,N_3777);
nand U5160 (N_5160,N_4001,N_4140);
xnor U5161 (N_5161,N_3626,N_4260);
nand U5162 (N_5162,N_4302,N_3726);
nor U5163 (N_5163,N_3646,N_3998);
nor U5164 (N_5164,N_3896,N_3851);
or U5165 (N_5165,N_3848,N_4142);
or U5166 (N_5166,N_4634,N_3922);
and U5167 (N_5167,N_4558,N_4295);
and U5168 (N_5168,N_4012,N_4331);
and U5169 (N_5169,N_4098,N_3914);
and U5170 (N_5170,N_4565,N_4752);
xnor U5171 (N_5171,N_4413,N_4704);
and U5172 (N_5172,N_3738,N_4076);
and U5173 (N_5173,N_3755,N_4610);
nand U5174 (N_5174,N_3953,N_4236);
or U5175 (N_5175,N_4402,N_4282);
nand U5176 (N_5176,N_4075,N_3911);
xnor U5177 (N_5177,N_4669,N_4434);
nor U5178 (N_5178,N_3737,N_4352);
and U5179 (N_5179,N_3844,N_4117);
and U5180 (N_5180,N_4343,N_4045);
and U5181 (N_5181,N_4060,N_3634);
and U5182 (N_5182,N_4759,N_4622);
nand U5183 (N_5183,N_4189,N_4384);
or U5184 (N_5184,N_3765,N_4601);
nand U5185 (N_5185,N_3961,N_4194);
nor U5186 (N_5186,N_4729,N_3733);
and U5187 (N_5187,N_4742,N_3663);
nand U5188 (N_5188,N_4014,N_3756);
xor U5189 (N_5189,N_4293,N_4141);
nand U5190 (N_5190,N_4585,N_3994);
or U5191 (N_5191,N_4545,N_4760);
nor U5192 (N_5192,N_4306,N_4480);
and U5193 (N_5193,N_4597,N_4005);
nor U5194 (N_5194,N_4782,N_3676);
nor U5195 (N_5195,N_4524,N_4714);
or U5196 (N_5196,N_4063,N_4277);
nand U5197 (N_5197,N_4226,N_4428);
nor U5198 (N_5198,N_4210,N_3904);
and U5199 (N_5199,N_4115,N_3608);
and U5200 (N_5200,N_4415,N_3696);
xnor U5201 (N_5201,N_4727,N_4623);
nor U5202 (N_5202,N_4489,N_4033);
or U5203 (N_5203,N_4482,N_3679);
xor U5204 (N_5204,N_4748,N_4517);
or U5205 (N_5205,N_4008,N_4684);
nor U5206 (N_5206,N_3615,N_4273);
xnor U5207 (N_5207,N_3969,N_3762);
and U5208 (N_5208,N_3973,N_4359);
and U5209 (N_5209,N_3678,N_3821);
and U5210 (N_5210,N_4043,N_3855);
nand U5211 (N_5211,N_4580,N_4526);
nand U5212 (N_5212,N_4787,N_4672);
xnor U5213 (N_5213,N_4365,N_3711);
xor U5214 (N_5214,N_3681,N_4318);
nor U5215 (N_5215,N_4197,N_4270);
or U5216 (N_5216,N_4391,N_4757);
and U5217 (N_5217,N_4382,N_3741);
or U5218 (N_5218,N_3644,N_4731);
nand U5219 (N_5219,N_4406,N_4304);
xor U5220 (N_5220,N_4114,N_3693);
and U5221 (N_5221,N_4792,N_3654);
and U5222 (N_5222,N_3631,N_3683);
or U5223 (N_5223,N_4203,N_4507);
nand U5224 (N_5224,N_4449,N_4371);
nor U5225 (N_5225,N_4654,N_4112);
or U5226 (N_5226,N_3955,N_3906);
nor U5227 (N_5227,N_4468,N_4397);
nor U5228 (N_5228,N_3806,N_4473);
or U5229 (N_5229,N_4340,N_3660);
xnor U5230 (N_5230,N_4168,N_3822);
and U5231 (N_5231,N_4533,N_4125);
or U5232 (N_5232,N_4275,N_3621);
nor U5233 (N_5233,N_4424,N_4354);
nor U5234 (N_5234,N_4085,N_3619);
nand U5235 (N_5235,N_4780,N_3889);
xor U5236 (N_5236,N_4048,N_3960);
and U5237 (N_5237,N_4348,N_4184);
nand U5238 (N_5238,N_4784,N_3876);
and U5239 (N_5239,N_4773,N_3805);
nand U5240 (N_5240,N_4430,N_3796);
or U5241 (N_5241,N_3638,N_3947);
nand U5242 (N_5242,N_3993,N_3672);
xor U5243 (N_5243,N_3754,N_3834);
and U5244 (N_5244,N_4096,N_4297);
nor U5245 (N_5245,N_4198,N_4307);
nand U5246 (N_5246,N_4763,N_3956);
nand U5247 (N_5247,N_4147,N_4056);
xor U5248 (N_5248,N_3845,N_4118);
or U5249 (N_5249,N_4110,N_4454);
nor U5250 (N_5250,N_4688,N_4167);
or U5251 (N_5251,N_3926,N_3836);
nand U5252 (N_5252,N_4252,N_4681);
xnor U5253 (N_5253,N_4245,N_4272);
nor U5254 (N_5254,N_4734,N_3779);
nand U5255 (N_5255,N_3941,N_4089);
nor U5256 (N_5256,N_4233,N_4501);
xor U5257 (N_5257,N_3829,N_3670);
xnor U5258 (N_5258,N_4274,N_4675);
nand U5259 (N_5259,N_4244,N_4338);
nor U5260 (N_5260,N_3913,N_3699);
and U5261 (N_5261,N_3792,N_4629);
nand U5262 (N_5262,N_3735,N_4469);
xnor U5263 (N_5263,N_4581,N_3720);
nand U5264 (N_5264,N_4720,N_4024);
xnor U5265 (N_5265,N_4738,N_4465);
nor U5266 (N_5266,N_4487,N_4682);
xnor U5267 (N_5267,N_3707,N_4551);
xnor U5268 (N_5268,N_3664,N_4132);
or U5269 (N_5269,N_4143,N_4458);
or U5270 (N_5270,N_4789,N_3723);
or U5271 (N_5271,N_4666,N_4335);
nor U5272 (N_5272,N_4450,N_4796);
xor U5273 (N_5273,N_4387,N_3921);
nand U5274 (N_5274,N_3625,N_3920);
or U5275 (N_5275,N_3651,N_4576);
nand U5276 (N_5276,N_4695,N_4170);
nor U5277 (N_5277,N_4618,N_4083);
or U5278 (N_5278,N_3709,N_4017);
nand U5279 (N_5279,N_4435,N_3752);
and U5280 (N_5280,N_4446,N_4717);
nor U5281 (N_5281,N_4228,N_3927);
or U5282 (N_5282,N_4685,N_3724);
and U5283 (N_5283,N_3946,N_3753);
xnor U5284 (N_5284,N_4109,N_3949);
and U5285 (N_5285,N_4765,N_4019);
or U5286 (N_5286,N_4456,N_3745);
and U5287 (N_5287,N_4287,N_4443);
nand U5288 (N_5288,N_4181,N_4705);
nand U5289 (N_5289,N_3750,N_4418);
nand U5290 (N_5290,N_3759,N_4256);
xor U5291 (N_5291,N_4790,N_3791);
and U5292 (N_5292,N_4461,N_3999);
and U5293 (N_5293,N_4408,N_4093);
nor U5294 (N_5294,N_4474,N_4174);
nor U5295 (N_5295,N_4419,N_4572);
nand U5296 (N_5296,N_4656,N_4021);
nand U5297 (N_5297,N_3614,N_3939);
and U5298 (N_5298,N_4064,N_4555);
or U5299 (N_5299,N_4028,N_3719);
and U5300 (N_5300,N_4737,N_3965);
or U5301 (N_5301,N_4679,N_4554);
nand U5302 (N_5302,N_4276,N_3648);
and U5303 (N_5303,N_3892,N_3749);
nor U5304 (N_5304,N_4559,N_4530);
nor U5305 (N_5305,N_4616,N_3722);
xnor U5306 (N_5306,N_3983,N_4144);
or U5307 (N_5307,N_3923,N_4081);
or U5308 (N_5308,N_4479,N_4246);
nand U5309 (N_5309,N_4134,N_3873);
xor U5310 (N_5310,N_4407,N_4235);
and U5311 (N_5311,N_4196,N_3936);
or U5312 (N_5312,N_4599,N_3761);
or U5313 (N_5313,N_4645,N_4240);
nand U5314 (N_5314,N_4232,N_4650);
nand U5315 (N_5315,N_4761,N_4149);
and U5316 (N_5316,N_4612,N_4798);
nor U5317 (N_5317,N_4694,N_4749);
nand U5318 (N_5318,N_4455,N_4590);
nor U5319 (N_5319,N_4133,N_3925);
and U5320 (N_5320,N_3747,N_3708);
or U5321 (N_5321,N_4157,N_4111);
xnor U5322 (N_5322,N_4131,N_4025);
and U5323 (N_5323,N_4515,N_3628);
and U5324 (N_5324,N_4750,N_4251);
or U5325 (N_5325,N_4403,N_3618);
nor U5326 (N_5326,N_4673,N_3803);
and U5327 (N_5327,N_3698,N_4778);
and U5328 (N_5328,N_4296,N_3630);
and U5329 (N_5329,N_4358,N_4733);
xnor U5330 (N_5330,N_3602,N_4316);
nand U5331 (N_5331,N_4660,N_3781);
and U5332 (N_5332,N_3912,N_4703);
nand U5333 (N_5333,N_3971,N_4191);
xnor U5334 (N_5334,N_3748,N_3669);
nor U5335 (N_5335,N_4278,N_4106);
and U5336 (N_5336,N_4736,N_4797);
xor U5337 (N_5337,N_4476,N_3823);
nand U5338 (N_5338,N_4319,N_3846);
nand U5339 (N_5339,N_4078,N_3622);
xnor U5340 (N_5340,N_4136,N_3832);
nand U5341 (N_5341,N_3816,N_4090);
xor U5342 (N_5342,N_4659,N_4638);
nor U5343 (N_5343,N_3647,N_4498);
nor U5344 (N_5344,N_3713,N_3635);
nand U5345 (N_5345,N_4180,N_4346);
xor U5346 (N_5346,N_4375,N_4627);
nor U5347 (N_5347,N_3935,N_4779);
and U5348 (N_5348,N_4238,N_4481);
or U5349 (N_5349,N_3788,N_4766);
and U5350 (N_5350,N_4148,N_3732);
and U5351 (N_5351,N_3760,N_3968);
nor U5352 (N_5352,N_4448,N_4635);
and U5353 (N_5353,N_3979,N_4539);
nor U5354 (N_5354,N_3928,N_4137);
xnor U5355 (N_5355,N_4360,N_4023);
nor U5356 (N_5356,N_4177,N_4574);
and U5357 (N_5357,N_4772,N_4771);
nand U5358 (N_5358,N_4221,N_3665);
xor U5359 (N_5359,N_4401,N_4002);
or U5360 (N_5360,N_3627,N_3690);
or U5361 (N_5361,N_4388,N_3826);
or U5362 (N_5362,N_3945,N_4129);
nand U5363 (N_5363,N_3815,N_3957);
nor U5364 (N_5364,N_4322,N_4431);
xnor U5365 (N_5365,N_4785,N_4596);
or U5366 (N_5366,N_3989,N_4292);
nor U5367 (N_5367,N_3706,N_4588);
or U5368 (N_5368,N_4088,N_3736);
xor U5369 (N_5369,N_3782,N_4389);
and U5370 (N_5370,N_4298,N_3986);
xor U5371 (N_5371,N_4592,N_4353);
nand U5372 (N_5372,N_4519,N_4165);
nor U5373 (N_5373,N_4022,N_4320);
or U5374 (N_5374,N_4072,N_4575);
xor U5375 (N_5375,N_4677,N_4692);
nand U5376 (N_5376,N_4721,N_4368);
or U5377 (N_5377,N_4776,N_4775);
nand U5378 (N_5378,N_4009,N_3860);
and U5379 (N_5379,N_4504,N_4224);
and U5380 (N_5380,N_4066,N_3909);
or U5381 (N_5381,N_3931,N_4104);
nor U5382 (N_5382,N_3610,N_4160);
nor U5383 (N_5383,N_4475,N_4051);
nor U5384 (N_5384,N_3605,N_4608);
nand U5385 (N_5385,N_4207,N_3700);
or U5386 (N_5386,N_4121,N_3811);
and U5387 (N_5387,N_4774,N_4055);
nor U5388 (N_5388,N_4628,N_3959);
nand U5389 (N_5389,N_4342,N_4744);
or U5390 (N_5390,N_3642,N_3944);
nor U5391 (N_5391,N_4042,N_3808);
or U5392 (N_5392,N_4291,N_4676);
nor U5393 (N_5393,N_4329,N_4364);
nand U5394 (N_5394,N_3981,N_4156);
nor U5395 (N_5395,N_3715,N_3819);
or U5396 (N_5396,N_3895,N_3785);
and U5397 (N_5397,N_4113,N_3641);
and U5398 (N_5398,N_3934,N_4039);
and U5399 (N_5399,N_4452,N_4697);
or U5400 (N_5400,N_4608,N_3993);
or U5401 (N_5401,N_4738,N_4311);
nor U5402 (N_5402,N_3805,N_3671);
xnor U5403 (N_5403,N_4793,N_4004);
nand U5404 (N_5404,N_4734,N_4033);
or U5405 (N_5405,N_4024,N_4776);
nor U5406 (N_5406,N_3913,N_3848);
or U5407 (N_5407,N_4636,N_3952);
nor U5408 (N_5408,N_4083,N_4724);
xor U5409 (N_5409,N_4614,N_4030);
xnor U5410 (N_5410,N_4480,N_4011);
xor U5411 (N_5411,N_4277,N_4018);
nand U5412 (N_5412,N_4061,N_4480);
nand U5413 (N_5413,N_4303,N_3625);
or U5414 (N_5414,N_4745,N_4523);
and U5415 (N_5415,N_3781,N_4515);
and U5416 (N_5416,N_4610,N_3632);
or U5417 (N_5417,N_4373,N_4097);
and U5418 (N_5418,N_3608,N_4282);
and U5419 (N_5419,N_4372,N_3816);
xnor U5420 (N_5420,N_3940,N_4040);
nand U5421 (N_5421,N_3782,N_4589);
nor U5422 (N_5422,N_4649,N_4521);
nand U5423 (N_5423,N_4113,N_4379);
nand U5424 (N_5424,N_3724,N_3649);
or U5425 (N_5425,N_4378,N_3847);
and U5426 (N_5426,N_4213,N_4219);
nand U5427 (N_5427,N_3819,N_4460);
nor U5428 (N_5428,N_4527,N_3853);
nand U5429 (N_5429,N_4346,N_3637);
or U5430 (N_5430,N_4395,N_4290);
or U5431 (N_5431,N_3623,N_3965);
or U5432 (N_5432,N_4049,N_4370);
xnor U5433 (N_5433,N_4569,N_4422);
and U5434 (N_5434,N_3827,N_4633);
and U5435 (N_5435,N_4284,N_4420);
nand U5436 (N_5436,N_3872,N_4110);
nor U5437 (N_5437,N_4006,N_4514);
or U5438 (N_5438,N_4554,N_3869);
nand U5439 (N_5439,N_3808,N_4675);
and U5440 (N_5440,N_3637,N_3951);
and U5441 (N_5441,N_4730,N_3670);
and U5442 (N_5442,N_4440,N_4378);
nand U5443 (N_5443,N_4526,N_3666);
nor U5444 (N_5444,N_4184,N_3799);
and U5445 (N_5445,N_4248,N_4071);
nand U5446 (N_5446,N_3672,N_3634);
and U5447 (N_5447,N_4065,N_4573);
or U5448 (N_5448,N_3730,N_4582);
and U5449 (N_5449,N_4480,N_4248);
nand U5450 (N_5450,N_3769,N_3984);
nand U5451 (N_5451,N_4612,N_4136);
nand U5452 (N_5452,N_3841,N_4077);
nor U5453 (N_5453,N_3740,N_4631);
xor U5454 (N_5454,N_4070,N_4064);
or U5455 (N_5455,N_4165,N_3935);
and U5456 (N_5456,N_4032,N_4591);
nor U5457 (N_5457,N_3866,N_4267);
and U5458 (N_5458,N_4345,N_3790);
nor U5459 (N_5459,N_3727,N_4136);
or U5460 (N_5460,N_4229,N_3671);
and U5461 (N_5461,N_3935,N_4555);
or U5462 (N_5462,N_4542,N_3634);
or U5463 (N_5463,N_4250,N_4625);
or U5464 (N_5464,N_4409,N_3658);
nor U5465 (N_5465,N_4709,N_4563);
nand U5466 (N_5466,N_3731,N_4185);
nand U5467 (N_5467,N_4747,N_4071);
xor U5468 (N_5468,N_4459,N_4435);
nor U5469 (N_5469,N_4317,N_4652);
nor U5470 (N_5470,N_4185,N_3891);
and U5471 (N_5471,N_4585,N_3969);
or U5472 (N_5472,N_4683,N_4765);
nand U5473 (N_5473,N_3823,N_4471);
and U5474 (N_5474,N_4131,N_3980);
nand U5475 (N_5475,N_4449,N_4137);
xnor U5476 (N_5476,N_4073,N_3839);
nand U5477 (N_5477,N_3628,N_3720);
nand U5478 (N_5478,N_4118,N_3718);
nor U5479 (N_5479,N_4115,N_3757);
nor U5480 (N_5480,N_4574,N_3974);
nor U5481 (N_5481,N_4667,N_4347);
or U5482 (N_5482,N_3708,N_3767);
and U5483 (N_5483,N_3990,N_3924);
xor U5484 (N_5484,N_4632,N_3858);
and U5485 (N_5485,N_4749,N_4011);
xnor U5486 (N_5486,N_4732,N_4027);
and U5487 (N_5487,N_4725,N_4330);
nor U5488 (N_5488,N_4524,N_4173);
or U5489 (N_5489,N_4530,N_4233);
nand U5490 (N_5490,N_4696,N_3981);
nand U5491 (N_5491,N_4149,N_4636);
nand U5492 (N_5492,N_3742,N_4276);
nand U5493 (N_5493,N_4193,N_4374);
nand U5494 (N_5494,N_3653,N_4235);
xor U5495 (N_5495,N_3926,N_3619);
nor U5496 (N_5496,N_4760,N_3659);
nor U5497 (N_5497,N_3965,N_4276);
and U5498 (N_5498,N_3938,N_4107);
and U5499 (N_5499,N_4447,N_3773);
and U5500 (N_5500,N_4454,N_3882);
or U5501 (N_5501,N_4348,N_4034);
nor U5502 (N_5502,N_4718,N_3963);
xor U5503 (N_5503,N_4289,N_4511);
or U5504 (N_5504,N_4519,N_3848);
xor U5505 (N_5505,N_4472,N_3661);
nand U5506 (N_5506,N_4253,N_4339);
nand U5507 (N_5507,N_4027,N_3783);
xnor U5508 (N_5508,N_4359,N_4227);
and U5509 (N_5509,N_4128,N_4575);
or U5510 (N_5510,N_3600,N_3774);
nand U5511 (N_5511,N_4624,N_3692);
xor U5512 (N_5512,N_4401,N_3860);
nor U5513 (N_5513,N_4037,N_4028);
or U5514 (N_5514,N_4345,N_3838);
and U5515 (N_5515,N_3736,N_4483);
xor U5516 (N_5516,N_3720,N_4124);
or U5517 (N_5517,N_4717,N_4263);
nand U5518 (N_5518,N_4170,N_4725);
or U5519 (N_5519,N_4741,N_3922);
and U5520 (N_5520,N_4105,N_3813);
nand U5521 (N_5521,N_4312,N_4069);
or U5522 (N_5522,N_3852,N_4189);
nor U5523 (N_5523,N_3989,N_4152);
xor U5524 (N_5524,N_4331,N_4256);
and U5525 (N_5525,N_3993,N_3866);
or U5526 (N_5526,N_3909,N_4792);
xnor U5527 (N_5527,N_4011,N_4075);
xnor U5528 (N_5528,N_4472,N_3726);
or U5529 (N_5529,N_4401,N_3996);
xor U5530 (N_5530,N_3837,N_3655);
or U5531 (N_5531,N_4039,N_3827);
and U5532 (N_5532,N_4557,N_3753);
or U5533 (N_5533,N_4367,N_4353);
nand U5534 (N_5534,N_3993,N_4503);
xor U5535 (N_5535,N_4385,N_4161);
nand U5536 (N_5536,N_4720,N_3678);
or U5537 (N_5537,N_4068,N_4398);
or U5538 (N_5538,N_3976,N_4656);
xor U5539 (N_5539,N_4193,N_4366);
or U5540 (N_5540,N_4207,N_4578);
xnor U5541 (N_5541,N_4300,N_4397);
or U5542 (N_5542,N_4307,N_4747);
nand U5543 (N_5543,N_3821,N_4624);
nand U5544 (N_5544,N_4748,N_4303);
nor U5545 (N_5545,N_4663,N_4376);
and U5546 (N_5546,N_3654,N_4368);
nand U5547 (N_5547,N_4755,N_3777);
xnor U5548 (N_5548,N_3921,N_3760);
nor U5549 (N_5549,N_4095,N_4664);
nor U5550 (N_5550,N_3806,N_4588);
and U5551 (N_5551,N_4109,N_4493);
and U5552 (N_5552,N_4733,N_4786);
and U5553 (N_5553,N_3751,N_3986);
xor U5554 (N_5554,N_4492,N_3806);
and U5555 (N_5555,N_4120,N_4757);
or U5556 (N_5556,N_4503,N_3826);
or U5557 (N_5557,N_4497,N_3913);
nor U5558 (N_5558,N_3977,N_3838);
nand U5559 (N_5559,N_4710,N_4517);
xor U5560 (N_5560,N_4662,N_3678);
and U5561 (N_5561,N_3648,N_3665);
nor U5562 (N_5562,N_3711,N_4667);
and U5563 (N_5563,N_4248,N_4106);
or U5564 (N_5564,N_4693,N_4523);
xnor U5565 (N_5565,N_3759,N_4262);
or U5566 (N_5566,N_3860,N_4509);
and U5567 (N_5567,N_4505,N_4704);
and U5568 (N_5568,N_4461,N_4579);
and U5569 (N_5569,N_4042,N_4056);
or U5570 (N_5570,N_3889,N_4688);
nand U5571 (N_5571,N_3655,N_4517);
xnor U5572 (N_5572,N_4596,N_4064);
or U5573 (N_5573,N_3739,N_3726);
and U5574 (N_5574,N_4078,N_4432);
or U5575 (N_5575,N_4444,N_4348);
nor U5576 (N_5576,N_4589,N_4570);
or U5577 (N_5577,N_4156,N_4085);
nor U5578 (N_5578,N_4202,N_4157);
or U5579 (N_5579,N_4205,N_4492);
and U5580 (N_5580,N_4434,N_3958);
nor U5581 (N_5581,N_3884,N_4213);
xnor U5582 (N_5582,N_4023,N_4190);
and U5583 (N_5583,N_4427,N_4611);
and U5584 (N_5584,N_4727,N_4018);
nor U5585 (N_5585,N_4348,N_4581);
and U5586 (N_5586,N_4312,N_4399);
nor U5587 (N_5587,N_3960,N_4330);
xnor U5588 (N_5588,N_3929,N_3612);
xor U5589 (N_5589,N_4294,N_4460);
nand U5590 (N_5590,N_4485,N_3809);
nor U5591 (N_5591,N_4130,N_4515);
nor U5592 (N_5592,N_3849,N_4487);
or U5593 (N_5593,N_3630,N_4212);
and U5594 (N_5594,N_4154,N_3941);
or U5595 (N_5595,N_3756,N_3945);
and U5596 (N_5596,N_3796,N_4731);
or U5597 (N_5597,N_4480,N_3757);
nor U5598 (N_5598,N_3760,N_3779);
xnor U5599 (N_5599,N_4540,N_4509);
xnor U5600 (N_5600,N_3906,N_3662);
and U5601 (N_5601,N_3796,N_3783);
xor U5602 (N_5602,N_4613,N_3748);
and U5603 (N_5603,N_4681,N_3643);
nor U5604 (N_5604,N_3670,N_4638);
nand U5605 (N_5605,N_4428,N_4746);
nor U5606 (N_5606,N_3826,N_4769);
or U5607 (N_5607,N_4354,N_4378);
nor U5608 (N_5608,N_4511,N_4768);
nand U5609 (N_5609,N_3717,N_4280);
nor U5610 (N_5610,N_4031,N_4092);
nor U5611 (N_5611,N_3997,N_3751);
and U5612 (N_5612,N_4231,N_3681);
or U5613 (N_5613,N_3744,N_4784);
xnor U5614 (N_5614,N_3783,N_3997);
or U5615 (N_5615,N_4097,N_3882);
and U5616 (N_5616,N_3627,N_4360);
or U5617 (N_5617,N_3737,N_4354);
xor U5618 (N_5618,N_3630,N_3964);
nand U5619 (N_5619,N_4458,N_4006);
and U5620 (N_5620,N_4708,N_4268);
and U5621 (N_5621,N_4766,N_3742);
nand U5622 (N_5622,N_3861,N_4152);
and U5623 (N_5623,N_3640,N_4776);
xnor U5624 (N_5624,N_4291,N_4635);
xnor U5625 (N_5625,N_4131,N_4214);
and U5626 (N_5626,N_3638,N_4066);
nand U5627 (N_5627,N_4090,N_3898);
xnor U5628 (N_5628,N_3784,N_4520);
and U5629 (N_5629,N_4178,N_3890);
and U5630 (N_5630,N_4202,N_3899);
or U5631 (N_5631,N_4014,N_3952);
or U5632 (N_5632,N_4544,N_3645);
or U5633 (N_5633,N_4794,N_4680);
or U5634 (N_5634,N_4363,N_4050);
or U5635 (N_5635,N_4262,N_4437);
or U5636 (N_5636,N_4535,N_4566);
and U5637 (N_5637,N_4481,N_4353);
nand U5638 (N_5638,N_4203,N_3658);
nor U5639 (N_5639,N_4015,N_4309);
nand U5640 (N_5640,N_3872,N_4636);
or U5641 (N_5641,N_4074,N_3774);
and U5642 (N_5642,N_4040,N_4376);
and U5643 (N_5643,N_4088,N_4688);
or U5644 (N_5644,N_3668,N_3896);
nor U5645 (N_5645,N_4096,N_3900);
nand U5646 (N_5646,N_3918,N_4633);
or U5647 (N_5647,N_4368,N_4793);
nand U5648 (N_5648,N_3602,N_3842);
xnor U5649 (N_5649,N_4700,N_3983);
or U5650 (N_5650,N_3725,N_4712);
xor U5651 (N_5651,N_4375,N_4321);
and U5652 (N_5652,N_4300,N_4579);
nor U5653 (N_5653,N_3936,N_3926);
or U5654 (N_5654,N_4229,N_4376);
nand U5655 (N_5655,N_3600,N_3700);
or U5656 (N_5656,N_4276,N_4065);
nor U5657 (N_5657,N_3929,N_3918);
nand U5658 (N_5658,N_3818,N_3751);
and U5659 (N_5659,N_4605,N_3940);
xor U5660 (N_5660,N_4119,N_3959);
or U5661 (N_5661,N_4095,N_4096);
nor U5662 (N_5662,N_3773,N_3996);
or U5663 (N_5663,N_4025,N_4333);
xor U5664 (N_5664,N_4543,N_3998);
nand U5665 (N_5665,N_3975,N_4242);
and U5666 (N_5666,N_4580,N_3602);
xnor U5667 (N_5667,N_4063,N_4280);
xor U5668 (N_5668,N_4455,N_4446);
or U5669 (N_5669,N_4150,N_3840);
and U5670 (N_5670,N_4252,N_3819);
xnor U5671 (N_5671,N_4550,N_3841);
nand U5672 (N_5672,N_3614,N_4285);
nor U5673 (N_5673,N_3831,N_4436);
or U5674 (N_5674,N_4527,N_3889);
or U5675 (N_5675,N_4141,N_4794);
xor U5676 (N_5676,N_4776,N_3959);
or U5677 (N_5677,N_4218,N_4723);
and U5678 (N_5678,N_4269,N_3643);
and U5679 (N_5679,N_4583,N_3665);
and U5680 (N_5680,N_4097,N_4167);
nor U5681 (N_5681,N_4103,N_4691);
nand U5682 (N_5682,N_3690,N_3955);
nor U5683 (N_5683,N_4111,N_4170);
and U5684 (N_5684,N_3748,N_4266);
and U5685 (N_5685,N_3697,N_3998);
or U5686 (N_5686,N_3931,N_4593);
nand U5687 (N_5687,N_3699,N_4121);
and U5688 (N_5688,N_4429,N_4315);
or U5689 (N_5689,N_4387,N_4684);
and U5690 (N_5690,N_4422,N_4652);
nand U5691 (N_5691,N_3696,N_4565);
or U5692 (N_5692,N_4263,N_3831);
nand U5693 (N_5693,N_4300,N_4311);
nor U5694 (N_5694,N_3642,N_3887);
xnor U5695 (N_5695,N_3856,N_3751);
nor U5696 (N_5696,N_4198,N_4727);
or U5697 (N_5697,N_4113,N_4756);
and U5698 (N_5698,N_3612,N_3828);
or U5699 (N_5699,N_3875,N_4014);
nand U5700 (N_5700,N_3886,N_3701);
nor U5701 (N_5701,N_4443,N_3917);
xor U5702 (N_5702,N_3604,N_3949);
and U5703 (N_5703,N_4769,N_4648);
nor U5704 (N_5704,N_3853,N_4696);
or U5705 (N_5705,N_4454,N_3985);
and U5706 (N_5706,N_4053,N_4132);
nand U5707 (N_5707,N_4226,N_4459);
nor U5708 (N_5708,N_4507,N_4509);
xnor U5709 (N_5709,N_4466,N_3665);
nor U5710 (N_5710,N_4414,N_3813);
xor U5711 (N_5711,N_4353,N_4344);
xnor U5712 (N_5712,N_4536,N_4377);
and U5713 (N_5713,N_3852,N_3700);
nor U5714 (N_5714,N_3604,N_4687);
or U5715 (N_5715,N_3916,N_3928);
and U5716 (N_5716,N_4141,N_3708);
and U5717 (N_5717,N_4276,N_3911);
nand U5718 (N_5718,N_4153,N_3620);
nor U5719 (N_5719,N_4707,N_4189);
nor U5720 (N_5720,N_3665,N_4640);
xnor U5721 (N_5721,N_3695,N_4749);
xnor U5722 (N_5722,N_4736,N_3835);
or U5723 (N_5723,N_4648,N_4414);
nand U5724 (N_5724,N_4358,N_3916);
xor U5725 (N_5725,N_3791,N_4531);
nor U5726 (N_5726,N_3743,N_4616);
nor U5727 (N_5727,N_4689,N_3773);
and U5728 (N_5728,N_3756,N_4557);
nor U5729 (N_5729,N_4279,N_3623);
or U5730 (N_5730,N_3694,N_4087);
and U5731 (N_5731,N_3900,N_3930);
or U5732 (N_5732,N_3601,N_4449);
nor U5733 (N_5733,N_3963,N_4085);
or U5734 (N_5734,N_4381,N_4626);
nor U5735 (N_5735,N_4100,N_4667);
or U5736 (N_5736,N_4260,N_4031);
or U5737 (N_5737,N_4766,N_3854);
or U5738 (N_5738,N_4204,N_4656);
nand U5739 (N_5739,N_4463,N_4393);
nor U5740 (N_5740,N_4330,N_4048);
and U5741 (N_5741,N_3757,N_4741);
xor U5742 (N_5742,N_4573,N_4436);
nor U5743 (N_5743,N_4689,N_4539);
xnor U5744 (N_5744,N_4673,N_4312);
xor U5745 (N_5745,N_4542,N_4061);
nand U5746 (N_5746,N_3771,N_4119);
nor U5747 (N_5747,N_4333,N_4176);
or U5748 (N_5748,N_4021,N_3636);
nand U5749 (N_5749,N_4072,N_4786);
or U5750 (N_5750,N_4411,N_4634);
nor U5751 (N_5751,N_4487,N_4275);
nand U5752 (N_5752,N_3852,N_4109);
xor U5753 (N_5753,N_4234,N_3915);
or U5754 (N_5754,N_4595,N_4010);
or U5755 (N_5755,N_4623,N_4049);
and U5756 (N_5756,N_4448,N_3979);
nor U5757 (N_5757,N_3959,N_3801);
and U5758 (N_5758,N_4129,N_4080);
nor U5759 (N_5759,N_4342,N_4110);
or U5760 (N_5760,N_4205,N_3733);
xor U5761 (N_5761,N_4202,N_3883);
and U5762 (N_5762,N_4161,N_4792);
and U5763 (N_5763,N_3909,N_4429);
xor U5764 (N_5764,N_3874,N_4557);
nor U5765 (N_5765,N_4198,N_3760);
and U5766 (N_5766,N_3738,N_4624);
and U5767 (N_5767,N_3833,N_4177);
and U5768 (N_5768,N_4200,N_4752);
nor U5769 (N_5769,N_3611,N_3981);
nand U5770 (N_5770,N_3888,N_3614);
xnor U5771 (N_5771,N_4028,N_4791);
or U5772 (N_5772,N_4553,N_4171);
xor U5773 (N_5773,N_4683,N_3896);
or U5774 (N_5774,N_4664,N_4572);
nand U5775 (N_5775,N_4633,N_3758);
nor U5776 (N_5776,N_3715,N_4698);
xnor U5777 (N_5777,N_4707,N_4513);
nor U5778 (N_5778,N_4165,N_3768);
or U5779 (N_5779,N_4774,N_4192);
xor U5780 (N_5780,N_4460,N_3663);
and U5781 (N_5781,N_4267,N_3721);
xnor U5782 (N_5782,N_4550,N_4622);
nand U5783 (N_5783,N_4574,N_4214);
and U5784 (N_5784,N_4762,N_4697);
or U5785 (N_5785,N_3851,N_4128);
and U5786 (N_5786,N_4663,N_4714);
nor U5787 (N_5787,N_4277,N_4263);
nor U5788 (N_5788,N_4488,N_4705);
or U5789 (N_5789,N_3830,N_3688);
nor U5790 (N_5790,N_3870,N_4236);
and U5791 (N_5791,N_3729,N_4175);
xnor U5792 (N_5792,N_4477,N_3891);
nand U5793 (N_5793,N_3938,N_3855);
nor U5794 (N_5794,N_3976,N_4346);
nand U5795 (N_5795,N_3687,N_3865);
and U5796 (N_5796,N_4081,N_4436);
nand U5797 (N_5797,N_4500,N_4166);
and U5798 (N_5798,N_4656,N_4052);
nand U5799 (N_5799,N_3995,N_4626);
xor U5800 (N_5800,N_4576,N_4144);
and U5801 (N_5801,N_3744,N_4238);
nor U5802 (N_5802,N_3920,N_4372);
nor U5803 (N_5803,N_4750,N_3939);
and U5804 (N_5804,N_4517,N_4405);
nand U5805 (N_5805,N_4547,N_4137);
nand U5806 (N_5806,N_4511,N_4233);
and U5807 (N_5807,N_4604,N_4629);
or U5808 (N_5808,N_3713,N_4514);
nand U5809 (N_5809,N_3605,N_4414);
and U5810 (N_5810,N_4713,N_3633);
nand U5811 (N_5811,N_4145,N_4737);
nand U5812 (N_5812,N_3697,N_3619);
xor U5813 (N_5813,N_3991,N_3844);
nand U5814 (N_5814,N_4671,N_4562);
nor U5815 (N_5815,N_3741,N_4191);
and U5816 (N_5816,N_4669,N_4403);
nor U5817 (N_5817,N_4796,N_3705);
or U5818 (N_5818,N_4632,N_3948);
and U5819 (N_5819,N_4610,N_4404);
xnor U5820 (N_5820,N_4207,N_4624);
nand U5821 (N_5821,N_4035,N_4149);
xor U5822 (N_5822,N_3766,N_3673);
or U5823 (N_5823,N_3813,N_4766);
nand U5824 (N_5824,N_4105,N_4758);
nand U5825 (N_5825,N_3865,N_3689);
nand U5826 (N_5826,N_3610,N_3656);
nor U5827 (N_5827,N_4196,N_3605);
nor U5828 (N_5828,N_4377,N_3744);
or U5829 (N_5829,N_4273,N_4294);
and U5830 (N_5830,N_4598,N_4647);
or U5831 (N_5831,N_4455,N_4690);
nand U5832 (N_5832,N_3692,N_3668);
xor U5833 (N_5833,N_3692,N_3707);
nand U5834 (N_5834,N_4680,N_3616);
and U5835 (N_5835,N_4103,N_4479);
and U5836 (N_5836,N_4299,N_4723);
xor U5837 (N_5837,N_3911,N_4572);
and U5838 (N_5838,N_3731,N_4239);
xor U5839 (N_5839,N_4078,N_4283);
nand U5840 (N_5840,N_4470,N_3662);
or U5841 (N_5841,N_4210,N_3975);
nand U5842 (N_5842,N_4385,N_4081);
nor U5843 (N_5843,N_3817,N_4126);
and U5844 (N_5844,N_3971,N_4130);
or U5845 (N_5845,N_3630,N_3707);
xnor U5846 (N_5846,N_4435,N_4403);
nand U5847 (N_5847,N_4571,N_4531);
xor U5848 (N_5848,N_3881,N_4615);
nand U5849 (N_5849,N_4226,N_4671);
or U5850 (N_5850,N_4620,N_4616);
or U5851 (N_5851,N_4184,N_4510);
xor U5852 (N_5852,N_4131,N_4549);
nand U5853 (N_5853,N_4180,N_4077);
or U5854 (N_5854,N_4343,N_3752);
and U5855 (N_5855,N_3810,N_4718);
and U5856 (N_5856,N_4352,N_3884);
xor U5857 (N_5857,N_3627,N_4301);
nand U5858 (N_5858,N_4737,N_4024);
xnor U5859 (N_5859,N_4545,N_4109);
nor U5860 (N_5860,N_4572,N_4713);
xnor U5861 (N_5861,N_4668,N_4640);
nor U5862 (N_5862,N_4412,N_4415);
and U5863 (N_5863,N_4605,N_4375);
or U5864 (N_5864,N_3713,N_4281);
nor U5865 (N_5865,N_4678,N_4268);
or U5866 (N_5866,N_4645,N_3807);
or U5867 (N_5867,N_4311,N_3734);
nand U5868 (N_5868,N_4787,N_4040);
or U5869 (N_5869,N_4406,N_3927);
and U5870 (N_5870,N_4362,N_4724);
nor U5871 (N_5871,N_4242,N_3732);
and U5872 (N_5872,N_4131,N_4014);
nand U5873 (N_5873,N_4233,N_4411);
or U5874 (N_5874,N_4292,N_4230);
or U5875 (N_5875,N_4227,N_4303);
nor U5876 (N_5876,N_3686,N_4077);
nor U5877 (N_5877,N_4604,N_3662);
nand U5878 (N_5878,N_4150,N_4003);
nor U5879 (N_5879,N_3601,N_4380);
or U5880 (N_5880,N_3823,N_4090);
or U5881 (N_5881,N_4744,N_4180);
or U5882 (N_5882,N_4608,N_4161);
nor U5883 (N_5883,N_4374,N_4340);
nor U5884 (N_5884,N_4497,N_4194);
or U5885 (N_5885,N_3881,N_4465);
nor U5886 (N_5886,N_3636,N_4709);
or U5887 (N_5887,N_4576,N_3817);
or U5888 (N_5888,N_4193,N_3868);
nand U5889 (N_5889,N_3943,N_4354);
and U5890 (N_5890,N_4675,N_4149);
nor U5891 (N_5891,N_4348,N_4380);
xnor U5892 (N_5892,N_3937,N_3882);
or U5893 (N_5893,N_4491,N_4279);
xnor U5894 (N_5894,N_4247,N_4002);
nand U5895 (N_5895,N_4512,N_4470);
and U5896 (N_5896,N_4392,N_4298);
or U5897 (N_5897,N_3747,N_3911);
nand U5898 (N_5898,N_3941,N_4043);
and U5899 (N_5899,N_3715,N_4649);
and U5900 (N_5900,N_4784,N_3937);
nand U5901 (N_5901,N_4221,N_4769);
and U5902 (N_5902,N_3697,N_4655);
and U5903 (N_5903,N_3889,N_4126);
or U5904 (N_5904,N_3933,N_3966);
or U5905 (N_5905,N_4187,N_4610);
nand U5906 (N_5906,N_3740,N_3743);
and U5907 (N_5907,N_4021,N_3621);
nor U5908 (N_5908,N_3785,N_4169);
nor U5909 (N_5909,N_4350,N_4051);
or U5910 (N_5910,N_3662,N_4399);
and U5911 (N_5911,N_4486,N_4246);
or U5912 (N_5912,N_3605,N_4682);
nor U5913 (N_5913,N_4542,N_4695);
xnor U5914 (N_5914,N_4269,N_3928);
and U5915 (N_5915,N_4397,N_3931);
nor U5916 (N_5916,N_4041,N_3752);
and U5917 (N_5917,N_4283,N_4150);
and U5918 (N_5918,N_4705,N_4137);
and U5919 (N_5919,N_4094,N_3623);
nor U5920 (N_5920,N_4178,N_3988);
nand U5921 (N_5921,N_4656,N_3715);
or U5922 (N_5922,N_4300,N_3649);
nor U5923 (N_5923,N_4023,N_3693);
or U5924 (N_5924,N_3865,N_4747);
or U5925 (N_5925,N_4609,N_3960);
nand U5926 (N_5926,N_4651,N_3777);
and U5927 (N_5927,N_4440,N_4223);
nand U5928 (N_5928,N_4264,N_3779);
and U5929 (N_5929,N_4435,N_4600);
and U5930 (N_5930,N_4194,N_4098);
nand U5931 (N_5931,N_4275,N_4261);
nand U5932 (N_5932,N_4282,N_3900);
nand U5933 (N_5933,N_4199,N_3670);
nor U5934 (N_5934,N_4058,N_3881);
and U5935 (N_5935,N_4034,N_3803);
or U5936 (N_5936,N_4736,N_3977);
and U5937 (N_5937,N_4407,N_4072);
or U5938 (N_5938,N_4592,N_3761);
nor U5939 (N_5939,N_4653,N_4764);
xor U5940 (N_5940,N_4061,N_4341);
and U5941 (N_5941,N_3632,N_4664);
nor U5942 (N_5942,N_4592,N_4065);
nor U5943 (N_5943,N_4605,N_4383);
nor U5944 (N_5944,N_4072,N_3791);
nand U5945 (N_5945,N_4395,N_3998);
or U5946 (N_5946,N_4786,N_4503);
and U5947 (N_5947,N_3828,N_4065);
xor U5948 (N_5948,N_4179,N_4273);
and U5949 (N_5949,N_3820,N_3713);
nor U5950 (N_5950,N_3813,N_3975);
and U5951 (N_5951,N_3911,N_4516);
nand U5952 (N_5952,N_3635,N_3732);
nor U5953 (N_5953,N_4353,N_4735);
nand U5954 (N_5954,N_4374,N_3944);
nor U5955 (N_5955,N_4075,N_3855);
and U5956 (N_5956,N_4416,N_4110);
xor U5957 (N_5957,N_4796,N_4580);
xor U5958 (N_5958,N_3950,N_4491);
nand U5959 (N_5959,N_3672,N_4324);
and U5960 (N_5960,N_4266,N_4727);
xor U5961 (N_5961,N_4384,N_4533);
and U5962 (N_5962,N_4495,N_4472);
and U5963 (N_5963,N_4213,N_4132);
nor U5964 (N_5964,N_3862,N_4527);
or U5965 (N_5965,N_3687,N_3685);
and U5966 (N_5966,N_4695,N_4020);
and U5967 (N_5967,N_3782,N_4769);
nor U5968 (N_5968,N_4399,N_4300);
or U5969 (N_5969,N_4265,N_4137);
xor U5970 (N_5970,N_4403,N_3654);
nor U5971 (N_5971,N_4275,N_4796);
xor U5972 (N_5972,N_3875,N_4180);
nor U5973 (N_5973,N_4702,N_4357);
xnor U5974 (N_5974,N_4170,N_4464);
nor U5975 (N_5975,N_3932,N_4629);
or U5976 (N_5976,N_4336,N_3810);
nor U5977 (N_5977,N_4591,N_4415);
nand U5978 (N_5978,N_4221,N_4577);
and U5979 (N_5979,N_4401,N_4561);
nor U5980 (N_5980,N_4687,N_3754);
nor U5981 (N_5981,N_3674,N_4247);
nand U5982 (N_5982,N_4252,N_3600);
nor U5983 (N_5983,N_4508,N_3960);
nor U5984 (N_5984,N_3758,N_3723);
and U5985 (N_5985,N_3660,N_3692);
and U5986 (N_5986,N_3983,N_4452);
or U5987 (N_5987,N_3921,N_4057);
xnor U5988 (N_5988,N_4358,N_3957);
and U5989 (N_5989,N_3637,N_4382);
nor U5990 (N_5990,N_4157,N_3703);
nor U5991 (N_5991,N_4200,N_3807);
nor U5992 (N_5992,N_3727,N_4397);
nor U5993 (N_5993,N_4744,N_4258);
nand U5994 (N_5994,N_3960,N_4626);
nor U5995 (N_5995,N_3931,N_3644);
or U5996 (N_5996,N_3815,N_4788);
nor U5997 (N_5997,N_3780,N_3812);
or U5998 (N_5998,N_4202,N_4297);
nor U5999 (N_5999,N_3719,N_4508);
nor U6000 (N_6000,N_5330,N_5967);
nor U6001 (N_6001,N_5001,N_4963);
nand U6002 (N_6002,N_5360,N_5431);
nand U6003 (N_6003,N_5249,N_5643);
or U6004 (N_6004,N_5925,N_5931);
nand U6005 (N_6005,N_5719,N_5484);
or U6006 (N_6006,N_5839,N_5971);
and U6007 (N_6007,N_4807,N_5645);
xnor U6008 (N_6008,N_5371,N_5050);
and U6009 (N_6009,N_5485,N_5392);
and U6010 (N_6010,N_5955,N_5912);
xor U6011 (N_6011,N_5059,N_5474);
nor U6012 (N_6012,N_5534,N_5283);
or U6013 (N_6013,N_5038,N_4856);
xor U6014 (N_6014,N_5374,N_5417);
or U6015 (N_6015,N_4932,N_5304);
xor U6016 (N_6016,N_4927,N_5650);
nor U6017 (N_6017,N_4829,N_5275);
nand U6018 (N_6018,N_5870,N_5129);
nor U6019 (N_6019,N_5286,N_5903);
xor U6020 (N_6020,N_5082,N_5506);
nand U6021 (N_6021,N_4813,N_5936);
nor U6022 (N_6022,N_5575,N_5873);
and U6023 (N_6023,N_5943,N_4959);
and U6024 (N_6024,N_5667,N_5227);
nor U6025 (N_6025,N_5364,N_4987);
nor U6026 (N_6026,N_5580,N_5174);
nor U6027 (N_6027,N_5015,N_5974);
nand U6028 (N_6028,N_5616,N_5133);
xnor U6029 (N_6029,N_5526,N_5994);
or U6030 (N_6030,N_5715,N_5421);
nand U6031 (N_6031,N_5297,N_5295);
and U6032 (N_6032,N_4960,N_4931);
or U6033 (N_6033,N_5085,N_5377);
and U6034 (N_6034,N_5866,N_5261);
or U6035 (N_6035,N_5656,N_5576);
nand U6036 (N_6036,N_5830,N_5333);
or U6037 (N_6037,N_5531,N_5503);
nand U6038 (N_6038,N_5411,N_5378);
and U6039 (N_6039,N_5871,N_5395);
or U6040 (N_6040,N_5666,N_5182);
or U6041 (N_6041,N_5770,N_5438);
nor U6042 (N_6042,N_5516,N_5710);
nand U6043 (N_6043,N_5141,N_5555);
nand U6044 (N_6044,N_5403,N_5525);
or U6045 (N_6045,N_5062,N_5434);
or U6046 (N_6046,N_5495,N_5224);
and U6047 (N_6047,N_5649,N_5184);
and U6048 (N_6048,N_5614,N_5535);
or U6049 (N_6049,N_5709,N_5189);
nor U6050 (N_6050,N_5891,N_5829);
or U6051 (N_6051,N_5468,N_5408);
nor U6052 (N_6052,N_4886,N_5047);
and U6053 (N_6053,N_5391,N_5442);
nand U6054 (N_6054,N_5569,N_5454);
nand U6055 (N_6055,N_5665,N_5479);
xnor U6056 (N_6056,N_5195,N_4824);
or U6057 (N_6057,N_5450,N_5633);
or U6058 (N_6058,N_5109,N_5087);
or U6059 (N_6059,N_5472,N_5733);
nand U6060 (N_6060,N_5996,N_4879);
nand U6061 (N_6061,N_5811,N_5150);
nand U6062 (N_6062,N_5852,N_5845);
nor U6063 (N_6063,N_5008,N_5499);
xnor U6064 (N_6064,N_5429,N_5396);
or U6065 (N_6065,N_5678,N_5383);
or U6066 (N_6066,N_5324,N_5142);
nand U6067 (N_6067,N_5316,N_5804);
and U6068 (N_6068,N_4921,N_5066);
and U6069 (N_6069,N_5581,N_5124);
or U6070 (N_6070,N_5307,N_5613);
xor U6071 (N_6071,N_5584,N_4998);
nor U6072 (N_6072,N_5798,N_5278);
nand U6073 (N_6073,N_5457,N_5545);
or U6074 (N_6074,N_5191,N_4945);
and U6075 (N_6075,N_5117,N_5522);
or U6076 (N_6076,N_5636,N_5158);
or U6077 (N_6077,N_5552,N_4869);
nand U6078 (N_6078,N_5606,N_5905);
nor U6079 (N_6079,N_5564,N_5361);
xor U6080 (N_6080,N_5147,N_5266);
xnor U6081 (N_6081,N_5847,N_5817);
nor U6082 (N_6082,N_5946,N_5076);
xor U6083 (N_6083,N_5044,N_5625);
nor U6084 (N_6084,N_5097,N_4968);
and U6085 (N_6085,N_5470,N_4833);
xnor U6086 (N_6086,N_5646,N_5493);
or U6087 (N_6087,N_5435,N_5951);
nand U6088 (N_6088,N_5730,N_5110);
xnor U6089 (N_6089,N_5599,N_5718);
nand U6090 (N_6090,N_5296,N_4967);
and U6091 (N_6091,N_5598,N_4804);
and U6092 (N_6092,N_5683,N_5366);
or U6093 (N_6093,N_5538,N_5441);
and U6094 (N_6094,N_4889,N_5746);
nor U6095 (N_6095,N_5353,N_5220);
and U6096 (N_6096,N_5600,N_5234);
and U6097 (N_6097,N_4914,N_5370);
nand U6098 (N_6098,N_5022,N_5563);
nand U6099 (N_6099,N_5623,N_5807);
nor U6100 (N_6100,N_5983,N_5835);
nand U6101 (N_6101,N_5618,N_5032);
xnor U6102 (N_6102,N_5963,N_5306);
and U6103 (N_6103,N_4903,N_5959);
nor U6104 (N_6104,N_5867,N_5458);
or U6105 (N_6105,N_5016,N_5610);
xor U6106 (N_6106,N_5664,N_5820);
nor U6107 (N_6107,N_5791,N_5273);
and U6108 (N_6108,N_5123,N_4993);
and U6109 (N_6109,N_5387,N_5877);
nand U6110 (N_6110,N_4839,N_5750);
nor U6111 (N_6111,N_5165,N_5476);
nand U6112 (N_6112,N_5897,N_5321);
nor U6113 (N_6113,N_5216,N_5009);
nand U6114 (N_6114,N_5005,N_5202);
nor U6115 (N_6115,N_4940,N_5337);
nor U6116 (N_6116,N_5887,N_5898);
and U6117 (N_6117,N_5146,N_5237);
and U6118 (N_6118,N_4958,N_5907);
or U6119 (N_6119,N_4939,N_5162);
xnor U6120 (N_6120,N_5761,N_4801);
and U6121 (N_6121,N_5632,N_5096);
and U6122 (N_6122,N_5194,N_4877);
or U6123 (N_6123,N_5230,N_5685);
and U6124 (N_6124,N_5111,N_5156);
nor U6125 (N_6125,N_5063,N_5399);
and U6126 (N_6126,N_4814,N_5676);
nor U6127 (N_6127,N_5390,N_5389);
and U6128 (N_6128,N_5995,N_5626);
nor U6129 (N_6129,N_4876,N_4866);
or U6130 (N_6130,N_5303,N_5058);
or U6131 (N_6131,N_5402,N_5318);
or U6132 (N_6132,N_5701,N_5192);
xnor U6133 (N_6133,N_5644,N_5968);
nand U6134 (N_6134,N_5838,N_5433);
xor U6135 (N_6135,N_5322,N_5265);
xor U6136 (N_6136,N_4859,N_4842);
nand U6137 (N_6137,N_5103,N_5257);
or U6138 (N_6138,N_5507,N_4844);
nor U6139 (N_6139,N_5821,N_5615);
or U6140 (N_6140,N_5823,N_4946);
and U6141 (N_6141,N_5100,N_5185);
nor U6142 (N_6142,N_4821,N_5879);
or U6143 (N_6143,N_5253,N_4865);
xor U6144 (N_6144,N_5874,N_5197);
nor U6145 (N_6145,N_5833,N_5126);
nor U6146 (N_6146,N_5211,N_5588);
and U6147 (N_6147,N_5724,N_5386);
and U6148 (N_6148,N_5177,N_5603);
xor U6149 (N_6149,N_5091,N_5589);
nor U6150 (N_6150,N_5621,N_5459);
nor U6151 (N_6151,N_5717,N_4902);
nor U6152 (N_6152,N_5842,N_5412);
xor U6153 (N_6153,N_5952,N_5148);
nor U6154 (N_6154,N_5751,N_5945);
nor U6155 (N_6155,N_5565,N_4944);
nor U6156 (N_6156,N_5671,N_5138);
or U6157 (N_6157,N_4990,N_5323);
or U6158 (N_6158,N_5487,N_5913);
xor U6159 (N_6159,N_5732,N_4898);
nor U6160 (N_6160,N_5699,N_4911);
or U6161 (N_6161,N_5794,N_4868);
or U6162 (N_6162,N_5011,N_5345);
xor U6163 (N_6163,N_5662,N_5289);
and U6164 (N_6164,N_5652,N_5551);
nand U6165 (N_6165,N_5934,N_5927);
and U6166 (N_6166,N_5209,N_4918);
xnor U6167 (N_6167,N_5759,N_5728);
or U6168 (N_6168,N_5357,N_4906);
nand U6169 (N_6169,N_5369,N_5035);
and U6170 (N_6170,N_5653,N_4895);
or U6171 (N_6171,N_5672,N_5801);
nor U6172 (N_6172,N_4892,N_4888);
nor U6173 (N_6173,N_5775,N_5233);
nand U6174 (N_6174,N_5579,N_4905);
nor U6175 (N_6175,N_5236,N_5583);
and U6176 (N_6176,N_4942,N_4857);
nand U6177 (N_6177,N_5027,N_5574);
nand U6178 (N_6178,N_5785,N_5068);
nand U6179 (N_6179,N_5269,N_5799);
nor U6180 (N_6180,N_5372,N_5542);
and U6181 (N_6181,N_5453,N_5228);
nand U6182 (N_6182,N_5836,N_5128);
nor U6183 (N_6183,N_5113,N_4860);
nand U6184 (N_6184,N_5570,N_5300);
xnor U6185 (N_6185,N_5053,N_4830);
nor U6186 (N_6186,N_5692,N_5642);
and U6187 (N_6187,N_4896,N_5171);
or U6188 (N_6188,N_5786,N_5231);
nand U6189 (N_6189,N_5602,N_4951);
and U6190 (N_6190,N_5325,N_4828);
or U6191 (N_6191,N_5203,N_4806);
and U6192 (N_6192,N_5781,N_5562);
xnor U6193 (N_6193,N_4955,N_4885);
and U6194 (N_6194,N_5972,N_5918);
xor U6195 (N_6195,N_5827,N_5302);
nor U6196 (N_6196,N_5074,N_4961);
nand U6197 (N_6197,N_5605,N_5463);
xnor U6198 (N_6198,N_5966,N_5594);
and U6199 (N_6199,N_4893,N_4949);
and U6200 (N_6200,N_5198,N_5217);
xor U6201 (N_6201,N_5512,N_4938);
and U6202 (N_6202,N_5766,N_5172);
and U6203 (N_6203,N_5819,N_5706);
xnor U6204 (N_6204,N_5334,N_5979);
nand U6205 (N_6205,N_5695,N_5893);
and U6206 (N_6206,N_5624,N_5002);
xnor U6207 (N_6207,N_5416,N_5862);
xor U6208 (N_6208,N_5726,N_5098);
nand U6209 (N_6209,N_5549,N_5406);
nand U6210 (N_6210,N_5868,N_4816);
or U6211 (N_6211,N_5277,N_5122);
and U6212 (N_6212,N_5883,N_4933);
nand U6213 (N_6213,N_5587,N_5067);
nor U6214 (N_6214,N_5341,N_5327);
xnor U6215 (N_6215,N_5631,N_5250);
or U6216 (N_6216,N_5081,N_5939);
or U6217 (N_6217,N_5385,N_5492);
nand U6218 (N_6218,N_4870,N_4965);
xnor U6219 (N_6219,N_5505,N_5166);
nand U6220 (N_6220,N_5439,N_5990);
and U6221 (N_6221,N_5550,N_5753);
and U6222 (N_6222,N_5875,N_4924);
and U6223 (N_6223,N_5338,N_5183);
xor U6224 (N_6224,N_5380,N_5376);
and U6225 (N_6225,N_5343,N_5677);
or U6226 (N_6226,N_5208,N_4917);
and U6227 (N_6227,N_4904,N_5301);
and U6228 (N_6228,N_5013,N_5886);
xnor U6229 (N_6229,N_5765,N_4972);
and U6230 (N_6230,N_5329,N_5478);
or U6231 (N_6231,N_5368,N_5070);
xor U6232 (N_6232,N_5577,N_5509);
and U6233 (N_6233,N_5263,N_5533);
nand U6234 (N_6234,N_5640,N_4997);
nor U6235 (N_6235,N_5657,N_5239);
nand U6236 (N_6236,N_5116,N_5312);
xnor U6237 (N_6237,N_5193,N_5687);
or U6238 (N_6238,N_5375,N_5860);
nor U6239 (N_6239,N_5524,N_5762);
and U6240 (N_6240,N_5517,N_5498);
and U6241 (N_6241,N_5373,N_5051);
nand U6242 (N_6242,N_5539,N_4884);
xnor U6243 (N_6243,N_5152,N_5536);
nand U6244 (N_6244,N_5452,N_5620);
nor U6245 (N_6245,N_5681,N_5557);
or U6246 (N_6246,N_4920,N_5086);
xor U6247 (N_6247,N_5986,N_5426);
or U6248 (N_6248,N_4846,N_5460);
nor U6249 (N_6249,N_5134,N_5713);
xnor U6250 (N_6250,N_5262,N_5161);
or U6251 (N_6251,N_5264,N_4831);
xor U6252 (N_6252,N_4956,N_5026);
and U6253 (N_6253,N_5168,N_5246);
nand U6254 (N_6254,N_4922,N_5639);
and U6255 (N_6255,N_5792,N_4957);
nand U6256 (N_6256,N_5741,N_5558);
xor U6257 (N_6257,N_5850,N_5359);
or U6258 (N_6258,N_4980,N_5175);
and U6259 (N_6259,N_5711,N_4851);
and U6260 (N_6260,N_4926,N_5083);
nor U6261 (N_6261,N_5365,N_5332);
xor U6262 (N_6262,N_5410,N_5419);
nand U6263 (N_6263,N_5440,N_5229);
and U6264 (N_6264,N_5409,N_4887);
xor U6265 (N_6265,N_5725,N_5714);
or U6266 (N_6266,N_4936,N_5832);
xnor U6267 (N_6267,N_5397,N_5856);
or U6268 (N_6268,N_5684,N_5401);
and U6269 (N_6269,N_5773,N_5101);
and U6270 (N_6270,N_4981,N_5328);
xor U6271 (N_6271,N_5004,N_5000);
or U6272 (N_6272,N_5553,N_5095);
xnor U6273 (N_6273,N_5747,N_5212);
nand U6274 (N_6274,N_4991,N_4923);
or U6275 (N_6275,N_5287,N_5331);
xor U6276 (N_6276,N_5556,N_5935);
or U6277 (N_6277,N_5696,N_5037);
xor U6278 (N_6278,N_5367,N_4954);
or U6279 (N_6279,N_4881,N_5446);
nor U6280 (N_6280,N_5888,N_5793);
nor U6281 (N_6281,N_5448,N_5055);
and U6282 (N_6282,N_5305,N_5119);
and U6283 (N_6283,N_5260,N_5423);
xor U6284 (N_6284,N_5885,N_5661);
xnor U6285 (N_6285,N_4871,N_4947);
and U6286 (N_6286,N_5077,N_5617);
and U6287 (N_6287,N_5754,N_4935);
nor U6288 (N_6288,N_5222,N_5447);
or U6289 (N_6289,N_5899,N_4973);
nor U6290 (N_6290,N_5069,N_5023);
and U6291 (N_6291,N_5863,N_5609);
or U6292 (N_6292,N_5796,N_5218);
nor U6293 (N_6293,N_5181,N_5675);
and U6294 (N_6294,N_5690,N_5572);
xnor U6295 (N_6295,N_5497,N_5244);
nand U6296 (N_6296,N_4894,N_5207);
nand U6297 (N_6297,N_5144,N_5957);
or U6298 (N_6298,N_4818,N_5169);
nor U6299 (N_6299,N_5561,N_5149);
and U6300 (N_6300,N_5480,N_5482);
xor U6301 (N_6301,N_5634,N_5991);
nor U6302 (N_6302,N_5586,N_5036);
nor U6303 (N_6303,N_5854,N_5483);
or U6304 (N_6304,N_5978,N_4934);
nor U6305 (N_6305,N_5929,N_4897);
nand U6306 (N_6306,N_5090,N_5720);
xor U6307 (N_6307,N_5407,N_4836);
nor U6308 (N_6308,N_5029,N_4812);
and U6309 (N_6309,N_5948,N_5544);
nand U6310 (N_6310,N_5201,N_5777);
nand U6311 (N_6311,N_4811,N_5938);
or U6312 (N_6312,N_5226,N_5464);
and U6313 (N_6313,N_5909,N_5735);
nor U6314 (N_6314,N_5099,N_5188);
and U6315 (N_6315,N_5471,N_5619);
nor U6316 (N_6316,N_5025,N_5500);
xnor U6317 (N_6317,N_4802,N_5810);
nor U6318 (N_6318,N_5094,N_5997);
xor U6319 (N_6319,N_4983,N_5659);
nor U6320 (N_6320,N_5756,N_4826);
xnor U6321 (N_6321,N_5573,N_4820);
and U6322 (N_6322,N_5924,N_5910);
or U6323 (N_6323,N_5637,N_5413);
or U6324 (N_6324,N_5560,N_5381);
or U6325 (N_6325,N_5048,N_5240);
xor U6326 (N_6326,N_5089,N_4929);
and U6327 (N_6327,N_5326,N_5477);
or U6328 (N_6328,N_5160,N_5846);
nand U6329 (N_6329,N_4841,N_5727);
or U6330 (N_6330,N_5200,N_5956);
nor U6331 (N_6331,N_4907,N_4978);
nor U6332 (N_6332,N_5906,N_4873);
nand U6333 (N_6333,N_4950,N_5030);
and U6334 (N_6334,N_5999,N_5881);
xnor U6335 (N_6335,N_5738,N_4919);
nor U6336 (N_6336,N_5213,N_5354);
xnor U6337 (N_6337,N_5797,N_5593);
or U6338 (N_6338,N_5436,N_5292);
nor U6339 (N_6339,N_5041,N_5242);
xnor U6340 (N_6340,N_5976,N_4872);
xor U6341 (N_6341,N_4823,N_5241);
nand U6342 (N_6342,N_4999,N_5186);
and U6343 (N_6343,N_5252,N_5774);
and U6344 (N_6344,N_4901,N_5179);
xnor U6345 (N_6345,N_5104,N_5187);
nor U6346 (N_6346,N_4874,N_5980);
or U6347 (N_6347,N_5744,N_5648);
nand U6348 (N_6348,N_5654,N_5540);
and U6349 (N_6349,N_5703,N_4937);
xnor U6350 (N_6350,N_5892,N_4912);
and U6351 (N_6351,N_5280,N_5582);
nand U6352 (N_6352,N_4855,N_5415);
nor U6353 (N_6353,N_4848,N_5060);
and U6354 (N_6354,N_5432,N_5020);
and U6355 (N_6355,N_5740,N_5592);
xnor U6356 (N_6356,N_5006,N_5221);
and U6357 (N_6357,N_4899,N_5255);
nand U6358 (N_6358,N_5849,N_5132);
nor U6359 (N_6359,N_5400,N_5554);
and U6360 (N_6360,N_5597,N_4916);
nand U6361 (N_6361,N_5748,N_5800);
and U6362 (N_6362,N_5443,N_5336);
nand U6363 (N_6363,N_5394,N_5546);
or U6364 (N_6364,N_5900,N_5114);
xnor U6365 (N_6365,N_4900,N_5837);
xnor U6366 (N_6366,N_4862,N_5521);
nor U6367 (N_6367,N_5056,N_5965);
nand U6368 (N_6368,N_5894,N_5831);
and U6369 (N_6369,N_5941,N_5812);
and U6370 (N_6370,N_5630,N_5567);
xnor U6371 (N_6371,N_4880,N_5151);
or U6372 (N_6372,N_5342,N_5347);
nor U6373 (N_6373,N_5749,N_4850);
nor U6374 (N_6374,N_4982,N_5075);
and U6375 (N_6375,N_5916,N_5734);
nand U6376 (N_6376,N_5818,N_5414);
xnor U6377 (N_6377,N_5697,N_5393);
or U6378 (N_6378,N_4827,N_5601);
xnor U6379 (N_6379,N_5694,N_5843);
or U6380 (N_6380,N_5789,N_4864);
xnor U6381 (N_6381,N_4952,N_5388);
nand U6382 (N_6382,N_5764,N_5828);
nor U6383 (N_6383,N_5315,N_5039);
or U6384 (N_6384,N_5758,N_4805);
and U6385 (N_6385,N_4988,N_5437);
xor U6386 (N_6386,N_5180,N_4863);
xor U6387 (N_6387,N_5520,N_5721);
nor U6388 (N_6388,N_5680,N_5281);
or U6389 (N_6389,N_5783,N_5813);
nand U6390 (N_6390,N_4835,N_5033);
nor U6391 (N_6391,N_4948,N_5308);
or U6392 (N_6392,N_5258,N_5723);
nand U6393 (N_6393,N_5272,N_5080);
xor U6394 (N_6394,N_5708,N_5298);
nor U6395 (N_6395,N_4803,N_5034);
or U6396 (N_6396,N_5571,N_5969);
or U6397 (N_6397,N_5019,N_5859);
or U6398 (N_6398,N_4822,N_5139);
nor U6399 (N_6399,N_5981,N_5455);
nor U6400 (N_6400,N_5073,N_5700);
and U6401 (N_6401,N_5093,N_5612);
xor U6402 (N_6402,N_5444,N_4966);
or U6403 (N_6403,N_4985,N_4890);
nor U6404 (N_6404,N_5362,N_4943);
nand U6405 (N_6405,N_5889,N_5890);
xor U6406 (N_6406,N_5848,N_5046);
or U6407 (N_6407,N_5808,N_5851);
xnor U6408 (N_6408,N_4975,N_4810);
xor U6409 (N_6409,N_5884,N_5496);
xnor U6410 (N_6410,N_5568,N_5908);
xor U6411 (N_6411,N_4875,N_5607);
or U6412 (N_6412,N_5864,N_5024);
nand U6413 (N_6413,N_5078,N_5882);
nand U6414 (N_6414,N_5379,N_5670);
nand U6415 (N_6415,N_5998,N_5079);
or U6416 (N_6416,N_5309,N_4913);
nand U6417 (N_6417,N_5214,N_4992);
or U6418 (N_6418,N_5243,N_4995);
and U6419 (N_6419,N_5205,N_5467);
or U6420 (N_6420,N_5752,N_5084);
and U6421 (N_6421,N_5313,N_5349);
nand U6422 (N_6422,N_5348,N_5473);
nand U6423 (N_6423,N_5031,N_5635);
xnor U6424 (N_6424,N_5755,N_4953);
and U6425 (N_6425,N_5422,N_5647);
or U6426 (N_6426,N_5673,N_5932);
nor U6427 (N_6427,N_5872,N_5809);
xor U6428 (N_6428,N_5988,N_5267);
nand U6429 (N_6429,N_5155,N_5543);
nor U6430 (N_6430,N_5491,N_5351);
nand U6431 (N_6431,N_5363,N_5153);
or U6432 (N_6432,N_5904,N_5973);
nand U6433 (N_6433,N_5961,N_5917);
nand U6434 (N_6434,N_5115,N_5712);
or U6435 (N_6435,N_5159,N_5815);
xor U6436 (N_6436,N_4891,N_5705);
and U6437 (N_6437,N_5515,N_5604);
nand U6438 (N_6438,N_5763,N_5944);
xnor U6439 (N_6439,N_4964,N_5949);
or U6440 (N_6440,N_5716,N_5356);
or U6441 (N_6441,N_5335,N_5737);
xnor U6442 (N_6442,N_5466,N_5494);
nand U6443 (N_6443,N_4984,N_5669);
or U6444 (N_6444,N_5923,N_5235);
or U6445 (N_6445,N_5853,N_5686);
xor U6446 (N_6446,N_5157,N_5043);
or U6447 (N_6447,N_5319,N_5247);
nand U6448 (N_6448,N_5427,N_5970);
xnor U6449 (N_6449,N_5501,N_5954);
or U6450 (N_6450,N_5461,N_5641);
nand U6451 (N_6451,N_5772,N_4977);
and U6452 (N_6452,N_5519,N_5805);
or U6453 (N_6453,N_5915,N_5049);
or U6454 (N_6454,N_4832,N_4915);
or U6455 (N_6455,N_5088,N_4861);
xor U6456 (N_6456,N_5779,N_5530);
or U6457 (N_6457,N_5490,N_5105);
nand U6458 (N_6458,N_5358,N_5707);
and U6459 (N_6459,N_5251,N_4996);
nor U6460 (N_6460,N_4969,N_4989);
and U6461 (N_6461,N_5841,N_5404);
or U6462 (N_6462,N_4808,N_5420);
xnor U6463 (N_6463,N_5288,N_5757);
nand U6464 (N_6464,N_5858,N_5537);
nand U6465 (N_6465,N_4800,N_5206);
nor U6466 (N_6466,N_4941,N_5219);
or U6467 (N_6467,N_4849,N_5962);
or U6468 (N_6468,N_5743,N_5010);
nand U6469 (N_6469,N_5294,N_5018);
nand U6470 (N_6470,N_5816,N_4883);
nor U6471 (N_6471,N_5745,N_5284);
nor U6472 (N_6472,N_5627,N_4825);
nand U6473 (N_6473,N_5173,N_5225);
and U6474 (N_6474,N_5911,N_4930);
xor U6475 (N_6475,N_5629,N_5481);
and U6476 (N_6476,N_5285,N_5107);
xnor U6477 (N_6477,N_4994,N_5803);
nand U6478 (N_6478,N_5784,N_5445);
and U6479 (N_6479,N_5840,N_5514);
xor U6480 (N_6480,N_5878,N_5984);
xnor U6481 (N_6481,N_5663,N_5947);
nor U6482 (N_6482,N_5121,N_5451);
and U6483 (N_6483,N_5350,N_5344);
nor U6484 (N_6484,N_5045,N_5131);
and U6485 (N_6485,N_5591,N_5989);
and U6486 (N_6486,N_5196,N_4852);
and U6487 (N_6487,N_5424,N_5204);
and U6488 (N_6488,N_5930,N_5430);
nand U6489 (N_6489,N_4979,N_5290);
xor U6490 (N_6490,N_5178,N_5143);
nand U6491 (N_6491,N_4882,N_5780);
xor U6492 (N_6492,N_5953,N_5992);
and U6493 (N_6493,N_5012,N_5689);
nand U6494 (N_6494,N_5154,N_5137);
nand U6495 (N_6495,N_5176,N_5547);
nand U6496 (N_6496,N_5822,N_5475);
nand U6497 (N_6497,N_5595,N_5017);
nor U6498 (N_6498,N_5778,N_5003);
xnor U6499 (N_6499,N_5960,N_4910);
nor U6500 (N_6500,N_5585,N_5674);
nor U6501 (N_6501,N_5655,N_5769);
xor U6502 (N_6502,N_5523,N_4847);
nand U6503 (N_6503,N_5428,N_5167);
nor U6504 (N_6504,N_5291,N_5254);
xnor U6505 (N_6505,N_5731,N_5488);
nand U6506 (N_6506,N_5061,N_5824);
nor U6507 (N_6507,N_5691,N_5861);
or U6508 (N_6508,N_5919,N_5541);
nand U6509 (N_6509,N_5072,N_5127);
nand U6510 (N_6510,N_5064,N_5806);
nand U6511 (N_6511,N_4867,N_5245);
xnor U6512 (N_6512,N_5937,N_4986);
or U6513 (N_6513,N_5274,N_5942);
or U6514 (N_6514,N_5276,N_5199);
or U6515 (N_6515,N_5135,N_5622);
or U6516 (N_6516,N_5042,N_5282);
or U6517 (N_6517,N_5355,N_5795);
or U6518 (N_6518,N_5742,N_5771);
and U6519 (N_6519,N_4970,N_5638);
and U6520 (N_6520,N_5902,N_4817);
nor U6521 (N_6521,N_5449,N_5528);
nand U6522 (N_6522,N_5628,N_5688);
xnor U6523 (N_6523,N_4837,N_5825);
and U6524 (N_6524,N_5977,N_5125);
nand U6525 (N_6525,N_5722,N_5928);
and U6526 (N_6526,N_5405,N_5130);
and U6527 (N_6527,N_5384,N_5418);
nor U6528 (N_6528,N_5223,N_5768);
and U6529 (N_6529,N_5190,N_5256);
and U6530 (N_6530,N_5529,N_5170);
xnor U6531 (N_6531,N_5346,N_4928);
nor U6532 (N_6532,N_4878,N_5660);
nor U6533 (N_6533,N_4834,N_5814);
nand U6534 (N_6534,N_5611,N_5982);
nand U6535 (N_6535,N_5040,N_5504);
or U6536 (N_6536,N_5513,N_5767);
xnor U6537 (N_6537,N_5985,N_5608);
nand U6538 (N_6538,N_5136,N_5926);
nand U6539 (N_6539,N_5311,N_5238);
and U6540 (N_6540,N_5993,N_5682);
xor U6541 (N_6541,N_5502,N_5651);
nand U6542 (N_6542,N_4974,N_5268);
or U6543 (N_6543,N_5790,N_5508);
nor U6544 (N_6544,N_5299,N_5548);
nand U6545 (N_6545,N_5729,N_4819);
nand U6546 (N_6546,N_5826,N_5469);
or U6547 (N_6547,N_5462,N_5210);
or U6548 (N_6548,N_5511,N_5950);
and U6549 (N_6549,N_5339,N_5352);
or U6550 (N_6550,N_5590,N_5559);
nor U6551 (N_6551,N_5510,N_5028);
xor U6552 (N_6552,N_5658,N_5855);
and U6553 (N_6553,N_5108,N_4909);
and U6554 (N_6554,N_5310,N_4971);
and U6555 (N_6555,N_5340,N_4853);
nor U6556 (N_6556,N_5456,N_5702);
xor U6557 (N_6557,N_4976,N_5920);
or U6558 (N_6558,N_5259,N_5054);
and U6559 (N_6559,N_5987,N_5518);
nand U6560 (N_6560,N_5102,N_5596);
xnor U6561 (N_6561,N_5092,N_5465);
and U6562 (N_6562,N_5880,N_4815);
xnor U6563 (N_6563,N_5052,N_4840);
and U6564 (N_6564,N_4845,N_4809);
and U6565 (N_6565,N_5398,N_5425);
or U6566 (N_6566,N_5698,N_4908);
nand U6567 (N_6567,N_5065,N_5895);
or U6568 (N_6568,N_5787,N_4925);
and U6569 (N_6569,N_5120,N_5802);
nand U6570 (N_6570,N_5566,N_5163);
or U6571 (N_6571,N_5164,N_5834);
nand U6572 (N_6572,N_5270,N_4962);
nand U6573 (N_6573,N_5382,N_5776);
xnor U6574 (N_6574,N_5922,N_4838);
nand U6575 (N_6575,N_5279,N_5704);
xnor U6576 (N_6576,N_5486,N_5933);
or U6577 (N_6577,N_5739,N_5857);
or U6578 (N_6578,N_5869,N_5112);
nor U6579 (N_6579,N_5248,N_5489);
nor U6580 (N_6580,N_5106,N_5693);
or U6581 (N_6581,N_5071,N_5668);
xnor U6582 (N_6582,N_5293,N_5021);
xor U6583 (N_6583,N_5320,N_4843);
nor U6584 (N_6584,N_5901,N_5527);
nor U6585 (N_6585,N_5057,N_5317);
xnor U6586 (N_6586,N_5532,N_5896);
nor U6587 (N_6587,N_5940,N_4858);
or U6588 (N_6588,N_5215,N_5736);
or U6589 (N_6589,N_5914,N_5865);
nand U6590 (N_6590,N_5314,N_5975);
or U6591 (N_6591,N_5140,N_4854);
or U6592 (N_6592,N_5578,N_5679);
nand U6593 (N_6593,N_5964,N_5844);
or U6594 (N_6594,N_5271,N_5007);
nand U6595 (N_6595,N_5118,N_5232);
and U6596 (N_6596,N_5014,N_5876);
nor U6597 (N_6597,N_5958,N_5782);
xor U6598 (N_6598,N_5921,N_5145);
nor U6599 (N_6599,N_5760,N_5788);
xor U6600 (N_6600,N_5470,N_5675);
xor U6601 (N_6601,N_5743,N_5386);
nor U6602 (N_6602,N_5400,N_4893);
nand U6603 (N_6603,N_5855,N_5659);
nor U6604 (N_6604,N_5929,N_4909);
nor U6605 (N_6605,N_5612,N_4890);
nor U6606 (N_6606,N_5273,N_4962);
nor U6607 (N_6607,N_5388,N_5152);
xnor U6608 (N_6608,N_5066,N_5030);
nor U6609 (N_6609,N_5761,N_5041);
nor U6610 (N_6610,N_5194,N_5705);
nor U6611 (N_6611,N_5929,N_5836);
nand U6612 (N_6612,N_5474,N_5774);
nor U6613 (N_6613,N_5866,N_5146);
nand U6614 (N_6614,N_5469,N_5210);
or U6615 (N_6615,N_5244,N_5453);
xnor U6616 (N_6616,N_5494,N_4937);
nand U6617 (N_6617,N_5659,N_5841);
nor U6618 (N_6618,N_5682,N_4928);
and U6619 (N_6619,N_5212,N_5961);
and U6620 (N_6620,N_5508,N_4914);
or U6621 (N_6621,N_5041,N_5741);
nor U6622 (N_6622,N_5071,N_5536);
nor U6623 (N_6623,N_5982,N_5845);
nand U6624 (N_6624,N_5946,N_4828);
and U6625 (N_6625,N_4817,N_5573);
nor U6626 (N_6626,N_5975,N_4970);
nor U6627 (N_6627,N_5737,N_5581);
nand U6628 (N_6628,N_5803,N_5833);
xnor U6629 (N_6629,N_5726,N_5638);
nor U6630 (N_6630,N_4813,N_5693);
and U6631 (N_6631,N_5707,N_5027);
nand U6632 (N_6632,N_5826,N_5635);
and U6633 (N_6633,N_5093,N_5330);
nand U6634 (N_6634,N_5430,N_4921);
nand U6635 (N_6635,N_5152,N_5471);
nand U6636 (N_6636,N_5825,N_5070);
nor U6637 (N_6637,N_5006,N_5687);
and U6638 (N_6638,N_5106,N_5431);
or U6639 (N_6639,N_5847,N_4869);
nand U6640 (N_6640,N_4884,N_5052);
or U6641 (N_6641,N_5273,N_4822);
xor U6642 (N_6642,N_5990,N_5240);
or U6643 (N_6643,N_5608,N_5190);
or U6644 (N_6644,N_5938,N_5286);
nor U6645 (N_6645,N_5224,N_5615);
or U6646 (N_6646,N_5252,N_4829);
xnor U6647 (N_6647,N_5419,N_5642);
nor U6648 (N_6648,N_5989,N_5125);
xor U6649 (N_6649,N_5320,N_5131);
and U6650 (N_6650,N_5126,N_5442);
or U6651 (N_6651,N_5494,N_5955);
and U6652 (N_6652,N_5486,N_5801);
nand U6653 (N_6653,N_5788,N_5230);
and U6654 (N_6654,N_5761,N_5537);
nor U6655 (N_6655,N_5662,N_5455);
nand U6656 (N_6656,N_5782,N_5729);
nand U6657 (N_6657,N_5580,N_4872);
or U6658 (N_6658,N_5408,N_4921);
xnor U6659 (N_6659,N_5089,N_5191);
and U6660 (N_6660,N_5874,N_5737);
and U6661 (N_6661,N_5656,N_5378);
and U6662 (N_6662,N_5271,N_5039);
xor U6663 (N_6663,N_5254,N_5421);
nor U6664 (N_6664,N_5634,N_5563);
and U6665 (N_6665,N_5109,N_4981);
or U6666 (N_6666,N_5079,N_5066);
or U6667 (N_6667,N_5513,N_5983);
xor U6668 (N_6668,N_5616,N_5456);
or U6669 (N_6669,N_5594,N_4981);
nor U6670 (N_6670,N_5644,N_5706);
and U6671 (N_6671,N_4873,N_5287);
nor U6672 (N_6672,N_5265,N_5493);
nand U6673 (N_6673,N_5352,N_5729);
nand U6674 (N_6674,N_5496,N_5054);
nand U6675 (N_6675,N_5297,N_5801);
xnor U6676 (N_6676,N_5297,N_5228);
or U6677 (N_6677,N_5005,N_4960);
nor U6678 (N_6678,N_5066,N_5179);
xnor U6679 (N_6679,N_5862,N_5512);
xnor U6680 (N_6680,N_5695,N_5026);
nor U6681 (N_6681,N_5400,N_4988);
nand U6682 (N_6682,N_5538,N_4815);
nor U6683 (N_6683,N_5978,N_5911);
or U6684 (N_6684,N_5319,N_5760);
nand U6685 (N_6685,N_4845,N_5081);
nor U6686 (N_6686,N_5186,N_5653);
nor U6687 (N_6687,N_5671,N_5907);
nand U6688 (N_6688,N_5582,N_5978);
or U6689 (N_6689,N_5340,N_4848);
or U6690 (N_6690,N_5012,N_5658);
xnor U6691 (N_6691,N_5503,N_5311);
or U6692 (N_6692,N_4901,N_5476);
nand U6693 (N_6693,N_5491,N_5823);
xnor U6694 (N_6694,N_5231,N_5837);
xnor U6695 (N_6695,N_5929,N_5827);
nand U6696 (N_6696,N_4882,N_5181);
nand U6697 (N_6697,N_5054,N_5732);
or U6698 (N_6698,N_5361,N_5621);
and U6699 (N_6699,N_5939,N_5911);
and U6700 (N_6700,N_5968,N_4876);
xor U6701 (N_6701,N_5486,N_5649);
nand U6702 (N_6702,N_5967,N_5740);
and U6703 (N_6703,N_4881,N_5492);
xor U6704 (N_6704,N_5757,N_5243);
and U6705 (N_6705,N_5948,N_5635);
or U6706 (N_6706,N_5579,N_4963);
nand U6707 (N_6707,N_5477,N_5530);
nand U6708 (N_6708,N_5744,N_5776);
or U6709 (N_6709,N_5079,N_4907);
nand U6710 (N_6710,N_5333,N_5133);
nor U6711 (N_6711,N_4833,N_5212);
or U6712 (N_6712,N_5548,N_5736);
xor U6713 (N_6713,N_5564,N_5486);
xor U6714 (N_6714,N_5915,N_5970);
or U6715 (N_6715,N_5220,N_5586);
nor U6716 (N_6716,N_5912,N_5559);
nand U6717 (N_6717,N_5780,N_5652);
nor U6718 (N_6718,N_5139,N_5352);
and U6719 (N_6719,N_4858,N_5818);
xor U6720 (N_6720,N_4806,N_5354);
or U6721 (N_6721,N_5217,N_4872);
nand U6722 (N_6722,N_5826,N_5926);
and U6723 (N_6723,N_4838,N_5872);
or U6724 (N_6724,N_5827,N_5517);
or U6725 (N_6725,N_4896,N_5975);
or U6726 (N_6726,N_5829,N_4815);
xnor U6727 (N_6727,N_5451,N_5242);
and U6728 (N_6728,N_5005,N_5831);
xor U6729 (N_6729,N_5420,N_5494);
nand U6730 (N_6730,N_5951,N_5857);
or U6731 (N_6731,N_5825,N_5456);
nand U6732 (N_6732,N_5100,N_5130);
or U6733 (N_6733,N_5956,N_5170);
and U6734 (N_6734,N_5553,N_5548);
or U6735 (N_6735,N_5121,N_5584);
xnor U6736 (N_6736,N_5715,N_5994);
and U6737 (N_6737,N_5107,N_5228);
nor U6738 (N_6738,N_5280,N_5446);
nor U6739 (N_6739,N_5766,N_5690);
and U6740 (N_6740,N_5120,N_5547);
nor U6741 (N_6741,N_5108,N_5585);
or U6742 (N_6742,N_5991,N_5840);
or U6743 (N_6743,N_5421,N_5264);
nand U6744 (N_6744,N_5339,N_5063);
xnor U6745 (N_6745,N_4884,N_4913);
and U6746 (N_6746,N_5594,N_5756);
nor U6747 (N_6747,N_5044,N_5172);
or U6748 (N_6748,N_5046,N_5977);
xnor U6749 (N_6749,N_4996,N_4828);
xor U6750 (N_6750,N_5081,N_4961);
nand U6751 (N_6751,N_4922,N_5013);
or U6752 (N_6752,N_5605,N_5876);
and U6753 (N_6753,N_5745,N_4905);
xnor U6754 (N_6754,N_5285,N_5932);
nand U6755 (N_6755,N_4962,N_5125);
and U6756 (N_6756,N_4955,N_5354);
nand U6757 (N_6757,N_5972,N_5612);
or U6758 (N_6758,N_5192,N_5567);
xnor U6759 (N_6759,N_5766,N_5078);
and U6760 (N_6760,N_5702,N_5760);
xor U6761 (N_6761,N_5392,N_5325);
xnor U6762 (N_6762,N_5667,N_5622);
xnor U6763 (N_6763,N_5427,N_5147);
xnor U6764 (N_6764,N_5194,N_5367);
nor U6765 (N_6765,N_5045,N_5284);
nand U6766 (N_6766,N_5064,N_4805);
nor U6767 (N_6767,N_5026,N_5597);
and U6768 (N_6768,N_5888,N_5904);
nand U6769 (N_6769,N_5174,N_5841);
nor U6770 (N_6770,N_5124,N_5430);
and U6771 (N_6771,N_5336,N_5379);
and U6772 (N_6772,N_4895,N_5196);
and U6773 (N_6773,N_4954,N_5465);
nand U6774 (N_6774,N_5819,N_4908);
or U6775 (N_6775,N_5777,N_5881);
xnor U6776 (N_6776,N_5973,N_5011);
xor U6777 (N_6777,N_5287,N_5884);
nor U6778 (N_6778,N_5429,N_5650);
nor U6779 (N_6779,N_4822,N_5773);
or U6780 (N_6780,N_5546,N_5488);
or U6781 (N_6781,N_4991,N_5408);
nand U6782 (N_6782,N_5690,N_5994);
or U6783 (N_6783,N_5947,N_5956);
or U6784 (N_6784,N_4828,N_4943);
and U6785 (N_6785,N_4963,N_5924);
nor U6786 (N_6786,N_5416,N_5986);
nand U6787 (N_6787,N_5256,N_5079);
or U6788 (N_6788,N_5453,N_5911);
nand U6789 (N_6789,N_5781,N_5008);
nand U6790 (N_6790,N_5991,N_5669);
nand U6791 (N_6791,N_5937,N_5224);
nor U6792 (N_6792,N_5340,N_5754);
and U6793 (N_6793,N_5821,N_4846);
nor U6794 (N_6794,N_5404,N_5175);
nor U6795 (N_6795,N_5523,N_4852);
nor U6796 (N_6796,N_4846,N_5364);
nor U6797 (N_6797,N_5338,N_5365);
and U6798 (N_6798,N_5278,N_5869);
and U6799 (N_6799,N_5437,N_5097);
or U6800 (N_6800,N_5222,N_4864);
xnor U6801 (N_6801,N_4845,N_5498);
nand U6802 (N_6802,N_5682,N_5895);
nor U6803 (N_6803,N_4934,N_4854);
and U6804 (N_6804,N_4892,N_5908);
or U6805 (N_6805,N_5448,N_5170);
or U6806 (N_6806,N_5293,N_5813);
xnor U6807 (N_6807,N_5188,N_5458);
nand U6808 (N_6808,N_4801,N_5774);
or U6809 (N_6809,N_5917,N_4939);
nand U6810 (N_6810,N_5251,N_5938);
and U6811 (N_6811,N_5094,N_5262);
nor U6812 (N_6812,N_5922,N_5940);
or U6813 (N_6813,N_5517,N_5793);
or U6814 (N_6814,N_5645,N_5870);
and U6815 (N_6815,N_5053,N_5422);
xnor U6816 (N_6816,N_5915,N_5434);
nand U6817 (N_6817,N_5111,N_5443);
nand U6818 (N_6818,N_5921,N_5742);
xnor U6819 (N_6819,N_5101,N_5304);
and U6820 (N_6820,N_4988,N_5206);
nand U6821 (N_6821,N_5845,N_5867);
nand U6822 (N_6822,N_5675,N_5249);
and U6823 (N_6823,N_5821,N_4963);
nor U6824 (N_6824,N_5790,N_4867);
and U6825 (N_6825,N_5620,N_5105);
and U6826 (N_6826,N_4985,N_5206);
xnor U6827 (N_6827,N_5980,N_5749);
xor U6828 (N_6828,N_5099,N_4874);
and U6829 (N_6829,N_5398,N_5971);
or U6830 (N_6830,N_5781,N_4891);
xor U6831 (N_6831,N_5160,N_5612);
and U6832 (N_6832,N_5624,N_5322);
or U6833 (N_6833,N_5580,N_5075);
or U6834 (N_6834,N_5749,N_5880);
or U6835 (N_6835,N_5887,N_5573);
or U6836 (N_6836,N_4930,N_4958);
and U6837 (N_6837,N_5717,N_5809);
and U6838 (N_6838,N_5343,N_4901);
nand U6839 (N_6839,N_5143,N_5304);
nand U6840 (N_6840,N_5353,N_4964);
xnor U6841 (N_6841,N_4953,N_5555);
nand U6842 (N_6842,N_5784,N_4917);
nor U6843 (N_6843,N_5934,N_5868);
and U6844 (N_6844,N_4939,N_5850);
and U6845 (N_6845,N_4907,N_4832);
or U6846 (N_6846,N_5660,N_5495);
or U6847 (N_6847,N_5949,N_5288);
nand U6848 (N_6848,N_5299,N_5698);
nor U6849 (N_6849,N_5154,N_5177);
nand U6850 (N_6850,N_5501,N_5725);
and U6851 (N_6851,N_5778,N_5805);
xnor U6852 (N_6852,N_5791,N_5404);
nand U6853 (N_6853,N_5115,N_5543);
nand U6854 (N_6854,N_5125,N_4935);
xor U6855 (N_6855,N_5706,N_5360);
and U6856 (N_6856,N_5942,N_4845);
and U6857 (N_6857,N_5267,N_5380);
and U6858 (N_6858,N_4932,N_5009);
or U6859 (N_6859,N_5148,N_5343);
or U6860 (N_6860,N_5412,N_5487);
and U6861 (N_6861,N_5130,N_4895);
and U6862 (N_6862,N_5223,N_5644);
and U6863 (N_6863,N_5265,N_5789);
or U6864 (N_6864,N_5125,N_5931);
or U6865 (N_6865,N_5264,N_5775);
nor U6866 (N_6866,N_5728,N_5371);
nor U6867 (N_6867,N_4807,N_5858);
or U6868 (N_6868,N_5156,N_5006);
xnor U6869 (N_6869,N_5056,N_4851);
and U6870 (N_6870,N_5736,N_5857);
or U6871 (N_6871,N_5985,N_5108);
nand U6872 (N_6872,N_5574,N_5652);
and U6873 (N_6873,N_4986,N_5341);
or U6874 (N_6874,N_5593,N_5870);
nand U6875 (N_6875,N_5691,N_5909);
and U6876 (N_6876,N_5304,N_5524);
or U6877 (N_6877,N_5034,N_5732);
or U6878 (N_6878,N_4977,N_5355);
or U6879 (N_6879,N_4866,N_5990);
nand U6880 (N_6880,N_5631,N_5179);
xnor U6881 (N_6881,N_5144,N_5638);
nand U6882 (N_6882,N_5515,N_5529);
and U6883 (N_6883,N_5730,N_5761);
and U6884 (N_6884,N_4961,N_5705);
and U6885 (N_6885,N_5100,N_5092);
or U6886 (N_6886,N_5614,N_5035);
xor U6887 (N_6887,N_5459,N_5918);
nor U6888 (N_6888,N_5353,N_5940);
nor U6889 (N_6889,N_4885,N_4875);
nand U6890 (N_6890,N_4883,N_5183);
nor U6891 (N_6891,N_5722,N_5035);
nand U6892 (N_6892,N_4917,N_5689);
nand U6893 (N_6893,N_4853,N_5536);
and U6894 (N_6894,N_4923,N_5748);
xnor U6895 (N_6895,N_5957,N_5284);
nand U6896 (N_6896,N_4810,N_5787);
nor U6897 (N_6897,N_5135,N_5513);
or U6898 (N_6898,N_5047,N_5467);
or U6899 (N_6899,N_5662,N_5603);
and U6900 (N_6900,N_4935,N_5572);
and U6901 (N_6901,N_5916,N_5614);
or U6902 (N_6902,N_5584,N_5442);
xor U6903 (N_6903,N_5205,N_5547);
nor U6904 (N_6904,N_5019,N_5707);
nor U6905 (N_6905,N_5857,N_5008);
or U6906 (N_6906,N_5716,N_5392);
nor U6907 (N_6907,N_5598,N_5956);
nand U6908 (N_6908,N_4823,N_5058);
nand U6909 (N_6909,N_5547,N_5124);
nor U6910 (N_6910,N_5876,N_5766);
nand U6911 (N_6911,N_5774,N_5778);
and U6912 (N_6912,N_5067,N_4870);
nand U6913 (N_6913,N_5003,N_5298);
xor U6914 (N_6914,N_5838,N_4943);
and U6915 (N_6915,N_5569,N_5950);
and U6916 (N_6916,N_5680,N_5834);
and U6917 (N_6917,N_5811,N_5447);
nor U6918 (N_6918,N_5123,N_5789);
nand U6919 (N_6919,N_4855,N_5459);
or U6920 (N_6920,N_4879,N_5556);
nor U6921 (N_6921,N_4912,N_5616);
and U6922 (N_6922,N_5139,N_5988);
xor U6923 (N_6923,N_4836,N_5709);
xor U6924 (N_6924,N_5411,N_4977);
and U6925 (N_6925,N_5133,N_4811);
and U6926 (N_6926,N_5649,N_5065);
nand U6927 (N_6927,N_5353,N_5118);
nor U6928 (N_6928,N_5763,N_5377);
and U6929 (N_6929,N_5575,N_5297);
and U6930 (N_6930,N_5370,N_5435);
and U6931 (N_6931,N_5789,N_5172);
and U6932 (N_6932,N_4863,N_5716);
xnor U6933 (N_6933,N_5734,N_5017);
nand U6934 (N_6934,N_4919,N_5627);
nor U6935 (N_6935,N_5438,N_5177);
and U6936 (N_6936,N_5236,N_5431);
xnor U6937 (N_6937,N_5737,N_5090);
xor U6938 (N_6938,N_5207,N_5580);
xor U6939 (N_6939,N_4877,N_5210);
xnor U6940 (N_6940,N_5029,N_5848);
nor U6941 (N_6941,N_5676,N_5037);
or U6942 (N_6942,N_5582,N_4933);
nand U6943 (N_6943,N_4910,N_5987);
xor U6944 (N_6944,N_5279,N_4897);
nor U6945 (N_6945,N_5899,N_4863);
and U6946 (N_6946,N_4875,N_5648);
xnor U6947 (N_6947,N_5766,N_5893);
and U6948 (N_6948,N_5775,N_5737);
nor U6949 (N_6949,N_5600,N_5630);
or U6950 (N_6950,N_5579,N_5940);
nor U6951 (N_6951,N_5551,N_5394);
nor U6952 (N_6952,N_5112,N_4995);
xnor U6953 (N_6953,N_5570,N_5152);
xor U6954 (N_6954,N_5515,N_5098);
xnor U6955 (N_6955,N_5917,N_4987);
or U6956 (N_6956,N_5870,N_5459);
and U6957 (N_6957,N_5332,N_5878);
nor U6958 (N_6958,N_5691,N_5074);
nor U6959 (N_6959,N_5395,N_4974);
and U6960 (N_6960,N_5576,N_4856);
xor U6961 (N_6961,N_5341,N_5649);
xnor U6962 (N_6962,N_5557,N_5451);
nand U6963 (N_6963,N_5964,N_5257);
nand U6964 (N_6964,N_5494,N_4822);
nand U6965 (N_6965,N_5302,N_5324);
or U6966 (N_6966,N_5022,N_5141);
xor U6967 (N_6967,N_5263,N_5668);
and U6968 (N_6968,N_5480,N_5521);
nand U6969 (N_6969,N_5505,N_5063);
and U6970 (N_6970,N_5036,N_5027);
nand U6971 (N_6971,N_5650,N_5313);
nand U6972 (N_6972,N_4990,N_5784);
nand U6973 (N_6973,N_5270,N_5259);
nand U6974 (N_6974,N_5592,N_5233);
nand U6975 (N_6975,N_5739,N_5938);
nor U6976 (N_6976,N_5357,N_5878);
nand U6977 (N_6977,N_5685,N_5504);
nor U6978 (N_6978,N_4815,N_5391);
nor U6979 (N_6979,N_4849,N_5919);
nor U6980 (N_6980,N_5056,N_5265);
and U6981 (N_6981,N_5422,N_5154);
or U6982 (N_6982,N_5561,N_5007);
or U6983 (N_6983,N_5900,N_5782);
or U6984 (N_6984,N_5915,N_5178);
nor U6985 (N_6985,N_5115,N_5927);
and U6986 (N_6986,N_5760,N_5851);
and U6987 (N_6987,N_5584,N_5406);
and U6988 (N_6988,N_5658,N_5791);
and U6989 (N_6989,N_4924,N_5021);
xor U6990 (N_6990,N_5481,N_5216);
nor U6991 (N_6991,N_5827,N_4864);
nand U6992 (N_6992,N_5472,N_5811);
or U6993 (N_6993,N_5933,N_5641);
xor U6994 (N_6994,N_5333,N_5218);
nand U6995 (N_6995,N_5490,N_5637);
or U6996 (N_6996,N_5842,N_4836);
and U6997 (N_6997,N_5097,N_5507);
nand U6998 (N_6998,N_5513,N_5208);
nand U6999 (N_6999,N_5044,N_5141);
xor U7000 (N_7000,N_4815,N_5241);
and U7001 (N_7001,N_5257,N_5631);
nand U7002 (N_7002,N_4817,N_4898);
or U7003 (N_7003,N_4837,N_5770);
and U7004 (N_7004,N_5197,N_5474);
and U7005 (N_7005,N_5830,N_5713);
xnor U7006 (N_7006,N_5739,N_5987);
nor U7007 (N_7007,N_4825,N_5369);
or U7008 (N_7008,N_5917,N_5438);
nand U7009 (N_7009,N_5815,N_4813);
nor U7010 (N_7010,N_5028,N_4950);
nand U7011 (N_7011,N_4923,N_5918);
nor U7012 (N_7012,N_5232,N_5679);
and U7013 (N_7013,N_5939,N_5704);
and U7014 (N_7014,N_5066,N_5083);
xor U7015 (N_7015,N_5668,N_5564);
xor U7016 (N_7016,N_5384,N_4809);
xnor U7017 (N_7017,N_4812,N_5014);
nand U7018 (N_7018,N_5805,N_5366);
nand U7019 (N_7019,N_5089,N_5941);
nand U7020 (N_7020,N_5539,N_5926);
nor U7021 (N_7021,N_4987,N_5274);
and U7022 (N_7022,N_5976,N_4803);
nand U7023 (N_7023,N_5981,N_5730);
nand U7024 (N_7024,N_5934,N_5439);
or U7025 (N_7025,N_5972,N_5377);
or U7026 (N_7026,N_5708,N_5972);
nor U7027 (N_7027,N_5579,N_5388);
xnor U7028 (N_7028,N_4961,N_5094);
and U7029 (N_7029,N_5513,N_4816);
nand U7030 (N_7030,N_5054,N_5583);
and U7031 (N_7031,N_4891,N_4944);
nand U7032 (N_7032,N_5119,N_5078);
xor U7033 (N_7033,N_5803,N_5157);
nand U7034 (N_7034,N_5053,N_5380);
xnor U7035 (N_7035,N_5776,N_5121);
or U7036 (N_7036,N_5579,N_5629);
nand U7037 (N_7037,N_5269,N_4935);
nand U7038 (N_7038,N_5713,N_4880);
nand U7039 (N_7039,N_5248,N_5613);
and U7040 (N_7040,N_5854,N_4925);
nor U7041 (N_7041,N_5944,N_5192);
or U7042 (N_7042,N_5331,N_5108);
and U7043 (N_7043,N_4824,N_5727);
nand U7044 (N_7044,N_4804,N_5474);
nand U7045 (N_7045,N_5588,N_5920);
and U7046 (N_7046,N_5257,N_5667);
and U7047 (N_7047,N_5048,N_4997);
or U7048 (N_7048,N_4907,N_5153);
or U7049 (N_7049,N_4962,N_5496);
or U7050 (N_7050,N_5961,N_5222);
nand U7051 (N_7051,N_5567,N_5258);
and U7052 (N_7052,N_4814,N_5407);
nand U7053 (N_7053,N_5447,N_5832);
nor U7054 (N_7054,N_5633,N_4917);
and U7055 (N_7055,N_5112,N_5546);
and U7056 (N_7056,N_5724,N_5830);
and U7057 (N_7057,N_5768,N_5952);
and U7058 (N_7058,N_5253,N_5214);
nor U7059 (N_7059,N_5131,N_5023);
or U7060 (N_7060,N_5616,N_5966);
xnor U7061 (N_7061,N_5716,N_5149);
nand U7062 (N_7062,N_5120,N_5018);
xnor U7063 (N_7063,N_5744,N_5014);
xnor U7064 (N_7064,N_5049,N_5177);
nor U7065 (N_7065,N_5605,N_5986);
nor U7066 (N_7066,N_5006,N_5483);
xor U7067 (N_7067,N_5180,N_5962);
xnor U7068 (N_7068,N_5647,N_4847);
or U7069 (N_7069,N_5358,N_5232);
nor U7070 (N_7070,N_5636,N_5549);
or U7071 (N_7071,N_4938,N_5197);
or U7072 (N_7072,N_5819,N_5754);
or U7073 (N_7073,N_5208,N_5897);
and U7074 (N_7074,N_5187,N_5416);
nor U7075 (N_7075,N_5589,N_5764);
or U7076 (N_7076,N_5522,N_5003);
nor U7077 (N_7077,N_5033,N_4918);
or U7078 (N_7078,N_5868,N_5858);
and U7079 (N_7079,N_5736,N_5832);
nand U7080 (N_7080,N_5412,N_5822);
nand U7081 (N_7081,N_5228,N_5873);
or U7082 (N_7082,N_5815,N_5749);
nor U7083 (N_7083,N_4834,N_4969);
nor U7084 (N_7084,N_5081,N_5042);
nor U7085 (N_7085,N_5485,N_5484);
and U7086 (N_7086,N_5371,N_4962);
nand U7087 (N_7087,N_5125,N_5794);
nand U7088 (N_7088,N_5822,N_4828);
nor U7089 (N_7089,N_5231,N_5497);
and U7090 (N_7090,N_5572,N_5171);
or U7091 (N_7091,N_5210,N_5429);
and U7092 (N_7092,N_5912,N_5056);
or U7093 (N_7093,N_5922,N_5904);
xor U7094 (N_7094,N_5200,N_5516);
or U7095 (N_7095,N_5698,N_5281);
nor U7096 (N_7096,N_5480,N_5224);
or U7097 (N_7097,N_5295,N_5195);
nand U7098 (N_7098,N_5771,N_5384);
nand U7099 (N_7099,N_5086,N_5011);
nand U7100 (N_7100,N_5561,N_5726);
nand U7101 (N_7101,N_5369,N_5129);
nand U7102 (N_7102,N_5477,N_5128);
or U7103 (N_7103,N_5222,N_5300);
or U7104 (N_7104,N_5166,N_5585);
nor U7105 (N_7105,N_5444,N_5741);
or U7106 (N_7106,N_5024,N_5590);
and U7107 (N_7107,N_5584,N_4956);
nor U7108 (N_7108,N_5524,N_5355);
or U7109 (N_7109,N_5419,N_5450);
and U7110 (N_7110,N_5456,N_5387);
nand U7111 (N_7111,N_5688,N_5935);
xor U7112 (N_7112,N_5223,N_4811);
nor U7113 (N_7113,N_5619,N_5568);
nor U7114 (N_7114,N_5062,N_5360);
and U7115 (N_7115,N_5464,N_5792);
nor U7116 (N_7116,N_5295,N_5098);
nand U7117 (N_7117,N_5981,N_5043);
or U7118 (N_7118,N_4949,N_5556);
and U7119 (N_7119,N_5430,N_4944);
and U7120 (N_7120,N_5714,N_4846);
and U7121 (N_7121,N_5028,N_5966);
nor U7122 (N_7122,N_5057,N_4860);
and U7123 (N_7123,N_5870,N_5160);
nor U7124 (N_7124,N_5273,N_5270);
or U7125 (N_7125,N_4983,N_4869);
xnor U7126 (N_7126,N_5577,N_5963);
xnor U7127 (N_7127,N_5102,N_5442);
xnor U7128 (N_7128,N_5219,N_5931);
nor U7129 (N_7129,N_5092,N_5801);
nand U7130 (N_7130,N_4818,N_5316);
nor U7131 (N_7131,N_5791,N_5968);
and U7132 (N_7132,N_5706,N_5879);
nand U7133 (N_7133,N_4902,N_4919);
nand U7134 (N_7134,N_5137,N_4830);
or U7135 (N_7135,N_5129,N_5032);
nand U7136 (N_7136,N_5856,N_4954);
nand U7137 (N_7137,N_4823,N_5286);
nand U7138 (N_7138,N_5502,N_5552);
nor U7139 (N_7139,N_5168,N_5927);
or U7140 (N_7140,N_5433,N_5488);
and U7141 (N_7141,N_5012,N_5822);
nand U7142 (N_7142,N_5181,N_4853);
nand U7143 (N_7143,N_5185,N_5711);
xor U7144 (N_7144,N_5251,N_5351);
nor U7145 (N_7145,N_5432,N_4889);
xnor U7146 (N_7146,N_5524,N_5777);
nand U7147 (N_7147,N_5825,N_4931);
nor U7148 (N_7148,N_5072,N_5456);
or U7149 (N_7149,N_5968,N_5748);
nor U7150 (N_7150,N_5690,N_5659);
xor U7151 (N_7151,N_5493,N_4843);
nand U7152 (N_7152,N_4967,N_5249);
or U7153 (N_7153,N_5402,N_5654);
nor U7154 (N_7154,N_5319,N_5323);
nand U7155 (N_7155,N_5063,N_4801);
nor U7156 (N_7156,N_5250,N_5006);
or U7157 (N_7157,N_4933,N_5349);
or U7158 (N_7158,N_5711,N_5265);
xnor U7159 (N_7159,N_5032,N_5174);
and U7160 (N_7160,N_5452,N_4985);
nor U7161 (N_7161,N_5554,N_5528);
nand U7162 (N_7162,N_5107,N_5220);
nor U7163 (N_7163,N_4942,N_5660);
nor U7164 (N_7164,N_5128,N_5947);
and U7165 (N_7165,N_4834,N_5617);
nand U7166 (N_7166,N_5984,N_5080);
nand U7167 (N_7167,N_5945,N_5604);
or U7168 (N_7168,N_4927,N_4935);
xor U7169 (N_7169,N_5942,N_5619);
nand U7170 (N_7170,N_5218,N_5548);
nor U7171 (N_7171,N_5394,N_5532);
nor U7172 (N_7172,N_5195,N_5033);
and U7173 (N_7173,N_5746,N_5505);
xor U7174 (N_7174,N_5237,N_4986);
nor U7175 (N_7175,N_5545,N_5347);
nand U7176 (N_7176,N_5074,N_5649);
or U7177 (N_7177,N_5102,N_5976);
xnor U7178 (N_7178,N_5021,N_5463);
or U7179 (N_7179,N_5901,N_5591);
nor U7180 (N_7180,N_5725,N_5769);
or U7181 (N_7181,N_5608,N_5238);
and U7182 (N_7182,N_5901,N_5392);
xnor U7183 (N_7183,N_5445,N_5519);
nor U7184 (N_7184,N_5031,N_5327);
and U7185 (N_7185,N_5754,N_5782);
xnor U7186 (N_7186,N_4985,N_5021);
or U7187 (N_7187,N_5932,N_4850);
nand U7188 (N_7188,N_5301,N_5382);
or U7189 (N_7189,N_5591,N_5059);
nor U7190 (N_7190,N_5401,N_5929);
or U7191 (N_7191,N_5430,N_5955);
nand U7192 (N_7192,N_5472,N_5685);
and U7193 (N_7193,N_5160,N_5292);
xor U7194 (N_7194,N_5035,N_5796);
and U7195 (N_7195,N_5111,N_5928);
nand U7196 (N_7196,N_5196,N_5640);
or U7197 (N_7197,N_5868,N_5552);
and U7198 (N_7198,N_4894,N_5254);
nor U7199 (N_7199,N_5989,N_5141);
nand U7200 (N_7200,N_6667,N_6716);
and U7201 (N_7201,N_6108,N_6597);
xnor U7202 (N_7202,N_6695,N_6913);
nor U7203 (N_7203,N_7066,N_6100);
xor U7204 (N_7204,N_6902,N_6816);
or U7205 (N_7205,N_6187,N_6367);
xor U7206 (N_7206,N_7123,N_6555);
and U7207 (N_7207,N_6068,N_7153);
nor U7208 (N_7208,N_6456,N_6674);
xnor U7209 (N_7209,N_6861,N_6118);
nor U7210 (N_7210,N_6749,N_6178);
nand U7211 (N_7211,N_6059,N_7142);
or U7212 (N_7212,N_6912,N_7107);
xor U7213 (N_7213,N_6755,N_6951);
or U7214 (N_7214,N_6840,N_6579);
or U7215 (N_7215,N_6741,N_7100);
and U7216 (N_7216,N_6857,N_6314);
nand U7217 (N_7217,N_6327,N_6705);
nor U7218 (N_7218,N_6486,N_6159);
nor U7219 (N_7219,N_6806,N_7037);
xor U7220 (N_7220,N_6039,N_7036);
nand U7221 (N_7221,N_6591,N_7167);
nor U7222 (N_7222,N_6265,N_6718);
and U7223 (N_7223,N_7012,N_6814);
and U7224 (N_7224,N_6169,N_6771);
nand U7225 (N_7225,N_6583,N_6623);
nand U7226 (N_7226,N_6246,N_7094);
xor U7227 (N_7227,N_6789,N_6150);
xor U7228 (N_7228,N_6323,N_6062);
nor U7229 (N_7229,N_6550,N_6981);
nor U7230 (N_7230,N_6375,N_6945);
nand U7231 (N_7231,N_6321,N_6934);
and U7232 (N_7232,N_6040,N_7067);
xor U7233 (N_7233,N_6032,N_6887);
nor U7234 (N_7234,N_6202,N_6878);
and U7235 (N_7235,N_6601,N_7166);
nor U7236 (N_7236,N_7060,N_6948);
or U7237 (N_7237,N_6698,N_6799);
or U7238 (N_7238,N_6443,N_7160);
nor U7239 (N_7239,N_6551,N_6368);
xor U7240 (N_7240,N_7186,N_6464);
and U7241 (N_7241,N_6885,N_6297);
xor U7242 (N_7242,N_6562,N_6292);
and U7243 (N_7243,N_6490,N_6166);
nor U7244 (N_7244,N_7175,N_6198);
or U7245 (N_7245,N_6004,N_6145);
nand U7246 (N_7246,N_6742,N_6659);
and U7247 (N_7247,N_6067,N_7120);
nand U7248 (N_7248,N_6684,N_6725);
xor U7249 (N_7249,N_7171,N_6071);
or U7250 (N_7250,N_6869,N_6179);
xor U7251 (N_7251,N_6495,N_6838);
and U7252 (N_7252,N_6304,N_6324);
xor U7253 (N_7253,N_6489,N_6434);
nor U7254 (N_7254,N_7141,N_6706);
xnor U7255 (N_7255,N_6989,N_6578);
or U7256 (N_7256,N_6964,N_6979);
xnor U7257 (N_7257,N_6011,N_6332);
xnor U7258 (N_7258,N_6310,N_6022);
or U7259 (N_7259,N_6263,N_6113);
nand U7260 (N_7260,N_6774,N_6135);
nand U7261 (N_7261,N_6782,N_6231);
nand U7262 (N_7262,N_6636,N_6300);
nor U7263 (N_7263,N_6326,N_6407);
or U7264 (N_7264,N_6256,N_6549);
nand U7265 (N_7265,N_6240,N_6573);
nand U7266 (N_7266,N_6439,N_7140);
xnor U7267 (N_7267,N_6516,N_6472);
xor U7268 (N_7268,N_6897,N_6270);
nor U7269 (N_7269,N_7097,N_6756);
xor U7270 (N_7270,N_7195,N_7013);
or U7271 (N_7271,N_6763,N_6946);
nor U7272 (N_7272,N_6491,N_6820);
xnor U7273 (N_7273,N_6156,N_6104);
or U7274 (N_7274,N_6947,N_7130);
nor U7275 (N_7275,N_6512,N_6365);
nand U7276 (N_7276,N_6037,N_6249);
or U7277 (N_7277,N_6079,N_6908);
and U7278 (N_7278,N_6160,N_6501);
nor U7279 (N_7279,N_6538,N_6959);
nand U7280 (N_7280,N_6590,N_6410);
and U7281 (N_7281,N_6053,N_6452);
nor U7282 (N_7282,N_6301,N_7178);
xnor U7283 (N_7283,N_6877,N_6691);
nor U7284 (N_7284,N_6313,N_6626);
and U7285 (N_7285,N_6128,N_6124);
xnor U7286 (N_7286,N_6349,N_6704);
nand U7287 (N_7287,N_6149,N_6077);
nand U7288 (N_7288,N_6228,N_6420);
and U7289 (N_7289,N_6517,N_7074);
nand U7290 (N_7290,N_6494,N_6248);
nand U7291 (N_7291,N_6033,N_6143);
nor U7292 (N_7292,N_6038,N_6086);
or U7293 (N_7293,N_6386,N_6261);
and U7294 (N_7294,N_6561,N_7154);
nand U7295 (N_7295,N_6405,N_6969);
xnor U7296 (N_7296,N_7000,N_6307);
xnor U7297 (N_7297,N_6835,N_6226);
xnor U7298 (N_7298,N_6459,N_6970);
or U7299 (N_7299,N_6176,N_6834);
and U7300 (N_7300,N_6640,N_7053);
xnor U7301 (N_7301,N_6660,N_6546);
nand U7302 (N_7302,N_7134,N_7043);
and U7303 (N_7303,N_6492,N_6938);
or U7304 (N_7304,N_6006,N_6708);
xnor U7305 (N_7305,N_6031,N_7073);
nor U7306 (N_7306,N_6556,N_6347);
or U7307 (N_7307,N_6144,N_7090);
xnor U7308 (N_7308,N_6302,N_6264);
and U7309 (N_7309,N_6414,N_6074);
nand U7310 (N_7310,N_6852,N_7092);
nand U7311 (N_7311,N_6277,N_6711);
or U7312 (N_7312,N_6670,N_7014);
nor U7313 (N_7313,N_6115,N_6847);
and U7314 (N_7314,N_6474,N_7185);
nand U7315 (N_7315,N_6273,N_7125);
and U7316 (N_7316,N_6880,N_6163);
nor U7317 (N_7317,N_6227,N_6987);
nand U7318 (N_7318,N_6889,N_7118);
or U7319 (N_7319,N_7006,N_6668);
or U7320 (N_7320,N_6268,N_6120);
or U7321 (N_7321,N_6453,N_6567);
nand U7322 (N_7322,N_6282,N_6728);
and U7323 (N_7323,N_7165,N_6131);
nor U7324 (N_7324,N_6041,N_6221);
xor U7325 (N_7325,N_6960,N_7001);
nand U7326 (N_7326,N_6823,N_6577);
xnor U7327 (N_7327,N_7071,N_6236);
nor U7328 (N_7328,N_6449,N_7061);
nor U7329 (N_7329,N_6648,N_6210);
nand U7330 (N_7330,N_6915,N_6543);
and U7331 (N_7331,N_6588,N_6418);
nand U7332 (N_7332,N_6585,N_6726);
nand U7333 (N_7333,N_6180,N_6436);
xnor U7334 (N_7334,N_6552,N_6493);
nor U7335 (N_7335,N_6213,N_6421);
nand U7336 (N_7336,N_6170,N_7148);
or U7337 (N_7337,N_6230,N_6614);
nor U7338 (N_7338,N_6111,N_6057);
nand U7339 (N_7339,N_6682,N_6744);
nor U7340 (N_7340,N_6023,N_6500);
xor U7341 (N_7341,N_6098,N_7193);
nor U7342 (N_7342,N_6865,N_7104);
xnor U7343 (N_7343,N_6557,N_6600);
nor U7344 (N_7344,N_6338,N_7045);
and U7345 (N_7345,N_6345,N_6630);
or U7346 (N_7346,N_7032,N_6027);
or U7347 (N_7347,N_6800,N_6048);
and U7348 (N_7348,N_6362,N_6566);
nand U7349 (N_7349,N_6432,N_6205);
or U7350 (N_7350,N_6101,N_6404);
or U7351 (N_7351,N_6563,N_6753);
nor U7352 (N_7352,N_6408,N_6446);
or U7353 (N_7353,N_7025,N_6141);
nor U7354 (N_7354,N_6433,N_6147);
or U7355 (N_7355,N_7190,N_6119);
and U7356 (N_7356,N_6978,N_6721);
nor U7357 (N_7357,N_6919,N_6707);
nand U7358 (N_7358,N_6528,N_6985);
nand U7359 (N_7359,N_6849,N_6051);
and U7360 (N_7360,N_6589,N_6424);
nor U7361 (N_7361,N_6322,N_7191);
and U7362 (N_7362,N_6672,N_6717);
or U7363 (N_7363,N_6503,N_6968);
nor U7364 (N_7364,N_7114,N_6036);
and U7365 (N_7365,N_6905,N_6003);
and U7366 (N_7366,N_6060,N_6758);
and U7367 (N_7367,N_6123,N_6233);
and U7368 (N_7368,N_7068,N_6117);
nor U7369 (N_7369,N_7021,N_6257);
or U7370 (N_7370,N_6457,N_6328);
xnor U7371 (N_7371,N_6883,N_6344);
nand U7372 (N_7372,N_6770,N_6351);
or U7373 (N_7373,N_6531,N_6625);
or U7374 (N_7374,N_6533,N_6653);
nand U7375 (N_7375,N_6211,N_6366);
nand U7376 (N_7376,N_7054,N_6502);
nor U7377 (N_7377,N_7170,N_6862);
and U7378 (N_7378,N_6102,N_7112);
nor U7379 (N_7379,N_6133,N_6958);
nor U7380 (N_7380,N_7151,N_7188);
nand U7381 (N_7381,N_6757,N_6088);
nand U7382 (N_7382,N_6631,N_6182);
nand U7383 (N_7383,N_6805,N_6988);
nor U7384 (N_7384,N_6406,N_6496);
nand U7385 (N_7385,N_6218,N_6423);
nor U7386 (N_7386,N_6641,N_6200);
and U7387 (N_7387,N_6786,N_7145);
and U7388 (N_7388,N_6899,N_6007);
nand U7389 (N_7389,N_6610,N_7059);
xor U7390 (N_7390,N_6678,N_6825);
xnor U7391 (N_7391,N_6188,N_6593);
xnor U7392 (N_7392,N_6854,N_6099);
nor U7393 (N_7393,N_7122,N_6035);
nand U7394 (N_7394,N_6642,N_6515);
xnor U7395 (N_7395,N_6925,N_6448);
nor U7396 (N_7396,N_6398,N_6943);
and U7397 (N_7397,N_7091,N_6542);
xor U7398 (N_7398,N_7124,N_6308);
xnor U7399 (N_7399,N_6703,N_7121);
and U7400 (N_7400,N_6372,N_6656);
nand U7401 (N_7401,N_7108,N_7144);
nand U7402 (N_7402,N_6910,N_6193);
xnor U7403 (N_7403,N_6477,N_6454);
xor U7404 (N_7404,N_7041,N_7087);
xnor U7405 (N_7405,N_7076,N_6204);
xnor U7406 (N_7406,N_6731,N_7176);
nand U7407 (N_7407,N_6613,N_6397);
or U7408 (N_7408,N_6941,N_6649);
nor U7409 (N_7409,N_7016,N_7005);
and U7410 (N_7410,N_6203,N_6252);
xnor U7411 (N_7411,N_6280,N_6030);
xor U7412 (N_7412,N_7198,N_6760);
nand U7413 (N_7413,N_7056,N_6339);
or U7414 (N_7414,N_6522,N_7040);
or U7415 (N_7415,N_6949,N_6821);
nand U7416 (N_7416,N_6441,N_7137);
nand U7417 (N_7417,N_6871,N_6956);
and U7418 (N_7418,N_6394,N_7046);
or U7419 (N_7419,N_6199,N_7075);
nand U7420 (N_7420,N_7180,N_7164);
and U7421 (N_7421,N_6914,N_6984);
and U7422 (N_7422,N_6173,N_6042);
nor U7423 (N_7423,N_6665,N_6009);
nor U7424 (N_7424,N_6330,N_6999);
nand U7425 (N_7425,N_7020,N_6831);
and U7426 (N_7426,N_7017,N_6860);
and U7427 (N_7427,N_7030,N_6291);
xor U7428 (N_7428,N_6629,N_7050);
or U7429 (N_7429,N_6076,N_6652);
nor U7430 (N_7430,N_6888,N_6468);
xnor U7431 (N_7431,N_6944,N_6891);
or U7432 (N_7432,N_6681,N_6957);
nor U7433 (N_7433,N_6244,N_6873);
nor U7434 (N_7434,N_6920,N_6875);
or U7435 (N_7435,N_7031,N_6982);
nand U7436 (N_7436,N_6829,N_6937);
xor U7437 (N_7437,N_7085,N_6019);
nor U7438 (N_7438,N_7058,N_7177);
nand U7439 (N_7439,N_6139,N_6933);
nand U7440 (N_7440,N_6499,N_6470);
xnor U7441 (N_7441,N_6797,N_6317);
nand U7442 (N_7442,N_6609,N_6377);
nor U7443 (N_7443,N_6824,N_6923);
and U7444 (N_7444,N_6810,N_6391);
nand U7445 (N_7445,N_6565,N_6225);
nor U7446 (N_7446,N_6052,N_7081);
or U7447 (N_7447,N_6673,N_6637);
nor U7448 (N_7448,N_7172,N_6378);
and U7449 (N_7449,N_6966,N_6991);
xor U7450 (N_7450,N_6392,N_6206);
or U7451 (N_7451,N_6016,N_6220);
or U7452 (N_7452,N_7182,N_6374);
nand U7453 (N_7453,N_6055,N_6662);
xnor U7454 (N_7454,N_6442,N_6903);
or U7455 (N_7455,N_6882,N_6622);
nor U7456 (N_7456,N_6005,N_6901);
and U7457 (N_7457,N_6851,N_7055);
or U7458 (N_7458,N_6801,N_7117);
xor U7459 (N_7459,N_6954,N_6632);
nand U7460 (N_7460,N_6222,N_6402);
or U7461 (N_7461,N_6780,N_6808);
xor U7462 (N_7462,N_6217,N_6072);
nand U7463 (N_7463,N_6788,N_6255);
xor U7464 (N_7464,N_6177,N_6535);
nor U7465 (N_7465,N_6661,N_6373);
nand U7466 (N_7466,N_6646,N_6769);
and U7467 (N_7467,N_6026,N_6034);
nand U7468 (N_7468,N_6395,N_6971);
and U7469 (N_7469,N_6025,N_6012);
nand U7470 (N_7470,N_6017,N_6754);
or U7471 (N_7471,N_6315,N_6603);
and U7472 (N_7472,N_6570,N_6895);
nand U7473 (N_7473,N_6858,N_6592);
nor U7474 (N_7474,N_6864,N_6109);
and U7475 (N_7475,N_6953,N_6384);
nor U7476 (N_7476,N_6643,N_6400);
nand U7477 (N_7477,N_6746,N_6275);
nor U7478 (N_7478,N_6605,N_6724);
or U7479 (N_7479,N_6267,N_6010);
or U7480 (N_7480,N_6709,N_6066);
and U7481 (N_7481,N_6689,N_7129);
or U7482 (N_7482,N_6548,N_6738);
nor U7483 (N_7483,N_7022,N_6606);
and U7484 (N_7484,N_6921,N_6096);
nand U7485 (N_7485,N_6740,N_6281);
nand U7486 (N_7486,N_6331,N_6276);
nor U7487 (N_7487,N_6319,N_6734);
and U7488 (N_7488,N_7103,N_6463);
nor U7489 (N_7489,N_6973,N_7086);
xnor U7490 (N_7490,N_6791,N_6475);
nor U7491 (N_7491,N_6369,N_6427);
or U7492 (N_7492,N_6986,N_6761);
or U7493 (N_7493,N_6942,N_6867);
and U7494 (N_7494,N_6993,N_6014);
nor U7495 (N_7495,N_6465,N_6998);
nand U7496 (N_7496,N_6142,N_6361);
nor U7497 (N_7497,N_6239,N_6584);
and U7498 (N_7498,N_7033,N_6803);
and U7499 (N_7499,N_6950,N_6827);
and U7500 (N_7500,N_6751,N_6994);
nand U7501 (N_7501,N_6795,N_6136);
and U7502 (N_7502,N_6461,N_6337);
xor U7503 (N_7503,N_7105,N_7136);
or U7504 (N_7504,N_6532,N_6214);
nand U7505 (N_7505,N_7065,N_7062);
and U7506 (N_7506,N_6116,N_6881);
nand U7507 (N_7507,N_6008,N_6965);
or U7508 (N_7508,N_6839,N_6259);
nand U7509 (N_7509,N_6747,N_6855);
nor U7510 (N_7510,N_6828,N_7199);
xor U7511 (N_7511,N_6476,N_6201);
nand U7512 (N_7512,N_6572,N_6483);
nor U7513 (N_7513,N_6272,N_6644);
nand U7514 (N_7514,N_6853,N_6967);
xnor U7515 (N_7515,N_7052,N_6168);
or U7516 (N_7516,N_6429,N_6929);
xnor U7517 (N_7517,N_6767,N_6049);
nand U7518 (N_7518,N_6237,N_6604);
nand U7519 (N_7519,N_6768,N_6254);
xnor U7520 (N_7520,N_6510,N_6387);
nor U7521 (N_7521,N_6872,N_7029);
xor U7522 (N_7522,N_6916,N_7133);
xnor U7523 (N_7523,N_6303,N_7039);
xnor U7524 (N_7524,N_6242,N_6155);
nor U7525 (N_7525,N_6093,N_6759);
or U7526 (N_7526,N_6107,N_6422);
or U7527 (N_7527,N_6262,N_6298);
nand U7528 (N_7528,N_6634,N_6061);
nor U7529 (N_7529,N_6320,N_6822);
xnor U7530 (N_7530,N_6364,N_7098);
and U7531 (N_7531,N_6140,N_6287);
and U7532 (N_7532,N_6930,N_6359);
and U7533 (N_7533,N_7146,N_6952);
nand U7534 (N_7534,N_6666,N_7174);
nor U7535 (N_7535,N_6787,N_6075);
nand U7536 (N_7536,N_6195,N_6935);
xor U7537 (N_7537,N_7027,N_6092);
nand U7538 (N_7538,N_7102,N_6018);
nand U7539 (N_7539,N_7109,N_6207);
xnor U7540 (N_7540,N_6876,N_6064);
or U7541 (N_7541,N_6393,N_6932);
xor U7542 (N_7542,N_6683,N_7083);
xnor U7543 (N_7543,N_6874,N_6779);
and U7544 (N_7544,N_6560,N_6306);
nand U7545 (N_7545,N_6348,N_6485);
or U7546 (N_7546,N_7111,N_6299);
nor U7547 (N_7547,N_6274,N_6411);
or U7548 (N_7548,N_6333,N_6258);
nor U7549 (N_7549,N_6480,N_7018);
or U7550 (N_7550,N_6545,N_6544);
nand U7551 (N_7551,N_6296,N_7082);
and U7552 (N_7552,N_6918,N_6574);
nor U7553 (N_7553,N_6358,N_7197);
nand U7554 (N_7554,N_6151,N_6190);
and U7555 (N_7555,N_7034,N_6680);
and U7556 (N_7556,N_6633,N_7077);
or U7557 (N_7557,N_6762,N_7064);
nor U7558 (N_7558,N_6430,N_7155);
or U7559 (N_7559,N_6509,N_6000);
nand U7560 (N_7560,N_6295,N_6450);
xor U7561 (N_7561,N_6167,N_7078);
or U7562 (N_7562,N_6841,N_6655);
xor U7563 (N_7563,N_6997,N_6677);
xor U7564 (N_7564,N_6154,N_6519);
and U7565 (N_7565,N_6352,N_6024);
and U7566 (N_7566,N_6524,N_7026);
and U7567 (N_7567,N_7179,N_6238);
xor U7568 (N_7568,N_6809,N_7156);
nor U7569 (N_7569,N_6158,N_6266);
or U7570 (N_7570,N_6701,N_6564);
and U7571 (N_7571,N_6288,N_7009);
nand U7572 (N_7572,N_6095,N_6571);
and U7573 (N_7573,N_6917,N_6325);
and U7574 (N_7574,N_6090,N_6900);
and U7575 (N_7575,N_6329,N_6341);
nor U7576 (N_7576,N_6581,N_6106);
nor U7577 (N_7577,N_6638,N_6316);
nand U7578 (N_7578,N_6664,N_6081);
and U7579 (N_7579,N_6044,N_6285);
and U7580 (N_7580,N_6558,N_6856);
and U7581 (N_7581,N_6063,N_6647);
nand U7582 (N_7582,N_6866,N_7115);
xor U7583 (N_7583,N_6690,N_6245);
and U7584 (N_7584,N_7088,N_7116);
or U7585 (N_7585,N_6833,N_6727);
xnor U7586 (N_7586,N_6184,N_6879);
xor U7587 (N_7587,N_6343,N_7023);
nor U7588 (N_7588,N_6215,N_6241);
xnor U7589 (N_7589,N_6576,N_6785);
nor U7590 (N_7590,N_6335,N_6381);
nor U7591 (N_7591,N_6694,N_6379);
nand U7592 (N_7592,N_7149,N_6181);
nand U7593 (N_7593,N_6540,N_6229);
nand U7594 (N_7594,N_7069,N_6687);
xnor U7595 (N_7595,N_6447,N_6013);
nor U7596 (N_7596,N_6482,N_6794);
or U7597 (N_7597,N_6992,N_6415);
xor U7598 (N_7598,N_6904,N_6621);
and U7599 (N_7599,N_6445,N_6893);
nand U7600 (N_7600,N_6554,N_6197);
xor U7601 (N_7601,N_6553,N_6783);
nand U7602 (N_7602,N_6186,N_6046);
nand U7603 (N_7603,N_6679,N_6983);
nand U7604 (N_7604,N_6183,N_6639);
nand U7605 (N_7605,N_6403,N_6253);
nand U7606 (N_7606,N_6425,N_6836);
and U7607 (N_7607,N_6431,N_6462);
nor U7608 (N_7608,N_7101,N_6657);
xnor U7609 (N_7609,N_6416,N_7161);
nor U7610 (N_7610,N_7169,N_6844);
nor U7611 (N_7611,N_6635,N_6846);
and U7612 (N_7612,N_6526,N_6162);
nor U7613 (N_7613,N_6105,N_6523);
and U7614 (N_7614,N_6409,N_6863);
nand U7615 (N_7615,N_6103,N_6790);
xor U7616 (N_7616,N_6353,N_6843);
nor U7617 (N_7617,N_7038,N_6611);
nand U7618 (N_7618,N_6342,N_6437);
or U7619 (N_7619,N_7051,N_6419);
nand U7620 (N_7620,N_6848,N_6235);
nor U7621 (N_7621,N_7048,N_6837);
nor U7622 (N_7622,N_6389,N_6702);
xnor U7623 (N_7623,N_6260,N_6289);
nor U7624 (N_7624,N_6525,N_6153);
or U7625 (N_7625,N_6191,N_6537);
xnor U7626 (N_7626,N_6487,N_6209);
or U7627 (N_7627,N_7047,N_7072);
or U7628 (N_7628,N_6311,N_7139);
xor U7629 (N_7629,N_6413,N_6232);
or U7630 (N_7630,N_6909,N_6216);
xor U7631 (N_7631,N_6284,N_6426);
xnor U7632 (N_7632,N_6796,N_7194);
or U7633 (N_7633,N_6700,N_6269);
nand U7634 (N_7634,N_6961,N_6481);
xnor U7635 (N_7635,N_6070,N_6157);
or U7636 (N_7636,N_6137,N_6804);
nand U7637 (N_7637,N_6498,N_6977);
and U7638 (N_7638,N_6043,N_6175);
and U7639 (N_7639,N_6078,N_6286);
xor U7640 (N_7640,N_6927,N_6870);
nor U7641 (N_7641,N_6624,N_6736);
xnor U7642 (N_7642,N_6091,N_7099);
nand U7643 (N_7643,N_6654,N_6627);
nor U7644 (N_7644,N_6618,N_6612);
or U7645 (N_7645,N_6826,N_6582);
xnor U7646 (N_7646,N_6130,N_6745);
xor U7647 (N_7647,N_7132,N_6164);
nor U7648 (N_7648,N_6906,N_6813);
and U7649 (N_7649,N_6224,N_6185);
nor U7650 (N_7650,N_6479,N_6743);
and U7651 (N_7651,N_6617,N_6765);
nor U7652 (N_7652,N_6511,N_7019);
or U7653 (N_7653,N_6305,N_6484);
nand U7654 (N_7654,N_6812,N_6174);
xor U7655 (N_7655,N_7181,N_6196);
and U7656 (N_7656,N_7159,N_6355);
xor U7657 (N_7657,N_6594,N_6506);
nor U7658 (N_7658,N_6972,N_6739);
xor U7659 (N_7659,N_6940,N_6974);
xor U7660 (N_7660,N_6460,N_6817);
and U7661 (N_7661,N_6792,N_7011);
xor U7662 (N_7662,N_6784,N_6294);
nor U7663 (N_7663,N_6663,N_7093);
nand U7664 (N_7664,N_6251,N_6455);
nand U7665 (N_7665,N_6645,N_6138);
nand U7666 (N_7666,N_7150,N_6884);
and U7667 (N_7667,N_7015,N_6886);
and U7668 (N_7668,N_6793,N_6931);
nor U7669 (N_7669,N_6363,N_6318);
and U7670 (N_7670,N_6697,N_7008);
nand U7671 (N_7671,N_6975,N_6161);
or U7672 (N_7672,N_7113,N_7044);
nand U7673 (N_7673,N_6309,N_7089);
xnor U7674 (N_7674,N_6212,N_6127);
or U7675 (N_7675,N_6507,N_6547);
and U7676 (N_7676,N_6370,N_6047);
xnor U7677 (N_7677,N_6148,N_6234);
or U7678 (N_7678,N_7168,N_6129);
xor U7679 (N_7679,N_6587,N_6710);
and U7680 (N_7680,N_6054,N_6080);
nand U7681 (N_7681,N_6383,N_6685);
and U7682 (N_7682,N_7096,N_6087);
or U7683 (N_7683,N_6766,N_6598);
nand U7684 (N_7684,N_7057,N_6995);
nand U7685 (N_7685,N_6699,N_6962);
nor U7686 (N_7686,N_6764,N_6777);
and U7687 (N_7687,N_6675,N_6776);
xnor U7688 (N_7688,N_6907,N_6508);
nand U7689 (N_7689,N_6223,N_6401);
xnor U7690 (N_7690,N_6467,N_6693);
and U7691 (N_7691,N_6868,N_6121);
nand U7692 (N_7692,N_7127,N_6541);
and U7693 (N_7693,N_6065,N_7063);
or U7694 (N_7694,N_6471,N_6720);
or U7695 (N_7695,N_7192,N_6748);
xor U7696 (N_7696,N_7135,N_6357);
and U7697 (N_7697,N_7035,N_6830);
nor U7698 (N_7698,N_7003,N_6165);
nand U7699 (N_7699,N_7162,N_6126);
and U7700 (N_7700,N_6842,N_6451);
xor U7701 (N_7701,N_6504,N_6513);
and U7702 (N_7702,N_6602,N_6911);
and U7703 (N_7703,N_6192,N_6599);
and U7704 (N_7704,N_6781,N_6001);
or U7705 (N_7705,N_6530,N_6334);
nand U7706 (N_7706,N_6290,N_6608);
nor U7707 (N_7707,N_7126,N_6020);
xnor U7708 (N_7708,N_6671,N_6775);
xor U7709 (N_7709,N_6271,N_6112);
nor U7710 (N_7710,N_7138,N_6083);
nor U7711 (N_7711,N_6478,N_6520);
and U7712 (N_7712,N_6505,N_7002);
nand U7713 (N_7713,N_6936,N_6850);
xnor U7714 (N_7714,N_6189,N_6514);
nand U7715 (N_7715,N_6473,N_7095);
xor U7716 (N_7716,N_7024,N_6586);
xor U7717 (N_7717,N_6926,N_6651);
nand U7718 (N_7718,N_6360,N_6058);
nand U7719 (N_7719,N_6713,N_6396);
and U7720 (N_7720,N_6412,N_7028);
and U7721 (N_7721,N_6845,N_6125);
nand U7722 (N_7722,N_6819,N_7147);
nand U7723 (N_7723,N_6980,N_6089);
or U7724 (N_7724,N_6752,N_6082);
nor U7725 (N_7725,N_6114,N_6773);
nor U7726 (N_7726,N_6438,N_7163);
nand U7727 (N_7727,N_7004,N_6469);
or U7728 (N_7728,N_6696,N_6219);
nor U7729 (N_7729,N_6778,N_6208);
xnor U7730 (N_7730,N_6029,N_6085);
or U7731 (N_7731,N_6084,N_7158);
xor U7732 (N_7732,N_6002,N_7131);
or U7733 (N_7733,N_6050,N_6712);
xnor U7734 (N_7734,N_6559,N_7173);
or U7735 (N_7735,N_6152,N_6815);
nor U7736 (N_7736,N_6056,N_6737);
or U7737 (N_7737,N_6293,N_6615);
or U7738 (N_7738,N_6015,N_6380);
nor U7739 (N_7739,N_6730,N_7007);
or U7740 (N_7740,N_6924,N_6732);
and U7741 (N_7741,N_6021,N_6045);
xor U7742 (N_7742,N_6466,N_7010);
and U7743 (N_7743,N_6110,N_6388);
or U7744 (N_7744,N_6518,N_6376);
nand U7745 (N_7745,N_6250,N_6278);
nor U7746 (N_7746,N_6428,N_6890);
or U7747 (N_7747,N_6569,N_6772);
nand U7748 (N_7748,N_7042,N_6818);
nor U7749 (N_7749,N_6676,N_6440);
or U7750 (N_7750,N_6279,N_6283);
nand U7751 (N_7751,N_6097,N_7119);
and U7752 (N_7752,N_6898,N_7187);
and U7753 (N_7753,N_6247,N_6688);
and U7754 (N_7754,N_6521,N_7128);
xnor U7755 (N_7755,N_6534,N_6650);
and U7756 (N_7756,N_6955,N_6619);
xor U7757 (N_7757,N_7143,N_6028);
xor U7758 (N_7758,N_6069,N_6385);
or U7759 (N_7759,N_6340,N_6539);
and U7760 (N_7760,N_6346,N_6568);
xnor U7761 (N_7761,N_6444,N_6580);
nor U7762 (N_7762,N_6729,N_6336);
xor U7763 (N_7763,N_6354,N_6892);
nor U7764 (N_7764,N_6536,N_6807);
or U7765 (N_7765,N_6976,N_6390);
nor U7766 (N_7766,N_6922,N_6723);
nand U7767 (N_7767,N_7070,N_7184);
or U7768 (N_7768,N_6996,N_7049);
xnor U7769 (N_7769,N_6896,N_6529);
nor U7770 (N_7770,N_7110,N_6073);
and U7771 (N_7771,N_6312,N_6735);
nor U7772 (N_7772,N_6715,N_7084);
and U7773 (N_7773,N_6371,N_6811);
xnor U7774 (N_7774,N_6399,N_6658);
and U7775 (N_7775,N_7106,N_6094);
nor U7776 (N_7776,N_6527,N_6458);
and U7777 (N_7777,N_7183,N_6669);
or U7778 (N_7778,N_6719,N_6798);
and U7779 (N_7779,N_6733,N_6607);
nand U7780 (N_7780,N_6616,N_6595);
xnor U7781 (N_7781,N_6750,N_6802);
xnor U7782 (N_7782,N_6356,N_6692);
and U7783 (N_7783,N_6628,N_7080);
and U7784 (N_7784,N_6894,N_7152);
or U7785 (N_7785,N_6350,N_6243);
nand U7786 (N_7786,N_6620,N_6686);
or U7787 (N_7787,N_7196,N_7079);
or U7788 (N_7788,N_6146,N_6134);
nand U7789 (N_7789,N_6722,N_6497);
nor U7790 (N_7790,N_6194,N_6832);
nor U7791 (N_7791,N_6122,N_6417);
and U7792 (N_7792,N_7157,N_6963);
xnor U7793 (N_7793,N_6382,N_6714);
nor U7794 (N_7794,N_6928,N_6435);
nand U7795 (N_7795,N_6939,N_6859);
or U7796 (N_7796,N_6488,N_6132);
and U7797 (N_7797,N_7189,N_6990);
nor U7798 (N_7798,N_6171,N_6575);
nand U7799 (N_7799,N_6596,N_6172);
or U7800 (N_7800,N_6862,N_6791);
and U7801 (N_7801,N_6275,N_7088);
xor U7802 (N_7802,N_7051,N_6795);
and U7803 (N_7803,N_6650,N_6508);
xnor U7804 (N_7804,N_6372,N_6867);
xor U7805 (N_7805,N_6830,N_6604);
and U7806 (N_7806,N_6727,N_6586);
nor U7807 (N_7807,N_6388,N_6202);
or U7808 (N_7808,N_7187,N_6347);
and U7809 (N_7809,N_6544,N_6826);
and U7810 (N_7810,N_6997,N_6465);
and U7811 (N_7811,N_6147,N_6326);
and U7812 (N_7812,N_6795,N_6804);
nor U7813 (N_7813,N_7194,N_6080);
and U7814 (N_7814,N_6556,N_7053);
nand U7815 (N_7815,N_6697,N_6690);
or U7816 (N_7816,N_6897,N_7110);
or U7817 (N_7817,N_6864,N_6967);
nand U7818 (N_7818,N_6538,N_6974);
xnor U7819 (N_7819,N_6652,N_7134);
and U7820 (N_7820,N_6657,N_6824);
xor U7821 (N_7821,N_6114,N_6590);
nand U7822 (N_7822,N_6192,N_6835);
nand U7823 (N_7823,N_7067,N_6997);
nor U7824 (N_7824,N_6750,N_7120);
nand U7825 (N_7825,N_7145,N_7150);
nand U7826 (N_7826,N_6916,N_7154);
nand U7827 (N_7827,N_6867,N_6254);
and U7828 (N_7828,N_6064,N_6018);
or U7829 (N_7829,N_6728,N_6414);
or U7830 (N_7830,N_6211,N_6229);
nor U7831 (N_7831,N_6710,N_7103);
xnor U7832 (N_7832,N_7061,N_6456);
xor U7833 (N_7833,N_6360,N_6137);
nand U7834 (N_7834,N_6266,N_6150);
and U7835 (N_7835,N_6070,N_6063);
nor U7836 (N_7836,N_6007,N_6654);
xnor U7837 (N_7837,N_6842,N_6042);
nor U7838 (N_7838,N_7008,N_6986);
and U7839 (N_7839,N_6788,N_7099);
nand U7840 (N_7840,N_6000,N_6544);
and U7841 (N_7841,N_7129,N_6778);
xnor U7842 (N_7842,N_6993,N_6172);
xor U7843 (N_7843,N_7041,N_7133);
and U7844 (N_7844,N_7194,N_6487);
and U7845 (N_7845,N_7138,N_6984);
nor U7846 (N_7846,N_6657,N_6036);
xnor U7847 (N_7847,N_6241,N_6316);
and U7848 (N_7848,N_6625,N_7077);
xnor U7849 (N_7849,N_6136,N_6975);
xor U7850 (N_7850,N_6976,N_6898);
and U7851 (N_7851,N_6962,N_7147);
nand U7852 (N_7852,N_6591,N_7139);
and U7853 (N_7853,N_6910,N_6033);
or U7854 (N_7854,N_6391,N_6807);
nand U7855 (N_7855,N_6720,N_6245);
nand U7856 (N_7856,N_7117,N_6161);
and U7857 (N_7857,N_6750,N_6556);
xor U7858 (N_7858,N_6339,N_6814);
nor U7859 (N_7859,N_6989,N_7177);
nor U7860 (N_7860,N_6485,N_6101);
and U7861 (N_7861,N_6244,N_7034);
or U7862 (N_7862,N_7196,N_6998);
nand U7863 (N_7863,N_6021,N_6290);
and U7864 (N_7864,N_7081,N_7021);
xor U7865 (N_7865,N_6488,N_6593);
and U7866 (N_7866,N_6555,N_6156);
xnor U7867 (N_7867,N_7100,N_6491);
xnor U7868 (N_7868,N_6677,N_6839);
nand U7869 (N_7869,N_6039,N_6596);
or U7870 (N_7870,N_7055,N_6609);
nand U7871 (N_7871,N_6919,N_6326);
nor U7872 (N_7872,N_7145,N_6172);
xnor U7873 (N_7873,N_6392,N_6518);
nand U7874 (N_7874,N_6875,N_6210);
nor U7875 (N_7875,N_6807,N_6162);
and U7876 (N_7876,N_6703,N_6038);
or U7877 (N_7877,N_6200,N_6247);
nor U7878 (N_7878,N_7027,N_6524);
and U7879 (N_7879,N_6055,N_6149);
and U7880 (N_7880,N_6768,N_6248);
xnor U7881 (N_7881,N_7180,N_6980);
nor U7882 (N_7882,N_6926,N_6326);
or U7883 (N_7883,N_6226,N_6875);
or U7884 (N_7884,N_6793,N_6597);
and U7885 (N_7885,N_7063,N_7053);
nor U7886 (N_7886,N_6452,N_6921);
and U7887 (N_7887,N_7103,N_7125);
or U7888 (N_7888,N_7061,N_6516);
nand U7889 (N_7889,N_7048,N_6191);
or U7890 (N_7890,N_6660,N_6801);
nor U7891 (N_7891,N_6883,N_6270);
xor U7892 (N_7892,N_7099,N_6519);
or U7893 (N_7893,N_6049,N_6953);
and U7894 (N_7894,N_6568,N_6444);
xor U7895 (N_7895,N_6851,N_6258);
xnor U7896 (N_7896,N_6267,N_6456);
nor U7897 (N_7897,N_6639,N_6238);
nor U7898 (N_7898,N_7185,N_6380);
xnor U7899 (N_7899,N_6887,N_6780);
nor U7900 (N_7900,N_6899,N_6205);
or U7901 (N_7901,N_6702,N_6295);
xor U7902 (N_7902,N_6097,N_6601);
and U7903 (N_7903,N_6922,N_6061);
xor U7904 (N_7904,N_6071,N_6409);
xor U7905 (N_7905,N_6266,N_6157);
nand U7906 (N_7906,N_6155,N_6597);
xor U7907 (N_7907,N_6106,N_6509);
nand U7908 (N_7908,N_6086,N_6656);
nor U7909 (N_7909,N_6374,N_7091);
nor U7910 (N_7910,N_7060,N_6114);
and U7911 (N_7911,N_6711,N_6780);
nand U7912 (N_7912,N_6322,N_6816);
nand U7913 (N_7913,N_6719,N_6555);
nor U7914 (N_7914,N_6990,N_6739);
and U7915 (N_7915,N_6114,N_6291);
and U7916 (N_7916,N_6022,N_6299);
xnor U7917 (N_7917,N_6353,N_7158);
or U7918 (N_7918,N_6218,N_6933);
xnor U7919 (N_7919,N_7102,N_6910);
and U7920 (N_7920,N_7184,N_6234);
nor U7921 (N_7921,N_6336,N_7127);
and U7922 (N_7922,N_7026,N_7148);
nor U7923 (N_7923,N_6457,N_6941);
or U7924 (N_7924,N_6109,N_6635);
and U7925 (N_7925,N_6862,N_6216);
and U7926 (N_7926,N_6542,N_6368);
and U7927 (N_7927,N_6126,N_6116);
nand U7928 (N_7928,N_7047,N_6466);
and U7929 (N_7929,N_6058,N_7119);
xnor U7930 (N_7930,N_6902,N_6265);
and U7931 (N_7931,N_6319,N_6924);
and U7932 (N_7932,N_6434,N_6435);
nand U7933 (N_7933,N_6326,N_6548);
nand U7934 (N_7934,N_6182,N_7143);
nand U7935 (N_7935,N_7070,N_6915);
or U7936 (N_7936,N_6008,N_6755);
xnor U7937 (N_7937,N_6940,N_6825);
and U7938 (N_7938,N_7163,N_6877);
or U7939 (N_7939,N_6454,N_6345);
nor U7940 (N_7940,N_6181,N_6585);
xor U7941 (N_7941,N_6884,N_6697);
nor U7942 (N_7942,N_6438,N_7197);
or U7943 (N_7943,N_6117,N_7021);
xnor U7944 (N_7944,N_6365,N_6223);
or U7945 (N_7945,N_7141,N_6087);
or U7946 (N_7946,N_6890,N_6536);
nor U7947 (N_7947,N_6649,N_7119);
nand U7948 (N_7948,N_6118,N_7058);
nand U7949 (N_7949,N_6171,N_6046);
or U7950 (N_7950,N_7166,N_6578);
xor U7951 (N_7951,N_6671,N_6898);
nand U7952 (N_7952,N_6542,N_7123);
nand U7953 (N_7953,N_6171,N_6314);
nor U7954 (N_7954,N_6292,N_6246);
nand U7955 (N_7955,N_7118,N_6263);
nand U7956 (N_7956,N_7030,N_6616);
xnor U7957 (N_7957,N_6571,N_6180);
nor U7958 (N_7958,N_6626,N_6554);
and U7959 (N_7959,N_6585,N_6618);
or U7960 (N_7960,N_7126,N_6361);
xor U7961 (N_7961,N_6451,N_6361);
and U7962 (N_7962,N_6951,N_6033);
xor U7963 (N_7963,N_6074,N_6446);
or U7964 (N_7964,N_6292,N_6839);
xnor U7965 (N_7965,N_6015,N_6381);
xnor U7966 (N_7966,N_6568,N_6321);
and U7967 (N_7967,N_6586,N_6866);
nand U7968 (N_7968,N_6703,N_6557);
nand U7969 (N_7969,N_6708,N_6224);
xnor U7970 (N_7970,N_6689,N_6835);
or U7971 (N_7971,N_6484,N_6502);
nand U7972 (N_7972,N_7174,N_6261);
nand U7973 (N_7973,N_6756,N_6349);
or U7974 (N_7974,N_6891,N_6943);
nand U7975 (N_7975,N_6483,N_6390);
or U7976 (N_7976,N_7020,N_6256);
nor U7977 (N_7977,N_6951,N_7130);
xor U7978 (N_7978,N_6380,N_6412);
nand U7979 (N_7979,N_6182,N_6353);
and U7980 (N_7980,N_6466,N_6100);
nand U7981 (N_7981,N_6873,N_6920);
xor U7982 (N_7982,N_6587,N_6843);
nand U7983 (N_7983,N_6514,N_6091);
xor U7984 (N_7984,N_6344,N_6007);
and U7985 (N_7985,N_7059,N_6482);
nor U7986 (N_7986,N_6959,N_6523);
and U7987 (N_7987,N_6023,N_6502);
or U7988 (N_7988,N_6221,N_6140);
or U7989 (N_7989,N_7130,N_6300);
nor U7990 (N_7990,N_6458,N_6030);
or U7991 (N_7991,N_6422,N_6467);
nor U7992 (N_7992,N_6199,N_6859);
and U7993 (N_7993,N_6438,N_6820);
and U7994 (N_7994,N_6385,N_7030);
and U7995 (N_7995,N_6452,N_6511);
nand U7996 (N_7996,N_6776,N_6347);
and U7997 (N_7997,N_6086,N_6083);
nor U7998 (N_7998,N_6877,N_6445);
or U7999 (N_7999,N_6299,N_6111);
nand U8000 (N_8000,N_6407,N_7018);
nor U8001 (N_8001,N_6468,N_6940);
nor U8002 (N_8002,N_6977,N_6731);
nand U8003 (N_8003,N_6058,N_6199);
or U8004 (N_8004,N_7173,N_6328);
or U8005 (N_8005,N_6916,N_6363);
and U8006 (N_8006,N_6536,N_6788);
xnor U8007 (N_8007,N_6871,N_6316);
xnor U8008 (N_8008,N_6366,N_6493);
and U8009 (N_8009,N_6805,N_6997);
and U8010 (N_8010,N_6088,N_6445);
or U8011 (N_8011,N_6488,N_6469);
nor U8012 (N_8012,N_6604,N_6074);
and U8013 (N_8013,N_7119,N_6315);
nand U8014 (N_8014,N_7040,N_6913);
or U8015 (N_8015,N_6873,N_7026);
and U8016 (N_8016,N_7144,N_6187);
xor U8017 (N_8017,N_6591,N_6935);
and U8018 (N_8018,N_6921,N_6245);
nand U8019 (N_8019,N_6843,N_6578);
nand U8020 (N_8020,N_6676,N_7011);
or U8021 (N_8021,N_6066,N_6635);
and U8022 (N_8022,N_6325,N_6802);
xor U8023 (N_8023,N_6896,N_6394);
xnor U8024 (N_8024,N_6667,N_6124);
xor U8025 (N_8025,N_6436,N_6738);
and U8026 (N_8026,N_6399,N_6837);
and U8027 (N_8027,N_6094,N_6711);
or U8028 (N_8028,N_6348,N_6400);
nand U8029 (N_8029,N_6775,N_6886);
and U8030 (N_8030,N_6660,N_6340);
nor U8031 (N_8031,N_6308,N_7055);
nor U8032 (N_8032,N_6503,N_6712);
and U8033 (N_8033,N_6266,N_6501);
xor U8034 (N_8034,N_6151,N_6263);
nand U8035 (N_8035,N_6549,N_6915);
or U8036 (N_8036,N_6946,N_6323);
and U8037 (N_8037,N_6488,N_7093);
nor U8038 (N_8038,N_6361,N_6307);
xor U8039 (N_8039,N_6826,N_6624);
xnor U8040 (N_8040,N_6322,N_6774);
nand U8041 (N_8041,N_6490,N_6088);
xnor U8042 (N_8042,N_6127,N_7192);
xor U8043 (N_8043,N_6306,N_6420);
nor U8044 (N_8044,N_6464,N_6860);
or U8045 (N_8045,N_6688,N_6270);
or U8046 (N_8046,N_6551,N_6528);
nor U8047 (N_8047,N_6077,N_6369);
xnor U8048 (N_8048,N_7057,N_6966);
or U8049 (N_8049,N_6192,N_6123);
and U8050 (N_8050,N_6353,N_6199);
and U8051 (N_8051,N_6490,N_6136);
nor U8052 (N_8052,N_6288,N_6936);
nand U8053 (N_8053,N_6417,N_6197);
nand U8054 (N_8054,N_6469,N_6565);
or U8055 (N_8055,N_6771,N_6760);
xor U8056 (N_8056,N_6880,N_6312);
and U8057 (N_8057,N_6497,N_7076);
nor U8058 (N_8058,N_6990,N_7009);
xor U8059 (N_8059,N_6575,N_6503);
xnor U8060 (N_8060,N_6876,N_6594);
xor U8061 (N_8061,N_6717,N_6554);
nor U8062 (N_8062,N_7073,N_6956);
xnor U8063 (N_8063,N_6074,N_6974);
nor U8064 (N_8064,N_7178,N_6688);
nand U8065 (N_8065,N_6239,N_6434);
xnor U8066 (N_8066,N_7081,N_6294);
or U8067 (N_8067,N_6581,N_7196);
xnor U8068 (N_8068,N_7124,N_6655);
xnor U8069 (N_8069,N_7037,N_7064);
and U8070 (N_8070,N_6651,N_6047);
xor U8071 (N_8071,N_6237,N_6797);
nand U8072 (N_8072,N_7093,N_6768);
nand U8073 (N_8073,N_6599,N_6296);
xnor U8074 (N_8074,N_6766,N_6299);
nand U8075 (N_8075,N_6458,N_6195);
or U8076 (N_8076,N_6315,N_6181);
nand U8077 (N_8077,N_6838,N_6320);
or U8078 (N_8078,N_6288,N_6534);
or U8079 (N_8079,N_7032,N_7191);
xnor U8080 (N_8080,N_6774,N_6236);
nand U8081 (N_8081,N_6893,N_7005);
nor U8082 (N_8082,N_6368,N_6846);
nor U8083 (N_8083,N_6354,N_7050);
nand U8084 (N_8084,N_7008,N_6357);
nand U8085 (N_8085,N_6320,N_6606);
or U8086 (N_8086,N_6779,N_7070);
nor U8087 (N_8087,N_6411,N_6122);
xnor U8088 (N_8088,N_6594,N_6907);
nand U8089 (N_8089,N_7168,N_7143);
nor U8090 (N_8090,N_6565,N_6826);
xor U8091 (N_8091,N_6436,N_6170);
or U8092 (N_8092,N_6011,N_6707);
and U8093 (N_8093,N_6032,N_6238);
and U8094 (N_8094,N_6567,N_7181);
or U8095 (N_8095,N_6464,N_6036);
and U8096 (N_8096,N_6978,N_6244);
nor U8097 (N_8097,N_6376,N_6764);
or U8098 (N_8098,N_6942,N_7173);
or U8099 (N_8099,N_6178,N_6851);
nor U8100 (N_8100,N_6644,N_6933);
nand U8101 (N_8101,N_6224,N_6324);
and U8102 (N_8102,N_7163,N_6042);
and U8103 (N_8103,N_6385,N_7083);
nand U8104 (N_8104,N_6232,N_6241);
or U8105 (N_8105,N_6625,N_6753);
or U8106 (N_8106,N_6690,N_6572);
or U8107 (N_8107,N_6185,N_6295);
nor U8108 (N_8108,N_6029,N_6772);
nor U8109 (N_8109,N_6065,N_6108);
and U8110 (N_8110,N_7027,N_6326);
or U8111 (N_8111,N_6793,N_6128);
nor U8112 (N_8112,N_6877,N_6270);
or U8113 (N_8113,N_6861,N_6241);
or U8114 (N_8114,N_6196,N_6122);
and U8115 (N_8115,N_6348,N_6795);
nand U8116 (N_8116,N_6285,N_6180);
nor U8117 (N_8117,N_7048,N_6404);
xnor U8118 (N_8118,N_6921,N_7174);
or U8119 (N_8119,N_6814,N_6377);
nand U8120 (N_8120,N_6608,N_6001);
nor U8121 (N_8121,N_6951,N_6563);
or U8122 (N_8122,N_6771,N_7155);
nand U8123 (N_8123,N_6207,N_6030);
or U8124 (N_8124,N_6942,N_6288);
xnor U8125 (N_8125,N_6793,N_6101);
xor U8126 (N_8126,N_6782,N_7145);
nand U8127 (N_8127,N_6960,N_6702);
xor U8128 (N_8128,N_6438,N_6406);
and U8129 (N_8129,N_6381,N_6767);
nor U8130 (N_8130,N_6465,N_6462);
nor U8131 (N_8131,N_6952,N_6044);
xnor U8132 (N_8132,N_6204,N_6072);
nor U8133 (N_8133,N_6243,N_6664);
or U8134 (N_8134,N_6624,N_6035);
nor U8135 (N_8135,N_6100,N_7031);
or U8136 (N_8136,N_6258,N_6344);
xor U8137 (N_8137,N_6182,N_6137);
nand U8138 (N_8138,N_7134,N_6681);
nand U8139 (N_8139,N_6505,N_7064);
xor U8140 (N_8140,N_6929,N_7088);
nand U8141 (N_8141,N_7087,N_6809);
xnor U8142 (N_8142,N_6127,N_6311);
nor U8143 (N_8143,N_6862,N_6411);
nand U8144 (N_8144,N_6411,N_6288);
or U8145 (N_8145,N_7055,N_6404);
nand U8146 (N_8146,N_7075,N_6015);
xor U8147 (N_8147,N_7080,N_6836);
nor U8148 (N_8148,N_6700,N_6106);
xor U8149 (N_8149,N_7173,N_6976);
nor U8150 (N_8150,N_6862,N_6945);
and U8151 (N_8151,N_6703,N_6309);
or U8152 (N_8152,N_6835,N_6932);
nor U8153 (N_8153,N_6085,N_7178);
xnor U8154 (N_8154,N_6143,N_6856);
nand U8155 (N_8155,N_6898,N_6436);
and U8156 (N_8156,N_6838,N_6243);
or U8157 (N_8157,N_6443,N_6692);
or U8158 (N_8158,N_6049,N_6372);
and U8159 (N_8159,N_6091,N_6079);
xor U8160 (N_8160,N_7117,N_6259);
xor U8161 (N_8161,N_6585,N_6683);
nor U8162 (N_8162,N_6766,N_7136);
nor U8163 (N_8163,N_6540,N_6096);
nor U8164 (N_8164,N_6484,N_6652);
and U8165 (N_8165,N_7035,N_6959);
and U8166 (N_8166,N_6515,N_6465);
or U8167 (N_8167,N_6349,N_6644);
nand U8168 (N_8168,N_6326,N_6009);
nor U8169 (N_8169,N_6580,N_6246);
or U8170 (N_8170,N_6384,N_6778);
nor U8171 (N_8171,N_6239,N_7164);
xor U8172 (N_8172,N_6336,N_6526);
xor U8173 (N_8173,N_7056,N_6936);
nor U8174 (N_8174,N_6897,N_6286);
nand U8175 (N_8175,N_6924,N_7025);
or U8176 (N_8176,N_6406,N_6050);
xnor U8177 (N_8177,N_7019,N_7072);
or U8178 (N_8178,N_6424,N_6051);
nor U8179 (N_8179,N_6316,N_6521);
or U8180 (N_8180,N_6999,N_6533);
nand U8181 (N_8181,N_7085,N_6245);
and U8182 (N_8182,N_6012,N_6009);
nor U8183 (N_8183,N_6697,N_6520);
and U8184 (N_8184,N_6390,N_6123);
xnor U8185 (N_8185,N_6713,N_6405);
xor U8186 (N_8186,N_6580,N_6680);
nor U8187 (N_8187,N_7170,N_6098);
and U8188 (N_8188,N_6389,N_6683);
or U8189 (N_8189,N_6775,N_6776);
nor U8190 (N_8190,N_6573,N_6625);
or U8191 (N_8191,N_6240,N_6737);
and U8192 (N_8192,N_6677,N_6693);
or U8193 (N_8193,N_6041,N_6341);
xor U8194 (N_8194,N_6226,N_6499);
xor U8195 (N_8195,N_6669,N_6778);
or U8196 (N_8196,N_6994,N_6070);
xnor U8197 (N_8197,N_7180,N_6128);
nand U8198 (N_8198,N_6169,N_6491);
nor U8199 (N_8199,N_6129,N_7011);
nor U8200 (N_8200,N_6653,N_6801);
nor U8201 (N_8201,N_6207,N_6368);
and U8202 (N_8202,N_6111,N_6531);
or U8203 (N_8203,N_6824,N_6910);
nor U8204 (N_8204,N_6296,N_6309);
and U8205 (N_8205,N_6084,N_7168);
or U8206 (N_8206,N_6745,N_7088);
xor U8207 (N_8207,N_6157,N_6770);
nand U8208 (N_8208,N_6310,N_6490);
and U8209 (N_8209,N_6894,N_6001);
and U8210 (N_8210,N_6981,N_6476);
xor U8211 (N_8211,N_6785,N_6374);
nor U8212 (N_8212,N_6232,N_7099);
nand U8213 (N_8213,N_6509,N_6287);
nor U8214 (N_8214,N_6877,N_7068);
or U8215 (N_8215,N_6496,N_6965);
and U8216 (N_8216,N_6932,N_6217);
nor U8217 (N_8217,N_6283,N_6030);
nand U8218 (N_8218,N_7073,N_6733);
xnor U8219 (N_8219,N_6788,N_6046);
xnor U8220 (N_8220,N_7062,N_6385);
nor U8221 (N_8221,N_6733,N_6693);
and U8222 (N_8222,N_6151,N_6376);
or U8223 (N_8223,N_6520,N_6302);
and U8224 (N_8224,N_6844,N_6669);
nor U8225 (N_8225,N_6608,N_7104);
nor U8226 (N_8226,N_6719,N_7065);
xor U8227 (N_8227,N_6635,N_6726);
or U8228 (N_8228,N_6903,N_6890);
and U8229 (N_8229,N_6549,N_6127);
nand U8230 (N_8230,N_6350,N_6463);
and U8231 (N_8231,N_6080,N_6711);
xnor U8232 (N_8232,N_6812,N_6810);
nor U8233 (N_8233,N_6767,N_6123);
and U8234 (N_8234,N_6546,N_6490);
xor U8235 (N_8235,N_6249,N_6118);
nor U8236 (N_8236,N_6483,N_6207);
and U8237 (N_8237,N_6318,N_6137);
nand U8238 (N_8238,N_6095,N_6984);
or U8239 (N_8239,N_6888,N_7084);
and U8240 (N_8240,N_6565,N_6235);
and U8241 (N_8241,N_6030,N_6224);
or U8242 (N_8242,N_6313,N_6483);
and U8243 (N_8243,N_6518,N_6925);
nor U8244 (N_8244,N_7074,N_6803);
nand U8245 (N_8245,N_6378,N_6101);
and U8246 (N_8246,N_6065,N_6781);
and U8247 (N_8247,N_6964,N_6491);
nand U8248 (N_8248,N_6626,N_7020);
and U8249 (N_8249,N_6308,N_6394);
or U8250 (N_8250,N_6154,N_6901);
xnor U8251 (N_8251,N_6781,N_6484);
nand U8252 (N_8252,N_6027,N_7165);
and U8253 (N_8253,N_6302,N_6184);
nand U8254 (N_8254,N_7109,N_6549);
nand U8255 (N_8255,N_6476,N_6466);
or U8256 (N_8256,N_6539,N_6413);
nand U8257 (N_8257,N_6792,N_6756);
nor U8258 (N_8258,N_6137,N_6983);
xnor U8259 (N_8259,N_6634,N_6563);
and U8260 (N_8260,N_6481,N_6690);
nand U8261 (N_8261,N_6454,N_6571);
or U8262 (N_8262,N_6161,N_6140);
xor U8263 (N_8263,N_6476,N_6985);
and U8264 (N_8264,N_6660,N_6276);
xnor U8265 (N_8265,N_6897,N_6888);
or U8266 (N_8266,N_6285,N_6368);
nand U8267 (N_8267,N_6708,N_6661);
or U8268 (N_8268,N_6894,N_7156);
nor U8269 (N_8269,N_6513,N_6313);
nand U8270 (N_8270,N_6828,N_6415);
and U8271 (N_8271,N_6673,N_6595);
or U8272 (N_8272,N_6665,N_6441);
nand U8273 (N_8273,N_7053,N_6401);
nor U8274 (N_8274,N_6475,N_6370);
xor U8275 (N_8275,N_6778,N_6692);
nand U8276 (N_8276,N_6657,N_7128);
and U8277 (N_8277,N_6603,N_7073);
nor U8278 (N_8278,N_6040,N_6297);
or U8279 (N_8279,N_6692,N_6896);
xor U8280 (N_8280,N_6716,N_6758);
and U8281 (N_8281,N_6278,N_6704);
nor U8282 (N_8282,N_6661,N_6743);
nand U8283 (N_8283,N_6074,N_6050);
or U8284 (N_8284,N_6376,N_6339);
and U8285 (N_8285,N_7131,N_6743);
and U8286 (N_8286,N_6336,N_6953);
xnor U8287 (N_8287,N_6529,N_6181);
xnor U8288 (N_8288,N_6532,N_6918);
nor U8289 (N_8289,N_6412,N_7157);
or U8290 (N_8290,N_6187,N_6309);
xnor U8291 (N_8291,N_6417,N_7019);
and U8292 (N_8292,N_6036,N_6556);
nor U8293 (N_8293,N_6846,N_6332);
and U8294 (N_8294,N_6382,N_7103);
nor U8295 (N_8295,N_6806,N_6878);
nand U8296 (N_8296,N_6132,N_6653);
and U8297 (N_8297,N_6148,N_6482);
nor U8298 (N_8298,N_6988,N_7106);
and U8299 (N_8299,N_6035,N_6788);
xnor U8300 (N_8300,N_6768,N_6398);
and U8301 (N_8301,N_6849,N_6936);
nand U8302 (N_8302,N_6389,N_6069);
nor U8303 (N_8303,N_7081,N_6483);
xor U8304 (N_8304,N_6658,N_6560);
xnor U8305 (N_8305,N_6187,N_6797);
or U8306 (N_8306,N_6074,N_6961);
nand U8307 (N_8307,N_7041,N_6891);
xnor U8308 (N_8308,N_6602,N_6921);
and U8309 (N_8309,N_6397,N_6152);
or U8310 (N_8310,N_7014,N_7107);
xnor U8311 (N_8311,N_6279,N_6452);
and U8312 (N_8312,N_6522,N_6929);
nand U8313 (N_8313,N_6716,N_6125);
and U8314 (N_8314,N_6104,N_6677);
nand U8315 (N_8315,N_6200,N_6937);
xnor U8316 (N_8316,N_6346,N_6725);
nand U8317 (N_8317,N_6202,N_6481);
nor U8318 (N_8318,N_6072,N_6451);
nand U8319 (N_8319,N_6967,N_6560);
nor U8320 (N_8320,N_6163,N_6486);
xnor U8321 (N_8321,N_6455,N_6384);
xnor U8322 (N_8322,N_6618,N_7169);
and U8323 (N_8323,N_6339,N_6486);
nand U8324 (N_8324,N_7179,N_6880);
nor U8325 (N_8325,N_6879,N_6372);
xnor U8326 (N_8326,N_6071,N_6313);
nand U8327 (N_8327,N_6731,N_6016);
nand U8328 (N_8328,N_6567,N_6781);
nor U8329 (N_8329,N_6184,N_6824);
nand U8330 (N_8330,N_6835,N_6492);
and U8331 (N_8331,N_6872,N_6302);
or U8332 (N_8332,N_7043,N_7186);
or U8333 (N_8333,N_6493,N_6790);
xnor U8334 (N_8334,N_6375,N_6768);
and U8335 (N_8335,N_6628,N_6884);
or U8336 (N_8336,N_6141,N_6498);
and U8337 (N_8337,N_6480,N_6602);
or U8338 (N_8338,N_6045,N_7008);
xor U8339 (N_8339,N_6019,N_7176);
xnor U8340 (N_8340,N_6505,N_6127);
and U8341 (N_8341,N_6821,N_6580);
xnor U8342 (N_8342,N_6911,N_6343);
nor U8343 (N_8343,N_6013,N_6534);
nand U8344 (N_8344,N_6981,N_6259);
nand U8345 (N_8345,N_6981,N_6386);
nor U8346 (N_8346,N_6064,N_6053);
nand U8347 (N_8347,N_6618,N_6739);
and U8348 (N_8348,N_7062,N_6282);
and U8349 (N_8349,N_6360,N_6271);
or U8350 (N_8350,N_6115,N_6260);
and U8351 (N_8351,N_6972,N_6425);
xnor U8352 (N_8352,N_7030,N_6052);
and U8353 (N_8353,N_7050,N_6062);
nor U8354 (N_8354,N_6637,N_6863);
xnor U8355 (N_8355,N_6642,N_6714);
nand U8356 (N_8356,N_6163,N_6181);
xnor U8357 (N_8357,N_6984,N_7105);
or U8358 (N_8358,N_6864,N_6448);
xor U8359 (N_8359,N_6967,N_6466);
and U8360 (N_8360,N_6206,N_6072);
or U8361 (N_8361,N_6119,N_7014);
nor U8362 (N_8362,N_6372,N_6899);
xnor U8363 (N_8363,N_6881,N_6314);
and U8364 (N_8364,N_6187,N_6120);
or U8365 (N_8365,N_7050,N_6472);
xor U8366 (N_8366,N_6638,N_6259);
and U8367 (N_8367,N_6493,N_6070);
nor U8368 (N_8368,N_6622,N_6113);
nand U8369 (N_8369,N_7185,N_6033);
and U8370 (N_8370,N_7124,N_6276);
or U8371 (N_8371,N_6968,N_6950);
and U8372 (N_8372,N_6404,N_6895);
nand U8373 (N_8373,N_6994,N_6246);
and U8374 (N_8374,N_6752,N_6022);
and U8375 (N_8375,N_6344,N_6284);
xnor U8376 (N_8376,N_6806,N_6957);
nand U8377 (N_8377,N_6701,N_6783);
nor U8378 (N_8378,N_6082,N_7086);
and U8379 (N_8379,N_6953,N_6309);
and U8380 (N_8380,N_6417,N_7067);
or U8381 (N_8381,N_6188,N_6658);
nand U8382 (N_8382,N_6313,N_6216);
or U8383 (N_8383,N_6486,N_6132);
and U8384 (N_8384,N_6926,N_6065);
xnor U8385 (N_8385,N_7159,N_6263);
nor U8386 (N_8386,N_7030,N_6506);
or U8387 (N_8387,N_6075,N_6364);
nand U8388 (N_8388,N_6532,N_6166);
or U8389 (N_8389,N_6010,N_6220);
or U8390 (N_8390,N_6030,N_6045);
nor U8391 (N_8391,N_6720,N_7056);
nand U8392 (N_8392,N_6555,N_6208);
and U8393 (N_8393,N_6975,N_6339);
and U8394 (N_8394,N_7164,N_6447);
or U8395 (N_8395,N_7030,N_6451);
nor U8396 (N_8396,N_6166,N_7081);
or U8397 (N_8397,N_6993,N_6870);
or U8398 (N_8398,N_6481,N_6511);
nor U8399 (N_8399,N_6952,N_6255);
nor U8400 (N_8400,N_7536,N_7974);
or U8401 (N_8401,N_7522,N_7574);
and U8402 (N_8402,N_8301,N_7677);
and U8403 (N_8403,N_7864,N_8378);
and U8404 (N_8404,N_7809,N_8299);
xnor U8405 (N_8405,N_7729,N_8153);
nand U8406 (N_8406,N_8159,N_7822);
nor U8407 (N_8407,N_7706,N_7892);
nand U8408 (N_8408,N_7816,N_7728);
nor U8409 (N_8409,N_7573,N_8147);
xor U8410 (N_8410,N_8317,N_7794);
nand U8411 (N_8411,N_7991,N_7317);
nor U8412 (N_8412,N_7430,N_7683);
or U8413 (N_8413,N_7965,N_7557);
nand U8414 (N_8414,N_7753,N_7339);
and U8415 (N_8415,N_7811,N_8243);
xnor U8416 (N_8416,N_7995,N_8007);
nand U8417 (N_8417,N_7603,N_7987);
nand U8418 (N_8418,N_7602,N_7943);
nor U8419 (N_8419,N_7423,N_7469);
nor U8420 (N_8420,N_8043,N_7748);
xnor U8421 (N_8421,N_8316,N_7321);
nor U8422 (N_8422,N_8157,N_8245);
and U8423 (N_8423,N_7242,N_7951);
xor U8424 (N_8424,N_8025,N_7261);
nand U8425 (N_8425,N_8106,N_7342);
nor U8426 (N_8426,N_7420,N_7688);
xnor U8427 (N_8427,N_7275,N_8031);
or U8428 (N_8428,N_7778,N_7689);
nor U8429 (N_8429,N_7986,N_7674);
xnor U8430 (N_8430,N_7203,N_7896);
and U8431 (N_8431,N_7703,N_7730);
nor U8432 (N_8432,N_7471,N_7801);
nor U8433 (N_8433,N_8366,N_8283);
nor U8434 (N_8434,N_7546,N_7608);
nor U8435 (N_8435,N_8331,N_7666);
nor U8436 (N_8436,N_8224,N_8201);
nor U8437 (N_8437,N_8122,N_7961);
and U8438 (N_8438,N_8078,N_7643);
and U8439 (N_8439,N_7627,N_7717);
nand U8440 (N_8440,N_7597,N_7854);
nand U8441 (N_8441,N_8327,N_8033);
nor U8442 (N_8442,N_7789,N_7806);
or U8443 (N_8443,N_8394,N_7929);
nand U8444 (N_8444,N_7518,N_8362);
nor U8445 (N_8445,N_8399,N_7397);
and U8446 (N_8446,N_8042,N_7247);
or U8447 (N_8447,N_8357,N_7464);
and U8448 (N_8448,N_7997,N_7364);
nand U8449 (N_8449,N_7226,N_7893);
nor U8450 (N_8450,N_7682,N_8053);
or U8451 (N_8451,N_7784,N_8375);
xor U8452 (N_8452,N_8143,N_7950);
or U8453 (N_8453,N_7972,N_7807);
nand U8454 (N_8454,N_7289,N_8087);
xor U8455 (N_8455,N_8238,N_7631);
and U8456 (N_8456,N_8295,N_7785);
nand U8457 (N_8457,N_7447,N_7402);
or U8458 (N_8458,N_8128,N_7322);
or U8459 (N_8459,N_8011,N_8195);
or U8460 (N_8460,N_7381,N_7818);
or U8461 (N_8461,N_7538,N_8352);
or U8462 (N_8462,N_7590,N_7907);
xnor U8463 (N_8463,N_7812,N_7216);
and U8464 (N_8464,N_7567,N_7359);
nor U8465 (N_8465,N_7527,N_7504);
or U8466 (N_8466,N_8109,N_7354);
xor U8467 (N_8467,N_7942,N_8267);
xnor U8468 (N_8468,N_7498,N_7213);
and U8469 (N_8469,N_8185,N_7960);
or U8470 (N_8470,N_7742,N_7551);
nand U8471 (N_8471,N_8155,N_8160);
and U8472 (N_8472,N_7982,N_7416);
or U8473 (N_8473,N_7768,N_7741);
xor U8474 (N_8474,N_7408,N_7422);
nand U8475 (N_8475,N_7790,N_7484);
or U8476 (N_8476,N_8003,N_8223);
nor U8477 (N_8477,N_7714,N_7284);
nor U8478 (N_8478,N_7883,N_8126);
nand U8479 (N_8479,N_7834,N_7312);
xnor U8480 (N_8480,N_7610,N_7502);
or U8481 (N_8481,N_8204,N_7862);
or U8482 (N_8482,N_7744,N_7882);
nor U8483 (N_8483,N_7800,N_7492);
and U8484 (N_8484,N_7468,N_7999);
and U8485 (N_8485,N_7957,N_7466);
nand U8486 (N_8486,N_7707,N_8151);
nand U8487 (N_8487,N_7911,N_7440);
nand U8488 (N_8488,N_7479,N_7959);
nand U8489 (N_8489,N_8354,N_8056);
and U8490 (N_8490,N_7325,N_7556);
nand U8491 (N_8491,N_8311,N_7214);
or U8492 (N_8492,N_7345,N_7539);
nor U8493 (N_8493,N_7413,N_8110);
nor U8494 (N_8494,N_8361,N_7238);
xor U8495 (N_8495,N_8288,N_7251);
and U8496 (N_8496,N_7441,N_8148);
and U8497 (N_8497,N_8373,N_7391);
nand U8498 (N_8498,N_8123,N_7827);
nand U8499 (N_8499,N_7316,N_7537);
or U8500 (N_8500,N_7727,N_7348);
nor U8501 (N_8501,N_7555,N_7825);
nand U8502 (N_8502,N_7710,N_7908);
and U8503 (N_8503,N_7726,N_7563);
and U8504 (N_8504,N_7228,N_7926);
and U8505 (N_8505,N_7411,N_8051);
nand U8506 (N_8506,N_7863,N_8213);
nor U8507 (N_8507,N_7534,N_7850);
xnor U8508 (N_8508,N_7781,N_8014);
xnor U8509 (N_8509,N_8228,N_7398);
nand U8510 (N_8510,N_8175,N_8065);
nor U8511 (N_8511,N_7699,N_7824);
and U8512 (N_8512,N_7234,N_7686);
nand U8513 (N_8513,N_7779,N_7552);
or U8514 (N_8514,N_8141,N_8358);
and U8515 (N_8515,N_7767,N_7799);
and U8516 (N_8516,N_8154,N_7891);
or U8517 (N_8517,N_7382,N_7501);
nor U8518 (N_8518,N_7765,N_8008);
or U8519 (N_8519,N_7980,N_8116);
nand U8520 (N_8520,N_7559,N_7988);
or U8521 (N_8521,N_7685,N_7246);
and U8522 (N_8522,N_8344,N_7692);
nor U8523 (N_8523,N_8231,N_7255);
nor U8524 (N_8524,N_8019,N_7346);
or U8525 (N_8525,N_7736,N_8196);
and U8526 (N_8526,N_7217,N_7334);
or U8527 (N_8527,N_7283,N_8194);
nand U8528 (N_8528,N_8144,N_7287);
and U8529 (N_8529,N_7244,N_8112);
xor U8530 (N_8530,N_7560,N_8114);
nor U8531 (N_8531,N_8265,N_8277);
nand U8532 (N_8532,N_7568,N_8377);
and U8533 (N_8533,N_7528,N_8315);
nand U8534 (N_8534,N_7973,N_7885);
nor U8535 (N_8535,N_8235,N_7503);
nor U8536 (N_8536,N_8297,N_7720);
xnor U8537 (N_8537,N_8009,N_8132);
xor U8538 (N_8538,N_7277,N_7507);
nor U8539 (N_8539,N_7482,N_7525);
nor U8540 (N_8540,N_8115,N_7327);
xor U8541 (N_8541,N_7586,N_7314);
nor U8542 (N_8542,N_8125,N_7587);
and U8543 (N_8543,N_8055,N_7329);
nor U8544 (N_8544,N_7403,N_8232);
and U8545 (N_8545,N_8341,N_8146);
or U8546 (N_8546,N_7656,N_7589);
nor U8547 (N_8547,N_7291,N_7731);
nor U8548 (N_8548,N_8119,N_7426);
nand U8549 (N_8549,N_7324,N_8092);
or U8550 (N_8550,N_7838,N_8161);
nor U8551 (N_8551,N_7265,N_7802);
xor U8552 (N_8552,N_8152,N_7887);
nor U8553 (N_8553,N_7695,N_7837);
xor U8554 (N_8554,N_7696,N_8039);
and U8555 (N_8555,N_7684,N_7598);
or U8556 (N_8556,N_7671,N_7776);
xnor U8557 (N_8557,N_7313,N_7902);
nand U8558 (N_8558,N_7996,N_7924);
and U8559 (N_8559,N_7947,N_8313);
nand U8560 (N_8560,N_8117,N_7296);
nor U8561 (N_8561,N_8212,N_7473);
nand U8562 (N_8562,N_7511,N_7544);
xor U8563 (N_8563,N_7497,N_7338);
and U8564 (N_8564,N_7820,N_7488);
nand U8565 (N_8565,N_7512,N_7712);
nand U8566 (N_8566,N_7739,N_7769);
xor U8567 (N_8567,N_8292,N_8108);
nor U8568 (N_8568,N_7526,N_7495);
or U8569 (N_8569,N_7798,N_8263);
nand U8570 (N_8570,N_7612,N_8398);
or U8571 (N_8571,N_8219,N_7585);
nand U8572 (N_8572,N_7901,N_8364);
nor U8573 (N_8573,N_8207,N_7480);
or U8574 (N_8574,N_7515,N_8272);
xnor U8575 (N_8575,N_7481,N_8047);
or U8576 (N_8576,N_7318,N_7897);
and U8577 (N_8577,N_7212,N_7379);
nand U8578 (N_8578,N_7766,N_7953);
nor U8579 (N_8579,N_7917,N_7904);
or U8580 (N_8580,N_8239,N_7207);
nand U8581 (N_8581,N_7675,N_7826);
and U8582 (N_8582,N_7638,N_7489);
nand U8583 (N_8583,N_7687,N_7762);
nor U8584 (N_8584,N_8333,N_7723);
xnor U8585 (N_8585,N_7757,N_7583);
or U8586 (N_8586,N_8329,N_8081);
nor U8587 (N_8587,N_8189,N_8356);
nor U8588 (N_8588,N_7575,N_8391);
and U8589 (N_8589,N_8323,N_8396);
and U8590 (N_8590,N_8050,N_7442);
or U8591 (N_8591,N_8041,N_8200);
or U8592 (N_8592,N_7465,N_7428);
nor U8593 (N_8593,N_7934,N_7360);
nand U8594 (N_8594,N_7852,N_7549);
nor U8595 (N_8595,N_8100,N_7380);
and U8596 (N_8596,N_8321,N_7400);
nor U8597 (N_8597,N_7830,N_7657);
and U8598 (N_8598,N_7362,N_8312);
nand U8599 (N_8599,N_8246,N_8138);
xnor U8600 (N_8600,N_7323,N_7620);
or U8601 (N_8601,N_8257,N_7530);
xor U8602 (N_8602,N_7335,N_7274);
and U8603 (N_8603,N_7264,N_7888);
nor U8604 (N_8604,N_8355,N_7754);
xor U8605 (N_8605,N_8156,N_8318);
nor U8606 (N_8606,N_7861,N_7404);
nand U8607 (N_8607,N_7294,N_8214);
xor U8608 (N_8608,N_8305,N_7709);
and U8609 (N_8609,N_8237,N_7860);
nand U8610 (N_8610,N_8163,N_7993);
nand U8611 (N_8611,N_7437,N_7259);
and U8612 (N_8612,N_7343,N_8229);
nand U8613 (N_8613,N_7865,N_8351);
nor U8614 (N_8614,N_7676,N_7743);
nand U8615 (N_8615,N_7376,N_8177);
nand U8616 (N_8616,N_7390,N_7414);
xnor U8617 (N_8617,N_7782,N_7434);
xnor U8618 (N_8618,N_7384,N_7763);
or U8619 (N_8619,N_7831,N_8113);
nor U8620 (N_8620,N_8310,N_7490);
and U8621 (N_8621,N_7662,N_8266);
nor U8622 (N_8622,N_8325,N_8222);
or U8623 (N_8623,N_7967,N_7293);
nand U8624 (N_8624,N_8024,N_8180);
xor U8625 (N_8625,N_7431,N_7415);
or U8626 (N_8626,N_7308,N_7793);
and U8627 (N_8627,N_7451,N_7910);
nand U8628 (N_8628,N_8379,N_8282);
or U8629 (N_8629,N_8133,N_7249);
or U8630 (N_8630,N_7697,N_7702);
nor U8631 (N_8631,N_8275,N_8320);
nand U8632 (N_8632,N_8057,N_7894);
xor U8633 (N_8633,N_7690,N_7459);
xor U8634 (N_8634,N_8192,N_7846);
nor U8635 (N_8635,N_7542,N_8287);
or U8636 (N_8636,N_7553,N_7278);
xnor U8637 (N_8637,N_7368,N_7315);
and U8638 (N_8638,N_7461,N_8359);
nand U8639 (N_8639,N_8045,N_7859);
xnor U8640 (N_8640,N_7272,N_8339);
xor U8641 (N_8641,N_7281,N_7208);
and U8642 (N_8642,N_7565,N_8016);
xor U8643 (N_8643,N_7646,N_8190);
nor U8644 (N_8644,N_8074,N_7716);
nor U8645 (N_8645,N_8086,N_7562);
nand U8646 (N_8646,N_7594,N_8096);
nand U8647 (N_8647,N_8094,N_8183);
or U8648 (N_8648,N_7460,N_7200);
nand U8649 (N_8649,N_8193,N_7252);
or U8650 (N_8650,N_8300,N_7976);
nand U8651 (N_8651,N_7349,N_8118);
nand U8652 (N_8652,N_7499,N_8062);
xnor U8653 (N_8653,N_8075,N_7796);
xnor U8654 (N_8654,N_8211,N_7641);
xnor U8655 (N_8655,N_7304,N_8169);
or U8656 (N_8656,N_7660,N_7601);
and U8657 (N_8657,N_8184,N_7344);
or U8658 (N_8658,N_7964,N_8000);
nor U8659 (N_8659,N_8080,N_8102);
or U8660 (N_8660,N_8089,N_8236);
nand U8661 (N_8661,N_7758,N_8264);
or U8662 (N_8662,N_8202,N_8386);
and U8663 (N_8663,N_8284,N_8170);
and U8664 (N_8664,N_7615,N_7446);
xnor U8665 (N_8665,N_7326,N_7302);
and U8666 (N_8666,N_7202,N_7418);
nand U8667 (N_8667,N_7791,N_8130);
nand U8668 (N_8668,N_7592,N_8077);
or U8669 (N_8669,N_8348,N_7625);
and U8670 (N_8670,N_7306,N_7337);
and U8671 (N_8671,N_7412,N_7843);
xnor U8672 (N_8672,N_7630,N_7889);
or U8673 (N_8673,N_7279,N_7670);
nand U8674 (N_8674,N_7698,N_7577);
nand U8675 (N_8675,N_8233,N_7652);
or U8676 (N_8676,N_7232,N_8067);
nand U8677 (N_8677,N_8261,N_8072);
and U8678 (N_8678,N_8307,N_7206);
nor U8679 (N_8679,N_7298,N_7572);
or U8680 (N_8680,N_8322,N_8208);
and U8681 (N_8681,N_7220,N_7250);
xnor U8682 (N_8682,N_7204,N_8336);
xor U8683 (N_8683,N_8028,N_7909);
xor U8684 (N_8684,N_7478,N_8218);
and U8685 (N_8685,N_8198,N_7808);
or U8686 (N_8686,N_7795,N_8145);
or U8687 (N_8687,N_7605,N_8091);
nand U8688 (N_8688,N_7474,N_7363);
nor U8689 (N_8689,N_7621,N_7550);
and U8690 (N_8690,N_7835,N_8247);
nand U8691 (N_8691,N_8254,N_8101);
xnor U8692 (N_8692,N_7305,N_8304);
nand U8693 (N_8693,N_7899,N_7230);
and U8694 (N_8694,N_8384,N_7906);
or U8695 (N_8695,N_7371,N_7328);
or U8696 (N_8696,N_7240,N_7813);
nand U8697 (N_8697,N_8191,N_7288);
nand U8698 (N_8698,N_7650,N_7506);
nor U8699 (N_8699,N_7956,N_7821);
nor U8700 (N_8700,N_7211,N_7958);
nor U8701 (N_8701,N_7462,N_7353);
or U8702 (N_8702,N_7836,N_7770);
and U8703 (N_8703,N_7694,N_8326);
nor U8704 (N_8704,N_8251,N_7425);
or U8705 (N_8705,N_7571,N_7623);
xor U8706 (N_8706,N_8279,N_7637);
nand U8707 (N_8707,N_7740,N_7399);
or U8708 (N_8708,N_7640,N_8381);
and U8709 (N_8709,N_7921,N_7596);
xnor U8710 (N_8710,N_7303,N_8027);
or U8711 (N_8711,N_7358,N_7475);
or U8712 (N_8712,N_7470,N_8020);
or U8713 (N_8713,N_8250,N_8234);
nand U8714 (N_8714,N_7633,N_8215);
xnor U8715 (N_8715,N_7734,N_7636);
nor U8716 (N_8716,N_8129,N_7248);
and U8717 (N_8717,N_8337,N_8054);
and U8718 (N_8718,N_8259,N_8380);
nand U8719 (N_8719,N_7639,N_8035);
xor U8720 (N_8720,N_8084,N_8392);
and U8721 (N_8721,N_7679,N_7450);
xor U8722 (N_8722,N_7448,N_7890);
or U8723 (N_8723,N_8149,N_7905);
nand U8724 (N_8724,N_7780,N_8269);
xnor U8725 (N_8725,N_7310,N_7300);
and U8726 (N_8726,N_7945,N_7604);
and U8727 (N_8727,N_7725,N_8085);
and U8728 (N_8728,N_8124,N_8274);
xnor U8729 (N_8729,N_7815,N_7547);
nand U8730 (N_8730,N_7994,N_8249);
and U8731 (N_8731,N_7580,N_7978);
nor U8732 (N_8732,N_7672,N_7787);
nand U8733 (N_8733,N_7245,N_7254);
nand U8734 (N_8734,N_8308,N_8225);
nand U8735 (N_8735,N_7606,N_7372);
nand U8736 (N_8736,N_7410,N_7472);
nor U8737 (N_8737,N_7500,N_7485);
xor U8738 (N_8738,N_7634,N_8029);
xnor U8739 (N_8739,N_7738,N_7872);
nand U8740 (N_8740,N_8199,N_7719);
nand U8741 (N_8741,N_7984,N_7355);
nor U8742 (N_8742,N_7406,N_7783);
nor U8743 (N_8743,N_7331,N_7952);
xor U8744 (N_8744,N_7494,N_8095);
nand U8745 (N_8745,N_8073,N_7309);
xnor U8746 (N_8746,N_7792,N_7444);
xnor U8747 (N_8747,N_8083,N_7533);
and U8748 (N_8748,N_7394,N_7881);
and U8749 (N_8749,N_7665,N_7223);
xnor U8750 (N_8750,N_8226,N_8167);
nand U8751 (N_8751,N_8064,N_7463);
and U8752 (N_8752,N_7595,N_7855);
or U8753 (N_8753,N_7333,N_7607);
or U8754 (N_8754,N_8388,N_8343);
and U8755 (N_8755,N_7844,N_7445);
or U8756 (N_8756,N_8176,N_7930);
or U8757 (N_8757,N_8290,N_7299);
xor U8758 (N_8758,N_7876,N_8069);
or U8759 (N_8759,N_7514,N_7803);
or U8760 (N_8760,N_7386,N_8273);
nand U8761 (N_8761,N_8382,N_7352);
and U8762 (N_8762,N_8136,N_8216);
nand U8763 (N_8763,N_8098,N_7336);
nand U8764 (N_8764,N_8303,N_7269);
nand U8765 (N_8765,N_8187,N_8017);
nor U8766 (N_8766,N_7427,N_7433);
xor U8767 (N_8767,N_7877,N_7593);
and U8768 (N_8768,N_8090,N_7401);
xnor U8769 (N_8769,N_8367,N_7616);
or U8770 (N_8770,N_7954,N_7624);
or U8771 (N_8771,N_8068,N_8032);
and U8772 (N_8772,N_7531,N_7396);
or U8773 (N_8773,N_8256,N_7405);
nor U8774 (N_8774,N_7759,N_7817);
xor U8775 (N_8775,N_7387,N_7383);
xor U8776 (N_8776,N_8034,N_7823);
or U8777 (N_8777,N_7949,N_7419);
or U8778 (N_8778,N_7975,N_7962);
or U8779 (N_8779,N_7483,N_7541);
or U8780 (N_8780,N_7409,N_7347);
xor U8781 (N_8781,N_7632,N_7523);
and U8782 (N_8782,N_7439,N_8262);
xnor U8783 (N_8783,N_7654,N_7218);
and U8784 (N_8784,N_7262,N_7365);
nand U8785 (N_8785,N_8171,N_8079);
and U8786 (N_8786,N_7366,N_7487);
nand U8787 (N_8787,N_7745,N_7224);
nand U8788 (N_8788,N_7201,N_7658);
or U8789 (N_8789,N_8023,N_7378);
and U8790 (N_8790,N_7516,N_7752);
and U8791 (N_8791,N_8059,N_7878);
and U8792 (N_8792,N_7449,N_7737);
nor U8793 (N_8793,N_7939,N_8241);
nand U8794 (N_8794,N_7773,N_8037);
or U8795 (N_8795,N_7966,N_7256);
and U8796 (N_8796,N_8006,N_7290);
nand U8797 (N_8797,N_7543,N_7626);
and U8798 (N_8798,N_7871,N_8197);
nor U8799 (N_8799,N_7319,N_7505);
or U8800 (N_8800,N_7257,N_7661);
or U8801 (N_8801,N_8107,N_7755);
nor U8802 (N_8802,N_8363,N_7642);
nand U8803 (N_8803,N_8076,N_7869);
nor U8804 (N_8804,N_7680,N_7285);
nand U8805 (N_8805,N_8010,N_7644);
and U8806 (N_8806,N_8030,N_8070);
and U8807 (N_8807,N_7311,N_7764);
or U8808 (N_8808,N_7569,N_7509);
or U8809 (N_8809,N_7868,N_8334);
xor U8810 (N_8810,N_7705,N_7476);
or U8811 (N_8811,N_7356,N_8105);
or U8812 (N_8812,N_7635,N_7867);
and U8813 (N_8813,N_7848,N_8150);
and U8814 (N_8814,N_7618,N_7267);
or U8815 (N_8815,N_8026,N_7969);
xor U8816 (N_8816,N_7307,N_7297);
nand U8817 (N_8817,N_7819,N_7842);
and U8818 (N_8818,N_8389,N_8046);
xnor U8819 (N_8819,N_7520,N_7678);
nand U8820 (N_8820,N_7613,N_8255);
and U8821 (N_8821,N_7351,N_7229);
or U8822 (N_8822,N_7900,N_8395);
nor U8823 (N_8823,N_8368,N_7558);
nand U8824 (N_8824,N_7369,N_7756);
nand U8825 (N_8825,N_7467,N_8178);
xor U8826 (N_8826,N_8135,N_8397);
and U8827 (N_8827,N_8209,N_8253);
xnor U8828 (N_8828,N_8314,N_7708);
nor U8829 (N_8829,N_8330,N_7922);
nor U8830 (N_8830,N_7271,N_7385);
nand U8831 (N_8831,N_7225,N_8103);
or U8832 (N_8832,N_8393,N_7839);
nand U8833 (N_8833,N_7421,N_7588);
nor U8834 (N_8834,N_8268,N_7513);
and U8835 (N_8835,N_7477,N_7940);
nand U8836 (N_8836,N_7711,N_8306);
nand U8837 (N_8837,N_7581,N_7937);
and U8838 (N_8838,N_8387,N_7651);
or U8839 (N_8839,N_7424,N_8012);
and U8840 (N_8840,N_7786,N_7829);
xnor U8841 (N_8841,N_8350,N_8174);
nand U8842 (N_8842,N_7373,N_8071);
and U8843 (N_8843,N_8099,N_7880);
nand U8844 (N_8844,N_7221,N_7946);
nand U8845 (N_8845,N_7375,N_7681);
nor U8846 (N_8846,N_7268,N_8013);
nor U8847 (N_8847,N_7669,N_7617);
and U8848 (N_8848,N_8302,N_7718);
xnor U8849 (N_8849,N_8104,N_7870);
or U8850 (N_8850,N_7751,N_7788);
and U8851 (N_8851,N_7395,N_7963);
nand U8852 (N_8852,N_7749,N_8340);
and U8853 (N_8853,N_7777,N_8210);
and U8854 (N_8854,N_7925,N_7866);
nor U8855 (N_8855,N_8347,N_7496);
or U8856 (N_8856,N_7851,N_7282);
or U8857 (N_8857,N_7205,N_8001);
or U8858 (N_8858,N_8390,N_7874);
xor U8859 (N_8859,N_7619,N_7438);
nor U8860 (N_8860,N_7895,N_7486);
nor U8861 (N_8861,N_7805,N_8280);
nand U8862 (N_8862,N_8142,N_7330);
or U8863 (N_8863,N_7241,N_7941);
or U8864 (N_8864,N_7760,N_7715);
nor U8865 (N_8865,N_8172,N_7320);
xnor U8866 (N_8866,N_7772,N_8040);
and U8867 (N_8867,N_8230,N_8294);
nor U8868 (N_8868,N_7582,N_8383);
nand U8869 (N_8869,N_8082,N_8060);
and U8870 (N_8870,N_7673,N_7903);
or U8871 (N_8871,N_7599,N_7611);
nand U8872 (N_8872,N_7774,N_8296);
nor U8873 (N_8873,N_8127,N_8182);
xnor U8874 (N_8874,N_7614,N_7578);
xor U8875 (N_8875,N_7432,N_7388);
nand U8876 (N_8876,N_7771,N_8221);
xor U8877 (N_8877,N_7840,N_7653);
or U8878 (N_8878,N_8058,N_7747);
nand U8879 (N_8879,N_8374,N_8286);
xnor U8880 (N_8880,N_7931,N_8158);
or U8881 (N_8881,N_7655,N_7227);
nor U8882 (N_8882,N_7933,N_7948);
xor U8883 (N_8883,N_8309,N_7667);
nand U8884 (N_8884,N_7301,N_7266);
xor U8885 (N_8885,N_8018,N_7928);
nand U8886 (N_8886,N_7913,N_7292);
and U8887 (N_8887,N_7732,N_7701);
or U8888 (N_8888,N_8371,N_7435);
and U8889 (N_8889,N_7253,N_7443);
nor U8890 (N_8890,N_7832,N_8186);
and U8891 (N_8891,N_7998,N_8240);
and U8892 (N_8892,N_7691,N_7458);
xnor U8893 (N_8893,N_8252,N_7389);
or U8894 (N_8894,N_7219,N_7532);
nor U8895 (N_8895,N_8137,N_8258);
nand U8896 (N_8896,N_8332,N_7704);
or U8897 (N_8897,N_7700,N_7992);
nor U8898 (N_8898,N_7341,N_7989);
and U8899 (N_8899,N_7237,N_8165);
nand U8900 (N_8900,N_7915,N_8140);
nand U8901 (N_8901,N_7833,N_8066);
nand U8902 (N_8902,N_7548,N_7566);
nand U8903 (N_8903,N_7576,N_8206);
nand U8904 (N_8904,N_7215,N_7417);
and U8905 (N_8905,N_7350,N_7436);
and U8906 (N_8906,N_8324,N_8015);
xnor U8907 (N_8907,N_8360,N_7236);
xnor U8908 (N_8908,N_8111,N_7454);
xnor U8909 (N_8909,N_8038,N_7280);
nor U8910 (N_8910,N_7828,N_7927);
or U8911 (N_8911,N_8022,N_7235);
xnor U8912 (N_8912,N_7629,N_7858);
xnor U8913 (N_8913,N_8205,N_7243);
and U8914 (N_8914,N_7920,N_7524);
nand U8915 (N_8915,N_7367,N_8063);
xnor U8916 (N_8916,N_7579,N_7263);
and U8917 (N_8917,N_8278,N_7209);
xnor U8918 (N_8918,N_7377,N_8270);
nand U8919 (N_8919,N_7239,N_7979);
or U8920 (N_8920,N_7649,N_7873);
xor U8921 (N_8921,N_7570,N_7273);
and U8922 (N_8922,N_7622,N_7457);
or U8923 (N_8923,N_8372,N_8342);
xor U8924 (N_8924,N_8335,N_7722);
or U8925 (N_8925,N_8097,N_7693);
nand U8926 (N_8926,N_7981,N_7944);
or U8927 (N_8927,N_8093,N_7600);
xnor U8928 (N_8928,N_7970,N_7735);
xnor U8929 (N_8929,N_7456,N_7374);
or U8930 (N_8930,N_7554,N_7370);
or U8931 (N_8931,N_7210,N_7797);
xnor U8932 (N_8932,N_8188,N_7985);
nor U8933 (N_8933,N_7628,N_8005);
nor U8934 (N_8934,N_7990,N_8166);
nand U8935 (N_8935,N_8134,N_7935);
and U8936 (N_8936,N_8328,N_7898);
nor U8937 (N_8937,N_7564,N_8291);
nand U8938 (N_8938,N_8173,N_8271);
or U8939 (N_8939,N_8242,N_7750);
nor U8940 (N_8940,N_8298,N_7932);
and U8941 (N_8941,N_7453,N_7286);
nor U8942 (N_8942,N_7968,N_8345);
nor U8943 (N_8943,N_7357,N_8203);
xor U8944 (N_8944,N_7493,N_8260);
xnor U8945 (N_8945,N_7761,N_7733);
nor U8946 (N_8946,N_7270,N_7529);
nand U8947 (N_8947,N_7659,N_7936);
and U8948 (N_8948,N_7648,N_7647);
nor U8949 (N_8949,N_8121,N_8179);
xor U8950 (N_8950,N_7340,N_7938);
and U8951 (N_8951,N_8293,N_8217);
or U8952 (N_8952,N_7517,N_8061);
xor U8953 (N_8953,N_8353,N_7918);
and U8954 (N_8954,N_7452,N_7923);
or U8955 (N_8955,N_8276,N_7853);
nor U8956 (N_8956,N_8044,N_7233);
nand U8957 (N_8957,N_7591,N_7664);
or U8958 (N_8958,N_8220,N_7724);
xor U8959 (N_8959,N_8088,N_7857);
nand U8960 (N_8960,N_7491,N_7584);
nand U8961 (N_8961,N_8244,N_8164);
xnor U8962 (N_8962,N_8004,N_7258);
xor U8963 (N_8963,N_8162,N_7609);
or U8964 (N_8964,N_7849,N_8289);
and U8965 (N_8965,N_8120,N_8285);
nand U8966 (N_8966,N_7804,N_7919);
xor U8967 (N_8967,N_7407,N_7260);
and U8968 (N_8968,N_7845,N_8049);
or U8969 (N_8969,N_7668,N_8370);
nor U8970 (N_8970,N_7875,N_8281);
or U8971 (N_8971,N_7540,N_8227);
nand U8972 (N_8972,N_7508,N_7392);
or U8973 (N_8973,N_7814,N_7841);
or U8974 (N_8974,N_7645,N_7810);
nor U8975 (N_8975,N_8369,N_7429);
and U8976 (N_8976,N_8021,N_8319);
and U8977 (N_8977,N_7231,N_8349);
or U8978 (N_8978,N_7519,N_7914);
xnor U8979 (N_8979,N_7535,N_7721);
nand U8980 (N_8980,N_8168,N_8338);
xnor U8981 (N_8981,N_7295,N_8181);
and U8982 (N_8982,N_7521,N_7561);
and U8983 (N_8983,N_7545,N_7713);
nand U8984 (N_8984,N_8139,N_8365);
and U8985 (N_8985,N_7361,N_7663);
nand U8986 (N_8986,N_8385,N_7955);
and U8987 (N_8987,N_7971,N_8248);
or U8988 (N_8988,N_8036,N_8002);
nor U8989 (N_8989,N_7912,N_7393);
or U8990 (N_8990,N_8131,N_7983);
nand U8991 (N_8991,N_7879,N_7222);
nand U8992 (N_8992,N_7746,N_7916);
xor U8993 (N_8993,N_7510,N_7332);
nor U8994 (N_8994,N_7856,N_7455);
or U8995 (N_8995,N_7847,N_7775);
or U8996 (N_8996,N_8052,N_8346);
and U8997 (N_8997,N_7884,N_7886);
or U8998 (N_8998,N_7276,N_8048);
xor U8999 (N_8999,N_7977,N_8376);
nand U9000 (N_9000,N_7925,N_7801);
xor U9001 (N_9001,N_8044,N_7902);
xor U9002 (N_9002,N_7373,N_8188);
xor U9003 (N_9003,N_7807,N_8252);
nor U9004 (N_9004,N_7351,N_7764);
or U9005 (N_9005,N_8350,N_7788);
and U9006 (N_9006,N_8252,N_7831);
xor U9007 (N_9007,N_7667,N_7646);
or U9008 (N_9008,N_7588,N_7959);
nand U9009 (N_9009,N_7792,N_7822);
and U9010 (N_9010,N_7635,N_7295);
xor U9011 (N_9011,N_7618,N_7497);
nor U9012 (N_9012,N_7351,N_7750);
nand U9013 (N_9013,N_7512,N_8033);
nand U9014 (N_9014,N_7995,N_7533);
nor U9015 (N_9015,N_7408,N_7613);
or U9016 (N_9016,N_7398,N_7720);
or U9017 (N_9017,N_8144,N_7480);
and U9018 (N_9018,N_7640,N_7420);
nand U9019 (N_9019,N_7983,N_7270);
xnor U9020 (N_9020,N_7790,N_8061);
xnor U9021 (N_9021,N_8272,N_7532);
nor U9022 (N_9022,N_8302,N_7407);
nor U9023 (N_9023,N_7380,N_7258);
or U9024 (N_9024,N_7485,N_7929);
and U9025 (N_9025,N_7316,N_7897);
nand U9026 (N_9026,N_7262,N_7250);
nor U9027 (N_9027,N_8237,N_8214);
and U9028 (N_9028,N_8118,N_8112);
or U9029 (N_9029,N_7611,N_8206);
nand U9030 (N_9030,N_7710,N_7671);
xnor U9031 (N_9031,N_7651,N_8085);
or U9032 (N_9032,N_7313,N_8060);
nand U9033 (N_9033,N_8295,N_8153);
and U9034 (N_9034,N_7292,N_7588);
nor U9035 (N_9035,N_7390,N_7849);
xnor U9036 (N_9036,N_7907,N_7868);
or U9037 (N_9037,N_7265,N_8252);
xor U9038 (N_9038,N_8154,N_7973);
xnor U9039 (N_9039,N_7338,N_8177);
or U9040 (N_9040,N_7276,N_8364);
or U9041 (N_9041,N_7314,N_7769);
or U9042 (N_9042,N_7704,N_7584);
and U9043 (N_9043,N_8376,N_7651);
and U9044 (N_9044,N_8251,N_7925);
nand U9045 (N_9045,N_8396,N_7769);
or U9046 (N_9046,N_8170,N_7371);
nor U9047 (N_9047,N_7833,N_8273);
or U9048 (N_9048,N_7899,N_8236);
nor U9049 (N_9049,N_7336,N_8201);
xnor U9050 (N_9050,N_7870,N_7207);
and U9051 (N_9051,N_7774,N_7966);
and U9052 (N_9052,N_7585,N_8068);
nand U9053 (N_9053,N_7622,N_7848);
xor U9054 (N_9054,N_7817,N_7969);
nand U9055 (N_9055,N_7969,N_8002);
and U9056 (N_9056,N_8228,N_7612);
or U9057 (N_9057,N_7383,N_7496);
or U9058 (N_9058,N_7694,N_7907);
nor U9059 (N_9059,N_7709,N_8387);
or U9060 (N_9060,N_7640,N_7706);
and U9061 (N_9061,N_8100,N_8131);
nand U9062 (N_9062,N_8135,N_8300);
or U9063 (N_9063,N_7400,N_7640);
xnor U9064 (N_9064,N_8045,N_7358);
xnor U9065 (N_9065,N_7724,N_8289);
nor U9066 (N_9066,N_8172,N_7525);
and U9067 (N_9067,N_7810,N_8366);
nand U9068 (N_9068,N_7889,N_7659);
or U9069 (N_9069,N_8368,N_8171);
nor U9070 (N_9070,N_7526,N_7971);
or U9071 (N_9071,N_7422,N_7628);
xor U9072 (N_9072,N_7855,N_7620);
and U9073 (N_9073,N_8064,N_7388);
nor U9074 (N_9074,N_7417,N_7893);
xor U9075 (N_9075,N_7504,N_7729);
nor U9076 (N_9076,N_7324,N_7586);
nand U9077 (N_9077,N_7934,N_8204);
and U9078 (N_9078,N_7722,N_7242);
nand U9079 (N_9079,N_8388,N_7628);
and U9080 (N_9080,N_7803,N_8029);
or U9081 (N_9081,N_7336,N_8102);
and U9082 (N_9082,N_7942,N_7202);
nor U9083 (N_9083,N_8130,N_7973);
nand U9084 (N_9084,N_7675,N_8354);
and U9085 (N_9085,N_7701,N_7583);
nand U9086 (N_9086,N_7355,N_7624);
and U9087 (N_9087,N_7469,N_7800);
and U9088 (N_9088,N_8303,N_7647);
nor U9089 (N_9089,N_7780,N_7384);
nor U9090 (N_9090,N_7659,N_8190);
and U9091 (N_9091,N_8228,N_7543);
nand U9092 (N_9092,N_8381,N_7936);
nor U9093 (N_9093,N_7831,N_7518);
and U9094 (N_9094,N_7346,N_7762);
or U9095 (N_9095,N_8238,N_7684);
and U9096 (N_9096,N_8188,N_7296);
nand U9097 (N_9097,N_7430,N_7288);
nand U9098 (N_9098,N_7920,N_8348);
nor U9099 (N_9099,N_7603,N_8188);
xnor U9100 (N_9100,N_7606,N_7592);
or U9101 (N_9101,N_8164,N_7862);
nor U9102 (N_9102,N_7222,N_8020);
and U9103 (N_9103,N_8001,N_7421);
nand U9104 (N_9104,N_7284,N_7235);
or U9105 (N_9105,N_7224,N_7955);
nor U9106 (N_9106,N_7605,N_7591);
nor U9107 (N_9107,N_7957,N_7902);
or U9108 (N_9108,N_7897,N_8363);
nand U9109 (N_9109,N_7950,N_7746);
or U9110 (N_9110,N_7738,N_7376);
and U9111 (N_9111,N_8326,N_8075);
or U9112 (N_9112,N_8302,N_7627);
nand U9113 (N_9113,N_8381,N_7326);
nand U9114 (N_9114,N_7859,N_8052);
xnor U9115 (N_9115,N_7495,N_8179);
xor U9116 (N_9116,N_7813,N_7793);
nand U9117 (N_9117,N_8331,N_7759);
nand U9118 (N_9118,N_7464,N_8342);
nor U9119 (N_9119,N_7999,N_7441);
nand U9120 (N_9120,N_7581,N_7218);
nor U9121 (N_9121,N_8231,N_7742);
nor U9122 (N_9122,N_7282,N_8169);
xnor U9123 (N_9123,N_7689,N_7269);
or U9124 (N_9124,N_8361,N_8287);
xor U9125 (N_9125,N_7483,N_7507);
nand U9126 (N_9126,N_7949,N_7561);
xor U9127 (N_9127,N_7497,N_7971);
or U9128 (N_9128,N_7742,N_7999);
xor U9129 (N_9129,N_7627,N_7573);
or U9130 (N_9130,N_8259,N_8226);
nor U9131 (N_9131,N_7268,N_7729);
and U9132 (N_9132,N_7465,N_7694);
or U9133 (N_9133,N_7685,N_8268);
or U9134 (N_9134,N_8372,N_7213);
nand U9135 (N_9135,N_8213,N_8184);
nand U9136 (N_9136,N_7871,N_7263);
and U9137 (N_9137,N_8197,N_7840);
and U9138 (N_9138,N_7769,N_7730);
and U9139 (N_9139,N_7791,N_7410);
nand U9140 (N_9140,N_7905,N_7351);
nand U9141 (N_9141,N_7797,N_7641);
xnor U9142 (N_9142,N_7360,N_7583);
xnor U9143 (N_9143,N_8038,N_7413);
nor U9144 (N_9144,N_7271,N_7381);
xnor U9145 (N_9145,N_7749,N_7909);
nand U9146 (N_9146,N_7252,N_8231);
or U9147 (N_9147,N_8374,N_8020);
nand U9148 (N_9148,N_7232,N_8266);
xnor U9149 (N_9149,N_7927,N_7877);
or U9150 (N_9150,N_7684,N_7731);
nor U9151 (N_9151,N_7653,N_7830);
nand U9152 (N_9152,N_7697,N_7489);
nor U9153 (N_9153,N_8091,N_7830);
nor U9154 (N_9154,N_7496,N_7946);
xor U9155 (N_9155,N_7855,N_7650);
and U9156 (N_9156,N_7397,N_8283);
nor U9157 (N_9157,N_8077,N_7220);
or U9158 (N_9158,N_7407,N_7457);
nand U9159 (N_9159,N_8121,N_7794);
nand U9160 (N_9160,N_7881,N_7935);
nor U9161 (N_9161,N_7518,N_8060);
nand U9162 (N_9162,N_7550,N_7739);
or U9163 (N_9163,N_7872,N_8347);
xnor U9164 (N_9164,N_7513,N_7704);
nor U9165 (N_9165,N_7535,N_7252);
nor U9166 (N_9166,N_7719,N_7740);
nor U9167 (N_9167,N_7226,N_7656);
and U9168 (N_9168,N_8179,N_7858);
or U9169 (N_9169,N_7909,N_7922);
and U9170 (N_9170,N_7544,N_7710);
xnor U9171 (N_9171,N_7941,N_8228);
xnor U9172 (N_9172,N_7350,N_7854);
nor U9173 (N_9173,N_7871,N_7443);
xnor U9174 (N_9174,N_7555,N_7856);
or U9175 (N_9175,N_7904,N_7316);
xor U9176 (N_9176,N_7395,N_7522);
or U9177 (N_9177,N_8028,N_7377);
or U9178 (N_9178,N_7796,N_7837);
nand U9179 (N_9179,N_7776,N_7621);
xnor U9180 (N_9180,N_7281,N_7249);
and U9181 (N_9181,N_8257,N_7490);
or U9182 (N_9182,N_7529,N_7740);
and U9183 (N_9183,N_7290,N_8291);
nand U9184 (N_9184,N_8132,N_8396);
xnor U9185 (N_9185,N_7284,N_7559);
nor U9186 (N_9186,N_7699,N_7830);
nor U9187 (N_9187,N_8191,N_7676);
xor U9188 (N_9188,N_8136,N_7716);
or U9189 (N_9189,N_8056,N_7757);
xnor U9190 (N_9190,N_7780,N_7311);
and U9191 (N_9191,N_7833,N_8068);
and U9192 (N_9192,N_8030,N_8167);
nor U9193 (N_9193,N_7279,N_7205);
nand U9194 (N_9194,N_7331,N_8231);
or U9195 (N_9195,N_7203,N_7716);
nand U9196 (N_9196,N_8037,N_8048);
xnor U9197 (N_9197,N_8081,N_8110);
or U9198 (N_9198,N_7535,N_8218);
xor U9199 (N_9199,N_8069,N_8093);
xor U9200 (N_9200,N_7803,N_7990);
or U9201 (N_9201,N_8292,N_8282);
xor U9202 (N_9202,N_7844,N_8195);
nor U9203 (N_9203,N_7932,N_8381);
nor U9204 (N_9204,N_7585,N_7842);
nor U9205 (N_9205,N_7940,N_7759);
nand U9206 (N_9206,N_7977,N_7818);
nand U9207 (N_9207,N_7927,N_7264);
nor U9208 (N_9208,N_7371,N_7224);
or U9209 (N_9209,N_7204,N_7300);
xor U9210 (N_9210,N_7324,N_7408);
or U9211 (N_9211,N_8276,N_7720);
or U9212 (N_9212,N_7511,N_7349);
or U9213 (N_9213,N_7717,N_8225);
xor U9214 (N_9214,N_8251,N_7698);
and U9215 (N_9215,N_7931,N_8231);
nand U9216 (N_9216,N_7713,N_7783);
nor U9217 (N_9217,N_8219,N_7775);
nand U9218 (N_9218,N_7778,N_8088);
xor U9219 (N_9219,N_7734,N_8031);
nand U9220 (N_9220,N_8010,N_8074);
and U9221 (N_9221,N_8190,N_7204);
and U9222 (N_9222,N_8387,N_7874);
or U9223 (N_9223,N_8353,N_7333);
and U9224 (N_9224,N_8398,N_8037);
nor U9225 (N_9225,N_8098,N_7341);
nand U9226 (N_9226,N_7827,N_8351);
or U9227 (N_9227,N_7505,N_7626);
and U9228 (N_9228,N_7902,N_8284);
nand U9229 (N_9229,N_7658,N_7900);
xor U9230 (N_9230,N_7551,N_7953);
nand U9231 (N_9231,N_7932,N_7891);
xor U9232 (N_9232,N_7807,N_7827);
or U9233 (N_9233,N_8041,N_7511);
xnor U9234 (N_9234,N_8347,N_7232);
xor U9235 (N_9235,N_7529,N_7591);
nor U9236 (N_9236,N_7458,N_8267);
and U9237 (N_9237,N_7873,N_8295);
nand U9238 (N_9238,N_8174,N_7403);
or U9239 (N_9239,N_7834,N_8191);
and U9240 (N_9240,N_7608,N_8160);
and U9241 (N_9241,N_7475,N_8203);
nand U9242 (N_9242,N_7754,N_8022);
nor U9243 (N_9243,N_8357,N_7605);
nand U9244 (N_9244,N_8124,N_7915);
nand U9245 (N_9245,N_7801,N_7941);
and U9246 (N_9246,N_8025,N_7219);
or U9247 (N_9247,N_8136,N_8162);
nand U9248 (N_9248,N_7930,N_7712);
nor U9249 (N_9249,N_8322,N_7766);
xnor U9250 (N_9250,N_7200,N_8003);
nor U9251 (N_9251,N_8181,N_7239);
xnor U9252 (N_9252,N_7377,N_8003);
xor U9253 (N_9253,N_7757,N_8321);
and U9254 (N_9254,N_7382,N_7412);
or U9255 (N_9255,N_7560,N_8095);
or U9256 (N_9256,N_8124,N_7660);
xnor U9257 (N_9257,N_8016,N_7528);
nor U9258 (N_9258,N_7277,N_7620);
nor U9259 (N_9259,N_7920,N_7394);
nor U9260 (N_9260,N_7819,N_8382);
nand U9261 (N_9261,N_8379,N_8215);
or U9262 (N_9262,N_7427,N_7777);
nand U9263 (N_9263,N_7219,N_7210);
nand U9264 (N_9264,N_8068,N_7256);
or U9265 (N_9265,N_7661,N_7874);
xor U9266 (N_9266,N_7259,N_7729);
or U9267 (N_9267,N_8100,N_8395);
nand U9268 (N_9268,N_7289,N_7564);
nand U9269 (N_9269,N_7925,N_7328);
or U9270 (N_9270,N_8043,N_8026);
nor U9271 (N_9271,N_7409,N_8200);
and U9272 (N_9272,N_7889,N_8164);
and U9273 (N_9273,N_7673,N_7860);
or U9274 (N_9274,N_7308,N_8232);
nor U9275 (N_9275,N_7605,N_7819);
nand U9276 (N_9276,N_7401,N_8120);
and U9277 (N_9277,N_8042,N_7506);
or U9278 (N_9278,N_7370,N_7814);
nor U9279 (N_9279,N_7884,N_7550);
and U9280 (N_9280,N_7514,N_8361);
nor U9281 (N_9281,N_7879,N_7482);
nand U9282 (N_9282,N_7919,N_7461);
xor U9283 (N_9283,N_8195,N_7828);
or U9284 (N_9284,N_7218,N_8153);
nor U9285 (N_9285,N_7726,N_7515);
or U9286 (N_9286,N_7363,N_7203);
nand U9287 (N_9287,N_7773,N_8297);
xnor U9288 (N_9288,N_7263,N_8366);
nor U9289 (N_9289,N_7783,N_7509);
xnor U9290 (N_9290,N_7394,N_8307);
nand U9291 (N_9291,N_7230,N_7688);
or U9292 (N_9292,N_7981,N_7636);
nor U9293 (N_9293,N_8074,N_7855);
xnor U9294 (N_9294,N_7644,N_7966);
xnor U9295 (N_9295,N_7275,N_7361);
xor U9296 (N_9296,N_7801,N_7824);
nor U9297 (N_9297,N_7478,N_7781);
xnor U9298 (N_9298,N_8188,N_7751);
nor U9299 (N_9299,N_7617,N_7384);
nand U9300 (N_9300,N_7732,N_7803);
or U9301 (N_9301,N_8108,N_7583);
and U9302 (N_9302,N_8151,N_8230);
nor U9303 (N_9303,N_7824,N_7728);
or U9304 (N_9304,N_8227,N_7771);
and U9305 (N_9305,N_7316,N_8097);
nand U9306 (N_9306,N_8103,N_7284);
and U9307 (N_9307,N_7531,N_7315);
xor U9308 (N_9308,N_7782,N_8288);
xor U9309 (N_9309,N_8143,N_7347);
nand U9310 (N_9310,N_7651,N_7512);
nor U9311 (N_9311,N_7432,N_7386);
or U9312 (N_9312,N_7400,N_7605);
and U9313 (N_9313,N_8240,N_7790);
or U9314 (N_9314,N_7865,N_7606);
or U9315 (N_9315,N_7745,N_7326);
xnor U9316 (N_9316,N_7286,N_7655);
and U9317 (N_9317,N_7243,N_7617);
nor U9318 (N_9318,N_8127,N_7262);
and U9319 (N_9319,N_8106,N_7219);
nand U9320 (N_9320,N_7880,N_7691);
xor U9321 (N_9321,N_7884,N_7289);
xnor U9322 (N_9322,N_8375,N_7733);
xor U9323 (N_9323,N_8073,N_7464);
nand U9324 (N_9324,N_8094,N_7925);
and U9325 (N_9325,N_7674,N_7893);
xor U9326 (N_9326,N_7718,N_7817);
and U9327 (N_9327,N_7910,N_7576);
and U9328 (N_9328,N_8106,N_7444);
and U9329 (N_9329,N_7971,N_8231);
or U9330 (N_9330,N_8140,N_7527);
nor U9331 (N_9331,N_8006,N_7643);
nand U9332 (N_9332,N_7539,N_8255);
and U9333 (N_9333,N_7298,N_7925);
nand U9334 (N_9334,N_7476,N_7569);
xor U9335 (N_9335,N_8368,N_7991);
or U9336 (N_9336,N_7684,N_7622);
nand U9337 (N_9337,N_7531,N_7606);
or U9338 (N_9338,N_7436,N_8331);
xnor U9339 (N_9339,N_7994,N_7222);
nand U9340 (N_9340,N_7397,N_7838);
or U9341 (N_9341,N_8391,N_7459);
nand U9342 (N_9342,N_7350,N_7965);
nand U9343 (N_9343,N_8208,N_8095);
nor U9344 (N_9344,N_7460,N_8141);
and U9345 (N_9345,N_7510,N_7278);
xnor U9346 (N_9346,N_7451,N_7341);
nor U9347 (N_9347,N_7738,N_8348);
and U9348 (N_9348,N_8131,N_7578);
or U9349 (N_9349,N_7966,N_8246);
and U9350 (N_9350,N_8048,N_7546);
and U9351 (N_9351,N_8074,N_7994);
nor U9352 (N_9352,N_8115,N_7864);
nand U9353 (N_9353,N_7588,N_7246);
and U9354 (N_9354,N_7962,N_7672);
nand U9355 (N_9355,N_7933,N_8294);
or U9356 (N_9356,N_7714,N_8298);
or U9357 (N_9357,N_7940,N_7372);
nand U9358 (N_9358,N_7647,N_7328);
or U9359 (N_9359,N_8113,N_7881);
and U9360 (N_9360,N_7345,N_7840);
nor U9361 (N_9361,N_7987,N_8050);
nand U9362 (N_9362,N_7869,N_7386);
or U9363 (N_9363,N_8251,N_7435);
xnor U9364 (N_9364,N_7688,N_7830);
and U9365 (N_9365,N_8314,N_7320);
xor U9366 (N_9366,N_8220,N_7880);
xor U9367 (N_9367,N_7768,N_7615);
nor U9368 (N_9368,N_7916,N_8382);
nor U9369 (N_9369,N_7442,N_8219);
and U9370 (N_9370,N_7993,N_7666);
or U9371 (N_9371,N_8014,N_7262);
nand U9372 (N_9372,N_7994,N_8313);
nor U9373 (N_9373,N_7334,N_7401);
or U9374 (N_9374,N_8104,N_7401);
or U9375 (N_9375,N_7318,N_8190);
or U9376 (N_9376,N_7722,N_8136);
xnor U9377 (N_9377,N_8375,N_7757);
nand U9378 (N_9378,N_8152,N_8057);
nor U9379 (N_9379,N_8174,N_8072);
or U9380 (N_9380,N_7787,N_8025);
nand U9381 (N_9381,N_8183,N_7391);
or U9382 (N_9382,N_8237,N_7729);
nor U9383 (N_9383,N_7352,N_7288);
xor U9384 (N_9384,N_7846,N_8366);
and U9385 (N_9385,N_7964,N_7585);
and U9386 (N_9386,N_7895,N_7645);
and U9387 (N_9387,N_8012,N_8178);
xor U9388 (N_9388,N_7394,N_7627);
nor U9389 (N_9389,N_7564,N_7863);
nor U9390 (N_9390,N_8369,N_8013);
nand U9391 (N_9391,N_7938,N_7945);
nor U9392 (N_9392,N_7797,N_7575);
nor U9393 (N_9393,N_8123,N_7657);
nor U9394 (N_9394,N_7522,N_7502);
xor U9395 (N_9395,N_8269,N_7731);
and U9396 (N_9396,N_7780,N_7699);
or U9397 (N_9397,N_8317,N_7924);
and U9398 (N_9398,N_8217,N_7916);
nor U9399 (N_9399,N_8148,N_7659);
nand U9400 (N_9400,N_7778,N_7727);
or U9401 (N_9401,N_7607,N_7603);
nor U9402 (N_9402,N_7612,N_8163);
or U9403 (N_9403,N_7620,N_7470);
nand U9404 (N_9404,N_7289,N_8190);
xor U9405 (N_9405,N_8244,N_8015);
xor U9406 (N_9406,N_7429,N_7549);
or U9407 (N_9407,N_7886,N_7955);
nor U9408 (N_9408,N_7626,N_8287);
nand U9409 (N_9409,N_8081,N_8262);
and U9410 (N_9410,N_8353,N_7700);
nand U9411 (N_9411,N_8225,N_7539);
nand U9412 (N_9412,N_7978,N_7611);
and U9413 (N_9413,N_7265,N_8187);
or U9414 (N_9414,N_7618,N_7226);
and U9415 (N_9415,N_7911,N_8041);
and U9416 (N_9416,N_8010,N_7426);
nand U9417 (N_9417,N_7285,N_7372);
nand U9418 (N_9418,N_7750,N_8394);
or U9419 (N_9419,N_7719,N_7834);
and U9420 (N_9420,N_7590,N_7905);
xor U9421 (N_9421,N_8393,N_7223);
or U9422 (N_9422,N_7371,N_8091);
nand U9423 (N_9423,N_7410,N_8375);
xor U9424 (N_9424,N_7975,N_8133);
and U9425 (N_9425,N_7861,N_7492);
nand U9426 (N_9426,N_7491,N_8257);
nor U9427 (N_9427,N_7860,N_7975);
nor U9428 (N_9428,N_7745,N_7578);
nor U9429 (N_9429,N_7477,N_7326);
or U9430 (N_9430,N_8381,N_7754);
nand U9431 (N_9431,N_8035,N_7619);
and U9432 (N_9432,N_8099,N_7609);
xor U9433 (N_9433,N_7505,N_8245);
or U9434 (N_9434,N_7804,N_7535);
and U9435 (N_9435,N_7476,N_8188);
nand U9436 (N_9436,N_8065,N_7871);
or U9437 (N_9437,N_8143,N_8379);
or U9438 (N_9438,N_8301,N_7784);
and U9439 (N_9439,N_7861,N_7727);
or U9440 (N_9440,N_7504,N_8312);
or U9441 (N_9441,N_8131,N_7962);
nand U9442 (N_9442,N_8136,N_7477);
or U9443 (N_9443,N_7958,N_7303);
xnor U9444 (N_9444,N_7822,N_8083);
and U9445 (N_9445,N_7440,N_7789);
or U9446 (N_9446,N_7324,N_7969);
or U9447 (N_9447,N_7209,N_7246);
and U9448 (N_9448,N_8313,N_7993);
or U9449 (N_9449,N_8018,N_7950);
or U9450 (N_9450,N_7267,N_8294);
nand U9451 (N_9451,N_8206,N_7277);
nor U9452 (N_9452,N_7202,N_7637);
and U9453 (N_9453,N_7676,N_7328);
xor U9454 (N_9454,N_8245,N_7383);
xor U9455 (N_9455,N_8375,N_8012);
nand U9456 (N_9456,N_7345,N_7255);
or U9457 (N_9457,N_7631,N_7888);
or U9458 (N_9458,N_8253,N_7666);
and U9459 (N_9459,N_7372,N_8162);
and U9460 (N_9460,N_7233,N_8236);
xnor U9461 (N_9461,N_7449,N_7233);
nor U9462 (N_9462,N_7277,N_7288);
nand U9463 (N_9463,N_7873,N_7522);
xnor U9464 (N_9464,N_8265,N_7893);
or U9465 (N_9465,N_8039,N_7693);
nor U9466 (N_9466,N_8340,N_7221);
nand U9467 (N_9467,N_7394,N_7243);
nor U9468 (N_9468,N_7364,N_8370);
nor U9469 (N_9469,N_7898,N_7465);
and U9470 (N_9470,N_7556,N_7336);
nand U9471 (N_9471,N_8119,N_7200);
or U9472 (N_9472,N_7637,N_7946);
nand U9473 (N_9473,N_8397,N_7500);
and U9474 (N_9474,N_8334,N_8225);
xnor U9475 (N_9475,N_7928,N_7225);
nand U9476 (N_9476,N_7961,N_7243);
xor U9477 (N_9477,N_7384,N_8259);
nand U9478 (N_9478,N_8316,N_8389);
xor U9479 (N_9479,N_7475,N_7957);
xor U9480 (N_9480,N_8196,N_8127);
or U9481 (N_9481,N_7437,N_7559);
xor U9482 (N_9482,N_7572,N_8369);
or U9483 (N_9483,N_7912,N_8146);
and U9484 (N_9484,N_7345,N_7492);
and U9485 (N_9485,N_7595,N_7636);
and U9486 (N_9486,N_8163,N_7565);
xor U9487 (N_9487,N_7564,N_8378);
nor U9488 (N_9488,N_7870,N_7266);
nand U9489 (N_9489,N_7998,N_7621);
xnor U9490 (N_9490,N_8377,N_7984);
or U9491 (N_9491,N_7439,N_8040);
or U9492 (N_9492,N_8180,N_8141);
nand U9493 (N_9493,N_8376,N_8225);
nand U9494 (N_9494,N_7329,N_7324);
or U9495 (N_9495,N_7674,N_8086);
nor U9496 (N_9496,N_7299,N_8008);
and U9497 (N_9497,N_8237,N_7579);
or U9498 (N_9498,N_7849,N_7756);
nand U9499 (N_9499,N_8081,N_8035);
xnor U9500 (N_9500,N_7983,N_7962);
nand U9501 (N_9501,N_7447,N_7292);
xnor U9502 (N_9502,N_7592,N_8022);
nor U9503 (N_9503,N_7407,N_7415);
xor U9504 (N_9504,N_7282,N_7784);
xor U9505 (N_9505,N_7973,N_7368);
nor U9506 (N_9506,N_7752,N_7818);
or U9507 (N_9507,N_8072,N_7234);
or U9508 (N_9508,N_7397,N_8381);
and U9509 (N_9509,N_7478,N_7658);
nand U9510 (N_9510,N_7859,N_7967);
nand U9511 (N_9511,N_7509,N_8071);
nor U9512 (N_9512,N_7836,N_8208);
nand U9513 (N_9513,N_7232,N_8058);
nand U9514 (N_9514,N_7538,N_7442);
or U9515 (N_9515,N_7576,N_7777);
nor U9516 (N_9516,N_8310,N_7695);
xnor U9517 (N_9517,N_8225,N_8371);
or U9518 (N_9518,N_7583,N_7250);
xnor U9519 (N_9519,N_7207,N_7282);
or U9520 (N_9520,N_8109,N_7281);
xor U9521 (N_9521,N_7969,N_7311);
xnor U9522 (N_9522,N_7217,N_7695);
or U9523 (N_9523,N_8300,N_7748);
or U9524 (N_9524,N_7792,N_7953);
nor U9525 (N_9525,N_8374,N_7752);
or U9526 (N_9526,N_7726,N_7745);
xnor U9527 (N_9527,N_7917,N_7398);
or U9528 (N_9528,N_8143,N_7744);
xor U9529 (N_9529,N_7561,N_8294);
xor U9530 (N_9530,N_7793,N_7764);
nor U9531 (N_9531,N_7579,N_7367);
or U9532 (N_9532,N_7485,N_8126);
nor U9533 (N_9533,N_7586,N_8175);
and U9534 (N_9534,N_8211,N_7374);
and U9535 (N_9535,N_8179,N_7783);
xor U9536 (N_9536,N_8249,N_8376);
or U9537 (N_9537,N_7627,N_8066);
xor U9538 (N_9538,N_8327,N_7300);
or U9539 (N_9539,N_7826,N_7332);
and U9540 (N_9540,N_7616,N_7705);
nor U9541 (N_9541,N_7455,N_7232);
or U9542 (N_9542,N_8314,N_7680);
and U9543 (N_9543,N_7307,N_7517);
nand U9544 (N_9544,N_8355,N_8108);
nand U9545 (N_9545,N_7715,N_8388);
nor U9546 (N_9546,N_8122,N_7217);
xor U9547 (N_9547,N_7232,N_7477);
and U9548 (N_9548,N_7928,N_7765);
or U9549 (N_9549,N_7336,N_8099);
xnor U9550 (N_9550,N_7963,N_7327);
xnor U9551 (N_9551,N_7716,N_7583);
xor U9552 (N_9552,N_8327,N_7829);
or U9553 (N_9553,N_7837,N_7375);
or U9554 (N_9554,N_7251,N_7769);
or U9555 (N_9555,N_7518,N_7593);
nand U9556 (N_9556,N_8031,N_7263);
nand U9557 (N_9557,N_7816,N_7604);
xnor U9558 (N_9558,N_7430,N_7405);
or U9559 (N_9559,N_7793,N_8125);
nand U9560 (N_9560,N_7567,N_8251);
xnor U9561 (N_9561,N_7249,N_7590);
or U9562 (N_9562,N_8116,N_7786);
or U9563 (N_9563,N_8023,N_7354);
and U9564 (N_9564,N_7217,N_8050);
or U9565 (N_9565,N_7595,N_8012);
or U9566 (N_9566,N_7669,N_7739);
or U9567 (N_9567,N_7768,N_7989);
nand U9568 (N_9568,N_7874,N_8281);
nand U9569 (N_9569,N_7984,N_7574);
nor U9570 (N_9570,N_7574,N_7343);
and U9571 (N_9571,N_7497,N_7313);
and U9572 (N_9572,N_7789,N_7487);
nor U9573 (N_9573,N_7772,N_8047);
nor U9574 (N_9574,N_8199,N_7813);
nand U9575 (N_9575,N_7402,N_7775);
nor U9576 (N_9576,N_7377,N_8017);
nor U9577 (N_9577,N_8027,N_7998);
nand U9578 (N_9578,N_7840,N_8215);
nand U9579 (N_9579,N_8265,N_7289);
and U9580 (N_9580,N_8076,N_8370);
or U9581 (N_9581,N_7972,N_8016);
nor U9582 (N_9582,N_7227,N_7890);
xnor U9583 (N_9583,N_7952,N_7612);
or U9584 (N_9584,N_8085,N_7730);
and U9585 (N_9585,N_7911,N_7437);
or U9586 (N_9586,N_7324,N_8093);
nand U9587 (N_9587,N_7522,N_8250);
or U9588 (N_9588,N_7295,N_7858);
nand U9589 (N_9589,N_7563,N_7291);
xor U9590 (N_9590,N_7411,N_8151);
and U9591 (N_9591,N_7681,N_7476);
xnor U9592 (N_9592,N_8224,N_8047);
xnor U9593 (N_9593,N_8342,N_7817);
xnor U9594 (N_9594,N_7996,N_7854);
xor U9595 (N_9595,N_7864,N_7789);
or U9596 (N_9596,N_7774,N_8174);
nand U9597 (N_9597,N_7713,N_7273);
nor U9598 (N_9598,N_7541,N_7846);
nand U9599 (N_9599,N_7583,N_7694);
nor U9600 (N_9600,N_9577,N_8966);
nor U9601 (N_9601,N_9395,N_9153);
and U9602 (N_9602,N_8791,N_8731);
and U9603 (N_9603,N_9090,N_9144);
xor U9604 (N_9604,N_8546,N_8543);
and U9605 (N_9605,N_8887,N_9214);
xnor U9606 (N_9606,N_8679,N_8490);
nand U9607 (N_9607,N_9010,N_9496);
or U9608 (N_9608,N_9277,N_9064);
nor U9609 (N_9609,N_8661,N_8693);
nand U9610 (N_9610,N_8676,N_8720);
xor U9611 (N_9611,N_9342,N_8770);
and U9612 (N_9612,N_8835,N_9231);
or U9613 (N_9613,N_8939,N_9505);
or U9614 (N_9614,N_8483,N_8715);
xor U9615 (N_9615,N_9523,N_8656);
nor U9616 (N_9616,N_9338,N_8618);
and U9617 (N_9617,N_8487,N_9442);
or U9618 (N_9618,N_8607,N_8511);
or U9619 (N_9619,N_8570,N_8517);
nand U9620 (N_9620,N_8502,N_8950);
or U9621 (N_9621,N_9202,N_9264);
or U9622 (N_9622,N_9100,N_8574);
xor U9623 (N_9623,N_9460,N_8523);
and U9624 (N_9624,N_9131,N_9288);
and U9625 (N_9625,N_9519,N_8752);
and U9626 (N_9626,N_9418,N_9016);
xnor U9627 (N_9627,N_8905,N_8562);
and U9628 (N_9628,N_9116,N_8444);
and U9629 (N_9629,N_8780,N_9278);
xnor U9630 (N_9630,N_9526,N_9066);
xnor U9631 (N_9631,N_8684,N_9017);
nor U9632 (N_9632,N_9268,N_8500);
xnor U9633 (N_9633,N_9472,N_9341);
or U9634 (N_9634,N_9004,N_9050);
and U9635 (N_9635,N_9025,N_8694);
nor U9636 (N_9636,N_8706,N_8530);
nand U9637 (N_9637,N_9498,N_9474);
xnor U9638 (N_9638,N_8832,N_9485);
or U9639 (N_9639,N_8536,N_8465);
and U9640 (N_9640,N_9229,N_9309);
and U9641 (N_9641,N_9493,N_9473);
nor U9642 (N_9642,N_9210,N_9522);
and U9643 (N_9643,N_8416,N_9404);
or U9644 (N_9644,N_9383,N_8827);
nor U9645 (N_9645,N_9329,N_8707);
nand U9646 (N_9646,N_8733,N_8912);
nand U9647 (N_9647,N_8995,N_8840);
nand U9648 (N_9648,N_8761,N_9562);
nor U9649 (N_9649,N_9195,N_8855);
nor U9650 (N_9650,N_8400,N_8479);
and U9651 (N_9651,N_8409,N_9495);
xnor U9652 (N_9652,N_9228,N_8973);
or U9653 (N_9653,N_8877,N_8998);
and U9654 (N_9654,N_9084,N_8503);
and U9655 (N_9655,N_9267,N_8726);
nor U9656 (N_9656,N_9431,N_9410);
nor U9657 (N_9657,N_9298,N_9054);
nor U9658 (N_9658,N_9104,N_9006);
nand U9659 (N_9659,N_8440,N_8804);
and U9660 (N_9660,N_8792,N_8514);
or U9661 (N_9661,N_8829,N_9174);
and U9662 (N_9662,N_8445,N_9572);
or U9663 (N_9663,N_9282,N_9112);
or U9664 (N_9664,N_8508,N_8519);
xnor U9665 (N_9665,N_8455,N_8669);
xor U9666 (N_9666,N_9076,N_9408);
and U9667 (N_9667,N_8558,N_9041);
xor U9668 (N_9668,N_9484,N_8878);
and U9669 (N_9669,N_8556,N_9110);
nand U9670 (N_9670,N_8639,N_8787);
or U9671 (N_9671,N_8708,N_9578);
or U9672 (N_9672,N_8499,N_9542);
xor U9673 (N_9673,N_9245,N_9290);
xnor U9674 (N_9674,N_9160,N_8725);
and U9675 (N_9675,N_8560,N_9412);
nor U9676 (N_9676,N_8781,N_8576);
nand U9677 (N_9677,N_8498,N_8621);
and U9678 (N_9678,N_9478,N_9322);
and U9679 (N_9679,N_8846,N_8789);
nor U9680 (N_9680,N_8753,N_8994);
and U9681 (N_9681,N_9363,N_8464);
nor U9682 (N_9682,N_8977,N_8833);
nor U9683 (N_9683,N_8990,N_9307);
nand U9684 (N_9684,N_8537,N_9462);
or U9685 (N_9685,N_8486,N_8493);
or U9686 (N_9686,N_9081,N_9065);
nor U9687 (N_9687,N_9087,N_8422);
nand U9688 (N_9688,N_8822,N_9294);
or U9689 (N_9689,N_9543,N_8704);
or U9690 (N_9690,N_9005,N_8431);
or U9691 (N_9691,N_8768,N_8442);
or U9692 (N_9692,N_8677,N_9052);
xnor U9693 (N_9693,N_9028,N_8630);
or U9694 (N_9694,N_9598,N_8535);
and U9695 (N_9695,N_9502,N_9058);
or U9696 (N_9696,N_8853,N_9142);
or U9697 (N_9697,N_8593,N_9082);
and U9698 (N_9698,N_9221,N_8754);
xor U9699 (N_9699,N_9218,N_8579);
or U9700 (N_9700,N_9428,N_8627);
xnor U9701 (N_9701,N_9500,N_8469);
nor U9702 (N_9702,N_9036,N_8880);
or U9703 (N_9703,N_9092,N_9149);
xnor U9704 (N_9704,N_8577,N_9553);
and U9705 (N_9705,N_9447,N_9102);
nor U9706 (N_9706,N_9416,N_8848);
nor U9707 (N_9707,N_9143,N_9306);
or U9708 (N_9708,N_8700,N_9070);
nand U9709 (N_9709,N_9475,N_9073);
nor U9710 (N_9710,N_8901,N_8923);
nor U9711 (N_9711,N_9217,N_9336);
nand U9712 (N_9712,N_8613,N_9467);
xor U9713 (N_9713,N_8643,N_8949);
or U9714 (N_9714,N_8935,N_9439);
and U9715 (N_9715,N_8606,N_9513);
or U9716 (N_9716,N_9300,N_9321);
nand U9717 (N_9717,N_9171,N_9330);
and U9718 (N_9718,N_9154,N_8433);
nor U9719 (N_9719,N_9566,N_8759);
and U9720 (N_9720,N_9072,N_9549);
and U9721 (N_9721,N_9456,N_8441);
nor U9722 (N_9722,N_8838,N_8467);
nand U9723 (N_9723,N_8485,N_8659);
or U9724 (N_9724,N_8857,N_9044);
nor U9725 (N_9725,N_8911,N_9097);
and U9726 (N_9726,N_9095,N_8472);
nand U9727 (N_9727,N_8929,N_9320);
xnor U9728 (N_9728,N_9129,N_9545);
and U9729 (N_9729,N_9083,N_8760);
xor U9730 (N_9730,N_8797,N_8631);
and U9731 (N_9731,N_8763,N_9417);
nand U9732 (N_9732,N_9436,N_9359);
nand U9733 (N_9733,N_9172,N_8671);
nand U9734 (N_9734,N_8646,N_8854);
and U9735 (N_9735,N_9305,N_8404);
nand U9736 (N_9736,N_9398,N_9069);
and U9737 (N_9737,N_8735,N_9509);
or U9738 (N_9738,N_9373,N_9173);
nor U9739 (N_9739,N_9554,N_8748);
or U9740 (N_9740,N_8425,N_8664);
nor U9741 (N_9741,N_9506,N_9433);
xnor U9742 (N_9742,N_8428,N_8852);
or U9743 (N_9743,N_8858,N_9165);
nand U9744 (N_9744,N_8524,N_8612);
nor U9745 (N_9745,N_9411,N_9540);
nand U9746 (N_9746,N_8497,N_8954);
xnor U9747 (N_9747,N_8452,N_8842);
nand U9748 (N_9748,N_9492,N_8713);
or U9749 (N_9749,N_8583,N_8757);
nand U9750 (N_9750,N_8430,N_8476);
nor U9751 (N_9751,N_9369,N_8897);
and U9752 (N_9752,N_9538,N_9008);
nand U9753 (N_9753,N_9077,N_9343);
nand U9754 (N_9754,N_8682,N_9029);
and U9755 (N_9755,N_9575,N_8978);
and U9756 (N_9756,N_9454,N_9579);
nor U9757 (N_9757,N_9501,N_9504);
and U9758 (N_9758,N_9521,N_9197);
xor U9759 (N_9759,N_8515,N_9515);
and U9760 (N_9760,N_9444,N_9062);
xor U9761 (N_9761,N_9440,N_9269);
xnor U9762 (N_9762,N_9536,N_8420);
and U9763 (N_9763,N_8495,N_9213);
xnor U9764 (N_9764,N_8443,N_8689);
and U9765 (N_9765,N_8640,N_8699);
nor U9766 (N_9766,N_8471,N_8913);
nand U9767 (N_9767,N_8432,N_9013);
nand U9768 (N_9768,N_9586,N_9511);
or U9769 (N_9769,N_9237,N_8811);
nor U9770 (N_9770,N_8569,N_8951);
nand U9771 (N_9771,N_8976,N_8605);
xor U9772 (N_9772,N_8866,N_8936);
or U9773 (N_9773,N_8925,N_8948);
xor U9774 (N_9774,N_8538,N_8403);
or U9775 (N_9775,N_8657,N_8642);
and U9776 (N_9776,N_8667,N_9266);
and U9777 (N_9777,N_8672,N_8969);
xnor U9778 (N_9778,N_9313,N_8819);
xnor U9779 (N_9779,N_8552,N_8889);
and U9780 (N_9780,N_9255,N_9466);
xnor U9781 (N_9781,N_8737,N_9120);
or U9782 (N_9782,N_8893,N_9164);
nor U9783 (N_9783,N_8739,N_9386);
or U9784 (N_9784,N_9333,N_8744);
nor U9785 (N_9785,N_8609,N_8419);
nor U9786 (N_9786,N_9361,N_9224);
nand U9787 (N_9787,N_9022,N_8685);
nand U9788 (N_9788,N_9158,N_9001);
xnor U9789 (N_9789,N_8963,N_8810);
xnor U9790 (N_9790,N_8686,N_9093);
nand U9791 (N_9791,N_8967,N_8899);
nand U9792 (N_9792,N_9130,N_9242);
nand U9793 (N_9793,N_9175,N_8553);
nor U9794 (N_9794,N_8587,N_9452);
or U9795 (N_9795,N_8695,N_8917);
xnor U9796 (N_9796,N_8421,N_8806);
nor U9797 (N_9797,N_9319,N_9079);
or U9798 (N_9798,N_8405,N_8534);
nand U9799 (N_9799,N_9257,N_9516);
nor U9800 (N_9800,N_8598,N_8635);
nand U9801 (N_9801,N_8462,N_8908);
nor U9802 (N_9802,N_9381,N_8510);
or U9803 (N_9803,N_8719,N_9252);
or U9804 (N_9804,N_9156,N_9459);
and U9805 (N_9805,N_8520,N_8983);
nor U9806 (N_9806,N_9375,N_9096);
nand U9807 (N_9807,N_9365,N_9114);
or U9808 (N_9808,N_9067,N_9275);
and U9809 (N_9809,N_9030,N_8703);
nor U9810 (N_9810,N_9358,N_8716);
and U9811 (N_9811,N_8996,N_8414);
xnor U9812 (N_9812,N_8888,N_8803);
and U9813 (N_9813,N_8919,N_8999);
xor U9814 (N_9814,N_8974,N_8603);
or U9815 (N_9815,N_9370,N_8769);
nand U9816 (N_9816,N_8815,N_9251);
nand U9817 (N_9817,N_9212,N_9399);
nor U9818 (N_9818,N_9366,N_9061);
nand U9819 (N_9819,N_8860,N_8937);
xnor U9820 (N_9820,N_9285,N_8454);
nand U9821 (N_9821,N_8824,N_9244);
nor U9822 (N_9822,N_9558,N_9227);
xor U9823 (N_9823,N_8764,N_8933);
nor U9824 (N_9824,N_9089,N_9510);
xnor U9825 (N_9825,N_8729,N_9397);
nand U9826 (N_9826,N_8828,N_8710);
and U9827 (N_9827,N_8542,N_8525);
or U9828 (N_9828,N_8683,N_9348);
nand U9829 (N_9829,N_9388,N_8952);
and U9830 (N_9830,N_9126,N_8745);
xor U9831 (N_9831,N_8450,N_8545);
or U9832 (N_9832,N_8799,N_9098);
nand U9833 (N_9833,N_8565,N_9565);
or U9834 (N_9834,N_8453,N_8741);
xnor U9835 (N_9835,N_8850,N_9512);
nor U9836 (N_9836,N_9133,N_9147);
xor U9837 (N_9837,N_9589,N_9563);
and U9838 (N_9838,N_9481,N_9378);
nor U9839 (N_9839,N_8932,N_9207);
and U9840 (N_9840,N_9405,N_8411);
nor U9841 (N_9841,N_8796,N_9470);
or U9842 (N_9842,N_8993,N_9380);
and U9843 (N_9843,N_9457,N_8924);
nand U9844 (N_9844,N_9243,N_9219);
or U9845 (N_9845,N_9374,N_8632);
nand U9846 (N_9846,N_9256,N_9135);
or U9847 (N_9847,N_8580,N_9537);
nor U9848 (N_9848,N_9489,N_9534);
nor U9849 (N_9849,N_9037,N_9503);
nand U9850 (N_9850,N_9203,N_8883);
nor U9851 (N_9851,N_8596,N_8805);
or U9852 (N_9852,N_9134,N_8834);
nor U9853 (N_9853,N_9150,N_9310);
nand U9854 (N_9854,N_9232,N_9101);
and U9855 (N_9855,N_8956,N_8915);
nor U9856 (N_9856,N_9592,N_9314);
and U9857 (N_9857,N_8724,N_8563);
and U9858 (N_9858,N_9420,N_8885);
or U9859 (N_9859,N_8849,N_8979);
nor U9860 (N_9860,N_9194,N_9587);
or U9861 (N_9861,N_8655,N_8909);
and U9862 (N_9862,N_9240,N_9051);
and U9863 (N_9863,N_9220,N_9038);
nor U9864 (N_9864,N_9132,N_9570);
nor U9865 (N_9865,N_8869,N_9024);
or U9866 (N_9866,N_8892,N_9488);
xor U9867 (N_9867,N_9302,N_9349);
nor U9868 (N_9868,N_8712,N_8448);
nor U9869 (N_9869,N_8673,N_9225);
xnor U9870 (N_9870,N_8597,N_8647);
xor U9871 (N_9871,N_9550,N_9469);
nand U9872 (N_9872,N_8417,N_9458);
or U9873 (N_9873,N_8548,N_8589);
or U9874 (N_9874,N_8900,N_9140);
xor U9875 (N_9875,N_9119,N_8876);
nor U9876 (N_9876,N_8489,N_8406);
xor U9877 (N_9877,N_8697,N_9497);
xnor U9878 (N_9878,N_8423,N_8491);
nand U9879 (N_9879,N_8732,N_8964);
or U9880 (N_9880,N_8412,N_9331);
nor U9881 (N_9881,N_9163,N_9196);
xnor U9882 (N_9882,N_8955,N_9190);
nand U9883 (N_9883,N_9259,N_9226);
nand U9884 (N_9884,N_9327,N_9393);
xor U9885 (N_9885,N_9045,N_9527);
xor U9886 (N_9886,N_8870,N_8959);
or U9887 (N_9887,N_8439,N_8567);
and U9888 (N_9888,N_8595,N_8528);
nand U9889 (N_9889,N_8641,N_8928);
nand U9890 (N_9890,N_9368,N_9429);
xor U9891 (N_9891,N_9274,N_9351);
or U9892 (N_9892,N_8991,N_9552);
nand U9893 (N_9893,N_8539,N_8687);
nand U9894 (N_9894,N_8782,N_9169);
or U9895 (N_9895,N_9146,N_8727);
or U9896 (N_9896,N_8943,N_8592);
xnor U9897 (N_9897,N_9170,N_9209);
nor U9898 (N_9898,N_9247,N_8920);
xnor U9899 (N_9899,N_8575,N_9569);
or U9900 (N_9900,N_9049,N_9317);
or U9901 (N_9901,N_9573,N_8634);
or U9902 (N_9902,N_9364,N_9222);
nor U9903 (N_9903,N_9128,N_8823);
nand U9904 (N_9904,N_8875,N_9443);
and U9905 (N_9905,N_8960,N_8831);
xnor U9906 (N_9906,N_9406,N_9020);
or U9907 (N_9907,N_8633,N_9326);
xnor U9908 (N_9908,N_8776,N_8461);
and U9909 (N_9909,N_8590,N_9352);
xnor U9910 (N_9910,N_8675,N_8701);
and U9911 (N_9911,N_9032,N_9031);
nand U9912 (N_9912,N_8826,N_9483);
nor U9913 (N_9913,N_8813,N_9528);
xnor U9914 (N_9914,N_9441,N_9585);
nor U9915 (N_9915,N_8692,N_8856);
nor U9916 (N_9916,N_8446,N_8814);
or U9917 (N_9917,N_9453,N_9402);
nand U9918 (N_9918,N_8944,N_8551);
nand U9919 (N_9919,N_9125,N_9353);
nand U9920 (N_9920,N_8494,N_8946);
and U9921 (N_9921,N_8847,N_9339);
nand U9922 (N_9922,N_8961,N_8460);
xor U9923 (N_9923,N_9490,N_9448);
and U9924 (N_9924,N_9253,N_9544);
and U9925 (N_9925,N_8985,N_8786);
nand U9926 (N_9926,N_8459,N_8424);
and U9927 (N_9927,N_9152,N_8788);
or U9928 (N_9928,N_8890,N_8617);
xor U9929 (N_9929,N_8561,N_8722);
and U9930 (N_9930,N_8550,N_9308);
nand U9931 (N_9931,N_8668,N_8865);
nand U9932 (N_9932,N_8426,N_9346);
or U9933 (N_9933,N_8625,N_9035);
nor U9934 (N_9934,N_9019,N_8622);
xor U9935 (N_9935,N_9533,N_9561);
and U9936 (N_9936,N_8859,N_9063);
nand U9937 (N_9937,N_9201,N_9299);
xor U9938 (N_9938,N_8772,N_8825);
nor U9939 (N_9939,N_8526,N_9324);
nand U9940 (N_9940,N_8907,N_9548);
and U9941 (N_9941,N_8968,N_8540);
or U9942 (N_9942,N_9099,N_9292);
and U9943 (N_9943,N_9479,N_8541);
xor U9944 (N_9944,N_8987,N_8555);
nor U9945 (N_9945,N_8918,N_9591);
nand U9946 (N_9946,N_9151,N_9139);
xor U9947 (N_9947,N_8965,N_9239);
and U9948 (N_9948,N_8896,N_8544);
nand U9949 (N_9949,N_8749,N_8506);
nand U9950 (N_9950,N_9507,N_9376);
nor U9951 (N_9951,N_9480,N_9223);
nor U9952 (N_9952,N_9461,N_9118);
nand U9953 (N_9953,N_9360,N_9234);
xor U9954 (N_9954,N_8658,N_8839);
nand U9955 (N_9955,N_9124,N_8578);
nor U9956 (N_9956,N_8972,N_9465);
or U9957 (N_9957,N_8941,N_8921);
nand U9958 (N_9958,N_8938,N_9047);
or U9959 (N_9959,N_9176,N_9254);
nor U9960 (N_9960,N_8554,N_9159);
or U9961 (N_9961,N_8730,N_9551);
or U9962 (N_9962,N_8619,N_9471);
and U9963 (N_9963,N_8678,N_8942);
nor U9964 (N_9964,N_8415,N_8820);
xnor U9965 (N_9965,N_9241,N_9074);
and U9966 (N_9966,N_8652,N_8705);
nor U9967 (N_9967,N_8649,N_9046);
nand U9968 (N_9968,N_9117,N_9574);
or U9969 (N_9969,N_9085,N_8594);
or U9970 (N_9970,N_8662,N_9568);
nor U9971 (N_9971,N_9188,N_9168);
or U9972 (N_9972,N_8475,N_8436);
nor U9973 (N_9973,N_9422,N_8573);
and U9974 (N_9974,N_9367,N_8767);
xor U9975 (N_9975,N_8926,N_8777);
xnor U9976 (N_9976,N_8568,N_8636);
nand U9977 (N_9977,N_8591,N_9508);
nor U9978 (N_9978,N_9250,N_8457);
and U9979 (N_9979,N_9057,N_8775);
or U9980 (N_9980,N_9328,N_8413);
nor U9981 (N_9981,N_9179,N_8614);
and U9982 (N_9982,N_9409,N_9377);
or U9983 (N_9983,N_9582,N_8435);
or U9984 (N_9984,N_9555,N_9425);
and U9985 (N_9985,N_8997,N_9027);
xor U9986 (N_9986,N_9446,N_8798);
or U9987 (N_9987,N_9419,N_8721);
and U9988 (N_9988,N_9583,N_8743);
and U9989 (N_9989,N_9039,N_9524);
nand U9990 (N_9990,N_9599,N_9012);
nor U9991 (N_9991,N_9021,N_8894);
nand U9992 (N_9992,N_9546,N_8751);
nor U9993 (N_9993,N_9105,N_9449);
and U9994 (N_9994,N_9034,N_8736);
nand U9995 (N_9995,N_8886,N_9597);
nor U9996 (N_9996,N_9557,N_9316);
nand U9997 (N_9997,N_8882,N_8532);
and U9998 (N_9998,N_8601,N_9260);
xnor U9999 (N_9999,N_9345,N_9181);
nor U10000 (N_10000,N_9136,N_9535);
nand U10001 (N_10001,N_8549,N_8910);
nor U10002 (N_10002,N_9111,N_9166);
and U10003 (N_10003,N_9560,N_9424);
xor U10004 (N_10004,N_9400,N_9262);
and U10005 (N_10005,N_8463,N_9438);
or U10006 (N_10006,N_8970,N_8620);
nand U10007 (N_10007,N_9434,N_8670);
nor U10008 (N_10008,N_8879,N_9468);
nand U10009 (N_10009,N_9463,N_8914);
nand U10010 (N_10010,N_8778,N_9427);
nand U10011 (N_10011,N_8666,N_9184);
xnor U10012 (N_10012,N_9182,N_9407);
nand U10013 (N_10013,N_8992,N_9335);
or U10014 (N_10014,N_9115,N_9340);
or U10015 (N_10015,N_9198,N_8711);
xor U10016 (N_10016,N_8586,N_8864);
and U10017 (N_10017,N_8758,N_8843);
xnor U10018 (N_10018,N_8518,N_8868);
xor U10019 (N_10019,N_8447,N_9078);
nand U10020 (N_10020,N_8779,N_8790);
and U10021 (N_10021,N_9514,N_9155);
nor U10022 (N_10022,N_9178,N_8728);
or U10023 (N_10023,N_9211,N_8971);
xor U10024 (N_10024,N_9088,N_9185);
nand U10025 (N_10025,N_8709,N_9435);
or U10026 (N_10026,N_9216,N_8484);
nor U10027 (N_10027,N_8891,N_9148);
nand U10028 (N_10028,N_8756,N_8698);
and U10029 (N_10029,N_8680,N_8945);
or U10030 (N_10030,N_9215,N_8650);
and U10031 (N_10031,N_9325,N_9531);
xor U10032 (N_10032,N_8505,N_9186);
or U10033 (N_10033,N_9281,N_8458);
xnor U10034 (N_10034,N_8504,N_8610);
nand U10035 (N_10035,N_8509,N_9167);
nor U10036 (N_10036,N_9265,N_8903);
nor U10037 (N_10037,N_9571,N_9137);
nand U10038 (N_10038,N_9014,N_9270);
nor U10039 (N_10039,N_8800,N_9520);
or U10040 (N_10040,N_8784,N_9385);
or U10041 (N_10041,N_8582,N_9121);
nand U10042 (N_10042,N_9391,N_8674);
or U10043 (N_10043,N_9432,N_9080);
xor U10044 (N_10044,N_8645,N_8638);
or U10045 (N_10045,N_9109,N_9517);
xnor U10046 (N_10046,N_8696,N_8470);
xor U10047 (N_10047,N_9199,N_9567);
and U10048 (N_10048,N_8615,N_8873);
and U10049 (N_10049,N_9539,N_8557);
and U10050 (N_10050,N_9284,N_8830);
nor U10051 (N_10051,N_8988,N_9055);
or U10052 (N_10052,N_8477,N_9499);
xor U10053 (N_10053,N_8738,N_8427);
xor U10054 (N_10054,N_8906,N_9396);
xnor U10055 (N_10055,N_9382,N_8407);
xnor U10056 (N_10056,N_9301,N_8785);
or U10057 (N_10057,N_9235,N_9423);
and U10058 (N_10058,N_8665,N_8660);
xnor U10059 (N_10059,N_8608,N_9162);
nand U10060 (N_10060,N_8718,N_9529);
or U10061 (N_10061,N_8602,N_8957);
nand U10062 (N_10062,N_9204,N_9390);
and U10063 (N_10063,N_9334,N_8817);
or U10064 (N_10064,N_9594,N_8521);
xor U10065 (N_10065,N_9248,N_9384);
nand U10066 (N_10066,N_9401,N_8585);
xor U10067 (N_10067,N_8773,N_9043);
nand U10068 (N_10068,N_8953,N_8931);
and U10069 (N_10069,N_8571,N_8401);
or U10070 (N_10070,N_8507,N_8482);
xnor U10071 (N_10071,N_9007,N_9015);
or U10072 (N_10072,N_9491,N_8581);
and U10073 (N_10073,N_8691,N_8794);
or U10074 (N_10074,N_9362,N_8559);
nand U10075 (N_10075,N_8747,N_9564);
nor U10076 (N_10076,N_8651,N_9056);
or U10077 (N_10077,N_8429,N_8975);
xor U10078 (N_10078,N_9426,N_9494);
nor U10079 (N_10079,N_9337,N_9487);
nand U10080 (N_10080,N_9291,N_8473);
nor U10081 (N_10081,N_8881,N_9091);
or U10082 (N_10082,N_9261,N_9177);
nand U10083 (N_10083,N_9584,N_8566);
or U10084 (N_10084,N_9541,N_8982);
xor U10085 (N_10085,N_8808,N_8895);
or U10086 (N_10086,N_8930,N_8904);
xnor U10087 (N_10087,N_8783,N_9205);
nand U10088 (N_10088,N_9026,N_8564);
or U10089 (N_10089,N_8962,N_8600);
or U10090 (N_10090,N_8654,N_8809);
or U10091 (N_10091,N_8527,N_9122);
and U10092 (N_10092,N_8807,N_9258);
nand U10093 (N_10093,N_9161,N_8688);
nand U10094 (N_10094,N_8841,N_9094);
or U10095 (N_10095,N_8750,N_8746);
xnor U10096 (N_10096,N_8531,N_9053);
xor U10097 (N_10097,N_8812,N_8434);
and U10098 (N_10098,N_9593,N_8492);
xor U10099 (N_10099,N_9437,N_9033);
and U10100 (N_10100,N_8616,N_9127);
xor U10101 (N_10101,N_9295,N_9113);
and U10102 (N_10102,N_9318,N_9464);
xor U10103 (N_10103,N_9413,N_9312);
or U10104 (N_10104,N_9415,N_9323);
or U10105 (N_10105,N_8940,N_8588);
xor U10106 (N_10106,N_8916,N_9233);
and U10107 (N_10107,N_9392,N_8947);
xnor U10108 (N_10108,N_9477,N_8410);
nor U10109 (N_10109,N_9354,N_8653);
nor U10110 (N_10110,N_9279,N_9556);
xor U10111 (N_10111,N_9315,N_9193);
or U10112 (N_10112,N_9230,N_8516);
or U10113 (N_10113,N_9372,N_9486);
nand U10114 (N_10114,N_8765,N_9208);
xnor U10115 (N_10115,N_8755,N_8795);
or U10116 (N_10116,N_9272,N_8702);
and U10117 (N_10117,N_8981,N_8898);
nand U10118 (N_10118,N_9011,N_8723);
and U10119 (N_10119,N_9086,N_8466);
nor U10120 (N_10120,N_9141,N_8862);
or U10121 (N_10121,N_9183,N_9482);
and U10122 (N_10122,N_9276,N_9347);
and U10123 (N_10123,N_9145,N_9576);
nor U10124 (N_10124,N_9138,N_9371);
or U10125 (N_10125,N_8861,N_9547);
or U10126 (N_10126,N_9287,N_8845);
nor U10127 (N_10127,N_8816,N_9379);
nand U10128 (N_10128,N_8774,N_9451);
xor U10129 (N_10129,N_9003,N_8762);
or U10130 (N_10130,N_9518,N_9580);
or U10131 (N_10131,N_9293,N_8522);
or U10132 (N_10132,N_8927,N_9002);
and U10133 (N_10133,N_9108,N_8644);
and U10134 (N_10134,N_9180,N_9023);
nand U10135 (N_10135,N_9106,N_8742);
nand U10136 (N_10136,N_8629,N_9476);
or U10137 (N_10137,N_9350,N_9191);
nor U10138 (N_10138,N_8871,N_9068);
or U10139 (N_10139,N_9040,N_9192);
nor U10140 (N_10140,N_8934,N_9581);
or U10141 (N_10141,N_8449,N_9187);
and U10142 (N_10142,N_8437,N_8496);
nand U10143 (N_10143,N_9421,N_8611);
nor U10144 (N_10144,N_9332,N_8771);
nor U10145 (N_10145,N_8844,N_8624);
nand U10146 (N_10146,N_8480,N_9304);
nand U10147 (N_10147,N_9271,N_9071);
xnor U10148 (N_10148,N_8501,N_9048);
xor U10149 (N_10149,N_8851,N_8547);
xor U10150 (N_10150,N_8474,N_9344);
nor U10151 (N_10151,N_8902,N_9455);
xor U10152 (N_10152,N_8648,N_8867);
xnor U10153 (N_10153,N_8740,N_9206);
and U10154 (N_10154,N_8958,N_8734);
xor U10155 (N_10155,N_9189,N_8821);
and U10156 (N_10156,N_8818,N_8628);
nor U10157 (N_10157,N_8681,N_9357);
or U10158 (N_10158,N_8402,N_9394);
nand U10159 (N_10159,N_9000,N_8408);
xnor U10160 (N_10160,N_8418,N_8766);
or U10161 (N_10161,N_8690,N_9107);
xnor U10162 (N_10162,N_9283,N_8584);
xnor U10163 (N_10163,N_9296,N_8989);
nor U10164 (N_10164,N_9414,N_9060);
or U10165 (N_10165,N_9297,N_8604);
nand U10166 (N_10166,N_8836,N_8481);
nand U10167 (N_10167,N_8533,N_8980);
xnor U10168 (N_10168,N_9103,N_9355);
and U10169 (N_10169,N_8529,N_8512);
or U10170 (N_10170,N_8513,N_8438);
nand U10171 (N_10171,N_8478,N_9273);
or U10172 (N_10172,N_8488,N_8837);
or U10173 (N_10173,N_9018,N_9588);
nand U10174 (N_10174,N_9236,N_9530);
nor U10175 (N_10175,N_9289,N_9123);
or U10176 (N_10176,N_8884,N_9200);
xnor U10177 (N_10177,N_9403,N_8874);
xor U10178 (N_10178,N_8793,N_9595);
xor U10179 (N_10179,N_8637,N_9532);
xor U10180 (N_10180,N_9075,N_8863);
nor U10181 (N_10181,N_8801,N_9157);
nor U10182 (N_10182,N_9286,N_8456);
or U10183 (N_10183,N_9059,N_9389);
nand U10184 (N_10184,N_8468,N_8451);
and U10185 (N_10185,N_9246,N_9596);
nor U10186 (N_10186,N_8922,N_9445);
nor U10187 (N_10187,N_9009,N_8717);
xnor U10188 (N_10188,N_8714,N_8872);
and U10189 (N_10189,N_9430,N_9042);
or U10190 (N_10190,N_9590,N_8663);
or U10191 (N_10191,N_9311,N_9238);
nand U10192 (N_10192,N_9280,N_9559);
or U10193 (N_10193,N_8984,N_9303);
xor U10194 (N_10194,N_9450,N_8599);
xor U10195 (N_10195,N_8572,N_9263);
or U10196 (N_10196,N_8626,N_9387);
or U10197 (N_10197,N_9249,N_9525);
nor U10198 (N_10198,N_8623,N_9356);
or U10199 (N_10199,N_8986,N_8802);
xnor U10200 (N_10200,N_8821,N_8457);
nor U10201 (N_10201,N_9458,N_8482);
and U10202 (N_10202,N_9351,N_8767);
or U10203 (N_10203,N_9493,N_9101);
and U10204 (N_10204,N_8861,N_9480);
nor U10205 (N_10205,N_9523,N_9305);
nor U10206 (N_10206,N_8724,N_9086);
xnor U10207 (N_10207,N_9546,N_8792);
and U10208 (N_10208,N_8763,N_8703);
and U10209 (N_10209,N_9486,N_9193);
and U10210 (N_10210,N_9360,N_8790);
nand U10211 (N_10211,N_8505,N_8778);
or U10212 (N_10212,N_8438,N_9417);
xor U10213 (N_10213,N_9494,N_8726);
nand U10214 (N_10214,N_8889,N_9422);
xor U10215 (N_10215,N_9312,N_9363);
nor U10216 (N_10216,N_9304,N_8623);
or U10217 (N_10217,N_9332,N_8438);
and U10218 (N_10218,N_8464,N_9093);
and U10219 (N_10219,N_9017,N_8409);
or U10220 (N_10220,N_8451,N_8630);
nand U10221 (N_10221,N_9445,N_9483);
and U10222 (N_10222,N_9208,N_8460);
and U10223 (N_10223,N_9147,N_8716);
nor U10224 (N_10224,N_9001,N_8641);
or U10225 (N_10225,N_9273,N_8710);
xor U10226 (N_10226,N_9084,N_8828);
nand U10227 (N_10227,N_9551,N_8614);
xnor U10228 (N_10228,N_9485,N_8975);
nand U10229 (N_10229,N_8569,N_8930);
xnor U10230 (N_10230,N_9194,N_9303);
nor U10231 (N_10231,N_8605,N_9516);
or U10232 (N_10232,N_8679,N_8966);
nor U10233 (N_10233,N_9084,N_9302);
or U10234 (N_10234,N_8751,N_9177);
xnor U10235 (N_10235,N_9018,N_8926);
or U10236 (N_10236,N_9340,N_9537);
nor U10237 (N_10237,N_8944,N_9147);
xor U10238 (N_10238,N_9232,N_9143);
or U10239 (N_10239,N_9165,N_8518);
and U10240 (N_10240,N_9563,N_9015);
nand U10241 (N_10241,N_8792,N_8420);
nor U10242 (N_10242,N_9099,N_9098);
nor U10243 (N_10243,N_8776,N_8570);
or U10244 (N_10244,N_8410,N_9413);
nor U10245 (N_10245,N_8739,N_9396);
nor U10246 (N_10246,N_8748,N_9260);
or U10247 (N_10247,N_8842,N_9033);
and U10248 (N_10248,N_9559,N_9379);
or U10249 (N_10249,N_9269,N_9157);
or U10250 (N_10250,N_8848,N_9503);
nand U10251 (N_10251,N_9314,N_9524);
xor U10252 (N_10252,N_9181,N_8814);
xnor U10253 (N_10253,N_9286,N_9391);
and U10254 (N_10254,N_8976,N_9360);
nor U10255 (N_10255,N_9563,N_8978);
or U10256 (N_10256,N_8683,N_8788);
nor U10257 (N_10257,N_8539,N_8586);
nand U10258 (N_10258,N_8517,N_8869);
nor U10259 (N_10259,N_8571,N_9059);
and U10260 (N_10260,N_8967,N_8848);
nor U10261 (N_10261,N_9275,N_8827);
xnor U10262 (N_10262,N_8632,N_9582);
nor U10263 (N_10263,N_8417,N_9115);
or U10264 (N_10264,N_8643,N_8536);
nor U10265 (N_10265,N_8549,N_9328);
or U10266 (N_10266,N_9504,N_9143);
xor U10267 (N_10267,N_8576,N_9125);
and U10268 (N_10268,N_9026,N_9032);
nor U10269 (N_10269,N_8789,N_9178);
and U10270 (N_10270,N_8644,N_9101);
and U10271 (N_10271,N_9479,N_8482);
xor U10272 (N_10272,N_9086,N_9523);
xnor U10273 (N_10273,N_8721,N_9136);
or U10274 (N_10274,N_9524,N_9112);
nand U10275 (N_10275,N_8836,N_9370);
nor U10276 (N_10276,N_8459,N_8613);
xnor U10277 (N_10277,N_8698,N_8675);
and U10278 (N_10278,N_9136,N_9133);
nor U10279 (N_10279,N_9575,N_9292);
and U10280 (N_10280,N_9593,N_9319);
xnor U10281 (N_10281,N_8796,N_8431);
and U10282 (N_10282,N_9211,N_9276);
or U10283 (N_10283,N_9284,N_8442);
nand U10284 (N_10284,N_8405,N_8783);
or U10285 (N_10285,N_9106,N_9498);
nand U10286 (N_10286,N_9434,N_9014);
or U10287 (N_10287,N_9400,N_9084);
or U10288 (N_10288,N_8517,N_9079);
nand U10289 (N_10289,N_8619,N_9579);
nand U10290 (N_10290,N_9570,N_8895);
xnor U10291 (N_10291,N_9189,N_9180);
xnor U10292 (N_10292,N_8652,N_9131);
nand U10293 (N_10293,N_8630,N_8991);
nor U10294 (N_10294,N_8436,N_9082);
nand U10295 (N_10295,N_9423,N_8755);
and U10296 (N_10296,N_9056,N_8751);
and U10297 (N_10297,N_8496,N_9512);
nor U10298 (N_10298,N_9010,N_9535);
xnor U10299 (N_10299,N_9353,N_8523);
nor U10300 (N_10300,N_9364,N_8973);
nor U10301 (N_10301,N_9598,N_9302);
or U10302 (N_10302,N_9412,N_9212);
xnor U10303 (N_10303,N_9054,N_8467);
nand U10304 (N_10304,N_9554,N_8513);
nand U10305 (N_10305,N_8856,N_9398);
and U10306 (N_10306,N_8525,N_8719);
and U10307 (N_10307,N_9536,N_9399);
or U10308 (N_10308,N_9155,N_9443);
nor U10309 (N_10309,N_8414,N_9000);
xor U10310 (N_10310,N_9285,N_8458);
or U10311 (N_10311,N_8513,N_9111);
nor U10312 (N_10312,N_9075,N_8780);
or U10313 (N_10313,N_9103,N_8605);
and U10314 (N_10314,N_8759,N_8665);
and U10315 (N_10315,N_9253,N_8863);
nor U10316 (N_10316,N_8472,N_9460);
nand U10317 (N_10317,N_8451,N_9319);
nor U10318 (N_10318,N_8852,N_9167);
nand U10319 (N_10319,N_8487,N_9436);
nor U10320 (N_10320,N_8451,N_9117);
and U10321 (N_10321,N_8730,N_9218);
nor U10322 (N_10322,N_8875,N_9114);
and U10323 (N_10323,N_9041,N_8829);
and U10324 (N_10324,N_9556,N_9354);
or U10325 (N_10325,N_8957,N_8927);
nand U10326 (N_10326,N_8868,N_9019);
or U10327 (N_10327,N_9430,N_9253);
and U10328 (N_10328,N_8465,N_9151);
nor U10329 (N_10329,N_9270,N_9174);
or U10330 (N_10330,N_8775,N_9142);
nor U10331 (N_10331,N_8694,N_8987);
and U10332 (N_10332,N_8957,N_9021);
nand U10333 (N_10333,N_8539,N_9500);
or U10334 (N_10334,N_9205,N_9046);
xnor U10335 (N_10335,N_9113,N_8969);
nand U10336 (N_10336,N_9137,N_9116);
nor U10337 (N_10337,N_9333,N_9381);
nand U10338 (N_10338,N_8822,N_9550);
or U10339 (N_10339,N_9201,N_8637);
or U10340 (N_10340,N_8546,N_9404);
nand U10341 (N_10341,N_8881,N_9190);
nand U10342 (N_10342,N_9446,N_9022);
and U10343 (N_10343,N_9169,N_8780);
xor U10344 (N_10344,N_9365,N_9482);
nor U10345 (N_10345,N_8430,N_8634);
or U10346 (N_10346,N_8527,N_9342);
or U10347 (N_10347,N_9269,N_9228);
or U10348 (N_10348,N_8645,N_8756);
or U10349 (N_10349,N_9142,N_8661);
nand U10350 (N_10350,N_8984,N_8797);
nand U10351 (N_10351,N_8965,N_9162);
and U10352 (N_10352,N_8912,N_8830);
and U10353 (N_10353,N_9070,N_8696);
xnor U10354 (N_10354,N_8748,N_8895);
xor U10355 (N_10355,N_9589,N_8482);
nand U10356 (N_10356,N_9195,N_9079);
nor U10357 (N_10357,N_8877,N_9273);
nor U10358 (N_10358,N_9087,N_9364);
or U10359 (N_10359,N_8742,N_9162);
xor U10360 (N_10360,N_9432,N_8937);
nor U10361 (N_10361,N_8727,N_9401);
xor U10362 (N_10362,N_9467,N_8860);
nor U10363 (N_10363,N_8583,N_8417);
nand U10364 (N_10364,N_9585,N_9047);
and U10365 (N_10365,N_9199,N_9206);
or U10366 (N_10366,N_8401,N_9077);
xnor U10367 (N_10367,N_8771,N_8405);
and U10368 (N_10368,N_9459,N_8702);
nand U10369 (N_10369,N_8745,N_8469);
and U10370 (N_10370,N_8875,N_8643);
nand U10371 (N_10371,N_9379,N_8546);
and U10372 (N_10372,N_8432,N_9572);
xor U10373 (N_10373,N_8997,N_8571);
and U10374 (N_10374,N_9335,N_8957);
or U10375 (N_10375,N_8476,N_8661);
nor U10376 (N_10376,N_9520,N_8660);
nand U10377 (N_10377,N_9415,N_8836);
nand U10378 (N_10378,N_8867,N_9290);
or U10379 (N_10379,N_9273,N_9178);
and U10380 (N_10380,N_8831,N_9550);
and U10381 (N_10381,N_8924,N_9094);
or U10382 (N_10382,N_8535,N_9362);
and U10383 (N_10383,N_8907,N_8747);
nor U10384 (N_10384,N_9242,N_8968);
and U10385 (N_10385,N_9587,N_8713);
or U10386 (N_10386,N_8851,N_8401);
nor U10387 (N_10387,N_8655,N_9338);
nand U10388 (N_10388,N_8710,N_9192);
and U10389 (N_10389,N_8627,N_8811);
nor U10390 (N_10390,N_9526,N_8697);
and U10391 (N_10391,N_9038,N_9504);
and U10392 (N_10392,N_8544,N_9516);
xnor U10393 (N_10393,N_9111,N_8461);
xnor U10394 (N_10394,N_9417,N_9562);
or U10395 (N_10395,N_8797,N_9365);
or U10396 (N_10396,N_8965,N_9331);
and U10397 (N_10397,N_8467,N_8826);
or U10398 (N_10398,N_9558,N_9104);
or U10399 (N_10399,N_9306,N_8795);
nand U10400 (N_10400,N_8660,N_9115);
nor U10401 (N_10401,N_9060,N_8693);
xnor U10402 (N_10402,N_8802,N_9425);
and U10403 (N_10403,N_8702,N_8708);
and U10404 (N_10404,N_8641,N_8515);
nand U10405 (N_10405,N_8684,N_9416);
nand U10406 (N_10406,N_9048,N_9470);
and U10407 (N_10407,N_8554,N_9431);
xor U10408 (N_10408,N_9309,N_9522);
xor U10409 (N_10409,N_8775,N_8650);
and U10410 (N_10410,N_9525,N_8926);
and U10411 (N_10411,N_9330,N_8420);
nor U10412 (N_10412,N_8712,N_9442);
and U10413 (N_10413,N_8910,N_9291);
nor U10414 (N_10414,N_9206,N_8790);
nand U10415 (N_10415,N_8560,N_8571);
nand U10416 (N_10416,N_8820,N_9485);
nand U10417 (N_10417,N_9474,N_9456);
and U10418 (N_10418,N_8804,N_9358);
nor U10419 (N_10419,N_9009,N_9108);
nand U10420 (N_10420,N_8508,N_9326);
xor U10421 (N_10421,N_8736,N_9005);
nor U10422 (N_10422,N_8668,N_9494);
nand U10423 (N_10423,N_9325,N_8908);
nand U10424 (N_10424,N_8913,N_8585);
or U10425 (N_10425,N_8766,N_8672);
nor U10426 (N_10426,N_9362,N_9242);
and U10427 (N_10427,N_8691,N_9507);
and U10428 (N_10428,N_9048,N_9427);
nor U10429 (N_10429,N_8772,N_9029);
nor U10430 (N_10430,N_8669,N_9480);
nor U10431 (N_10431,N_9156,N_9090);
or U10432 (N_10432,N_9332,N_9142);
nor U10433 (N_10433,N_9341,N_9039);
nand U10434 (N_10434,N_9492,N_9143);
nor U10435 (N_10435,N_9215,N_9411);
xor U10436 (N_10436,N_8751,N_8988);
nand U10437 (N_10437,N_8764,N_8591);
and U10438 (N_10438,N_8530,N_9356);
and U10439 (N_10439,N_9040,N_8839);
or U10440 (N_10440,N_9474,N_8692);
xnor U10441 (N_10441,N_8468,N_9028);
nor U10442 (N_10442,N_8515,N_8720);
nor U10443 (N_10443,N_9300,N_9191);
or U10444 (N_10444,N_8828,N_8600);
and U10445 (N_10445,N_9449,N_8856);
nor U10446 (N_10446,N_8671,N_8684);
or U10447 (N_10447,N_8940,N_8924);
nand U10448 (N_10448,N_9350,N_9083);
nor U10449 (N_10449,N_8546,N_8436);
nor U10450 (N_10450,N_8402,N_8731);
xnor U10451 (N_10451,N_8521,N_8789);
nand U10452 (N_10452,N_8455,N_8921);
and U10453 (N_10453,N_9358,N_8840);
nand U10454 (N_10454,N_8830,N_8730);
or U10455 (N_10455,N_9279,N_9205);
and U10456 (N_10456,N_8449,N_8724);
nand U10457 (N_10457,N_8712,N_8832);
and U10458 (N_10458,N_8890,N_9148);
and U10459 (N_10459,N_8616,N_8660);
xnor U10460 (N_10460,N_9497,N_9210);
and U10461 (N_10461,N_9291,N_8524);
nor U10462 (N_10462,N_9452,N_8990);
xnor U10463 (N_10463,N_9381,N_9263);
xor U10464 (N_10464,N_9097,N_9315);
nor U10465 (N_10465,N_8765,N_9128);
nor U10466 (N_10466,N_9353,N_9390);
nor U10467 (N_10467,N_9279,N_9000);
and U10468 (N_10468,N_8655,N_8801);
nor U10469 (N_10469,N_8965,N_8700);
and U10470 (N_10470,N_9168,N_9289);
nand U10471 (N_10471,N_8436,N_8996);
xor U10472 (N_10472,N_8835,N_8871);
and U10473 (N_10473,N_9001,N_8827);
nand U10474 (N_10474,N_8945,N_9076);
nor U10475 (N_10475,N_9386,N_9528);
and U10476 (N_10476,N_9371,N_9011);
nand U10477 (N_10477,N_9463,N_9263);
nor U10478 (N_10478,N_9422,N_8992);
nor U10479 (N_10479,N_8494,N_9191);
or U10480 (N_10480,N_8802,N_8549);
and U10481 (N_10481,N_9156,N_9255);
nand U10482 (N_10482,N_8540,N_8741);
or U10483 (N_10483,N_8991,N_8833);
or U10484 (N_10484,N_9028,N_8433);
xor U10485 (N_10485,N_8754,N_9103);
or U10486 (N_10486,N_9375,N_9183);
nor U10487 (N_10487,N_8606,N_9116);
and U10488 (N_10488,N_8420,N_8482);
xor U10489 (N_10489,N_9528,N_8730);
xnor U10490 (N_10490,N_9320,N_9352);
nor U10491 (N_10491,N_9539,N_9282);
nand U10492 (N_10492,N_9088,N_9585);
xnor U10493 (N_10493,N_9226,N_8680);
and U10494 (N_10494,N_9368,N_8420);
xor U10495 (N_10495,N_8824,N_9004);
nand U10496 (N_10496,N_8984,N_9338);
or U10497 (N_10497,N_8958,N_8794);
nor U10498 (N_10498,N_8920,N_9184);
xnor U10499 (N_10499,N_9501,N_9379);
nand U10500 (N_10500,N_9288,N_9102);
nand U10501 (N_10501,N_8926,N_8737);
or U10502 (N_10502,N_9569,N_8734);
nor U10503 (N_10503,N_8945,N_8905);
and U10504 (N_10504,N_8416,N_9478);
nor U10505 (N_10505,N_9035,N_8487);
nand U10506 (N_10506,N_8946,N_9130);
nor U10507 (N_10507,N_8578,N_9408);
nand U10508 (N_10508,N_9193,N_8893);
nor U10509 (N_10509,N_9594,N_9476);
xor U10510 (N_10510,N_8836,N_9122);
and U10511 (N_10511,N_8573,N_8470);
and U10512 (N_10512,N_8503,N_8521);
and U10513 (N_10513,N_9584,N_9389);
or U10514 (N_10514,N_9041,N_8813);
or U10515 (N_10515,N_9145,N_8832);
nand U10516 (N_10516,N_8677,N_9224);
xor U10517 (N_10517,N_8627,N_8593);
xnor U10518 (N_10518,N_8540,N_8624);
and U10519 (N_10519,N_9008,N_8466);
nor U10520 (N_10520,N_8466,N_8899);
nand U10521 (N_10521,N_9150,N_9128);
or U10522 (N_10522,N_9232,N_8552);
nand U10523 (N_10523,N_9429,N_8600);
or U10524 (N_10524,N_9179,N_8924);
and U10525 (N_10525,N_8917,N_9535);
nor U10526 (N_10526,N_9123,N_8677);
or U10527 (N_10527,N_9023,N_8908);
xor U10528 (N_10528,N_9021,N_8953);
or U10529 (N_10529,N_8700,N_8841);
and U10530 (N_10530,N_8845,N_8906);
and U10531 (N_10531,N_8518,N_8573);
or U10532 (N_10532,N_9224,N_9594);
nand U10533 (N_10533,N_8832,N_9052);
nor U10534 (N_10534,N_9505,N_9310);
xor U10535 (N_10535,N_8820,N_9383);
and U10536 (N_10536,N_9320,N_8685);
nor U10537 (N_10537,N_8408,N_9303);
and U10538 (N_10538,N_9572,N_9168);
xor U10539 (N_10539,N_8641,N_9549);
nor U10540 (N_10540,N_9502,N_8934);
or U10541 (N_10541,N_9051,N_8916);
nor U10542 (N_10542,N_8498,N_9414);
nand U10543 (N_10543,N_9497,N_9089);
nor U10544 (N_10544,N_9146,N_9382);
nor U10545 (N_10545,N_9480,N_9499);
nor U10546 (N_10546,N_8765,N_8773);
xor U10547 (N_10547,N_9206,N_8850);
nand U10548 (N_10548,N_8782,N_8545);
and U10549 (N_10549,N_8427,N_9331);
or U10550 (N_10550,N_8683,N_9422);
and U10551 (N_10551,N_8889,N_9335);
nand U10552 (N_10552,N_9058,N_9104);
nor U10553 (N_10553,N_8852,N_9357);
nand U10554 (N_10554,N_8493,N_8794);
or U10555 (N_10555,N_9455,N_8551);
or U10556 (N_10556,N_8917,N_8418);
or U10557 (N_10557,N_8859,N_8611);
or U10558 (N_10558,N_9574,N_9061);
or U10559 (N_10559,N_9054,N_9443);
and U10560 (N_10560,N_9183,N_8478);
or U10561 (N_10561,N_8572,N_8784);
nor U10562 (N_10562,N_9414,N_9469);
nor U10563 (N_10563,N_9066,N_8863);
nor U10564 (N_10564,N_9070,N_9490);
and U10565 (N_10565,N_9266,N_8604);
nor U10566 (N_10566,N_9236,N_8703);
nor U10567 (N_10567,N_9551,N_9338);
nor U10568 (N_10568,N_8670,N_9441);
or U10569 (N_10569,N_8935,N_8620);
and U10570 (N_10570,N_9487,N_9264);
xnor U10571 (N_10571,N_9574,N_8856);
nor U10572 (N_10572,N_9543,N_9077);
or U10573 (N_10573,N_9126,N_8608);
nor U10574 (N_10574,N_9150,N_8663);
and U10575 (N_10575,N_8876,N_8442);
nand U10576 (N_10576,N_8633,N_8832);
nand U10577 (N_10577,N_8724,N_9450);
nand U10578 (N_10578,N_9435,N_8447);
xnor U10579 (N_10579,N_9302,N_8810);
or U10580 (N_10580,N_9056,N_8518);
or U10581 (N_10581,N_9149,N_9048);
xnor U10582 (N_10582,N_9387,N_8832);
xnor U10583 (N_10583,N_8914,N_9217);
nand U10584 (N_10584,N_9075,N_8403);
nand U10585 (N_10585,N_8832,N_9348);
nor U10586 (N_10586,N_9469,N_8531);
nand U10587 (N_10587,N_8448,N_9370);
nand U10588 (N_10588,N_8794,N_9426);
and U10589 (N_10589,N_9459,N_9487);
nor U10590 (N_10590,N_9175,N_8740);
or U10591 (N_10591,N_9529,N_9261);
nand U10592 (N_10592,N_8625,N_9229);
and U10593 (N_10593,N_9183,N_8410);
and U10594 (N_10594,N_9001,N_9411);
or U10595 (N_10595,N_9390,N_8787);
nand U10596 (N_10596,N_9293,N_8401);
nor U10597 (N_10597,N_9451,N_9198);
nand U10598 (N_10598,N_8682,N_8796);
and U10599 (N_10599,N_8887,N_8457);
xor U10600 (N_10600,N_9413,N_8911);
xnor U10601 (N_10601,N_9080,N_9474);
or U10602 (N_10602,N_8833,N_9495);
nand U10603 (N_10603,N_9219,N_8610);
and U10604 (N_10604,N_9138,N_8868);
xor U10605 (N_10605,N_9049,N_9118);
or U10606 (N_10606,N_8734,N_9289);
or U10607 (N_10607,N_8470,N_9251);
or U10608 (N_10608,N_9036,N_8829);
or U10609 (N_10609,N_9014,N_9157);
or U10610 (N_10610,N_8615,N_8739);
xor U10611 (N_10611,N_9434,N_9187);
xnor U10612 (N_10612,N_9325,N_9057);
xor U10613 (N_10613,N_9359,N_9165);
xor U10614 (N_10614,N_8598,N_9200);
xnor U10615 (N_10615,N_9109,N_9542);
nor U10616 (N_10616,N_9060,N_9479);
nor U10617 (N_10617,N_8653,N_9345);
or U10618 (N_10618,N_9344,N_9523);
and U10619 (N_10619,N_8623,N_8802);
and U10620 (N_10620,N_9369,N_9072);
and U10621 (N_10621,N_8559,N_9175);
nor U10622 (N_10622,N_8533,N_8702);
nor U10623 (N_10623,N_9297,N_9138);
nand U10624 (N_10624,N_8830,N_8753);
nand U10625 (N_10625,N_8897,N_9538);
xnor U10626 (N_10626,N_8636,N_8404);
nand U10627 (N_10627,N_8481,N_9348);
or U10628 (N_10628,N_8418,N_9035);
nand U10629 (N_10629,N_8558,N_9368);
and U10630 (N_10630,N_9212,N_9181);
nand U10631 (N_10631,N_9188,N_8966);
and U10632 (N_10632,N_9242,N_9392);
or U10633 (N_10633,N_9198,N_9185);
or U10634 (N_10634,N_8588,N_9013);
and U10635 (N_10635,N_8620,N_9384);
xnor U10636 (N_10636,N_9191,N_9169);
xnor U10637 (N_10637,N_9411,N_8809);
xor U10638 (N_10638,N_9393,N_8930);
nor U10639 (N_10639,N_9232,N_9059);
and U10640 (N_10640,N_8823,N_8606);
nor U10641 (N_10641,N_9105,N_9241);
nor U10642 (N_10642,N_9239,N_9180);
nor U10643 (N_10643,N_8416,N_9380);
nand U10644 (N_10644,N_9293,N_9504);
nor U10645 (N_10645,N_8503,N_8783);
nor U10646 (N_10646,N_8635,N_9190);
nand U10647 (N_10647,N_9584,N_9238);
nand U10648 (N_10648,N_8868,N_9397);
or U10649 (N_10649,N_9026,N_8727);
nand U10650 (N_10650,N_8598,N_9469);
or U10651 (N_10651,N_8969,N_8548);
and U10652 (N_10652,N_8795,N_9565);
nor U10653 (N_10653,N_8928,N_9333);
xnor U10654 (N_10654,N_8739,N_9406);
or U10655 (N_10655,N_9254,N_8478);
nand U10656 (N_10656,N_8795,N_9286);
nand U10657 (N_10657,N_9372,N_8719);
nor U10658 (N_10658,N_8940,N_8512);
xor U10659 (N_10659,N_8478,N_8699);
or U10660 (N_10660,N_8796,N_9213);
nand U10661 (N_10661,N_8990,N_8582);
xnor U10662 (N_10662,N_8895,N_9173);
or U10663 (N_10663,N_8488,N_9573);
and U10664 (N_10664,N_9047,N_8539);
xor U10665 (N_10665,N_9586,N_8839);
nor U10666 (N_10666,N_8931,N_9046);
nor U10667 (N_10667,N_8891,N_8762);
xnor U10668 (N_10668,N_9138,N_9372);
nor U10669 (N_10669,N_8697,N_9321);
nor U10670 (N_10670,N_9500,N_9304);
and U10671 (N_10671,N_8832,N_9135);
and U10672 (N_10672,N_8966,N_9415);
xnor U10673 (N_10673,N_8571,N_8480);
xor U10674 (N_10674,N_9366,N_9229);
and U10675 (N_10675,N_9346,N_9206);
or U10676 (N_10676,N_8803,N_9407);
and U10677 (N_10677,N_8999,N_9282);
and U10678 (N_10678,N_8411,N_8683);
or U10679 (N_10679,N_8744,N_8626);
xnor U10680 (N_10680,N_8682,N_8420);
xnor U10681 (N_10681,N_8831,N_9115);
and U10682 (N_10682,N_8871,N_8704);
and U10683 (N_10683,N_8868,N_9096);
or U10684 (N_10684,N_8766,N_9502);
or U10685 (N_10685,N_8449,N_9205);
and U10686 (N_10686,N_8684,N_9291);
and U10687 (N_10687,N_9218,N_9143);
nand U10688 (N_10688,N_8726,N_9120);
nand U10689 (N_10689,N_9255,N_8585);
nand U10690 (N_10690,N_8466,N_9365);
or U10691 (N_10691,N_8700,N_9068);
xnor U10692 (N_10692,N_8806,N_8633);
and U10693 (N_10693,N_8448,N_9226);
nand U10694 (N_10694,N_9508,N_8870);
nand U10695 (N_10695,N_8797,N_9183);
xor U10696 (N_10696,N_9412,N_8538);
nand U10697 (N_10697,N_9255,N_9035);
xor U10698 (N_10698,N_8553,N_9407);
nor U10699 (N_10699,N_8591,N_9331);
nand U10700 (N_10700,N_8770,N_9468);
or U10701 (N_10701,N_9336,N_9523);
nor U10702 (N_10702,N_8882,N_9022);
and U10703 (N_10703,N_8839,N_9354);
nand U10704 (N_10704,N_8707,N_8703);
or U10705 (N_10705,N_8453,N_9592);
and U10706 (N_10706,N_8991,N_8551);
nor U10707 (N_10707,N_9159,N_8459);
xor U10708 (N_10708,N_9180,N_9337);
or U10709 (N_10709,N_8618,N_8890);
nor U10710 (N_10710,N_8495,N_9375);
nand U10711 (N_10711,N_9073,N_8940);
and U10712 (N_10712,N_8723,N_9317);
nor U10713 (N_10713,N_9108,N_8511);
and U10714 (N_10714,N_8418,N_8996);
nor U10715 (N_10715,N_8819,N_9077);
nand U10716 (N_10716,N_8515,N_9426);
nand U10717 (N_10717,N_8634,N_8641);
or U10718 (N_10718,N_9018,N_9159);
or U10719 (N_10719,N_9061,N_8623);
or U10720 (N_10720,N_9356,N_9482);
nor U10721 (N_10721,N_9199,N_8491);
xnor U10722 (N_10722,N_8819,N_9509);
and U10723 (N_10723,N_9124,N_9487);
nor U10724 (N_10724,N_8615,N_9290);
nor U10725 (N_10725,N_8926,N_8795);
xor U10726 (N_10726,N_8548,N_8514);
xnor U10727 (N_10727,N_9212,N_9486);
nor U10728 (N_10728,N_9130,N_9486);
or U10729 (N_10729,N_9248,N_8455);
nand U10730 (N_10730,N_9198,N_8657);
or U10731 (N_10731,N_8547,N_9314);
or U10732 (N_10732,N_8470,N_9452);
and U10733 (N_10733,N_9037,N_9560);
and U10734 (N_10734,N_8904,N_8965);
xor U10735 (N_10735,N_9303,N_8686);
nand U10736 (N_10736,N_8570,N_8717);
nor U10737 (N_10737,N_9193,N_9233);
xnor U10738 (N_10738,N_8505,N_8687);
or U10739 (N_10739,N_9131,N_9587);
nor U10740 (N_10740,N_9370,N_9129);
xnor U10741 (N_10741,N_8875,N_9588);
nand U10742 (N_10742,N_8762,N_9077);
xor U10743 (N_10743,N_8822,N_8800);
and U10744 (N_10744,N_9087,N_9271);
nand U10745 (N_10745,N_8918,N_9029);
nand U10746 (N_10746,N_9331,N_8485);
nand U10747 (N_10747,N_8647,N_8819);
nand U10748 (N_10748,N_9519,N_9161);
and U10749 (N_10749,N_8906,N_8633);
and U10750 (N_10750,N_9130,N_9433);
xnor U10751 (N_10751,N_8677,N_8784);
or U10752 (N_10752,N_8479,N_8750);
and U10753 (N_10753,N_8424,N_8766);
xor U10754 (N_10754,N_8501,N_9105);
nand U10755 (N_10755,N_8624,N_8575);
and U10756 (N_10756,N_9286,N_8834);
xnor U10757 (N_10757,N_8474,N_8834);
or U10758 (N_10758,N_9487,N_9518);
xnor U10759 (N_10759,N_9284,N_8925);
or U10760 (N_10760,N_9466,N_9509);
and U10761 (N_10761,N_8466,N_8691);
and U10762 (N_10762,N_8794,N_9050);
and U10763 (N_10763,N_8952,N_9531);
and U10764 (N_10764,N_9291,N_8946);
and U10765 (N_10765,N_8508,N_8805);
nand U10766 (N_10766,N_8953,N_9228);
xor U10767 (N_10767,N_9557,N_8783);
nand U10768 (N_10768,N_9075,N_9225);
or U10769 (N_10769,N_8591,N_8625);
and U10770 (N_10770,N_9209,N_8823);
xor U10771 (N_10771,N_8859,N_8410);
xnor U10772 (N_10772,N_9316,N_9061);
nor U10773 (N_10773,N_8999,N_9563);
xnor U10774 (N_10774,N_9491,N_9206);
nor U10775 (N_10775,N_9004,N_8930);
nand U10776 (N_10776,N_8694,N_9083);
and U10777 (N_10777,N_8618,N_9296);
nor U10778 (N_10778,N_9594,N_8545);
nor U10779 (N_10779,N_9521,N_9429);
nor U10780 (N_10780,N_8651,N_8969);
nor U10781 (N_10781,N_8442,N_8883);
and U10782 (N_10782,N_8640,N_9299);
or U10783 (N_10783,N_9569,N_9572);
xnor U10784 (N_10784,N_8712,N_8633);
nor U10785 (N_10785,N_9392,N_9222);
or U10786 (N_10786,N_9132,N_8583);
or U10787 (N_10787,N_8679,N_8748);
and U10788 (N_10788,N_8646,N_8936);
or U10789 (N_10789,N_8602,N_8535);
and U10790 (N_10790,N_8831,N_8577);
nor U10791 (N_10791,N_9219,N_9122);
and U10792 (N_10792,N_8443,N_9396);
xor U10793 (N_10793,N_9598,N_8979);
xor U10794 (N_10794,N_9454,N_9083);
nand U10795 (N_10795,N_8525,N_8608);
or U10796 (N_10796,N_9398,N_8949);
nor U10797 (N_10797,N_8490,N_8651);
and U10798 (N_10798,N_8756,N_9310);
xnor U10799 (N_10799,N_9135,N_9208);
and U10800 (N_10800,N_9828,N_10005);
or U10801 (N_10801,N_9698,N_9771);
nand U10802 (N_10802,N_10471,N_10002);
and U10803 (N_10803,N_10590,N_9864);
xor U10804 (N_10804,N_10658,N_9774);
nand U10805 (N_10805,N_9815,N_10742);
nand U10806 (N_10806,N_9999,N_9764);
nand U10807 (N_10807,N_10546,N_9773);
or U10808 (N_10808,N_10366,N_10328);
or U10809 (N_10809,N_10577,N_10374);
nor U10810 (N_10810,N_10682,N_10461);
or U10811 (N_10811,N_10357,N_10406);
nor U10812 (N_10812,N_9693,N_9796);
nor U10813 (N_10813,N_9637,N_10215);
and U10814 (N_10814,N_9869,N_9681);
nand U10815 (N_10815,N_10660,N_10695);
and U10816 (N_10816,N_9664,N_10148);
or U10817 (N_10817,N_9959,N_10584);
and U10818 (N_10818,N_9762,N_10063);
nor U10819 (N_10819,N_10319,N_10330);
nor U10820 (N_10820,N_10015,N_10012);
nand U10821 (N_10821,N_10007,N_9997);
and U10822 (N_10822,N_10073,N_9895);
nor U10823 (N_10823,N_10227,N_10340);
nor U10824 (N_10824,N_9735,N_9642);
xnor U10825 (N_10825,N_9628,N_10723);
xnor U10826 (N_10826,N_10788,N_10503);
and U10827 (N_10827,N_10204,N_10626);
nor U10828 (N_10828,N_10468,N_9643);
or U10829 (N_10829,N_10728,N_9650);
nand U10830 (N_10830,N_10191,N_10244);
or U10831 (N_10831,N_10190,N_10708);
and U10832 (N_10832,N_9622,N_9662);
xor U10833 (N_10833,N_10659,N_10674);
nand U10834 (N_10834,N_10194,N_9884);
nand U10835 (N_10835,N_10782,N_10383);
nor U10836 (N_10836,N_10218,N_10131);
xor U10837 (N_10837,N_10716,N_9956);
xnor U10838 (N_10838,N_10569,N_10100);
xnor U10839 (N_10839,N_10416,N_10405);
and U10840 (N_10840,N_9675,N_10663);
and U10841 (N_10841,N_10135,N_9836);
nand U10842 (N_10842,N_10394,N_10538);
and U10843 (N_10843,N_10678,N_10795);
or U10844 (N_10844,N_9854,N_10500);
xnor U10845 (N_10845,N_9678,N_10562);
and U10846 (N_10846,N_10236,N_9974);
and U10847 (N_10847,N_9683,N_10447);
xor U10848 (N_10848,N_9964,N_10243);
and U10849 (N_10849,N_9738,N_10566);
and U10850 (N_10850,N_9900,N_10565);
nand U10851 (N_10851,N_10303,N_9891);
and U10852 (N_10852,N_10113,N_10532);
nand U10853 (N_10853,N_10142,N_10107);
or U10854 (N_10854,N_10152,N_9640);
nor U10855 (N_10855,N_10008,N_10269);
or U10856 (N_10856,N_10645,N_10765);
or U10857 (N_10857,N_10010,N_10624);
xor U10858 (N_10858,N_10267,N_9962);
and U10859 (N_10859,N_10230,N_9667);
nor U10860 (N_10860,N_10030,N_10282);
or U10861 (N_10861,N_10455,N_10757);
xnor U10862 (N_10862,N_10472,N_10280);
and U10863 (N_10863,N_9690,N_10259);
nor U10864 (N_10864,N_10398,N_9811);
and U10865 (N_10865,N_10619,N_10484);
or U10866 (N_10866,N_10085,N_9679);
or U10867 (N_10867,N_9813,N_10410);
xor U10868 (N_10868,N_10032,N_10104);
nand U10869 (N_10869,N_10119,N_9990);
xnor U10870 (N_10870,N_9792,N_10247);
or U10871 (N_10871,N_9928,N_10163);
and U10872 (N_10872,N_9732,N_10601);
xnor U10873 (N_10873,N_10598,N_9927);
nor U10874 (N_10874,N_10384,N_10180);
nor U10875 (N_10875,N_10222,N_10497);
and U10876 (N_10876,N_9718,N_10697);
xnor U10877 (N_10877,N_10046,N_10099);
and U10878 (N_10878,N_10603,N_9783);
and U10879 (N_10879,N_10196,N_9987);
and U10880 (N_10880,N_9801,N_10050);
nor U10881 (N_10881,N_9803,N_10480);
nor U10882 (N_10882,N_9908,N_10754);
nand U10883 (N_10883,N_10375,N_10710);
and U10884 (N_10884,N_10111,N_10289);
and U10885 (N_10885,N_10534,N_10078);
xor U10886 (N_10886,N_10593,N_10517);
nor U10887 (N_10887,N_10225,N_9670);
and U10888 (N_10888,N_10140,N_9686);
or U10889 (N_10889,N_10199,N_9863);
xnor U10890 (N_10890,N_9739,N_10278);
or U10891 (N_10891,N_10096,N_10595);
xor U10892 (N_10892,N_10787,N_10509);
or U10893 (N_10893,N_10181,N_10769);
and U10894 (N_10894,N_10064,N_10501);
or U10895 (N_10895,N_10414,N_9697);
nor U10896 (N_10896,N_10570,N_10198);
or U10897 (N_10897,N_10102,N_9761);
nor U10898 (N_10898,N_10161,N_10170);
and U10899 (N_10899,N_9791,N_10691);
or U10900 (N_10900,N_10537,N_10056);
or U10901 (N_10901,N_10698,N_10790);
nor U10902 (N_10902,N_9782,N_10356);
and U10903 (N_10903,N_9763,N_9871);
xor U10904 (N_10904,N_10287,N_10126);
xnor U10905 (N_10905,N_10429,N_10117);
and U10906 (N_10906,N_10744,N_10689);
or U10907 (N_10907,N_9798,N_10144);
nor U10908 (N_10908,N_9949,N_10530);
nor U10909 (N_10909,N_9754,N_10427);
nor U10910 (N_10910,N_10178,N_9714);
nand U10911 (N_10911,N_10389,N_10137);
nand U10912 (N_10912,N_10737,N_10632);
nor U10913 (N_10913,N_9883,N_9867);
xor U10914 (N_10914,N_9753,N_9818);
xnor U10915 (N_10915,N_9940,N_10256);
xnor U10916 (N_10916,N_9725,N_10388);
and U10917 (N_10917,N_9674,N_10642);
nor U10918 (N_10918,N_9760,N_10029);
or U10919 (N_10919,N_10585,N_10460);
xor U10920 (N_10920,N_9847,N_9979);
nor U10921 (N_10921,N_10575,N_10223);
xnor U10922 (N_10922,N_9971,N_10034);
nand U10923 (N_10923,N_9817,N_10224);
nand U10924 (N_10924,N_10512,N_9939);
xnor U10925 (N_10925,N_10295,N_10294);
nor U10926 (N_10926,N_10004,N_10221);
and U10927 (N_10927,N_9861,N_10554);
xor U10928 (N_10928,N_10798,N_10553);
nor U10929 (N_10929,N_9776,N_10229);
or U10930 (N_10930,N_10138,N_10035);
and U10931 (N_10931,N_9743,N_10362);
nand U10932 (N_10932,N_10636,N_10611);
nor U10933 (N_10933,N_10367,N_9638);
and U10934 (N_10934,N_10618,N_9882);
and U10935 (N_10935,N_10783,N_9772);
and U10936 (N_10936,N_10132,N_10077);
and U10937 (N_10937,N_10671,N_10515);
nand U10938 (N_10938,N_9937,N_10616);
xnor U10939 (N_10939,N_9768,N_10571);
nor U10940 (N_10940,N_10157,N_10764);
xor U10941 (N_10941,N_10239,N_10321);
xor U10942 (N_10942,N_10628,N_10466);
nand U10943 (N_10943,N_10653,N_9832);
or U10944 (N_10944,N_10597,N_10298);
xnor U10945 (N_10945,N_9926,N_10122);
xor U10946 (N_10946,N_10232,N_10361);
xnor U10947 (N_10947,N_10607,N_9834);
nor U10948 (N_10948,N_9759,N_10150);
nor U10949 (N_10949,N_10345,N_9898);
and U10950 (N_10950,N_10589,N_10045);
and U10951 (N_10951,N_10341,N_10290);
and U10952 (N_10952,N_10772,N_9621);
xor U10953 (N_10953,N_9777,N_10508);
nand U10954 (N_10954,N_10605,N_9845);
xnor U10955 (N_10955,N_9737,N_10778);
and U10956 (N_10956,N_10439,N_10770);
and U10957 (N_10957,N_9914,N_9934);
and U10958 (N_10958,N_10792,N_10037);
nor U10959 (N_10959,N_9618,N_10060);
xor U10960 (N_10960,N_10520,N_10338);
nand U10961 (N_10961,N_9989,N_9862);
nand U10962 (N_10962,N_10610,N_9750);
and U10963 (N_10963,N_10041,N_10525);
nor U10964 (N_10964,N_10552,N_10775);
nor U10965 (N_10965,N_10291,N_10097);
nand U10966 (N_10966,N_10756,N_9850);
xnor U10967 (N_10967,N_9660,N_10453);
nand U10968 (N_10968,N_10668,N_10066);
and U10969 (N_10969,N_10648,N_9881);
xor U10970 (N_10970,N_9986,N_10071);
nand U10971 (N_10971,N_10160,N_10103);
nand U10972 (N_10972,N_10039,N_9631);
xnor U10973 (N_10973,N_9837,N_10110);
or U10974 (N_10974,N_10370,N_9703);
and U10975 (N_10975,N_9961,N_9710);
or U10976 (N_10976,N_10317,N_9938);
xor U10977 (N_10977,N_10780,N_9692);
or U10978 (N_10978,N_9919,N_9705);
nor U10979 (N_10979,N_10408,N_10167);
or U10980 (N_10980,N_9902,N_9767);
nor U10981 (N_10981,N_10544,N_10721);
and U10982 (N_10982,N_9838,N_10752);
and U10983 (N_10983,N_10040,N_10784);
or U10984 (N_10984,N_10320,N_10136);
or U10985 (N_10985,N_10694,N_9634);
and U10986 (N_10986,N_9985,N_9611);
xor U10987 (N_10987,N_9833,N_10048);
or U10988 (N_10988,N_10342,N_10479);
nor U10989 (N_10989,N_9757,N_9878);
and U10990 (N_10990,N_10664,N_9655);
or U10991 (N_10991,N_10271,N_10089);
and U10992 (N_10992,N_10067,N_10513);
xor U10993 (N_10993,N_9696,N_10255);
or U10994 (N_10994,N_10188,N_10623);
nand U10995 (N_10995,N_10358,N_10437);
and U10996 (N_10996,N_10718,N_10604);
nand U10997 (N_10997,N_10379,N_10675);
nand U10998 (N_10998,N_9819,N_10210);
nand U10999 (N_10999,N_10680,N_9633);
xnor U11000 (N_11000,N_10699,N_10692);
and U11001 (N_11001,N_10318,N_9712);
and U11002 (N_11002,N_10000,N_9676);
or U11003 (N_11003,N_10360,N_10331);
nand U11004 (N_11004,N_10419,N_9746);
nand U11005 (N_11005,N_9946,N_10730);
xor U11006 (N_11006,N_10541,N_10420);
and U11007 (N_11007,N_10677,N_10094);
nor U11008 (N_11008,N_10310,N_10777);
xor U11009 (N_11009,N_10643,N_10305);
nor U11010 (N_11010,N_10124,N_10667);
and U11011 (N_11011,N_10202,N_10095);
nor U11012 (N_11012,N_10545,N_10396);
and U11013 (N_11013,N_9765,N_10573);
nand U11014 (N_11014,N_9730,N_9831);
or U11015 (N_11015,N_10302,N_10175);
nor U11016 (N_11016,N_10679,N_9930);
xnor U11017 (N_11017,N_10174,N_9616);
nor U11018 (N_11018,N_9614,N_10558);
and U11019 (N_11019,N_9810,N_10033);
nor U11020 (N_11020,N_10147,N_9694);
xor U11021 (N_11021,N_10141,N_10038);
nor U11022 (N_11022,N_10314,N_9879);
nand U11023 (N_11023,N_9972,N_10169);
xor U11024 (N_11024,N_9913,N_9733);
nor U11025 (N_11025,N_10108,N_10514);
xor U11026 (N_11026,N_10324,N_10596);
xor U11027 (N_11027,N_9748,N_10153);
or U11028 (N_11028,N_10542,N_10703);
xnor U11029 (N_11029,N_9952,N_10380);
or U11030 (N_11030,N_10608,N_9708);
nand U11031 (N_11031,N_9687,N_9639);
nand U11032 (N_11032,N_10003,N_9797);
nand U11033 (N_11033,N_9843,N_10307);
nor U11034 (N_11034,N_10347,N_10673);
nand U11035 (N_11035,N_9865,N_10081);
xnor U11036 (N_11036,N_9886,N_10452);
nor U11037 (N_11037,N_10751,N_10650);
and U11038 (N_11038,N_9799,N_9994);
xnor U11039 (N_11039,N_10759,N_10794);
or U11040 (N_11040,N_10106,N_10092);
nor U11041 (N_11041,N_9852,N_9713);
or U11042 (N_11042,N_10485,N_9669);
nor U11043 (N_11043,N_10011,N_10434);
or U11044 (N_11044,N_10502,N_10241);
and U11045 (N_11045,N_10683,N_9947);
and U11046 (N_11046,N_9800,N_10425);
and U11047 (N_11047,N_9704,N_10154);
and U11048 (N_11048,N_10422,N_10519);
or U11049 (N_11049,N_10771,N_9756);
and U11050 (N_11050,N_10171,N_10395);
or U11051 (N_11051,N_9641,N_10696);
nor U11052 (N_11052,N_10183,N_9781);
nor U11053 (N_11053,N_10237,N_9630);
nand U11054 (N_11054,N_10109,N_10490);
or U11055 (N_11055,N_10327,N_10062);
nand U11056 (N_11056,N_10495,N_10409);
xnor U11057 (N_11057,N_10768,N_9721);
and U11058 (N_11058,N_10676,N_10024);
nor U11059 (N_11059,N_10638,N_10785);
xor U11060 (N_11060,N_10368,N_9917);
and U11061 (N_11061,N_10612,N_10155);
xor U11062 (N_11062,N_10214,N_10172);
nor U11063 (N_11063,N_10690,N_10505);
and U11064 (N_11064,N_10450,N_9996);
nor U11065 (N_11065,N_10745,N_10657);
xor U11066 (N_11066,N_10749,N_10572);
nor U11067 (N_11067,N_10776,N_10615);
nor U11068 (N_11068,N_10344,N_10209);
xnor U11069 (N_11069,N_9691,N_9876);
or U11070 (N_11070,N_10234,N_9602);
xnor U11071 (N_11071,N_9720,N_10293);
nor U11072 (N_11072,N_10235,N_10350);
xnor U11073 (N_11073,N_10426,N_9846);
xor U11074 (N_11074,N_10463,N_10684);
nand U11075 (N_11075,N_9751,N_10755);
or U11076 (N_11076,N_10335,N_9632);
xnor U11077 (N_11077,N_10753,N_10264);
nor U11078 (N_11078,N_9849,N_9855);
nand U11079 (N_11079,N_10630,N_9809);
nand U11080 (N_11080,N_10220,N_10299);
nor U11081 (N_11081,N_10579,N_9734);
and U11082 (N_11082,N_10702,N_9982);
and U11083 (N_11083,N_9646,N_10424);
or U11084 (N_11084,N_9950,N_10149);
xnor U11085 (N_11085,N_10740,N_10313);
xnor U11086 (N_11086,N_10528,N_10477);
nor U11087 (N_11087,N_10219,N_10296);
and U11088 (N_11088,N_10134,N_9857);
xor U11089 (N_11089,N_10655,N_10581);
and U11090 (N_11090,N_9840,N_10326);
or U11091 (N_11091,N_9620,N_9976);
nand U11092 (N_11092,N_10348,N_10057);
nand U11093 (N_11093,N_10251,N_10182);
or U11094 (N_11094,N_10486,N_10334);
nand U11095 (N_11095,N_10205,N_10779);
nand U11096 (N_11096,N_10462,N_10731);
xnor U11097 (N_11097,N_10189,N_10760);
nor U11098 (N_11098,N_9995,N_10014);
or U11099 (N_11099,N_10233,N_10028);
xor U11100 (N_11100,N_10079,N_9823);
nand U11101 (N_11101,N_10726,N_10415);
nand U11102 (N_11102,N_10401,N_9603);
nor U11103 (N_11103,N_9715,N_10614);
or U11104 (N_11104,N_10750,N_9775);
nor U11105 (N_11105,N_9766,N_9711);
nand U11106 (N_11106,N_10563,N_10662);
xor U11107 (N_11107,N_10261,N_10083);
nand U11108 (N_11108,N_10719,N_10449);
or U11109 (N_11109,N_9923,N_10253);
and U11110 (N_11110,N_9780,N_10279);
nor U11111 (N_11111,N_10043,N_9741);
nand U11112 (N_11112,N_10504,N_10164);
nand U11113 (N_11113,N_10550,N_9835);
xnor U11114 (N_11114,N_9787,N_9851);
and U11115 (N_11115,N_10114,N_10635);
nor U11116 (N_11116,N_9747,N_10070);
or U11117 (N_11117,N_10743,N_10533);
xnor U11118 (N_11118,N_10793,N_9924);
nand U11119 (N_11119,N_10337,N_10454);
nand U11120 (N_11120,N_10187,N_9680);
and U11121 (N_11121,N_10378,N_10052);
nor U11122 (N_11122,N_10574,N_10524);
nor U11123 (N_11123,N_9910,N_10438);
or U11124 (N_11124,N_9903,N_10156);
nand U11125 (N_11125,N_9856,N_10591);
xor U11126 (N_11126,N_9794,N_10588);
nor U11127 (N_11127,N_10580,N_9647);
and U11128 (N_11128,N_9727,N_10311);
nand U11129 (N_11129,N_9933,N_9617);
xnor U11130 (N_11130,N_10207,N_10712);
and U11131 (N_11131,N_10376,N_10457);
nor U11132 (N_11132,N_10464,N_10786);
or U11133 (N_11133,N_10470,N_10625);
or U11134 (N_11134,N_9812,N_10561);
nor U11135 (N_11135,N_10799,N_10088);
xnor U11136 (N_11136,N_10309,N_10392);
nor U11137 (N_11137,N_9899,N_10065);
nor U11138 (N_11138,N_10536,N_9954);
and U11139 (N_11139,N_10036,N_10701);
nor U11140 (N_11140,N_10443,N_9790);
nor U11141 (N_11141,N_9609,N_10143);
or U11142 (N_11142,N_9804,N_9607);
nand U11143 (N_11143,N_10606,N_9625);
and U11144 (N_11144,N_10781,N_9844);
nor U11145 (N_11145,N_9916,N_9935);
or U11146 (N_11146,N_10640,N_10411);
nand U11147 (N_11147,N_10578,N_9969);
nor U11148 (N_11148,N_9918,N_9793);
nand U11149 (N_11149,N_10487,N_10185);
and U11150 (N_11150,N_10158,N_10260);
xnor U11151 (N_11151,N_9877,N_10206);
xnor U11152 (N_11152,N_10281,N_9841);
or U11153 (N_11153,N_10019,N_10724);
nor U11154 (N_11154,N_10707,N_10200);
nand U11155 (N_11155,N_9728,N_10483);
xnor U11156 (N_11156,N_10300,N_9752);
nor U11157 (N_11157,N_10074,N_10404);
nor U11158 (N_11158,N_9889,N_10539);
nor U11159 (N_11159,N_10061,N_10633);
or U11160 (N_11160,N_10722,N_10531);
xnor U11161 (N_11161,N_9859,N_10284);
nand U11162 (N_11162,N_9839,N_9953);
nor U11163 (N_11163,N_10093,N_9717);
and U11164 (N_11164,N_9610,N_10120);
xnor U11165 (N_11165,N_10700,N_10308);
and U11166 (N_11166,N_10343,N_10322);
xor U11167 (N_11167,N_10613,N_9984);
xnor U11168 (N_11168,N_10417,N_9932);
or U11169 (N_11169,N_9821,N_9661);
or U11170 (N_11170,N_10166,N_10423);
and U11171 (N_11171,N_9740,N_10262);
or U11172 (N_11172,N_10709,N_10400);
nand U11173 (N_11173,N_9673,N_10016);
xor U11174 (N_11174,N_10118,N_9853);
and U11175 (N_11175,N_10725,N_10516);
and U11176 (N_11176,N_9880,N_10339);
nand U11177 (N_11177,N_9677,N_10403);
nor U11178 (N_11178,N_9684,N_10129);
xnor U11179 (N_11179,N_10448,N_10518);
and U11180 (N_11180,N_10796,N_10714);
xnor U11181 (N_11181,N_9649,N_9967);
nand U11182 (N_11182,N_9612,N_10734);
nor U11183 (N_11183,N_10482,N_10639);
nand U11184 (N_11184,N_10025,N_10767);
nor U11185 (N_11185,N_10249,N_10669);
or U11186 (N_11186,N_10521,N_10201);
or U11187 (N_11187,N_10494,N_10706);
nor U11188 (N_11188,N_10741,N_10681);
or U11189 (N_11189,N_10257,N_10576);
xnor U11190 (N_11190,N_10058,N_10001);
or U11191 (N_11191,N_9770,N_10369);
and U11192 (N_11192,N_10746,N_10715);
or U11193 (N_11193,N_9860,N_10240);
xor U11194 (N_11194,N_9826,N_10727);
nand U11195 (N_11195,N_10192,N_10090);
xnor U11196 (N_11196,N_10456,N_10548);
nand U11197 (N_11197,N_10285,N_9873);
and U11198 (N_11198,N_10254,N_10351);
nor U11199 (N_11199,N_10634,N_9755);
and U11200 (N_11200,N_10499,N_10023);
or U11201 (N_11201,N_10665,N_10125);
or U11202 (N_11202,N_10274,N_10474);
or U11203 (N_11203,N_9742,N_10560);
xnor U11204 (N_11204,N_9601,N_10087);
nor U11205 (N_11205,N_9719,N_10130);
nor U11206 (N_11206,N_10250,N_10549);
nand U11207 (N_11207,N_10353,N_9744);
xor U11208 (N_11208,N_9868,N_10146);
nor U11209 (N_11209,N_9626,N_10373);
and U11210 (N_11210,N_10355,N_9991);
xnor U11211 (N_11211,N_10162,N_9897);
or U11212 (N_11212,N_10622,N_10761);
or U11213 (N_11213,N_9769,N_10594);
or U11214 (N_11214,N_10364,N_9929);
nand U11215 (N_11215,N_10333,N_9842);
or U11216 (N_11216,N_9890,N_10082);
and U11217 (N_11217,N_10688,N_10276);
or U11218 (N_11218,N_10323,N_10748);
and U11219 (N_11219,N_9920,N_10245);
or U11220 (N_11220,N_9870,N_10432);
nor U11221 (N_11221,N_10197,N_10105);
or U11222 (N_11222,N_10489,N_10349);
nand U11223 (N_11223,N_10583,N_10458);
nor U11224 (N_11224,N_9945,N_10133);
or U11225 (N_11225,N_10672,N_10602);
nor U11226 (N_11226,N_10265,N_9825);
xnor U11227 (N_11227,N_9805,N_9659);
xor U11228 (N_11228,N_10145,N_9906);
or U11229 (N_11229,N_10195,N_9701);
xnor U11230 (N_11230,N_10592,N_9668);
xnor U11231 (N_11231,N_10151,N_10713);
or U11232 (N_11232,N_10582,N_10733);
nand U11233 (N_11233,N_10231,N_9973);
nor U11234 (N_11234,N_10084,N_10435);
or U11235 (N_11235,N_10354,N_9955);
and U11236 (N_11236,N_9722,N_9830);
xnor U11237 (N_11237,N_10022,N_10051);
and U11238 (N_11238,N_10018,N_10661);
or U11239 (N_11239,N_10292,N_10412);
and U11240 (N_11240,N_9784,N_10629);
xnor U11241 (N_11241,N_10059,N_9915);
xnor U11242 (N_11242,N_9905,N_10522);
or U11243 (N_11243,N_10551,N_10047);
xnor U11244 (N_11244,N_10399,N_10773);
xor U11245 (N_11245,N_10381,N_10316);
or U11246 (N_11246,N_10476,N_10248);
xor U11247 (N_11247,N_10031,N_10556);
or U11248 (N_11248,N_10213,N_10127);
nand U11249 (N_11249,N_10228,N_10736);
xor U11250 (N_11250,N_10054,N_10526);
and U11251 (N_11251,N_10547,N_9957);
nand U11252 (N_11252,N_10270,N_9789);
nand U11253 (N_11253,N_9613,N_9778);
nand U11254 (N_11254,N_10382,N_9688);
nor U11255 (N_11255,N_10325,N_10115);
xor U11256 (N_11256,N_10735,N_10493);
xor U11257 (N_11257,N_10179,N_10072);
nand U11258 (N_11258,N_9981,N_10555);
and U11259 (N_11259,N_10272,N_10217);
nand U11260 (N_11260,N_10444,N_10397);
or U11261 (N_11261,N_10193,N_10128);
xor U11262 (N_11262,N_10445,N_10617);
nor U11263 (N_11263,N_10586,N_9758);
xnor U11264 (N_11264,N_9716,N_9975);
or U11265 (N_11265,N_10069,N_9808);
nand U11266 (N_11266,N_9875,N_10506);
nor U11267 (N_11267,N_10766,N_9922);
and U11268 (N_11268,N_9912,N_9963);
nor U11269 (N_11269,N_10268,N_9998);
xor U11270 (N_11270,N_10621,N_10242);
nand U11271 (N_11271,N_10371,N_9885);
nor U11272 (N_11272,N_9911,N_10101);
xor U11273 (N_11273,N_10017,N_10705);
nand U11274 (N_11274,N_9665,N_10091);
nor U11275 (N_11275,N_10184,N_10332);
nor U11276 (N_11276,N_9731,N_9700);
nand U11277 (N_11277,N_9779,N_9635);
nor U11278 (N_11278,N_10386,N_10246);
nor U11279 (N_11279,N_10631,N_9689);
nor U11280 (N_11280,N_9606,N_10440);
or U11281 (N_11281,N_9695,N_10263);
or U11282 (N_11282,N_10402,N_9785);
and U11283 (N_11283,N_10644,N_9887);
and U11284 (N_11284,N_10704,N_10465);
nand U11285 (N_11285,N_9663,N_10226);
nor U11286 (N_11286,N_9824,N_9644);
and U11287 (N_11287,N_10666,N_9723);
nand U11288 (N_11288,N_10080,N_10637);
nor U11289 (N_11289,N_9645,N_10027);
and U11290 (N_11290,N_10738,N_10732);
and U11291 (N_11291,N_10407,N_10567);
xor U11292 (N_11292,N_10646,N_10442);
xnor U11293 (N_11293,N_9827,N_9672);
xnor U11294 (N_11294,N_10055,N_10729);
nor U11295 (N_11295,N_10053,N_9909);
and U11296 (N_11296,N_10433,N_10687);
xnor U11297 (N_11297,N_9992,N_10441);
and U11298 (N_11298,N_10009,N_10491);
xnor U11299 (N_11299,N_10098,N_10436);
nand U11300 (N_11300,N_9894,N_9699);
xnor U11301 (N_11301,N_9671,N_10315);
xor U11302 (N_11302,N_10359,N_10609);
xnor U11303 (N_11303,N_10301,N_10564);
nand U11304 (N_11304,N_9858,N_10762);
and U11305 (N_11305,N_10075,N_10176);
nor U11306 (N_11306,N_9685,N_9872);
nand U11307 (N_11307,N_9627,N_9951);
or U11308 (N_11308,N_9749,N_10720);
and U11309 (N_11309,N_9709,N_10159);
or U11310 (N_11310,N_9608,N_9653);
nand U11311 (N_11311,N_10076,N_9619);
nand U11312 (N_11312,N_10620,N_9978);
nor U11313 (N_11313,N_10116,N_10372);
nor U11314 (N_11314,N_9965,N_10747);
nor U11315 (N_11315,N_9706,N_10418);
nand U11316 (N_11316,N_9624,N_9904);
or U11317 (N_11317,N_10275,N_10599);
nand U11318 (N_11318,N_10459,N_10654);
nor U11319 (N_11319,N_10121,N_10177);
and U11320 (N_11320,N_10496,N_10510);
xor U11321 (N_11321,N_9893,N_10006);
xor U11322 (N_11322,N_9666,N_10670);
xor U11323 (N_11323,N_9814,N_10488);
and U11324 (N_11324,N_10469,N_9829);
xor U11325 (N_11325,N_10211,N_10173);
and U11326 (N_11326,N_9977,N_9848);
and U11327 (N_11327,N_10641,N_10789);
and U11328 (N_11328,N_9966,N_9600);
nor U11329 (N_11329,N_9941,N_10428);
xnor U11330 (N_11330,N_9656,N_10329);
and U11331 (N_11331,N_10523,N_9958);
or U11332 (N_11332,N_9948,N_9943);
or U11333 (N_11333,N_9896,N_9795);
xnor U11334 (N_11334,N_10686,N_10086);
xnor U11335 (N_11335,N_10273,N_10559);
or U11336 (N_11336,N_10208,N_10252);
or U11337 (N_11337,N_9892,N_9866);
nand U11338 (N_11338,N_10478,N_10306);
nand U11339 (N_11339,N_10390,N_10112);
xor U11340 (N_11340,N_10431,N_10774);
nand U11341 (N_11341,N_10346,N_9605);
and U11342 (N_11342,N_9925,N_9980);
or U11343 (N_11343,N_10791,N_9724);
nor U11344 (N_11344,N_9907,N_10283);
nor U11345 (N_11345,N_10527,N_10498);
nand U11346 (N_11346,N_9745,N_10363);
or U11347 (N_11347,N_10068,N_10451);
and U11348 (N_11348,N_10413,N_10186);
xor U11349 (N_11349,N_10352,N_10168);
and U11350 (N_11350,N_10763,N_10385);
or U11351 (N_11351,N_9942,N_9652);
nand U11352 (N_11352,N_10026,N_10277);
and U11353 (N_11353,N_10568,N_10758);
or U11354 (N_11354,N_10651,N_9983);
nand U11355 (N_11355,N_10266,N_10507);
and U11356 (N_11356,N_10717,N_9788);
or U11357 (N_11357,N_10020,N_9726);
nand U11358 (N_11358,N_9636,N_10649);
xor U11359 (N_11359,N_10492,N_10377);
nor U11360 (N_11360,N_10238,N_10475);
xor U11361 (N_11361,N_10013,N_10557);
or U11362 (N_11362,N_9654,N_10365);
xor U11363 (N_11363,N_9615,N_10627);
nor U11364 (N_11364,N_9707,N_9806);
and U11365 (N_11365,N_10421,N_10165);
nand U11366 (N_11366,N_9786,N_10511);
nor U11367 (N_11367,N_9729,N_10391);
nand U11368 (N_11368,N_10312,N_10387);
or U11369 (N_11369,N_10693,N_10656);
or U11370 (N_11370,N_10473,N_10467);
nand U11371 (N_11371,N_10647,N_10203);
nor U11372 (N_11372,N_10739,N_10258);
nand U11373 (N_11373,N_10286,N_9648);
nand U11374 (N_11374,N_10430,N_10797);
nand U11375 (N_11375,N_10600,N_10685);
xnor U11376 (N_11376,N_10042,N_9651);
xnor U11377 (N_11377,N_9623,N_9629);
and U11378 (N_11378,N_9657,N_9736);
and U11379 (N_11379,N_10044,N_9921);
and U11380 (N_11380,N_10540,N_9901);
and U11381 (N_11381,N_10529,N_9970);
xor U11382 (N_11382,N_9822,N_9820);
nand U11383 (N_11383,N_9682,N_10049);
or U11384 (N_11384,N_9988,N_10021);
xnor U11385 (N_11385,N_9931,N_10481);
and U11386 (N_11386,N_10216,N_9936);
xnor U11387 (N_11387,N_9944,N_9874);
nor U11388 (N_11388,N_10587,N_9658);
nor U11389 (N_11389,N_10297,N_10139);
nor U11390 (N_11390,N_9968,N_10535);
and U11391 (N_11391,N_9604,N_9802);
or U11392 (N_11392,N_9888,N_10212);
and U11393 (N_11393,N_10336,N_10393);
or U11394 (N_11394,N_10711,N_9993);
nand U11395 (N_11395,N_10288,N_9816);
nor U11396 (N_11396,N_9960,N_10543);
or U11397 (N_11397,N_9807,N_10304);
nand U11398 (N_11398,N_10446,N_9702);
nand U11399 (N_11399,N_10652,N_10123);
or U11400 (N_11400,N_10192,N_9981);
xnor U11401 (N_11401,N_10097,N_9737);
and U11402 (N_11402,N_9660,N_9864);
nor U11403 (N_11403,N_10001,N_10587);
or U11404 (N_11404,N_10561,N_10157);
nor U11405 (N_11405,N_10271,N_10189);
nor U11406 (N_11406,N_10249,N_10752);
nand U11407 (N_11407,N_10247,N_10352);
or U11408 (N_11408,N_10208,N_10561);
xor U11409 (N_11409,N_10042,N_9665);
xnor U11410 (N_11410,N_10523,N_9858);
and U11411 (N_11411,N_10065,N_10317);
nand U11412 (N_11412,N_10377,N_10628);
nand U11413 (N_11413,N_9955,N_10018);
nor U11414 (N_11414,N_9882,N_9734);
xnor U11415 (N_11415,N_10386,N_9729);
or U11416 (N_11416,N_10297,N_9647);
xnor U11417 (N_11417,N_10084,N_10795);
nand U11418 (N_11418,N_9721,N_10222);
xor U11419 (N_11419,N_10714,N_10219);
xor U11420 (N_11420,N_10540,N_10793);
or U11421 (N_11421,N_10266,N_10128);
nand U11422 (N_11422,N_10482,N_9989);
and U11423 (N_11423,N_10107,N_10342);
and U11424 (N_11424,N_10078,N_10122);
or U11425 (N_11425,N_10403,N_10737);
or U11426 (N_11426,N_10110,N_9710);
nor U11427 (N_11427,N_9653,N_10359);
and U11428 (N_11428,N_10441,N_9931);
xnor U11429 (N_11429,N_10691,N_10130);
nor U11430 (N_11430,N_10291,N_9636);
nor U11431 (N_11431,N_10256,N_10686);
nand U11432 (N_11432,N_10319,N_9977);
and U11433 (N_11433,N_9970,N_9749);
nand U11434 (N_11434,N_9786,N_9601);
nand U11435 (N_11435,N_10284,N_10635);
nand U11436 (N_11436,N_9945,N_9746);
nor U11437 (N_11437,N_10130,N_10053);
nand U11438 (N_11438,N_9869,N_10613);
nand U11439 (N_11439,N_10064,N_10022);
nor U11440 (N_11440,N_10068,N_10006);
and U11441 (N_11441,N_9970,N_9834);
or U11442 (N_11442,N_10308,N_10657);
nor U11443 (N_11443,N_10356,N_9751);
nor U11444 (N_11444,N_10469,N_10763);
or U11445 (N_11445,N_9869,N_10514);
nand U11446 (N_11446,N_10231,N_9851);
or U11447 (N_11447,N_9899,N_9765);
or U11448 (N_11448,N_10423,N_9780);
or U11449 (N_11449,N_9803,N_10551);
xnor U11450 (N_11450,N_9868,N_10057);
nor U11451 (N_11451,N_10352,N_10681);
or U11452 (N_11452,N_9865,N_10077);
nand U11453 (N_11453,N_10465,N_10059);
nor U11454 (N_11454,N_10063,N_10765);
xor U11455 (N_11455,N_10346,N_9710);
nor U11456 (N_11456,N_10435,N_9635);
and U11457 (N_11457,N_10534,N_10662);
nor U11458 (N_11458,N_9930,N_9840);
xnor U11459 (N_11459,N_10695,N_10475);
nand U11460 (N_11460,N_9641,N_10416);
xnor U11461 (N_11461,N_9868,N_9802);
nand U11462 (N_11462,N_10464,N_10241);
xor U11463 (N_11463,N_10668,N_9995);
xor U11464 (N_11464,N_10144,N_10471);
nor U11465 (N_11465,N_9757,N_10771);
nor U11466 (N_11466,N_9725,N_10436);
nand U11467 (N_11467,N_9832,N_10045);
or U11468 (N_11468,N_10659,N_9796);
xnor U11469 (N_11469,N_10740,N_10751);
and U11470 (N_11470,N_10107,N_10736);
nor U11471 (N_11471,N_10131,N_9749);
xnor U11472 (N_11472,N_10323,N_9925);
nor U11473 (N_11473,N_9908,N_10552);
nor U11474 (N_11474,N_9863,N_9660);
and U11475 (N_11475,N_10534,N_10471);
and U11476 (N_11476,N_9889,N_9878);
nand U11477 (N_11477,N_9788,N_9649);
xnor U11478 (N_11478,N_10282,N_10622);
xor U11479 (N_11479,N_10427,N_10508);
xor U11480 (N_11480,N_10744,N_10424);
xnor U11481 (N_11481,N_10164,N_9649);
xnor U11482 (N_11482,N_10234,N_10668);
xnor U11483 (N_11483,N_10230,N_9856);
xor U11484 (N_11484,N_10215,N_10111);
nor U11485 (N_11485,N_10051,N_10172);
xor U11486 (N_11486,N_9864,N_9665);
nor U11487 (N_11487,N_10239,N_10219);
nor U11488 (N_11488,N_10255,N_10557);
nand U11489 (N_11489,N_9862,N_10253);
nand U11490 (N_11490,N_9820,N_9957);
nor U11491 (N_11491,N_10582,N_10707);
nor U11492 (N_11492,N_9992,N_10056);
xnor U11493 (N_11493,N_10221,N_9743);
or U11494 (N_11494,N_10706,N_10611);
xor U11495 (N_11495,N_9897,N_10697);
xor U11496 (N_11496,N_10118,N_10737);
or U11497 (N_11497,N_10378,N_10167);
and U11498 (N_11498,N_10755,N_10327);
xor U11499 (N_11499,N_10711,N_9844);
and U11500 (N_11500,N_10271,N_9601);
and U11501 (N_11501,N_10632,N_10072);
nand U11502 (N_11502,N_9850,N_10244);
and U11503 (N_11503,N_10294,N_9670);
xnor U11504 (N_11504,N_10023,N_10508);
and U11505 (N_11505,N_10764,N_10096);
nand U11506 (N_11506,N_10243,N_10305);
xor U11507 (N_11507,N_10487,N_10601);
nor U11508 (N_11508,N_10498,N_10699);
xor U11509 (N_11509,N_10305,N_9777);
and U11510 (N_11510,N_9888,N_10197);
or U11511 (N_11511,N_9856,N_10179);
or U11512 (N_11512,N_9725,N_10761);
nor U11513 (N_11513,N_10243,N_9858);
nand U11514 (N_11514,N_10525,N_9900);
or U11515 (N_11515,N_9824,N_10299);
xnor U11516 (N_11516,N_9673,N_10048);
nand U11517 (N_11517,N_10358,N_9669);
or U11518 (N_11518,N_10169,N_9715);
nor U11519 (N_11519,N_10004,N_10306);
and U11520 (N_11520,N_10648,N_9919);
xnor U11521 (N_11521,N_10774,N_9972);
nor U11522 (N_11522,N_10018,N_10657);
or U11523 (N_11523,N_10248,N_10186);
and U11524 (N_11524,N_10319,N_9992);
nor U11525 (N_11525,N_10112,N_10391);
xor U11526 (N_11526,N_9788,N_9889);
and U11527 (N_11527,N_10183,N_10085);
nand U11528 (N_11528,N_10070,N_10455);
or U11529 (N_11529,N_10286,N_9853);
xor U11530 (N_11530,N_10722,N_9854);
nand U11531 (N_11531,N_10628,N_10069);
xnor U11532 (N_11532,N_10312,N_10779);
nor U11533 (N_11533,N_10690,N_10173);
or U11534 (N_11534,N_10483,N_10361);
and U11535 (N_11535,N_10389,N_10639);
nand U11536 (N_11536,N_9919,N_9765);
or U11537 (N_11537,N_10101,N_10704);
and U11538 (N_11538,N_10408,N_10552);
nor U11539 (N_11539,N_10529,N_10302);
xor U11540 (N_11540,N_10425,N_9885);
and U11541 (N_11541,N_10243,N_10388);
nand U11542 (N_11542,N_9856,N_9916);
nor U11543 (N_11543,N_10766,N_10181);
xnor U11544 (N_11544,N_10525,N_10306);
and U11545 (N_11545,N_10135,N_9683);
nand U11546 (N_11546,N_10561,N_10588);
nor U11547 (N_11547,N_9643,N_10733);
xor U11548 (N_11548,N_9856,N_9748);
nand U11549 (N_11549,N_10202,N_10772);
xor U11550 (N_11550,N_10551,N_9709);
xnor U11551 (N_11551,N_9878,N_10686);
or U11552 (N_11552,N_10293,N_9763);
nor U11553 (N_11553,N_10423,N_10231);
xor U11554 (N_11554,N_9916,N_10313);
nor U11555 (N_11555,N_10217,N_9929);
or U11556 (N_11556,N_10444,N_9624);
xor U11557 (N_11557,N_10463,N_10608);
xor U11558 (N_11558,N_10014,N_10286);
nor U11559 (N_11559,N_10120,N_10145);
nand U11560 (N_11560,N_10078,N_10096);
nor U11561 (N_11561,N_9899,N_10564);
nor U11562 (N_11562,N_9931,N_10350);
or U11563 (N_11563,N_9614,N_10088);
and U11564 (N_11564,N_10278,N_10478);
xor U11565 (N_11565,N_9827,N_10416);
xor U11566 (N_11566,N_10013,N_10608);
nor U11567 (N_11567,N_10251,N_10188);
nand U11568 (N_11568,N_9751,N_10062);
or U11569 (N_11569,N_9741,N_9877);
or U11570 (N_11570,N_10072,N_10513);
and U11571 (N_11571,N_10726,N_10364);
and U11572 (N_11572,N_10648,N_10547);
and U11573 (N_11573,N_9806,N_10550);
nor U11574 (N_11574,N_9899,N_10449);
nor U11575 (N_11575,N_10476,N_10046);
xor U11576 (N_11576,N_10445,N_10654);
xor U11577 (N_11577,N_9824,N_9624);
xnor U11578 (N_11578,N_10141,N_9797);
nor U11579 (N_11579,N_10094,N_9880);
and U11580 (N_11580,N_10739,N_10081);
or U11581 (N_11581,N_9684,N_10140);
or U11582 (N_11582,N_9842,N_10761);
or U11583 (N_11583,N_10177,N_10433);
or U11584 (N_11584,N_9900,N_10475);
and U11585 (N_11585,N_10196,N_10625);
and U11586 (N_11586,N_10404,N_9622);
xnor U11587 (N_11587,N_10669,N_9671);
and U11588 (N_11588,N_10647,N_9695);
or U11589 (N_11589,N_10306,N_10684);
xor U11590 (N_11590,N_10606,N_9939);
or U11591 (N_11591,N_9825,N_10045);
or U11592 (N_11592,N_9997,N_10087);
or U11593 (N_11593,N_10798,N_9768);
or U11594 (N_11594,N_10496,N_9931);
and U11595 (N_11595,N_10089,N_10071);
or U11596 (N_11596,N_9912,N_10758);
xor U11597 (N_11597,N_10589,N_10070);
and U11598 (N_11598,N_10646,N_10490);
xnor U11599 (N_11599,N_10579,N_9937);
and U11600 (N_11600,N_10426,N_10311);
nor U11601 (N_11601,N_9825,N_9652);
or U11602 (N_11602,N_10328,N_10125);
nand U11603 (N_11603,N_10186,N_9834);
and U11604 (N_11604,N_10445,N_9965);
nor U11605 (N_11605,N_9972,N_9825);
and U11606 (N_11606,N_10324,N_10419);
nand U11607 (N_11607,N_10319,N_10358);
or U11608 (N_11608,N_10098,N_9713);
nand U11609 (N_11609,N_9701,N_9696);
nand U11610 (N_11610,N_10015,N_9643);
or U11611 (N_11611,N_9746,N_9811);
xor U11612 (N_11612,N_9604,N_10373);
nor U11613 (N_11613,N_10742,N_10639);
nor U11614 (N_11614,N_10349,N_10213);
or U11615 (N_11615,N_9782,N_10149);
or U11616 (N_11616,N_10539,N_10545);
xor U11617 (N_11617,N_10161,N_10634);
nand U11618 (N_11618,N_10414,N_10379);
or U11619 (N_11619,N_10544,N_10621);
and U11620 (N_11620,N_10509,N_10401);
nand U11621 (N_11621,N_10588,N_10164);
and U11622 (N_11622,N_10630,N_9767);
and U11623 (N_11623,N_10114,N_9673);
or U11624 (N_11624,N_9787,N_10176);
or U11625 (N_11625,N_10685,N_10453);
and U11626 (N_11626,N_10428,N_10038);
nand U11627 (N_11627,N_10107,N_10217);
and U11628 (N_11628,N_9703,N_10278);
nand U11629 (N_11629,N_10199,N_10785);
and U11630 (N_11630,N_10365,N_9923);
xor U11631 (N_11631,N_10551,N_9893);
or U11632 (N_11632,N_10703,N_9967);
nor U11633 (N_11633,N_10163,N_10499);
xor U11634 (N_11634,N_9809,N_10034);
nor U11635 (N_11635,N_9917,N_10544);
nor U11636 (N_11636,N_10695,N_10572);
and U11637 (N_11637,N_10577,N_9870);
or U11638 (N_11638,N_10278,N_10497);
or U11639 (N_11639,N_10609,N_9668);
nand U11640 (N_11640,N_10136,N_9845);
and U11641 (N_11641,N_10158,N_9801);
xor U11642 (N_11642,N_9919,N_9736);
or U11643 (N_11643,N_10284,N_10492);
xor U11644 (N_11644,N_9780,N_9636);
and U11645 (N_11645,N_10500,N_10709);
nor U11646 (N_11646,N_9786,N_9779);
or U11647 (N_11647,N_10598,N_9604);
and U11648 (N_11648,N_10628,N_10436);
or U11649 (N_11649,N_10506,N_9846);
or U11650 (N_11650,N_9978,N_10042);
or U11651 (N_11651,N_10657,N_10645);
and U11652 (N_11652,N_10518,N_10697);
nor U11653 (N_11653,N_9659,N_10288);
xor U11654 (N_11654,N_10180,N_10681);
nor U11655 (N_11655,N_10272,N_10132);
or U11656 (N_11656,N_10493,N_10178);
nor U11657 (N_11657,N_10584,N_10006);
or U11658 (N_11658,N_9971,N_9704);
nand U11659 (N_11659,N_9701,N_10253);
nor U11660 (N_11660,N_10281,N_10782);
nor U11661 (N_11661,N_10226,N_10408);
xnor U11662 (N_11662,N_9630,N_10130);
nand U11663 (N_11663,N_10767,N_10515);
nor U11664 (N_11664,N_9909,N_10473);
nand U11665 (N_11665,N_9797,N_9996);
nand U11666 (N_11666,N_10284,N_10007);
xnor U11667 (N_11667,N_10210,N_10097);
xor U11668 (N_11668,N_10662,N_10229);
and U11669 (N_11669,N_9825,N_10622);
xnor U11670 (N_11670,N_10196,N_10423);
nor U11671 (N_11671,N_10206,N_9633);
or U11672 (N_11672,N_10124,N_10290);
nand U11673 (N_11673,N_9791,N_9886);
and U11674 (N_11674,N_9602,N_10059);
nand U11675 (N_11675,N_10376,N_10723);
nand U11676 (N_11676,N_10279,N_9954);
or U11677 (N_11677,N_10673,N_10180);
nor U11678 (N_11678,N_10391,N_10632);
nand U11679 (N_11679,N_10208,N_9876);
nand U11680 (N_11680,N_9907,N_9664);
nand U11681 (N_11681,N_10743,N_10099);
nor U11682 (N_11682,N_10014,N_9892);
and U11683 (N_11683,N_10284,N_10102);
or U11684 (N_11684,N_10626,N_10631);
nand U11685 (N_11685,N_10126,N_9731);
or U11686 (N_11686,N_10045,N_9867);
nor U11687 (N_11687,N_10663,N_10745);
nand U11688 (N_11688,N_9901,N_10636);
and U11689 (N_11689,N_10273,N_9901);
xor U11690 (N_11690,N_10039,N_9775);
and U11691 (N_11691,N_10637,N_9873);
or U11692 (N_11692,N_9826,N_10307);
xor U11693 (N_11693,N_9884,N_10341);
xnor U11694 (N_11694,N_10156,N_10124);
xnor U11695 (N_11695,N_10541,N_10547);
nor U11696 (N_11696,N_10424,N_9943);
nand U11697 (N_11697,N_10072,N_9601);
or U11698 (N_11698,N_10385,N_9662);
xnor U11699 (N_11699,N_9606,N_10607);
nor U11700 (N_11700,N_10437,N_9818);
nand U11701 (N_11701,N_10761,N_10063);
xor U11702 (N_11702,N_9633,N_10723);
xnor U11703 (N_11703,N_10638,N_9621);
xnor U11704 (N_11704,N_9681,N_9754);
xor U11705 (N_11705,N_10783,N_9842);
nor U11706 (N_11706,N_10002,N_10630);
and U11707 (N_11707,N_10190,N_9780);
or U11708 (N_11708,N_9699,N_10600);
or U11709 (N_11709,N_9857,N_9672);
nand U11710 (N_11710,N_9601,N_9746);
xnor U11711 (N_11711,N_9671,N_9847);
or U11712 (N_11712,N_10289,N_9901);
nor U11713 (N_11713,N_10589,N_9673);
or U11714 (N_11714,N_9653,N_10746);
or U11715 (N_11715,N_9646,N_9839);
or U11716 (N_11716,N_10113,N_10642);
nor U11717 (N_11717,N_10112,N_9894);
xor U11718 (N_11718,N_9989,N_9903);
nor U11719 (N_11719,N_9780,N_10663);
or U11720 (N_11720,N_10258,N_10646);
and U11721 (N_11721,N_9617,N_10770);
nor U11722 (N_11722,N_9971,N_10388);
or U11723 (N_11723,N_9818,N_9605);
or U11724 (N_11724,N_10581,N_10096);
xnor U11725 (N_11725,N_10416,N_10257);
or U11726 (N_11726,N_10459,N_10144);
and U11727 (N_11727,N_9888,N_10663);
xor U11728 (N_11728,N_10034,N_10017);
or U11729 (N_11729,N_10138,N_10478);
or U11730 (N_11730,N_10655,N_10467);
nor U11731 (N_11731,N_9809,N_9982);
and U11732 (N_11732,N_10229,N_10321);
nand U11733 (N_11733,N_10721,N_10136);
nor U11734 (N_11734,N_9851,N_10443);
nor U11735 (N_11735,N_10126,N_10271);
xor U11736 (N_11736,N_10403,N_9908);
xnor U11737 (N_11737,N_10460,N_9668);
xnor U11738 (N_11738,N_10169,N_10189);
xnor U11739 (N_11739,N_10285,N_10650);
and U11740 (N_11740,N_10036,N_9903);
or U11741 (N_11741,N_9983,N_10086);
or U11742 (N_11742,N_9679,N_10510);
nor U11743 (N_11743,N_10529,N_10724);
and U11744 (N_11744,N_10573,N_10239);
xor U11745 (N_11745,N_9676,N_10238);
or U11746 (N_11746,N_9744,N_10331);
nand U11747 (N_11747,N_10423,N_9700);
nand U11748 (N_11748,N_10779,N_9900);
or U11749 (N_11749,N_9989,N_10488);
xor U11750 (N_11750,N_10712,N_10441);
nor U11751 (N_11751,N_9869,N_10694);
and U11752 (N_11752,N_9876,N_10427);
nor U11753 (N_11753,N_9621,N_9941);
xor U11754 (N_11754,N_9981,N_10421);
nor U11755 (N_11755,N_10659,N_10130);
and U11756 (N_11756,N_9792,N_10221);
xnor U11757 (N_11757,N_10202,N_9681);
nor U11758 (N_11758,N_9685,N_10736);
nand U11759 (N_11759,N_10058,N_10182);
nor U11760 (N_11760,N_10528,N_10054);
and U11761 (N_11761,N_10649,N_10729);
nor U11762 (N_11762,N_9664,N_10624);
or U11763 (N_11763,N_9856,N_10557);
and U11764 (N_11764,N_10018,N_10603);
or U11765 (N_11765,N_10013,N_10227);
nand U11766 (N_11766,N_9637,N_10046);
nor U11767 (N_11767,N_9671,N_10089);
nor U11768 (N_11768,N_9745,N_9927);
and U11769 (N_11769,N_10182,N_10196);
or U11770 (N_11770,N_10261,N_10720);
nand U11771 (N_11771,N_9696,N_10524);
xnor U11772 (N_11772,N_9923,N_10230);
or U11773 (N_11773,N_9742,N_10798);
or U11774 (N_11774,N_9884,N_9651);
or U11775 (N_11775,N_10134,N_10458);
and U11776 (N_11776,N_10299,N_9611);
nand U11777 (N_11777,N_9757,N_10184);
xnor U11778 (N_11778,N_10284,N_10383);
nand U11779 (N_11779,N_10193,N_9885);
nor U11780 (N_11780,N_10205,N_10708);
xnor U11781 (N_11781,N_9965,N_10725);
nor U11782 (N_11782,N_9903,N_10314);
nor U11783 (N_11783,N_9846,N_10011);
nor U11784 (N_11784,N_10792,N_10142);
xnor U11785 (N_11785,N_10031,N_10476);
or U11786 (N_11786,N_10389,N_10411);
nor U11787 (N_11787,N_10461,N_10631);
nand U11788 (N_11788,N_10785,N_10788);
and U11789 (N_11789,N_10461,N_10347);
and U11790 (N_11790,N_10409,N_10008);
and U11791 (N_11791,N_10140,N_10227);
xor U11792 (N_11792,N_9865,N_10761);
and U11793 (N_11793,N_10436,N_10768);
nand U11794 (N_11794,N_10201,N_10172);
or U11795 (N_11795,N_10453,N_9846);
or U11796 (N_11796,N_10023,N_10189);
nand U11797 (N_11797,N_9981,N_10464);
nand U11798 (N_11798,N_9883,N_10517);
xnor U11799 (N_11799,N_9881,N_10204);
or U11800 (N_11800,N_9858,N_10111);
or U11801 (N_11801,N_10281,N_10505);
and U11802 (N_11802,N_9762,N_10574);
and U11803 (N_11803,N_9921,N_10516);
or U11804 (N_11804,N_10353,N_10566);
nor U11805 (N_11805,N_10677,N_9902);
xor U11806 (N_11806,N_9841,N_10023);
and U11807 (N_11807,N_10130,N_9912);
xor U11808 (N_11808,N_9869,N_9849);
nor U11809 (N_11809,N_10480,N_10427);
and U11810 (N_11810,N_9784,N_10221);
nor U11811 (N_11811,N_10200,N_9860);
and U11812 (N_11812,N_10451,N_9771);
xor U11813 (N_11813,N_9732,N_10608);
nand U11814 (N_11814,N_9970,N_10747);
xnor U11815 (N_11815,N_9799,N_9720);
or U11816 (N_11816,N_10106,N_9774);
nor U11817 (N_11817,N_10354,N_10338);
or U11818 (N_11818,N_10076,N_10660);
nor U11819 (N_11819,N_10365,N_10041);
nor U11820 (N_11820,N_10317,N_9680);
xnor U11821 (N_11821,N_10736,N_10077);
and U11822 (N_11822,N_9893,N_9648);
xnor U11823 (N_11823,N_10756,N_9727);
nand U11824 (N_11824,N_10027,N_10271);
nor U11825 (N_11825,N_9714,N_10786);
xnor U11826 (N_11826,N_9745,N_10673);
xnor U11827 (N_11827,N_9978,N_9716);
xnor U11828 (N_11828,N_9816,N_9653);
or U11829 (N_11829,N_10185,N_10300);
nand U11830 (N_11830,N_10680,N_9962);
nand U11831 (N_11831,N_10139,N_9969);
nand U11832 (N_11832,N_10765,N_10684);
and U11833 (N_11833,N_10168,N_10073);
nand U11834 (N_11834,N_10054,N_9806);
xor U11835 (N_11835,N_9983,N_9607);
or U11836 (N_11836,N_10648,N_10191);
or U11837 (N_11837,N_10119,N_10124);
xnor U11838 (N_11838,N_9902,N_10280);
or U11839 (N_11839,N_10279,N_10678);
or U11840 (N_11840,N_10476,N_10298);
and U11841 (N_11841,N_9913,N_10109);
and U11842 (N_11842,N_10702,N_10701);
nor U11843 (N_11843,N_10697,N_10339);
nand U11844 (N_11844,N_10609,N_9897);
nor U11845 (N_11845,N_9934,N_10701);
xor U11846 (N_11846,N_9617,N_10583);
xor U11847 (N_11847,N_9995,N_10131);
and U11848 (N_11848,N_9931,N_10505);
xor U11849 (N_11849,N_10723,N_9813);
nand U11850 (N_11850,N_10585,N_9714);
or U11851 (N_11851,N_10639,N_10705);
xor U11852 (N_11852,N_10654,N_9900);
xnor U11853 (N_11853,N_9799,N_10282);
or U11854 (N_11854,N_10136,N_10588);
nor U11855 (N_11855,N_10520,N_10649);
or U11856 (N_11856,N_9607,N_9819);
and U11857 (N_11857,N_9673,N_10523);
nand U11858 (N_11858,N_10515,N_10252);
nor U11859 (N_11859,N_10304,N_10765);
and U11860 (N_11860,N_10409,N_10206);
or U11861 (N_11861,N_10374,N_10519);
nand U11862 (N_11862,N_9679,N_9770);
nand U11863 (N_11863,N_10364,N_9984);
and U11864 (N_11864,N_10211,N_9886);
or U11865 (N_11865,N_10776,N_10461);
nor U11866 (N_11866,N_9827,N_9983);
nand U11867 (N_11867,N_10212,N_9987);
and U11868 (N_11868,N_9946,N_10259);
xor U11869 (N_11869,N_10122,N_10510);
or U11870 (N_11870,N_10008,N_10677);
or U11871 (N_11871,N_10112,N_9806);
nand U11872 (N_11872,N_10259,N_10121);
and U11873 (N_11873,N_9953,N_10176);
nand U11874 (N_11874,N_10741,N_10221);
nand U11875 (N_11875,N_10552,N_9933);
nor U11876 (N_11876,N_10010,N_9909);
or U11877 (N_11877,N_9865,N_9831);
xnor U11878 (N_11878,N_10140,N_9720);
and U11879 (N_11879,N_10732,N_10766);
nand U11880 (N_11880,N_10701,N_10646);
nor U11881 (N_11881,N_10617,N_10056);
or U11882 (N_11882,N_10438,N_9660);
nor U11883 (N_11883,N_10065,N_10669);
or U11884 (N_11884,N_10373,N_9640);
xor U11885 (N_11885,N_10790,N_10771);
xnor U11886 (N_11886,N_9738,N_9898);
nor U11887 (N_11887,N_10531,N_9970);
nor U11888 (N_11888,N_9940,N_10557);
and U11889 (N_11889,N_9774,N_9741);
or U11890 (N_11890,N_9755,N_10670);
xor U11891 (N_11891,N_10013,N_10682);
xnor U11892 (N_11892,N_10530,N_10773);
and U11893 (N_11893,N_10416,N_10259);
nor U11894 (N_11894,N_10183,N_9752);
xnor U11895 (N_11895,N_10140,N_10019);
and U11896 (N_11896,N_10288,N_9942);
nor U11897 (N_11897,N_9892,N_9792);
xnor U11898 (N_11898,N_9792,N_10057);
nand U11899 (N_11899,N_10326,N_10263);
nor U11900 (N_11900,N_10014,N_10529);
xnor U11901 (N_11901,N_10449,N_10344);
and U11902 (N_11902,N_9861,N_10042);
nor U11903 (N_11903,N_9995,N_10149);
or U11904 (N_11904,N_10676,N_10725);
or U11905 (N_11905,N_10595,N_9720);
and U11906 (N_11906,N_9968,N_10490);
and U11907 (N_11907,N_9684,N_9677);
nand U11908 (N_11908,N_9750,N_10464);
and U11909 (N_11909,N_10678,N_10100);
nand U11910 (N_11910,N_9913,N_10240);
or U11911 (N_11911,N_10607,N_9800);
nand U11912 (N_11912,N_9808,N_9731);
and U11913 (N_11913,N_10775,N_10299);
nor U11914 (N_11914,N_10235,N_10756);
nand U11915 (N_11915,N_10454,N_9794);
and U11916 (N_11916,N_10609,N_9835);
xnor U11917 (N_11917,N_10638,N_9670);
nand U11918 (N_11918,N_10554,N_10642);
or U11919 (N_11919,N_9969,N_9643);
or U11920 (N_11920,N_10636,N_10107);
and U11921 (N_11921,N_9838,N_10214);
nor U11922 (N_11922,N_10440,N_10562);
nand U11923 (N_11923,N_9611,N_10363);
nor U11924 (N_11924,N_9948,N_10182);
nand U11925 (N_11925,N_10561,N_10377);
nand U11926 (N_11926,N_9881,N_9979);
xor U11927 (N_11927,N_9950,N_9737);
nor U11928 (N_11928,N_9600,N_10378);
or U11929 (N_11929,N_10697,N_10039);
nor U11930 (N_11930,N_10685,N_10727);
or U11931 (N_11931,N_9692,N_10702);
or U11932 (N_11932,N_10465,N_9625);
xor U11933 (N_11933,N_10024,N_10288);
nand U11934 (N_11934,N_10656,N_9602);
and U11935 (N_11935,N_10449,N_9825);
and U11936 (N_11936,N_10218,N_10354);
nor U11937 (N_11937,N_10415,N_10518);
or U11938 (N_11938,N_10474,N_9899);
nor U11939 (N_11939,N_10124,N_10557);
nand U11940 (N_11940,N_9737,N_9796);
and U11941 (N_11941,N_9925,N_10699);
and U11942 (N_11942,N_9957,N_10687);
nand U11943 (N_11943,N_10038,N_10254);
xnor U11944 (N_11944,N_9844,N_10090);
or U11945 (N_11945,N_9893,N_9972);
xnor U11946 (N_11946,N_9661,N_10345);
nand U11947 (N_11947,N_9865,N_10079);
xnor U11948 (N_11948,N_10097,N_10693);
and U11949 (N_11949,N_10724,N_10346);
and U11950 (N_11950,N_9821,N_10612);
nand U11951 (N_11951,N_10243,N_9680);
nand U11952 (N_11952,N_9941,N_10158);
and U11953 (N_11953,N_10477,N_9709);
xnor U11954 (N_11954,N_10414,N_10718);
xor U11955 (N_11955,N_10179,N_9796);
or U11956 (N_11956,N_9711,N_10391);
or U11957 (N_11957,N_10584,N_10173);
or U11958 (N_11958,N_9825,N_10487);
or U11959 (N_11959,N_10460,N_10368);
nor U11960 (N_11960,N_9742,N_10112);
xnor U11961 (N_11961,N_10190,N_10262);
nand U11962 (N_11962,N_10515,N_10139);
nand U11963 (N_11963,N_9775,N_9734);
xnor U11964 (N_11964,N_10571,N_9671);
and U11965 (N_11965,N_10503,N_9922);
and U11966 (N_11966,N_9735,N_9978);
nand U11967 (N_11967,N_10251,N_10015);
xnor U11968 (N_11968,N_10075,N_10184);
or U11969 (N_11969,N_10537,N_10556);
and U11970 (N_11970,N_10612,N_9840);
nand U11971 (N_11971,N_10455,N_9708);
or U11972 (N_11972,N_10171,N_9758);
and U11973 (N_11973,N_10627,N_9861);
or U11974 (N_11974,N_10734,N_9767);
xor U11975 (N_11975,N_9660,N_10047);
or U11976 (N_11976,N_10732,N_9811);
nor U11977 (N_11977,N_9807,N_10102);
nor U11978 (N_11978,N_10176,N_9733);
and U11979 (N_11979,N_10767,N_10110);
nor U11980 (N_11980,N_10242,N_10051);
nand U11981 (N_11981,N_10241,N_9688);
nand U11982 (N_11982,N_9669,N_10223);
or U11983 (N_11983,N_10618,N_9965);
nand U11984 (N_11984,N_9888,N_10192);
nor U11985 (N_11985,N_10468,N_10096);
and U11986 (N_11986,N_9643,N_9669);
nand U11987 (N_11987,N_9687,N_9939);
nand U11988 (N_11988,N_10444,N_10476);
and U11989 (N_11989,N_10439,N_9968);
nor U11990 (N_11990,N_9651,N_10795);
nand U11991 (N_11991,N_10044,N_10582);
xor U11992 (N_11992,N_9614,N_9927);
and U11993 (N_11993,N_10681,N_9987);
nor U11994 (N_11994,N_10666,N_10712);
nor U11995 (N_11995,N_10418,N_10674);
nand U11996 (N_11996,N_10026,N_10742);
nor U11997 (N_11997,N_9901,N_9739);
nor U11998 (N_11998,N_10176,N_9768);
nor U11999 (N_11999,N_10774,N_10729);
nor U12000 (N_12000,N_10870,N_11367);
nand U12001 (N_12001,N_10810,N_10998);
or U12002 (N_12002,N_11306,N_11038);
nand U12003 (N_12003,N_10853,N_11819);
nor U12004 (N_12004,N_11220,N_11424);
nand U12005 (N_12005,N_11432,N_11611);
or U12006 (N_12006,N_11155,N_11666);
xor U12007 (N_12007,N_10817,N_11057);
or U12008 (N_12008,N_11095,N_11735);
nand U12009 (N_12009,N_11516,N_11435);
and U12010 (N_12010,N_11518,N_11282);
xnor U12011 (N_12011,N_11201,N_11903);
nor U12012 (N_12012,N_11817,N_11189);
or U12013 (N_12013,N_11450,N_11795);
and U12014 (N_12014,N_11254,N_11778);
and U12015 (N_12015,N_11953,N_11608);
and U12016 (N_12016,N_10949,N_10940);
and U12017 (N_12017,N_11933,N_11899);
nand U12018 (N_12018,N_11105,N_11579);
and U12019 (N_12019,N_10936,N_11229);
xnor U12020 (N_12020,N_11618,N_11074);
or U12021 (N_12021,N_11131,N_11414);
or U12022 (N_12022,N_11524,N_10830);
nand U12023 (N_12023,N_11695,N_10878);
nand U12024 (N_12024,N_11909,N_11571);
and U12025 (N_12025,N_11764,N_11122);
or U12026 (N_12026,N_10967,N_11931);
and U12027 (N_12027,N_11321,N_11939);
nand U12028 (N_12028,N_11420,N_11697);
or U12029 (N_12029,N_11183,N_11228);
and U12030 (N_12030,N_11827,N_11556);
and U12031 (N_12031,N_11001,N_11459);
nand U12032 (N_12032,N_11896,N_11215);
xnor U12033 (N_12033,N_11015,N_11716);
nor U12034 (N_12034,N_11974,N_10952);
xnor U12035 (N_12035,N_11784,N_11096);
nor U12036 (N_12036,N_11411,N_11945);
and U12037 (N_12037,N_11777,N_11685);
nand U12038 (N_12038,N_11438,N_11062);
and U12039 (N_12039,N_10814,N_10816);
xnor U12040 (N_12040,N_11546,N_11822);
nand U12041 (N_12041,N_10825,N_11493);
xor U12042 (N_12042,N_11690,N_11728);
and U12043 (N_12043,N_11508,N_11651);
and U12044 (N_12044,N_10843,N_10927);
nor U12045 (N_12045,N_10903,N_11068);
xor U12046 (N_12046,N_11686,N_11146);
and U12047 (N_12047,N_11761,N_11341);
xnor U12048 (N_12048,N_10954,N_11710);
nor U12049 (N_12049,N_11515,N_11967);
and U12050 (N_12050,N_11045,N_11835);
or U12051 (N_12051,N_11482,N_11771);
xor U12052 (N_12052,N_11117,N_11989);
nand U12053 (N_12053,N_11499,N_11732);
xor U12054 (N_12054,N_11924,N_11354);
nand U12055 (N_12055,N_11997,N_10989);
and U12056 (N_12056,N_11553,N_11998);
xor U12057 (N_12057,N_11335,N_11665);
nor U12058 (N_12058,N_11512,N_11090);
xor U12059 (N_12059,N_11600,N_11312);
xnor U12060 (N_12060,N_11613,N_11153);
nor U12061 (N_12061,N_10812,N_10963);
xnor U12062 (N_12062,N_11136,N_10898);
xor U12063 (N_12063,N_11169,N_11980);
nor U12064 (N_12064,N_11339,N_10871);
nor U12065 (N_12065,N_11483,N_11452);
xnor U12066 (N_12066,N_10934,N_11680);
and U12067 (N_12067,N_11102,N_11806);
xnor U12068 (N_12068,N_11921,N_11112);
and U12069 (N_12069,N_11663,N_10834);
nand U12070 (N_12070,N_11872,N_11789);
nor U12071 (N_12071,N_11564,N_11058);
nor U12072 (N_12072,N_11689,N_11907);
or U12073 (N_12073,N_11776,N_11317);
and U12074 (N_12074,N_10938,N_11113);
and U12075 (N_12075,N_11679,N_10953);
nand U12076 (N_12076,N_10966,N_11867);
and U12077 (N_12077,N_11384,N_11466);
and U12078 (N_12078,N_11478,N_11328);
or U12079 (N_12079,N_10857,N_10986);
nand U12080 (N_12080,N_11506,N_10991);
and U12081 (N_12081,N_10947,N_11467);
xnor U12082 (N_12082,N_10976,N_11233);
nand U12083 (N_12083,N_11104,N_11902);
xnor U12084 (N_12084,N_10868,N_11079);
xnor U12085 (N_12085,N_11775,N_11623);
and U12086 (N_12086,N_11368,N_11133);
and U12087 (N_12087,N_11440,N_10961);
nor U12088 (N_12088,N_11536,N_11436);
xnor U12089 (N_12089,N_11575,N_11390);
and U12090 (N_12090,N_11831,N_10856);
or U12091 (N_12091,N_11444,N_11533);
and U12092 (N_12092,N_11805,N_11917);
nor U12093 (N_12093,N_10841,N_11069);
nor U12094 (N_12094,N_11260,N_11812);
and U12095 (N_12095,N_11358,N_11299);
xnor U12096 (N_12096,N_11446,N_11811);
xnor U12097 (N_12097,N_11044,N_11346);
and U12098 (N_12098,N_11619,N_11401);
xor U12099 (N_12099,N_11007,N_11056);
nor U12100 (N_12100,N_11036,N_11176);
or U12101 (N_12101,N_10854,N_10877);
and U12102 (N_12102,N_11668,N_11486);
nor U12103 (N_12103,N_11570,N_10839);
xor U12104 (N_12104,N_10836,N_11647);
or U12105 (N_12105,N_11398,N_11863);
and U12106 (N_12106,N_10804,N_11930);
and U12107 (N_12107,N_11983,N_11362);
and U12108 (N_12108,N_11743,N_11754);
nor U12109 (N_12109,N_11519,N_11677);
xnor U12110 (N_12110,N_11675,N_11239);
nor U12111 (N_12111,N_11526,N_11272);
and U12112 (N_12112,N_11294,N_11204);
nor U12113 (N_12113,N_11409,N_11264);
and U12114 (N_12114,N_11563,N_11203);
or U12115 (N_12115,N_11151,N_11433);
nor U12116 (N_12116,N_10892,N_11923);
and U12117 (N_12117,N_11916,N_11365);
and U12118 (N_12118,N_10888,N_11985);
and U12119 (N_12119,N_10842,N_11373);
or U12120 (N_12120,N_11938,N_11879);
nand U12121 (N_12121,N_11502,N_11807);
nand U12122 (N_12122,N_11005,N_11455);
xnor U12123 (N_12123,N_11972,N_11262);
and U12124 (N_12124,N_11332,N_11150);
xor U12125 (N_12125,N_11173,N_11091);
nor U12126 (N_12126,N_11491,N_11253);
nand U12127 (N_12127,N_11824,N_11361);
nand U12128 (N_12128,N_11773,N_11925);
nand U12129 (N_12129,N_11108,N_11061);
nand U12130 (N_12130,N_11947,N_10815);
or U12131 (N_12131,N_10968,N_11785);
xor U12132 (N_12132,N_11142,N_11576);
nor U12133 (N_12133,N_11936,N_11656);
or U12134 (N_12134,N_11664,N_11298);
or U12135 (N_12135,N_11525,N_11520);
or U12136 (N_12136,N_10926,N_11223);
or U12137 (N_12137,N_11303,N_11587);
or U12138 (N_12138,N_11674,N_11628);
and U12139 (N_12139,N_11219,N_10801);
and U12140 (N_12140,N_11441,N_11696);
nand U12141 (N_12141,N_11759,N_11029);
xnor U12142 (N_12142,N_10981,N_11760);
nor U12143 (N_12143,N_10914,N_11190);
xor U12144 (N_12144,N_11964,N_11503);
or U12145 (N_12145,N_11406,N_11024);
nor U12146 (N_12146,N_11393,N_11713);
nand U12147 (N_12147,N_11999,N_11198);
or U12148 (N_12148,N_11707,N_10946);
and U12149 (N_12149,N_11946,N_11137);
nand U12150 (N_12150,N_11145,N_10880);
xnor U12151 (N_12151,N_10941,N_11315);
and U12152 (N_12152,N_11577,N_11046);
xor U12153 (N_12153,N_11331,N_11227);
xor U12154 (N_12154,N_11720,N_11510);
and U12155 (N_12155,N_11369,N_10851);
nor U12156 (N_12156,N_11605,N_11192);
xor U12157 (N_12157,N_11070,N_11421);
or U12158 (N_12158,N_11359,N_11217);
nor U12159 (N_12159,N_10932,N_11606);
nand U12160 (N_12160,N_11681,N_11382);
nor U12161 (N_12161,N_11084,N_10866);
or U12162 (N_12162,N_11087,N_11181);
or U12163 (N_12163,N_11555,N_11366);
xor U12164 (N_12164,N_11951,N_10979);
or U12165 (N_12165,N_11395,N_11729);
and U12166 (N_12166,N_11780,N_11292);
or U12167 (N_12167,N_11767,N_10884);
nor U12168 (N_12168,N_11174,N_11672);
nor U12169 (N_12169,N_11415,N_11265);
nand U12170 (N_12170,N_11968,N_11639);
or U12171 (N_12171,N_11742,N_11170);
nand U12172 (N_12172,N_11871,N_11197);
and U12173 (N_12173,N_11635,N_11314);
and U12174 (N_12174,N_10919,N_11073);
or U12175 (N_12175,N_11320,N_11988);
nor U12176 (N_12176,N_11374,N_11900);
xor U12177 (N_12177,N_11866,N_11032);
xnor U12178 (N_12178,N_11127,N_11528);
nand U12179 (N_12179,N_11285,N_11881);
and U12180 (N_12180,N_11347,N_11271);
xnor U12181 (N_12181,N_11781,N_11590);
xnor U12182 (N_12182,N_10827,N_11574);
xnor U12183 (N_12183,N_11402,N_11592);
xnor U12184 (N_12184,N_11910,N_11251);
xnor U12185 (N_12185,N_11869,N_11706);
xnor U12186 (N_12186,N_11667,N_10855);
nand U12187 (N_12187,N_11929,N_11678);
xor U12188 (N_12188,N_11256,N_11427);
or U12189 (N_12189,N_11698,N_11889);
or U12190 (N_12190,N_10901,N_11744);
and U12191 (N_12191,N_11818,N_11165);
and U12192 (N_12192,N_11230,N_11969);
and U12193 (N_12193,N_11753,N_10803);
nor U12194 (N_12194,N_11158,N_11934);
and U12195 (N_12195,N_11786,N_11034);
nand U12196 (N_12196,N_11263,N_11476);
nor U12197 (N_12197,N_11085,N_11031);
or U12198 (N_12198,N_11614,N_11283);
nand U12199 (N_12199,N_10974,N_11166);
nor U12200 (N_12200,N_11652,N_11477);
and U12201 (N_12201,N_11211,N_11385);
and U12202 (N_12202,N_11210,N_11958);
or U12203 (N_12203,N_11304,N_11751);
nor U12204 (N_12204,N_11003,N_11645);
nand U12205 (N_12205,N_10905,N_11126);
nand U12206 (N_12206,N_10860,N_11100);
or U12207 (N_12207,N_11948,N_11157);
nor U12208 (N_12208,N_11193,N_11319);
xnor U12209 (N_12209,N_11877,N_11952);
xnor U12210 (N_12210,N_11991,N_11589);
or U12211 (N_12211,N_11124,N_11171);
or U12212 (N_12212,N_11699,N_10820);
or U12213 (N_12213,N_11722,N_11023);
and U12214 (N_12214,N_11487,N_11457);
nand U12215 (N_12215,N_11966,N_10818);
nand U12216 (N_12216,N_11177,N_11008);
or U12217 (N_12217,N_11631,N_11880);
and U12218 (N_12218,N_11638,N_11212);
or U12219 (N_12219,N_10959,N_11248);
xnor U12220 (N_12220,N_11572,N_11990);
or U12221 (N_12221,N_11655,N_11268);
and U12222 (N_12222,N_11598,N_10844);
xor U12223 (N_12223,N_11801,N_11858);
nor U12224 (N_12224,N_11730,N_11957);
xnor U12225 (N_12225,N_11609,N_11116);
or U12226 (N_12226,N_11965,N_11118);
nand U12227 (N_12227,N_11098,N_10945);
and U12228 (N_12228,N_11996,N_11379);
and U12229 (N_12229,N_11800,N_10918);
xnor U12230 (N_12230,N_11511,N_11794);
nand U12231 (N_12231,N_11372,N_11599);
and U12232 (N_12232,N_10806,N_11097);
nand U12233 (N_12233,N_11883,N_11154);
or U12234 (N_12234,N_11344,N_11002);
and U12235 (N_12235,N_11757,N_11531);
or U12236 (N_12236,N_11895,N_11718);
and U12237 (N_12237,N_11026,N_11629);
and U12238 (N_12238,N_11654,N_11963);
nor U12239 (N_12239,N_11391,N_11245);
xor U12240 (N_12240,N_11027,N_11237);
or U12241 (N_12241,N_11746,N_10916);
nor U12242 (N_12242,N_11509,N_11465);
nor U12243 (N_12243,N_11621,N_11121);
xor U12244 (N_12244,N_11033,N_11540);
or U12245 (N_12245,N_11364,N_11261);
xnor U12246 (N_12246,N_11030,N_11363);
nor U12247 (N_12247,N_11567,N_11529);
xnor U12248 (N_12248,N_11669,N_11496);
nand U12249 (N_12249,N_11135,N_11139);
xnor U12250 (N_12250,N_10802,N_11394);
nand U12251 (N_12251,N_11000,N_11025);
nor U12252 (N_12252,N_11642,N_11782);
nand U12253 (N_12253,N_11184,N_11982);
nor U12254 (N_12254,N_11423,N_11724);
xor U12255 (N_12255,N_11080,N_11114);
nor U12256 (N_12256,N_11843,N_10873);
xor U12257 (N_12257,N_10811,N_11826);
nor U12258 (N_12258,N_10931,N_11439);
and U12259 (N_12259,N_11717,N_11047);
nor U12260 (N_12260,N_11736,N_10890);
nand U12261 (N_12261,N_11325,N_11397);
nand U12262 (N_12262,N_11296,N_11469);
nor U12263 (N_12263,N_11016,N_11560);
or U12264 (N_12264,N_11186,N_11492);
nand U12265 (N_12265,N_11521,N_11453);
xnor U12266 (N_12266,N_11961,N_11882);
or U12267 (N_12267,N_11284,N_11954);
xor U12268 (N_12268,N_11099,N_11756);
xor U12269 (N_12269,N_11497,N_11351);
or U12270 (N_12270,N_11582,N_11875);
and U12271 (N_12271,N_11081,N_11830);
or U12272 (N_12272,N_11049,N_11425);
nand U12273 (N_12273,N_11650,N_10900);
nor U12274 (N_12274,N_11232,N_11646);
nand U12275 (N_12275,N_11891,N_10970);
xnor U12276 (N_12276,N_10912,N_11376);
nor U12277 (N_12277,N_11101,N_10891);
and U12278 (N_12278,N_11235,N_11740);
or U12279 (N_12279,N_10973,N_10993);
xor U12280 (N_12280,N_11986,N_11326);
or U12281 (N_12281,N_11489,N_11813);
or U12282 (N_12282,N_10982,N_10838);
nor U12283 (N_12283,N_10956,N_11886);
and U12284 (N_12284,N_10987,N_11313);
nor U12285 (N_12285,N_10800,N_11468);
xnor U12286 (N_12286,N_11224,N_10955);
xnor U12287 (N_12287,N_11694,N_11993);
nor U12288 (N_12288,N_11148,N_10902);
xnor U12289 (N_12289,N_11648,N_11593);
or U12290 (N_12290,N_11216,N_11750);
or U12291 (N_12291,N_11859,N_11396);
or U12292 (N_12292,N_11463,N_11662);
and U12293 (N_12293,N_10889,N_11218);
nor U12294 (N_12294,N_11267,N_11448);
or U12295 (N_12295,N_11275,N_11714);
or U12296 (N_12296,N_11544,N_11625);
nor U12297 (N_12297,N_10992,N_11490);
and U12298 (N_12298,N_11597,N_11701);
nand U12299 (N_12299,N_11636,N_11532);
or U12300 (N_12300,N_11380,N_10933);
nor U12301 (N_12301,N_10983,N_10999);
xnor U12302 (N_12302,N_11857,N_10923);
nand U12303 (N_12303,N_11630,N_10847);
xor U12304 (N_12304,N_11012,N_11180);
nand U12305 (N_12305,N_10852,N_11584);
and U12306 (N_12306,N_11702,N_11734);
nand U12307 (N_12307,N_11833,N_11110);
and U12308 (N_12308,N_10997,N_11334);
or U12309 (N_12309,N_10823,N_11839);
nand U12310 (N_12310,N_11474,N_10929);
and U12311 (N_12311,N_11422,N_11092);
xor U12312 (N_12312,N_11844,N_11763);
nand U12313 (N_12313,N_11692,N_11984);
and U12314 (N_12314,N_11207,N_11851);
nor U12315 (N_12315,N_11333,N_11783);
or U12316 (N_12316,N_11289,N_10829);
or U12317 (N_12317,N_11552,N_11060);
xnor U12318 (N_12318,N_11302,N_10887);
nor U12319 (N_12319,N_11616,N_11340);
nand U12320 (N_12320,N_11622,N_11021);
and U12321 (N_12321,N_11808,N_10907);
nor U12322 (N_12322,N_11255,N_11222);
and U12323 (N_12323,N_11213,N_10960);
xor U12324 (N_12324,N_11653,N_11048);
or U12325 (N_12325,N_10809,N_11853);
nand U12326 (N_12326,N_10917,N_10928);
nand U12327 (N_12327,N_11274,N_11042);
or U12328 (N_12328,N_11887,N_11911);
nor U12329 (N_12329,N_10881,N_11484);
nor U12330 (N_12330,N_11796,N_11300);
or U12331 (N_12331,N_11799,N_11920);
nand U12332 (N_12332,N_11278,N_11175);
and U12333 (N_12333,N_11658,N_11562);
or U12334 (N_12334,N_11270,N_11551);
or U12335 (N_12335,N_10948,N_11956);
and U12336 (N_12336,N_11083,N_11103);
nand U12337 (N_12337,N_10835,N_11330);
or U12338 (N_12338,N_11381,N_11693);
nor U12339 (N_12339,N_11814,N_11399);
xor U12340 (N_12340,N_11078,N_11660);
or U12341 (N_12341,N_11410,N_11093);
and U12342 (N_12342,N_11307,N_11854);
nand U12343 (N_12343,N_11485,N_11727);
and U12344 (N_12344,N_11387,N_11684);
nor U12345 (N_12345,N_11129,N_10985);
nor U12346 (N_12346,N_11981,N_11187);
nor U12347 (N_12347,N_11975,N_11141);
nor U12348 (N_12348,N_10950,N_11733);
nor U12349 (N_12349,N_11748,N_10831);
or U12350 (N_12350,N_11052,N_11941);
and U12351 (N_12351,N_11200,N_11370);
nand U12352 (N_12352,N_11573,N_11774);
and U12353 (N_12353,N_11243,N_11534);
nor U12354 (N_12354,N_11231,N_10951);
or U12355 (N_12355,N_11168,N_10859);
nand U12356 (N_12356,N_11676,N_11726);
and U12357 (N_12357,N_11202,N_11400);
xnor U12358 (N_12358,N_11585,N_10915);
xnor U12359 (N_12359,N_11971,N_11206);
nor U12360 (N_12360,N_11244,N_11815);
nor U12361 (N_12361,N_10957,N_10893);
nand U12362 (N_12362,N_11994,N_11094);
nand U12363 (N_12363,N_11182,N_11017);
nor U12364 (N_12364,N_11741,N_11035);
or U12365 (N_12365,N_10922,N_10894);
and U12366 (N_12366,N_11357,N_11739);
nand U12367 (N_12367,N_11451,N_11310);
nand U12368 (N_12368,N_11731,N_11792);
nor U12369 (N_12369,N_10895,N_11928);
or U12370 (N_12370,N_11517,N_11594);
nor U12371 (N_12371,N_11657,N_11915);
nor U12372 (N_12372,N_11904,N_11603);
or U12373 (N_12373,N_11987,N_11935);
or U12374 (N_12374,N_11040,N_11355);
and U12375 (N_12375,N_10975,N_11138);
xnor U12376 (N_12376,N_11259,N_11067);
xnor U12377 (N_12377,N_11802,N_11225);
or U12378 (N_12378,N_11279,N_11721);
and U12379 (N_12379,N_11416,N_11063);
nor U12380 (N_12380,N_10910,N_11862);
nor U12381 (N_12381,N_11688,N_11542);
nor U12382 (N_12382,N_11336,N_11565);
or U12383 (N_12383,N_10867,N_11447);
nand U12384 (N_12384,N_11538,N_11281);
nand U12385 (N_12385,N_10813,N_10863);
nand U12386 (N_12386,N_11064,N_10861);
xnor U12387 (N_12387,N_11481,N_11790);
nand U12388 (N_12388,N_11758,N_11247);
xnor U12389 (N_12389,N_11637,N_11338);
nor U12390 (N_12390,N_11803,N_11152);
xnor U12391 (N_12391,N_11888,N_10924);
nor U12392 (N_12392,N_11712,N_11196);
or U12393 (N_12393,N_11120,N_11293);
nand U12394 (N_12394,N_11462,N_10977);
or U12395 (N_12395,N_11906,N_11345);
or U12396 (N_12396,N_11352,N_11940);
nand U12397 (N_12397,N_11290,N_10882);
or U12398 (N_12398,N_11890,N_11295);
and U12399 (N_12399,N_11445,N_11860);
or U12400 (N_12400,N_11973,N_11615);
and U12401 (N_12401,N_11456,N_10904);
nor U12402 (N_12402,N_11864,N_11075);
nor U12403 (N_12403,N_10872,N_11832);
nand U12404 (N_12404,N_11429,N_10925);
xnor U12405 (N_12405,N_10886,N_11849);
xor U12406 (N_12406,N_11149,N_11995);
or U12407 (N_12407,N_11797,N_11766);
nor U12408 (N_12408,N_11188,N_11992);
nor U12409 (N_12409,N_11897,N_11670);
xnor U12410 (N_12410,N_10906,N_11234);
or U12411 (N_12411,N_11065,N_11185);
nor U12412 (N_12412,N_11106,N_11905);
and U12413 (N_12413,N_11829,N_11318);
or U12414 (N_12414,N_11322,N_11745);
nand U12415 (N_12415,N_11348,N_11705);
and U12416 (N_12416,N_11559,N_11054);
and U12417 (N_12417,N_11874,N_11834);
and U12418 (N_12418,N_11488,N_11970);
nand U12419 (N_12419,N_11252,N_11053);
nand U12420 (N_12420,N_11641,N_11144);
or U12421 (N_12421,N_10808,N_10994);
or U12422 (N_12422,N_10876,N_11236);
or U12423 (N_12423,N_11109,N_11885);
and U12424 (N_12424,N_10846,N_11013);
and U12425 (N_12425,N_11172,N_11737);
nand U12426 (N_12426,N_11164,N_11009);
xnor U12427 (N_12427,N_10909,N_11527);
nor U12428 (N_12428,N_10920,N_10978);
and U12429 (N_12429,N_11309,N_11578);
nor U12430 (N_12430,N_11840,N_11134);
xnor U12431 (N_12431,N_10883,N_11549);
xor U12432 (N_12432,N_11942,N_11111);
and U12433 (N_12433,N_11147,N_11816);
and U12434 (N_12434,N_11226,N_11671);
nor U12435 (N_12435,N_11979,N_11434);
or U12436 (N_12436,N_11823,N_11828);
xnor U12437 (N_12437,N_10921,N_11128);
and U12438 (N_12438,N_11140,N_11848);
xnor U12439 (N_12439,N_11798,N_11386);
nor U12440 (N_12440,N_11250,N_11350);
nor U12441 (N_12441,N_11055,N_11020);
nand U12442 (N_12442,N_11494,N_11955);
nand U12443 (N_12443,N_11195,N_11537);
and U12444 (N_12444,N_11632,N_11460);
and U12445 (N_12445,N_11010,N_11943);
and U12446 (N_12446,N_10869,N_11550);
xor U12447 (N_12447,N_11554,N_11568);
xnor U12448 (N_12448,N_10805,N_11473);
nor U12449 (N_12449,N_10913,N_11051);
nor U12450 (N_12450,N_11464,N_11768);
nand U12451 (N_12451,N_10828,N_11011);
nand U12452 (N_12452,N_11107,N_11865);
nand U12453 (N_12453,N_11130,N_11119);
nor U12454 (N_12454,N_11311,N_11837);
nand U12455 (N_12455,N_11356,N_11836);
xor U12456 (N_12456,N_11076,N_11962);
nor U12457 (N_12457,N_11316,N_11868);
or U12458 (N_12458,N_11349,N_11082);
xnor U12459 (N_12459,N_11715,N_11884);
nor U12460 (N_12460,N_11431,N_11249);
xor U12461 (N_12461,N_11498,N_11583);
nand U12462 (N_12462,N_11709,N_11557);
or U12463 (N_12463,N_11847,N_11301);
xnor U12464 (N_12464,N_11541,N_11163);
and U12465 (N_12465,N_11028,N_11545);
or U12466 (N_12466,N_11626,N_10840);
or U12467 (N_12467,N_11308,N_11944);
xnor U12468 (N_12468,N_11437,N_11769);
xnor U12469 (N_12469,N_11479,N_11960);
nor U12470 (N_12470,N_11413,N_11779);
nor U12471 (N_12471,N_11530,N_11926);
and U12472 (N_12472,N_11329,N_11132);
nor U12473 (N_12473,N_11418,N_10821);
nand U12474 (N_12474,N_11949,N_11793);
nand U12475 (N_12475,N_11850,N_11738);
or U12476 (N_12476,N_11649,N_11755);
and U12477 (N_12477,N_11711,N_11612);
nand U12478 (N_12478,N_10874,N_11620);
nand U12479 (N_12479,N_11371,N_10897);
or U12480 (N_12480,N_11375,N_10995);
xor U12481 (N_12481,N_11809,N_11442);
and U12482 (N_12482,N_11687,N_11006);
xnor U12483 (N_12483,N_11586,N_11089);
nand U12484 (N_12484,N_11077,N_10879);
and U12485 (N_12485,N_11461,N_10944);
and U12486 (N_12486,N_11595,N_11159);
nand U12487 (N_12487,N_11004,N_10875);
and U12488 (N_12488,N_11430,N_11209);
and U12489 (N_12489,N_11821,N_10939);
nor U12490 (N_12490,N_11700,N_11634);
or U12491 (N_12491,N_11919,N_11072);
or U12492 (N_12492,N_11125,N_10833);
or U12493 (N_12493,N_11810,N_11428);
nor U12494 (N_12494,N_11022,N_11288);
xnor U12495 (N_12495,N_11561,N_11258);
xnor U12496 (N_12496,N_11353,N_11894);
nand U12497 (N_12497,N_11950,N_11602);
nand U12498 (N_12498,N_11276,N_11405);
nand U12499 (N_12499,N_11591,N_11238);
xnor U12500 (N_12500,N_10865,N_11914);
nor U12501 (N_12501,N_11199,N_11762);
nor U12502 (N_12502,N_10911,N_11403);
or U12503 (N_12503,N_11327,N_10819);
or U12504 (N_12504,N_11342,N_11426);
or U12505 (N_12505,N_11604,N_11392);
xnor U12506 (N_12506,N_11543,N_11846);
and U12507 (N_12507,N_11558,N_10969);
nand U12508 (N_12508,N_11208,N_11178);
xor U12509 (N_12509,N_10832,N_10845);
and U12510 (N_12510,N_11143,N_11581);
or U12511 (N_12511,N_11898,N_11507);
nand U12512 (N_12512,N_11977,N_11838);
and U12513 (N_12513,N_10996,N_11845);
nand U12514 (N_12514,N_11240,N_11901);
nor U12515 (N_12515,N_11037,N_11043);
or U12516 (N_12516,N_11673,N_11257);
xor U12517 (N_12517,N_10984,N_11160);
nand U12518 (N_12518,N_11305,N_11378);
nor U12519 (N_12519,N_10885,N_10824);
xor U12520 (N_12520,N_11870,N_11504);
and U12521 (N_12521,N_11588,N_11404);
nor U12522 (N_12522,N_10958,N_11856);
and U12523 (N_12523,N_11214,N_11324);
or U12524 (N_12524,N_11205,N_11412);
and U12525 (N_12525,N_11708,N_11388);
or U12526 (N_12526,N_11682,N_11873);
and U12527 (N_12527,N_11343,N_11918);
nor U12528 (N_12528,N_11547,N_11855);
and U12529 (N_12529,N_11765,N_10848);
or U12530 (N_12530,N_11480,N_11221);
xnor U12531 (N_12531,N_10837,N_10849);
nand U12532 (N_12532,N_11976,N_11513);
nand U12533 (N_12533,N_11419,N_11601);
nand U12534 (N_12534,N_11723,N_11912);
nand U12535 (N_12535,N_11162,N_11323);
and U12536 (N_12536,N_11514,N_10972);
nor U12537 (N_12537,N_10937,N_11280);
nor U12538 (N_12538,N_10962,N_10980);
nor U12539 (N_12539,N_11337,N_11683);
nor U12540 (N_12540,N_10971,N_11161);
xor U12541 (N_12541,N_10864,N_11389);
or U12542 (N_12542,N_11627,N_11841);
nor U12543 (N_12543,N_11842,N_11019);
nor U12544 (N_12544,N_11913,N_11286);
or U12545 (N_12545,N_11408,N_11861);
nand U12546 (N_12546,N_11937,N_11580);
xor U12547 (N_12547,N_11471,N_11458);
or U12548 (N_12548,N_11500,N_11643);
xor U12549 (N_12549,N_11659,N_11495);
or U12550 (N_12550,N_11978,N_11908);
or U12551 (N_12551,N_10822,N_11041);
nor U12552 (N_12552,N_11246,N_10930);
xnor U12553 (N_12553,N_11523,N_11569);
xor U12554 (N_12554,N_11644,N_11266);
or U12555 (N_12555,N_11661,N_11505);
nand U12556 (N_12556,N_11066,N_11548);
and U12557 (N_12557,N_11539,N_11804);
or U12558 (N_12558,N_11624,N_11059);
nor U12559 (N_12559,N_11820,N_11825);
nor U12560 (N_12560,N_11242,N_11535);
or U12561 (N_12561,N_11454,N_11273);
or U12562 (N_12562,N_11269,N_11014);
and U12563 (N_12563,N_11788,N_11691);
or U12564 (N_12564,N_11522,N_11179);
and U12565 (N_12565,N_10899,N_11704);
nand U12566 (N_12566,N_11610,N_11417);
xnor U12567 (N_12567,N_11115,N_11018);
and U12568 (N_12568,N_11852,N_11241);
xnor U12569 (N_12569,N_11893,N_11039);
xnor U12570 (N_12570,N_10935,N_11156);
and U12571 (N_12571,N_10896,N_11291);
or U12572 (N_12572,N_11922,N_11640);
nor U12573 (N_12573,N_10942,N_11297);
nor U12574 (N_12574,N_10807,N_11703);
or U12575 (N_12575,N_11607,N_11772);
nor U12576 (N_12576,N_11123,N_11407);
and U12577 (N_12577,N_11787,N_11360);
and U12578 (N_12578,N_10908,N_11277);
or U12579 (N_12579,N_11770,N_11566);
and U12580 (N_12580,N_10858,N_10990);
and U12581 (N_12581,N_11377,N_11050);
nor U12582 (N_12582,N_10862,N_11475);
nand U12583 (N_12583,N_11596,N_11747);
or U12584 (N_12584,N_11191,N_11501);
xnor U12585 (N_12585,N_11167,N_11470);
and U12586 (N_12586,N_11383,N_11194);
nor U12587 (N_12587,N_11633,N_11725);
nand U12588 (N_12588,N_10965,N_11892);
or U12589 (N_12589,N_11071,N_11719);
xnor U12590 (N_12590,N_10943,N_11927);
xnor U12591 (N_12591,N_11876,N_11878);
or U12592 (N_12592,N_11959,N_10826);
nand U12593 (N_12593,N_11287,N_11443);
or U12594 (N_12594,N_11472,N_11932);
and U12595 (N_12595,N_10964,N_11752);
or U12596 (N_12596,N_11449,N_11617);
and U12597 (N_12597,N_10850,N_11088);
nor U12598 (N_12598,N_11749,N_11791);
nand U12599 (N_12599,N_10988,N_11086);
or U12600 (N_12600,N_10933,N_11779);
and U12601 (N_12601,N_11878,N_11798);
nand U12602 (N_12602,N_11946,N_11503);
nor U12603 (N_12603,N_10970,N_11219);
nor U12604 (N_12604,N_11348,N_11418);
nand U12605 (N_12605,N_10823,N_11723);
and U12606 (N_12606,N_11145,N_11026);
nand U12607 (N_12607,N_11373,N_11799);
nor U12608 (N_12608,N_10905,N_10976);
or U12609 (N_12609,N_11484,N_11637);
nor U12610 (N_12610,N_11721,N_11222);
nand U12611 (N_12611,N_11355,N_11058);
nand U12612 (N_12612,N_11866,N_11375);
nand U12613 (N_12613,N_11113,N_11631);
or U12614 (N_12614,N_11098,N_11679);
or U12615 (N_12615,N_11516,N_11247);
xnor U12616 (N_12616,N_11168,N_11377);
or U12617 (N_12617,N_11952,N_11321);
and U12618 (N_12618,N_11372,N_11822);
and U12619 (N_12619,N_11866,N_11123);
nor U12620 (N_12620,N_10920,N_11357);
nand U12621 (N_12621,N_10923,N_11577);
xor U12622 (N_12622,N_11015,N_11069);
or U12623 (N_12623,N_11821,N_10933);
and U12624 (N_12624,N_11678,N_11662);
or U12625 (N_12625,N_11450,N_11899);
xor U12626 (N_12626,N_10988,N_10914);
or U12627 (N_12627,N_10962,N_11375);
xor U12628 (N_12628,N_11894,N_11363);
nand U12629 (N_12629,N_11869,N_11369);
xor U12630 (N_12630,N_11281,N_11698);
or U12631 (N_12631,N_11125,N_11635);
or U12632 (N_12632,N_11309,N_10893);
nand U12633 (N_12633,N_11903,N_11289);
or U12634 (N_12634,N_11458,N_11320);
or U12635 (N_12635,N_11775,N_11149);
or U12636 (N_12636,N_11874,N_11465);
or U12637 (N_12637,N_11982,N_10962);
xnor U12638 (N_12638,N_11300,N_11748);
nand U12639 (N_12639,N_11309,N_11771);
and U12640 (N_12640,N_11106,N_11656);
nand U12641 (N_12641,N_11007,N_11839);
xnor U12642 (N_12642,N_11705,N_11771);
xor U12643 (N_12643,N_10857,N_11477);
nand U12644 (N_12644,N_11440,N_11606);
and U12645 (N_12645,N_11220,N_11527);
and U12646 (N_12646,N_11508,N_11176);
nor U12647 (N_12647,N_11877,N_11019);
and U12648 (N_12648,N_11901,N_11478);
xor U12649 (N_12649,N_11398,N_10843);
nand U12650 (N_12650,N_11619,N_11847);
and U12651 (N_12651,N_11708,N_11006);
and U12652 (N_12652,N_11046,N_11732);
and U12653 (N_12653,N_11667,N_10969);
nand U12654 (N_12654,N_11625,N_11382);
xnor U12655 (N_12655,N_11023,N_11308);
nor U12656 (N_12656,N_11670,N_10964);
xor U12657 (N_12657,N_10853,N_11175);
and U12658 (N_12658,N_11880,N_11363);
nand U12659 (N_12659,N_11798,N_11421);
nor U12660 (N_12660,N_10841,N_11952);
or U12661 (N_12661,N_11933,N_11434);
nor U12662 (N_12662,N_11378,N_11384);
or U12663 (N_12663,N_11689,N_10948);
and U12664 (N_12664,N_11810,N_11639);
and U12665 (N_12665,N_11418,N_11590);
nand U12666 (N_12666,N_11127,N_11497);
nor U12667 (N_12667,N_11600,N_11346);
xnor U12668 (N_12668,N_11464,N_11796);
nor U12669 (N_12669,N_11397,N_11312);
xor U12670 (N_12670,N_11711,N_11367);
xnor U12671 (N_12671,N_11340,N_11984);
or U12672 (N_12672,N_11896,N_11617);
nor U12673 (N_12673,N_11057,N_11667);
xnor U12674 (N_12674,N_11294,N_11965);
and U12675 (N_12675,N_11901,N_11006);
xnor U12676 (N_12676,N_11428,N_11136);
or U12677 (N_12677,N_11508,N_11656);
nand U12678 (N_12678,N_10981,N_10879);
nand U12679 (N_12679,N_11951,N_11903);
nand U12680 (N_12680,N_10954,N_11681);
and U12681 (N_12681,N_10873,N_10887);
nand U12682 (N_12682,N_11880,N_10911);
xor U12683 (N_12683,N_11330,N_11873);
or U12684 (N_12684,N_11231,N_10986);
xnor U12685 (N_12685,N_11578,N_11987);
nor U12686 (N_12686,N_11401,N_11515);
nand U12687 (N_12687,N_11352,N_11175);
xnor U12688 (N_12688,N_10824,N_11976);
xnor U12689 (N_12689,N_11981,N_11713);
or U12690 (N_12690,N_10889,N_11525);
nor U12691 (N_12691,N_11980,N_11567);
nand U12692 (N_12692,N_11820,N_11964);
nor U12693 (N_12693,N_11680,N_10942);
xor U12694 (N_12694,N_11510,N_11702);
or U12695 (N_12695,N_11673,N_10938);
nand U12696 (N_12696,N_11053,N_11179);
and U12697 (N_12697,N_11169,N_11956);
xor U12698 (N_12698,N_11315,N_11106);
or U12699 (N_12699,N_11262,N_11918);
nor U12700 (N_12700,N_11312,N_11014);
or U12701 (N_12701,N_11946,N_11013);
or U12702 (N_12702,N_11190,N_11892);
or U12703 (N_12703,N_11199,N_11715);
or U12704 (N_12704,N_11599,N_11402);
xor U12705 (N_12705,N_11166,N_11518);
nor U12706 (N_12706,N_11005,N_11746);
and U12707 (N_12707,N_11042,N_11184);
or U12708 (N_12708,N_11408,N_11488);
nor U12709 (N_12709,N_11759,N_11199);
nor U12710 (N_12710,N_11949,N_10981);
nor U12711 (N_12711,N_11857,N_11957);
or U12712 (N_12712,N_10888,N_11676);
xnor U12713 (N_12713,N_11960,N_11625);
nor U12714 (N_12714,N_11547,N_11903);
or U12715 (N_12715,N_10889,N_11463);
nand U12716 (N_12716,N_11582,N_11176);
or U12717 (N_12717,N_11812,N_11024);
or U12718 (N_12718,N_11536,N_11055);
nor U12719 (N_12719,N_11201,N_11523);
nor U12720 (N_12720,N_10966,N_11264);
nor U12721 (N_12721,N_11347,N_10801);
xnor U12722 (N_12722,N_11640,N_10845);
nor U12723 (N_12723,N_10818,N_11247);
nor U12724 (N_12724,N_11293,N_11656);
nor U12725 (N_12725,N_11117,N_11717);
nand U12726 (N_12726,N_11883,N_10880);
nand U12727 (N_12727,N_11378,N_10875);
nand U12728 (N_12728,N_11293,N_11428);
xnor U12729 (N_12729,N_11461,N_11864);
and U12730 (N_12730,N_11624,N_11751);
and U12731 (N_12731,N_11059,N_11138);
xor U12732 (N_12732,N_10967,N_11893);
and U12733 (N_12733,N_10931,N_10913);
xor U12734 (N_12734,N_11692,N_11691);
xnor U12735 (N_12735,N_11658,N_11778);
xnor U12736 (N_12736,N_11272,N_11065);
and U12737 (N_12737,N_10907,N_10914);
and U12738 (N_12738,N_11478,N_11552);
xnor U12739 (N_12739,N_11454,N_11823);
xor U12740 (N_12740,N_11857,N_11362);
nor U12741 (N_12741,N_10834,N_10925);
or U12742 (N_12742,N_11944,N_10885);
nand U12743 (N_12743,N_10957,N_11620);
nor U12744 (N_12744,N_11503,N_11497);
nor U12745 (N_12745,N_11371,N_11368);
xor U12746 (N_12746,N_11691,N_10866);
nor U12747 (N_12747,N_11270,N_11959);
xnor U12748 (N_12748,N_11409,N_11607);
nand U12749 (N_12749,N_11506,N_11388);
or U12750 (N_12750,N_10838,N_11176);
nand U12751 (N_12751,N_11865,N_11219);
nand U12752 (N_12752,N_11966,N_10808);
or U12753 (N_12753,N_11245,N_11440);
xor U12754 (N_12754,N_11889,N_11973);
and U12755 (N_12755,N_11594,N_10823);
xor U12756 (N_12756,N_11509,N_11513);
nor U12757 (N_12757,N_11149,N_11054);
nand U12758 (N_12758,N_11454,N_11620);
nor U12759 (N_12759,N_11260,N_11655);
nor U12760 (N_12760,N_11277,N_10883);
or U12761 (N_12761,N_11180,N_11631);
or U12762 (N_12762,N_11497,N_11363);
or U12763 (N_12763,N_11029,N_10889);
nor U12764 (N_12764,N_11911,N_11254);
or U12765 (N_12765,N_10867,N_10949);
and U12766 (N_12766,N_11382,N_11648);
nand U12767 (N_12767,N_11914,N_11318);
nand U12768 (N_12768,N_11295,N_11966);
nor U12769 (N_12769,N_10866,N_11741);
nor U12770 (N_12770,N_11234,N_11283);
nor U12771 (N_12771,N_11572,N_11141);
nor U12772 (N_12772,N_11702,N_11402);
nand U12773 (N_12773,N_11910,N_11401);
and U12774 (N_12774,N_11813,N_11374);
nand U12775 (N_12775,N_11502,N_10879);
or U12776 (N_12776,N_11207,N_11276);
xor U12777 (N_12777,N_11598,N_11449);
nor U12778 (N_12778,N_11264,N_11833);
and U12779 (N_12779,N_11380,N_11063);
xor U12780 (N_12780,N_11704,N_11234);
and U12781 (N_12781,N_10889,N_11867);
and U12782 (N_12782,N_11752,N_11206);
nor U12783 (N_12783,N_11110,N_11351);
nand U12784 (N_12784,N_11575,N_10810);
nand U12785 (N_12785,N_11122,N_11825);
nand U12786 (N_12786,N_11968,N_11867);
nor U12787 (N_12787,N_11310,N_11598);
nor U12788 (N_12788,N_10963,N_11698);
or U12789 (N_12789,N_11669,N_11571);
nor U12790 (N_12790,N_11870,N_11880);
or U12791 (N_12791,N_11745,N_11586);
and U12792 (N_12792,N_11748,N_11168);
nor U12793 (N_12793,N_11192,N_11072);
nor U12794 (N_12794,N_11793,N_11320);
or U12795 (N_12795,N_11601,N_11691);
or U12796 (N_12796,N_11003,N_11778);
nand U12797 (N_12797,N_11162,N_11835);
or U12798 (N_12798,N_11568,N_11183);
nor U12799 (N_12799,N_11063,N_11043);
and U12800 (N_12800,N_11342,N_11826);
nand U12801 (N_12801,N_11159,N_11073);
nor U12802 (N_12802,N_11086,N_10809);
or U12803 (N_12803,N_11471,N_11455);
nor U12804 (N_12804,N_11614,N_11040);
nand U12805 (N_12805,N_11076,N_11086);
and U12806 (N_12806,N_11424,N_11504);
nand U12807 (N_12807,N_10834,N_11213);
xnor U12808 (N_12808,N_11277,N_11241);
nand U12809 (N_12809,N_11141,N_11073);
nand U12810 (N_12810,N_11785,N_11294);
nand U12811 (N_12811,N_11541,N_11492);
xnor U12812 (N_12812,N_11155,N_11582);
xor U12813 (N_12813,N_11009,N_11195);
nor U12814 (N_12814,N_11920,N_10976);
nor U12815 (N_12815,N_10961,N_11620);
nor U12816 (N_12816,N_11218,N_11765);
xor U12817 (N_12817,N_11881,N_11601);
nor U12818 (N_12818,N_11764,N_11178);
and U12819 (N_12819,N_11076,N_11985);
and U12820 (N_12820,N_10891,N_11024);
nor U12821 (N_12821,N_11452,N_11600);
or U12822 (N_12822,N_11594,N_11257);
and U12823 (N_12823,N_11657,N_11547);
nor U12824 (N_12824,N_11806,N_11209);
and U12825 (N_12825,N_11885,N_11443);
xor U12826 (N_12826,N_11296,N_11510);
and U12827 (N_12827,N_11446,N_10913);
and U12828 (N_12828,N_11374,N_11365);
and U12829 (N_12829,N_10977,N_11847);
nand U12830 (N_12830,N_11255,N_11896);
xnor U12831 (N_12831,N_11277,N_10942);
nand U12832 (N_12832,N_11160,N_11327);
nand U12833 (N_12833,N_11958,N_11898);
nor U12834 (N_12834,N_11083,N_10832);
xnor U12835 (N_12835,N_11035,N_11059);
nand U12836 (N_12836,N_11584,N_11989);
nor U12837 (N_12837,N_11395,N_11619);
and U12838 (N_12838,N_11009,N_11882);
xor U12839 (N_12839,N_11741,N_10977);
xnor U12840 (N_12840,N_11816,N_11023);
or U12841 (N_12841,N_11383,N_11404);
or U12842 (N_12842,N_11775,N_11963);
or U12843 (N_12843,N_11676,N_10995);
nand U12844 (N_12844,N_11472,N_11304);
or U12845 (N_12845,N_10868,N_11185);
or U12846 (N_12846,N_11540,N_11194);
xnor U12847 (N_12847,N_11602,N_11263);
or U12848 (N_12848,N_11139,N_11434);
nor U12849 (N_12849,N_11886,N_10816);
nor U12850 (N_12850,N_11381,N_11234);
nand U12851 (N_12851,N_11275,N_11089);
xnor U12852 (N_12852,N_11140,N_10800);
and U12853 (N_12853,N_11330,N_11461);
and U12854 (N_12854,N_11272,N_10814);
or U12855 (N_12855,N_11491,N_11144);
and U12856 (N_12856,N_11482,N_10997);
and U12857 (N_12857,N_11988,N_10843);
nand U12858 (N_12858,N_11148,N_11656);
nand U12859 (N_12859,N_11758,N_10838);
or U12860 (N_12860,N_11805,N_11101);
nor U12861 (N_12861,N_10832,N_11947);
nor U12862 (N_12862,N_11520,N_11116);
nand U12863 (N_12863,N_11749,N_11911);
and U12864 (N_12864,N_11247,N_11642);
nand U12865 (N_12865,N_10806,N_11915);
and U12866 (N_12866,N_11246,N_11368);
xnor U12867 (N_12867,N_10848,N_11398);
nor U12868 (N_12868,N_11541,N_11420);
or U12869 (N_12869,N_11119,N_11141);
and U12870 (N_12870,N_11428,N_10842);
nand U12871 (N_12871,N_10819,N_11854);
nand U12872 (N_12872,N_11702,N_11499);
and U12873 (N_12873,N_11987,N_10918);
nor U12874 (N_12874,N_11406,N_11686);
nand U12875 (N_12875,N_11671,N_11408);
nor U12876 (N_12876,N_11434,N_11744);
or U12877 (N_12877,N_11768,N_11920);
or U12878 (N_12878,N_11774,N_11858);
or U12879 (N_12879,N_11556,N_11513);
nor U12880 (N_12880,N_11292,N_11229);
and U12881 (N_12881,N_11051,N_11876);
nor U12882 (N_12882,N_11643,N_11878);
nand U12883 (N_12883,N_11974,N_11792);
and U12884 (N_12884,N_11064,N_11727);
nand U12885 (N_12885,N_11624,N_11428);
and U12886 (N_12886,N_11983,N_11494);
or U12887 (N_12887,N_11784,N_11418);
nand U12888 (N_12888,N_11673,N_11743);
or U12889 (N_12889,N_11235,N_11805);
xnor U12890 (N_12890,N_11791,N_11015);
xnor U12891 (N_12891,N_11562,N_11065);
or U12892 (N_12892,N_11818,N_11428);
or U12893 (N_12893,N_10883,N_11901);
and U12894 (N_12894,N_10964,N_11142);
xnor U12895 (N_12895,N_11878,N_11213);
or U12896 (N_12896,N_10832,N_10917);
nor U12897 (N_12897,N_11332,N_11222);
nor U12898 (N_12898,N_11211,N_11366);
xor U12899 (N_12899,N_10816,N_11224);
and U12900 (N_12900,N_11781,N_11269);
or U12901 (N_12901,N_11728,N_11171);
nor U12902 (N_12902,N_11652,N_10857);
nand U12903 (N_12903,N_10860,N_11702);
nand U12904 (N_12904,N_11266,N_11919);
xor U12905 (N_12905,N_11239,N_10963);
nand U12906 (N_12906,N_11702,N_11466);
nor U12907 (N_12907,N_10957,N_11477);
nand U12908 (N_12908,N_11058,N_11543);
xor U12909 (N_12909,N_11825,N_11280);
xnor U12910 (N_12910,N_11513,N_11481);
and U12911 (N_12911,N_11379,N_11228);
nand U12912 (N_12912,N_11584,N_11369);
or U12913 (N_12913,N_11286,N_11438);
or U12914 (N_12914,N_11385,N_10839);
xor U12915 (N_12915,N_11148,N_11581);
nand U12916 (N_12916,N_11077,N_11950);
nor U12917 (N_12917,N_10842,N_11042);
or U12918 (N_12918,N_11264,N_11003);
nand U12919 (N_12919,N_11404,N_11029);
or U12920 (N_12920,N_11946,N_11641);
or U12921 (N_12921,N_11784,N_11641);
nand U12922 (N_12922,N_11341,N_11236);
or U12923 (N_12923,N_11187,N_11514);
xor U12924 (N_12924,N_11120,N_11117);
xnor U12925 (N_12925,N_11918,N_11483);
or U12926 (N_12926,N_11774,N_10859);
nor U12927 (N_12927,N_11497,N_10808);
nor U12928 (N_12928,N_10818,N_11767);
xnor U12929 (N_12929,N_11783,N_11003);
and U12930 (N_12930,N_11020,N_11989);
nor U12931 (N_12931,N_11004,N_11470);
xnor U12932 (N_12932,N_11269,N_11227);
nand U12933 (N_12933,N_11720,N_11694);
or U12934 (N_12934,N_11131,N_10957);
nand U12935 (N_12935,N_11412,N_11564);
or U12936 (N_12936,N_11984,N_11004);
or U12937 (N_12937,N_11756,N_10973);
nor U12938 (N_12938,N_11326,N_11926);
nor U12939 (N_12939,N_11559,N_11175);
and U12940 (N_12940,N_11367,N_11713);
nand U12941 (N_12941,N_11924,N_10852);
nand U12942 (N_12942,N_11124,N_11464);
and U12943 (N_12943,N_10895,N_11546);
nand U12944 (N_12944,N_11958,N_11442);
xnor U12945 (N_12945,N_11102,N_11711);
nor U12946 (N_12946,N_10995,N_11832);
and U12947 (N_12947,N_11552,N_11339);
xnor U12948 (N_12948,N_11804,N_10906);
nor U12949 (N_12949,N_11606,N_11979);
or U12950 (N_12950,N_11968,N_11371);
nor U12951 (N_12951,N_11574,N_11882);
nand U12952 (N_12952,N_11897,N_11448);
or U12953 (N_12953,N_11604,N_11301);
xor U12954 (N_12954,N_10836,N_11922);
nor U12955 (N_12955,N_10849,N_10954);
xor U12956 (N_12956,N_11667,N_11828);
xor U12957 (N_12957,N_11978,N_11730);
or U12958 (N_12958,N_11038,N_11300);
or U12959 (N_12959,N_10953,N_11658);
nor U12960 (N_12960,N_11893,N_11555);
nand U12961 (N_12961,N_11448,N_11406);
nand U12962 (N_12962,N_11442,N_11322);
or U12963 (N_12963,N_10854,N_11326);
and U12964 (N_12964,N_11209,N_11295);
nand U12965 (N_12965,N_10865,N_10864);
nand U12966 (N_12966,N_11076,N_11415);
xnor U12967 (N_12967,N_11293,N_11500);
and U12968 (N_12968,N_10992,N_10933);
and U12969 (N_12969,N_11696,N_11885);
nand U12970 (N_12970,N_11545,N_11709);
or U12971 (N_12971,N_11708,N_11335);
or U12972 (N_12972,N_11667,N_11801);
and U12973 (N_12973,N_11368,N_11122);
and U12974 (N_12974,N_10802,N_11994);
and U12975 (N_12975,N_10855,N_11694);
and U12976 (N_12976,N_11435,N_11813);
and U12977 (N_12977,N_10945,N_11526);
nand U12978 (N_12978,N_11046,N_11862);
or U12979 (N_12979,N_11921,N_11297);
xor U12980 (N_12980,N_11335,N_11375);
nor U12981 (N_12981,N_11046,N_11173);
nor U12982 (N_12982,N_10953,N_11400);
and U12983 (N_12983,N_11037,N_11878);
xnor U12984 (N_12984,N_11901,N_11120);
nor U12985 (N_12985,N_11919,N_10950);
xor U12986 (N_12986,N_11096,N_11196);
nand U12987 (N_12987,N_11650,N_11494);
and U12988 (N_12988,N_10938,N_11038);
or U12989 (N_12989,N_11315,N_11921);
nand U12990 (N_12990,N_11529,N_11560);
and U12991 (N_12991,N_11565,N_11200);
nor U12992 (N_12992,N_11867,N_11265);
and U12993 (N_12993,N_11344,N_10947);
nand U12994 (N_12994,N_11599,N_11767);
nor U12995 (N_12995,N_11220,N_11089);
or U12996 (N_12996,N_10837,N_11206);
nor U12997 (N_12997,N_10806,N_11856);
or U12998 (N_12998,N_11572,N_11630);
and U12999 (N_12999,N_11475,N_10983);
nor U13000 (N_13000,N_10919,N_11980);
xor U13001 (N_13001,N_11187,N_11325);
nor U13002 (N_13002,N_11191,N_11044);
nor U13003 (N_13003,N_11140,N_11638);
xnor U13004 (N_13004,N_11745,N_11682);
nor U13005 (N_13005,N_11988,N_11033);
xor U13006 (N_13006,N_11473,N_11300);
or U13007 (N_13007,N_11183,N_11833);
nand U13008 (N_13008,N_10908,N_11786);
nand U13009 (N_13009,N_11099,N_11172);
or U13010 (N_13010,N_11765,N_11131);
nor U13011 (N_13011,N_11463,N_11914);
xor U13012 (N_13012,N_11477,N_11507);
and U13013 (N_13013,N_11128,N_11357);
or U13014 (N_13014,N_11033,N_10835);
nand U13015 (N_13015,N_11048,N_11386);
nand U13016 (N_13016,N_11859,N_11391);
or U13017 (N_13017,N_11582,N_11670);
xor U13018 (N_13018,N_11948,N_10878);
nor U13019 (N_13019,N_11554,N_11495);
xor U13020 (N_13020,N_11204,N_11159);
nor U13021 (N_13021,N_11845,N_11313);
nand U13022 (N_13022,N_11310,N_11822);
or U13023 (N_13023,N_11256,N_11257);
nor U13024 (N_13024,N_11221,N_10931);
xnor U13025 (N_13025,N_11500,N_11925);
or U13026 (N_13026,N_10817,N_11448);
and U13027 (N_13027,N_11531,N_11720);
nor U13028 (N_13028,N_11441,N_11844);
or U13029 (N_13029,N_11258,N_11052);
and U13030 (N_13030,N_11559,N_11572);
nand U13031 (N_13031,N_11106,N_11314);
xor U13032 (N_13032,N_11068,N_11630);
nand U13033 (N_13033,N_11531,N_11439);
nor U13034 (N_13034,N_11676,N_11814);
and U13035 (N_13035,N_11834,N_11401);
xor U13036 (N_13036,N_11670,N_11609);
xnor U13037 (N_13037,N_11312,N_11990);
nor U13038 (N_13038,N_11216,N_10808);
or U13039 (N_13039,N_11580,N_10968);
and U13040 (N_13040,N_11208,N_11670);
or U13041 (N_13041,N_11745,N_11282);
or U13042 (N_13042,N_11679,N_10965);
or U13043 (N_13043,N_10952,N_10911);
and U13044 (N_13044,N_11969,N_11125);
or U13045 (N_13045,N_11576,N_11530);
and U13046 (N_13046,N_11535,N_11229);
xor U13047 (N_13047,N_11831,N_11584);
nand U13048 (N_13048,N_11034,N_11173);
and U13049 (N_13049,N_11143,N_10936);
nand U13050 (N_13050,N_11868,N_10964);
and U13051 (N_13051,N_11812,N_11650);
xnor U13052 (N_13052,N_11883,N_11804);
nor U13053 (N_13053,N_11563,N_11361);
nand U13054 (N_13054,N_11621,N_10830);
xor U13055 (N_13055,N_10959,N_11506);
and U13056 (N_13056,N_10928,N_11059);
xnor U13057 (N_13057,N_11872,N_11403);
xor U13058 (N_13058,N_11360,N_11392);
nand U13059 (N_13059,N_11155,N_10865);
nor U13060 (N_13060,N_11325,N_11808);
nand U13061 (N_13061,N_11729,N_10854);
nand U13062 (N_13062,N_11120,N_11469);
nand U13063 (N_13063,N_11571,N_11135);
and U13064 (N_13064,N_10802,N_11912);
or U13065 (N_13065,N_11472,N_11785);
xor U13066 (N_13066,N_11574,N_11291);
xnor U13067 (N_13067,N_11945,N_11066);
or U13068 (N_13068,N_10884,N_11042);
or U13069 (N_13069,N_11147,N_11009);
or U13070 (N_13070,N_11214,N_11349);
or U13071 (N_13071,N_10945,N_11612);
xnor U13072 (N_13072,N_11494,N_11091);
and U13073 (N_13073,N_11125,N_11407);
and U13074 (N_13074,N_11734,N_10970);
xnor U13075 (N_13075,N_11265,N_11497);
nor U13076 (N_13076,N_11093,N_11123);
nand U13077 (N_13077,N_11186,N_11344);
or U13078 (N_13078,N_11246,N_10987);
nand U13079 (N_13079,N_11169,N_11740);
or U13080 (N_13080,N_11991,N_11510);
nor U13081 (N_13081,N_11533,N_11337);
and U13082 (N_13082,N_11178,N_11959);
nand U13083 (N_13083,N_10937,N_10992);
and U13084 (N_13084,N_11830,N_11273);
and U13085 (N_13085,N_11331,N_10840);
xnor U13086 (N_13086,N_10840,N_11179);
nand U13087 (N_13087,N_10953,N_11739);
or U13088 (N_13088,N_11339,N_11420);
or U13089 (N_13089,N_11558,N_11071);
nor U13090 (N_13090,N_11699,N_10858);
xnor U13091 (N_13091,N_11851,N_11689);
or U13092 (N_13092,N_11405,N_10996);
or U13093 (N_13093,N_11939,N_11193);
nand U13094 (N_13094,N_10854,N_11247);
and U13095 (N_13095,N_11161,N_11111);
nor U13096 (N_13096,N_11745,N_11725);
xnor U13097 (N_13097,N_11474,N_11338);
xnor U13098 (N_13098,N_11091,N_11507);
or U13099 (N_13099,N_11166,N_11787);
nor U13100 (N_13100,N_11845,N_11780);
or U13101 (N_13101,N_11910,N_11662);
nor U13102 (N_13102,N_11103,N_11753);
xnor U13103 (N_13103,N_11238,N_11550);
and U13104 (N_13104,N_11841,N_11192);
or U13105 (N_13105,N_11557,N_11402);
and U13106 (N_13106,N_10829,N_11756);
nand U13107 (N_13107,N_10954,N_11365);
or U13108 (N_13108,N_11290,N_11682);
nand U13109 (N_13109,N_11507,N_11197);
nand U13110 (N_13110,N_11881,N_10967);
xor U13111 (N_13111,N_11289,N_11116);
and U13112 (N_13112,N_11706,N_11786);
nor U13113 (N_13113,N_11137,N_11385);
nand U13114 (N_13114,N_11829,N_11441);
nor U13115 (N_13115,N_11723,N_11763);
and U13116 (N_13116,N_11242,N_11915);
and U13117 (N_13117,N_11274,N_11915);
nand U13118 (N_13118,N_11996,N_10936);
xnor U13119 (N_13119,N_10932,N_11361);
or U13120 (N_13120,N_10882,N_11947);
nor U13121 (N_13121,N_11488,N_11339);
nand U13122 (N_13122,N_11386,N_11257);
xor U13123 (N_13123,N_11628,N_11474);
or U13124 (N_13124,N_10841,N_11593);
and U13125 (N_13125,N_11329,N_11008);
or U13126 (N_13126,N_11620,N_10808);
nand U13127 (N_13127,N_11582,N_11551);
and U13128 (N_13128,N_11823,N_11047);
or U13129 (N_13129,N_11218,N_11322);
nand U13130 (N_13130,N_11712,N_10830);
or U13131 (N_13131,N_11329,N_11217);
xnor U13132 (N_13132,N_11986,N_11754);
and U13133 (N_13133,N_10912,N_11009);
and U13134 (N_13134,N_11145,N_11382);
nand U13135 (N_13135,N_11215,N_11634);
and U13136 (N_13136,N_11108,N_11621);
and U13137 (N_13137,N_11032,N_11456);
and U13138 (N_13138,N_11710,N_11035);
nor U13139 (N_13139,N_11504,N_11550);
nand U13140 (N_13140,N_11407,N_11413);
nor U13141 (N_13141,N_11898,N_11150);
or U13142 (N_13142,N_11527,N_11973);
and U13143 (N_13143,N_11078,N_11545);
nand U13144 (N_13144,N_10901,N_11021);
and U13145 (N_13145,N_11572,N_11040);
nor U13146 (N_13146,N_10977,N_11931);
or U13147 (N_13147,N_11906,N_11532);
nor U13148 (N_13148,N_10873,N_11076);
or U13149 (N_13149,N_10808,N_11054);
nand U13150 (N_13150,N_11706,N_10814);
nor U13151 (N_13151,N_11469,N_11906);
and U13152 (N_13152,N_10862,N_11332);
and U13153 (N_13153,N_11944,N_11216);
xnor U13154 (N_13154,N_11689,N_10873);
nor U13155 (N_13155,N_11487,N_11524);
or U13156 (N_13156,N_11764,N_10924);
and U13157 (N_13157,N_11993,N_10871);
xnor U13158 (N_13158,N_11286,N_11079);
nand U13159 (N_13159,N_10905,N_11371);
xnor U13160 (N_13160,N_11130,N_11992);
nand U13161 (N_13161,N_11276,N_11250);
nand U13162 (N_13162,N_11392,N_11960);
nand U13163 (N_13163,N_10991,N_11333);
nand U13164 (N_13164,N_11589,N_11437);
nand U13165 (N_13165,N_11006,N_11382);
nand U13166 (N_13166,N_11431,N_10862);
xnor U13167 (N_13167,N_11713,N_11343);
xnor U13168 (N_13168,N_11704,N_10892);
and U13169 (N_13169,N_11288,N_11005);
nand U13170 (N_13170,N_11297,N_11333);
xor U13171 (N_13171,N_11052,N_11766);
nand U13172 (N_13172,N_11014,N_11812);
and U13173 (N_13173,N_11559,N_11943);
xor U13174 (N_13174,N_11529,N_11717);
and U13175 (N_13175,N_11657,N_11646);
or U13176 (N_13176,N_11798,N_11156);
xor U13177 (N_13177,N_11292,N_11211);
and U13178 (N_13178,N_11325,N_11083);
nand U13179 (N_13179,N_11992,N_11455);
or U13180 (N_13180,N_11845,N_11708);
and U13181 (N_13181,N_11623,N_10883);
nor U13182 (N_13182,N_11422,N_11419);
or U13183 (N_13183,N_10822,N_11308);
xnor U13184 (N_13184,N_10866,N_11375);
nand U13185 (N_13185,N_11877,N_11430);
xor U13186 (N_13186,N_11317,N_10921);
nand U13187 (N_13187,N_10969,N_10880);
xor U13188 (N_13188,N_11793,N_11254);
nand U13189 (N_13189,N_11199,N_11672);
xnor U13190 (N_13190,N_11792,N_11826);
xnor U13191 (N_13191,N_11512,N_11861);
xnor U13192 (N_13192,N_11574,N_11794);
and U13193 (N_13193,N_11741,N_11574);
or U13194 (N_13194,N_11154,N_11419);
or U13195 (N_13195,N_11951,N_11971);
xor U13196 (N_13196,N_11536,N_11298);
and U13197 (N_13197,N_11949,N_11958);
and U13198 (N_13198,N_11775,N_10838);
or U13199 (N_13199,N_11248,N_11333);
or U13200 (N_13200,N_12962,N_12468);
or U13201 (N_13201,N_13170,N_12982);
nand U13202 (N_13202,N_13111,N_12067);
xnor U13203 (N_13203,N_12193,N_12224);
xor U13204 (N_13204,N_12876,N_12145);
and U13205 (N_13205,N_13089,N_12394);
and U13206 (N_13206,N_12754,N_12586);
nand U13207 (N_13207,N_12363,N_12778);
nor U13208 (N_13208,N_12292,N_12133);
and U13209 (N_13209,N_12179,N_12889);
xnor U13210 (N_13210,N_12895,N_13073);
nand U13211 (N_13211,N_12213,N_13077);
or U13212 (N_13212,N_12742,N_12178);
nand U13213 (N_13213,N_13080,N_12555);
xnor U13214 (N_13214,N_12558,N_12910);
nand U13215 (N_13215,N_12485,N_13085);
xnor U13216 (N_13216,N_12746,N_12384);
nor U13217 (N_13217,N_12286,N_12704);
or U13218 (N_13218,N_12376,N_13125);
and U13219 (N_13219,N_12294,N_13024);
and U13220 (N_13220,N_12620,N_13019);
nand U13221 (N_13221,N_13044,N_12272);
nand U13222 (N_13222,N_12152,N_12391);
or U13223 (N_13223,N_12758,N_12393);
nand U13224 (N_13224,N_12734,N_12119);
or U13225 (N_13225,N_12091,N_12388);
and U13226 (N_13226,N_12601,N_12209);
or U13227 (N_13227,N_13193,N_12281);
and U13228 (N_13228,N_12873,N_13128);
nand U13229 (N_13229,N_13109,N_12549);
nor U13230 (N_13230,N_12414,N_13122);
nand U13231 (N_13231,N_12317,N_12865);
xor U13232 (N_13232,N_12680,N_12148);
xnor U13233 (N_13233,N_12052,N_12408);
xnor U13234 (N_13234,N_12733,N_12086);
and U13235 (N_13235,N_12990,N_13078);
nand U13236 (N_13236,N_12029,N_12154);
and U13237 (N_13237,N_13000,N_12832);
nand U13238 (N_13238,N_12600,N_12320);
xnor U13239 (N_13239,N_12277,N_13174);
or U13240 (N_13240,N_13033,N_13067);
or U13241 (N_13241,N_12419,N_12382);
xor U13242 (N_13242,N_12437,N_12532);
nand U13243 (N_13243,N_12476,N_12167);
xnor U13244 (N_13244,N_12821,N_12663);
and U13245 (N_13245,N_12624,N_12313);
and U13246 (N_13246,N_12137,N_12748);
and U13247 (N_13247,N_12981,N_12235);
nor U13248 (N_13248,N_12329,N_12176);
or U13249 (N_13249,N_13003,N_13163);
xnor U13250 (N_13250,N_12379,N_12037);
or U13251 (N_13251,N_12736,N_12813);
xor U13252 (N_13252,N_12852,N_13062);
nand U13253 (N_13253,N_13123,N_12797);
xnor U13254 (N_13254,N_12378,N_12039);
nand U13255 (N_13255,N_13135,N_12205);
nand U13256 (N_13256,N_12270,N_12578);
nor U13257 (N_13257,N_13127,N_12349);
xnor U13258 (N_13258,N_12573,N_12793);
xnor U13259 (N_13259,N_12315,N_12418);
xnor U13260 (N_13260,N_12773,N_12653);
and U13261 (N_13261,N_13095,N_12513);
or U13262 (N_13262,N_13016,N_12407);
xor U13263 (N_13263,N_13188,N_12735);
nor U13264 (N_13264,N_12498,N_12073);
xnor U13265 (N_13265,N_12948,N_12059);
nand U13266 (N_13266,N_12569,N_12759);
xor U13267 (N_13267,N_12714,N_13194);
nor U13268 (N_13268,N_12931,N_13094);
nand U13269 (N_13269,N_12946,N_12168);
and U13270 (N_13270,N_12968,N_12766);
nor U13271 (N_13271,N_12085,N_13146);
or U13272 (N_13272,N_12061,N_12880);
and U13273 (N_13273,N_12642,N_12135);
xor U13274 (N_13274,N_12301,N_12731);
and U13275 (N_13275,N_12449,N_12475);
and U13276 (N_13276,N_12482,N_12446);
and U13277 (N_13277,N_12093,N_12678);
nand U13278 (N_13278,N_12927,N_12131);
nand U13279 (N_13279,N_12868,N_13001);
or U13280 (N_13280,N_12023,N_12361);
nor U13281 (N_13281,N_12357,N_12201);
and U13282 (N_13282,N_12441,N_13172);
nor U13283 (N_13283,N_12013,N_12132);
xnor U13284 (N_13284,N_12582,N_12283);
nor U13285 (N_13285,N_12256,N_12830);
nor U13286 (N_13286,N_12715,N_12303);
nor U13287 (N_13287,N_12563,N_12929);
or U13288 (N_13288,N_12196,N_12583);
or U13289 (N_13289,N_12025,N_12877);
and U13290 (N_13290,N_13008,N_12151);
and U13291 (N_13291,N_13051,N_12916);
and U13292 (N_13292,N_12275,N_12011);
or U13293 (N_13293,N_12447,N_13047);
nor U13294 (N_13294,N_12829,N_12375);
nand U13295 (N_13295,N_12352,N_12814);
or U13296 (N_13296,N_13040,N_12238);
or U13297 (N_13297,N_12108,N_12187);
xnor U13298 (N_13298,N_12616,N_12707);
nand U13299 (N_13299,N_12040,N_12888);
nor U13300 (N_13300,N_12463,N_13184);
xnor U13301 (N_13301,N_12918,N_13186);
nor U13302 (N_13302,N_12323,N_12136);
or U13303 (N_13303,N_13107,N_13190);
or U13304 (N_13304,N_12791,N_12355);
nor U13305 (N_13305,N_12531,N_12621);
xor U13306 (N_13306,N_12522,N_12480);
or U13307 (N_13307,N_12041,N_12543);
nor U13308 (N_13308,N_12316,N_13011);
or U13309 (N_13309,N_13156,N_12157);
xnor U13310 (N_13310,N_12412,N_12785);
and U13311 (N_13311,N_12683,N_12649);
xor U13312 (N_13312,N_12423,N_12699);
nor U13313 (N_13313,N_12626,N_12138);
xnor U13314 (N_13314,N_13074,N_12765);
and U13315 (N_13315,N_12156,N_12777);
nand U13316 (N_13316,N_12637,N_12116);
nand U13317 (N_13317,N_12677,N_12420);
xnor U13318 (N_13318,N_12994,N_12459);
nor U13319 (N_13319,N_12980,N_12882);
nand U13320 (N_13320,N_12208,N_12950);
and U13321 (N_13321,N_12872,N_12076);
xor U13322 (N_13322,N_12967,N_12163);
nor U13323 (N_13323,N_12805,N_13117);
xnor U13324 (N_13324,N_13010,N_12327);
nor U13325 (N_13325,N_12692,N_12454);
xnor U13326 (N_13326,N_12634,N_12853);
nand U13327 (N_13327,N_12756,N_12698);
and U13328 (N_13328,N_12338,N_12198);
nand U13329 (N_13329,N_12744,N_12280);
nand U13330 (N_13330,N_12346,N_12779);
nand U13331 (N_13331,N_12460,N_12727);
xor U13332 (N_13332,N_12986,N_12243);
nor U13333 (N_13333,N_12373,N_12644);
nor U13334 (N_13334,N_12126,N_12033);
nor U13335 (N_13335,N_12892,N_12548);
and U13336 (N_13336,N_12599,N_12691);
and U13337 (N_13337,N_12870,N_12703);
xor U13338 (N_13338,N_12668,N_12380);
nor U13339 (N_13339,N_12854,N_12836);
xor U13340 (N_13340,N_12804,N_12142);
xnor U13341 (N_13341,N_12488,N_12232);
xnor U13342 (N_13342,N_12858,N_12058);
and U13343 (N_13343,N_12730,N_12713);
xor U13344 (N_13344,N_12075,N_12180);
xor U13345 (N_13345,N_12539,N_12887);
or U13346 (N_13346,N_13139,N_12786);
xnor U13347 (N_13347,N_12263,N_12080);
nor U13348 (N_13348,N_12121,N_13118);
and U13349 (N_13349,N_12939,N_12367);
nor U13350 (N_13350,N_13090,N_13081);
nor U13351 (N_13351,N_12847,N_12690);
or U13352 (N_13352,N_12435,N_12619);
and U13353 (N_13353,N_12045,N_13178);
nand U13354 (N_13354,N_12110,N_12987);
nor U13355 (N_13355,N_12099,N_12300);
nand U13356 (N_13356,N_12056,N_12122);
and U13357 (N_13357,N_12359,N_13088);
or U13358 (N_13358,N_12672,N_12752);
xnor U13359 (N_13359,N_12491,N_12124);
nor U13360 (N_13360,N_12751,N_12789);
xnor U13361 (N_13361,N_12996,N_12696);
nor U13362 (N_13362,N_12974,N_12207);
and U13363 (N_13363,N_12452,N_12705);
nor U13364 (N_13364,N_12060,N_12762);
xnor U13365 (N_13365,N_12335,N_12815);
or U13366 (N_13366,N_12949,N_12031);
nor U13367 (N_13367,N_12693,N_13169);
xnor U13368 (N_13368,N_12016,N_12845);
nand U13369 (N_13369,N_12422,N_12371);
nor U13370 (N_13370,N_12258,N_12340);
and U13371 (N_13371,N_12020,N_12726);
nand U13372 (N_13372,N_12771,N_12034);
nand U13373 (N_13373,N_12190,N_13141);
or U13374 (N_13374,N_12528,N_12926);
or U13375 (N_13375,N_13105,N_13110);
or U13376 (N_13376,N_13161,N_12776);
nor U13377 (N_13377,N_12947,N_12319);
nor U13378 (N_13378,N_12965,N_12386);
xor U13379 (N_13379,N_12251,N_12161);
or U13380 (N_13380,N_12643,N_12661);
and U13381 (N_13381,N_12557,N_12392);
nor U13382 (N_13382,N_12141,N_12943);
nor U13383 (N_13383,N_12622,N_13093);
xnor U13384 (N_13384,N_12239,N_12679);
and U13385 (N_13385,N_12720,N_13198);
or U13386 (N_13386,N_13012,N_12800);
nor U13387 (N_13387,N_12433,N_12267);
or U13388 (N_13388,N_12749,N_13175);
or U13389 (N_13389,N_12848,N_12509);
nand U13390 (N_13390,N_12591,N_12757);
nand U13391 (N_13391,N_12567,N_12240);
or U13392 (N_13392,N_12527,N_12385);
nand U13393 (N_13393,N_12851,N_12417);
nor U13394 (N_13394,N_12884,N_12761);
or U13395 (N_13395,N_13070,N_12606);
nor U13396 (N_13396,N_12684,N_12183);
and U13397 (N_13397,N_12553,N_12768);
xor U13398 (N_13398,N_12117,N_12487);
nor U13399 (N_13399,N_12216,N_12299);
nand U13400 (N_13400,N_12724,N_12869);
xnor U13401 (N_13401,N_12186,N_12722);
nand U13402 (N_13402,N_13082,N_12885);
nor U13403 (N_13403,N_12900,N_13021);
xor U13404 (N_13404,N_12217,N_12100);
and U13405 (N_13405,N_13179,N_12347);
or U13406 (N_13406,N_12005,N_13049);
nand U13407 (N_13407,N_12398,N_12369);
or U13408 (N_13408,N_12304,N_12508);
nand U13409 (N_13409,N_13042,N_12901);
and U13410 (N_13410,N_12928,N_12958);
and U13411 (N_13411,N_12657,N_12496);
and U13412 (N_13412,N_12101,N_12656);
or U13413 (N_13413,N_12220,N_12257);
and U13414 (N_13414,N_12844,N_13195);
or U13415 (N_13415,N_13187,N_12955);
or U13416 (N_13416,N_13140,N_12662);
and U13417 (N_13417,N_12397,N_12185);
nor U13418 (N_13418,N_12125,N_12597);
and U13419 (N_13419,N_13086,N_12002);
nor U13420 (N_13420,N_12760,N_13191);
and U13421 (N_13421,N_13035,N_13029);
and U13422 (N_13422,N_12500,N_12353);
and U13423 (N_13423,N_12495,N_12617);
xnor U13424 (N_13424,N_12465,N_13171);
nor U13425 (N_13425,N_12451,N_12194);
nor U13426 (N_13426,N_12381,N_12835);
or U13427 (N_13427,N_12360,N_12350);
nand U13428 (N_13428,N_12064,N_13166);
and U13429 (N_13429,N_12175,N_12218);
nand U13430 (N_13430,N_12801,N_12159);
xnor U13431 (N_13431,N_12556,N_12741);
nand U13432 (N_13432,N_12787,N_13134);
nor U13433 (N_13433,N_13143,N_12206);
or U13434 (N_13434,N_12229,N_12000);
and U13435 (N_13435,N_12524,N_12436);
and U13436 (N_13436,N_12992,N_12112);
or U13437 (N_13437,N_12262,N_12022);
xor U13438 (N_13438,N_13046,N_12134);
and U13439 (N_13439,N_12561,N_12658);
nand U13440 (N_13440,N_12402,N_12051);
and U13441 (N_13441,N_12828,N_12111);
nand U13442 (N_13442,N_12211,N_12226);
or U13443 (N_13443,N_12523,N_12989);
and U13444 (N_13444,N_13018,N_12769);
and U13445 (N_13445,N_12004,N_12344);
nor U13446 (N_13446,N_13177,N_12214);
and U13447 (N_13447,N_13069,N_12809);
and U13448 (N_13448,N_12747,N_12694);
or U13449 (N_13449,N_12172,N_12538);
nand U13450 (N_13450,N_12298,N_12442);
or U13451 (N_13451,N_13145,N_12611);
and U13452 (N_13452,N_13102,N_12332);
nor U13453 (N_13453,N_12063,N_13059);
and U13454 (N_13454,N_12307,N_13197);
nand U13455 (N_13455,N_12489,N_12646);
nand U13456 (N_13456,N_12254,N_12590);
or U13457 (N_13457,N_12952,N_13071);
nor U13458 (N_13458,N_12484,N_12246);
and U13459 (N_13459,N_12984,N_12841);
nand U13460 (N_13460,N_12291,N_12577);
nor U13461 (N_13461,N_13189,N_12906);
or U13462 (N_13462,N_12651,N_12035);
nor U13463 (N_13463,N_12675,N_12973);
and U13464 (N_13464,N_12954,N_12351);
nand U13465 (N_13465,N_12914,N_12983);
and U13466 (N_13466,N_12648,N_12972);
or U13467 (N_13467,N_12631,N_12941);
nand U13468 (N_13468,N_12118,N_12505);
nor U13469 (N_13469,N_12700,N_12147);
or U13470 (N_13470,N_13013,N_12874);
nor U13471 (N_13471,N_12784,N_12937);
or U13472 (N_13472,N_12047,N_12507);
xor U13473 (N_13473,N_12166,N_13176);
and U13474 (N_13474,N_12993,N_12146);
or U13475 (N_13475,N_12922,N_12288);
or U13476 (N_13476,N_12718,N_12660);
and U13477 (N_13477,N_12105,N_12077);
nand U13478 (N_13478,N_13014,N_12667);
nor U13479 (N_13479,N_12079,N_12158);
xor U13480 (N_13480,N_12788,N_12623);
or U13481 (N_13481,N_12795,N_12820);
and U13482 (N_13482,N_12354,N_12015);
xnor U13483 (N_13483,N_12195,N_12825);
and U13484 (N_13484,N_12883,N_12470);
xnor U13485 (N_13485,N_12160,N_12979);
or U13486 (N_13486,N_12740,N_12840);
nand U13487 (N_13487,N_12875,N_12399);
or U13488 (N_13488,N_12861,N_12439);
nor U13489 (N_13489,N_12405,N_12794);
or U13490 (N_13490,N_12745,N_12130);
nand U13491 (N_13491,N_12222,N_13101);
xor U13492 (N_13492,N_12839,N_12753);
and U13493 (N_13493,N_12721,N_13114);
nor U13494 (N_13494,N_13154,N_12309);
nand U13495 (N_13495,N_12846,N_13048);
nor U13496 (N_13496,N_12324,N_12409);
xor U13497 (N_13497,N_12372,N_12526);
or U13498 (N_13498,N_12472,N_12919);
nand U13499 (N_13499,N_12200,N_12615);
xnor U13500 (N_13500,N_13061,N_12387);
nor U13501 (N_13501,N_13155,N_12995);
and U13502 (N_13502,N_12737,N_12636);
or U13503 (N_13503,N_12911,N_13096);
and U13504 (N_13504,N_12072,N_12976);
nand U13505 (N_13505,N_12518,N_12236);
or U13506 (N_13506,N_12650,N_12799);
or U13507 (N_13507,N_12671,N_13153);
or U13508 (N_13508,N_12571,N_12424);
nor U13509 (N_13509,N_13037,N_12331);
nand U13510 (N_13510,N_13142,N_12455);
and U13511 (N_13511,N_12010,N_12803);
and U13512 (N_13512,N_13181,N_13043);
and U13513 (N_13513,N_12530,N_13130);
xnor U13514 (N_13514,N_13038,N_12891);
nand U13515 (N_13515,N_12991,N_12711);
xor U13516 (N_13516,N_12203,N_12434);
or U13517 (N_13517,N_12501,N_12271);
xor U13518 (N_13518,N_13005,N_12878);
nand U13519 (N_13519,N_13100,N_13152);
and U13520 (N_13520,N_13065,N_12341);
xnor U13521 (N_13521,N_13157,N_12796);
nor U13522 (N_13522,N_12961,N_12629);
xnor U13523 (N_13523,N_12311,N_12572);
nor U13524 (N_13524,N_12782,N_12602);
nand U13525 (N_13525,N_12276,N_12170);
nand U13526 (N_13526,N_12425,N_13165);
nand U13527 (N_13527,N_12542,N_12570);
xnor U13528 (N_13528,N_12348,N_12006);
nor U13529 (N_13529,N_12462,N_13092);
nor U13530 (N_13530,N_12610,N_13026);
nor U13531 (N_13531,N_12400,N_12242);
xnor U13532 (N_13532,N_12227,N_13052);
and U13533 (N_13533,N_13004,N_12411);
or U13534 (N_13534,N_12001,N_12595);
xnor U13535 (N_13535,N_12358,N_12934);
nor U13536 (N_13536,N_12550,N_12009);
nand U13537 (N_13537,N_12702,N_13034);
nor U13538 (N_13538,N_12413,N_12585);
or U13539 (N_13539,N_13091,N_12816);
nand U13540 (N_13540,N_12915,N_12826);
nand U13541 (N_13541,N_12325,N_12956);
nand U13542 (N_13542,N_12255,N_12781);
nor U13543 (N_13543,N_12849,N_12598);
or U13544 (N_13544,N_12429,N_12871);
nor U13545 (N_13545,N_13199,N_12043);
xor U13546 (N_13546,N_12410,N_12655);
or U13547 (N_13547,N_12625,N_12647);
and U13548 (N_13548,N_13066,N_12997);
or U13549 (N_13549,N_12129,N_12028);
and U13550 (N_13550,N_12665,N_13133);
nor U13551 (N_13551,N_13124,N_12917);
nand U13552 (N_13552,N_12248,N_12428);
and U13553 (N_13553,N_12945,N_12977);
or U13554 (N_13554,N_12297,N_12312);
or U13555 (N_13555,N_12305,N_12739);
and U13556 (N_13556,N_12516,N_12609);
xnor U13557 (N_13557,N_12823,N_13020);
xnor U13558 (N_13558,N_12894,N_12512);
nor U13559 (N_13559,N_13054,N_12287);
nor U13560 (N_13560,N_12908,N_12342);
and U13561 (N_13561,N_12716,N_12030);
or U13562 (N_13562,N_12109,N_12310);
xnor U13563 (N_13563,N_12219,N_12850);
nand U13564 (N_13564,N_12525,N_12710);
nand U13565 (N_13565,N_12529,N_12453);
nor U13566 (N_13566,N_12971,N_12438);
nor U13567 (N_13567,N_12898,N_12065);
or U13568 (N_13568,N_12202,N_12461);
nand U13569 (N_13569,N_12688,N_13138);
xnor U13570 (N_13570,N_12071,N_12807);
xnor U13571 (N_13571,N_12842,N_12775);
and U13572 (N_13572,N_12942,N_12204);
and U13573 (N_13573,N_12810,N_12604);
xnor U13574 (N_13574,N_12265,N_12709);
nand U13575 (N_13575,N_12467,N_13076);
and U13576 (N_13576,N_12389,N_13017);
and U13577 (N_13577,N_12920,N_12456);
and U13578 (N_13578,N_12416,N_12492);
nor U13579 (N_13579,N_12899,N_12806);
and U13580 (N_13580,N_13055,N_12123);
or U13581 (N_13581,N_12564,N_12450);
nand U13582 (N_13582,N_12554,N_13173);
nand U13583 (N_13583,N_12120,N_12223);
or U13584 (N_13584,N_12964,N_12448);
and U13585 (N_13585,N_12081,N_12103);
nand U13586 (N_13586,N_12293,N_12431);
and U13587 (N_13587,N_12537,N_13075);
nand U13588 (N_13588,N_12473,N_12466);
or U13589 (N_13589,N_12048,N_12261);
nand U13590 (N_13590,N_12681,N_13182);
nor U13591 (N_13591,N_12290,N_12812);
nand U13592 (N_13592,N_12562,N_13072);
nor U13593 (N_13593,N_12231,N_12362);
and U13594 (N_13594,N_13168,N_12088);
and U13595 (N_13595,N_12932,N_12188);
and U13596 (N_13596,N_12139,N_12032);
nand U13597 (N_13597,N_12144,N_12174);
nand U13598 (N_13598,N_13180,N_13056);
nor U13599 (N_13599,N_12959,N_13112);
and U13600 (N_13600,N_12933,N_12689);
xnor U13601 (N_13601,N_12007,N_13132);
nand U13602 (N_13602,N_12614,N_12269);
nor U13603 (N_13603,N_12477,N_13137);
and U13604 (N_13604,N_12930,N_13030);
or U13605 (N_13605,N_12695,N_12886);
and U13606 (N_13606,N_13126,N_13032);
xor U13607 (N_13607,N_12966,N_13084);
or U13608 (N_13608,N_12855,N_12102);
and U13609 (N_13609,N_12066,N_12864);
xor U13610 (N_13610,N_13045,N_12483);
nor U13611 (N_13611,N_12421,N_12924);
xnor U13612 (N_13612,N_12594,N_12115);
nor U13613 (N_13613,N_12587,N_13098);
nor U13614 (N_13614,N_12486,N_12780);
or U13615 (N_13615,N_12012,N_12579);
and U13616 (N_13616,N_12514,N_12545);
nand U13617 (N_13617,N_12822,N_12560);
and U13618 (N_13618,N_13183,N_12923);
or U13619 (N_13619,N_12343,N_12515);
or U13620 (N_13620,N_12764,N_12503);
nor U13621 (N_13621,N_13068,N_12936);
and U13622 (N_13622,N_12774,N_12199);
nand U13623 (N_13623,N_12763,N_12957);
nand U13624 (N_13624,N_12426,N_12540);
nor U13625 (N_13625,N_12314,N_12469);
nand U13626 (N_13626,N_12738,N_12302);
nor U13627 (N_13627,N_12798,N_12057);
nor U13628 (N_13628,N_12259,N_12905);
or U13629 (N_13629,N_12627,N_12169);
or U13630 (N_13630,N_13025,N_12478);
or U13631 (N_13631,N_12228,N_12859);
nor U13632 (N_13632,N_13159,N_13023);
nand U13633 (N_13633,N_12499,N_12592);
and U13634 (N_13634,N_12274,N_12940);
nor U13635 (N_13635,N_12306,N_12330);
nand U13636 (N_13636,N_12403,N_12879);
nor U13637 (N_13637,N_12988,N_12443);
nor U13638 (N_13638,N_12322,N_12042);
and U13639 (N_13639,N_12106,N_12212);
nand U13640 (N_13640,N_12638,N_13057);
or U13641 (N_13641,N_13041,N_12328);
xor U13642 (N_13642,N_12440,N_12652);
nor U13643 (N_13643,N_13060,N_13136);
or U13644 (N_13644,N_12003,N_12069);
xor U13645 (N_13645,N_12377,N_12641);
or U13646 (N_13646,N_12589,N_13147);
nand U13647 (N_13647,N_12345,N_13131);
or U13648 (N_13648,N_13002,N_12862);
nor U13649 (N_13649,N_12171,N_13115);
xor U13650 (N_13650,N_12321,N_12921);
nor U13651 (N_13651,N_12107,N_12092);
and U13652 (N_13652,N_12802,N_12368);
nand U13653 (N_13653,N_12427,N_12728);
nor U13654 (N_13654,N_12365,N_12502);
or U13655 (N_13655,N_13106,N_13064);
and U13656 (N_13656,N_12944,N_12279);
and U13657 (N_13657,N_12951,N_12580);
and U13658 (N_13658,N_12143,N_13006);
xor U13659 (N_13659,N_12860,N_12581);
or U13660 (N_13660,N_13050,N_12252);
nand U13661 (N_13661,N_12613,N_12070);
nor U13662 (N_13662,N_12506,N_12520);
xor U13663 (N_13663,N_13151,N_12113);
nor U13664 (N_13664,N_12493,N_12676);
xnor U13665 (N_13665,N_12444,N_12266);
and U13666 (N_13666,N_12863,N_12019);
nor U13667 (N_13667,N_12364,N_13083);
nor U13668 (N_13668,N_12881,N_12925);
and U13669 (N_13669,N_12114,N_12104);
xnor U13670 (N_13670,N_12673,N_12588);
and U13671 (N_13671,N_12162,N_12666);
and U13672 (N_13672,N_13063,N_12605);
nand U13673 (N_13673,N_12999,N_12985);
nand U13674 (N_13674,N_12576,N_12790);
or U13675 (N_13675,N_12127,N_12767);
or U13676 (N_13676,N_12837,N_12632);
or U13677 (N_13677,N_12907,N_12755);
nand U13678 (N_13678,N_12253,N_12318);
nor U13679 (N_13679,N_12723,N_12356);
xnor U13680 (N_13680,N_12819,N_12497);
xor U13681 (N_13681,N_12233,N_13022);
nand U13682 (N_13682,N_12049,N_12128);
or U13683 (N_13683,N_12308,N_12062);
or U13684 (N_13684,N_12708,N_12670);
or U13685 (N_13685,N_13120,N_12458);
xnor U13686 (N_13686,N_12511,N_12396);
or U13687 (N_13687,N_12953,N_12181);
and U13688 (N_13688,N_12479,N_12094);
nor U13689 (N_13689,N_13099,N_12659);
and U13690 (N_13690,N_13158,N_13149);
nor U13691 (N_13691,N_12824,N_12544);
nand U13692 (N_13692,N_12719,N_12536);
nand U13693 (N_13693,N_12024,N_13150);
nor U13694 (N_13694,N_12404,N_12334);
and U13695 (N_13695,N_12559,N_12374);
and U13696 (N_13696,N_12401,N_12164);
nand U13697 (N_13697,N_12140,N_12021);
or U13698 (N_13698,N_12743,N_12682);
nand U13699 (N_13699,N_12260,N_13162);
nor U13700 (N_13700,N_12237,N_12481);
xor U13701 (N_13701,N_12054,N_12568);
and U13702 (N_13702,N_12909,N_12551);
and U13703 (N_13703,N_12014,N_12628);
and U13704 (N_13704,N_12893,N_12078);
nand U13705 (N_13705,N_13121,N_12184);
xor U13706 (N_13706,N_12517,N_12474);
xnor U13707 (N_13707,N_12264,N_12017);
xor U13708 (N_13708,N_12296,N_12811);
xnor U13709 (N_13709,N_12896,N_13113);
or U13710 (N_13710,N_12027,N_12913);
or U13711 (N_13711,N_12008,N_12792);
and U13712 (N_13712,N_13185,N_12096);
xnor U13713 (N_13713,N_12831,N_12732);
xnor U13714 (N_13714,N_12333,N_12082);
or U13715 (N_13715,N_12221,N_12250);
and U13716 (N_13716,N_12827,N_12173);
xor U13717 (N_13717,N_13164,N_12717);
nand U13718 (N_13718,N_12406,N_12669);
nor U13719 (N_13719,N_12445,N_12247);
nand U13720 (N_13720,N_12182,N_12395);
and U13721 (N_13721,N_12969,N_12772);
or U13722 (N_13722,N_12191,N_13053);
and U13723 (N_13723,N_12018,N_12654);
and U13724 (N_13724,N_12165,N_12575);
nor U13725 (N_13725,N_13031,N_12038);
or U13726 (N_13726,N_12603,N_12215);
or U13727 (N_13727,N_12084,N_13079);
or U13728 (N_13728,N_12273,N_12090);
nand U13729 (N_13729,N_12457,N_12432);
nor U13730 (N_13730,N_13036,N_12225);
nor U13731 (N_13731,N_12050,N_12685);
nand U13732 (N_13732,N_13192,N_12975);
and U13733 (N_13733,N_12415,N_13119);
or U13734 (N_13734,N_12230,N_12095);
or U13735 (N_13735,N_12519,N_12770);
or U13736 (N_13736,N_12464,N_13144);
and U13737 (N_13737,N_12097,N_13028);
xnor U13738 (N_13738,N_12664,N_12535);
or U13739 (N_13739,N_12750,N_12285);
and U13740 (N_13740,N_12645,N_12686);
and U13741 (N_13741,N_12902,N_12593);
nor U13742 (N_13742,N_13116,N_12903);
and U13743 (N_13743,N_12541,N_12633);
and U13744 (N_13744,N_12640,N_13108);
nand U13745 (N_13745,N_12370,N_12808);
and U13746 (N_13746,N_12074,N_12574);
and U13747 (N_13747,N_12053,N_13058);
and U13748 (N_13748,N_13160,N_12533);
or U13749 (N_13749,N_12244,N_12268);
nand U13750 (N_13750,N_12978,N_12890);
and U13751 (N_13751,N_12838,N_13167);
or U13752 (N_13752,N_12960,N_12857);
nor U13753 (N_13753,N_12639,N_12026);
xnor U13754 (N_13754,N_12295,N_12150);
or U13755 (N_13755,N_13104,N_12818);
xor U13756 (N_13756,N_12055,N_12630);
or U13757 (N_13757,N_12089,N_12904);
and U13758 (N_13758,N_13027,N_12867);
nand U13759 (N_13759,N_12729,N_12608);
or U13760 (N_13760,N_12783,N_12044);
nand U13761 (N_13761,N_12390,N_12326);
and U13762 (N_13762,N_12430,N_12210);
and U13763 (N_13763,N_12935,N_12046);
nor U13764 (N_13764,N_12635,N_12241);
or U13765 (N_13765,N_12833,N_12938);
nor U13766 (N_13766,N_12189,N_12337);
xor U13767 (N_13767,N_12970,N_12607);
or U13768 (N_13768,N_13148,N_12897);
nor U13769 (N_13769,N_12697,N_12547);
xnor U13770 (N_13770,N_12912,N_12177);
or U13771 (N_13771,N_12155,N_12383);
nand U13772 (N_13772,N_12701,N_12494);
nand U13773 (N_13773,N_12843,N_12471);
xor U13774 (N_13774,N_12149,N_12618);
xor U13775 (N_13775,N_12963,N_12083);
xor U13776 (N_13776,N_12249,N_12068);
and U13777 (N_13777,N_13015,N_12336);
or U13778 (N_13778,N_12674,N_12552);
xnor U13779 (N_13779,N_12566,N_12866);
nor U13780 (N_13780,N_12192,N_12612);
and U13781 (N_13781,N_12856,N_13007);
nor U13782 (N_13782,N_12245,N_12289);
and U13783 (N_13783,N_13097,N_12712);
and U13784 (N_13784,N_12234,N_12504);
nand U13785 (N_13785,N_12725,N_12282);
xnor U13786 (N_13786,N_12510,N_12817);
nand U13787 (N_13787,N_13196,N_12339);
nor U13788 (N_13788,N_12706,N_13039);
nand U13789 (N_13789,N_13009,N_12998);
and U13790 (N_13790,N_12534,N_12584);
nand U13791 (N_13791,N_12490,N_12153);
and U13792 (N_13792,N_13129,N_12366);
xor U13793 (N_13793,N_12521,N_12036);
xnor U13794 (N_13794,N_12278,N_12565);
xor U13795 (N_13795,N_12596,N_13103);
xor U13796 (N_13796,N_12197,N_12087);
or U13797 (N_13797,N_12834,N_12098);
and U13798 (N_13798,N_12284,N_12546);
nand U13799 (N_13799,N_13087,N_12687);
nor U13800 (N_13800,N_12058,N_12846);
or U13801 (N_13801,N_12258,N_12085);
and U13802 (N_13802,N_12169,N_12205);
nor U13803 (N_13803,N_12908,N_12548);
nor U13804 (N_13804,N_12615,N_12185);
or U13805 (N_13805,N_12324,N_12485);
xor U13806 (N_13806,N_13060,N_12998);
nor U13807 (N_13807,N_12719,N_12950);
xnor U13808 (N_13808,N_12465,N_12561);
xor U13809 (N_13809,N_12834,N_12156);
nor U13810 (N_13810,N_13039,N_12361);
and U13811 (N_13811,N_12933,N_12681);
xor U13812 (N_13812,N_12865,N_13063);
nor U13813 (N_13813,N_12872,N_12433);
nand U13814 (N_13814,N_12973,N_12059);
or U13815 (N_13815,N_12294,N_12553);
nand U13816 (N_13816,N_12679,N_12252);
and U13817 (N_13817,N_12688,N_12720);
and U13818 (N_13818,N_12266,N_12777);
or U13819 (N_13819,N_12644,N_13062);
nand U13820 (N_13820,N_12693,N_12962);
and U13821 (N_13821,N_12112,N_12545);
and U13822 (N_13822,N_12979,N_13109);
nor U13823 (N_13823,N_12859,N_12245);
nor U13824 (N_13824,N_13195,N_12308);
xor U13825 (N_13825,N_12968,N_12938);
xnor U13826 (N_13826,N_12925,N_13141);
nand U13827 (N_13827,N_12333,N_12867);
nand U13828 (N_13828,N_12045,N_13090);
nor U13829 (N_13829,N_12925,N_12261);
and U13830 (N_13830,N_12068,N_12139);
and U13831 (N_13831,N_12828,N_13128);
nor U13832 (N_13832,N_12044,N_13109);
or U13833 (N_13833,N_13107,N_12587);
nand U13834 (N_13834,N_12279,N_12206);
nand U13835 (N_13835,N_12648,N_13028);
nor U13836 (N_13836,N_12518,N_12003);
nor U13837 (N_13837,N_12782,N_12343);
or U13838 (N_13838,N_12996,N_13069);
nand U13839 (N_13839,N_12677,N_12893);
or U13840 (N_13840,N_12411,N_12396);
nand U13841 (N_13841,N_12632,N_13089);
or U13842 (N_13842,N_12389,N_12463);
or U13843 (N_13843,N_12519,N_12614);
xnor U13844 (N_13844,N_12745,N_12583);
nor U13845 (N_13845,N_12592,N_12835);
or U13846 (N_13846,N_12020,N_12524);
nor U13847 (N_13847,N_12897,N_12761);
or U13848 (N_13848,N_13177,N_13076);
xor U13849 (N_13849,N_12118,N_12959);
nor U13850 (N_13850,N_12081,N_13023);
nand U13851 (N_13851,N_12729,N_12206);
nand U13852 (N_13852,N_13086,N_12247);
or U13853 (N_13853,N_13050,N_12325);
and U13854 (N_13854,N_12310,N_12228);
nand U13855 (N_13855,N_13032,N_13021);
or U13856 (N_13856,N_12332,N_12454);
nand U13857 (N_13857,N_13029,N_13114);
and U13858 (N_13858,N_12606,N_12766);
nor U13859 (N_13859,N_12276,N_12473);
or U13860 (N_13860,N_12949,N_12069);
or U13861 (N_13861,N_12151,N_13035);
or U13862 (N_13862,N_12512,N_12418);
or U13863 (N_13863,N_12937,N_12430);
and U13864 (N_13864,N_12305,N_12558);
nor U13865 (N_13865,N_12959,N_12562);
and U13866 (N_13866,N_12314,N_12159);
and U13867 (N_13867,N_12112,N_12761);
or U13868 (N_13868,N_12724,N_12638);
xnor U13869 (N_13869,N_12170,N_12346);
nand U13870 (N_13870,N_12187,N_12659);
or U13871 (N_13871,N_12388,N_12364);
and U13872 (N_13872,N_12905,N_12916);
and U13873 (N_13873,N_12396,N_12403);
nor U13874 (N_13874,N_12012,N_12466);
or U13875 (N_13875,N_12719,N_12341);
nand U13876 (N_13876,N_12907,N_12675);
and U13877 (N_13877,N_12994,N_12473);
xor U13878 (N_13878,N_12373,N_13180);
nand U13879 (N_13879,N_12192,N_12146);
xor U13880 (N_13880,N_12008,N_12442);
xor U13881 (N_13881,N_12278,N_12804);
and U13882 (N_13882,N_13170,N_12352);
nand U13883 (N_13883,N_12136,N_12649);
or U13884 (N_13884,N_12817,N_12137);
nor U13885 (N_13885,N_12361,N_12608);
nor U13886 (N_13886,N_13132,N_13163);
or U13887 (N_13887,N_12600,N_12960);
nor U13888 (N_13888,N_13166,N_12961);
xor U13889 (N_13889,N_12892,N_12311);
nand U13890 (N_13890,N_12638,N_12389);
nor U13891 (N_13891,N_12667,N_12748);
nor U13892 (N_13892,N_13145,N_12798);
xor U13893 (N_13893,N_12965,N_12606);
or U13894 (N_13894,N_12789,N_12794);
and U13895 (N_13895,N_12455,N_12116);
or U13896 (N_13896,N_12278,N_13015);
nand U13897 (N_13897,N_12469,N_12189);
or U13898 (N_13898,N_12771,N_12117);
xnor U13899 (N_13899,N_13124,N_12706);
nand U13900 (N_13900,N_13091,N_12665);
nor U13901 (N_13901,N_12287,N_13009);
or U13902 (N_13902,N_12865,N_13108);
xnor U13903 (N_13903,N_13132,N_13181);
xnor U13904 (N_13904,N_12478,N_12171);
nand U13905 (N_13905,N_12932,N_12399);
nand U13906 (N_13906,N_12456,N_12057);
xor U13907 (N_13907,N_12912,N_12869);
or U13908 (N_13908,N_13162,N_12531);
nor U13909 (N_13909,N_12276,N_12086);
nand U13910 (N_13910,N_12361,N_12133);
nor U13911 (N_13911,N_12923,N_12773);
or U13912 (N_13912,N_12370,N_12113);
nand U13913 (N_13913,N_12245,N_12992);
and U13914 (N_13914,N_12003,N_12153);
nand U13915 (N_13915,N_12489,N_12160);
nor U13916 (N_13916,N_12257,N_12054);
or U13917 (N_13917,N_12395,N_13101);
nor U13918 (N_13918,N_13176,N_12806);
nor U13919 (N_13919,N_13052,N_12964);
nand U13920 (N_13920,N_12279,N_12258);
xnor U13921 (N_13921,N_13110,N_12069);
nor U13922 (N_13922,N_12916,N_12267);
nor U13923 (N_13923,N_12810,N_12838);
nand U13924 (N_13924,N_12098,N_12368);
nand U13925 (N_13925,N_12179,N_13141);
or U13926 (N_13926,N_13068,N_12974);
nor U13927 (N_13927,N_12254,N_12762);
and U13928 (N_13928,N_12019,N_13031);
xnor U13929 (N_13929,N_12344,N_12876);
or U13930 (N_13930,N_12299,N_12018);
nor U13931 (N_13931,N_13022,N_12292);
or U13932 (N_13932,N_12180,N_12080);
and U13933 (N_13933,N_12224,N_12335);
xnor U13934 (N_13934,N_12547,N_12167);
and U13935 (N_13935,N_12714,N_12754);
and U13936 (N_13936,N_13173,N_12047);
or U13937 (N_13937,N_12766,N_12259);
nor U13938 (N_13938,N_12557,N_13085);
nor U13939 (N_13939,N_13166,N_12456);
or U13940 (N_13940,N_13174,N_12361);
nor U13941 (N_13941,N_13191,N_12702);
and U13942 (N_13942,N_12172,N_13196);
or U13943 (N_13943,N_12446,N_12738);
and U13944 (N_13944,N_12445,N_12297);
or U13945 (N_13945,N_12956,N_13116);
and U13946 (N_13946,N_12797,N_13125);
nand U13947 (N_13947,N_12490,N_13102);
nand U13948 (N_13948,N_12362,N_12965);
nor U13949 (N_13949,N_12187,N_12031);
and U13950 (N_13950,N_12256,N_12995);
nand U13951 (N_13951,N_12878,N_12780);
and U13952 (N_13952,N_12561,N_12148);
nand U13953 (N_13953,N_12807,N_12886);
xnor U13954 (N_13954,N_12606,N_13012);
nand U13955 (N_13955,N_12560,N_12218);
and U13956 (N_13956,N_12235,N_12744);
xor U13957 (N_13957,N_12221,N_12148);
nand U13958 (N_13958,N_12597,N_12448);
nand U13959 (N_13959,N_12599,N_13189);
or U13960 (N_13960,N_12076,N_13059);
nor U13961 (N_13961,N_12219,N_12758);
xor U13962 (N_13962,N_12311,N_12110);
nand U13963 (N_13963,N_12971,N_12565);
nand U13964 (N_13964,N_12097,N_12131);
nor U13965 (N_13965,N_12128,N_12074);
nand U13966 (N_13966,N_13114,N_12971);
and U13967 (N_13967,N_12370,N_13092);
and U13968 (N_13968,N_12490,N_12521);
and U13969 (N_13969,N_12499,N_12159);
nand U13970 (N_13970,N_12663,N_12787);
and U13971 (N_13971,N_12711,N_13032);
nand U13972 (N_13972,N_13082,N_12730);
or U13973 (N_13973,N_12859,N_12086);
xnor U13974 (N_13974,N_12123,N_13027);
xnor U13975 (N_13975,N_12205,N_12994);
and U13976 (N_13976,N_12014,N_12261);
or U13977 (N_13977,N_12154,N_12963);
xnor U13978 (N_13978,N_12149,N_12102);
xor U13979 (N_13979,N_12588,N_12742);
xor U13980 (N_13980,N_12833,N_12149);
nand U13981 (N_13981,N_12266,N_12865);
and U13982 (N_13982,N_12451,N_12066);
nor U13983 (N_13983,N_12436,N_12483);
xor U13984 (N_13984,N_13153,N_13137);
nor U13985 (N_13985,N_12532,N_12719);
or U13986 (N_13986,N_12573,N_12758);
nand U13987 (N_13987,N_12629,N_12505);
xnor U13988 (N_13988,N_13159,N_12246);
nand U13989 (N_13989,N_12505,N_13099);
or U13990 (N_13990,N_12997,N_12586);
and U13991 (N_13991,N_13178,N_12071);
nor U13992 (N_13992,N_12928,N_12460);
xnor U13993 (N_13993,N_12076,N_12829);
or U13994 (N_13994,N_12142,N_12007);
nand U13995 (N_13995,N_12096,N_12333);
nand U13996 (N_13996,N_13077,N_13026);
and U13997 (N_13997,N_12554,N_12568);
xor U13998 (N_13998,N_12688,N_12841);
and U13999 (N_13999,N_12913,N_12698);
nor U14000 (N_14000,N_12807,N_13020);
xor U14001 (N_14001,N_12323,N_12188);
and U14002 (N_14002,N_13027,N_12353);
nor U14003 (N_14003,N_12280,N_12364);
nor U14004 (N_14004,N_12447,N_12768);
and U14005 (N_14005,N_12653,N_12588);
and U14006 (N_14006,N_12924,N_12526);
nor U14007 (N_14007,N_12000,N_12663);
or U14008 (N_14008,N_12194,N_12433);
xor U14009 (N_14009,N_13094,N_12225);
xor U14010 (N_14010,N_12818,N_12726);
nand U14011 (N_14011,N_12807,N_12709);
nand U14012 (N_14012,N_12468,N_12670);
or U14013 (N_14013,N_12459,N_12925);
xor U14014 (N_14014,N_12399,N_12386);
xor U14015 (N_14015,N_13099,N_12733);
nand U14016 (N_14016,N_12949,N_12535);
xor U14017 (N_14017,N_12415,N_12417);
nand U14018 (N_14018,N_13071,N_12803);
xnor U14019 (N_14019,N_12866,N_12198);
nand U14020 (N_14020,N_12302,N_12258);
nor U14021 (N_14021,N_12193,N_12961);
nor U14022 (N_14022,N_12541,N_12913);
or U14023 (N_14023,N_12797,N_12740);
and U14024 (N_14024,N_12864,N_12790);
nand U14025 (N_14025,N_12950,N_12293);
nand U14026 (N_14026,N_12900,N_13197);
and U14027 (N_14027,N_13005,N_12733);
or U14028 (N_14028,N_13173,N_12258);
and U14029 (N_14029,N_12248,N_12864);
nand U14030 (N_14030,N_12764,N_13164);
and U14031 (N_14031,N_12585,N_13031);
nor U14032 (N_14032,N_12075,N_12623);
nor U14033 (N_14033,N_12197,N_13131);
and U14034 (N_14034,N_13083,N_13035);
xor U14035 (N_14035,N_12783,N_12407);
or U14036 (N_14036,N_12776,N_12276);
xnor U14037 (N_14037,N_12903,N_12043);
and U14038 (N_14038,N_12124,N_12186);
nor U14039 (N_14039,N_12284,N_12177);
xor U14040 (N_14040,N_12472,N_12108);
and U14041 (N_14041,N_12384,N_12324);
nor U14042 (N_14042,N_13043,N_13050);
and U14043 (N_14043,N_13104,N_13046);
and U14044 (N_14044,N_12442,N_12720);
or U14045 (N_14045,N_13184,N_13005);
or U14046 (N_14046,N_12542,N_12786);
xnor U14047 (N_14047,N_12044,N_12626);
and U14048 (N_14048,N_12261,N_12150);
xnor U14049 (N_14049,N_12044,N_12411);
nor U14050 (N_14050,N_12877,N_12099);
and U14051 (N_14051,N_12724,N_12946);
xor U14052 (N_14052,N_12320,N_12940);
and U14053 (N_14053,N_13116,N_12144);
and U14054 (N_14054,N_12678,N_12212);
nand U14055 (N_14055,N_12414,N_12861);
nor U14056 (N_14056,N_13130,N_12361);
and U14057 (N_14057,N_13017,N_12630);
xor U14058 (N_14058,N_12506,N_12776);
nor U14059 (N_14059,N_12443,N_13121);
and U14060 (N_14060,N_12443,N_12381);
and U14061 (N_14061,N_12684,N_12481);
nand U14062 (N_14062,N_12683,N_13039);
or U14063 (N_14063,N_12153,N_12408);
nor U14064 (N_14064,N_12177,N_12832);
and U14065 (N_14065,N_12719,N_12455);
nand U14066 (N_14066,N_12890,N_12061);
and U14067 (N_14067,N_13185,N_12297);
nand U14068 (N_14068,N_12506,N_12006);
xnor U14069 (N_14069,N_12884,N_12610);
xor U14070 (N_14070,N_12816,N_12193);
and U14071 (N_14071,N_12366,N_12089);
or U14072 (N_14072,N_13089,N_13189);
xnor U14073 (N_14073,N_12998,N_12913);
xor U14074 (N_14074,N_12410,N_12774);
and U14075 (N_14075,N_12641,N_12719);
xnor U14076 (N_14076,N_12419,N_12176);
nand U14077 (N_14077,N_12968,N_12903);
nand U14078 (N_14078,N_12696,N_12004);
nand U14079 (N_14079,N_12409,N_12343);
nand U14080 (N_14080,N_12991,N_12346);
nor U14081 (N_14081,N_13083,N_12247);
xnor U14082 (N_14082,N_12686,N_13077);
nor U14083 (N_14083,N_12024,N_12522);
and U14084 (N_14084,N_13007,N_12854);
nand U14085 (N_14085,N_13069,N_12345);
or U14086 (N_14086,N_12161,N_12561);
nand U14087 (N_14087,N_12853,N_12579);
nor U14088 (N_14088,N_12692,N_12408);
or U14089 (N_14089,N_12962,N_12863);
nand U14090 (N_14090,N_13092,N_12778);
and U14091 (N_14091,N_12912,N_12446);
and U14092 (N_14092,N_12864,N_13153);
xnor U14093 (N_14093,N_13153,N_12965);
nor U14094 (N_14094,N_12812,N_12341);
and U14095 (N_14095,N_12355,N_12535);
xnor U14096 (N_14096,N_13196,N_12421);
and U14097 (N_14097,N_12409,N_12448);
or U14098 (N_14098,N_12642,N_13000);
xnor U14099 (N_14099,N_13101,N_12001);
and U14100 (N_14100,N_12341,N_12901);
nand U14101 (N_14101,N_12942,N_13058);
and U14102 (N_14102,N_13093,N_12005);
nor U14103 (N_14103,N_12912,N_12862);
and U14104 (N_14104,N_12529,N_12202);
and U14105 (N_14105,N_12404,N_12269);
and U14106 (N_14106,N_12687,N_13122);
xor U14107 (N_14107,N_12868,N_12790);
nor U14108 (N_14108,N_12587,N_13124);
or U14109 (N_14109,N_12015,N_12723);
nor U14110 (N_14110,N_12302,N_13179);
xnor U14111 (N_14111,N_12050,N_12880);
nand U14112 (N_14112,N_12336,N_13083);
and U14113 (N_14113,N_12274,N_12779);
nor U14114 (N_14114,N_12677,N_12279);
xor U14115 (N_14115,N_12720,N_13067);
xnor U14116 (N_14116,N_12851,N_12004);
nand U14117 (N_14117,N_12112,N_12981);
nand U14118 (N_14118,N_13199,N_12114);
xor U14119 (N_14119,N_12645,N_12510);
and U14120 (N_14120,N_13199,N_13039);
xnor U14121 (N_14121,N_12099,N_12004);
nor U14122 (N_14122,N_12873,N_13003);
nand U14123 (N_14123,N_12023,N_13064);
nand U14124 (N_14124,N_12430,N_13051);
and U14125 (N_14125,N_13087,N_12139);
nor U14126 (N_14126,N_12272,N_12227);
nand U14127 (N_14127,N_13103,N_12976);
nor U14128 (N_14128,N_12740,N_12332);
or U14129 (N_14129,N_12333,N_12782);
nand U14130 (N_14130,N_12587,N_12584);
or U14131 (N_14131,N_12181,N_12212);
or U14132 (N_14132,N_12133,N_12890);
or U14133 (N_14133,N_12036,N_12896);
xor U14134 (N_14134,N_12160,N_13000);
or U14135 (N_14135,N_13014,N_12085);
and U14136 (N_14136,N_12801,N_12985);
and U14137 (N_14137,N_12680,N_12715);
and U14138 (N_14138,N_13072,N_12554);
nand U14139 (N_14139,N_12881,N_12278);
or U14140 (N_14140,N_12988,N_12676);
or U14141 (N_14141,N_12447,N_12959);
nor U14142 (N_14142,N_12438,N_12426);
or U14143 (N_14143,N_12518,N_12912);
nor U14144 (N_14144,N_12269,N_12899);
xor U14145 (N_14145,N_12196,N_12214);
nor U14146 (N_14146,N_12134,N_12116);
nor U14147 (N_14147,N_12550,N_12438);
and U14148 (N_14148,N_12644,N_12719);
xnor U14149 (N_14149,N_13040,N_12665);
xnor U14150 (N_14150,N_12425,N_12206);
xor U14151 (N_14151,N_12863,N_12625);
nor U14152 (N_14152,N_12352,N_12263);
nand U14153 (N_14153,N_12754,N_12582);
or U14154 (N_14154,N_12581,N_12234);
xor U14155 (N_14155,N_12601,N_12262);
xnor U14156 (N_14156,N_12096,N_13091);
or U14157 (N_14157,N_12743,N_12496);
nor U14158 (N_14158,N_12677,N_12968);
nor U14159 (N_14159,N_13140,N_12553);
or U14160 (N_14160,N_12651,N_13064);
xor U14161 (N_14161,N_12180,N_12730);
and U14162 (N_14162,N_12826,N_12493);
or U14163 (N_14163,N_12368,N_12970);
and U14164 (N_14164,N_12028,N_12997);
and U14165 (N_14165,N_13141,N_12176);
or U14166 (N_14166,N_12837,N_12825);
nand U14167 (N_14167,N_12589,N_12014);
and U14168 (N_14168,N_12949,N_12581);
nor U14169 (N_14169,N_13097,N_12742);
nand U14170 (N_14170,N_12208,N_12118);
and U14171 (N_14171,N_12148,N_13106);
xor U14172 (N_14172,N_12792,N_12935);
nor U14173 (N_14173,N_12349,N_12554);
xor U14174 (N_14174,N_13077,N_13066);
or U14175 (N_14175,N_12471,N_12710);
and U14176 (N_14176,N_12111,N_12327);
or U14177 (N_14177,N_12528,N_12324);
nand U14178 (N_14178,N_12547,N_12648);
and U14179 (N_14179,N_12203,N_12122);
and U14180 (N_14180,N_12091,N_12896);
xnor U14181 (N_14181,N_12155,N_12165);
or U14182 (N_14182,N_12800,N_12312);
xnor U14183 (N_14183,N_12986,N_12547);
or U14184 (N_14184,N_12423,N_12046);
or U14185 (N_14185,N_12883,N_13010);
nand U14186 (N_14186,N_12560,N_12065);
and U14187 (N_14187,N_12207,N_12398);
xnor U14188 (N_14188,N_12052,N_13159);
nand U14189 (N_14189,N_12074,N_12046);
and U14190 (N_14190,N_12636,N_12843);
nor U14191 (N_14191,N_12744,N_12406);
and U14192 (N_14192,N_12558,N_12264);
or U14193 (N_14193,N_12801,N_12010);
and U14194 (N_14194,N_12923,N_12436);
and U14195 (N_14195,N_12005,N_12047);
nor U14196 (N_14196,N_12554,N_13149);
nor U14197 (N_14197,N_12657,N_12844);
nor U14198 (N_14198,N_12116,N_13180);
nand U14199 (N_14199,N_12654,N_12832);
nor U14200 (N_14200,N_12332,N_12598);
and U14201 (N_14201,N_13032,N_13056);
nand U14202 (N_14202,N_12755,N_12618);
nor U14203 (N_14203,N_12280,N_12681);
nand U14204 (N_14204,N_12613,N_12686);
and U14205 (N_14205,N_12578,N_12812);
nor U14206 (N_14206,N_12365,N_12293);
or U14207 (N_14207,N_13073,N_13082);
xor U14208 (N_14208,N_12521,N_12531);
nand U14209 (N_14209,N_12974,N_12187);
or U14210 (N_14210,N_12547,N_12691);
nor U14211 (N_14211,N_12416,N_12172);
nor U14212 (N_14212,N_12339,N_12501);
and U14213 (N_14213,N_12088,N_12675);
xor U14214 (N_14214,N_12864,N_13123);
or U14215 (N_14215,N_13001,N_12236);
and U14216 (N_14216,N_12972,N_12021);
nand U14217 (N_14217,N_12037,N_13124);
and U14218 (N_14218,N_12726,N_12986);
and U14219 (N_14219,N_12506,N_12137);
or U14220 (N_14220,N_12782,N_12394);
xnor U14221 (N_14221,N_12448,N_12411);
nand U14222 (N_14222,N_12220,N_12169);
nor U14223 (N_14223,N_12519,N_12019);
nor U14224 (N_14224,N_12436,N_12795);
nor U14225 (N_14225,N_12762,N_12655);
xor U14226 (N_14226,N_12626,N_12410);
or U14227 (N_14227,N_13176,N_13024);
nand U14228 (N_14228,N_12601,N_12614);
and U14229 (N_14229,N_12270,N_12809);
nor U14230 (N_14230,N_12082,N_12499);
or U14231 (N_14231,N_12974,N_12878);
nand U14232 (N_14232,N_12634,N_13098);
nand U14233 (N_14233,N_12375,N_12288);
or U14234 (N_14234,N_12324,N_12028);
or U14235 (N_14235,N_12737,N_12141);
nand U14236 (N_14236,N_12197,N_12617);
xnor U14237 (N_14237,N_12867,N_13082);
nor U14238 (N_14238,N_12605,N_12440);
nor U14239 (N_14239,N_13181,N_13143);
nand U14240 (N_14240,N_12822,N_13192);
and U14241 (N_14241,N_12037,N_12197);
or U14242 (N_14242,N_12680,N_12139);
nand U14243 (N_14243,N_12389,N_12686);
nor U14244 (N_14244,N_13111,N_12299);
or U14245 (N_14245,N_12015,N_12235);
nand U14246 (N_14246,N_12534,N_13113);
nor U14247 (N_14247,N_12904,N_12256);
nor U14248 (N_14248,N_12657,N_12201);
xor U14249 (N_14249,N_12174,N_12009);
nand U14250 (N_14250,N_12361,N_12704);
nand U14251 (N_14251,N_13132,N_12887);
nand U14252 (N_14252,N_12974,N_12655);
nand U14253 (N_14253,N_12333,N_12649);
or U14254 (N_14254,N_12248,N_12727);
nor U14255 (N_14255,N_13175,N_12680);
nand U14256 (N_14256,N_13000,N_12178);
xor U14257 (N_14257,N_12928,N_12043);
nand U14258 (N_14258,N_12780,N_12400);
nand U14259 (N_14259,N_12500,N_12952);
nor U14260 (N_14260,N_12684,N_12660);
xor U14261 (N_14261,N_12728,N_12687);
and U14262 (N_14262,N_12239,N_12692);
nor U14263 (N_14263,N_13102,N_12690);
nor U14264 (N_14264,N_12240,N_13146);
nor U14265 (N_14265,N_12062,N_12973);
xnor U14266 (N_14266,N_12007,N_12933);
or U14267 (N_14267,N_12830,N_12351);
nand U14268 (N_14268,N_12194,N_12011);
nor U14269 (N_14269,N_12114,N_12638);
nand U14270 (N_14270,N_12359,N_12807);
xor U14271 (N_14271,N_12441,N_12554);
nor U14272 (N_14272,N_12204,N_12812);
or U14273 (N_14273,N_12750,N_12434);
nor U14274 (N_14274,N_12938,N_12782);
xnor U14275 (N_14275,N_12063,N_12308);
or U14276 (N_14276,N_12294,N_12099);
or U14277 (N_14277,N_13019,N_12371);
and U14278 (N_14278,N_12993,N_12204);
nor U14279 (N_14279,N_12139,N_13107);
or U14280 (N_14280,N_12255,N_12880);
xor U14281 (N_14281,N_12962,N_12339);
nor U14282 (N_14282,N_12219,N_12398);
or U14283 (N_14283,N_12498,N_12964);
nor U14284 (N_14284,N_12396,N_13096);
nand U14285 (N_14285,N_12062,N_12680);
xnor U14286 (N_14286,N_12585,N_12136);
or U14287 (N_14287,N_12165,N_12354);
xnor U14288 (N_14288,N_12632,N_12136);
nand U14289 (N_14289,N_13151,N_12570);
xor U14290 (N_14290,N_13179,N_12446);
nor U14291 (N_14291,N_12016,N_12574);
and U14292 (N_14292,N_12628,N_12430);
and U14293 (N_14293,N_13199,N_13169);
or U14294 (N_14294,N_13142,N_12072);
nand U14295 (N_14295,N_12479,N_12551);
xor U14296 (N_14296,N_12001,N_12258);
and U14297 (N_14297,N_13023,N_12805);
or U14298 (N_14298,N_12164,N_12712);
xnor U14299 (N_14299,N_12306,N_12844);
or U14300 (N_14300,N_12540,N_12938);
and U14301 (N_14301,N_12796,N_12430);
xnor U14302 (N_14302,N_12905,N_12311);
nand U14303 (N_14303,N_12856,N_12779);
or U14304 (N_14304,N_13019,N_13110);
xor U14305 (N_14305,N_13032,N_12581);
nor U14306 (N_14306,N_12295,N_13037);
and U14307 (N_14307,N_12939,N_12045);
or U14308 (N_14308,N_12288,N_12962);
or U14309 (N_14309,N_12564,N_12806);
or U14310 (N_14310,N_13039,N_13055);
nand U14311 (N_14311,N_12863,N_12954);
xnor U14312 (N_14312,N_12963,N_12696);
and U14313 (N_14313,N_12355,N_12702);
xnor U14314 (N_14314,N_12642,N_12157);
and U14315 (N_14315,N_13125,N_12490);
or U14316 (N_14316,N_12579,N_13176);
and U14317 (N_14317,N_13039,N_12494);
xnor U14318 (N_14318,N_12166,N_12906);
nor U14319 (N_14319,N_12286,N_12503);
and U14320 (N_14320,N_13070,N_12641);
nand U14321 (N_14321,N_12509,N_12969);
or U14322 (N_14322,N_12495,N_12221);
or U14323 (N_14323,N_12386,N_12314);
nor U14324 (N_14324,N_12678,N_12458);
and U14325 (N_14325,N_13090,N_12268);
xor U14326 (N_14326,N_13169,N_12567);
and U14327 (N_14327,N_12800,N_13143);
nor U14328 (N_14328,N_12180,N_12361);
and U14329 (N_14329,N_12487,N_12464);
and U14330 (N_14330,N_12238,N_12656);
or U14331 (N_14331,N_12866,N_13072);
xnor U14332 (N_14332,N_12604,N_12497);
nand U14333 (N_14333,N_12670,N_12887);
nand U14334 (N_14334,N_12887,N_12939);
xor U14335 (N_14335,N_12846,N_12798);
or U14336 (N_14336,N_12853,N_12192);
and U14337 (N_14337,N_12803,N_12189);
nor U14338 (N_14338,N_13105,N_12297);
or U14339 (N_14339,N_12643,N_12859);
xor U14340 (N_14340,N_13054,N_13183);
and U14341 (N_14341,N_12667,N_12585);
nor U14342 (N_14342,N_13106,N_12391);
xor U14343 (N_14343,N_12579,N_12693);
xnor U14344 (N_14344,N_12694,N_12533);
and U14345 (N_14345,N_13034,N_12187);
nor U14346 (N_14346,N_12206,N_12401);
nor U14347 (N_14347,N_12221,N_12788);
nand U14348 (N_14348,N_12486,N_13164);
xor U14349 (N_14349,N_12351,N_12563);
and U14350 (N_14350,N_12656,N_12403);
nand U14351 (N_14351,N_12372,N_13069);
xor U14352 (N_14352,N_12743,N_12193);
xnor U14353 (N_14353,N_12356,N_13157);
or U14354 (N_14354,N_12740,N_13034);
nand U14355 (N_14355,N_12085,N_12318);
or U14356 (N_14356,N_13140,N_13010);
nand U14357 (N_14357,N_12345,N_12809);
nand U14358 (N_14358,N_12601,N_13083);
or U14359 (N_14359,N_12847,N_13057);
and U14360 (N_14360,N_12609,N_12631);
nor U14361 (N_14361,N_13196,N_12497);
nor U14362 (N_14362,N_12371,N_12488);
nor U14363 (N_14363,N_12056,N_12267);
nor U14364 (N_14364,N_12595,N_12718);
or U14365 (N_14365,N_12640,N_12114);
xor U14366 (N_14366,N_12308,N_12750);
or U14367 (N_14367,N_12001,N_12351);
nand U14368 (N_14368,N_12281,N_12017);
xor U14369 (N_14369,N_12392,N_12358);
or U14370 (N_14370,N_12779,N_12656);
nor U14371 (N_14371,N_12408,N_12053);
nor U14372 (N_14372,N_12323,N_12632);
nand U14373 (N_14373,N_12084,N_12652);
nor U14374 (N_14374,N_12081,N_12893);
or U14375 (N_14375,N_12860,N_12794);
or U14376 (N_14376,N_12312,N_12597);
nor U14377 (N_14377,N_13156,N_12113);
nor U14378 (N_14378,N_12640,N_13155);
nor U14379 (N_14379,N_12452,N_13030);
and U14380 (N_14380,N_12150,N_12417);
and U14381 (N_14381,N_13020,N_12505);
nor U14382 (N_14382,N_12793,N_12691);
or U14383 (N_14383,N_12260,N_12203);
nand U14384 (N_14384,N_12664,N_13116);
or U14385 (N_14385,N_12833,N_12012);
xnor U14386 (N_14386,N_12709,N_12495);
and U14387 (N_14387,N_12453,N_12137);
xor U14388 (N_14388,N_12534,N_12996);
or U14389 (N_14389,N_13161,N_12834);
and U14390 (N_14390,N_12800,N_12604);
or U14391 (N_14391,N_12579,N_12708);
or U14392 (N_14392,N_12816,N_12615);
and U14393 (N_14393,N_12950,N_12688);
or U14394 (N_14394,N_12003,N_12915);
nor U14395 (N_14395,N_12733,N_12272);
nor U14396 (N_14396,N_12177,N_12085);
and U14397 (N_14397,N_13062,N_12376);
and U14398 (N_14398,N_12145,N_12483);
nand U14399 (N_14399,N_13151,N_12250);
nor U14400 (N_14400,N_14118,N_14239);
or U14401 (N_14401,N_14259,N_13406);
and U14402 (N_14402,N_13980,N_13833);
or U14403 (N_14403,N_14278,N_13596);
and U14404 (N_14404,N_13299,N_13958);
nand U14405 (N_14405,N_13289,N_13531);
nor U14406 (N_14406,N_13354,N_14097);
nor U14407 (N_14407,N_14133,N_13592);
or U14408 (N_14408,N_14395,N_13840);
or U14409 (N_14409,N_13766,N_14075);
xnor U14410 (N_14410,N_13381,N_13878);
nand U14411 (N_14411,N_14169,N_13557);
or U14412 (N_14412,N_13251,N_13454);
xnor U14413 (N_14413,N_14328,N_13721);
nand U14414 (N_14414,N_14099,N_13260);
nor U14415 (N_14415,N_13527,N_14024);
nor U14416 (N_14416,N_13226,N_14195);
nand U14417 (N_14417,N_14076,N_14321);
and U14418 (N_14418,N_14369,N_13642);
xnor U14419 (N_14419,N_13464,N_14373);
nor U14420 (N_14420,N_13990,N_14359);
or U14421 (N_14421,N_13987,N_13881);
nand U14422 (N_14422,N_13385,N_14265);
and U14423 (N_14423,N_14202,N_13800);
or U14424 (N_14424,N_14150,N_13220);
or U14425 (N_14425,N_14055,N_14082);
nor U14426 (N_14426,N_13329,N_14261);
or U14427 (N_14427,N_14086,N_13972);
nand U14428 (N_14428,N_13819,N_13262);
xnor U14429 (N_14429,N_13858,N_13886);
xor U14430 (N_14430,N_14019,N_13222);
or U14431 (N_14431,N_13829,N_13818);
and U14432 (N_14432,N_13919,N_13261);
nor U14433 (N_14433,N_13509,N_13871);
xnor U14434 (N_14434,N_13974,N_13484);
nor U14435 (N_14435,N_14013,N_13643);
or U14436 (N_14436,N_13201,N_14098);
nor U14437 (N_14437,N_14111,N_13439);
xnor U14438 (N_14438,N_14052,N_14384);
or U14439 (N_14439,N_13541,N_13554);
xor U14440 (N_14440,N_13914,N_13637);
xnor U14441 (N_14441,N_13761,N_13892);
and U14442 (N_14442,N_13981,N_14290);
nand U14443 (N_14443,N_13434,N_13920);
nand U14444 (N_14444,N_13614,N_14388);
or U14445 (N_14445,N_14138,N_13380);
or U14446 (N_14446,N_14152,N_14192);
xnor U14447 (N_14447,N_14029,N_13444);
or U14448 (N_14448,N_14092,N_14326);
and U14449 (N_14449,N_13896,N_14208);
and U14450 (N_14450,N_13340,N_13518);
nand U14451 (N_14451,N_14054,N_13505);
or U14452 (N_14452,N_13535,N_14323);
and U14453 (N_14453,N_13310,N_13238);
or U14454 (N_14454,N_14318,N_14053);
nor U14455 (N_14455,N_13760,N_13901);
xor U14456 (N_14456,N_13695,N_13243);
xnor U14457 (N_14457,N_13232,N_13301);
nand U14458 (N_14458,N_13269,N_13536);
nand U14459 (N_14459,N_13514,N_14116);
nor U14460 (N_14460,N_14088,N_14377);
xnor U14461 (N_14461,N_14194,N_14007);
nor U14462 (N_14462,N_14205,N_13580);
or U14463 (N_14463,N_13248,N_14238);
nand U14464 (N_14464,N_14347,N_13864);
and U14465 (N_14465,N_13801,N_13868);
or U14466 (N_14466,N_13526,N_13334);
nor U14467 (N_14467,N_13587,N_13319);
nand U14468 (N_14468,N_13317,N_13324);
nand U14469 (N_14469,N_13994,N_13652);
xnor U14470 (N_14470,N_14008,N_13433);
and U14471 (N_14471,N_13883,N_13409);
xnor U14472 (N_14472,N_14064,N_13333);
or U14473 (N_14473,N_13362,N_14067);
nand U14474 (N_14474,N_13750,N_13615);
and U14475 (N_14475,N_13784,N_13335);
xnor U14476 (N_14476,N_14301,N_13962);
nor U14477 (N_14477,N_13223,N_13459);
nor U14478 (N_14478,N_14394,N_13523);
nand U14479 (N_14479,N_13879,N_13537);
xnor U14480 (N_14480,N_14363,N_14317);
xor U14481 (N_14481,N_13744,N_14014);
nand U14482 (N_14482,N_13658,N_14002);
nand U14483 (N_14483,N_14083,N_14016);
or U14484 (N_14484,N_14179,N_13428);
and U14485 (N_14485,N_14050,N_13339);
nand U14486 (N_14486,N_13612,N_13233);
and U14487 (N_14487,N_14268,N_13870);
or U14488 (N_14488,N_13702,N_13715);
nand U14489 (N_14489,N_13641,N_13574);
nor U14490 (N_14490,N_14135,N_14140);
or U14491 (N_14491,N_14351,N_13672);
nand U14492 (N_14492,N_13487,N_14249);
or U14493 (N_14493,N_13613,N_13500);
nor U14494 (N_14494,N_13511,N_13465);
and U14495 (N_14495,N_13741,N_13777);
nor U14496 (N_14496,N_13899,N_14070);
nor U14497 (N_14497,N_13813,N_13968);
nor U14498 (N_14498,N_13351,N_13595);
and U14499 (N_14499,N_14187,N_14314);
nand U14500 (N_14500,N_13255,N_13869);
or U14501 (N_14501,N_14170,N_13325);
or U14502 (N_14502,N_13649,N_13298);
xnor U14503 (N_14503,N_13492,N_13372);
nor U14504 (N_14504,N_13679,N_13431);
xnor U14505 (N_14505,N_13735,N_13314);
nand U14506 (N_14506,N_14324,N_13685);
or U14507 (N_14507,N_13689,N_13982);
nor U14508 (N_14508,N_13258,N_14391);
nand U14509 (N_14509,N_13359,N_14224);
xor U14510 (N_14510,N_13648,N_13900);
nand U14511 (N_14511,N_14038,N_13476);
nor U14512 (N_14512,N_13483,N_14119);
xnor U14513 (N_14513,N_13722,N_13418);
xnor U14514 (N_14514,N_13585,N_14085);
or U14515 (N_14515,N_13664,N_13543);
or U14516 (N_14516,N_13323,N_13215);
nand U14517 (N_14517,N_14344,N_13307);
xnor U14518 (N_14518,N_13217,N_13618);
xnor U14519 (N_14519,N_13635,N_13558);
nand U14520 (N_14520,N_13657,N_13674);
nor U14521 (N_14521,N_13802,N_13731);
or U14522 (N_14522,N_13562,N_13403);
and U14523 (N_14523,N_14376,N_13769);
nand U14524 (N_14524,N_13793,N_13396);
or U14525 (N_14525,N_14298,N_13929);
xnor U14526 (N_14526,N_13302,N_13716);
xnor U14527 (N_14527,N_14327,N_13676);
nor U14528 (N_14528,N_13283,N_13330);
nand U14529 (N_14529,N_13320,N_13336);
nor U14530 (N_14530,N_14343,N_14236);
and U14531 (N_14531,N_13873,N_13321);
and U14532 (N_14532,N_13742,N_13771);
nand U14533 (N_14533,N_13825,N_14188);
and U14534 (N_14534,N_14059,N_14313);
and U14535 (N_14535,N_14158,N_14003);
xor U14536 (N_14536,N_14386,N_13416);
nor U14537 (N_14537,N_13862,N_13895);
or U14538 (N_14538,N_13304,N_14330);
and U14539 (N_14539,N_14271,N_14137);
or U14540 (N_14540,N_14307,N_14229);
and U14541 (N_14541,N_13457,N_14399);
and U14542 (N_14542,N_14032,N_14235);
and U14543 (N_14543,N_14272,N_14043);
or U14544 (N_14544,N_14030,N_13882);
nand U14545 (N_14545,N_14385,N_13593);
xor U14546 (N_14546,N_14335,N_13207);
or U14547 (N_14547,N_13315,N_13377);
or U14548 (N_14548,N_13241,N_14380);
xnor U14549 (N_14549,N_13728,N_14291);
nor U14550 (N_14550,N_14247,N_14181);
nand U14551 (N_14551,N_13538,N_13610);
nand U14552 (N_14552,N_13291,N_13564);
nor U14553 (N_14553,N_14215,N_13775);
nor U14554 (N_14554,N_13216,N_14129);
and U14555 (N_14555,N_14080,N_14371);
nor U14556 (N_14556,N_13639,N_13525);
and U14557 (N_14557,N_13252,N_14035);
or U14558 (N_14558,N_13256,N_14046);
nor U14559 (N_14559,N_14387,N_13502);
nor U14560 (N_14560,N_13270,N_13203);
xnor U14561 (N_14561,N_13979,N_13874);
nand U14562 (N_14562,N_13601,N_13908);
nand U14563 (N_14563,N_13210,N_13382);
xnor U14564 (N_14564,N_13563,N_14182);
nor U14565 (N_14565,N_13369,N_13582);
and U14566 (N_14566,N_13988,N_13897);
or U14567 (N_14567,N_13785,N_13350);
nor U14568 (N_14568,N_14203,N_13508);
or U14569 (N_14569,N_14154,N_13296);
and U14570 (N_14570,N_13844,N_13237);
and U14571 (N_14571,N_14364,N_13501);
nor U14572 (N_14572,N_14322,N_13532);
xnor U14573 (N_14573,N_14079,N_13719);
nor U14574 (N_14574,N_14090,N_14176);
or U14575 (N_14575,N_14036,N_14108);
nand U14576 (N_14576,N_14257,N_14393);
and U14577 (N_14577,N_14222,N_14153);
or U14578 (N_14578,N_14381,N_13933);
xor U14579 (N_14579,N_13423,N_14213);
or U14580 (N_14580,N_14355,N_13412);
nor U14581 (N_14581,N_14284,N_13673);
nand U14582 (N_14582,N_13277,N_13206);
nor U14583 (N_14583,N_14103,N_13746);
and U14584 (N_14584,N_14311,N_13947);
and U14585 (N_14585,N_13907,N_13992);
or U14586 (N_14586,N_13460,N_13725);
xnor U14587 (N_14587,N_14071,N_14066);
or U14588 (N_14588,N_13584,N_14360);
or U14589 (N_14589,N_13455,N_13628);
nand U14590 (N_14590,N_14214,N_13821);
or U14591 (N_14591,N_14254,N_14146);
nor U14592 (N_14592,N_13572,N_14274);
xor U14593 (N_14593,N_13687,N_13281);
or U14594 (N_14594,N_13627,N_13653);
xnor U14595 (N_14595,N_14042,N_13265);
xnor U14596 (N_14596,N_13569,N_13540);
nor U14597 (N_14597,N_14012,N_13948);
nand U14598 (N_14598,N_13686,N_14379);
nand U14599 (N_14599,N_13857,N_13565);
and U14600 (N_14600,N_13512,N_13791);
nand U14601 (N_14601,N_14011,N_13834);
and U14602 (N_14602,N_13597,N_13453);
xor U14603 (N_14603,N_13747,N_13544);
nor U14604 (N_14604,N_14068,N_13282);
or U14605 (N_14605,N_14025,N_13472);
nor U14606 (N_14606,N_13338,N_13894);
nor U14607 (N_14607,N_13309,N_14173);
and U14608 (N_14608,N_13401,N_13630);
nand U14609 (N_14609,N_13959,N_13488);
and U14610 (N_14610,N_14230,N_14287);
nand U14611 (N_14611,N_13799,N_14329);
and U14612 (N_14612,N_13790,N_13524);
nand U14613 (N_14613,N_13634,N_14006);
nor U14614 (N_14614,N_14056,N_14017);
nor U14615 (N_14615,N_13528,N_13481);
nor U14616 (N_14616,N_13814,N_13400);
xor U14617 (N_14617,N_14275,N_13780);
nand U14618 (N_14618,N_13954,N_14115);
and U14619 (N_14619,N_13545,N_14362);
or U14620 (N_14620,N_13724,N_13713);
nand U14621 (N_14621,N_13579,N_13463);
and U14622 (N_14622,N_14094,N_13665);
or U14623 (N_14623,N_14340,N_14241);
xor U14624 (N_14624,N_14382,N_13890);
nand U14625 (N_14625,N_13495,N_13342);
xor U14626 (N_14626,N_13397,N_13430);
nor U14627 (N_14627,N_13683,N_13930);
xor U14628 (N_14628,N_14201,N_14288);
xnor U14629 (N_14629,N_14005,N_13424);
xnor U14630 (N_14630,N_13837,N_14034);
or U14631 (N_14631,N_13308,N_13690);
xor U14632 (N_14632,N_13231,N_14246);
xnor U14633 (N_14633,N_14104,N_14061);
nor U14634 (N_14634,N_14352,N_14296);
xnor U14635 (N_14635,N_13976,N_13473);
nor U14636 (N_14636,N_13998,N_13957);
nand U14637 (N_14637,N_13697,N_13675);
or U14638 (N_14638,N_13244,N_13263);
xor U14639 (N_14639,N_13313,N_13221);
nand U14640 (N_14640,N_14255,N_13559);
nor U14641 (N_14641,N_13969,N_14087);
xnor U14642 (N_14642,N_14252,N_13376);
or U14643 (N_14643,N_13842,N_13264);
or U14644 (N_14644,N_13922,N_14081);
nor U14645 (N_14645,N_14200,N_14357);
or U14646 (N_14646,N_13816,N_14130);
nor U14647 (N_14647,N_14027,N_13576);
xnor U14648 (N_14648,N_14175,N_14000);
and U14649 (N_14649,N_13305,N_13796);
xor U14650 (N_14650,N_13848,N_13529);
nor U14651 (N_14651,N_13978,N_13876);
nor U14652 (N_14652,N_14033,N_13577);
nor U14653 (N_14653,N_14009,N_14049);
nor U14654 (N_14654,N_13451,N_14292);
nor U14655 (N_14655,N_13971,N_14190);
or U14656 (N_14656,N_14375,N_13462);
nor U14657 (N_14657,N_13865,N_13357);
nand U14658 (N_14658,N_13918,N_13290);
nand U14659 (N_14659,N_13708,N_13950);
xor U14660 (N_14660,N_13271,N_13245);
xor U14661 (N_14661,N_13347,N_14223);
nor U14662 (N_14662,N_13847,N_13754);
nand U14663 (N_14663,N_13999,N_13975);
nor U14664 (N_14664,N_13411,N_14279);
and U14665 (N_14665,N_13547,N_13375);
or U14666 (N_14666,N_13694,N_14171);
or U14667 (N_14667,N_14177,N_14073);
and U14668 (N_14668,N_13311,N_13696);
or U14669 (N_14669,N_14167,N_14302);
or U14670 (N_14670,N_13611,N_13989);
nor U14671 (N_14671,N_13405,N_13352);
and U14672 (N_14672,N_14240,N_13358);
or U14673 (N_14673,N_13925,N_13909);
nand U14674 (N_14674,N_14101,N_13651);
xnor U14675 (N_14675,N_13752,N_13966);
and U14676 (N_14676,N_14178,N_13884);
nor U14677 (N_14677,N_13360,N_14022);
or U14678 (N_14678,N_13860,N_13927);
and U14679 (N_14679,N_13578,N_13437);
or U14680 (N_14680,N_13893,N_13661);
or U14681 (N_14681,N_13568,N_14227);
or U14682 (N_14682,N_13407,N_13867);
nor U14683 (N_14683,N_14132,N_13205);
xnor U14684 (N_14684,N_13475,N_13445);
nand U14685 (N_14685,N_14112,N_13489);
nor U14686 (N_14686,N_14004,N_14157);
and U14687 (N_14687,N_13300,N_13733);
or U14688 (N_14688,N_13371,N_14370);
nor U14689 (N_14689,N_13419,N_13240);
xor U14690 (N_14690,N_14131,N_13964);
or U14691 (N_14691,N_13792,N_14039);
nor U14692 (N_14692,N_13285,N_14295);
nand U14693 (N_14693,N_13831,N_13436);
nand U14694 (N_14694,N_13940,N_14361);
or U14695 (N_14695,N_13478,N_14297);
nand U14696 (N_14696,N_13705,N_13700);
nor U14697 (N_14697,N_13200,N_13228);
or U14698 (N_14698,N_13316,N_14306);
nor U14699 (N_14699,N_13448,N_13822);
xor U14700 (N_14700,N_13655,N_13779);
and U14701 (N_14701,N_13743,N_13951);
and U14702 (N_14702,N_13880,N_13588);
xor U14703 (N_14703,N_14078,N_13917);
nand U14704 (N_14704,N_13905,N_13830);
or U14705 (N_14705,N_14122,N_13506);
nand U14706 (N_14706,N_14262,N_14256);
nand U14707 (N_14707,N_14114,N_14031);
and U14708 (N_14708,N_14172,N_13803);
or U14709 (N_14709,N_14069,N_14197);
xnor U14710 (N_14710,N_14305,N_14156);
xnor U14711 (N_14711,N_14209,N_13961);
nor U14712 (N_14712,N_13985,N_14077);
and U14713 (N_14713,N_13332,N_13392);
nor U14714 (N_14714,N_13727,N_13364);
nor U14715 (N_14715,N_13759,N_13275);
or U14716 (N_14716,N_13219,N_14220);
nand U14717 (N_14717,N_13622,N_14123);
nor U14718 (N_14718,N_13303,N_13758);
and U14719 (N_14719,N_13234,N_13402);
nand U14720 (N_14720,N_13770,N_13503);
or U14721 (N_14721,N_13935,N_14163);
nor U14722 (N_14722,N_13534,N_14372);
and U14723 (N_14723,N_13671,N_13680);
or U14724 (N_14724,N_13812,N_14285);
and U14725 (N_14725,N_13608,N_13660);
nor U14726 (N_14726,N_13707,N_13517);
nor U14727 (N_14727,N_13349,N_14196);
or U14728 (N_14728,N_13212,N_13942);
and U14729 (N_14729,N_14367,N_13482);
nand U14730 (N_14730,N_14392,N_13768);
or U14731 (N_14731,N_13274,N_14155);
nand U14732 (N_14732,N_13328,N_13549);
or U14733 (N_14733,N_13516,N_13753);
and U14734 (N_14734,N_13997,N_13717);
nor U14735 (N_14735,N_14147,N_14001);
and U14736 (N_14736,N_14183,N_13539);
or U14737 (N_14737,N_13378,N_13471);
nor U14738 (N_14738,N_13945,N_13776);
nor U14739 (N_14739,N_13726,N_14164);
nand U14740 (N_14740,N_13678,N_14126);
nand U14741 (N_14741,N_14339,N_13730);
nand U14742 (N_14742,N_13710,N_13810);
xor U14743 (N_14743,N_13924,N_13936);
nor U14744 (N_14744,N_13772,N_14331);
xnor U14745 (N_14745,N_14342,N_13513);
or U14746 (N_14746,N_13845,N_13941);
and U14747 (N_14747,N_13370,N_14110);
or U14748 (N_14748,N_14136,N_14269);
and U14749 (N_14749,N_14251,N_13943);
and U14750 (N_14750,N_13607,N_13640);
and U14751 (N_14751,N_13806,N_13440);
or U14752 (N_14752,N_14300,N_13395);
nor U14753 (N_14753,N_13751,N_14020);
nand U14754 (N_14754,N_13490,N_14266);
or U14755 (N_14755,N_14180,N_14219);
nand U14756 (N_14756,N_13225,N_13394);
or U14757 (N_14757,N_13877,N_13254);
nor U14758 (N_14758,N_14141,N_13497);
or U14759 (N_14759,N_13452,N_13645);
or U14760 (N_14760,N_14121,N_14037);
nor U14761 (N_14761,N_13820,N_14289);
xnor U14762 (N_14762,N_13838,N_14160);
nand U14763 (N_14763,N_13561,N_14074);
and U14764 (N_14764,N_14159,N_13684);
nand U14765 (N_14765,N_13552,N_13781);
nor U14766 (N_14766,N_14354,N_13599);
nor U14767 (N_14767,N_14293,N_13422);
nand U14768 (N_14768,N_13404,N_13938);
nor U14769 (N_14769,N_13590,N_13594);
nor U14770 (N_14770,N_14117,N_13361);
nand U14771 (N_14771,N_14063,N_13573);
and U14772 (N_14772,N_13408,N_13732);
nand U14773 (N_14773,N_13811,N_13609);
or U14774 (N_14774,N_13923,N_14162);
or U14775 (N_14775,N_14089,N_13835);
xor U14776 (N_14776,N_13331,N_13209);
nor U14777 (N_14777,N_14198,N_13934);
xor U14778 (N_14778,N_13662,N_13327);
nand U14779 (N_14779,N_13783,N_13738);
and U14780 (N_14780,N_13773,N_13891);
or U14781 (N_14781,N_14283,N_14148);
and U14782 (N_14782,N_13712,N_13571);
xnor U14783 (N_14783,N_13774,N_14258);
nor U14784 (N_14784,N_13853,N_14026);
or U14785 (N_14785,N_13787,N_13602);
or U14786 (N_14786,N_14174,N_13931);
nor U14787 (N_14787,N_13242,N_14028);
nor U14788 (N_14788,N_13953,N_13496);
xnor U14789 (N_14789,N_14319,N_13861);
xor U14790 (N_14790,N_14398,N_14109);
and U14791 (N_14791,N_13236,N_14270);
and U14792 (N_14792,N_13669,N_14096);
or U14793 (N_14793,N_13619,N_13211);
nor U14794 (N_14794,N_13967,N_13863);
nand U14795 (N_14795,N_14366,N_13729);
nand U14796 (N_14796,N_13677,N_13856);
nand U14797 (N_14797,N_14310,N_13485);
xor U14798 (N_14798,N_14397,N_13410);
nand U14799 (N_14799,N_13912,N_13704);
and U14800 (N_14800,N_14166,N_13970);
nand U14801 (N_14801,N_13949,N_14231);
nor U14802 (N_14802,N_14084,N_14184);
and U14803 (N_14803,N_13701,N_14228);
nor U14804 (N_14804,N_13295,N_13698);
or U14805 (N_14805,N_14165,N_13583);
and U14806 (N_14806,N_14294,N_13515);
or U14807 (N_14807,N_13447,N_13986);
nand U14808 (N_14808,N_13548,N_13956);
nor U14809 (N_14809,N_13960,N_13996);
nand U14810 (N_14810,N_13441,N_13467);
or U14811 (N_14811,N_13429,N_13550);
and U14812 (N_14812,N_14018,N_13762);
xor U14813 (N_14813,N_13326,N_13581);
or U14814 (N_14814,N_13510,N_13629);
and U14815 (N_14815,N_13763,N_13356);
and U14816 (N_14816,N_13626,N_14334);
nor U14817 (N_14817,N_14142,N_13341);
or U14818 (N_14818,N_13851,N_14374);
nand U14819 (N_14819,N_13991,N_13681);
xnor U14820 (N_14820,N_13383,N_14124);
and U14821 (N_14821,N_13693,N_13470);
nand U14822 (N_14822,N_14341,N_13832);
and U14823 (N_14823,N_14045,N_13239);
or U14824 (N_14824,N_13827,N_13213);
nor U14825 (N_14825,N_13666,N_13414);
and U14826 (N_14826,N_13692,N_13656);
or U14827 (N_14827,N_13556,N_13723);
nor U14828 (N_14828,N_13415,N_13287);
nand U14829 (N_14829,N_13253,N_14051);
nand U14830 (N_14830,N_13426,N_14368);
nand U14831 (N_14831,N_14041,N_13390);
nor U14832 (N_14832,N_14396,N_13343);
and U14833 (N_14833,N_13667,N_13247);
nand U14834 (N_14834,N_13363,N_14100);
nor U14835 (N_14835,N_13450,N_13788);
xor U14836 (N_14836,N_13946,N_13278);
xor U14837 (N_14837,N_13284,N_13650);
nand U14838 (N_14838,N_13519,N_13420);
nor U14839 (N_14839,N_14226,N_13826);
nor U14840 (N_14840,N_13560,N_13566);
xor U14841 (N_14841,N_13855,N_14149);
and U14842 (N_14842,N_14057,N_13469);
or U14843 (N_14843,N_14023,N_14242);
nor U14844 (N_14844,N_14316,N_14207);
or U14845 (N_14845,N_13765,N_13898);
nor U14846 (N_14846,N_14102,N_13542);
xnor U14847 (N_14847,N_14345,N_13983);
nand U14848 (N_14848,N_14062,N_13466);
nand U14849 (N_14849,N_14212,N_13663);
nand U14850 (N_14850,N_13312,N_13911);
or U14851 (N_14851,N_13745,N_13259);
and U14852 (N_14852,N_13734,N_14048);
or U14853 (N_14853,N_13872,N_13421);
or U14854 (N_14854,N_14337,N_13794);
xnor U14855 (N_14855,N_13276,N_13963);
or U14856 (N_14856,N_14346,N_13366);
nor U14857 (N_14857,N_13555,N_13798);
and U14858 (N_14858,N_13913,N_13229);
or U14859 (N_14859,N_13432,N_14145);
xnor U14860 (N_14860,N_13944,N_13984);
nand U14861 (N_14861,N_13399,N_14134);
and U14862 (N_14862,N_13670,N_14234);
and U14863 (N_14863,N_13435,N_13250);
or U14864 (N_14864,N_13266,N_13644);
nand U14865 (N_14865,N_13346,N_13633);
and U14866 (N_14866,N_13995,N_13294);
or U14867 (N_14867,N_13740,N_13617);
and U14868 (N_14868,N_14253,N_14325);
and U14869 (N_14869,N_13218,N_13417);
nor U14870 (N_14870,N_13442,N_13965);
nand U14871 (N_14871,N_13368,N_13293);
xnor U14872 (N_14872,N_13606,N_14303);
or U14873 (N_14873,N_13272,N_13230);
xnor U14874 (N_14874,N_13720,N_13688);
xnor U14875 (N_14875,N_13507,N_13711);
and U14876 (N_14876,N_13279,N_13456);
xor U14877 (N_14877,N_13739,N_14093);
xnor U14878 (N_14878,N_13443,N_13621);
nand U14879 (N_14879,N_13374,N_14065);
xnor U14880 (N_14880,N_13393,N_14333);
and U14881 (N_14881,N_13446,N_13292);
nor U14882 (N_14882,N_13498,N_14193);
nand U14883 (N_14883,N_14199,N_13849);
nor U14884 (N_14884,N_14273,N_13480);
or U14885 (N_14885,N_13915,N_13389);
nor U14886 (N_14886,N_14233,N_13932);
or U14887 (N_14887,N_13224,N_14365);
and U14888 (N_14888,N_13468,N_14204);
nor U14889 (N_14889,N_13551,N_13714);
nor U14890 (N_14890,N_13204,N_14245);
nand U14891 (N_14891,N_14315,N_13386);
and U14892 (N_14892,N_14106,N_13921);
or U14893 (N_14893,N_13208,N_13438);
or U14894 (N_14894,N_13257,N_14021);
nor U14895 (N_14895,N_14383,N_13477);
xnor U14896 (N_14896,N_14277,N_14047);
and U14897 (N_14897,N_14095,N_13504);
xnor U14898 (N_14898,N_14358,N_13249);
nand U14899 (N_14899,N_14232,N_13993);
and U14900 (N_14900,N_13553,N_13699);
xor U14901 (N_14901,N_13227,N_14151);
and U14902 (N_14902,N_13384,N_13246);
or U14903 (N_14903,N_13398,N_13767);
and U14904 (N_14904,N_13928,N_13631);
or U14905 (N_14905,N_13839,N_13906);
xnor U14906 (N_14906,N_13479,N_13808);
xnor U14907 (N_14907,N_13952,N_13598);
nor U14908 (N_14908,N_13904,N_14091);
nor U14909 (N_14909,N_13567,N_13373);
nor U14910 (N_14910,N_13636,N_13625);
and U14911 (N_14911,N_14304,N_13824);
and U14912 (N_14912,N_13691,N_14389);
xnor U14913 (N_14913,N_14264,N_13903);
or U14914 (N_14914,N_13388,N_14143);
xnor U14915 (N_14915,N_14010,N_13854);
nor U14916 (N_14916,N_13570,N_13910);
nor U14917 (N_14917,N_14216,N_13977);
xnor U14918 (N_14918,N_13875,N_13709);
and U14919 (N_14919,N_14186,N_13591);
or U14920 (N_14920,N_13782,N_13344);
and U14921 (N_14921,N_14237,N_13306);
or U14922 (N_14922,N_14015,N_13520);
nor U14923 (N_14923,N_13926,N_14282);
nand U14924 (N_14924,N_13586,N_13297);
nor U14925 (N_14925,N_14225,N_13843);
or U14926 (N_14926,N_14040,N_13797);
nand U14927 (N_14927,N_14105,N_13322);
and U14928 (N_14928,N_13850,N_13624);
nand U14929 (N_14929,N_14308,N_13391);
and U14930 (N_14930,N_13286,N_14125);
nor U14931 (N_14931,N_13682,N_13805);
xor U14932 (N_14932,N_13888,N_13387);
nor U14933 (N_14933,N_14072,N_13846);
xor U14934 (N_14934,N_14243,N_14144);
or U14935 (N_14935,N_14353,N_13623);
nand U14936 (N_14936,N_14338,N_13647);
and U14937 (N_14937,N_13499,N_14349);
xor U14938 (N_14938,N_13546,N_13638);
xor U14939 (N_14939,N_13795,N_14332);
nand U14940 (N_14940,N_13337,N_14286);
and U14941 (N_14941,N_13522,N_13887);
nand U14942 (N_14942,N_14107,N_14210);
nand U14943 (N_14943,N_13267,N_13807);
and U14944 (N_14944,N_13449,N_13916);
xor U14945 (N_14945,N_14267,N_13703);
xnor U14946 (N_14946,N_14320,N_14250);
and U14947 (N_14947,N_13786,N_13425);
or U14948 (N_14948,N_13575,N_14263);
nand U14949 (N_14949,N_14299,N_13836);
nor U14950 (N_14950,N_14189,N_13804);
or U14951 (N_14951,N_13273,N_13737);
and U14952 (N_14952,N_13789,N_13474);
nand U14953 (N_14953,N_13603,N_14350);
and U14954 (N_14954,N_13530,N_14113);
nor U14955 (N_14955,N_13491,N_14206);
xnor U14956 (N_14956,N_14248,N_13706);
and U14957 (N_14957,N_13600,N_13268);
and U14958 (N_14958,N_13458,N_14218);
nor U14959 (N_14959,N_13736,N_13748);
and U14960 (N_14960,N_14161,N_14336);
xnor U14961 (N_14961,N_14260,N_13866);
nand U14962 (N_14962,N_13202,N_14390);
or U14963 (N_14963,N_13345,N_14191);
xor U14964 (N_14964,N_14058,N_13214);
nand U14965 (N_14965,N_14221,N_14168);
or U14966 (N_14966,N_14128,N_13756);
and U14967 (N_14967,N_14280,N_13486);
nor U14968 (N_14968,N_13280,N_13521);
nor U14969 (N_14969,N_14120,N_13604);
or U14970 (N_14970,N_13620,N_13764);
nor U14971 (N_14971,N_14139,N_14217);
xor U14972 (N_14972,N_13427,N_13605);
xnor U14973 (N_14973,N_13817,N_13646);
or U14974 (N_14974,N_13902,N_13348);
nor U14975 (N_14975,N_13859,N_13955);
xor U14976 (N_14976,N_14185,N_14312);
xnor U14977 (N_14977,N_13757,N_13885);
xor U14978 (N_14978,N_13318,N_14244);
or U14979 (N_14979,N_13823,N_13533);
or U14980 (N_14980,N_14378,N_13589);
nor U14981 (N_14981,N_14060,N_13632);
xor U14982 (N_14982,N_13828,N_14127);
nand U14983 (N_14983,N_13288,N_13939);
nor U14984 (N_14984,N_13718,N_13668);
nand U14985 (N_14985,N_13937,N_13778);
and U14986 (N_14986,N_13494,N_13616);
nand U14987 (N_14987,N_13379,N_14276);
nor U14988 (N_14988,N_13413,N_13654);
or U14989 (N_14989,N_13659,N_13367);
nand U14990 (N_14990,N_13889,N_13852);
and U14991 (N_14991,N_14281,N_14309);
nand U14992 (N_14992,N_13749,N_14348);
nor U14993 (N_14993,N_13355,N_13841);
or U14994 (N_14994,N_13353,N_14356);
and U14995 (N_14995,N_13973,N_13755);
nand U14996 (N_14996,N_13493,N_13815);
nand U14997 (N_14997,N_13365,N_13809);
nand U14998 (N_14998,N_14211,N_13235);
or U14999 (N_14999,N_13461,N_14044);
xnor U15000 (N_15000,N_14209,N_13732);
xnor U15001 (N_15001,N_13215,N_14162);
or U15002 (N_15002,N_13895,N_14308);
nor U15003 (N_15003,N_13861,N_13557);
nor U15004 (N_15004,N_13643,N_14393);
xor U15005 (N_15005,N_13397,N_13445);
and U15006 (N_15006,N_13864,N_14139);
and U15007 (N_15007,N_13358,N_13547);
and U15008 (N_15008,N_13954,N_13505);
nand U15009 (N_15009,N_13235,N_13809);
nor U15010 (N_15010,N_13636,N_13213);
nor U15011 (N_15011,N_13395,N_13312);
nand U15012 (N_15012,N_13526,N_14378);
and U15013 (N_15013,N_13982,N_14252);
and U15014 (N_15014,N_14294,N_13366);
or U15015 (N_15015,N_13446,N_13645);
nor U15016 (N_15016,N_13796,N_13496);
xnor U15017 (N_15017,N_13311,N_13270);
and U15018 (N_15018,N_13260,N_13528);
or U15019 (N_15019,N_13651,N_13475);
and U15020 (N_15020,N_14195,N_13878);
nor U15021 (N_15021,N_13939,N_13242);
or U15022 (N_15022,N_13884,N_13659);
or U15023 (N_15023,N_14019,N_14132);
nand U15024 (N_15024,N_14037,N_13364);
nor U15025 (N_15025,N_13779,N_14030);
xor U15026 (N_15026,N_14010,N_13964);
and U15027 (N_15027,N_13926,N_13609);
xnor U15028 (N_15028,N_13679,N_14215);
xor U15029 (N_15029,N_13455,N_13618);
xor U15030 (N_15030,N_13447,N_13837);
or U15031 (N_15031,N_13246,N_13484);
and U15032 (N_15032,N_14085,N_13804);
nor U15033 (N_15033,N_14333,N_14392);
and U15034 (N_15034,N_14053,N_14155);
xnor U15035 (N_15035,N_13606,N_13925);
and U15036 (N_15036,N_13891,N_13565);
and U15037 (N_15037,N_14212,N_14284);
xnor U15038 (N_15038,N_13412,N_13678);
or U15039 (N_15039,N_13379,N_13871);
xnor U15040 (N_15040,N_14100,N_13452);
and U15041 (N_15041,N_14295,N_13937);
or U15042 (N_15042,N_13744,N_13943);
nor U15043 (N_15043,N_14149,N_13868);
and U15044 (N_15044,N_13826,N_13848);
nand U15045 (N_15045,N_13557,N_13277);
and U15046 (N_15046,N_14004,N_13768);
xor U15047 (N_15047,N_13467,N_13710);
nand U15048 (N_15048,N_13746,N_13649);
or U15049 (N_15049,N_14251,N_13691);
nand U15050 (N_15050,N_13587,N_13387);
xnor U15051 (N_15051,N_13224,N_14088);
nor U15052 (N_15052,N_13895,N_13412);
and U15053 (N_15053,N_13610,N_13286);
nor U15054 (N_15054,N_14098,N_13485);
or U15055 (N_15055,N_13222,N_13287);
nor U15056 (N_15056,N_14141,N_13293);
and U15057 (N_15057,N_14313,N_14007);
nor U15058 (N_15058,N_13398,N_13691);
nor U15059 (N_15059,N_13715,N_13352);
nand U15060 (N_15060,N_13910,N_14235);
or U15061 (N_15061,N_13861,N_13992);
nand U15062 (N_15062,N_13394,N_13511);
xor U15063 (N_15063,N_13211,N_13462);
nor U15064 (N_15064,N_13271,N_13694);
and U15065 (N_15065,N_14174,N_14043);
nand U15066 (N_15066,N_13427,N_14340);
or U15067 (N_15067,N_14107,N_13819);
or U15068 (N_15068,N_13813,N_14302);
or U15069 (N_15069,N_14279,N_14330);
nor U15070 (N_15070,N_13788,N_14229);
or U15071 (N_15071,N_13891,N_13652);
xnor U15072 (N_15072,N_13617,N_13328);
nand U15073 (N_15073,N_14307,N_14087);
nand U15074 (N_15074,N_14068,N_13782);
nor U15075 (N_15075,N_13668,N_13624);
xnor U15076 (N_15076,N_13885,N_14155);
xnor U15077 (N_15077,N_13206,N_14391);
or U15078 (N_15078,N_13825,N_13979);
or U15079 (N_15079,N_13379,N_13539);
and U15080 (N_15080,N_13333,N_13708);
or U15081 (N_15081,N_14309,N_14299);
and U15082 (N_15082,N_13551,N_14110);
and U15083 (N_15083,N_13370,N_14081);
and U15084 (N_15084,N_13646,N_14126);
nand U15085 (N_15085,N_14371,N_13264);
nand U15086 (N_15086,N_14213,N_13853);
xor U15087 (N_15087,N_13870,N_13758);
nor U15088 (N_15088,N_13232,N_14141);
nand U15089 (N_15089,N_14126,N_13613);
and U15090 (N_15090,N_14394,N_14398);
nand U15091 (N_15091,N_13591,N_13831);
and U15092 (N_15092,N_13405,N_13719);
nor U15093 (N_15093,N_13390,N_13217);
nor U15094 (N_15094,N_13570,N_13544);
xnor U15095 (N_15095,N_14105,N_13978);
and U15096 (N_15096,N_13635,N_13454);
nor U15097 (N_15097,N_13993,N_13318);
nor U15098 (N_15098,N_13615,N_14370);
and U15099 (N_15099,N_13436,N_14218);
xor U15100 (N_15100,N_13702,N_13374);
nand U15101 (N_15101,N_14385,N_14227);
and U15102 (N_15102,N_13767,N_14025);
nand U15103 (N_15103,N_13580,N_13665);
nor U15104 (N_15104,N_13629,N_13807);
or U15105 (N_15105,N_13477,N_13975);
xor U15106 (N_15106,N_14077,N_13234);
nand U15107 (N_15107,N_14092,N_14266);
nor U15108 (N_15108,N_13411,N_14039);
xor U15109 (N_15109,N_14393,N_14103);
and U15110 (N_15110,N_13821,N_13595);
nand U15111 (N_15111,N_13238,N_14050);
and U15112 (N_15112,N_14090,N_13336);
nand U15113 (N_15113,N_14243,N_13264);
or U15114 (N_15114,N_13908,N_13962);
nand U15115 (N_15115,N_13751,N_13289);
nand U15116 (N_15116,N_13885,N_13479);
nand U15117 (N_15117,N_13277,N_14095);
or U15118 (N_15118,N_13651,N_13949);
or U15119 (N_15119,N_14220,N_13849);
nor U15120 (N_15120,N_14131,N_14388);
nand U15121 (N_15121,N_13566,N_13915);
nor U15122 (N_15122,N_14339,N_13926);
and U15123 (N_15123,N_14322,N_13405);
or U15124 (N_15124,N_14091,N_13474);
nand U15125 (N_15125,N_13669,N_14178);
or U15126 (N_15126,N_14205,N_13204);
nand U15127 (N_15127,N_13206,N_14091);
and U15128 (N_15128,N_13639,N_13814);
or U15129 (N_15129,N_14360,N_13916);
and U15130 (N_15130,N_13796,N_13232);
nor U15131 (N_15131,N_14370,N_14082);
xor U15132 (N_15132,N_13614,N_14034);
nor U15133 (N_15133,N_13742,N_13265);
and U15134 (N_15134,N_14310,N_13349);
nor U15135 (N_15135,N_13829,N_13852);
nor U15136 (N_15136,N_13385,N_14220);
xor U15137 (N_15137,N_13255,N_13989);
nand U15138 (N_15138,N_14131,N_13731);
nand U15139 (N_15139,N_13569,N_13488);
or U15140 (N_15140,N_13505,N_13335);
nor U15141 (N_15141,N_14288,N_13546);
nor U15142 (N_15142,N_13579,N_13646);
nor U15143 (N_15143,N_13495,N_13767);
or U15144 (N_15144,N_13812,N_13372);
or U15145 (N_15145,N_14274,N_13710);
and U15146 (N_15146,N_14022,N_14115);
and U15147 (N_15147,N_13211,N_13333);
xor U15148 (N_15148,N_13277,N_14215);
and U15149 (N_15149,N_13281,N_13479);
nor U15150 (N_15150,N_13542,N_13750);
xor U15151 (N_15151,N_14135,N_13633);
nor U15152 (N_15152,N_14184,N_13544);
and U15153 (N_15153,N_14288,N_14082);
or U15154 (N_15154,N_14225,N_14190);
xor U15155 (N_15155,N_13530,N_14085);
and U15156 (N_15156,N_13715,N_13357);
nand U15157 (N_15157,N_13639,N_14163);
and U15158 (N_15158,N_14096,N_13377);
and U15159 (N_15159,N_13338,N_14193);
and U15160 (N_15160,N_14072,N_13955);
nand U15161 (N_15161,N_14187,N_13230);
and U15162 (N_15162,N_14204,N_14366);
nor U15163 (N_15163,N_14396,N_14020);
nor U15164 (N_15164,N_13550,N_13513);
and U15165 (N_15165,N_13970,N_14339);
nand U15166 (N_15166,N_14333,N_13573);
nand U15167 (N_15167,N_14344,N_13320);
and U15168 (N_15168,N_13301,N_13325);
xnor U15169 (N_15169,N_14202,N_14274);
or U15170 (N_15170,N_13379,N_13788);
or U15171 (N_15171,N_14233,N_13975);
nand U15172 (N_15172,N_13684,N_13383);
xor U15173 (N_15173,N_13704,N_13237);
nand U15174 (N_15174,N_13857,N_13664);
and U15175 (N_15175,N_13467,N_13611);
xnor U15176 (N_15176,N_13389,N_13512);
nand U15177 (N_15177,N_13656,N_13470);
or U15178 (N_15178,N_13988,N_14280);
nand U15179 (N_15179,N_13640,N_13305);
xor U15180 (N_15180,N_13547,N_13377);
xnor U15181 (N_15181,N_14131,N_14374);
or U15182 (N_15182,N_13488,N_13704);
and U15183 (N_15183,N_14319,N_13318);
xor U15184 (N_15184,N_13974,N_13640);
nor U15185 (N_15185,N_14381,N_14103);
and U15186 (N_15186,N_13259,N_13590);
or U15187 (N_15187,N_13335,N_14041);
xor U15188 (N_15188,N_14180,N_13426);
and U15189 (N_15189,N_13638,N_14142);
nor U15190 (N_15190,N_13456,N_13775);
nor U15191 (N_15191,N_13525,N_13933);
nor U15192 (N_15192,N_13544,N_13677);
nor U15193 (N_15193,N_14285,N_13354);
nor U15194 (N_15194,N_13334,N_14354);
and U15195 (N_15195,N_13667,N_13558);
or U15196 (N_15196,N_13488,N_14193);
nor U15197 (N_15197,N_14207,N_13616);
xnor U15198 (N_15198,N_13338,N_14236);
and U15199 (N_15199,N_13350,N_13417);
and U15200 (N_15200,N_13656,N_13813);
or U15201 (N_15201,N_13926,N_14224);
and U15202 (N_15202,N_14231,N_13253);
xnor U15203 (N_15203,N_13649,N_14226);
nor U15204 (N_15204,N_13907,N_13244);
and U15205 (N_15205,N_13874,N_14161);
and U15206 (N_15206,N_13542,N_14284);
or U15207 (N_15207,N_13602,N_13374);
nor U15208 (N_15208,N_13441,N_13291);
or U15209 (N_15209,N_14241,N_13743);
nor U15210 (N_15210,N_14165,N_14100);
and U15211 (N_15211,N_13697,N_13253);
or U15212 (N_15212,N_14051,N_13357);
nand U15213 (N_15213,N_14017,N_14010);
nor U15214 (N_15214,N_13232,N_14150);
or U15215 (N_15215,N_13752,N_13202);
nor U15216 (N_15216,N_13617,N_13764);
xnor U15217 (N_15217,N_13574,N_13463);
and U15218 (N_15218,N_13967,N_14219);
nor U15219 (N_15219,N_13809,N_13276);
or U15220 (N_15220,N_13726,N_13962);
nor U15221 (N_15221,N_14010,N_13314);
and U15222 (N_15222,N_14210,N_13648);
xnor U15223 (N_15223,N_14317,N_14087);
xor U15224 (N_15224,N_14376,N_13660);
or U15225 (N_15225,N_13755,N_13619);
and U15226 (N_15226,N_14202,N_13655);
xnor U15227 (N_15227,N_13223,N_13928);
or U15228 (N_15228,N_13788,N_14144);
nand U15229 (N_15229,N_13326,N_13411);
and U15230 (N_15230,N_13219,N_14311);
or U15231 (N_15231,N_14100,N_13573);
and U15232 (N_15232,N_13813,N_14336);
xor U15233 (N_15233,N_13276,N_13474);
nor U15234 (N_15234,N_13297,N_13822);
or U15235 (N_15235,N_13744,N_13538);
or U15236 (N_15236,N_14185,N_13344);
nor U15237 (N_15237,N_13534,N_13779);
and U15238 (N_15238,N_13687,N_13916);
and U15239 (N_15239,N_14084,N_14034);
nor U15240 (N_15240,N_13485,N_13661);
and U15241 (N_15241,N_13714,N_13685);
xnor U15242 (N_15242,N_14315,N_14308);
nand U15243 (N_15243,N_14099,N_14350);
xnor U15244 (N_15244,N_13477,N_14243);
or U15245 (N_15245,N_13680,N_13393);
and U15246 (N_15246,N_14330,N_13761);
and U15247 (N_15247,N_14019,N_13387);
nor U15248 (N_15248,N_14282,N_14055);
or U15249 (N_15249,N_13438,N_14311);
or U15250 (N_15250,N_13937,N_14262);
xnor U15251 (N_15251,N_13884,N_13934);
nor U15252 (N_15252,N_13720,N_14257);
nor U15253 (N_15253,N_14336,N_14079);
and U15254 (N_15254,N_13677,N_13505);
nor U15255 (N_15255,N_13520,N_14225);
nand U15256 (N_15256,N_13942,N_14299);
nand U15257 (N_15257,N_13722,N_14074);
nand U15258 (N_15258,N_13609,N_14016);
nor U15259 (N_15259,N_13743,N_13482);
nand U15260 (N_15260,N_13800,N_13867);
nand U15261 (N_15261,N_14296,N_13860);
and U15262 (N_15262,N_13323,N_13902);
nor U15263 (N_15263,N_13581,N_13495);
xnor U15264 (N_15264,N_14180,N_13307);
nor U15265 (N_15265,N_13855,N_13201);
xor U15266 (N_15266,N_14178,N_13495);
nor U15267 (N_15267,N_13775,N_13906);
nor U15268 (N_15268,N_13345,N_13391);
nand U15269 (N_15269,N_13711,N_14171);
or U15270 (N_15270,N_13606,N_13856);
or U15271 (N_15271,N_14178,N_13277);
or U15272 (N_15272,N_13838,N_14278);
nand U15273 (N_15273,N_14341,N_13208);
nor U15274 (N_15274,N_13202,N_14159);
xor U15275 (N_15275,N_13324,N_14047);
and U15276 (N_15276,N_14198,N_13875);
nor U15277 (N_15277,N_14030,N_14298);
xnor U15278 (N_15278,N_13822,N_13688);
and U15279 (N_15279,N_14375,N_13597);
and U15280 (N_15280,N_14374,N_13282);
and U15281 (N_15281,N_14041,N_13464);
nor U15282 (N_15282,N_14120,N_14363);
nand U15283 (N_15283,N_13494,N_13554);
and U15284 (N_15284,N_13409,N_13942);
and U15285 (N_15285,N_13396,N_13471);
and U15286 (N_15286,N_13671,N_13772);
nor U15287 (N_15287,N_13587,N_13495);
xnor U15288 (N_15288,N_13570,N_13475);
and U15289 (N_15289,N_13569,N_13210);
nor U15290 (N_15290,N_13294,N_13270);
nand U15291 (N_15291,N_14223,N_13668);
or U15292 (N_15292,N_14182,N_13831);
or U15293 (N_15293,N_14372,N_13406);
xor U15294 (N_15294,N_13376,N_14150);
nand U15295 (N_15295,N_13573,N_13728);
nand U15296 (N_15296,N_13292,N_14108);
nand U15297 (N_15297,N_14317,N_14321);
nor U15298 (N_15298,N_14019,N_13980);
nand U15299 (N_15299,N_13213,N_14193);
or U15300 (N_15300,N_13352,N_13505);
nand U15301 (N_15301,N_13276,N_13773);
or U15302 (N_15302,N_13630,N_14309);
nand U15303 (N_15303,N_14240,N_13321);
or U15304 (N_15304,N_13323,N_13842);
nand U15305 (N_15305,N_13575,N_13618);
nand U15306 (N_15306,N_13285,N_13325);
or U15307 (N_15307,N_13202,N_13937);
and U15308 (N_15308,N_13821,N_14031);
xnor U15309 (N_15309,N_13658,N_13856);
xor U15310 (N_15310,N_14326,N_14020);
and U15311 (N_15311,N_14215,N_13644);
nor U15312 (N_15312,N_13211,N_13563);
nand U15313 (N_15313,N_14182,N_13879);
nor U15314 (N_15314,N_13690,N_13652);
nand U15315 (N_15315,N_13244,N_13839);
nor U15316 (N_15316,N_14372,N_13655);
nor U15317 (N_15317,N_14124,N_14010);
and U15318 (N_15318,N_13644,N_13637);
or U15319 (N_15319,N_14173,N_14084);
xnor U15320 (N_15320,N_13343,N_14142);
nor U15321 (N_15321,N_13564,N_14157);
nand U15322 (N_15322,N_14367,N_14240);
xnor U15323 (N_15323,N_13980,N_14302);
xnor U15324 (N_15324,N_13648,N_13833);
or U15325 (N_15325,N_13850,N_13686);
or U15326 (N_15326,N_13251,N_14320);
and U15327 (N_15327,N_13447,N_13483);
xor U15328 (N_15328,N_13791,N_13377);
nor U15329 (N_15329,N_13903,N_13423);
nand U15330 (N_15330,N_14001,N_13834);
xor U15331 (N_15331,N_13294,N_13306);
nand U15332 (N_15332,N_13909,N_13426);
and U15333 (N_15333,N_14082,N_13671);
xor U15334 (N_15334,N_13958,N_13563);
or U15335 (N_15335,N_13412,N_14192);
nand U15336 (N_15336,N_13350,N_13450);
and U15337 (N_15337,N_13999,N_14000);
nand U15338 (N_15338,N_14236,N_14132);
nand U15339 (N_15339,N_13956,N_13467);
nand U15340 (N_15340,N_13884,N_14343);
and U15341 (N_15341,N_14334,N_13300);
xnor U15342 (N_15342,N_13476,N_13552);
or U15343 (N_15343,N_13241,N_13808);
or U15344 (N_15344,N_13696,N_13903);
or U15345 (N_15345,N_13805,N_14085);
nor U15346 (N_15346,N_14387,N_13273);
or U15347 (N_15347,N_14247,N_13331);
or U15348 (N_15348,N_13926,N_14399);
and U15349 (N_15349,N_13937,N_13939);
xnor U15350 (N_15350,N_13443,N_13363);
nand U15351 (N_15351,N_14315,N_13707);
or U15352 (N_15352,N_14034,N_13258);
and U15353 (N_15353,N_14145,N_13268);
nor U15354 (N_15354,N_13553,N_13350);
nor U15355 (N_15355,N_13349,N_14094);
or U15356 (N_15356,N_14032,N_13905);
xnor U15357 (N_15357,N_13975,N_13430);
xor U15358 (N_15358,N_14073,N_14058);
xnor U15359 (N_15359,N_13721,N_13831);
and U15360 (N_15360,N_14273,N_13590);
nand U15361 (N_15361,N_13933,N_13602);
or U15362 (N_15362,N_13298,N_13774);
and U15363 (N_15363,N_14377,N_13723);
xnor U15364 (N_15364,N_13659,N_13365);
and U15365 (N_15365,N_13218,N_13227);
and U15366 (N_15366,N_13607,N_14351);
nand U15367 (N_15367,N_13360,N_13300);
and U15368 (N_15368,N_13882,N_14289);
nand U15369 (N_15369,N_14167,N_14351);
xor U15370 (N_15370,N_14259,N_14350);
nand U15371 (N_15371,N_13872,N_14248);
and U15372 (N_15372,N_13300,N_14228);
and U15373 (N_15373,N_14020,N_13843);
nor U15374 (N_15374,N_13828,N_13994);
xnor U15375 (N_15375,N_13383,N_14346);
nand U15376 (N_15376,N_13709,N_13364);
nor U15377 (N_15377,N_13913,N_14113);
nor U15378 (N_15378,N_13711,N_13569);
xnor U15379 (N_15379,N_13219,N_14102);
or U15380 (N_15380,N_13506,N_14205);
xnor U15381 (N_15381,N_13591,N_13740);
nand U15382 (N_15382,N_14269,N_13898);
or U15383 (N_15383,N_14380,N_13522);
or U15384 (N_15384,N_13744,N_14148);
or U15385 (N_15385,N_13821,N_13251);
nand U15386 (N_15386,N_13710,N_14153);
and U15387 (N_15387,N_13476,N_14129);
nor U15388 (N_15388,N_14158,N_13873);
nor U15389 (N_15389,N_13973,N_13777);
nand U15390 (N_15390,N_13390,N_14346);
and U15391 (N_15391,N_14361,N_13405);
and U15392 (N_15392,N_13923,N_13695);
nor U15393 (N_15393,N_13412,N_13974);
xor U15394 (N_15394,N_13804,N_14220);
nand U15395 (N_15395,N_14332,N_13915);
or U15396 (N_15396,N_13677,N_14213);
nor U15397 (N_15397,N_13580,N_13633);
nor U15398 (N_15398,N_14033,N_13268);
and U15399 (N_15399,N_14364,N_14285);
xor U15400 (N_15400,N_13657,N_13501);
nor U15401 (N_15401,N_14231,N_13832);
xnor U15402 (N_15402,N_13369,N_13766);
nand U15403 (N_15403,N_14212,N_14318);
and U15404 (N_15404,N_13499,N_14360);
or U15405 (N_15405,N_13314,N_13496);
and U15406 (N_15406,N_13495,N_13728);
nand U15407 (N_15407,N_13430,N_13223);
nor U15408 (N_15408,N_13553,N_13597);
xor U15409 (N_15409,N_13802,N_14330);
nand U15410 (N_15410,N_13352,N_14349);
or U15411 (N_15411,N_13529,N_13342);
or U15412 (N_15412,N_13219,N_13282);
nand U15413 (N_15413,N_14073,N_14239);
xnor U15414 (N_15414,N_14289,N_13825);
or U15415 (N_15415,N_13682,N_14001);
nor U15416 (N_15416,N_13615,N_13756);
nand U15417 (N_15417,N_13567,N_14336);
nor U15418 (N_15418,N_13989,N_14034);
nor U15419 (N_15419,N_13853,N_13777);
or U15420 (N_15420,N_13709,N_13660);
or U15421 (N_15421,N_13839,N_13635);
nor U15422 (N_15422,N_14187,N_13839);
nand U15423 (N_15423,N_13994,N_13216);
xor U15424 (N_15424,N_13934,N_14293);
xnor U15425 (N_15425,N_13318,N_14040);
nor U15426 (N_15426,N_13987,N_14260);
nor U15427 (N_15427,N_14396,N_13624);
nand U15428 (N_15428,N_13309,N_13546);
and U15429 (N_15429,N_14240,N_13958);
or U15430 (N_15430,N_13461,N_13425);
nor U15431 (N_15431,N_13538,N_14077);
and U15432 (N_15432,N_13250,N_13997);
nand U15433 (N_15433,N_13305,N_13925);
xor U15434 (N_15434,N_13774,N_13537);
nand U15435 (N_15435,N_13672,N_14393);
nor U15436 (N_15436,N_13621,N_13415);
and U15437 (N_15437,N_14335,N_13605);
nor U15438 (N_15438,N_13411,N_13827);
nor U15439 (N_15439,N_14102,N_13476);
or U15440 (N_15440,N_14392,N_14244);
nand U15441 (N_15441,N_13303,N_13272);
and U15442 (N_15442,N_13679,N_13574);
xnor U15443 (N_15443,N_13808,N_13314);
nor U15444 (N_15444,N_13244,N_14167);
and U15445 (N_15445,N_14180,N_13522);
nand U15446 (N_15446,N_13348,N_13589);
nor U15447 (N_15447,N_13561,N_14324);
and U15448 (N_15448,N_13917,N_14036);
or U15449 (N_15449,N_13401,N_13365);
nor U15450 (N_15450,N_14391,N_13580);
and U15451 (N_15451,N_13426,N_13268);
xor U15452 (N_15452,N_14058,N_13338);
and U15453 (N_15453,N_13917,N_13968);
nand U15454 (N_15454,N_13231,N_13713);
nand U15455 (N_15455,N_13374,N_13470);
nor U15456 (N_15456,N_14080,N_14372);
nand U15457 (N_15457,N_14370,N_13632);
nand U15458 (N_15458,N_14043,N_13628);
or U15459 (N_15459,N_13592,N_14190);
xnor U15460 (N_15460,N_14074,N_14305);
xor U15461 (N_15461,N_13978,N_13800);
or U15462 (N_15462,N_13861,N_14284);
nor U15463 (N_15463,N_13540,N_13848);
nand U15464 (N_15464,N_14027,N_14380);
and U15465 (N_15465,N_13615,N_14126);
or U15466 (N_15466,N_13688,N_13280);
xnor U15467 (N_15467,N_13854,N_14030);
or U15468 (N_15468,N_13553,N_14139);
nand U15469 (N_15469,N_14180,N_13958);
and U15470 (N_15470,N_13753,N_14036);
nor U15471 (N_15471,N_13676,N_13960);
nand U15472 (N_15472,N_14025,N_13645);
or U15473 (N_15473,N_14376,N_13236);
and U15474 (N_15474,N_14065,N_13385);
or U15475 (N_15475,N_14370,N_13603);
nand U15476 (N_15476,N_14138,N_13854);
and U15477 (N_15477,N_13470,N_13295);
or U15478 (N_15478,N_14170,N_14101);
and U15479 (N_15479,N_13900,N_14361);
xnor U15480 (N_15480,N_14066,N_13817);
xnor U15481 (N_15481,N_14199,N_13341);
nand U15482 (N_15482,N_13223,N_13361);
nand U15483 (N_15483,N_13930,N_14339);
nand U15484 (N_15484,N_14158,N_13707);
nand U15485 (N_15485,N_14390,N_13592);
xor U15486 (N_15486,N_14233,N_13885);
and U15487 (N_15487,N_14023,N_13956);
xnor U15488 (N_15488,N_14150,N_13762);
nor U15489 (N_15489,N_13649,N_13886);
and U15490 (N_15490,N_13237,N_13402);
nor U15491 (N_15491,N_13692,N_14301);
or U15492 (N_15492,N_13374,N_13690);
or U15493 (N_15493,N_13695,N_13953);
xnor U15494 (N_15494,N_13720,N_13511);
nand U15495 (N_15495,N_13761,N_14247);
or U15496 (N_15496,N_14028,N_13620);
or U15497 (N_15497,N_13211,N_13548);
and U15498 (N_15498,N_13711,N_13698);
or U15499 (N_15499,N_14333,N_14043);
or U15500 (N_15500,N_13287,N_13378);
nand U15501 (N_15501,N_13488,N_13584);
nor U15502 (N_15502,N_13572,N_14179);
and U15503 (N_15503,N_13541,N_13523);
nor U15504 (N_15504,N_14307,N_13754);
nor U15505 (N_15505,N_14084,N_13480);
xor U15506 (N_15506,N_13420,N_13397);
and U15507 (N_15507,N_14056,N_13266);
and U15508 (N_15508,N_13969,N_13723);
nor U15509 (N_15509,N_13235,N_14194);
xor U15510 (N_15510,N_14385,N_13589);
xor U15511 (N_15511,N_13276,N_13686);
nor U15512 (N_15512,N_14343,N_13943);
and U15513 (N_15513,N_13475,N_13806);
xnor U15514 (N_15514,N_14038,N_13263);
or U15515 (N_15515,N_13575,N_14007);
xor U15516 (N_15516,N_13224,N_14153);
or U15517 (N_15517,N_13950,N_14036);
nand U15518 (N_15518,N_13699,N_14277);
nand U15519 (N_15519,N_13461,N_14088);
or U15520 (N_15520,N_13657,N_13255);
xnor U15521 (N_15521,N_14151,N_13941);
or U15522 (N_15522,N_13791,N_13721);
or U15523 (N_15523,N_13550,N_14200);
or U15524 (N_15524,N_13404,N_14226);
and U15525 (N_15525,N_13828,N_14038);
nor U15526 (N_15526,N_13474,N_13212);
or U15527 (N_15527,N_13291,N_13206);
xnor U15528 (N_15528,N_13891,N_13819);
nand U15529 (N_15529,N_14265,N_14310);
nand U15530 (N_15530,N_13877,N_14164);
xor U15531 (N_15531,N_13662,N_13885);
nor U15532 (N_15532,N_13939,N_13859);
or U15533 (N_15533,N_13477,N_13212);
xnor U15534 (N_15534,N_14123,N_14301);
nand U15535 (N_15535,N_14193,N_14229);
and U15536 (N_15536,N_13628,N_13432);
nor U15537 (N_15537,N_13615,N_13940);
xor U15538 (N_15538,N_13947,N_13629);
nor U15539 (N_15539,N_14104,N_14378);
nor U15540 (N_15540,N_13861,N_13680);
nor U15541 (N_15541,N_13997,N_14385);
nor U15542 (N_15542,N_13612,N_13699);
nor U15543 (N_15543,N_13902,N_14017);
xor U15544 (N_15544,N_13426,N_13557);
nand U15545 (N_15545,N_13952,N_13685);
nand U15546 (N_15546,N_13748,N_13534);
or U15547 (N_15547,N_14158,N_13994);
or U15548 (N_15548,N_14182,N_13653);
nor U15549 (N_15549,N_14099,N_13208);
xnor U15550 (N_15550,N_13905,N_13257);
xnor U15551 (N_15551,N_13927,N_13325);
or U15552 (N_15552,N_13938,N_14169);
and U15553 (N_15553,N_13520,N_14322);
or U15554 (N_15554,N_13856,N_13666);
or U15555 (N_15555,N_14337,N_13740);
nor U15556 (N_15556,N_14039,N_13303);
and U15557 (N_15557,N_14388,N_13759);
nor U15558 (N_15558,N_13272,N_14238);
and U15559 (N_15559,N_13553,N_13816);
nand U15560 (N_15560,N_13777,N_13228);
and U15561 (N_15561,N_14005,N_13308);
and U15562 (N_15562,N_13716,N_14384);
nor U15563 (N_15563,N_13206,N_13213);
xnor U15564 (N_15564,N_14139,N_14026);
xnor U15565 (N_15565,N_13567,N_13684);
and U15566 (N_15566,N_13419,N_13462);
or U15567 (N_15567,N_13871,N_14205);
and U15568 (N_15568,N_13909,N_13420);
nand U15569 (N_15569,N_14151,N_14093);
and U15570 (N_15570,N_13254,N_13204);
and U15571 (N_15571,N_14319,N_13607);
xnor U15572 (N_15572,N_13788,N_13321);
nor U15573 (N_15573,N_14346,N_14199);
or U15574 (N_15574,N_13779,N_14154);
and U15575 (N_15575,N_13903,N_13393);
xnor U15576 (N_15576,N_14298,N_14025);
or U15577 (N_15577,N_14325,N_13435);
and U15578 (N_15578,N_14312,N_13486);
nand U15579 (N_15579,N_14029,N_14119);
or U15580 (N_15580,N_13352,N_13296);
xnor U15581 (N_15581,N_13558,N_13393);
or U15582 (N_15582,N_13291,N_13543);
or U15583 (N_15583,N_13309,N_14358);
xor U15584 (N_15584,N_14368,N_13915);
nor U15585 (N_15585,N_13839,N_13319);
or U15586 (N_15586,N_13879,N_14322);
or U15587 (N_15587,N_13871,N_13529);
nand U15588 (N_15588,N_13277,N_14266);
nand U15589 (N_15589,N_14317,N_14139);
xnor U15590 (N_15590,N_14036,N_13356);
or U15591 (N_15591,N_14375,N_14399);
nand U15592 (N_15592,N_13528,N_14304);
xnor U15593 (N_15593,N_14121,N_14185);
or U15594 (N_15594,N_14332,N_13293);
nor U15595 (N_15595,N_13613,N_13714);
xor U15596 (N_15596,N_13579,N_13709);
nand U15597 (N_15597,N_13973,N_13289);
or U15598 (N_15598,N_13475,N_13239);
xor U15599 (N_15599,N_14236,N_14201);
xor U15600 (N_15600,N_15282,N_14814);
xnor U15601 (N_15601,N_15104,N_14674);
xor U15602 (N_15602,N_15048,N_14872);
xnor U15603 (N_15603,N_15483,N_15235);
and U15604 (N_15604,N_14542,N_14488);
nor U15605 (N_15605,N_15592,N_15301);
or U15606 (N_15606,N_14682,N_15459);
and U15607 (N_15607,N_14708,N_14857);
or U15608 (N_15608,N_14628,N_15144);
nand U15609 (N_15609,N_14519,N_14873);
nor U15610 (N_15610,N_14869,N_15234);
or U15611 (N_15611,N_15380,N_15574);
or U15612 (N_15612,N_14851,N_15310);
or U15613 (N_15613,N_14957,N_15154);
xnor U15614 (N_15614,N_15428,N_14701);
and U15615 (N_15615,N_15449,N_15315);
nor U15616 (N_15616,N_15458,N_15180);
xnor U15617 (N_15617,N_14409,N_14978);
and U15618 (N_15618,N_15441,N_15107);
xor U15619 (N_15619,N_14921,N_15448);
nand U15620 (N_15620,N_15488,N_14992);
nor U15621 (N_15621,N_14412,N_14579);
or U15622 (N_15622,N_14877,N_15462);
or U15623 (N_15623,N_14833,N_14989);
nor U15624 (N_15624,N_15548,N_14463);
nand U15625 (N_15625,N_14681,N_14726);
xor U15626 (N_15626,N_14443,N_15078);
or U15627 (N_15627,N_14467,N_15581);
nor U15628 (N_15628,N_14808,N_15351);
nor U15629 (N_15629,N_14754,N_15011);
and U15630 (N_15630,N_15464,N_14604);
and U15631 (N_15631,N_15190,N_14440);
xnor U15632 (N_15632,N_14817,N_14920);
xor U15633 (N_15633,N_15576,N_15418);
or U15634 (N_15634,N_15225,N_15049);
or U15635 (N_15635,N_15314,N_14600);
nor U15636 (N_15636,N_14632,N_15500);
nor U15637 (N_15637,N_15421,N_15480);
nor U15638 (N_15638,N_15504,N_15528);
nor U15639 (N_15639,N_15260,N_15207);
nor U15640 (N_15640,N_14786,N_15281);
or U15641 (N_15641,N_14820,N_14635);
nor U15642 (N_15642,N_15187,N_15128);
and U15643 (N_15643,N_14479,N_15465);
nand U15644 (N_15644,N_14717,N_14909);
xnor U15645 (N_15645,N_15105,N_15439);
nand U15646 (N_15646,N_14575,N_14780);
xnor U15647 (N_15647,N_15437,N_15212);
or U15648 (N_15648,N_14751,N_15403);
xor U15649 (N_15649,N_15531,N_15346);
and U15650 (N_15650,N_15491,N_14511);
xnor U15651 (N_15651,N_15111,N_14993);
and U15652 (N_15652,N_14777,N_14637);
nand U15653 (N_15653,N_15426,N_14973);
and U15654 (N_15654,N_14522,N_14969);
nor U15655 (N_15655,N_14531,N_15097);
nor U15656 (N_15656,N_15295,N_14465);
and U15657 (N_15657,N_14854,N_15200);
and U15658 (N_15658,N_14775,N_14796);
xor U15659 (N_15659,N_14594,N_15161);
nor U15660 (N_15660,N_15397,N_14764);
and U15661 (N_15661,N_14549,N_14995);
nor U15662 (N_15662,N_15412,N_14602);
or U15663 (N_15663,N_14415,N_14406);
and U15664 (N_15664,N_15422,N_14578);
nor U15665 (N_15665,N_14444,N_14848);
xor U15666 (N_15666,N_14580,N_14929);
or U15667 (N_15667,N_14893,N_15575);
or U15668 (N_15668,N_15184,N_14642);
nor U15669 (N_15669,N_15517,N_14928);
or U15670 (N_15670,N_14662,N_15408);
and U15671 (N_15671,N_15329,N_14474);
or U15672 (N_15672,N_14477,N_15194);
and U15673 (N_15673,N_15446,N_15123);
nand U15674 (N_15674,N_14844,N_14539);
xnor U15675 (N_15675,N_15168,N_15062);
nor U15676 (N_15676,N_14723,N_14693);
and U15677 (N_15677,N_14952,N_14791);
xor U15678 (N_15678,N_14900,N_15580);
and U15679 (N_15679,N_14449,N_14582);
nor U15680 (N_15680,N_15519,N_14798);
xnor U15681 (N_15681,N_14448,N_14459);
nor U15682 (N_15682,N_14789,N_14876);
and U15683 (N_15683,N_15126,N_15246);
or U15684 (N_15684,N_15125,N_14910);
xnor U15685 (N_15685,N_15475,N_14736);
or U15686 (N_15686,N_15599,N_15502);
nor U15687 (N_15687,N_14475,N_14932);
nor U15688 (N_15688,N_15169,N_14901);
or U15689 (N_15689,N_15455,N_15223);
nand U15690 (N_15690,N_14953,N_15457);
or U15691 (N_15691,N_14863,N_14613);
or U15692 (N_15692,N_14783,N_14428);
nand U15693 (N_15693,N_14499,N_14585);
and U15694 (N_15694,N_14512,N_14664);
xnor U15695 (N_15695,N_15537,N_14945);
xnor U15696 (N_15696,N_14566,N_15362);
nor U15697 (N_15697,N_15101,N_14842);
nand U15698 (N_15698,N_15036,N_15151);
nand U15699 (N_15699,N_15160,N_15514);
nand U15700 (N_15700,N_15086,N_15170);
or U15701 (N_15701,N_15066,N_15538);
nor U15702 (N_15702,N_15313,N_15092);
nand U15703 (N_15703,N_14420,N_15023);
nor U15704 (N_15704,N_15269,N_14748);
and U15705 (N_15705,N_14405,N_14562);
or U15706 (N_15706,N_14418,N_14698);
or U15707 (N_15707,N_14419,N_14556);
nand U15708 (N_15708,N_15479,N_14981);
or U15709 (N_15709,N_14554,N_14934);
xnor U15710 (N_15710,N_14725,N_15245);
nor U15711 (N_15711,N_14828,N_14907);
or U15712 (N_15712,N_15179,N_15192);
nor U15713 (N_15713,N_15469,N_14410);
nand U15714 (N_15714,N_15454,N_15134);
nand U15715 (N_15715,N_14906,N_14912);
or U15716 (N_15716,N_15486,N_15567);
and U15717 (N_15717,N_14850,N_14926);
and U15718 (N_15718,N_15198,N_14862);
or U15719 (N_15719,N_14899,N_14716);
xor U15720 (N_15720,N_15414,N_14644);
and U15721 (N_15721,N_15091,N_15142);
or U15722 (N_15722,N_14913,N_15132);
nor U15723 (N_15723,N_14773,N_14584);
xnor U15724 (N_15724,N_15562,N_15213);
xnor U15725 (N_15725,N_14871,N_14441);
xnor U15726 (N_15726,N_15396,N_14818);
and U15727 (N_15727,N_15555,N_14831);
and U15728 (N_15728,N_15098,N_14771);
nor U15729 (N_15729,N_15355,N_14822);
and U15730 (N_15730,N_15415,N_15423);
nor U15731 (N_15731,N_15365,N_14675);
nor U15732 (N_15732,N_15229,N_14506);
nand U15733 (N_15733,N_14691,N_14638);
nand U15734 (N_15734,N_15432,N_14655);
nor U15735 (N_15735,N_15472,N_15335);
nor U15736 (N_15736,N_14983,N_15337);
or U15737 (N_15737,N_14744,N_15109);
and U15738 (N_15738,N_15560,N_14571);
nand U15739 (N_15739,N_14927,N_14841);
xnor U15740 (N_15740,N_15197,N_15326);
or U15741 (N_15741,N_15589,N_14625);
nand U15742 (N_15742,N_14446,N_15591);
nand U15743 (N_15743,N_15383,N_15040);
and U15744 (N_15744,N_14572,N_14533);
nor U15745 (N_15745,N_15309,N_15585);
nor U15746 (N_15746,N_15060,N_14843);
xor U15747 (N_15747,N_14936,N_14507);
xor U15748 (N_15748,N_15178,N_14481);
nand U15749 (N_15749,N_14498,N_15435);
nand U15750 (N_15750,N_14733,N_15113);
nor U15751 (N_15751,N_15006,N_14942);
nor U15752 (N_15752,N_15220,N_15541);
nand U15753 (N_15753,N_15453,N_15022);
nor U15754 (N_15754,N_14879,N_14940);
and U15755 (N_15755,N_15378,N_14917);
or U15756 (N_15756,N_15595,N_14776);
nand U15757 (N_15757,N_15185,N_14669);
and U15758 (N_15758,N_15390,N_15028);
nand U15759 (N_15759,N_15577,N_15413);
xnor U15760 (N_15760,N_15262,N_14422);
and U15761 (N_15761,N_14944,N_14960);
or U15762 (N_15762,N_15094,N_15565);
xnor U15763 (N_15763,N_14532,N_15367);
nand U15764 (N_15764,N_15119,N_15004);
xor U15765 (N_15765,N_14670,N_14971);
and U15766 (N_15766,N_15391,N_15143);
xnor U15767 (N_15767,N_15039,N_14659);
nor U15768 (N_15768,N_15416,N_14830);
and U15769 (N_15769,N_15171,N_15348);
or U15770 (N_15770,N_15073,N_14557);
nand U15771 (N_15771,N_14816,N_15230);
or U15772 (N_15772,N_14961,N_15007);
xor U15773 (N_15773,N_15138,N_14977);
nor U15774 (N_15774,N_15024,N_14486);
or U15775 (N_15775,N_15047,N_14483);
nor U15776 (N_15776,N_14437,N_14429);
nor U15777 (N_15777,N_14541,N_14704);
or U15778 (N_15778,N_15382,N_15117);
nand U15779 (N_15779,N_15196,N_14517);
nor U15780 (N_15780,N_15015,N_14760);
or U15781 (N_15781,N_15553,N_14643);
and U15782 (N_15782,N_14634,N_14787);
and U15783 (N_15783,N_15300,N_15546);
nand U15784 (N_15784,N_15545,N_15405);
or U15785 (N_15785,N_14985,N_14782);
nor U15786 (N_15786,N_14502,N_14658);
xnor U15787 (N_15787,N_14892,N_14938);
or U15788 (N_15788,N_14724,N_15122);
and U15789 (N_15789,N_15100,N_14838);
nor U15790 (N_15790,N_15343,N_14561);
or U15791 (N_15791,N_15487,N_14809);
or U15792 (N_15792,N_15000,N_14414);
nor U15793 (N_15793,N_15236,N_14812);
or U15794 (N_15794,N_15505,N_14472);
or U15795 (N_15795,N_15195,N_15532);
xor U15796 (N_15796,N_15241,N_15191);
nand U15797 (N_15797,N_15108,N_14813);
xnor U15798 (N_15798,N_15189,N_14805);
and U15799 (N_15799,N_15571,N_15593);
nand U15800 (N_15800,N_14515,N_15496);
nand U15801 (N_15801,N_15008,N_15360);
and U15802 (N_15802,N_15076,N_15278);
xor U15803 (N_15803,N_15003,N_14930);
xor U15804 (N_15804,N_14593,N_15244);
xnor U15805 (N_15805,N_15019,N_15254);
xnor U15806 (N_15806,N_15419,N_14874);
and U15807 (N_15807,N_14622,N_14469);
nor U15808 (N_15808,N_14962,N_15510);
nand U15809 (N_15809,N_15276,N_15485);
nor U15810 (N_15810,N_15385,N_15042);
nor U15811 (N_15811,N_14417,N_15050);
and U15812 (N_15812,N_15087,N_15334);
nand U15813 (N_15813,N_15588,N_15120);
nand U15814 (N_15814,N_15218,N_15037);
xnor U15815 (N_15815,N_15165,N_14870);
or U15816 (N_15816,N_14702,N_14774);
and U15817 (N_15817,N_14987,N_14866);
or U15818 (N_15818,N_14645,N_14599);
xor U15819 (N_15819,N_14480,N_14972);
or U15820 (N_15820,N_14997,N_15251);
xor U15821 (N_15821,N_14721,N_15158);
xor U15822 (N_15822,N_14490,N_15102);
xnor U15823 (N_15823,N_15359,N_15096);
or U15824 (N_15824,N_14804,N_14553);
nor U15825 (N_15825,N_15299,N_15427);
nand U15826 (N_15826,N_15221,N_15085);
nor U15827 (N_15827,N_15172,N_14758);
xor U15828 (N_15828,N_15393,N_14759);
xor U15829 (N_15829,N_14471,N_15384);
nor U15830 (N_15830,N_14657,N_15539);
xnor U15831 (N_15831,N_14954,N_15074);
xnor U15832 (N_15832,N_15399,N_15075);
xor U15833 (N_15833,N_15392,N_15162);
and U15834 (N_15834,N_15228,N_14445);
nor U15835 (N_15835,N_15358,N_14948);
nor U15836 (N_15836,N_15084,N_15253);
xor U15837 (N_15837,N_14476,N_15470);
nand U15838 (N_15838,N_14891,N_15507);
xnor U15839 (N_15839,N_15090,N_14695);
xor U15840 (N_15840,N_15202,N_14767);
nand U15841 (N_15841,N_15381,N_15305);
xnor U15842 (N_15842,N_14516,N_14668);
nor U15843 (N_15843,N_14705,N_14685);
and U15844 (N_15844,N_15494,N_14886);
nand U15845 (N_15845,N_15492,N_15280);
and U15846 (N_15846,N_14826,N_14959);
or U15847 (N_15847,N_15072,N_15148);
nor U15848 (N_15848,N_14807,N_15330);
and U15849 (N_15849,N_15400,N_14795);
or U15850 (N_15850,N_14588,N_14661);
xor U15851 (N_15851,N_14464,N_15534);
nand U15852 (N_15852,N_15316,N_14425);
and U15853 (N_15853,N_14855,N_14606);
and U15854 (N_15854,N_14407,N_15174);
and U15855 (N_15855,N_15298,N_14860);
nand U15856 (N_15856,N_15093,N_15018);
nor U15857 (N_15857,N_15121,N_14457);
nand U15858 (N_15858,N_15516,N_14679);
or U15859 (N_15859,N_15156,N_15157);
nand U15860 (N_15860,N_15069,N_15175);
nand U15861 (N_15861,N_15478,N_14895);
nand U15862 (N_15862,N_15127,N_14530);
xor U15863 (N_15863,N_14694,N_15318);
and U15864 (N_15864,N_15193,N_15252);
and U15865 (N_15865,N_14750,N_15594);
xor U15866 (N_15866,N_15058,N_15079);
or U15867 (N_15867,N_14727,N_15370);
xnor U15868 (N_15868,N_15530,N_15371);
nand U15869 (N_15869,N_15533,N_15064);
or U15870 (N_15870,N_14458,N_14713);
and U15871 (N_15871,N_14646,N_14770);
nor U15872 (N_15872,N_14496,N_14801);
and U15873 (N_15873,N_14856,N_15250);
xnor U15874 (N_15874,N_15511,N_14683);
xor U15875 (N_15875,N_14460,N_15369);
nor U15876 (N_15876,N_14666,N_14741);
xnor U15877 (N_15877,N_14603,N_14663);
and U15878 (N_15878,N_14896,N_14528);
nor U15879 (N_15879,N_14621,N_14875);
or U15880 (N_15880,N_14489,N_15286);
or U15881 (N_15881,N_15590,N_15354);
or U15882 (N_15882,N_14615,N_14840);
and U15883 (N_15883,N_14933,N_15095);
nand U15884 (N_15884,N_15082,N_14686);
nand U15885 (N_15885,N_15292,N_14494);
nand U15886 (N_15886,N_15474,N_15340);
and U15887 (N_15887,N_15044,N_15032);
xor U15888 (N_15888,N_15341,N_15131);
and U15889 (N_15889,N_15319,N_14688);
nor U15890 (N_15890,N_14797,N_15304);
and U15891 (N_15891,N_14649,N_14802);
or U15892 (N_15892,N_15338,N_14610);
xnor U15893 (N_15893,N_15322,N_15002);
and U15894 (N_15894,N_15248,N_15523);
xnor U15895 (N_15895,N_15243,N_14509);
nor U15896 (N_15896,N_14853,N_15265);
and U15897 (N_15897,N_14624,N_14641);
and U15898 (N_15898,N_14423,N_14715);
nand U15899 (N_15899,N_15249,N_14676);
or U15900 (N_15900,N_15268,N_15339);
nor U15901 (N_15901,N_15434,N_15274);
nor U15902 (N_15902,N_14990,N_15201);
or U15903 (N_15903,N_15140,N_15543);
xnor U15904 (N_15904,N_14763,N_14629);
nor U15905 (N_15905,N_14803,N_14501);
nand U15906 (N_15906,N_14825,N_14894);
and U15907 (N_15907,N_14925,N_14521);
and U15908 (N_15908,N_15137,N_14970);
nand U15909 (N_15909,N_15311,N_15556);
nor U15910 (N_15910,N_15345,N_14966);
or U15911 (N_15911,N_14689,N_15145);
xnor U15912 (N_15912,N_15052,N_14881);
and U15913 (N_15913,N_15374,N_15264);
nor U15914 (N_15914,N_15325,N_14651);
or U15915 (N_15915,N_14815,N_15386);
nand U15916 (N_15916,N_14432,N_15153);
nor U15917 (N_15917,N_14518,N_15509);
or U15918 (N_15918,N_14994,N_15372);
xnor U15919 (N_15919,N_14495,N_15493);
nand U15920 (N_15920,N_14707,N_14508);
nor U15921 (N_15921,N_14746,N_14887);
and U15922 (N_15922,N_15363,N_15027);
nor U15923 (N_15923,N_14627,N_14793);
and U15924 (N_15924,N_15222,N_14618);
and U15925 (N_15925,N_14762,N_15130);
and U15926 (N_15926,N_14535,N_15373);
nor U15927 (N_15927,N_15321,N_14678);
xnor U15928 (N_15928,N_15526,N_15293);
and U15929 (N_15929,N_15217,N_15081);
nand U15930 (N_15930,N_14982,N_15557);
or U15931 (N_15931,N_14967,N_15336);
nand U15932 (N_15932,N_14740,N_15320);
and U15933 (N_15933,N_15489,N_14570);
and U15934 (N_15934,N_14607,N_14491);
nand U15935 (N_15935,N_14598,N_14577);
or U15936 (N_15936,N_14609,N_14950);
and U15937 (N_15937,N_14447,N_14546);
and U15938 (N_15938,N_14847,N_14520);
xor U15939 (N_15939,N_15349,N_15468);
or U15940 (N_15940,N_14747,N_14485);
and U15941 (N_15941,N_14772,N_14623);
xor U15942 (N_15942,N_14540,N_14536);
or U15943 (N_15943,N_14996,N_15368);
nor U15944 (N_15944,N_15508,N_14473);
nor U15945 (N_15945,N_14845,N_15561);
or U15946 (N_15946,N_15513,N_14742);
nand U15947 (N_15947,N_14720,N_15233);
or U15948 (N_15948,N_14563,N_15477);
or U15949 (N_15949,N_15598,N_14964);
nor U15950 (N_15950,N_14810,N_14792);
or U15951 (N_15951,N_14849,N_15306);
xor U15952 (N_15952,N_15518,N_14728);
and U15953 (N_15953,N_15041,N_15570);
nor U15954 (N_15954,N_14956,N_14461);
or U15955 (N_15955,N_14431,N_15021);
and U15956 (N_15956,N_15498,N_14769);
nand U15957 (N_15957,N_14980,N_14790);
xor U15958 (N_15958,N_15232,N_15499);
nand U15959 (N_15959,N_15552,N_14550);
and U15960 (N_15960,N_15331,N_15307);
or U15961 (N_15961,N_15110,N_15159);
xor U15962 (N_15962,N_15389,N_14665);
and U15963 (N_15963,N_15017,N_14650);
xnor U15964 (N_15964,N_14731,N_14527);
nand U15965 (N_15965,N_14633,N_14951);
nand U15966 (N_15966,N_15379,N_15255);
nand U15967 (N_15967,N_14587,N_15226);
or U15968 (N_15968,N_15106,N_15182);
or U15969 (N_15969,N_15398,N_14424);
and U15970 (N_15970,N_15114,N_14558);
nand U15971 (N_15971,N_15256,N_15317);
nor U15972 (N_15972,N_15308,N_15332);
xor U15973 (N_15973,N_14779,N_15551);
and U15974 (N_15974,N_14573,N_14735);
xor U15975 (N_15975,N_14614,N_15167);
nand U15976 (N_15976,N_15054,N_14974);
or U15977 (N_15977,N_14478,N_15239);
nor U15978 (N_15978,N_15214,N_15088);
and U15979 (N_15979,N_15536,N_15558);
and U15980 (N_15980,N_14719,N_14697);
nor U15981 (N_15981,N_14756,N_14703);
nand U15982 (N_15982,N_14411,N_15290);
nand U15983 (N_15983,N_14710,N_14864);
xor U15984 (N_15984,N_15521,N_15524);
nand U15985 (N_15985,N_14543,N_15053);
nand U15986 (N_15986,N_15442,N_14470);
nor U15987 (N_15987,N_15067,N_14616);
nand U15988 (N_15988,N_15240,N_15387);
nand U15989 (N_15989,N_14636,N_15020);
nand U15990 (N_15990,N_15296,N_14656);
nor U15991 (N_15991,N_14597,N_15231);
and U15992 (N_15992,N_14560,N_14700);
and U15993 (N_15993,N_15559,N_14529);
or U15994 (N_15994,N_15279,N_14867);
nor U15995 (N_15995,N_14421,N_14824);
nor U15996 (N_15996,N_15471,N_15238);
nand U15997 (N_15997,N_15080,N_15569);
or U15998 (N_15998,N_14452,N_15447);
nor U15999 (N_15999,N_14868,N_14439);
or U16000 (N_16000,N_14505,N_14538);
nand U16001 (N_16001,N_14592,N_15150);
nand U16002 (N_16002,N_14880,N_15204);
and U16003 (N_16003,N_14684,N_14890);
and U16004 (N_16004,N_14821,N_15476);
and U16005 (N_16005,N_15544,N_15512);
or U16006 (N_16006,N_14898,N_15582);
xnor U16007 (N_16007,N_15267,N_15327);
nor U16008 (N_16008,N_15436,N_15164);
and U16009 (N_16009,N_15323,N_15404);
or U16010 (N_16010,N_15055,N_14513);
nor U16011 (N_16011,N_14548,N_15342);
nor U16012 (N_16012,N_15014,N_15025);
nand U16013 (N_16013,N_14564,N_14914);
nor U16014 (N_16014,N_14752,N_15409);
nand U16015 (N_16015,N_15501,N_14976);
xor U16016 (N_16016,N_14800,N_15010);
nor U16017 (N_16017,N_14749,N_15333);
or U16018 (N_16018,N_14537,N_15535);
and U16019 (N_16019,N_14545,N_14626);
nand U16020 (N_16020,N_15353,N_15433);
or U16021 (N_16021,N_15438,N_14630);
nand U16022 (N_16022,N_15467,N_14468);
xnor U16023 (N_16023,N_15350,N_14569);
nor U16024 (N_16024,N_14839,N_14504);
or U16025 (N_16025,N_15057,N_14552);
xor U16026 (N_16026,N_14619,N_15257);
nand U16027 (N_16027,N_14743,N_15112);
nor U16028 (N_16028,N_14908,N_14555);
and U16029 (N_16029,N_14963,N_14781);
and U16030 (N_16030,N_15473,N_15139);
nand U16031 (N_16031,N_14837,N_15155);
nor U16032 (N_16032,N_14836,N_14450);
nor U16033 (N_16033,N_15579,N_15583);
and U16034 (N_16034,N_15012,N_15445);
nand U16035 (N_16035,N_14524,N_15456);
xnor U16036 (N_16036,N_15034,N_14559);
nor U16037 (N_16037,N_15401,N_15026);
nand U16038 (N_16038,N_14631,N_14732);
and U16039 (N_16039,N_15407,N_14918);
and U16040 (N_16040,N_14433,N_15273);
and U16041 (N_16041,N_15206,N_15277);
or U16042 (N_16042,N_14915,N_15224);
or U16043 (N_16043,N_14696,N_15586);
or U16044 (N_16044,N_15210,N_15063);
nor U16045 (N_16045,N_14904,N_14699);
xnor U16046 (N_16046,N_14514,N_15135);
and U16047 (N_16047,N_15247,N_14975);
xnor U16048 (N_16048,N_14986,N_15572);
nand U16049 (N_16049,N_15219,N_15303);
nor U16050 (N_16050,N_14709,N_15173);
nand U16051 (N_16051,N_14671,N_15291);
nand U16052 (N_16052,N_14827,N_15068);
xor U16053 (N_16053,N_14492,N_15406);
nand U16054 (N_16054,N_14738,N_14984);
xnor U16055 (N_16055,N_15124,N_14753);
nor U16056 (N_16056,N_15361,N_14576);
nand U16057 (N_16057,N_15216,N_15115);
and U16058 (N_16058,N_15118,N_14617);
and U16059 (N_16059,N_15578,N_14503);
xnor U16060 (N_16060,N_15554,N_15070);
and U16061 (N_16061,N_14785,N_15484);
xnor U16062 (N_16062,N_14859,N_15352);
nor U16063 (N_16063,N_14806,N_14601);
nor U16064 (N_16064,N_15550,N_14568);
or U16065 (N_16065,N_15056,N_15417);
xnor U16066 (N_16066,N_14999,N_14712);
and U16067 (N_16067,N_15258,N_14861);
nand U16068 (N_16068,N_15227,N_14858);
nor U16069 (N_16069,N_15215,N_15287);
or U16070 (N_16070,N_15522,N_14852);
nand U16071 (N_16071,N_14430,N_14882);
and U16072 (N_16072,N_15263,N_15099);
or U16073 (N_16073,N_14998,N_14919);
nand U16074 (N_16074,N_15357,N_15038);
nor U16075 (N_16075,N_15288,N_15547);
or U16076 (N_16076,N_14487,N_14436);
nor U16077 (N_16077,N_14905,N_14639);
and U16078 (N_16078,N_14761,N_14690);
or U16079 (N_16079,N_14922,N_14739);
xor U16080 (N_16080,N_15183,N_14583);
or U16081 (N_16081,N_14943,N_14692);
or U16082 (N_16082,N_14955,N_14965);
or U16083 (N_16083,N_14648,N_14523);
or U16084 (N_16084,N_15395,N_15272);
xor U16085 (N_16085,N_15065,N_14435);
nor U16086 (N_16086,N_14667,N_15420);
nor U16087 (N_16087,N_14551,N_14931);
xor U16088 (N_16088,N_15452,N_14878);
nor U16089 (N_16089,N_14958,N_14788);
nand U16090 (N_16090,N_15549,N_14734);
and U16091 (N_16091,N_15181,N_15466);
nor U16092 (N_16092,N_14653,N_15297);
or U16093 (N_16093,N_15103,N_15440);
and U16094 (N_16094,N_14916,N_15564);
nand U16095 (N_16095,N_14510,N_14427);
xnor U16096 (N_16096,N_15203,N_14640);
nor U16097 (N_16097,N_15242,N_15497);
nand U16098 (N_16098,N_15188,N_14402);
nand U16099 (N_16099,N_14454,N_15031);
or U16100 (N_16100,N_15402,N_14968);
xnor U16101 (N_16101,N_14722,N_14526);
nand U16102 (N_16102,N_14652,N_14883);
xnor U16103 (N_16103,N_14946,N_14819);
nand U16104 (N_16104,N_14947,N_14608);
nor U16105 (N_16105,N_14590,N_15133);
xnor U16106 (N_16106,N_15377,N_15503);
xnor U16107 (N_16107,N_14574,N_14401);
nor U16108 (N_16108,N_15444,N_14647);
xnor U16109 (N_16109,N_15045,N_14596);
nand U16110 (N_16110,N_15166,N_14778);
nor U16111 (N_16111,N_14829,N_14482);
or U16112 (N_16112,N_15443,N_14654);
and U16113 (N_16113,N_15525,N_14442);
nor U16114 (N_16114,N_15460,N_14484);
or U16115 (N_16115,N_15573,N_15566);
and U16116 (N_16116,N_15284,N_15176);
or U16117 (N_16117,N_14832,N_15376);
xnor U16118 (N_16118,N_14408,N_14612);
nand U16119 (N_16119,N_14897,N_15046);
or U16120 (N_16120,N_14846,N_15289);
or U16121 (N_16121,N_14404,N_15270);
and U16122 (N_16122,N_15461,N_15033);
nor U16123 (N_16123,N_15366,N_14567);
and U16124 (N_16124,N_15271,N_14581);
xnor U16125 (N_16125,N_15059,N_15344);
nand U16126 (N_16126,N_14493,N_14784);
and U16127 (N_16127,N_14888,N_15266);
nand U16128 (N_16128,N_15587,N_14937);
xor U16129 (N_16129,N_14988,N_14434);
xnor U16130 (N_16130,N_15199,N_14660);
nor U16131 (N_16131,N_14547,N_15141);
xor U16132 (N_16132,N_14902,N_15285);
or U16133 (N_16133,N_14884,N_15450);
or U16134 (N_16134,N_14438,N_14757);
xor U16135 (N_16135,N_14687,N_14718);
nand U16136 (N_16136,N_14706,N_15388);
nor U16137 (N_16137,N_14451,N_15451);
xor U16138 (N_16138,N_14413,N_14589);
nand U16139 (N_16139,N_15152,N_14835);
xnor U16140 (N_16140,N_14620,N_15540);
nand U16141 (N_16141,N_15424,N_14714);
nor U16142 (N_16142,N_14711,N_14455);
nand U16143 (N_16143,N_14935,N_15146);
or U16144 (N_16144,N_14497,N_15495);
and U16145 (N_16145,N_15596,N_15237);
and U16146 (N_16146,N_14885,N_15312);
or U16147 (N_16147,N_14903,N_14729);
or U16148 (N_16148,N_15411,N_15205);
or U16149 (N_16149,N_15527,N_14766);
nor U16150 (N_16150,N_14745,N_15597);
and U16151 (N_16151,N_15147,N_15177);
and U16152 (N_16152,N_14765,N_15463);
and U16153 (N_16153,N_14834,N_15013);
and U16154 (N_16154,N_14911,N_15209);
xnor U16155 (N_16155,N_14949,N_15009);
nand U16156 (N_16156,N_14939,N_15030);
nand U16157 (N_16157,N_15211,N_14672);
xnor U16158 (N_16158,N_14991,N_14565);
nor U16159 (N_16159,N_14403,N_14823);
nor U16160 (N_16160,N_15568,N_15430);
and U16161 (N_16161,N_15529,N_14979);
nor U16162 (N_16162,N_15375,N_15163);
xnor U16163 (N_16163,N_14923,N_15542);
and U16164 (N_16164,N_14924,N_14595);
or U16165 (N_16165,N_14811,N_14534);
nor U16166 (N_16166,N_14680,N_14456);
and U16167 (N_16167,N_14677,N_14794);
nor U16168 (N_16168,N_14416,N_14755);
nand U16169 (N_16169,N_15077,N_15515);
and U16170 (N_16170,N_14500,N_15071);
or U16171 (N_16171,N_15001,N_15584);
or U16172 (N_16172,N_15506,N_14889);
or U16173 (N_16173,N_15481,N_15394);
xor U16174 (N_16174,N_15302,N_14768);
nand U16175 (N_16175,N_15035,N_15347);
nand U16176 (N_16176,N_14737,N_15275);
nand U16177 (N_16177,N_14466,N_15051);
and U16178 (N_16178,N_15294,N_15520);
nor U16179 (N_16179,N_15043,N_15490);
xnor U16180 (N_16180,N_15083,N_15029);
or U16181 (N_16181,N_15129,N_14941);
and U16182 (N_16182,N_15324,N_15283);
or U16183 (N_16183,N_15410,N_15186);
nand U16184 (N_16184,N_14611,N_14730);
nand U16185 (N_16185,N_15089,N_14426);
nor U16186 (N_16186,N_15208,N_14591);
xnor U16187 (N_16187,N_15261,N_15482);
nor U16188 (N_16188,N_14400,N_15429);
and U16189 (N_16189,N_15563,N_15016);
and U16190 (N_16190,N_14462,N_15061);
xor U16191 (N_16191,N_15425,N_14605);
xnor U16192 (N_16192,N_14586,N_15149);
nand U16193 (N_16193,N_15328,N_15364);
nor U16194 (N_16194,N_14799,N_15259);
xor U16195 (N_16195,N_15116,N_15431);
nand U16196 (N_16196,N_14865,N_14673);
nor U16197 (N_16197,N_15356,N_14525);
nor U16198 (N_16198,N_14544,N_15136);
nand U16199 (N_16199,N_14453,N_15005);
or U16200 (N_16200,N_15414,N_14776);
nand U16201 (N_16201,N_14464,N_15203);
xor U16202 (N_16202,N_14845,N_15529);
and U16203 (N_16203,N_14576,N_14961);
xor U16204 (N_16204,N_15022,N_14976);
and U16205 (N_16205,N_15559,N_14985);
nor U16206 (N_16206,N_14752,N_15338);
and U16207 (N_16207,N_15135,N_15569);
or U16208 (N_16208,N_14810,N_14754);
xnor U16209 (N_16209,N_14523,N_14647);
xor U16210 (N_16210,N_15561,N_14930);
or U16211 (N_16211,N_15539,N_14899);
nand U16212 (N_16212,N_15392,N_14540);
nor U16213 (N_16213,N_14854,N_15147);
and U16214 (N_16214,N_15059,N_15408);
xnor U16215 (N_16215,N_14569,N_15377);
nand U16216 (N_16216,N_14703,N_14404);
and U16217 (N_16217,N_14806,N_15564);
nor U16218 (N_16218,N_15046,N_15316);
xnor U16219 (N_16219,N_15121,N_14993);
nor U16220 (N_16220,N_15225,N_14743);
nand U16221 (N_16221,N_15236,N_15552);
or U16222 (N_16222,N_14683,N_15500);
or U16223 (N_16223,N_14637,N_15012);
or U16224 (N_16224,N_15233,N_15416);
nor U16225 (N_16225,N_14819,N_14857);
nand U16226 (N_16226,N_14699,N_15500);
nand U16227 (N_16227,N_15453,N_14591);
nand U16228 (N_16228,N_15030,N_15441);
nand U16229 (N_16229,N_14767,N_14605);
nand U16230 (N_16230,N_14401,N_14512);
or U16231 (N_16231,N_15428,N_14581);
nor U16232 (N_16232,N_15232,N_14462);
xor U16233 (N_16233,N_15232,N_14961);
nand U16234 (N_16234,N_14879,N_14950);
nand U16235 (N_16235,N_15293,N_15039);
xor U16236 (N_16236,N_15016,N_14555);
and U16237 (N_16237,N_15258,N_14607);
and U16238 (N_16238,N_15074,N_15310);
nand U16239 (N_16239,N_15074,N_14908);
or U16240 (N_16240,N_14558,N_14919);
nor U16241 (N_16241,N_14520,N_15198);
xor U16242 (N_16242,N_15063,N_14663);
nand U16243 (N_16243,N_14422,N_14941);
nand U16244 (N_16244,N_14508,N_15405);
nand U16245 (N_16245,N_14727,N_15525);
and U16246 (N_16246,N_15088,N_14839);
nor U16247 (N_16247,N_14948,N_14588);
or U16248 (N_16248,N_14514,N_15229);
xor U16249 (N_16249,N_15311,N_14823);
nand U16250 (N_16250,N_15480,N_14647);
nor U16251 (N_16251,N_14979,N_15185);
and U16252 (N_16252,N_15360,N_15511);
or U16253 (N_16253,N_14931,N_14506);
or U16254 (N_16254,N_14660,N_14815);
and U16255 (N_16255,N_15420,N_15231);
nor U16256 (N_16256,N_15083,N_14652);
nor U16257 (N_16257,N_14678,N_14462);
xor U16258 (N_16258,N_14762,N_14416);
and U16259 (N_16259,N_14897,N_15213);
xor U16260 (N_16260,N_15446,N_15285);
and U16261 (N_16261,N_15320,N_14653);
or U16262 (N_16262,N_15588,N_15255);
xor U16263 (N_16263,N_14503,N_15238);
and U16264 (N_16264,N_14895,N_15451);
or U16265 (N_16265,N_14802,N_14426);
nor U16266 (N_16266,N_14916,N_15280);
and U16267 (N_16267,N_15027,N_14527);
or U16268 (N_16268,N_14757,N_14609);
nand U16269 (N_16269,N_15502,N_15141);
nor U16270 (N_16270,N_15152,N_14459);
and U16271 (N_16271,N_14676,N_15152);
xor U16272 (N_16272,N_15416,N_15253);
nor U16273 (N_16273,N_15163,N_15357);
and U16274 (N_16274,N_14565,N_15150);
nor U16275 (N_16275,N_14733,N_14590);
nor U16276 (N_16276,N_15508,N_14970);
nor U16277 (N_16277,N_14573,N_15038);
or U16278 (N_16278,N_14592,N_15452);
and U16279 (N_16279,N_14938,N_15393);
and U16280 (N_16280,N_15442,N_14587);
xor U16281 (N_16281,N_15285,N_15587);
or U16282 (N_16282,N_15064,N_14790);
nand U16283 (N_16283,N_15269,N_15053);
xor U16284 (N_16284,N_15045,N_14855);
xnor U16285 (N_16285,N_14798,N_14412);
and U16286 (N_16286,N_15011,N_15488);
nand U16287 (N_16287,N_15105,N_15053);
nor U16288 (N_16288,N_14462,N_15330);
xor U16289 (N_16289,N_15437,N_14996);
nand U16290 (N_16290,N_15481,N_15147);
or U16291 (N_16291,N_14987,N_15025);
nor U16292 (N_16292,N_15302,N_15454);
xor U16293 (N_16293,N_14763,N_14958);
nand U16294 (N_16294,N_15073,N_15524);
nor U16295 (N_16295,N_14588,N_15259);
or U16296 (N_16296,N_14533,N_15338);
nand U16297 (N_16297,N_14505,N_14780);
or U16298 (N_16298,N_15501,N_14844);
nand U16299 (N_16299,N_14678,N_15290);
nand U16300 (N_16300,N_14723,N_14912);
xor U16301 (N_16301,N_15546,N_15240);
nand U16302 (N_16302,N_15121,N_14678);
xnor U16303 (N_16303,N_15514,N_14437);
nor U16304 (N_16304,N_14873,N_15405);
nand U16305 (N_16305,N_14904,N_15482);
xor U16306 (N_16306,N_15041,N_14461);
and U16307 (N_16307,N_15465,N_14659);
or U16308 (N_16308,N_15048,N_15106);
xor U16309 (N_16309,N_14627,N_14970);
nor U16310 (N_16310,N_15518,N_14819);
nand U16311 (N_16311,N_15258,N_15193);
nand U16312 (N_16312,N_15181,N_14934);
nor U16313 (N_16313,N_14896,N_14660);
xnor U16314 (N_16314,N_15420,N_15365);
nor U16315 (N_16315,N_14740,N_14462);
nor U16316 (N_16316,N_14493,N_14908);
and U16317 (N_16317,N_15334,N_15485);
and U16318 (N_16318,N_15467,N_15531);
and U16319 (N_16319,N_14564,N_15149);
and U16320 (N_16320,N_15460,N_15180);
nor U16321 (N_16321,N_14714,N_14937);
or U16322 (N_16322,N_15556,N_15037);
or U16323 (N_16323,N_15422,N_15139);
nand U16324 (N_16324,N_14733,N_15003);
or U16325 (N_16325,N_14954,N_15429);
nor U16326 (N_16326,N_15543,N_14714);
nand U16327 (N_16327,N_15154,N_14496);
nor U16328 (N_16328,N_15431,N_14471);
nor U16329 (N_16329,N_14650,N_14557);
xor U16330 (N_16330,N_14840,N_14900);
nand U16331 (N_16331,N_15290,N_14554);
nand U16332 (N_16332,N_15135,N_15193);
xnor U16333 (N_16333,N_15506,N_14946);
nor U16334 (N_16334,N_14591,N_14988);
xnor U16335 (N_16335,N_14942,N_14853);
or U16336 (N_16336,N_15406,N_14928);
or U16337 (N_16337,N_14678,N_14744);
nand U16338 (N_16338,N_15440,N_14628);
xor U16339 (N_16339,N_15239,N_15009);
xnor U16340 (N_16340,N_15389,N_15543);
or U16341 (N_16341,N_15469,N_14505);
nor U16342 (N_16342,N_14697,N_14842);
or U16343 (N_16343,N_14829,N_14889);
and U16344 (N_16344,N_15008,N_15165);
nand U16345 (N_16345,N_15539,N_15499);
or U16346 (N_16346,N_15170,N_15497);
or U16347 (N_16347,N_15430,N_15527);
or U16348 (N_16348,N_14576,N_14616);
or U16349 (N_16349,N_15485,N_15521);
nand U16350 (N_16350,N_15237,N_15064);
and U16351 (N_16351,N_15211,N_15326);
or U16352 (N_16352,N_15456,N_14773);
and U16353 (N_16353,N_15452,N_14410);
nand U16354 (N_16354,N_14947,N_15561);
and U16355 (N_16355,N_15172,N_15322);
nor U16356 (N_16356,N_14774,N_14962);
or U16357 (N_16357,N_14586,N_15094);
or U16358 (N_16358,N_15329,N_14939);
and U16359 (N_16359,N_15133,N_14795);
nand U16360 (N_16360,N_14754,N_15232);
xnor U16361 (N_16361,N_14704,N_14424);
nand U16362 (N_16362,N_15209,N_14752);
xnor U16363 (N_16363,N_15520,N_15498);
nor U16364 (N_16364,N_15580,N_15051);
and U16365 (N_16365,N_15596,N_15121);
nand U16366 (N_16366,N_15479,N_14958);
xor U16367 (N_16367,N_14661,N_15521);
nand U16368 (N_16368,N_14746,N_14445);
or U16369 (N_16369,N_15085,N_15545);
and U16370 (N_16370,N_14664,N_15195);
and U16371 (N_16371,N_15198,N_14631);
nand U16372 (N_16372,N_14524,N_14875);
nand U16373 (N_16373,N_14501,N_14985);
and U16374 (N_16374,N_14495,N_14950);
or U16375 (N_16375,N_14806,N_14551);
nor U16376 (N_16376,N_15098,N_15111);
xor U16377 (N_16377,N_15546,N_14426);
nor U16378 (N_16378,N_15212,N_15533);
or U16379 (N_16379,N_15577,N_14580);
nand U16380 (N_16380,N_15161,N_15000);
nand U16381 (N_16381,N_14436,N_14907);
or U16382 (N_16382,N_15000,N_14742);
xnor U16383 (N_16383,N_14914,N_15554);
or U16384 (N_16384,N_15357,N_15096);
nand U16385 (N_16385,N_14642,N_15594);
and U16386 (N_16386,N_14424,N_15214);
and U16387 (N_16387,N_15490,N_15041);
and U16388 (N_16388,N_14553,N_14546);
and U16389 (N_16389,N_14668,N_14997);
or U16390 (N_16390,N_15212,N_15234);
and U16391 (N_16391,N_15152,N_15270);
nand U16392 (N_16392,N_15152,N_14911);
and U16393 (N_16393,N_14985,N_15025);
nand U16394 (N_16394,N_14750,N_15584);
nor U16395 (N_16395,N_14820,N_14708);
xnor U16396 (N_16396,N_14599,N_15235);
or U16397 (N_16397,N_14791,N_14515);
or U16398 (N_16398,N_15474,N_14521);
or U16399 (N_16399,N_15287,N_14469);
xnor U16400 (N_16400,N_15366,N_15362);
and U16401 (N_16401,N_14939,N_14855);
xor U16402 (N_16402,N_14476,N_14667);
nor U16403 (N_16403,N_15489,N_15027);
or U16404 (N_16404,N_14515,N_15124);
nor U16405 (N_16405,N_14838,N_15336);
nand U16406 (N_16406,N_14988,N_15172);
or U16407 (N_16407,N_15294,N_15244);
xnor U16408 (N_16408,N_14738,N_15495);
and U16409 (N_16409,N_15087,N_15494);
and U16410 (N_16410,N_14480,N_15440);
xor U16411 (N_16411,N_15332,N_14735);
nand U16412 (N_16412,N_15337,N_15203);
and U16413 (N_16413,N_15368,N_15184);
nor U16414 (N_16414,N_14406,N_15346);
nor U16415 (N_16415,N_14443,N_14990);
nand U16416 (N_16416,N_14863,N_15241);
xor U16417 (N_16417,N_15474,N_14979);
xor U16418 (N_16418,N_15599,N_15538);
nand U16419 (N_16419,N_15449,N_15521);
nor U16420 (N_16420,N_14931,N_14555);
nand U16421 (N_16421,N_15333,N_14969);
xor U16422 (N_16422,N_15318,N_15092);
nor U16423 (N_16423,N_15058,N_14835);
or U16424 (N_16424,N_14863,N_14852);
nand U16425 (N_16425,N_14594,N_14519);
xnor U16426 (N_16426,N_14458,N_14910);
nand U16427 (N_16427,N_14831,N_14594);
nor U16428 (N_16428,N_15093,N_14645);
xnor U16429 (N_16429,N_15081,N_15334);
or U16430 (N_16430,N_15176,N_14918);
or U16431 (N_16431,N_14402,N_15352);
or U16432 (N_16432,N_15096,N_15487);
nor U16433 (N_16433,N_15364,N_14664);
and U16434 (N_16434,N_14989,N_14761);
nor U16435 (N_16435,N_14549,N_14660);
or U16436 (N_16436,N_15573,N_14679);
xnor U16437 (N_16437,N_14856,N_14826);
nor U16438 (N_16438,N_14952,N_14764);
xnor U16439 (N_16439,N_14910,N_14865);
nand U16440 (N_16440,N_14855,N_14720);
or U16441 (N_16441,N_15033,N_15227);
and U16442 (N_16442,N_15314,N_14700);
xor U16443 (N_16443,N_14480,N_14963);
xnor U16444 (N_16444,N_15341,N_15583);
xor U16445 (N_16445,N_14788,N_14882);
or U16446 (N_16446,N_14758,N_15227);
or U16447 (N_16447,N_14516,N_14688);
and U16448 (N_16448,N_15437,N_14879);
and U16449 (N_16449,N_15247,N_14789);
nor U16450 (N_16450,N_15503,N_15381);
and U16451 (N_16451,N_14434,N_15445);
nor U16452 (N_16452,N_15201,N_14880);
nor U16453 (N_16453,N_14918,N_15437);
nand U16454 (N_16454,N_14500,N_15055);
xor U16455 (N_16455,N_14843,N_14458);
or U16456 (N_16456,N_14984,N_14406);
nand U16457 (N_16457,N_14870,N_14425);
and U16458 (N_16458,N_14755,N_15435);
or U16459 (N_16459,N_14644,N_15353);
nand U16460 (N_16460,N_15273,N_14839);
xnor U16461 (N_16461,N_15470,N_14774);
nor U16462 (N_16462,N_15129,N_14601);
and U16463 (N_16463,N_15342,N_14639);
and U16464 (N_16464,N_14463,N_15111);
nor U16465 (N_16465,N_14735,N_15439);
and U16466 (N_16466,N_15027,N_15180);
and U16467 (N_16467,N_15088,N_15400);
or U16468 (N_16468,N_15528,N_14710);
and U16469 (N_16469,N_15004,N_15171);
xnor U16470 (N_16470,N_15593,N_15312);
nand U16471 (N_16471,N_14998,N_14792);
xnor U16472 (N_16472,N_15315,N_15543);
nand U16473 (N_16473,N_15320,N_14669);
nor U16474 (N_16474,N_14941,N_14938);
xor U16475 (N_16475,N_15031,N_14736);
or U16476 (N_16476,N_14685,N_14576);
or U16477 (N_16477,N_15247,N_14997);
xor U16478 (N_16478,N_14750,N_14781);
or U16479 (N_16479,N_14558,N_15487);
or U16480 (N_16480,N_14989,N_15379);
xnor U16481 (N_16481,N_15457,N_15477);
or U16482 (N_16482,N_15534,N_14480);
or U16483 (N_16483,N_15320,N_15017);
nor U16484 (N_16484,N_15461,N_14637);
nor U16485 (N_16485,N_15211,N_14593);
xor U16486 (N_16486,N_15508,N_14553);
or U16487 (N_16487,N_15088,N_15371);
nand U16488 (N_16488,N_14891,N_15142);
nand U16489 (N_16489,N_15340,N_14956);
xor U16490 (N_16490,N_14701,N_14885);
xnor U16491 (N_16491,N_14583,N_15470);
nand U16492 (N_16492,N_14641,N_15499);
and U16493 (N_16493,N_15104,N_15191);
nor U16494 (N_16494,N_14805,N_14443);
nor U16495 (N_16495,N_15227,N_14486);
or U16496 (N_16496,N_14653,N_15146);
and U16497 (N_16497,N_14961,N_14652);
nand U16498 (N_16498,N_15570,N_14525);
nor U16499 (N_16499,N_15217,N_15343);
nand U16500 (N_16500,N_15296,N_15040);
or U16501 (N_16501,N_15078,N_14472);
or U16502 (N_16502,N_15319,N_14916);
nand U16503 (N_16503,N_14740,N_14796);
nor U16504 (N_16504,N_15420,N_15559);
nand U16505 (N_16505,N_14608,N_15477);
nand U16506 (N_16506,N_14544,N_15422);
xor U16507 (N_16507,N_14495,N_14460);
nor U16508 (N_16508,N_15043,N_15374);
and U16509 (N_16509,N_15188,N_14442);
and U16510 (N_16510,N_14607,N_15302);
xnor U16511 (N_16511,N_14677,N_14722);
nor U16512 (N_16512,N_15500,N_15387);
nor U16513 (N_16513,N_14423,N_14592);
or U16514 (N_16514,N_15094,N_14589);
or U16515 (N_16515,N_14953,N_15177);
nand U16516 (N_16516,N_15367,N_14817);
nor U16517 (N_16517,N_14881,N_15504);
nor U16518 (N_16518,N_15121,N_15203);
nand U16519 (N_16519,N_15344,N_14826);
or U16520 (N_16520,N_15334,N_14614);
and U16521 (N_16521,N_15452,N_15236);
or U16522 (N_16522,N_15312,N_14492);
nor U16523 (N_16523,N_15455,N_14417);
nor U16524 (N_16524,N_15086,N_15359);
or U16525 (N_16525,N_15318,N_15027);
xor U16526 (N_16526,N_14617,N_15110);
nand U16527 (N_16527,N_14840,N_14439);
nor U16528 (N_16528,N_14942,N_14790);
xnor U16529 (N_16529,N_15048,N_15558);
nand U16530 (N_16530,N_15200,N_15369);
xor U16531 (N_16531,N_15397,N_14559);
and U16532 (N_16532,N_15460,N_15341);
nand U16533 (N_16533,N_14652,N_15064);
or U16534 (N_16534,N_15137,N_15553);
or U16535 (N_16535,N_14989,N_15255);
and U16536 (N_16536,N_14528,N_14559);
nand U16537 (N_16537,N_14486,N_14920);
and U16538 (N_16538,N_15395,N_15067);
xnor U16539 (N_16539,N_15088,N_15112);
or U16540 (N_16540,N_14861,N_14939);
nand U16541 (N_16541,N_14666,N_15555);
nand U16542 (N_16542,N_15316,N_15532);
and U16543 (N_16543,N_15369,N_15391);
nand U16544 (N_16544,N_15152,N_14986);
nor U16545 (N_16545,N_14624,N_14796);
nand U16546 (N_16546,N_14977,N_15454);
xor U16547 (N_16547,N_14530,N_15562);
nor U16548 (N_16548,N_15336,N_15009);
or U16549 (N_16549,N_14706,N_14723);
nor U16550 (N_16550,N_15160,N_14605);
nor U16551 (N_16551,N_14692,N_15522);
and U16552 (N_16552,N_15191,N_14472);
xnor U16553 (N_16553,N_14963,N_14802);
xor U16554 (N_16554,N_15330,N_15005);
or U16555 (N_16555,N_14460,N_14738);
xnor U16556 (N_16556,N_15525,N_15246);
nand U16557 (N_16557,N_14829,N_14629);
and U16558 (N_16558,N_14513,N_14872);
or U16559 (N_16559,N_14954,N_14633);
or U16560 (N_16560,N_14569,N_14779);
and U16561 (N_16561,N_14405,N_14864);
nor U16562 (N_16562,N_14427,N_15031);
nand U16563 (N_16563,N_15435,N_15280);
nor U16564 (N_16564,N_14489,N_15116);
xnor U16565 (N_16565,N_14682,N_14993);
nand U16566 (N_16566,N_14846,N_15407);
nor U16567 (N_16567,N_15433,N_15049);
nand U16568 (N_16568,N_15192,N_14662);
and U16569 (N_16569,N_14848,N_15113);
and U16570 (N_16570,N_14468,N_14588);
and U16571 (N_16571,N_15070,N_15248);
nor U16572 (N_16572,N_14593,N_15489);
xnor U16573 (N_16573,N_15430,N_14639);
xor U16574 (N_16574,N_14449,N_14547);
xor U16575 (N_16575,N_14555,N_14758);
nor U16576 (N_16576,N_15167,N_14480);
xnor U16577 (N_16577,N_15222,N_15512);
or U16578 (N_16578,N_14465,N_14867);
nand U16579 (N_16579,N_14536,N_15117);
or U16580 (N_16580,N_15342,N_15390);
nor U16581 (N_16581,N_14417,N_14717);
and U16582 (N_16582,N_14750,N_14935);
xor U16583 (N_16583,N_14715,N_14476);
nand U16584 (N_16584,N_15090,N_15127);
nor U16585 (N_16585,N_15341,N_14568);
or U16586 (N_16586,N_15113,N_15149);
xnor U16587 (N_16587,N_15196,N_14534);
or U16588 (N_16588,N_14478,N_14849);
nor U16589 (N_16589,N_15546,N_14513);
xnor U16590 (N_16590,N_15302,N_14866);
or U16591 (N_16591,N_15144,N_14826);
nor U16592 (N_16592,N_14976,N_15327);
nand U16593 (N_16593,N_15456,N_14963);
nor U16594 (N_16594,N_14464,N_15275);
nor U16595 (N_16595,N_15314,N_14543);
and U16596 (N_16596,N_14852,N_15138);
nand U16597 (N_16597,N_14559,N_14923);
or U16598 (N_16598,N_15239,N_14877);
nand U16599 (N_16599,N_14952,N_15366);
xnor U16600 (N_16600,N_15505,N_14966);
nor U16601 (N_16601,N_14470,N_15371);
nor U16602 (N_16602,N_15006,N_14625);
xor U16603 (N_16603,N_15204,N_15570);
nand U16604 (N_16604,N_15005,N_15279);
and U16605 (N_16605,N_15573,N_14735);
nand U16606 (N_16606,N_14536,N_14855);
or U16607 (N_16607,N_14976,N_15349);
or U16608 (N_16608,N_14573,N_14782);
xnor U16609 (N_16609,N_15483,N_14606);
nor U16610 (N_16610,N_14753,N_15458);
or U16611 (N_16611,N_14704,N_15216);
nand U16612 (N_16612,N_14997,N_14888);
and U16613 (N_16613,N_14636,N_14522);
nor U16614 (N_16614,N_14612,N_14850);
nor U16615 (N_16615,N_14746,N_15044);
nand U16616 (N_16616,N_15329,N_15271);
nand U16617 (N_16617,N_15432,N_15028);
nand U16618 (N_16618,N_14605,N_15513);
and U16619 (N_16619,N_15505,N_15174);
xnor U16620 (N_16620,N_14883,N_14787);
and U16621 (N_16621,N_15250,N_14546);
or U16622 (N_16622,N_14831,N_15399);
nor U16623 (N_16623,N_15440,N_14705);
and U16624 (N_16624,N_14871,N_15571);
or U16625 (N_16625,N_15241,N_15387);
nor U16626 (N_16626,N_15200,N_14677);
nor U16627 (N_16627,N_14893,N_15491);
xnor U16628 (N_16628,N_15594,N_15257);
and U16629 (N_16629,N_15069,N_15488);
or U16630 (N_16630,N_15358,N_15559);
xnor U16631 (N_16631,N_14532,N_14465);
nand U16632 (N_16632,N_14494,N_14633);
nand U16633 (N_16633,N_15279,N_14499);
or U16634 (N_16634,N_14487,N_15383);
and U16635 (N_16635,N_14839,N_15291);
xor U16636 (N_16636,N_14940,N_15475);
nand U16637 (N_16637,N_15293,N_14441);
or U16638 (N_16638,N_14621,N_15250);
and U16639 (N_16639,N_14906,N_14437);
xor U16640 (N_16640,N_15031,N_14469);
or U16641 (N_16641,N_14754,N_15279);
and U16642 (N_16642,N_15049,N_14434);
xor U16643 (N_16643,N_14630,N_14725);
nand U16644 (N_16644,N_15548,N_14642);
xnor U16645 (N_16645,N_15451,N_15354);
and U16646 (N_16646,N_14630,N_15114);
nand U16647 (N_16647,N_14437,N_14723);
and U16648 (N_16648,N_15095,N_14751);
or U16649 (N_16649,N_15054,N_14880);
xnor U16650 (N_16650,N_14714,N_14590);
nor U16651 (N_16651,N_14995,N_14596);
nand U16652 (N_16652,N_14538,N_15275);
nor U16653 (N_16653,N_14471,N_14831);
or U16654 (N_16654,N_15288,N_14903);
xnor U16655 (N_16655,N_14838,N_14444);
nand U16656 (N_16656,N_14712,N_14752);
or U16657 (N_16657,N_15407,N_14996);
nor U16658 (N_16658,N_15435,N_14764);
nand U16659 (N_16659,N_15269,N_15122);
nor U16660 (N_16660,N_15152,N_15506);
xor U16661 (N_16661,N_15594,N_15394);
xnor U16662 (N_16662,N_15375,N_15555);
xor U16663 (N_16663,N_15350,N_14756);
nand U16664 (N_16664,N_15360,N_14805);
xor U16665 (N_16665,N_14761,N_15233);
nand U16666 (N_16666,N_14415,N_14905);
and U16667 (N_16667,N_14456,N_15099);
and U16668 (N_16668,N_15285,N_15536);
xnor U16669 (N_16669,N_14941,N_14457);
and U16670 (N_16670,N_14439,N_15507);
xnor U16671 (N_16671,N_15100,N_14775);
nand U16672 (N_16672,N_15332,N_15298);
nand U16673 (N_16673,N_14553,N_14712);
nor U16674 (N_16674,N_15340,N_14673);
nor U16675 (N_16675,N_14843,N_15559);
and U16676 (N_16676,N_15519,N_15159);
xnor U16677 (N_16677,N_14662,N_15127);
xor U16678 (N_16678,N_14434,N_14507);
and U16679 (N_16679,N_15528,N_14794);
or U16680 (N_16680,N_14419,N_14486);
or U16681 (N_16681,N_14593,N_15299);
xnor U16682 (N_16682,N_14939,N_14405);
or U16683 (N_16683,N_14401,N_14830);
and U16684 (N_16684,N_15311,N_14518);
or U16685 (N_16685,N_14589,N_14441);
xor U16686 (N_16686,N_15100,N_14817);
nor U16687 (N_16687,N_14665,N_15148);
nand U16688 (N_16688,N_15058,N_14670);
and U16689 (N_16689,N_15486,N_15471);
or U16690 (N_16690,N_14609,N_14998);
and U16691 (N_16691,N_14936,N_15231);
xnor U16692 (N_16692,N_14486,N_15199);
or U16693 (N_16693,N_15474,N_15342);
xnor U16694 (N_16694,N_15262,N_15031);
nor U16695 (N_16695,N_15077,N_14772);
xnor U16696 (N_16696,N_14615,N_15010);
nor U16697 (N_16697,N_15510,N_15582);
or U16698 (N_16698,N_14873,N_14518);
xnor U16699 (N_16699,N_15094,N_14727);
or U16700 (N_16700,N_14947,N_14491);
nand U16701 (N_16701,N_14773,N_15278);
xnor U16702 (N_16702,N_15052,N_14541);
and U16703 (N_16703,N_14493,N_14951);
xor U16704 (N_16704,N_15378,N_15058);
or U16705 (N_16705,N_14500,N_15349);
nor U16706 (N_16706,N_14529,N_14798);
nand U16707 (N_16707,N_15259,N_14529);
xnor U16708 (N_16708,N_14600,N_14963);
nor U16709 (N_16709,N_14844,N_14591);
and U16710 (N_16710,N_14736,N_15110);
nor U16711 (N_16711,N_14644,N_14607);
or U16712 (N_16712,N_15551,N_15531);
nor U16713 (N_16713,N_14473,N_15442);
nand U16714 (N_16714,N_15509,N_14769);
and U16715 (N_16715,N_15102,N_14730);
nor U16716 (N_16716,N_15517,N_15537);
nand U16717 (N_16717,N_14726,N_14578);
nor U16718 (N_16718,N_14981,N_14597);
or U16719 (N_16719,N_15551,N_14623);
or U16720 (N_16720,N_14952,N_14796);
nor U16721 (N_16721,N_15083,N_14790);
or U16722 (N_16722,N_14532,N_15165);
or U16723 (N_16723,N_14723,N_15582);
and U16724 (N_16724,N_14929,N_14767);
or U16725 (N_16725,N_14844,N_15166);
nand U16726 (N_16726,N_15499,N_14990);
xor U16727 (N_16727,N_14672,N_14703);
or U16728 (N_16728,N_15391,N_14553);
or U16729 (N_16729,N_14754,N_14574);
or U16730 (N_16730,N_14704,N_14769);
nand U16731 (N_16731,N_15217,N_14422);
or U16732 (N_16732,N_14618,N_15005);
and U16733 (N_16733,N_15533,N_15182);
and U16734 (N_16734,N_15012,N_14919);
xor U16735 (N_16735,N_14599,N_15355);
xnor U16736 (N_16736,N_14845,N_14551);
nand U16737 (N_16737,N_15145,N_15330);
nor U16738 (N_16738,N_15459,N_14457);
nor U16739 (N_16739,N_15035,N_15444);
nor U16740 (N_16740,N_15267,N_14465);
nand U16741 (N_16741,N_15451,N_14418);
and U16742 (N_16742,N_14528,N_15099);
and U16743 (N_16743,N_15158,N_14515);
and U16744 (N_16744,N_15158,N_14827);
nand U16745 (N_16745,N_14405,N_14464);
xnor U16746 (N_16746,N_14663,N_14755);
nor U16747 (N_16747,N_15400,N_15061);
nand U16748 (N_16748,N_15528,N_14461);
and U16749 (N_16749,N_14730,N_14600);
and U16750 (N_16750,N_15122,N_14418);
nand U16751 (N_16751,N_14746,N_15432);
or U16752 (N_16752,N_15295,N_15081);
or U16753 (N_16753,N_14465,N_14732);
nand U16754 (N_16754,N_14821,N_15129);
xor U16755 (N_16755,N_15407,N_15589);
or U16756 (N_16756,N_14761,N_15119);
nand U16757 (N_16757,N_15143,N_15154);
xnor U16758 (N_16758,N_14602,N_14995);
or U16759 (N_16759,N_15498,N_15070);
or U16760 (N_16760,N_14629,N_14960);
and U16761 (N_16761,N_15479,N_15139);
xor U16762 (N_16762,N_15255,N_15290);
and U16763 (N_16763,N_15458,N_14544);
and U16764 (N_16764,N_15486,N_15329);
xor U16765 (N_16765,N_14915,N_14637);
nand U16766 (N_16766,N_15308,N_14615);
or U16767 (N_16767,N_14650,N_14695);
xor U16768 (N_16768,N_14732,N_15397);
xor U16769 (N_16769,N_15107,N_14806);
and U16770 (N_16770,N_15591,N_14458);
nor U16771 (N_16771,N_14862,N_14758);
and U16772 (N_16772,N_14962,N_14420);
or U16773 (N_16773,N_14909,N_15174);
xor U16774 (N_16774,N_14441,N_15310);
or U16775 (N_16775,N_14791,N_15455);
or U16776 (N_16776,N_15470,N_15585);
xor U16777 (N_16777,N_15490,N_14680);
or U16778 (N_16778,N_15115,N_14903);
nor U16779 (N_16779,N_14970,N_15005);
nand U16780 (N_16780,N_15099,N_15003);
xor U16781 (N_16781,N_15439,N_15547);
or U16782 (N_16782,N_15290,N_15473);
xor U16783 (N_16783,N_15599,N_15576);
nor U16784 (N_16784,N_15171,N_15413);
nand U16785 (N_16785,N_15379,N_14506);
nand U16786 (N_16786,N_14816,N_15507);
and U16787 (N_16787,N_15226,N_14882);
and U16788 (N_16788,N_15018,N_15478);
xnor U16789 (N_16789,N_14961,N_14429);
xor U16790 (N_16790,N_14741,N_15309);
nand U16791 (N_16791,N_15469,N_15529);
or U16792 (N_16792,N_15448,N_15079);
nor U16793 (N_16793,N_14553,N_14548);
nor U16794 (N_16794,N_14445,N_14945);
xnor U16795 (N_16795,N_15592,N_15234);
and U16796 (N_16796,N_14477,N_14417);
nor U16797 (N_16797,N_15068,N_15046);
xnor U16798 (N_16798,N_15159,N_14425);
nand U16799 (N_16799,N_15567,N_15558);
or U16800 (N_16800,N_16093,N_16259);
nand U16801 (N_16801,N_15992,N_16261);
xor U16802 (N_16802,N_16598,N_15814);
xor U16803 (N_16803,N_16303,N_16051);
and U16804 (N_16804,N_15903,N_16284);
nor U16805 (N_16805,N_16160,N_16139);
xor U16806 (N_16806,N_16782,N_16256);
and U16807 (N_16807,N_15648,N_15916);
nand U16808 (N_16808,N_15717,N_16476);
nand U16809 (N_16809,N_16527,N_16566);
or U16810 (N_16810,N_16709,N_16528);
or U16811 (N_16811,N_16588,N_16411);
nor U16812 (N_16812,N_16216,N_16014);
and U16813 (N_16813,N_16656,N_15969);
and U16814 (N_16814,N_15966,N_15973);
nor U16815 (N_16815,N_15637,N_16280);
or U16816 (N_16816,N_16100,N_16475);
and U16817 (N_16817,N_15993,N_15659);
or U16818 (N_16818,N_16773,N_16300);
nor U16819 (N_16819,N_16186,N_16045);
xnor U16820 (N_16820,N_16589,N_15693);
and U16821 (N_16821,N_16645,N_16163);
nand U16822 (N_16822,N_15673,N_16655);
nor U16823 (N_16823,N_16473,N_16370);
and U16824 (N_16824,N_16550,N_16771);
and U16825 (N_16825,N_15641,N_15758);
xor U16826 (N_16826,N_16657,N_15664);
nor U16827 (N_16827,N_15628,N_16615);
or U16828 (N_16828,N_15729,N_16237);
nand U16829 (N_16829,N_16480,N_16437);
and U16830 (N_16830,N_16441,N_15981);
and U16831 (N_16831,N_16315,N_15854);
nand U16832 (N_16832,N_16459,N_16125);
or U16833 (N_16833,N_15788,N_16152);
or U16834 (N_16834,N_15895,N_16096);
xnor U16835 (N_16835,N_15864,N_15978);
nand U16836 (N_16836,N_15802,N_16376);
nor U16837 (N_16837,N_15679,N_16583);
xor U16838 (N_16838,N_16552,N_15710);
nand U16839 (N_16839,N_16135,N_15619);
xor U16840 (N_16840,N_16224,N_16623);
nand U16841 (N_16841,N_16688,N_16357);
or U16842 (N_16842,N_16503,N_16166);
xor U16843 (N_16843,N_16714,N_15774);
or U16844 (N_16844,N_16724,N_16121);
or U16845 (N_16845,N_15736,N_15761);
or U16846 (N_16846,N_15707,N_16639);
nor U16847 (N_16847,N_15692,N_16056);
nand U16848 (N_16848,N_16225,N_15951);
nand U16849 (N_16849,N_16016,N_16708);
nor U16850 (N_16850,N_16103,N_16454);
nand U16851 (N_16851,N_16472,N_16223);
or U16852 (N_16852,N_16696,N_16666);
xor U16853 (N_16853,N_16187,N_16307);
nand U16854 (N_16854,N_15826,N_15672);
nor U16855 (N_16855,N_16784,N_15605);
xnor U16856 (N_16856,N_16567,N_15747);
xnor U16857 (N_16857,N_16742,N_15732);
or U16858 (N_16858,N_16294,N_15714);
nand U16859 (N_16859,N_16629,N_16047);
nor U16860 (N_16860,N_16574,N_16424);
nand U16861 (N_16861,N_16579,N_16003);
and U16862 (N_16862,N_15680,N_15794);
nand U16863 (N_16863,N_16283,N_15769);
xor U16864 (N_16864,N_15937,N_16366);
xnor U16865 (N_16865,N_15909,N_16272);
nand U16866 (N_16866,N_15793,N_16354);
or U16867 (N_16867,N_15810,N_15801);
and U16868 (N_16868,N_16442,N_15789);
nand U16869 (N_16869,N_16532,N_16618);
or U16870 (N_16870,N_16250,N_16607);
or U16871 (N_16871,N_16034,N_15811);
and U16872 (N_16872,N_16154,N_16597);
nor U16873 (N_16873,N_16642,N_16520);
xnor U16874 (N_16874,N_16342,N_15927);
nand U16875 (N_16875,N_15816,N_16543);
and U16876 (N_16876,N_16146,N_16698);
nand U16877 (N_16877,N_16388,N_16221);
nor U16878 (N_16878,N_16327,N_16478);
xnor U16879 (N_16879,N_15636,N_16514);
and U16880 (N_16880,N_16384,N_16195);
nor U16881 (N_16881,N_16505,N_15625);
nand U16882 (N_16882,N_16368,N_15829);
xnor U16883 (N_16883,N_15936,N_16251);
or U16884 (N_16884,N_15611,N_16627);
nor U16885 (N_16885,N_15799,N_16364);
and U16886 (N_16886,N_15866,N_15959);
and U16887 (N_16887,N_16767,N_16020);
nand U16888 (N_16888,N_16752,N_16274);
and U16889 (N_16889,N_15630,N_16290);
xor U16890 (N_16890,N_15610,N_16746);
xnor U16891 (N_16891,N_16390,N_15975);
xor U16892 (N_16892,N_16559,N_15721);
xnor U16893 (N_16893,N_15681,N_15887);
xnor U16894 (N_16894,N_15857,N_16205);
xnor U16895 (N_16895,N_15674,N_15771);
nor U16896 (N_16896,N_16270,N_16030);
nor U16897 (N_16897,N_15735,N_15930);
nor U16898 (N_16898,N_16293,N_16423);
nand U16899 (N_16899,N_16621,N_16391);
xnor U16900 (N_16900,N_16078,N_16076);
or U16901 (N_16901,N_16636,N_16153);
nor U16902 (N_16902,N_15827,N_16281);
nand U16903 (N_16903,N_16510,N_16455);
xnor U16904 (N_16904,N_16622,N_16780);
nand U16905 (N_16905,N_16105,N_16386);
nand U16906 (N_16906,N_16491,N_16634);
nand U16907 (N_16907,N_15698,N_15987);
nand U16908 (N_16908,N_16213,N_15911);
nor U16909 (N_16909,N_15748,N_15656);
and U16910 (N_16910,N_16687,N_16501);
xor U16911 (N_16911,N_16433,N_16027);
nor U16912 (N_16912,N_16207,N_16718);
xor U16913 (N_16913,N_16155,N_16490);
nand U16914 (N_16914,N_15878,N_15668);
and U16915 (N_16915,N_15686,N_16333);
and U16916 (N_16916,N_15932,N_15704);
and U16917 (N_16917,N_16568,N_16326);
nand U16918 (N_16918,N_16264,N_15730);
nand U16919 (N_16919,N_15902,N_16551);
nand U16920 (N_16920,N_15905,N_15614);
nor U16921 (N_16921,N_15928,N_15782);
nand U16922 (N_16922,N_16091,N_16233);
and U16923 (N_16923,N_16791,N_16422);
nor U16924 (N_16924,N_16576,N_16499);
xor U16925 (N_16925,N_16596,N_16081);
and U16926 (N_16926,N_16498,N_16113);
nor U16927 (N_16927,N_16603,N_16608);
nand U16928 (N_16928,N_16434,N_16012);
xor U16929 (N_16929,N_16164,N_15888);
nand U16930 (N_16930,N_16547,N_16753);
xnor U16931 (N_16931,N_16005,N_16601);
xnor U16932 (N_16932,N_15785,N_15926);
nand U16933 (N_16933,N_16173,N_16244);
and U16934 (N_16934,N_16074,N_15696);
nand U16935 (N_16935,N_15723,N_15892);
or U16936 (N_16936,N_15792,N_15777);
nand U16937 (N_16937,N_15703,N_16789);
and U16938 (N_16938,N_16319,N_16339);
nor U16939 (N_16939,N_16040,N_16446);
and U16940 (N_16940,N_16352,N_15775);
nor U16941 (N_16941,N_16479,N_15861);
nor U16942 (N_16942,N_16408,N_16720);
nor U16943 (N_16943,N_16196,N_16123);
nand U16944 (N_16944,N_15868,N_15832);
and U16945 (N_16945,N_16594,N_15876);
and U16946 (N_16946,N_16521,N_16534);
xnor U16947 (N_16947,N_15813,N_16675);
and U16948 (N_16948,N_15918,N_15970);
nand U16949 (N_16949,N_16204,N_15746);
and U16950 (N_16950,N_15889,N_15634);
and U16951 (N_16951,N_16697,N_16353);
and U16952 (N_16952,N_16108,N_15778);
and U16953 (N_16953,N_15645,N_15865);
nand U16954 (N_16954,N_16212,N_16757);
nand U16955 (N_16955,N_16329,N_16763);
nand U16956 (N_16956,N_16430,N_16343);
nand U16957 (N_16957,N_16402,N_15952);
xor U16958 (N_16958,N_16448,N_16723);
xnor U16959 (N_16959,N_16147,N_16018);
and U16960 (N_16960,N_16144,N_16725);
xor U16961 (N_16961,N_15665,N_15867);
and U16962 (N_16962,N_15862,N_16631);
and U16963 (N_16963,N_16511,N_16744);
xnor U16964 (N_16964,N_16109,N_15961);
and U16965 (N_16965,N_16316,N_16513);
or U16966 (N_16966,N_15609,N_15731);
nor U16967 (N_16967,N_16586,N_16120);
nor U16968 (N_16968,N_15727,N_15694);
xnor U16969 (N_16969,N_16277,N_15880);
or U16970 (N_16970,N_16545,N_16082);
or U16971 (N_16971,N_16592,N_16463);
and U16972 (N_16972,N_15820,N_15818);
and U16973 (N_16973,N_16200,N_16575);
and U16974 (N_16974,N_15950,N_15910);
or U16975 (N_16975,N_16361,N_16776);
nand U16976 (N_16976,N_15836,N_16711);
xor U16977 (N_16977,N_16359,N_16395);
nor U16978 (N_16978,N_16796,N_16462);
or U16979 (N_16979,N_16477,N_16418);
xor U16980 (N_16980,N_16273,N_16112);
nor U16981 (N_16981,N_16383,N_16682);
and U16982 (N_16982,N_15660,N_16584);
or U16983 (N_16983,N_16210,N_15995);
or U16984 (N_16984,N_16786,N_16614);
or U16985 (N_16985,N_16322,N_16255);
and U16986 (N_16986,N_15702,N_15881);
nand U16987 (N_16987,N_16132,N_16755);
nor U16988 (N_16988,N_16214,N_15741);
nor U16989 (N_16989,N_15671,N_16149);
nor U16990 (N_16990,N_16556,N_16457);
xor U16991 (N_16991,N_15850,N_16136);
nor U16992 (N_16992,N_15804,N_16063);
or U16993 (N_16993,N_16525,N_15682);
or U16994 (N_16994,N_16737,N_16138);
xor U16995 (N_16995,N_15651,N_15815);
nand U16996 (N_16996,N_16181,N_16247);
nand U16997 (N_16997,N_15797,N_15808);
nor U16998 (N_16998,N_16208,N_15765);
nand U16999 (N_16999,N_16407,N_16193);
nor U17000 (N_17000,N_16695,N_15786);
and U17001 (N_17001,N_16538,N_16308);
nand U17002 (N_17002,N_15945,N_16038);
xor U17003 (N_17003,N_15980,N_16335);
xor U17004 (N_17004,N_16373,N_16481);
and U17005 (N_17005,N_15776,N_15608);
or U17006 (N_17006,N_15967,N_16661);
nand U17007 (N_17007,N_16450,N_16468);
and U17008 (N_17008,N_16649,N_16070);
and U17009 (N_17009,N_16232,N_15644);
xor U17010 (N_17010,N_15824,N_15766);
or U17011 (N_17011,N_16190,N_16516);
nand U17012 (N_17012,N_16385,N_16346);
nand U17013 (N_17013,N_16297,N_16797);
or U17014 (N_17014,N_15849,N_16793);
nor U17015 (N_17015,N_16119,N_16330);
nor U17016 (N_17016,N_15896,N_16569);
or U17017 (N_17017,N_16654,N_16600);
xor U17018 (N_17018,N_16519,N_15873);
xnor U17019 (N_17019,N_16350,N_15718);
nor U17020 (N_17020,N_16658,N_16461);
and U17021 (N_17021,N_15997,N_16409);
and U17022 (N_17022,N_16496,N_16241);
nor U17023 (N_17023,N_16648,N_15649);
and U17024 (N_17024,N_16664,N_15715);
nand U17025 (N_17025,N_16443,N_16474);
nand U17026 (N_17026,N_16775,N_16515);
and U17027 (N_17027,N_16660,N_15760);
nor U17028 (N_17028,N_16309,N_15779);
xnor U17029 (N_17029,N_16577,N_15601);
and U17030 (N_17030,N_16122,N_15953);
nor U17031 (N_17031,N_15946,N_16022);
and U17032 (N_17032,N_15844,N_15940);
or U17033 (N_17033,N_16142,N_15684);
xnor U17034 (N_17034,N_16504,N_15752);
or U17035 (N_17035,N_16392,N_16777);
nor U17036 (N_17036,N_16262,N_15709);
nand U17037 (N_17037,N_16029,N_16042);
nand U17038 (N_17038,N_16302,N_15879);
or U17039 (N_17039,N_16317,N_16587);
nand U17040 (N_17040,N_16535,N_16458);
nand U17041 (N_17041,N_16760,N_16637);
or U17042 (N_17042,N_16175,N_16150);
nand U17043 (N_17043,N_15893,N_16628);
nand U17044 (N_17044,N_16218,N_15929);
xor U17045 (N_17045,N_15787,N_16268);
xor U17046 (N_17046,N_16674,N_16143);
nor U17047 (N_17047,N_16509,N_15982);
or U17048 (N_17048,N_16305,N_15699);
or U17049 (N_17049,N_15968,N_16097);
xnor U17050 (N_17050,N_15988,N_15843);
or U17051 (N_17051,N_16117,N_16304);
nand U17052 (N_17052,N_16089,N_16371);
nor U17053 (N_17053,N_16662,N_16469);
nor U17054 (N_17054,N_16471,N_16148);
xor U17055 (N_17055,N_16276,N_15908);
nand U17056 (N_17056,N_16134,N_15923);
and U17057 (N_17057,N_15943,N_16727);
nor U17058 (N_17058,N_15965,N_15652);
and U17059 (N_17059,N_15859,N_16440);
or U17060 (N_17060,N_16704,N_15984);
and U17061 (N_17061,N_15976,N_16745);
nand U17062 (N_17062,N_16736,N_15757);
nand U17063 (N_17063,N_15620,N_16374);
and U17064 (N_17064,N_15763,N_16131);
xnor U17065 (N_17065,N_16690,N_15958);
or U17066 (N_17066,N_15841,N_16372);
and U17067 (N_17067,N_16179,N_16772);
nand U17068 (N_17068,N_16092,N_16764);
or U17069 (N_17069,N_16663,N_16717);
xnor U17070 (N_17070,N_16253,N_16162);
xnor U17071 (N_17071,N_16396,N_15678);
nand U17072 (N_17072,N_16470,N_15842);
nand U17073 (N_17073,N_16397,N_15901);
nor U17074 (N_17074,N_16019,N_16114);
and U17075 (N_17075,N_16778,N_16158);
nor U17076 (N_17076,N_15657,N_15885);
xnor U17077 (N_17077,N_16336,N_16537);
nand U17078 (N_17078,N_16382,N_16313);
or U17079 (N_17079,N_16129,N_16328);
xor U17080 (N_17080,N_16495,N_15998);
nand U17081 (N_17081,N_16406,N_16617);
xor U17082 (N_17082,N_16610,N_15606);
nand U17083 (N_17083,N_16188,N_16287);
or U17084 (N_17084,N_15640,N_16743);
or U17085 (N_17085,N_16482,N_15607);
nand U17086 (N_17086,N_16009,N_16799);
nand U17087 (N_17087,N_15897,N_15985);
nor U17088 (N_17088,N_15695,N_15661);
nand U17089 (N_17089,N_16367,N_16311);
and U17090 (N_17090,N_16578,N_16644);
xnor U17091 (N_17091,N_16419,N_15638);
nand U17092 (N_17092,N_16403,N_15848);
or U17093 (N_17093,N_16184,N_16400);
xnor U17094 (N_17094,N_16013,N_15670);
or U17095 (N_17095,N_15855,N_16088);
xor U17096 (N_17096,N_15886,N_16591);
nor U17097 (N_17097,N_16380,N_15711);
xnor U17098 (N_17098,N_15662,N_15600);
nor U17099 (N_17099,N_15615,N_15904);
nand U17100 (N_17100,N_16377,N_16215);
xor U17101 (N_17101,N_16235,N_15784);
nor U17102 (N_17102,N_16258,N_16781);
nand U17103 (N_17103,N_16220,N_15972);
xor U17104 (N_17104,N_15805,N_16604);
nor U17105 (N_17105,N_15890,N_16414);
and U17106 (N_17106,N_15739,N_15817);
nor U17107 (N_17107,N_16068,N_15705);
and U17108 (N_17108,N_16243,N_15914);
and U17109 (N_17109,N_16729,N_16405);
or U17110 (N_17110,N_16291,N_15840);
nand U17111 (N_17111,N_15623,N_16689);
or U17112 (N_17112,N_16531,N_15963);
nor U17113 (N_17113,N_15921,N_16228);
and U17114 (N_17114,N_15875,N_16032);
nand U17115 (N_17115,N_16060,N_15856);
and U17116 (N_17116,N_16750,N_15796);
and U17117 (N_17117,N_16732,N_16719);
xor U17118 (N_17118,N_16792,N_16118);
and U17119 (N_17119,N_16249,N_15957);
xnor U17120 (N_17120,N_16066,N_16416);
and U17121 (N_17121,N_16606,N_16127);
and U17122 (N_17122,N_16325,N_16602);
and U17123 (N_17123,N_16762,N_16739);
or U17124 (N_17124,N_15616,N_15837);
and U17125 (N_17125,N_15871,N_16023);
and U17126 (N_17126,N_16095,N_15839);
or U17127 (N_17127,N_16044,N_16116);
nand U17128 (N_17128,N_15690,N_16191);
or U17129 (N_17129,N_16500,N_16705);
and U17130 (N_17130,N_15643,N_16766);
nand U17131 (N_17131,N_16381,N_16102);
nand U17132 (N_17132,N_15942,N_15663);
or U17133 (N_17133,N_16389,N_15750);
or U17134 (N_17134,N_16770,N_15754);
nor U17135 (N_17135,N_16493,N_16387);
xnor U17136 (N_17136,N_16176,N_16508);
nand U17137 (N_17137,N_15745,N_16094);
and U17138 (N_17138,N_16542,N_15915);
xor U17139 (N_17139,N_16435,N_16137);
or U17140 (N_17140,N_16570,N_15999);
or U17141 (N_17141,N_16252,N_15917);
nand U17142 (N_17142,N_16180,N_16759);
nand U17143 (N_17143,N_15954,N_16748);
xnor U17144 (N_17144,N_16314,N_15983);
or U17145 (N_17145,N_16561,N_15906);
nand U17146 (N_17146,N_16072,N_16726);
and U17147 (N_17147,N_16572,N_15728);
and U17148 (N_17148,N_15706,N_16399);
xor U17149 (N_17149,N_16197,N_16055);
and U17150 (N_17150,N_16242,N_16774);
xnor U17151 (N_17151,N_16630,N_16185);
or U17152 (N_17152,N_16348,N_16590);
nand U17153 (N_17153,N_16710,N_16580);
xor U17154 (N_17154,N_15689,N_16684);
nand U17155 (N_17155,N_16269,N_16605);
or U17156 (N_17156,N_15650,N_15955);
nand U17157 (N_17157,N_16375,N_15604);
xor U17158 (N_17158,N_16783,N_16156);
nor U17159 (N_17159,N_15846,N_16310);
or U17160 (N_17160,N_16452,N_16699);
nor U17161 (N_17161,N_16263,N_15977);
or U17162 (N_17162,N_16098,N_16680);
xor U17163 (N_17163,N_15724,N_16512);
and U17164 (N_17164,N_16706,N_16126);
nor U17165 (N_17165,N_16299,N_16151);
xor U17166 (N_17166,N_16716,N_16703);
or U17167 (N_17167,N_16417,N_15639);
nand U17168 (N_17168,N_16445,N_15812);
nor U17169 (N_17169,N_16090,N_16420);
nor U17170 (N_17170,N_15956,N_16369);
or U17171 (N_17171,N_16431,N_16393);
nand U17172 (N_17172,N_16404,N_16360);
nand U17173 (N_17173,N_16128,N_16157);
or U17174 (N_17174,N_16523,N_16075);
or U17175 (N_17175,N_16564,N_16141);
xnor U17176 (N_17176,N_16692,N_16238);
nor U17177 (N_17177,N_16069,N_16236);
nor U17178 (N_17178,N_15726,N_16756);
and U17179 (N_17179,N_16323,N_16585);
xor U17180 (N_17180,N_15960,N_15964);
nand U17181 (N_17181,N_16178,N_15733);
and U17182 (N_17182,N_16145,N_16643);
nand U17183 (N_17183,N_15898,N_16483);
and U17184 (N_17184,N_15767,N_16616);
nand U17185 (N_17185,N_16084,N_16059);
nor U17186 (N_17186,N_16735,N_16106);
nand U17187 (N_17187,N_16625,N_16230);
and U17188 (N_17188,N_16669,N_16279);
nand U17189 (N_17189,N_16432,N_16079);
nor U17190 (N_17190,N_16460,N_15869);
or U17191 (N_17191,N_16008,N_16340);
xnor U17192 (N_17192,N_15831,N_16334);
nor U17193 (N_17193,N_15762,N_15919);
nand U17194 (N_17194,N_16593,N_16741);
nand U17195 (N_17195,N_16275,N_15845);
or U17196 (N_17196,N_15626,N_16033);
or U17197 (N_17197,N_16167,N_16707);
nand U17198 (N_17198,N_16749,N_15899);
and U17199 (N_17199,N_16609,N_16306);
and U17200 (N_17200,N_16347,N_16700);
or U17201 (N_17201,N_16659,N_16524);
xnor U17202 (N_17202,N_16246,N_16239);
nand U17203 (N_17203,N_16282,N_16086);
nor U17204 (N_17204,N_16011,N_16506);
xnor U17205 (N_17205,N_16161,N_16562);
and U17206 (N_17206,N_15691,N_16497);
or U17207 (N_17207,N_16083,N_16638);
and U17208 (N_17208,N_16712,N_16558);
nor U17209 (N_17209,N_15828,N_15734);
or U17210 (N_17210,N_16635,N_16231);
and U17211 (N_17211,N_15996,N_16110);
nand U17212 (N_17212,N_16254,N_16331);
or U17213 (N_17213,N_15962,N_16694);
xnor U17214 (N_17214,N_15803,N_16099);
xnor U17215 (N_17215,N_15632,N_16573);
nor U17216 (N_17216,N_16421,N_15891);
or U17217 (N_17217,N_15986,N_15768);
nor U17218 (N_17218,N_16549,N_16321);
xnor U17219 (N_17219,N_16245,N_16679);
nand U17220 (N_17220,N_16362,N_15685);
or U17221 (N_17221,N_16464,N_16626);
xor U17222 (N_17222,N_16554,N_16324);
or U17223 (N_17223,N_16183,N_16104);
and U17224 (N_17224,N_16209,N_15979);
nand U17225 (N_17225,N_16581,N_16466);
and U17226 (N_17226,N_16077,N_16017);
or U17227 (N_17227,N_16668,N_16227);
nor U17228 (N_17228,N_16676,N_16555);
and U17229 (N_17229,N_16219,N_16673);
xor U17230 (N_17230,N_15894,N_16758);
xnor U17231 (N_17231,N_16641,N_15822);
and U17232 (N_17232,N_15825,N_15838);
nand U17233 (N_17233,N_16769,N_16701);
nor U17234 (N_17234,N_16427,N_15806);
nor U17235 (N_17235,N_16341,N_15603);
and U17236 (N_17236,N_16358,N_16665);
nand U17237 (N_17237,N_16734,N_15612);
nand U17238 (N_17238,N_16492,N_15751);
xor U17239 (N_17239,N_16702,N_16085);
and U17240 (N_17240,N_16413,N_16488);
or U17241 (N_17241,N_15617,N_16266);
nand U17242 (N_17242,N_16165,N_16507);
nor U17243 (N_17243,N_15990,N_16115);
xnor U17244 (N_17244,N_16288,N_16240);
or U17245 (N_17245,N_15877,N_16015);
and U17246 (N_17246,N_16670,N_16260);
and U17247 (N_17247,N_16039,N_16170);
and U17248 (N_17248,N_16779,N_16429);
nor U17249 (N_17249,N_16541,N_16351);
xnor U17250 (N_17250,N_15989,N_16312);
nor U17251 (N_17251,N_15944,N_16651);
and U17252 (N_17252,N_16456,N_16049);
xnor U17253 (N_17253,N_15655,N_15870);
nand U17254 (N_17254,N_16206,N_16107);
and U17255 (N_17255,N_15697,N_16054);
or U17256 (N_17256,N_16439,N_16465);
or U17257 (N_17257,N_16026,N_15743);
nand U17258 (N_17258,N_16787,N_16248);
and U17259 (N_17259,N_16043,N_16192);
nand U17260 (N_17260,N_15949,N_15931);
xor U17261 (N_17261,N_15753,N_16332);
xnor U17262 (N_17262,N_15647,N_16057);
nor U17263 (N_17263,N_16067,N_16048);
nand U17264 (N_17264,N_16728,N_16761);
or U17265 (N_17265,N_15790,N_16037);
nor U17266 (N_17266,N_16453,N_16087);
nor U17267 (N_17267,N_15716,N_15974);
nand U17268 (N_17268,N_16672,N_15835);
nand U17269 (N_17269,N_15791,N_16686);
xnor U17270 (N_17270,N_15883,N_15688);
and U17271 (N_17271,N_15913,N_16344);
and U17272 (N_17272,N_16530,N_16633);
nand U17273 (N_17273,N_16061,N_16794);
nor U17274 (N_17274,N_16599,N_15712);
or U17275 (N_17275,N_16536,N_16058);
nand U17276 (N_17276,N_15687,N_15618);
nand U17277 (N_17277,N_16349,N_16595);
and U17278 (N_17278,N_15621,N_16544);
xnor U17279 (N_17279,N_15740,N_16345);
or U17280 (N_17280,N_15635,N_16751);
xnor U17281 (N_17281,N_16517,N_15759);
xor U17282 (N_17282,N_16451,N_16024);
xnor U17283 (N_17283,N_16647,N_16740);
and U17284 (N_17284,N_16271,N_16002);
xnor U17285 (N_17285,N_16486,N_15800);
nand U17286 (N_17286,N_16733,N_15613);
nand U17287 (N_17287,N_16721,N_16412);
or U17288 (N_17288,N_16010,N_16071);
or U17289 (N_17289,N_15622,N_15780);
nor U17290 (N_17290,N_16640,N_16394);
or U17291 (N_17291,N_15935,N_16285);
or U17292 (N_17292,N_16785,N_16021);
nand U17293 (N_17293,N_15666,N_15933);
nor U17294 (N_17294,N_16229,N_15720);
or U17295 (N_17295,N_15654,N_16065);
nand U17296 (N_17296,N_16226,N_16006);
nor U17297 (N_17297,N_15809,N_16194);
nor U17298 (N_17298,N_16548,N_15653);
xnor U17299 (N_17299,N_15658,N_16234);
and U17300 (N_17300,N_16278,N_15713);
and U17301 (N_17301,N_16050,N_16563);
xor U17302 (N_17302,N_16356,N_15683);
and U17303 (N_17303,N_15749,N_16612);
and U17304 (N_17304,N_16355,N_16320);
or U17305 (N_17305,N_16667,N_16035);
xor U17306 (N_17306,N_16487,N_15772);
and U17307 (N_17307,N_16169,N_15646);
and U17308 (N_17308,N_16182,N_15939);
nor U17309 (N_17309,N_16337,N_16080);
xor U17310 (N_17310,N_15912,N_16053);
xor U17311 (N_17311,N_16788,N_16624);
nor U17312 (N_17312,N_15631,N_15925);
and U17313 (N_17313,N_15807,N_16518);
or U17314 (N_17314,N_15676,N_16398);
nor U17315 (N_17315,N_16619,N_16546);
xnor U17316 (N_17316,N_15781,N_15677);
or U17317 (N_17317,N_16678,N_16467);
nor U17318 (N_17318,N_16526,N_16485);
or U17319 (N_17319,N_15708,N_16425);
or U17320 (N_17320,N_15833,N_16683);
nor U17321 (N_17321,N_15627,N_15851);
and U17322 (N_17322,N_16140,N_15667);
and U17323 (N_17323,N_15675,N_15852);
xnor U17324 (N_17324,N_16177,N_15924);
or U17325 (N_17325,N_16073,N_16295);
and U17326 (N_17326,N_15669,N_15629);
xor U17327 (N_17327,N_16447,N_16265);
xnor U17328 (N_17328,N_16653,N_16111);
or U17329 (N_17329,N_15872,N_15602);
nor U17330 (N_17330,N_16489,N_16298);
nor U17331 (N_17331,N_15920,N_16677);
or U17332 (N_17332,N_16790,N_16174);
or U17333 (N_17333,N_16130,N_16052);
or U17334 (N_17334,N_15884,N_15764);
xor U17335 (N_17335,N_16484,N_16529);
nand U17336 (N_17336,N_16379,N_16571);
xor U17337 (N_17337,N_16410,N_15830);
or U17338 (N_17338,N_16041,N_15783);
nor U17339 (N_17339,N_16171,N_16036);
or U17340 (N_17340,N_15633,N_16795);
or U17341 (N_17341,N_16798,N_16257);
xnor U17342 (N_17342,N_16289,N_16046);
xnor U17343 (N_17343,N_15624,N_15738);
or U17344 (N_17344,N_16553,N_15823);
or U17345 (N_17345,N_15948,N_16211);
xnor U17346 (N_17346,N_16620,N_16133);
and U17347 (N_17347,N_16201,N_16001);
nor U17348 (N_17348,N_16582,N_15742);
nand U17349 (N_17349,N_16222,N_16426);
and U17350 (N_17350,N_16738,N_16681);
nand U17351 (N_17351,N_15773,N_15737);
and U17352 (N_17352,N_15941,N_15821);
and U17353 (N_17353,N_15756,N_16286);
and U17354 (N_17354,N_15700,N_15863);
and U17355 (N_17355,N_16768,N_16632);
and U17356 (N_17356,N_16000,N_16540);
or U17357 (N_17357,N_15907,N_16296);
xor U17358 (N_17358,N_16444,N_16713);
or U17359 (N_17359,N_16202,N_15770);
nor U17360 (N_17360,N_16338,N_15795);
or U17361 (N_17361,N_16731,N_16502);
xor U17362 (N_17362,N_15971,N_15819);
or U17363 (N_17363,N_16292,N_15722);
nor U17364 (N_17364,N_15834,N_16172);
nor U17365 (N_17365,N_15991,N_15701);
or U17366 (N_17366,N_15994,N_16449);
or U17367 (N_17367,N_16730,N_16722);
or U17368 (N_17368,N_15934,N_16693);
nand U17369 (N_17369,N_15744,N_16646);
xnor U17370 (N_17370,N_16539,N_16438);
or U17371 (N_17371,N_15642,N_16611);
nor U17372 (N_17372,N_16522,N_16401);
nand U17373 (N_17373,N_16189,N_16533);
nor U17374 (N_17374,N_15900,N_16363);
nand U17375 (N_17375,N_16267,N_16203);
nor U17376 (N_17376,N_16613,N_16494);
nand U17377 (N_17377,N_16198,N_15938);
and U17378 (N_17378,N_16007,N_16671);
nor U17379 (N_17379,N_15719,N_16754);
xnor U17380 (N_17380,N_16652,N_16318);
or U17381 (N_17381,N_16557,N_15725);
nor U17382 (N_17382,N_16004,N_16378);
or U17383 (N_17383,N_15847,N_16031);
and U17384 (N_17384,N_15860,N_16365);
nor U17385 (N_17385,N_16565,N_16747);
xor U17386 (N_17386,N_15922,N_16199);
or U17387 (N_17387,N_16217,N_16025);
nand U17388 (N_17388,N_16124,N_15874);
nor U17389 (N_17389,N_16062,N_15947);
nor U17390 (N_17390,N_16064,N_16159);
and U17391 (N_17391,N_16560,N_16650);
or U17392 (N_17392,N_16168,N_15853);
xor U17393 (N_17393,N_16415,N_15755);
nor U17394 (N_17394,N_15858,N_16691);
nand U17395 (N_17395,N_16436,N_15882);
and U17396 (N_17396,N_16715,N_15798);
xnor U17397 (N_17397,N_16428,N_16765);
nand U17398 (N_17398,N_16301,N_16685);
nor U17399 (N_17399,N_16101,N_16028);
nor U17400 (N_17400,N_16197,N_16219);
and U17401 (N_17401,N_15853,N_16670);
and U17402 (N_17402,N_15709,N_16693);
or U17403 (N_17403,N_15645,N_15749);
and U17404 (N_17404,N_15936,N_15741);
nor U17405 (N_17405,N_16046,N_15908);
nand U17406 (N_17406,N_16588,N_16102);
and U17407 (N_17407,N_16226,N_16129);
and U17408 (N_17408,N_16490,N_16065);
or U17409 (N_17409,N_16047,N_16703);
nor U17410 (N_17410,N_16644,N_16037);
nand U17411 (N_17411,N_16747,N_16098);
nand U17412 (N_17412,N_16625,N_16767);
nand U17413 (N_17413,N_16069,N_16279);
or U17414 (N_17414,N_16180,N_16498);
or U17415 (N_17415,N_16637,N_16231);
or U17416 (N_17416,N_16327,N_16371);
nor U17417 (N_17417,N_16064,N_16615);
or U17418 (N_17418,N_16640,N_15799);
nor U17419 (N_17419,N_15795,N_16138);
xnor U17420 (N_17420,N_15682,N_15912);
and U17421 (N_17421,N_16589,N_16267);
xor U17422 (N_17422,N_16650,N_15804);
or U17423 (N_17423,N_15940,N_15618);
xnor U17424 (N_17424,N_15600,N_15711);
nor U17425 (N_17425,N_15753,N_16347);
or U17426 (N_17426,N_16788,N_16095);
nor U17427 (N_17427,N_16528,N_16577);
nand U17428 (N_17428,N_16779,N_16507);
or U17429 (N_17429,N_16072,N_16190);
and U17430 (N_17430,N_16463,N_16173);
nand U17431 (N_17431,N_16403,N_16143);
or U17432 (N_17432,N_16670,N_16564);
nor U17433 (N_17433,N_16307,N_16184);
and U17434 (N_17434,N_16023,N_15953);
xnor U17435 (N_17435,N_15750,N_16639);
nand U17436 (N_17436,N_15866,N_16013);
xnor U17437 (N_17437,N_16117,N_15913);
nor U17438 (N_17438,N_15915,N_16551);
nand U17439 (N_17439,N_16637,N_15745);
and U17440 (N_17440,N_15716,N_15956);
nand U17441 (N_17441,N_15806,N_15620);
and U17442 (N_17442,N_15739,N_15731);
nand U17443 (N_17443,N_16649,N_15760);
nor U17444 (N_17444,N_15775,N_15754);
or U17445 (N_17445,N_15969,N_15739);
nand U17446 (N_17446,N_15778,N_16052);
xnor U17447 (N_17447,N_16630,N_15927);
nor U17448 (N_17448,N_16558,N_15746);
or U17449 (N_17449,N_16184,N_15898);
or U17450 (N_17450,N_15790,N_15743);
xnor U17451 (N_17451,N_16322,N_16303);
xor U17452 (N_17452,N_16302,N_15811);
xor U17453 (N_17453,N_15957,N_16442);
xor U17454 (N_17454,N_16380,N_16045);
and U17455 (N_17455,N_15953,N_15817);
nor U17456 (N_17456,N_15822,N_15872);
nand U17457 (N_17457,N_15754,N_16133);
and U17458 (N_17458,N_16091,N_15972);
and U17459 (N_17459,N_15934,N_16485);
xnor U17460 (N_17460,N_16378,N_15731);
xor U17461 (N_17461,N_16248,N_16241);
and U17462 (N_17462,N_16618,N_16793);
nor U17463 (N_17463,N_15962,N_16059);
nor U17464 (N_17464,N_16085,N_16473);
nor U17465 (N_17465,N_15982,N_15806);
nand U17466 (N_17466,N_16013,N_15965);
xor U17467 (N_17467,N_15945,N_16096);
and U17468 (N_17468,N_16351,N_15609);
or U17469 (N_17469,N_15986,N_16062);
nand U17470 (N_17470,N_16159,N_16033);
nand U17471 (N_17471,N_16060,N_15790);
nor U17472 (N_17472,N_16237,N_15854);
xor U17473 (N_17473,N_16569,N_15656);
xnor U17474 (N_17474,N_16064,N_15652);
or U17475 (N_17475,N_15796,N_16126);
nor U17476 (N_17476,N_15939,N_15853);
or U17477 (N_17477,N_16626,N_16433);
and U17478 (N_17478,N_16199,N_16211);
or U17479 (N_17479,N_16766,N_16057);
nor U17480 (N_17480,N_16106,N_15829);
and U17481 (N_17481,N_16627,N_15761);
or U17482 (N_17482,N_16499,N_16008);
or U17483 (N_17483,N_16320,N_15957);
or U17484 (N_17484,N_16003,N_16217);
nand U17485 (N_17485,N_16359,N_16314);
nand U17486 (N_17486,N_16139,N_15712);
and U17487 (N_17487,N_16419,N_16337);
xor U17488 (N_17488,N_16388,N_15870);
or U17489 (N_17489,N_16388,N_15900);
and U17490 (N_17490,N_15683,N_15828);
xnor U17491 (N_17491,N_15730,N_16410);
and U17492 (N_17492,N_16369,N_16452);
xnor U17493 (N_17493,N_15972,N_16646);
nand U17494 (N_17494,N_16121,N_15994);
or U17495 (N_17495,N_16545,N_15770);
nand U17496 (N_17496,N_16774,N_15960);
nor U17497 (N_17497,N_16317,N_16038);
xnor U17498 (N_17498,N_16785,N_16655);
nand U17499 (N_17499,N_16074,N_16344);
nor U17500 (N_17500,N_16732,N_16061);
nor U17501 (N_17501,N_15897,N_15653);
nand U17502 (N_17502,N_16415,N_16148);
nor U17503 (N_17503,N_16797,N_16431);
nor U17504 (N_17504,N_16043,N_16375);
nor U17505 (N_17505,N_16412,N_16308);
nand U17506 (N_17506,N_15786,N_16371);
xnor U17507 (N_17507,N_16750,N_16731);
nor U17508 (N_17508,N_16133,N_16658);
xnor U17509 (N_17509,N_16057,N_15837);
xor U17510 (N_17510,N_15762,N_15942);
or U17511 (N_17511,N_16138,N_16617);
or U17512 (N_17512,N_15702,N_16759);
nor U17513 (N_17513,N_15687,N_15682);
or U17514 (N_17514,N_16706,N_16287);
nand U17515 (N_17515,N_15891,N_16790);
nand U17516 (N_17516,N_16343,N_16084);
and U17517 (N_17517,N_15652,N_15832);
nand U17518 (N_17518,N_16479,N_16678);
nand U17519 (N_17519,N_16613,N_15653);
nand U17520 (N_17520,N_15692,N_16537);
nor U17521 (N_17521,N_15953,N_15675);
nor U17522 (N_17522,N_16737,N_16291);
nor U17523 (N_17523,N_15767,N_16285);
xnor U17524 (N_17524,N_16443,N_16275);
and U17525 (N_17525,N_16204,N_16201);
and U17526 (N_17526,N_15743,N_15638);
and U17527 (N_17527,N_15745,N_16398);
and U17528 (N_17528,N_16449,N_15629);
xor U17529 (N_17529,N_15636,N_16319);
xor U17530 (N_17530,N_16031,N_16134);
nor U17531 (N_17531,N_16699,N_15880);
nand U17532 (N_17532,N_15765,N_16196);
or U17533 (N_17533,N_16344,N_15828);
and U17534 (N_17534,N_16101,N_16387);
or U17535 (N_17535,N_15843,N_16656);
xnor U17536 (N_17536,N_16362,N_16277);
and U17537 (N_17537,N_16130,N_16678);
xnor U17538 (N_17538,N_16405,N_15939);
nand U17539 (N_17539,N_16429,N_16076);
nor U17540 (N_17540,N_16571,N_15624);
and U17541 (N_17541,N_16633,N_16787);
xnor U17542 (N_17542,N_15655,N_15703);
nand U17543 (N_17543,N_16637,N_16751);
and U17544 (N_17544,N_15792,N_15704);
and U17545 (N_17545,N_16254,N_15629);
xor U17546 (N_17546,N_16218,N_16428);
nand U17547 (N_17547,N_15843,N_15841);
nand U17548 (N_17548,N_16681,N_15659);
xor U17549 (N_17549,N_16443,N_16352);
and U17550 (N_17550,N_15650,N_16685);
nand U17551 (N_17551,N_16373,N_15601);
xnor U17552 (N_17552,N_16385,N_16719);
nor U17553 (N_17553,N_16626,N_16365);
and U17554 (N_17554,N_15732,N_15910);
xor U17555 (N_17555,N_16131,N_16072);
nand U17556 (N_17556,N_15978,N_16451);
nor U17557 (N_17557,N_16600,N_16063);
and U17558 (N_17558,N_15756,N_15652);
nand U17559 (N_17559,N_15931,N_15667);
and U17560 (N_17560,N_16530,N_16484);
and U17561 (N_17561,N_15880,N_15842);
and U17562 (N_17562,N_16037,N_16083);
nand U17563 (N_17563,N_15714,N_16029);
nor U17564 (N_17564,N_16317,N_15890);
nand U17565 (N_17565,N_16025,N_16478);
and U17566 (N_17566,N_16322,N_16447);
nor U17567 (N_17567,N_16326,N_16784);
or U17568 (N_17568,N_16203,N_16101);
or U17569 (N_17569,N_16417,N_15845);
xnor U17570 (N_17570,N_16072,N_15665);
xor U17571 (N_17571,N_16104,N_16300);
xnor U17572 (N_17572,N_16532,N_16092);
or U17573 (N_17573,N_15878,N_16384);
xnor U17574 (N_17574,N_15694,N_16495);
nor U17575 (N_17575,N_15758,N_15677);
xnor U17576 (N_17576,N_16213,N_16653);
nor U17577 (N_17577,N_16408,N_16331);
nand U17578 (N_17578,N_16761,N_16158);
and U17579 (N_17579,N_15873,N_16723);
and U17580 (N_17580,N_15673,N_15978);
nand U17581 (N_17581,N_16470,N_16292);
nor U17582 (N_17582,N_15734,N_16160);
or U17583 (N_17583,N_15802,N_16453);
nor U17584 (N_17584,N_15607,N_16483);
xor U17585 (N_17585,N_16273,N_16202);
xnor U17586 (N_17586,N_15608,N_16799);
nor U17587 (N_17587,N_15830,N_16244);
nor U17588 (N_17588,N_15739,N_15638);
nand U17589 (N_17589,N_16772,N_16446);
nand U17590 (N_17590,N_15823,N_15910);
nor U17591 (N_17591,N_15768,N_16656);
nand U17592 (N_17592,N_15606,N_16166);
nor U17593 (N_17593,N_16491,N_16469);
and U17594 (N_17594,N_15986,N_16069);
nand U17595 (N_17595,N_16309,N_16417);
nand U17596 (N_17596,N_15869,N_16534);
and U17597 (N_17597,N_16085,N_16382);
nor U17598 (N_17598,N_16384,N_15732);
and U17599 (N_17599,N_16730,N_16519);
nand U17600 (N_17600,N_16094,N_16309);
or U17601 (N_17601,N_16498,N_16077);
and U17602 (N_17602,N_15976,N_16178);
or U17603 (N_17603,N_16071,N_15626);
and U17604 (N_17604,N_16274,N_15878);
xor U17605 (N_17605,N_16741,N_15700);
nand U17606 (N_17606,N_16527,N_16283);
xor U17607 (N_17607,N_15732,N_15896);
nand U17608 (N_17608,N_16248,N_16060);
nand U17609 (N_17609,N_16769,N_15875);
nor U17610 (N_17610,N_15798,N_16775);
nor U17611 (N_17611,N_15885,N_16170);
nor U17612 (N_17612,N_16627,N_16469);
and U17613 (N_17613,N_15987,N_15984);
nor U17614 (N_17614,N_15820,N_15614);
or U17615 (N_17615,N_15821,N_16721);
or U17616 (N_17616,N_16710,N_16208);
and U17617 (N_17617,N_16209,N_15960);
xor U17618 (N_17618,N_16583,N_15902);
nand U17619 (N_17619,N_16783,N_16771);
or U17620 (N_17620,N_16703,N_15677);
xnor U17621 (N_17621,N_16616,N_15698);
and U17622 (N_17622,N_15880,N_16637);
nand U17623 (N_17623,N_16381,N_16632);
xor U17624 (N_17624,N_15611,N_16697);
nand U17625 (N_17625,N_16191,N_15935);
xor U17626 (N_17626,N_15864,N_16332);
xor U17627 (N_17627,N_15687,N_15916);
nand U17628 (N_17628,N_15752,N_16647);
nand U17629 (N_17629,N_15917,N_16004);
xnor U17630 (N_17630,N_16032,N_16230);
and U17631 (N_17631,N_16122,N_16345);
or U17632 (N_17632,N_15810,N_16406);
xnor U17633 (N_17633,N_15908,N_16054);
nor U17634 (N_17634,N_16254,N_16233);
or U17635 (N_17635,N_16530,N_16123);
or U17636 (N_17636,N_15740,N_15710);
or U17637 (N_17637,N_16487,N_16354);
nand U17638 (N_17638,N_16383,N_15755);
nor U17639 (N_17639,N_16143,N_16545);
or U17640 (N_17640,N_16485,N_15665);
and U17641 (N_17641,N_15821,N_16727);
or U17642 (N_17642,N_16305,N_16592);
nand U17643 (N_17643,N_16745,N_15779);
or U17644 (N_17644,N_15845,N_16284);
nor U17645 (N_17645,N_16751,N_16500);
xor U17646 (N_17646,N_15644,N_16342);
nor U17647 (N_17647,N_16132,N_15979);
or U17648 (N_17648,N_16425,N_15690);
and U17649 (N_17649,N_16322,N_16755);
xnor U17650 (N_17650,N_15698,N_16768);
nor U17651 (N_17651,N_16194,N_16495);
or U17652 (N_17652,N_15779,N_16623);
xor U17653 (N_17653,N_16144,N_15631);
xnor U17654 (N_17654,N_15786,N_16676);
nand U17655 (N_17655,N_16775,N_16101);
nand U17656 (N_17656,N_16548,N_15794);
or U17657 (N_17657,N_16340,N_15651);
or U17658 (N_17658,N_16266,N_16058);
and U17659 (N_17659,N_16309,N_15972);
xnor U17660 (N_17660,N_16159,N_15936);
and U17661 (N_17661,N_15898,N_16428);
nor U17662 (N_17662,N_15646,N_16499);
nand U17663 (N_17663,N_16364,N_16059);
nand U17664 (N_17664,N_16789,N_16041);
xnor U17665 (N_17665,N_15782,N_16466);
or U17666 (N_17666,N_16250,N_16768);
and U17667 (N_17667,N_15710,N_16602);
or U17668 (N_17668,N_15938,N_16539);
or U17669 (N_17669,N_16660,N_15692);
and U17670 (N_17670,N_15862,N_15968);
nor U17671 (N_17671,N_15841,N_15698);
xnor U17672 (N_17672,N_15980,N_16269);
and U17673 (N_17673,N_15765,N_16537);
nand U17674 (N_17674,N_15620,N_16303);
xnor U17675 (N_17675,N_15695,N_15836);
nor U17676 (N_17676,N_15724,N_15870);
nor U17677 (N_17677,N_16703,N_16470);
or U17678 (N_17678,N_16525,N_16601);
or U17679 (N_17679,N_15671,N_15822);
nand U17680 (N_17680,N_15991,N_15923);
xnor U17681 (N_17681,N_15935,N_16192);
nor U17682 (N_17682,N_16489,N_16589);
and U17683 (N_17683,N_15846,N_16457);
and U17684 (N_17684,N_15845,N_15864);
xnor U17685 (N_17685,N_16063,N_16207);
nand U17686 (N_17686,N_15835,N_16167);
or U17687 (N_17687,N_16133,N_16656);
nor U17688 (N_17688,N_15859,N_16083);
or U17689 (N_17689,N_16581,N_15607);
xnor U17690 (N_17690,N_16211,N_15922);
nor U17691 (N_17691,N_16016,N_15653);
and U17692 (N_17692,N_15703,N_15995);
xnor U17693 (N_17693,N_15625,N_16511);
and U17694 (N_17694,N_15674,N_15955);
xnor U17695 (N_17695,N_16271,N_16150);
and U17696 (N_17696,N_16012,N_16310);
xor U17697 (N_17697,N_16707,N_16512);
nand U17698 (N_17698,N_15754,N_16589);
nor U17699 (N_17699,N_16475,N_16204);
nand U17700 (N_17700,N_16035,N_15822);
nor U17701 (N_17701,N_16052,N_16184);
nand U17702 (N_17702,N_15892,N_16263);
xnor U17703 (N_17703,N_16161,N_15902);
and U17704 (N_17704,N_16525,N_15971);
nand U17705 (N_17705,N_15631,N_16201);
xnor U17706 (N_17706,N_15940,N_16132);
xor U17707 (N_17707,N_15704,N_16009);
or U17708 (N_17708,N_16065,N_16786);
nand U17709 (N_17709,N_16661,N_16715);
xnor U17710 (N_17710,N_16687,N_16521);
nor U17711 (N_17711,N_15880,N_15995);
nor U17712 (N_17712,N_16125,N_16173);
and U17713 (N_17713,N_16324,N_15678);
or U17714 (N_17714,N_15739,N_16360);
xnor U17715 (N_17715,N_16207,N_16431);
xor U17716 (N_17716,N_16091,N_16332);
and U17717 (N_17717,N_16768,N_16252);
or U17718 (N_17718,N_15601,N_16038);
nand U17719 (N_17719,N_15680,N_16126);
nor U17720 (N_17720,N_16402,N_16001);
and U17721 (N_17721,N_15684,N_16414);
nand U17722 (N_17722,N_15799,N_16776);
nor U17723 (N_17723,N_15852,N_16360);
nor U17724 (N_17724,N_15854,N_15715);
and U17725 (N_17725,N_15620,N_16737);
or U17726 (N_17726,N_16456,N_15927);
or U17727 (N_17727,N_16353,N_16450);
nor U17728 (N_17728,N_15882,N_15736);
nand U17729 (N_17729,N_16192,N_15875);
xnor U17730 (N_17730,N_16792,N_16554);
xnor U17731 (N_17731,N_16217,N_15873);
nor U17732 (N_17732,N_16035,N_16781);
nand U17733 (N_17733,N_16080,N_16422);
nor U17734 (N_17734,N_16094,N_15822);
or U17735 (N_17735,N_15679,N_15692);
nor U17736 (N_17736,N_16319,N_16166);
nor U17737 (N_17737,N_16133,N_15641);
nor U17738 (N_17738,N_16693,N_16143);
or U17739 (N_17739,N_15961,N_15645);
or U17740 (N_17740,N_16344,N_16120);
nand U17741 (N_17741,N_15658,N_16194);
xor U17742 (N_17742,N_16246,N_15920);
xor U17743 (N_17743,N_16299,N_16655);
nor U17744 (N_17744,N_15629,N_15949);
nor U17745 (N_17745,N_16294,N_16780);
or U17746 (N_17746,N_15690,N_15762);
nand U17747 (N_17747,N_16653,N_15942);
xor U17748 (N_17748,N_16373,N_16110);
or U17749 (N_17749,N_15895,N_16005);
xor U17750 (N_17750,N_16284,N_15874);
and U17751 (N_17751,N_16521,N_15660);
or U17752 (N_17752,N_15866,N_15729);
nor U17753 (N_17753,N_16444,N_15721);
nor U17754 (N_17754,N_16567,N_16759);
nand U17755 (N_17755,N_16502,N_16541);
or U17756 (N_17756,N_16503,N_16733);
or U17757 (N_17757,N_16561,N_16685);
and U17758 (N_17758,N_16059,N_16717);
nor U17759 (N_17759,N_16650,N_15614);
nand U17760 (N_17760,N_16085,N_16745);
nor U17761 (N_17761,N_16292,N_15626);
nor U17762 (N_17762,N_16257,N_16132);
or U17763 (N_17763,N_16069,N_16652);
xnor U17764 (N_17764,N_15873,N_15913);
nor U17765 (N_17765,N_16736,N_16076);
xnor U17766 (N_17766,N_16384,N_16192);
nand U17767 (N_17767,N_16354,N_15834);
xor U17768 (N_17768,N_15969,N_16208);
nor U17769 (N_17769,N_16587,N_16055);
nor U17770 (N_17770,N_16580,N_16010);
xnor U17771 (N_17771,N_16125,N_16527);
nand U17772 (N_17772,N_16468,N_16110);
and U17773 (N_17773,N_16102,N_15768);
and U17774 (N_17774,N_16749,N_16012);
or U17775 (N_17775,N_16474,N_16082);
or U17776 (N_17776,N_16303,N_15603);
xor U17777 (N_17777,N_16034,N_15750);
and U17778 (N_17778,N_16390,N_16471);
xor U17779 (N_17779,N_16399,N_16660);
nand U17780 (N_17780,N_16562,N_16398);
xnor U17781 (N_17781,N_15872,N_16026);
and U17782 (N_17782,N_16139,N_15773);
nand U17783 (N_17783,N_16385,N_15917);
and U17784 (N_17784,N_16449,N_16138);
or U17785 (N_17785,N_15856,N_16136);
nand U17786 (N_17786,N_16220,N_15736);
or U17787 (N_17787,N_16266,N_15812);
nor U17788 (N_17788,N_15702,N_16252);
nor U17789 (N_17789,N_16256,N_16131);
xnor U17790 (N_17790,N_15717,N_16271);
xnor U17791 (N_17791,N_15869,N_15858);
xor U17792 (N_17792,N_15825,N_15755);
nand U17793 (N_17793,N_16536,N_16480);
or U17794 (N_17794,N_16742,N_16731);
nand U17795 (N_17795,N_15989,N_15906);
nor U17796 (N_17796,N_15715,N_15645);
or U17797 (N_17797,N_16474,N_16304);
xnor U17798 (N_17798,N_16058,N_16199);
xor U17799 (N_17799,N_16222,N_16522);
or U17800 (N_17800,N_16590,N_16119);
or U17801 (N_17801,N_15609,N_16456);
nor U17802 (N_17802,N_16286,N_16684);
xor U17803 (N_17803,N_15861,N_16033);
nand U17804 (N_17804,N_16159,N_16002);
xor U17805 (N_17805,N_15907,N_16371);
nor U17806 (N_17806,N_15687,N_15883);
nor U17807 (N_17807,N_16205,N_15691);
or U17808 (N_17808,N_16581,N_16073);
nand U17809 (N_17809,N_16713,N_15830);
or U17810 (N_17810,N_15926,N_15660);
xnor U17811 (N_17811,N_15735,N_16309);
and U17812 (N_17812,N_16077,N_15653);
xor U17813 (N_17813,N_16725,N_16779);
nand U17814 (N_17814,N_16165,N_16187);
xnor U17815 (N_17815,N_16642,N_16146);
or U17816 (N_17816,N_16765,N_15693);
nand U17817 (N_17817,N_16002,N_15868);
nor U17818 (N_17818,N_15739,N_16481);
nand U17819 (N_17819,N_16241,N_15993);
and U17820 (N_17820,N_16358,N_15960);
nor U17821 (N_17821,N_16620,N_16257);
nor U17822 (N_17822,N_15939,N_15931);
nand U17823 (N_17823,N_16741,N_16148);
or U17824 (N_17824,N_15683,N_16375);
nor U17825 (N_17825,N_16735,N_16269);
and U17826 (N_17826,N_15745,N_15688);
and U17827 (N_17827,N_15801,N_16288);
nand U17828 (N_17828,N_16263,N_16012);
xor U17829 (N_17829,N_16262,N_15769);
nand U17830 (N_17830,N_16466,N_16357);
or U17831 (N_17831,N_16776,N_15798);
xor U17832 (N_17832,N_16411,N_16553);
nand U17833 (N_17833,N_16409,N_15851);
nor U17834 (N_17834,N_15671,N_16508);
xnor U17835 (N_17835,N_15982,N_16396);
or U17836 (N_17836,N_15613,N_15919);
or U17837 (N_17837,N_16018,N_16461);
xnor U17838 (N_17838,N_16578,N_15685);
nand U17839 (N_17839,N_15849,N_16432);
and U17840 (N_17840,N_16305,N_16259);
or U17841 (N_17841,N_15956,N_16095);
xor U17842 (N_17842,N_15961,N_16341);
nand U17843 (N_17843,N_15966,N_16611);
or U17844 (N_17844,N_16306,N_15853);
nand U17845 (N_17845,N_16256,N_15860);
xnor U17846 (N_17846,N_16784,N_16082);
or U17847 (N_17847,N_16656,N_16349);
nor U17848 (N_17848,N_16534,N_16048);
nand U17849 (N_17849,N_16788,N_15848);
or U17850 (N_17850,N_16359,N_16735);
or U17851 (N_17851,N_16462,N_15829);
or U17852 (N_17852,N_16234,N_16718);
and U17853 (N_17853,N_16764,N_16411);
or U17854 (N_17854,N_16462,N_15935);
nor U17855 (N_17855,N_16363,N_15872);
nor U17856 (N_17856,N_16003,N_16359);
nor U17857 (N_17857,N_16183,N_16396);
or U17858 (N_17858,N_15684,N_15753);
nor U17859 (N_17859,N_16266,N_16230);
or U17860 (N_17860,N_16041,N_16695);
xor U17861 (N_17861,N_16046,N_16747);
nor U17862 (N_17862,N_16656,N_15740);
xor U17863 (N_17863,N_15663,N_16484);
xor U17864 (N_17864,N_16751,N_15697);
nor U17865 (N_17865,N_16721,N_16700);
and U17866 (N_17866,N_16432,N_16414);
nor U17867 (N_17867,N_16678,N_15826);
and U17868 (N_17868,N_16273,N_16417);
xor U17869 (N_17869,N_15959,N_15636);
or U17870 (N_17870,N_16571,N_15620);
nand U17871 (N_17871,N_15667,N_15683);
nor U17872 (N_17872,N_16652,N_16332);
nand U17873 (N_17873,N_16688,N_16201);
or U17874 (N_17874,N_16639,N_15736);
nand U17875 (N_17875,N_16563,N_16464);
nand U17876 (N_17876,N_15738,N_16037);
and U17877 (N_17877,N_16514,N_16473);
and U17878 (N_17878,N_16058,N_16436);
nand U17879 (N_17879,N_15620,N_16404);
xnor U17880 (N_17880,N_15638,N_16417);
nor U17881 (N_17881,N_15657,N_16593);
xor U17882 (N_17882,N_16700,N_15802);
or U17883 (N_17883,N_16215,N_16497);
xnor U17884 (N_17884,N_15912,N_16778);
or U17885 (N_17885,N_15857,N_16286);
and U17886 (N_17886,N_16548,N_16732);
or U17887 (N_17887,N_16174,N_15979);
nand U17888 (N_17888,N_15685,N_16272);
and U17889 (N_17889,N_15853,N_16108);
and U17890 (N_17890,N_16243,N_15880);
or U17891 (N_17891,N_16312,N_16131);
or U17892 (N_17892,N_15675,N_16644);
nor U17893 (N_17893,N_15933,N_16570);
and U17894 (N_17894,N_16374,N_16799);
xor U17895 (N_17895,N_16496,N_16066);
or U17896 (N_17896,N_16354,N_16707);
or U17897 (N_17897,N_16319,N_16165);
nand U17898 (N_17898,N_16356,N_16459);
nand U17899 (N_17899,N_16092,N_16744);
xor U17900 (N_17900,N_15721,N_15718);
nand U17901 (N_17901,N_15728,N_16717);
nand U17902 (N_17902,N_16457,N_16389);
nor U17903 (N_17903,N_15936,N_16058);
xor U17904 (N_17904,N_15781,N_16227);
xnor U17905 (N_17905,N_16301,N_15789);
xnor U17906 (N_17906,N_16630,N_15944);
and U17907 (N_17907,N_16211,N_16446);
and U17908 (N_17908,N_16738,N_16424);
nand U17909 (N_17909,N_15760,N_15685);
nand U17910 (N_17910,N_15684,N_15841);
and U17911 (N_17911,N_16369,N_16212);
nand U17912 (N_17912,N_16726,N_16501);
nand U17913 (N_17913,N_16561,N_16364);
nand U17914 (N_17914,N_16490,N_16528);
or U17915 (N_17915,N_16633,N_15738);
nor U17916 (N_17916,N_15616,N_15809);
or U17917 (N_17917,N_16427,N_16442);
or U17918 (N_17918,N_15720,N_16337);
nor U17919 (N_17919,N_15681,N_15634);
xor U17920 (N_17920,N_15696,N_16395);
and U17921 (N_17921,N_15618,N_16657);
nor U17922 (N_17922,N_16087,N_15714);
xnor U17923 (N_17923,N_15821,N_16423);
xor U17924 (N_17924,N_15955,N_16325);
and U17925 (N_17925,N_16590,N_16409);
or U17926 (N_17926,N_16510,N_15939);
and U17927 (N_17927,N_16668,N_16565);
nand U17928 (N_17928,N_15922,N_15727);
nand U17929 (N_17929,N_15640,N_16644);
or U17930 (N_17930,N_16189,N_15854);
and U17931 (N_17931,N_16579,N_16798);
and U17932 (N_17932,N_16583,N_16405);
nor U17933 (N_17933,N_16732,N_16019);
or U17934 (N_17934,N_16345,N_16724);
or U17935 (N_17935,N_16452,N_15892);
xor U17936 (N_17936,N_16373,N_16138);
xor U17937 (N_17937,N_16043,N_16074);
and U17938 (N_17938,N_16391,N_16037);
nand U17939 (N_17939,N_15625,N_16407);
or U17940 (N_17940,N_16481,N_16434);
or U17941 (N_17941,N_16368,N_15940);
and U17942 (N_17942,N_16329,N_16082);
and U17943 (N_17943,N_16557,N_15858);
nor U17944 (N_17944,N_15721,N_16073);
xor U17945 (N_17945,N_16760,N_15664);
nand U17946 (N_17946,N_16538,N_15980);
or U17947 (N_17947,N_15788,N_15768);
nand U17948 (N_17948,N_16010,N_15655);
or U17949 (N_17949,N_16400,N_16158);
nand U17950 (N_17950,N_16743,N_16659);
and U17951 (N_17951,N_16708,N_16536);
xnor U17952 (N_17952,N_16444,N_15933);
nand U17953 (N_17953,N_15916,N_16405);
nor U17954 (N_17954,N_16746,N_16535);
xnor U17955 (N_17955,N_15697,N_16593);
nand U17956 (N_17956,N_16764,N_15916);
xnor U17957 (N_17957,N_16588,N_16230);
or U17958 (N_17958,N_15667,N_15901);
xnor U17959 (N_17959,N_15621,N_16283);
nor U17960 (N_17960,N_16781,N_16097);
nand U17961 (N_17961,N_16738,N_16017);
xnor U17962 (N_17962,N_16136,N_16468);
and U17963 (N_17963,N_15648,N_16553);
or U17964 (N_17964,N_16038,N_15734);
xnor U17965 (N_17965,N_16175,N_16257);
and U17966 (N_17966,N_15858,N_16310);
xnor U17967 (N_17967,N_15698,N_15683);
and U17968 (N_17968,N_15734,N_16494);
nor U17969 (N_17969,N_15837,N_15777);
nor U17970 (N_17970,N_16235,N_15757);
or U17971 (N_17971,N_16334,N_16649);
nor U17972 (N_17972,N_16002,N_16260);
xnor U17973 (N_17973,N_16531,N_16341);
nand U17974 (N_17974,N_16172,N_16463);
nor U17975 (N_17975,N_16703,N_16313);
or U17976 (N_17976,N_16188,N_15959);
or U17977 (N_17977,N_16571,N_16373);
xor U17978 (N_17978,N_16718,N_16341);
nor U17979 (N_17979,N_15694,N_15790);
and U17980 (N_17980,N_16721,N_16103);
or U17981 (N_17981,N_15688,N_15832);
nor U17982 (N_17982,N_15910,N_15846);
and U17983 (N_17983,N_16698,N_15613);
nor U17984 (N_17984,N_15655,N_15833);
xnor U17985 (N_17985,N_16561,N_16636);
or U17986 (N_17986,N_16656,N_16397);
xor U17987 (N_17987,N_15802,N_16287);
nor U17988 (N_17988,N_15830,N_16286);
xnor U17989 (N_17989,N_16159,N_16481);
nor U17990 (N_17990,N_16758,N_15853);
or U17991 (N_17991,N_15932,N_16220);
nand U17992 (N_17992,N_16675,N_16394);
nor U17993 (N_17993,N_15983,N_16569);
or U17994 (N_17994,N_16698,N_15787);
nand U17995 (N_17995,N_15946,N_16139);
and U17996 (N_17996,N_16608,N_15624);
or U17997 (N_17997,N_16234,N_16273);
or U17998 (N_17998,N_16208,N_16662);
xnor U17999 (N_17999,N_16172,N_15676);
or U18000 (N_18000,N_17535,N_17827);
nor U18001 (N_18001,N_17625,N_17167);
and U18002 (N_18002,N_17998,N_17201);
nand U18003 (N_18003,N_17174,N_17377);
or U18004 (N_18004,N_17960,N_17101);
nor U18005 (N_18005,N_17527,N_17733);
nand U18006 (N_18006,N_17037,N_17066);
nand U18007 (N_18007,N_17104,N_17283);
nand U18008 (N_18008,N_17515,N_17562);
xnor U18009 (N_18009,N_16803,N_17962);
xnor U18010 (N_18010,N_17788,N_16932);
nor U18011 (N_18011,N_17442,N_17819);
nor U18012 (N_18012,N_17516,N_17248);
xor U18013 (N_18013,N_17540,N_17006);
xnor U18014 (N_18014,N_16863,N_17492);
nor U18015 (N_18015,N_17900,N_16879);
and U18016 (N_18016,N_17461,N_17479);
nand U18017 (N_18017,N_17996,N_16826);
nor U18018 (N_18018,N_17302,N_17400);
xnor U18019 (N_18019,N_17877,N_16994);
nand U18020 (N_18020,N_17022,N_17452);
nor U18021 (N_18021,N_17495,N_17500);
or U18022 (N_18022,N_17117,N_17431);
or U18023 (N_18023,N_16978,N_17241);
or U18024 (N_18024,N_17284,N_17858);
nand U18025 (N_18025,N_17281,N_16969);
or U18026 (N_18026,N_17624,N_16975);
nand U18027 (N_18027,N_17252,N_17586);
and U18028 (N_18028,N_17993,N_16875);
and U18029 (N_18029,N_17246,N_17350);
nor U18030 (N_18030,N_17895,N_17790);
and U18031 (N_18031,N_17646,N_17756);
or U18032 (N_18032,N_17694,N_16937);
or U18033 (N_18033,N_17047,N_17940);
nor U18034 (N_18034,N_16801,N_17726);
nand U18035 (N_18035,N_17340,N_17390);
nor U18036 (N_18036,N_17845,N_17432);
xor U18037 (N_18037,N_16970,N_17210);
and U18038 (N_18038,N_17202,N_17472);
xnor U18039 (N_18039,N_17667,N_17575);
xor U18040 (N_18040,N_17100,N_17948);
or U18041 (N_18041,N_17093,N_16914);
xnor U18042 (N_18042,N_17884,N_17129);
and U18043 (N_18043,N_17588,N_17517);
nand U18044 (N_18044,N_17089,N_17091);
or U18045 (N_18045,N_17567,N_17449);
nor U18046 (N_18046,N_16841,N_17125);
nor U18047 (N_18047,N_17342,N_17383);
or U18048 (N_18048,N_16956,N_17822);
and U18049 (N_18049,N_16981,N_17863);
nor U18050 (N_18050,N_17685,N_17676);
nor U18051 (N_18051,N_17274,N_17956);
or U18052 (N_18052,N_17551,N_17207);
or U18053 (N_18053,N_17208,N_16849);
or U18054 (N_18054,N_17912,N_17634);
nand U18055 (N_18055,N_17490,N_17553);
and U18056 (N_18056,N_17847,N_17010);
nor U18057 (N_18057,N_16816,N_17769);
or U18058 (N_18058,N_17850,N_16878);
nor U18059 (N_18059,N_17236,N_17357);
and U18060 (N_18060,N_17149,N_17152);
or U18061 (N_18061,N_17581,N_16854);
and U18062 (N_18062,N_17361,N_17780);
or U18063 (N_18063,N_17489,N_17640);
nor U18064 (N_18064,N_17666,N_17007);
nand U18065 (N_18065,N_17249,N_17140);
nand U18066 (N_18066,N_17478,N_16870);
and U18067 (N_18067,N_17043,N_17166);
nor U18068 (N_18068,N_17306,N_17381);
or U18069 (N_18069,N_16943,N_17525);
nand U18070 (N_18070,N_17224,N_17052);
xor U18071 (N_18071,N_17983,N_17460);
nor U18072 (N_18072,N_17691,N_16961);
xnor U18073 (N_18073,N_17905,N_17650);
nand U18074 (N_18074,N_17784,N_17565);
or U18075 (N_18075,N_17740,N_17990);
nor U18076 (N_18076,N_17183,N_17739);
nor U18077 (N_18077,N_17402,N_16842);
nand U18078 (N_18078,N_17641,N_16967);
and U18079 (N_18079,N_17407,N_17215);
nand U18080 (N_18080,N_17404,N_17995);
xnor U18081 (N_18081,N_17734,N_17752);
and U18082 (N_18082,N_17419,N_17338);
nor U18083 (N_18083,N_17312,N_17760);
nand U18084 (N_18084,N_16954,N_17800);
nor U18085 (N_18085,N_17941,N_17865);
or U18086 (N_18086,N_17398,N_17664);
and U18087 (N_18087,N_17360,N_17929);
xor U18088 (N_18088,N_17409,N_16818);
nor U18089 (N_18089,N_17481,N_16944);
xnor U18090 (N_18090,N_17268,N_17805);
nand U18091 (N_18091,N_17602,N_17512);
xnor U18092 (N_18092,N_17391,N_17572);
or U18093 (N_18093,N_17121,N_16952);
or U18094 (N_18094,N_17566,N_17514);
nor U18095 (N_18095,N_17480,N_17485);
xnor U18096 (N_18096,N_17318,N_17766);
nand U18097 (N_18097,N_17065,N_16919);
xnor U18098 (N_18098,N_17373,N_16860);
or U18099 (N_18099,N_16844,N_17233);
or U18100 (N_18100,N_17534,N_17315);
or U18101 (N_18101,N_16977,N_17628);
or U18102 (N_18102,N_17656,N_17808);
xnor U18103 (N_18103,N_17272,N_17005);
and U18104 (N_18104,N_16899,N_16908);
xnor U18105 (N_18105,N_17055,N_17552);
or U18106 (N_18106,N_17722,N_17580);
xor U18107 (N_18107,N_16985,N_17486);
nand U18108 (N_18108,N_17613,N_17465);
xnor U18109 (N_18109,N_16928,N_17751);
or U18110 (N_18110,N_17818,N_17687);
or U18111 (N_18111,N_17802,N_17019);
xnor U18112 (N_18112,N_17369,N_17439);
xor U18113 (N_18113,N_17068,N_17292);
nor U18114 (N_18114,N_17874,N_17059);
or U18115 (N_18115,N_17343,N_17976);
nor U18116 (N_18116,N_17475,N_16855);
and U18117 (N_18117,N_17684,N_17522);
nand U18118 (N_18118,N_17111,N_17699);
or U18119 (N_18119,N_17882,N_17978);
xor U18120 (N_18120,N_16804,N_16809);
or U18121 (N_18121,N_17298,N_16976);
nand U18122 (N_18122,N_17584,N_17794);
xnor U18123 (N_18123,N_16993,N_17749);
xor U18124 (N_18124,N_17179,N_17075);
or U18125 (N_18125,N_16845,N_17310);
nor U18126 (N_18126,N_17484,N_17659);
xnor U18127 (N_18127,N_16979,N_17401);
and U18128 (N_18128,N_17108,N_17672);
xnor U18129 (N_18129,N_17754,N_17028);
xnor U18130 (N_18130,N_17970,N_17119);
or U18131 (N_18131,N_17366,N_17238);
nand U18132 (N_18132,N_17464,N_17928);
nor U18133 (N_18133,N_17275,N_17290);
nor U18134 (N_18134,N_17714,N_17943);
nand U18135 (N_18135,N_17798,N_17118);
nor U18136 (N_18136,N_17169,N_17771);
or U18137 (N_18137,N_17331,N_17741);
or U18138 (N_18138,N_17508,N_17840);
nand U18139 (N_18139,N_16988,N_17200);
xor U18140 (N_18140,N_17192,N_17384);
and U18141 (N_18141,N_17772,N_17999);
xnor U18142 (N_18142,N_17603,N_17707);
nand U18143 (N_18143,N_17397,N_17762);
xor U18144 (N_18144,N_17239,N_17335);
xnor U18145 (N_18145,N_17622,N_16945);
xor U18146 (N_18146,N_17765,N_16831);
xnor U18147 (N_18147,N_17244,N_17738);
or U18148 (N_18148,N_17795,N_16972);
xor U18149 (N_18149,N_17326,N_16906);
xor U18150 (N_18150,N_17499,N_17546);
or U18151 (N_18151,N_16865,N_17496);
xor U18152 (N_18152,N_17045,N_17520);
nand U18153 (N_18153,N_16847,N_17637);
nor U18154 (N_18154,N_17148,N_17387);
nor U18155 (N_18155,N_16987,N_17447);
or U18156 (N_18156,N_17730,N_17194);
nor U18157 (N_18157,N_17614,N_17151);
nand U18158 (N_18158,N_17632,N_17177);
nand U18159 (N_18159,N_16901,N_16857);
xor U18160 (N_18160,N_17959,N_17336);
nor U18161 (N_18161,N_17189,N_17955);
nor U18162 (N_18162,N_16931,N_17187);
nor U18163 (N_18163,N_17846,N_16839);
nand U18164 (N_18164,N_17203,N_17245);
and U18165 (N_18165,N_16866,N_16828);
xnor U18166 (N_18166,N_16838,N_16861);
and U18167 (N_18167,N_17792,N_17706);
or U18168 (N_18168,N_16827,N_16984);
nand U18169 (N_18169,N_17106,N_17297);
nor U18170 (N_18170,N_17643,N_17470);
and U18171 (N_18171,N_16902,N_17420);
xor U18172 (N_18172,N_16949,N_17090);
xor U18173 (N_18173,N_16966,N_16800);
nand U18174 (N_18174,N_17303,N_17930);
xnor U18175 (N_18175,N_17251,N_17997);
nor U18176 (N_18176,N_17523,N_17971);
nor U18177 (N_18177,N_17354,N_17809);
nor U18178 (N_18178,N_17209,N_17337);
xnor U18179 (N_18179,N_17592,N_17237);
or U18180 (N_18180,N_17261,N_17791);
and U18181 (N_18181,N_17597,N_17693);
nor U18182 (N_18182,N_17899,N_17559);
and U18183 (N_18183,N_16856,N_17473);
xor U18184 (N_18184,N_17957,N_17758);
and U18185 (N_18185,N_17204,N_17226);
and U18186 (N_18186,N_16836,N_17102);
xor U18187 (N_18187,N_17072,N_17185);
xor U18188 (N_18188,N_17058,N_17061);
or U18189 (N_18189,N_17103,N_17647);
or U18190 (N_18190,N_16884,N_17982);
xor U18191 (N_18191,N_17213,N_17083);
xnor U18192 (N_18192,N_17084,N_16903);
or U18193 (N_18193,N_17018,N_17026);
and U18194 (N_18194,N_17304,N_17405);
xor U18195 (N_18195,N_16889,N_17669);
or U18196 (N_18196,N_17184,N_17160);
nand U18197 (N_18197,N_17839,N_17864);
and U18198 (N_18198,N_16922,N_17892);
or U18199 (N_18199,N_16867,N_17379);
or U18200 (N_18200,N_16892,N_16980);
xnor U18201 (N_18201,N_17105,N_17688);
and U18202 (N_18202,N_17502,N_17265);
nor U18203 (N_18203,N_16874,N_17132);
xor U18204 (N_18204,N_17014,N_17073);
nor U18205 (N_18205,N_16999,N_17560);
xnor U18206 (N_18206,N_17901,N_17513);
or U18207 (N_18207,N_17175,N_17785);
or U18208 (N_18208,N_17074,N_17469);
nor U18209 (N_18209,N_17606,N_17848);
and U18210 (N_18210,N_17768,N_17168);
and U18211 (N_18211,N_17347,N_17674);
nor U18212 (N_18212,N_17456,N_17307);
nor U18213 (N_18213,N_17728,N_16876);
and U18214 (N_18214,N_17595,N_17974);
nor U18215 (N_18215,N_17044,N_16971);
and U18216 (N_18216,N_17723,N_17568);
nand U18217 (N_18217,N_17372,N_17986);
nand U18218 (N_18218,N_17935,N_17933);
and U18219 (N_18219,N_17334,N_17878);
nand U18220 (N_18220,N_17747,N_16881);
and U18221 (N_18221,N_17333,N_17182);
xor U18222 (N_18222,N_17138,N_16883);
or U18223 (N_18223,N_17443,N_17824);
or U18224 (N_18224,N_17040,N_16934);
nand U18225 (N_18225,N_17761,N_17231);
nand U18226 (N_18226,N_17109,N_17977);
or U18227 (N_18227,N_17851,N_17288);
or U18228 (N_18228,N_17036,N_17786);
or U18229 (N_18229,N_17041,N_17199);
xor U18230 (N_18230,N_17198,N_17910);
nor U18231 (N_18231,N_16930,N_17703);
nand U18232 (N_18232,N_16929,N_17164);
nand U18233 (N_18233,N_17378,N_17926);
xnor U18234 (N_18234,N_17423,N_16834);
or U18235 (N_18235,N_17911,N_17570);
xor U18236 (N_18236,N_17399,N_17356);
xnor U18237 (N_18237,N_17524,N_17627);
and U18238 (N_18238,N_17590,N_17596);
xnor U18239 (N_18239,N_17804,N_17287);
and U18240 (N_18240,N_17857,N_16888);
xor U18241 (N_18241,N_17985,N_17713);
xor U18242 (N_18242,N_17973,N_17776);
or U18243 (N_18243,N_16926,N_17020);
nor U18244 (N_18244,N_17406,N_16959);
and U18245 (N_18245,N_17085,N_17963);
nand U18246 (N_18246,N_17266,N_17147);
nor U18247 (N_18247,N_17435,N_16963);
xor U18248 (N_18248,N_16852,N_17725);
or U18249 (N_18249,N_17532,N_17433);
xor U18250 (N_18250,N_17374,N_17743);
xor U18251 (N_18251,N_17434,N_17662);
and U18252 (N_18252,N_17813,N_16858);
nor U18253 (N_18253,N_17587,N_17130);
or U18254 (N_18254,N_17427,N_17777);
or U18255 (N_18255,N_17339,N_17582);
nor U18256 (N_18256,N_17621,N_16933);
and U18257 (N_18257,N_17411,N_16864);
and U18258 (N_18258,N_16958,N_16895);
nand U18259 (N_18259,N_17981,N_17188);
nor U18260 (N_18260,N_17299,N_17161);
xor U18261 (N_18261,N_17697,N_16885);
nor U18262 (N_18262,N_17968,N_17050);
or U18263 (N_18263,N_17501,N_17852);
nand U18264 (N_18264,N_17345,N_16824);
nor U18265 (N_18265,N_17530,N_17269);
nand U18266 (N_18266,N_17285,N_17806);
xnor U18267 (N_18267,N_17143,N_17436);
xnor U18268 (N_18268,N_17114,N_17259);
nor U18269 (N_18269,N_17810,N_17867);
and U18270 (N_18270,N_16904,N_17894);
or U18271 (N_18271,N_17098,N_17416);
and U18272 (N_18272,N_16825,N_16806);
nor U18273 (N_18273,N_17086,N_17389);
xor U18274 (N_18274,N_17729,N_17746);
xnor U18275 (N_18275,N_17422,N_17654);
xnor U18276 (N_18276,N_16846,N_17604);
xor U18277 (N_18277,N_17529,N_17919);
xnor U18278 (N_18278,N_17126,N_17712);
nand U18279 (N_18279,N_17016,N_17942);
xor U18280 (N_18280,N_17979,N_17459);
and U18281 (N_18281,N_17498,N_17414);
or U18282 (N_18282,N_17171,N_17257);
or U18283 (N_18283,N_17577,N_16894);
xnor U18284 (N_18284,N_17113,N_17382);
and U18285 (N_18285,N_16869,N_17564);
nand U18286 (N_18286,N_17951,N_16820);
nor U18287 (N_18287,N_17885,N_17444);
and U18288 (N_18288,N_16940,N_17362);
xor U18289 (N_18289,N_16974,N_17950);
or U18290 (N_18290,N_17451,N_17814);
nor U18291 (N_18291,N_17250,N_17327);
nand U18292 (N_18292,N_17834,N_17286);
and U18293 (N_18293,N_17695,N_16942);
xnor U18294 (N_18294,N_17793,N_16813);
nor U18295 (N_18295,N_17533,N_17071);
or U18296 (N_18296,N_17150,N_17932);
nand U18297 (N_18297,N_17871,N_17629);
or U18298 (N_18298,N_17651,N_17528);
or U18299 (N_18299,N_17396,N_17773);
xor U18300 (N_18300,N_17032,N_17253);
and U18301 (N_18301,N_17745,N_17753);
nand U18302 (N_18302,N_17386,N_17862);
nor U18303 (N_18303,N_17004,N_17914);
nor U18304 (N_18304,N_17737,N_17679);
nand U18305 (N_18305,N_17711,N_17649);
nor U18306 (N_18306,N_17305,N_17294);
nand U18307 (N_18307,N_17821,N_17843);
xnor U18308 (N_18308,N_17178,N_17906);
or U18309 (N_18309,N_17365,N_17096);
nor U18310 (N_18310,N_17293,N_16909);
or U18311 (N_18311,N_17571,N_16819);
xnor U18312 (N_18312,N_17067,N_17173);
and U18313 (N_18313,N_17410,N_17046);
or U18314 (N_18314,N_17750,N_17057);
nor U18315 (N_18315,N_17056,N_17158);
nand U18316 (N_18316,N_17218,N_16814);
nor U18317 (N_18317,N_17353,N_17049);
and U18318 (N_18318,N_17537,N_16890);
and U18319 (N_18319,N_17035,N_17593);
and U18320 (N_18320,N_17142,N_16953);
or U18321 (N_18321,N_17759,N_17254);
nand U18322 (N_18322,N_17988,N_16882);
nor U18323 (N_18323,N_16998,N_17619);
nor U18324 (N_18324,N_17673,N_17958);
nor U18325 (N_18325,N_17736,N_17300);
or U18326 (N_18326,N_17547,N_17886);
nand U18327 (N_18327,N_16925,N_17011);
and U18328 (N_18328,N_17415,N_17817);
xnor U18329 (N_18329,N_16862,N_17205);
xnor U18330 (N_18330,N_17193,N_17506);
nor U18331 (N_18331,N_17618,N_17364);
xor U18332 (N_18332,N_16873,N_17324);
and U18333 (N_18333,N_17159,N_17869);
nand U18334 (N_18334,N_17346,N_16950);
xnor U18335 (N_18335,N_17242,N_16913);
or U18336 (N_18336,N_17328,N_16851);
xor U18337 (N_18337,N_17081,N_17270);
and U18338 (N_18338,N_17023,N_17429);
nand U18339 (N_18339,N_17042,N_17027);
nand U18340 (N_18340,N_17038,N_17991);
nand U18341 (N_18341,N_17891,N_17836);
and U18342 (N_18342,N_17927,N_17724);
nor U18343 (N_18343,N_17088,N_17898);
and U18344 (N_18344,N_17428,N_17062);
or U18345 (N_18345,N_17594,N_17934);
and U18346 (N_18346,N_17000,N_17380);
and U18347 (N_18347,N_17320,N_17609);
or U18348 (N_18348,N_17709,N_17137);
nand U18349 (N_18349,N_17191,N_17421);
nand U18350 (N_18350,N_17576,N_17296);
nand U18351 (N_18351,N_16939,N_17658);
or U18352 (N_18352,N_17015,N_17466);
xnor U18353 (N_18353,N_16920,N_17890);
or U18354 (N_18354,N_17639,N_17221);
and U18355 (N_18355,N_17116,N_17838);
or U18356 (N_18356,N_17219,N_17550);
nor U18357 (N_18357,N_17949,N_17363);
and U18358 (N_18358,N_16989,N_17260);
and U18359 (N_18359,N_16960,N_17543);
nor U18360 (N_18360,N_17868,N_17229);
nor U18361 (N_18361,N_17823,N_16853);
nand U18362 (N_18362,N_17860,N_17225);
nand U18363 (N_18363,N_17467,N_17033);
or U18364 (N_18364,N_17235,N_16887);
xor U18365 (N_18365,N_17494,N_17313);
nand U18366 (N_18366,N_17854,N_16923);
nand U18367 (N_18367,N_17921,N_17842);
xor U18368 (N_18368,N_16997,N_17180);
xor U18369 (N_18369,N_17938,N_17644);
nand U18370 (N_18370,N_17655,N_17917);
nor U18371 (N_18371,N_17853,N_16837);
or U18372 (N_18372,N_17170,N_17816);
nor U18373 (N_18373,N_17471,N_17789);
xor U18374 (N_18374,N_17003,N_17557);
nor U18375 (N_18375,N_16995,N_16891);
nor U18376 (N_18376,N_17220,N_17176);
and U18377 (N_18377,N_17732,N_17393);
nand U18378 (N_18378,N_17698,N_17457);
xnor U18379 (N_18379,N_17903,N_17539);
nor U18380 (N_18380,N_17031,N_17279);
nor U18381 (N_18381,N_17488,N_17563);
and U18382 (N_18382,N_17849,N_17329);
nor U18383 (N_18383,N_17855,N_17830);
or U18384 (N_18384,N_17441,N_17511);
nor U18385 (N_18385,N_17321,N_17141);
or U18386 (N_18386,N_17600,N_17653);
xnor U18387 (N_18387,N_17700,N_17538);
and U18388 (N_18388,N_17696,N_17888);
xor U18389 (N_18389,N_17352,N_16936);
xnor U18390 (N_18390,N_17526,N_17770);
nor U18391 (N_18391,N_16898,N_17051);
nand U18392 (N_18392,N_17787,N_17273);
nand U18393 (N_18393,N_17240,N_17394);
nand U18394 (N_18394,N_17944,N_17156);
or U18395 (N_18395,N_17607,N_17774);
or U18396 (N_18396,N_17797,N_17463);
and U18397 (N_18397,N_17799,N_17675);
xor U18398 (N_18398,N_17972,N_17230);
or U18399 (N_18399,N_16877,N_16948);
xnor U18400 (N_18400,N_17453,N_17545);
nor U18401 (N_18401,N_17418,N_17837);
xor U18402 (N_18402,N_17718,N_17682);
and U18403 (N_18403,N_17701,N_17316);
nor U18404 (N_18404,N_17332,N_17491);
or U18405 (N_18405,N_17154,N_17223);
or U18406 (N_18406,N_17680,N_16808);
nor U18407 (N_18407,N_17017,N_17112);
nand U18408 (N_18408,N_17692,N_16812);
and U18409 (N_18409,N_17965,N_16821);
nand U18410 (N_18410,N_16921,N_17438);
xor U18411 (N_18411,N_17217,N_17779);
nor U18412 (N_18412,N_17355,N_17476);
nand U18413 (N_18413,N_17907,N_16986);
nor U18414 (N_18414,N_17660,N_16835);
nand U18415 (N_18415,N_16924,N_17638);
nand U18416 (N_18416,N_17579,N_16905);
and U18417 (N_18417,N_17755,N_17358);
or U18418 (N_18418,N_17206,N_16871);
nand U18419 (N_18419,N_16927,N_17678);
nand U18420 (N_18420,N_17630,N_17987);
nor U18421 (N_18421,N_17216,N_17426);
nand U18422 (N_18422,N_17964,N_16805);
xor U18423 (N_18423,N_17897,N_17831);
and U18424 (N_18424,N_17348,N_17946);
xor U18425 (N_18425,N_17054,N_17136);
nor U18426 (N_18426,N_17908,N_17531);
nand U18427 (N_18427,N_17626,N_17896);
or U18428 (N_18428,N_17642,N_17359);
xor U18429 (N_18429,N_17146,N_17092);
and U18430 (N_18430,N_17705,N_17070);
and U18431 (N_18431,N_17195,N_17131);
or U18432 (N_18432,N_17992,N_17856);
and U18433 (N_18433,N_17462,N_17487);
or U18434 (N_18434,N_17681,N_17727);
xor U18435 (N_18435,N_17953,N_17504);
or U18436 (N_18436,N_17021,N_17835);
and U18437 (N_18437,N_17569,N_17145);
and U18438 (N_18438,N_16859,N_17255);
or U18439 (N_18439,N_17861,N_17893);
or U18440 (N_18440,N_17127,N_17889);
nor U18441 (N_18441,N_17120,N_16872);
nor U18442 (N_18442,N_17322,N_17617);
or U18443 (N_18443,N_17351,N_17735);
nand U18444 (N_18444,N_17317,N_17271);
and U18445 (N_18445,N_17228,N_17196);
xor U18446 (N_18446,N_17716,N_17128);
xnor U18447 (N_18447,N_17832,N_17913);
xor U18448 (N_18448,N_17731,N_17425);
and U18449 (N_18449,N_17099,N_17803);
nor U18450 (N_18450,N_17657,N_17757);
xnor U18451 (N_18451,N_16823,N_17599);
nand U18452 (N_18452,N_17967,N_17227);
nor U18453 (N_18453,N_17605,N_17468);
nand U18454 (N_18454,N_17833,N_17277);
nand U18455 (N_18455,N_17591,N_17264);
and U18456 (N_18456,N_17954,N_17197);
or U18457 (N_18457,N_17616,N_17243);
nor U18458 (N_18458,N_17034,N_17918);
nor U18459 (N_18459,N_17370,N_17133);
nand U18460 (N_18460,N_17087,N_17214);
and U18461 (N_18461,N_17686,N_17620);
and U18462 (N_18462,N_17039,N_17704);
or U18463 (N_18463,N_16915,N_17165);
nand U18464 (N_18464,N_17585,N_17875);
or U18465 (N_18465,N_17153,N_16810);
xor U18466 (N_18466,N_17162,N_17721);
nor U18467 (N_18467,N_17601,N_17232);
or U18468 (N_18468,N_17053,N_16996);
nor U18469 (N_18469,N_17069,N_17190);
or U18470 (N_18470,N_17222,N_16983);
nor U18471 (N_18471,N_16982,N_17872);
xnor U18472 (N_18472,N_16830,N_17916);
and U18473 (N_18473,N_17446,N_17135);
nand U18474 (N_18474,N_17902,N_17966);
nand U18475 (N_18475,N_17767,N_17163);
and U18476 (N_18476,N_17060,N_17445);
nand U18477 (N_18477,N_17608,N_17880);
xnor U18478 (N_18478,N_17134,N_17671);
and U18479 (N_18479,N_17385,N_17936);
nor U18480 (N_18480,N_16955,N_17289);
nand U18481 (N_18481,N_16910,N_17764);
or U18482 (N_18482,N_17536,N_17258);
xor U18483 (N_18483,N_17668,N_17826);
xnor U18484 (N_18484,N_17980,N_17841);
xor U18485 (N_18485,N_16918,N_17717);
nor U18486 (N_18486,N_16968,N_17424);
or U18487 (N_18487,N_17984,N_17989);
and U18488 (N_18488,N_17598,N_17388);
nand U18489 (N_18489,N_17825,N_17095);
nand U18490 (N_18490,N_17969,N_17078);
nor U18491 (N_18491,N_16900,N_17574);
and U18492 (N_18492,N_16951,N_17781);
xor U18493 (N_18493,N_16907,N_17403);
xor U18494 (N_18494,N_17859,N_17952);
or U18495 (N_18495,N_16850,N_16811);
nor U18496 (N_18496,N_17811,N_17482);
and U18497 (N_18497,N_17308,N_17742);
nor U18498 (N_18498,N_16822,N_17812);
and U18499 (N_18499,N_17048,N_17030);
xor U18500 (N_18500,N_17578,N_17412);
and U18501 (N_18501,N_17323,N_17110);
nor U18502 (N_18502,N_17807,N_17309);
nor U18503 (N_18503,N_17139,N_17262);
and U18504 (N_18504,N_17503,N_17931);
xor U18505 (N_18505,N_17458,N_17879);
and U18506 (N_18506,N_17631,N_17172);
and U18507 (N_18507,N_17395,N_17454);
nor U18508 (N_18508,N_17922,N_17212);
xor U18509 (N_18509,N_17677,N_16973);
xor U18510 (N_18510,N_16947,N_17583);
nor U18511 (N_18511,N_17325,N_17079);
xor U18512 (N_18512,N_17263,N_17077);
and U18513 (N_18513,N_16965,N_16832);
nand U18514 (N_18514,N_16991,N_17702);
or U18515 (N_18515,N_17611,N_17828);
or U18516 (N_18516,N_17663,N_17652);
and U18517 (N_18517,N_16964,N_17247);
xnor U18518 (N_18518,N_17815,N_17301);
nor U18519 (N_18519,N_17612,N_17124);
and U18520 (N_18520,N_17549,N_16886);
and U18521 (N_18521,N_17544,N_17648);
nand U18522 (N_18522,N_16912,N_16916);
xor U18523 (N_18523,N_17763,N_17276);
nor U18524 (N_18524,N_17645,N_17437);
nand U18525 (N_18525,N_17234,N_17368);
xnor U18526 (N_18526,N_17844,N_17211);
nand U18527 (N_18527,N_17720,N_17291);
nand U18528 (N_18528,N_17947,N_17558);
xnor U18529 (N_18529,N_17589,N_16829);
xor U18530 (N_18530,N_16896,N_16941);
nand U18531 (N_18531,N_17282,N_17904);
or U18532 (N_18532,N_17076,N_17330);
or U18533 (N_18533,N_16911,N_17923);
or U18534 (N_18534,N_17493,N_17521);
xnor U18535 (N_18535,N_17280,N_16938);
nor U18536 (N_18536,N_17939,N_16897);
xor U18537 (N_18537,N_17518,N_17556);
nor U18538 (N_18538,N_17873,N_16815);
nand U18539 (N_18539,N_17107,N_16946);
nor U18540 (N_18540,N_17554,N_17915);
xor U18541 (N_18541,N_17080,N_17349);
and U18542 (N_18542,N_17689,N_17367);
or U18543 (N_18543,N_17115,N_17341);
or U18544 (N_18544,N_17392,N_16880);
nor U18545 (N_18545,N_17267,N_17507);
nor U18546 (N_18546,N_17690,N_16990);
or U18547 (N_18547,N_17483,N_17881);
nor U18548 (N_18548,N_17024,N_17820);
or U18549 (N_18549,N_17455,N_17796);
or U18550 (N_18550,N_17295,N_17635);
and U18551 (N_18551,N_17314,N_17430);
nor U18552 (N_18552,N_17413,N_16917);
xnor U18553 (N_18553,N_16962,N_17477);
xor U18554 (N_18554,N_17920,N_17775);
or U18555 (N_18555,N_17748,N_17008);
nand U18556 (N_18556,N_17665,N_17887);
nor U18557 (N_18557,N_17541,N_17623);
or U18558 (N_18558,N_17801,N_17573);
and U18559 (N_18559,N_16833,N_17375);
and U18560 (N_18560,N_17876,N_17683);
nand U18561 (N_18561,N_17448,N_16935);
nand U18562 (N_18562,N_16802,N_17376);
and U18563 (N_18563,N_17924,N_16868);
nand U18564 (N_18564,N_17155,N_17440);
or U18565 (N_18565,N_16807,N_17013);
and U18566 (N_18566,N_17001,N_17122);
and U18567 (N_18567,N_17344,N_17025);
or U18568 (N_18568,N_16843,N_17719);
nand U18569 (N_18569,N_17909,N_17925);
and U18570 (N_18570,N_17715,N_17636);
or U18571 (N_18571,N_17181,N_17945);
nor U18572 (N_18572,N_17661,N_17542);
xor U18573 (N_18573,N_17783,N_17610);
and U18574 (N_18574,N_17311,N_17937);
nor U18575 (N_18575,N_17866,N_17256);
nor U18576 (N_18576,N_17097,N_16848);
or U18577 (N_18577,N_17474,N_17561);
nand U18578 (N_18578,N_17029,N_17510);
and U18579 (N_18579,N_17778,N_17064);
nor U18580 (N_18580,N_17123,N_17555);
and U18581 (N_18581,N_17009,N_17497);
and U18582 (N_18582,N_17186,N_17157);
xor U18583 (N_18583,N_16817,N_17883);
or U18584 (N_18584,N_17144,N_17870);
nor U18585 (N_18585,N_17505,N_17417);
and U18586 (N_18586,N_17519,N_17782);
and U18587 (N_18587,N_17708,N_17450);
and U18588 (N_18588,N_17278,N_17994);
nand U18589 (N_18589,N_17548,N_17371);
or U18590 (N_18590,N_17744,N_17094);
nand U18591 (N_18591,N_17082,N_17063);
or U18592 (N_18592,N_17961,N_16893);
or U18593 (N_18593,N_17509,N_17670);
nor U18594 (N_18594,N_17408,N_17615);
xnor U18595 (N_18595,N_17319,N_16957);
and U18596 (N_18596,N_17975,N_17633);
or U18597 (N_18597,N_17012,N_17710);
nor U18598 (N_18598,N_16992,N_17829);
nand U18599 (N_18599,N_16840,N_17002);
or U18600 (N_18600,N_17818,N_17441);
and U18601 (N_18601,N_16813,N_17811);
nor U18602 (N_18602,N_17123,N_17200);
nand U18603 (N_18603,N_17912,N_17593);
nand U18604 (N_18604,N_17480,N_16919);
nand U18605 (N_18605,N_17565,N_17403);
nor U18606 (N_18606,N_17446,N_17829);
xnor U18607 (N_18607,N_17554,N_16899);
nor U18608 (N_18608,N_17623,N_17781);
xor U18609 (N_18609,N_16966,N_16974);
nor U18610 (N_18610,N_16849,N_17624);
and U18611 (N_18611,N_17284,N_17921);
nand U18612 (N_18612,N_17375,N_16968);
nor U18613 (N_18613,N_17500,N_17109);
nor U18614 (N_18614,N_17805,N_17935);
and U18615 (N_18615,N_17682,N_17296);
nand U18616 (N_18616,N_17428,N_17787);
nand U18617 (N_18617,N_17873,N_16875);
or U18618 (N_18618,N_17391,N_17860);
and U18619 (N_18619,N_16954,N_16987);
nand U18620 (N_18620,N_17597,N_17123);
or U18621 (N_18621,N_17160,N_17939);
xnor U18622 (N_18622,N_17109,N_17973);
or U18623 (N_18623,N_16846,N_17739);
and U18624 (N_18624,N_17848,N_17923);
xnor U18625 (N_18625,N_17617,N_17078);
nand U18626 (N_18626,N_17094,N_17506);
nor U18627 (N_18627,N_17039,N_17371);
nand U18628 (N_18628,N_16968,N_17133);
nor U18629 (N_18629,N_17160,N_17206);
or U18630 (N_18630,N_17020,N_17155);
and U18631 (N_18631,N_17184,N_17622);
or U18632 (N_18632,N_17861,N_17230);
nor U18633 (N_18633,N_16938,N_17740);
nand U18634 (N_18634,N_17543,N_17504);
and U18635 (N_18635,N_17233,N_16960);
or U18636 (N_18636,N_16880,N_17576);
nor U18637 (N_18637,N_17632,N_17190);
nor U18638 (N_18638,N_17125,N_17668);
nand U18639 (N_18639,N_17334,N_17864);
nor U18640 (N_18640,N_17121,N_17230);
xnor U18641 (N_18641,N_17061,N_17856);
nand U18642 (N_18642,N_17563,N_17791);
or U18643 (N_18643,N_17446,N_17703);
and U18644 (N_18644,N_17549,N_17235);
or U18645 (N_18645,N_16846,N_17615);
nor U18646 (N_18646,N_17752,N_17738);
and U18647 (N_18647,N_17125,N_17233);
and U18648 (N_18648,N_17375,N_17478);
xnor U18649 (N_18649,N_17463,N_16869);
xor U18650 (N_18650,N_17297,N_17795);
xor U18651 (N_18651,N_17241,N_17881);
nand U18652 (N_18652,N_17165,N_17569);
and U18653 (N_18653,N_17298,N_17156);
and U18654 (N_18654,N_17468,N_17357);
or U18655 (N_18655,N_16965,N_16929);
or U18656 (N_18656,N_16817,N_17637);
nor U18657 (N_18657,N_17425,N_17438);
or U18658 (N_18658,N_17857,N_17253);
xor U18659 (N_18659,N_17256,N_16909);
or U18660 (N_18660,N_17168,N_17028);
nor U18661 (N_18661,N_16847,N_17754);
xor U18662 (N_18662,N_16932,N_16878);
nand U18663 (N_18663,N_17087,N_17508);
and U18664 (N_18664,N_17259,N_17771);
or U18665 (N_18665,N_17771,N_17516);
nand U18666 (N_18666,N_17728,N_16883);
or U18667 (N_18667,N_17538,N_17719);
xor U18668 (N_18668,N_17757,N_17867);
xor U18669 (N_18669,N_17295,N_16887);
and U18670 (N_18670,N_17939,N_17719);
nand U18671 (N_18671,N_17161,N_16851);
and U18672 (N_18672,N_17413,N_17752);
xnor U18673 (N_18673,N_17350,N_17635);
nand U18674 (N_18674,N_16944,N_17072);
xnor U18675 (N_18675,N_17307,N_17697);
nor U18676 (N_18676,N_16805,N_17974);
nor U18677 (N_18677,N_17747,N_17253);
xor U18678 (N_18678,N_17979,N_17429);
xor U18679 (N_18679,N_17858,N_16883);
nor U18680 (N_18680,N_17550,N_16959);
xor U18681 (N_18681,N_17992,N_16923);
xnor U18682 (N_18682,N_17948,N_16917);
nor U18683 (N_18683,N_17455,N_16986);
nor U18684 (N_18684,N_16930,N_17046);
xor U18685 (N_18685,N_17516,N_17154);
and U18686 (N_18686,N_17078,N_17411);
and U18687 (N_18687,N_17474,N_17458);
or U18688 (N_18688,N_17106,N_16922);
nor U18689 (N_18689,N_16820,N_17985);
nor U18690 (N_18690,N_17910,N_17370);
xnor U18691 (N_18691,N_17700,N_17225);
and U18692 (N_18692,N_17546,N_17989);
xor U18693 (N_18693,N_17071,N_16858);
or U18694 (N_18694,N_17257,N_17298);
xor U18695 (N_18695,N_17385,N_17371);
and U18696 (N_18696,N_17137,N_17864);
or U18697 (N_18697,N_17331,N_17593);
and U18698 (N_18698,N_17265,N_16869);
and U18699 (N_18699,N_16868,N_17477);
xnor U18700 (N_18700,N_17867,N_17554);
nor U18701 (N_18701,N_17214,N_17014);
xnor U18702 (N_18702,N_17670,N_17901);
nand U18703 (N_18703,N_17710,N_17150);
or U18704 (N_18704,N_17721,N_17843);
nor U18705 (N_18705,N_17696,N_17234);
and U18706 (N_18706,N_17349,N_17962);
xnor U18707 (N_18707,N_17122,N_17374);
nor U18708 (N_18708,N_17057,N_17789);
nor U18709 (N_18709,N_17536,N_17574);
xnor U18710 (N_18710,N_17896,N_16980);
nand U18711 (N_18711,N_17270,N_17656);
nand U18712 (N_18712,N_17857,N_17903);
or U18713 (N_18713,N_17603,N_17659);
nor U18714 (N_18714,N_17470,N_17837);
and U18715 (N_18715,N_16938,N_16811);
nor U18716 (N_18716,N_17067,N_17812);
or U18717 (N_18717,N_17676,N_17930);
xnor U18718 (N_18718,N_17262,N_17960);
xnor U18719 (N_18719,N_17935,N_17603);
nand U18720 (N_18720,N_17577,N_16930);
or U18721 (N_18721,N_17847,N_17921);
nor U18722 (N_18722,N_16964,N_17647);
nand U18723 (N_18723,N_17334,N_17503);
or U18724 (N_18724,N_16817,N_16922);
nor U18725 (N_18725,N_17196,N_17446);
or U18726 (N_18726,N_17488,N_17972);
or U18727 (N_18727,N_17326,N_17758);
xor U18728 (N_18728,N_17656,N_16875);
and U18729 (N_18729,N_17514,N_16862);
or U18730 (N_18730,N_17851,N_17036);
nand U18731 (N_18731,N_16960,N_17193);
or U18732 (N_18732,N_16909,N_17891);
nor U18733 (N_18733,N_17312,N_17295);
or U18734 (N_18734,N_17765,N_17059);
nand U18735 (N_18735,N_17790,N_17658);
and U18736 (N_18736,N_17279,N_17142);
xor U18737 (N_18737,N_17142,N_17403);
nand U18738 (N_18738,N_17253,N_17599);
xnor U18739 (N_18739,N_17879,N_16985);
or U18740 (N_18740,N_17195,N_17027);
or U18741 (N_18741,N_17016,N_16878);
nand U18742 (N_18742,N_17014,N_17622);
or U18743 (N_18743,N_17196,N_17922);
xnor U18744 (N_18744,N_17092,N_17920);
xor U18745 (N_18745,N_17313,N_16923);
nor U18746 (N_18746,N_17189,N_17256);
xor U18747 (N_18747,N_17504,N_17007);
xor U18748 (N_18748,N_17702,N_16956);
xor U18749 (N_18749,N_17236,N_17295);
xnor U18750 (N_18750,N_16938,N_17660);
xor U18751 (N_18751,N_17703,N_17885);
xnor U18752 (N_18752,N_16811,N_17622);
or U18753 (N_18753,N_17458,N_17283);
nor U18754 (N_18754,N_17678,N_17210);
and U18755 (N_18755,N_17479,N_17335);
or U18756 (N_18756,N_17793,N_17026);
xnor U18757 (N_18757,N_16923,N_17120);
or U18758 (N_18758,N_17146,N_17496);
nor U18759 (N_18759,N_17598,N_17507);
nor U18760 (N_18760,N_17005,N_17207);
and U18761 (N_18761,N_17867,N_16967);
nand U18762 (N_18762,N_17006,N_17170);
nand U18763 (N_18763,N_17616,N_17880);
nand U18764 (N_18764,N_17240,N_17271);
nand U18765 (N_18765,N_16911,N_17183);
nand U18766 (N_18766,N_17412,N_17367);
xnor U18767 (N_18767,N_17191,N_17658);
or U18768 (N_18768,N_17045,N_17295);
nor U18769 (N_18769,N_17609,N_16927);
and U18770 (N_18770,N_17383,N_16981);
nor U18771 (N_18771,N_17767,N_17647);
nand U18772 (N_18772,N_17879,N_17446);
xnor U18773 (N_18773,N_17716,N_16871);
nand U18774 (N_18774,N_17770,N_16833);
or U18775 (N_18775,N_17076,N_17526);
and U18776 (N_18776,N_16884,N_17437);
and U18777 (N_18777,N_17628,N_17198);
or U18778 (N_18778,N_17176,N_17039);
and U18779 (N_18779,N_17038,N_17639);
xnor U18780 (N_18780,N_17042,N_17690);
nor U18781 (N_18781,N_17648,N_17342);
xor U18782 (N_18782,N_16943,N_17633);
nand U18783 (N_18783,N_17795,N_16960);
xor U18784 (N_18784,N_17401,N_17997);
nand U18785 (N_18785,N_17281,N_17443);
nor U18786 (N_18786,N_17186,N_17172);
and U18787 (N_18787,N_17810,N_17423);
and U18788 (N_18788,N_17717,N_17393);
xnor U18789 (N_18789,N_17076,N_17434);
nand U18790 (N_18790,N_17526,N_17112);
and U18791 (N_18791,N_16903,N_17365);
nor U18792 (N_18792,N_17476,N_16816);
xnor U18793 (N_18793,N_17506,N_17119);
or U18794 (N_18794,N_17582,N_17405);
xor U18795 (N_18795,N_17292,N_17094);
nand U18796 (N_18796,N_16868,N_17908);
xnor U18797 (N_18797,N_17230,N_17965);
nand U18798 (N_18798,N_16999,N_16906);
or U18799 (N_18799,N_16803,N_17218);
and U18800 (N_18800,N_17569,N_17987);
nand U18801 (N_18801,N_17896,N_16858);
nand U18802 (N_18802,N_17739,N_17471);
xnor U18803 (N_18803,N_16953,N_17272);
nor U18804 (N_18804,N_16891,N_16848);
and U18805 (N_18805,N_17973,N_17132);
xor U18806 (N_18806,N_17567,N_17342);
or U18807 (N_18807,N_17103,N_16863);
nor U18808 (N_18808,N_17150,N_17613);
xnor U18809 (N_18809,N_17984,N_17682);
or U18810 (N_18810,N_17020,N_16825);
nor U18811 (N_18811,N_17537,N_17998);
or U18812 (N_18812,N_17143,N_17453);
nor U18813 (N_18813,N_17355,N_17969);
and U18814 (N_18814,N_17585,N_17577);
and U18815 (N_18815,N_17184,N_16968);
nor U18816 (N_18816,N_17807,N_17004);
and U18817 (N_18817,N_17855,N_17840);
nor U18818 (N_18818,N_17193,N_17851);
or U18819 (N_18819,N_17764,N_17659);
or U18820 (N_18820,N_17948,N_17983);
and U18821 (N_18821,N_17967,N_16871);
nand U18822 (N_18822,N_16943,N_17401);
or U18823 (N_18823,N_17286,N_17216);
and U18824 (N_18824,N_16805,N_17225);
xor U18825 (N_18825,N_16805,N_17057);
and U18826 (N_18826,N_17027,N_16918);
or U18827 (N_18827,N_17535,N_17244);
nand U18828 (N_18828,N_17670,N_17408);
xnor U18829 (N_18829,N_17089,N_17906);
nand U18830 (N_18830,N_16824,N_17695);
or U18831 (N_18831,N_17671,N_17041);
or U18832 (N_18832,N_17641,N_17919);
and U18833 (N_18833,N_17066,N_16920);
nand U18834 (N_18834,N_17189,N_17761);
and U18835 (N_18835,N_17783,N_17159);
xnor U18836 (N_18836,N_17043,N_17497);
nand U18837 (N_18837,N_16839,N_17177);
or U18838 (N_18838,N_16870,N_17904);
or U18839 (N_18839,N_17957,N_16922);
nor U18840 (N_18840,N_17094,N_17627);
or U18841 (N_18841,N_17485,N_17179);
or U18842 (N_18842,N_17315,N_17535);
xnor U18843 (N_18843,N_17448,N_17979);
nor U18844 (N_18844,N_17067,N_17904);
nor U18845 (N_18845,N_16867,N_17083);
xor U18846 (N_18846,N_17277,N_16861);
xnor U18847 (N_18847,N_17431,N_17596);
nand U18848 (N_18848,N_17298,N_17976);
or U18849 (N_18849,N_17518,N_17125);
xor U18850 (N_18850,N_17201,N_17767);
and U18851 (N_18851,N_17724,N_17169);
nor U18852 (N_18852,N_17313,N_17674);
nor U18853 (N_18853,N_17872,N_16850);
xnor U18854 (N_18854,N_17927,N_17315);
or U18855 (N_18855,N_17592,N_17971);
nand U18856 (N_18856,N_17000,N_17037);
and U18857 (N_18857,N_17550,N_17691);
or U18858 (N_18858,N_17820,N_17199);
nor U18859 (N_18859,N_16850,N_16859);
nand U18860 (N_18860,N_16804,N_17234);
xnor U18861 (N_18861,N_16956,N_16951);
or U18862 (N_18862,N_17577,N_17174);
or U18863 (N_18863,N_17631,N_17940);
xnor U18864 (N_18864,N_17339,N_17326);
nand U18865 (N_18865,N_16867,N_17483);
xor U18866 (N_18866,N_17935,N_16831);
xnor U18867 (N_18867,N_17143,N_17325);
or U18868 (N_18868,N_17079,N_17549);
and U18869 (N_18869,N_17689,N_17636);
or U18870 (N_18870,N_17885,N_17690);
nand U18871 (N_18871,N_17518,N_17969);
nor U18872 (N_18872,N_17679,N_17280);
nor U18873 (N_18873,N_16974,N_16992);
nand U18874 (N_18874,N_17058,N_17465);
nand U18875 (N_18875,N_16903,N_17388);
or U18876 (N_18876,N_17240,N_17350);
nor U18877 (N_18877,N_17306,N_17477);
or U18878 (N_18878,N_17230,N_17696);
nor U18879 (N_18879,N_17290,N_17302);
and U18880 (N_18880,N_17949,N_17369);
xnor U18881 (N_18881,N_17336,N_17226);
and U18882 (N_18882,N_16944,N_17841);
nor U18883 (N_18883,N_17710,N_17225);
and U18884 (N_18884,N_17132,N_17606);
or U18885 (N_18885,N_17161,N_17573);
xnor U18886 (N_18886,N_17557,N_16990);
nand U18887 (N_18887,N_17651,N_17319);
xor U18888 (N_18888,N_17029,N_17121);
nand U18889 (N_18889,N_17650,N_17187);
xor U18890 (N_18890,N_17012,N_17309);
nand U18891 (N_18891,N_17418,N_17389);
nor U18892 (N_18892,N_17627,N_16845);
xor U18893 (N_18893,N_17380,N_17725);
nand U18894 (N_18894,N_17791,N_16946);
and U18895 (N_18895,N_17321,N_17545);
nor U18896 (N_18896,N_17228,N_16886);
and U18897 (N_18897,N_17610,N_17859);
nand U18898 (N_18898,N_16868,N_17991);
and U18899 (N_18899,N_16944,N_17385);
nor U18900 (N_18900,N_16965,N_16902);
or U18901 (N_18901,N_17647,N_17298);
xor U18902 (N_18902,N_17600,N_17039);
nor U18903 (N_18903,N_17169,N_17461);
or U18904 (N_18904,N_17022,N_17212);
xor U18905 (N_18905,N_17236,N_17559);
nor U18906 (N_18906,N_17965,N_17589);
nand U18907 (N_18907,N_17742,N_17084);
xnor U18908 (N_18908,N_17878,N_16976);
nor U18909 (N_18909,N_17275,N_16835);
nand U18910 (N_18910,N_17416,N_17614);
xnor U18911 (N_18911,N_17512,N_17593);
and U18912 (N_18912,N_16864,N_17091);
nor U18913 (N_18913,N_17864,N_17299);
nand U18914 (N_18914,N_17518,N_17052);
xor U18915 (N_18915,N_17901,N_17984);
xor U18916 (N_18916,N_17023,N_17049);
nand U18917 (N_18917,N_17387,N_17768);
nand U18918 (N_18918,N_17404,N_17807);
nand U18919 (N_18919,N_17901,N_17621);
or U18920 (N_18920,N_17072,N_17194);
or U18921 (N_18921,N_17439,N_17506);
nor U18922 (N_18922,N_17178,N_16962);
nor U18923 (N_18923,N_17964,N_17514);
or U18924 (N_18924,N_17423,N_17766);
nand U18925 (N_18925,N_17885,N_17124);
or U18926 (N_18926,N_16988,N_16989);
and U18927 (N_18927,N_17534,N_17946);
nor U18928 (N_18928,N_16891,N_17745);
nand U18929 (N_18929,N_17144,N_17024);
xnor U18930 (N_18930,N_17433,N_17985);
nor U18931 (N_18931,N_17794,N_17546);
and U18932 (N_18932,N_17528,N_17090);
nand U18933 (N_18933,N_17752,N_17641);
nand U18934 (N_18934,N_17380,N_16801);
or U18935 (N_18935,N_17038,N_17961);
nor U18936 (N_18936,N_17089,N_17268);
or U18937 (N_18937,N_17396,N_17665);
nor U18938 (N_18938,N_17655,N_17185);
or U18939 (N_18939,N_17235,N_17952);
or U18940 (N_18940,N_17082,N_17112);
and U18941 (N_18941,N_17260,N_17848);
nand U18942 (N_18942,N_16883,N_17311);
nand U18943 (N_18943,N_17146,N_17205);
nand U18944 (N_18944,N_17512,N_17830);
xnor U18945 (N_18945,N_17921,N_17773);
nand U18946 (N_18946,N_17749,N_17729);
nor U18947 (N_18947,N_17133,N_17632);
nand U18948 (N_18948,N_17979,N_17832);
nor U18949 (N_18949,N_17271,N_17186);
or U18950 (N_18950,N_17205,N_17658);
and U18951 (N_18951,N_17296,N_17588);
nor U18952 (N_18952,N_17174,N_17401);
nor U18953 (N_18953,N_17672,N_17256);
nand U18954 (N_18954,N_16961,N_17860);
nor U18955 (N_18955,N_17481,N_17349);
nor U18956 (N_18956,N_16885,N_17580);
and U18957 (N_18957,N_16822,N_17150);
and U18958 (N_18958,N_17957,N_17290);
nor U18959 (N_18959,N_17819,N_17499);
xor U18960 (N_18960,N_17588,N_17167);
and U18961 (N_18961,N_17211,N_16908);
and U18962 (N_18962,N_17122,N_17985);
nand U18963 (N_18963,N_17068,N_16805);
and U18964 (N_18964,N_17338,N_17328);
nand U18965 (N_18965,N_17257,N_17684);
or U18966 (N_18966,N_17277,N_17438);
nor U18967 (N_18967,N_17811,N_17484);
nor U18968 (N_18968,N_17537,N_17562);
and U18969 (N_18969,N_16833,N_17136);
and U18970 (N_18970,N_17137,N_17913);
and U18971 (N_18971,N_17336,N_17503);
or U18972 (N_18972,N_17052,N_16972);
and U18973 (N_18973,N_17830,N_17587);
and U18974 (N_18974,N_17598,N_17917);
or U18975 (N_18975,N_17637,N_17657);
and U18976 (N_18976,N_17259,N_17086);
and U18977 (N_18977,N_16986,N_17650);
xnor U18978 (N_18978,N_17415,N_17160);
or U18979 (N_18979,N_16956,N_17490);
or U18980 (N_18980,N_16908,N_17228);
xor U18981 (N_18981,N_17490,N_17828);
xor U18982 (N_18982,N_16972,N_17632);
and U18983 (N_18983,N_17206,N_17779);
nand U18984 (N_18984,N_17245,N_17290);
and U18985 (N_18985,N_17826,N_17735);
nor U18986 (N_18986,N_17950,N_17159);
xor U18987 (N_18987,N_17208,N_17221);
nor U18988 (N_18988,N_17514,N_16963);
xor U18989 (N_18989,N_17868,N_17098);
or U18990 (N_18990,N_17723,N_17605);
nand U18991 (N_18991,N_17308,N_16837);
xor U18992 (N_18992,N_17528,N_16927);
nor U18993 (N_18993,N_17677,N_17683);
nor U18994 (N_18994,N_17624,N_17405);
or U18995 (N_18995,N_17272,N_17834);
or U18996 (N_18996,N_17001,N_17873);
nand U18997 (N_18997,N_17112,N_17558);
nand U18998 (N_18998,N_17803,N_17316);
nor U18999 (N_18999,N_17611,N_17279);
nand U19000 (N_19000,N_17731,N_17909);
xor U19001 (N_19001,N_16862,N_17656);
nor U19002 (N_19002,N_16849,N_17180);
or U19003 (N_19003,N_17563,N_17764);
and U19004 (N_19004,N_17126,N_16932);
and U19005 (N_19005,N_17574,N_17228);
or U19006 (N_19006,N_17007,N_17067);
and U19007 (N_19007,N_17919,N_17907);
nand U19008 (N_19008,N_17948,N_17858);
xor U19009 (N_19009,N_17209,N_17651);
xnor U19010 (N_19010,N_16943,N_17521);
and U19011 (N_19011,N_17489,N_16950);
and U19012 (N_19012,N_17479,N_17483);
nor U19013 (N_19013,N_17620,N_17899);
and U19014 (N_19014,N_16891,N_17181);
nand U19015 (N_19015,N_16882,N_17162);
or U19016 (N_19016,N_17124,N_17796);
and U19017 (N_19017,N_17752,N_17809);
and U19018 (N_19018,N_17686,N_17805);
or U19019 (N_19019,N_17985,N_17360);
xor U19020 (N_19020,N_17483,N_16919);
or U19021 (N_19021,N_17421,N_16975);
or U19022 (N_19022,N_17790,N_17488);
and U19023 (N_19023,N_17833,N_17906);
and U19024 (N_19024,N_17120,N_16809);
or U19025 (N_19025,N_17625,N_17084);
and U19026 (N_19026,N_17906,N_17995);
and U19027 (N_19027,N_17176,N_16817);
and U19028 (N_19028,N_17676,N_17439);
and U19029 (N_19029,N_17316,N_17105);
nor U19030 (N_19030,N_16840,N_17434);
nand U19031 (N_19031,N_17597,N_17538);
xor U19032 (N_19032,N_17793,N_17395);
or U19033 (N_19033,N_16948,N_17950);
nand U19034 (N_19034,N_17153,N_17754);
nor U19035 (N_19035,N_16996,N_17097);
nor U19036 (N_19036,N_16960,N_17212);
nand U19037 (N_19037,N_17157,N_17831);
or U19038 (N_19038,N_17817,N_17506);
xnor U19039 (N_19039,N_17393,N_17055);
or U19040 (N_19040,N_17518,N_17274);
nand U19041 (N_19041,N_17226,N_17679);
nor U19042 (N_19042,N_17575,N_17187);
and U19043 (N_19043,N_17789,N_16905);
nand U19044 (N_19044,N_17934,N_17653);
or U19045 (N_19045,N_16899,N_17298);
or U19046 (N_19046,N_17661,N_17654);
nand U19047 (N_19047,N_17951,N_17990);
or U19048 (N_19048,N_17232,N_17514);
and U19049 (N_19049,N_17292,N_17882);
xnor U19050 (N_19050,N_17910,N_17369);
and U19051 (N_19051,N_16845,N_17095);
or U19052 (N_19052,N_17472,N_17804);
nand U19053 (N_19053,N_17116,N_17154);
nor U19054 (N_19054,N_17418,N_17967);
nand U19055 (N_19055,N_17866,N_17126);
nand U19056 (N_19056,N_17457,N_17497);
xor U19057 (N_19057,N_17630,N_17788);
xnor U19058 (N_19058,N_17482,N_17071);
or U19059 (N_19059,N_17261,N_17942);
xnor U19060 (N_19060,N_17183,N_17089);
xnor U19061 (N_19061,N_17138,N_17872);
xor U19062 (N_19062,N_17647,N_17075);
xnor U19063 (N_19063,N_17087,N_16933);
nand U19064 (N_19064,N_17111,N_17002);
xnor U19065 (N_19065,N_17884,N_17998);
and U19066 (N_19066,N_17805,N_16888);
nand U19067 (N_19067,N_17058,N_17607);
xor U19068 (N_19068,N_17743,N_17580);
and U19069 (N_19069,N_17771,N_17970);
nor U19070 (N_19070,N_16854,N_17908);
or U19071 (N_19071,N_17053,N_17662);
nor U19072 (N_19072,N_17420,N_16927);
xor U19073 (N_19073,N_17121,N_17619);
or U19074 (N_19074,N_17675,N_17889);
nor U19075 (N_19075,N_17190,N_17334);
or U19076 (N_19076,N_16958,N_17219);
nand U19077 (N_19077,N_17462,N_17215);
nand U19078 (N_19078,N_17966,N_17325);
nand U19079 (N_19079,N_16983,N_17028);
nand U19080 (N_19080,N_17799,N_17036);
nand U19081 (N_19081,N_17209,N_17492);
nand U19082 (N_19082,N_17217,N_17762);
and U19083 (N_19083,N_17952,N_17531);
and U19084 (N_19084,N_17967,N_17904);
xor U19085 (N_19085,N_17399,N_17004);
nand U19086 (N_19086,N_17927,N_17302);
xor U19087 (N_19087,N_17834,N_17191);
xor U19088 (N_19088,N_17366,N_17683);
nand U19089 (N_19089,N_17896,N_17825);
xnor U19090 (N_19090,N_16829,N_16894);
nand U19091 (N_19091,N_17300,N_17919);
xnor U19092 (N_19092,N_17889,N_16945);
or U19093 (N_19093,N_17720,N_17692);
xor U19094 (N_19094,N_17499,N_16856);
xor U19095 (N_19095,N_17878,N_17927);
or U19096 (N_19096,N_17773,N_16944);
xnor U19097 (N_19097,N_17264,N_17015);
nand U19098 (N_19098,N_17500,N_17499);
or U19099 (N_19099,N_17118,N_17454);
and U19100 (N_19100,N_17873,N_16943);
nor U19101 (N_19101,N_17882,N_17599);
or U19102 (N_19102,N_17113,N_16878);
xor U19103 (N_19103,N_17251,N_17643);
xor U19104 (N_19104,N_17226,N_17109);
xnor U19105 (N_19105,N_16968,N_17213);
nor U19106 (N_19106,N_17930,N_17213);
nand U19107 (N_19107,N_17095,N_17094);
xnor U19108 (N_19108,N_17423,N_16832);
nand U19109 (N_19109,N_17146,N_17557);
or U19110 (N_19110,N_17607,N_17826);
nand U19111 (N_19111,N_16865,N_17607);
nor U19112 (N_19112,N_17821,N_16992);
xnor U19113 (N_19113,N_17967,N_17700);
nor U19114 (N_19114,N_17697,N_17459);
or U19115 (N_19115,N_17106,N_16928);
xnor U19116 (N_19116,N_17646,N_17202);
xor U19117 (N_19117,N_17163,N_16895);
xnor U19118 (N_19118,N_17849,N_17953);
nand U19119 (N_19119,N_17865,N_17284);
nor U19120 (N_19120,N_17146,N_17938);
or U19121 (N_19121,N_17716,N_17127);
nand U19122 (N_19122,N_17105,N_17063);
and U19123 (N_19123,N_17564,N_17201);
nor U19124 (N_19124,N_17427,N_17716);
or U19125 (N_19125,N_17459,N_17197);
or U19126 (N_19126,N_17006,N_17556);
nand U19127 (N_19127,N_17995,N_17684);
xnor U19128 (N_19128,N_17432,N_17442);
xor U19129 (N_19129,N_16932,N_17306);
nand U19130 (N_19130,N_16889,N_17257);
nand U19131 (N_19131,N_17905,N_16894);
nor U19132 (N_19132,N_17724,N_17554);
nand U19133 (N_19133,N_17375,N_17855);
and U19134 (N_19134,N_17226,N_17585);
xor U19135 (N_19135,N_17038,N_17337);
and U19136 (N_19136,N_17143,N_17800);
or U19137 (N_19137,N_17699,N_17210);
or U19138 (N_19138,N_17067,N_17295);
nand U19139 (N_19139,N_17434,N_17704);
or U19140 (N_19140,N_17765,N_17556);
nand U19141 (N_19141,N_16948,N_17753);
or U19142 (N_19142,N_16898,N_17045);
nand U19143 (N_19143,N_17493,N_17602);
and U19144 (N_19144,N_17240,N_16804);
nand U19145 (N_19145,N_17753,N_17836);
xnor U19146 (N_19146,N_17481,N_17625);
or U19147 (N_19147,N_17881,N_17820);
and U19148 (N_19148,N_17208,N_17876);
nand U19149 (N_19149,N_17080,N_17378);
xnor U19150 (N_19150,N_17634,N_16842);
xor U19151 (N_19151,N_17983,N_17875);
or U19152 (N_19152,N_17563,N_17915);
and U19153 (N_19153,N_17950,N_16988);
and U19154 (N_19154,N_17356,N_17297);
nand U19155 (N_19155,N_17371,N_17640);
nor U19156 (N_19156,N_17481,N_17999);
nand U19157 (N_19157,N_17982,N_17104);
nand U19158 (N_19158,N_17088,N_17208);
xnor U19159 (N_19159,N_17535,N_16918);
nand U19160 (N_19160,N_16853,N_17719);
and U19161 (N_19161,N_16882,N_17208);
nand U19162 (N_19162,N_16896,N_17034);
or U19163 (N_19163,N_17248,N_17356);
nand U19164 (N_19164,N_17380,N_17814);
nor U19165 (N_19165,N_17410,N_17484);
nor U19166 (N_19166,N_16835,N_17312);
nor U19167 (N_19167,N_17466,N_17853);
xor U19168 (N_19168,N_17171,N_17913);
nor U19169 (N_19169,N_17288,N_17603);
xnor U19170 (N_19170,N_17375,N_17055);
xor U19171 (N_19171,N_17448,N_17050);
nand U19172 (N_19172,N_17524,N_17919);
or U19173 (N_19173,N_17795,N_17876);
xnor U19174 (N_19174,N_17340,N_17280);
nand U19175 (N_19175,N_17061,N_17789);
and U19176 (N_19176,N_17090,N_17897);
xor U19177 (N_19177,N_17448,N_16972);
nand U19178 (N_19178,N_16961,N_16941);
xnor U19179 (N_19179,N_17617,N_17742);
nor U19180 (N_19180,N_16818,N_17112);
nand U19181 (N_19181,N_16878,N_17211);
or U19182 (N_19182,N_17595,N_17357);
or U19183 (N_19183,N_16947,N_16884);
nand U19184 (N_19184,N_16999,N_17559);
and U19185 (N_19185,N_17229,N_17228);
nand U19186 (N_19186,N_17860,N_17566);
nor U19187 (N_19187,N_17256,N_17276);
or U19188 (N_19188,N_17440,N_17834);
or U19189 (N_19189,N_17367,N_16906);
nand U19190 (N_19190,N_17222,N_17240);
and U19191 (N_19191,N_16953,N_17006);
nor U19192 (N_19192,N_17066,N_17337);
or U19193 (N_19193,N_17264,N_17583);
nor U19194 (N_19194,N_17161,N_17260);
or U19195 (N_19195,N_17877,N_17890);
nor U19196 (N_19196,N_16919,N_16824);
xor U19197 (N_19197,N_17249,N_17352);
or U19198 (N_19198,N_16818,N_17880);
nand U19199 (N_19199,N_17145,N_17352);
or U19200 (N_19200,N_19161,N_18644);
nor U19201 (N_19201,N_19001,N_18773);
nand U19202 (N_19202,N_18530,N_18790);
nor U19203 (N_19203,N_19084,N_18088);
nor U19204 (N_19204,N_19171,N_18330);
or U19205 (N_19205,N_18923,N_18612);
nor U19206 (N_19206,N_19131,N_18982);
xor U19207 (N_19207,N_18004,N_18523);
and U19208 (N_19208,N_18502,N_18978);
nand U19209 (N_19209,N_18558,N_19125);
and U19210 (N_19210,N_19118,N_19085);
or U19211 (N_19211,N_18957,N_19182);
nor U19212 (N_19212,N_18181,N_18304);
nor U19213 (N_19213,N_18439,N_18730);
and U19214 (N_19214,N_18930,N_18598);
nor U19215 (N_19215,N_18036,N_19005);
or U19216 (N_19216,N_18652,N_18246);
xor U19217 (N_19217,N_18283,N_19073);
nand U19218 (N_19218,N_18293,N_19071);
or U19219 (N_19219,N_18749,N_18678);
xnor U19220 (N_19220,N_19098,N_18389);
or U19221 (N_19221,N_18115,N_18259);
nor U19222 (N_19222,N_18161,N_18569);
nor U19223 (N_19223,N_18023,N_18087);
nor U19224 (N_19224,N_18603,N_19153);
or U19225 (N_19225,N_19176,N_18463);
and U19226 (N_19226,N_18511,N_18508);
or U19227 (N_19227,N_18316,N_18820);
nor U19228 (N_19228,N_18369,N_18366);
xor U19229 (N_19229,N_18766,N_18361);
and U19230 (N_19230,N_18617,N_18094);
nand U19231 (N_19231,N_19061,N_18198);
nor U19232 (N_19232,N_18725,N_19045);
xnor U19233 (N_19233,N_18012,N_18716);
nand U19234 (N_19234,N_18131,N_18141);
nor U19235 (N_19235,N_18086,N_18883);
xnor U19236 (N_19236,N_18997,N_18777);
nand U19237 (N_19237,N_18681,N_18714);
nor U19238 (N_19238,N_19057,N_18514);
xor U19239 (N_19239,N_19157,N_18970);
and U19240 (N_19240,N_19049,N_18459);
and U19241 (N_19241,N_18256,N_18029);
or U19242 (N_19242,N_19197,N_18679);
nand U19243 (N_19243,N_18143,N_19065);
or U19244 (N_19244,N_18104,N_18755);
nand U19245 (N_19245,N_19166,N_18601);
nor U19246 (N_19246,N_18680,N_18428);
and U19247 (N_19247,N_18183,N_18560);
nor U19248 (N_19248,N_18845,N_18564);
or U19249 (N_19249,N_18000,N_18693);
or U19250 (N_19250,N_18224,N_19081);
xor U19251 (N_19251,N_18656,N_18448);
and U19252 (N_19252,N_18182,N_18387);
nor U19253 (N_19253,N_18265,N_19079);
nor U19254 (N_19254,N_18364,N_18007);
nand U19255 (N_19255,N_19068,N_18362);
or U19256 (N_19256,N_18055,N_18819);
and U19257 (N_19257,N_19123,N_18760);
nand U19258 (N_19258,N_18746,N_18020);
or U19259 (N_19259,N_18273,N_18798);
or U19260 (N_19260,N_18825,N_18894);
nor U19261 (N_19261,N_18778,N_19179);
nor U19262 (N_19262,N_18989,N_18669);
nand U19263 (N_19263,N_18105,N_18724);
nand U19264 (N_19264,N_18675,N_18609);
and U19265 (N_19265,N_18196,N_18538);
nand U19266 (N_19266,N_18578,N_18084);
or U19267 (N_19267,N_18484,N_19192);
nor U19268 (N_19268,N_18706,N_18736);
nor U19269 (N_19269,N_18419,N_18019);
xnor U19270 (N_19270,N_18215,N_18818);
and U19271 (N_19271,N_18945,N_18847);
xnor U19272 (N_19272,N_18791,N_18768);
xor U19273 (N_19273,N_19121,N_18253);
and U19274 (N_19274,N_19052,N_18994);
or U19275 (N_19275,N_19097,N_18507);
nor U19276 (N_19276,N_18067,N_18902);
nor U19277 (N_19277,N_18545,N_18295);
xor U19278 (N_19278,N_18713,N_18535);
nand U19279 (N_19279,N_18310,N_18638);
nor U19280 (N_19280,N_18043,N_18437);
or U19281 (N_19281,N_18835,N_18187);
nand U19282 (N_19282,N_18116,N_18481);
nand U19283 (N_19283,N_18286,N_18103);
or U19284 (N_19284,N_18621,N_18080);
nor U19285 (N_19285,N_18465,N_18026);
and U19286 (N_19286,N_18596,N_19172);
or U19287 (N_19287,N_18168,N_18150);
or U19288 (N_19288,N_18824,N_18261);
nand U19289 (N_19289,N_18301,N_18968);
xor U19290 (N_19290,N_19159,N_19129);
nor U19291 (N_19291,N_18868,N_18738);
xor U19292 (N_19292,N_18775,N_18816);
or U19293 (N_19293,N_18956,N_18157);
or U19294 (N_19294,N_18723,N_18817);
nand U19295 (N_19295,N_18311,N_19195);
or U19296 (N_19296,N_18971,N_18155);
or U19297 (N_19297,N_19196,N_18331);
and U19298 (N_19298,N_19050,N_18173);
and U19299 (N_19299,N_19011,N_18434);
nor U19300 (N_19300,N_18585,N_18660);
xnor U19301 (N_19301,N_18841,N_18472);
and U19302 (N_19302,N_18045,N_18312);
and U19303 (N_19303,N_18221,N_18473);
xor U19304 (N_19304,N_18346,N_18138);
nor U19305 (N_19305,N_19155,N_18061);
nand U19306 (N_19306,N_18489,N_18418);
nor U19307 (N_19307,N_18920,N_18477);
or U19308 (N_19308,N_18880,N_18610);
nand U19309 (N_19309,N_18668,N_18891);
nand U19310 (N_19310,N_19072,N_19189);
nand U19311 (N_19311,N_18344,N_18941);
or U19312 (N_19312,N_18262,N_19037);
nand U19313 (N_19313,N_18862,N_18125);
or U19314 (N_19314,N_18275,N_18276);
or U19315 (N_19315,N_18388,N_18541);
and U19316 (N_19316,N_18915,N_18748);
and U19317 (N_19317,N_18132,N_18258);
nor U19318 (N_19318,N_18497,N_18589);
or U19319 (N_19319,N_18667,N_18453);
or U19320 (N_19320,N_18822,N_18030);
and U19321 (N_19321,N_18436,N_19111);
or U19322 (N_19322,N_18499,N_18355);
nor U19323 (N_19323,N_18863,N_18426);
or U19324 (N_19324,N_19029,N_19027);
nor U19325 (N_19325,N_18544,N_18857);
xor U19326 (N_19326,N_18145,N_18339);
nor U19327 (N_19327,N_19141,N_18254);
nor U19328 (N_19328,N_19115,N_18114);
nor U19329 (N_19329,N_18367,N_18102);
nand U19330 (N_19330,N_19120,N_18573);
xnor U19331 (N_19331,N_18509,N_18600);
nand U19332 (N_19332,N_18995,N_18852);
or U19333 (N_19333,N_19107,N_18910);
nand U19334 (N_19334,N_18397,N_18916);
and U19335 (N_19335,N_18417,N_18976);
nand U19336 (N_19336,N_18718,N_18285);
xor U19337 (N_19337,N_18504,N_18614);
or U19338 (N_19338,N_18303,N_18909);
or U19339 (N_19339,N_19112,N_18129);
nor U19340 (N_19340,N_18851,N_18528);
xor U19341 (N_19341,N_18826,N_18281);
nor U19342 (N_19342,N_18914,N_18540);
or U19343 (N_19343,N_18815,N_18811);
and U19344 (N_19344,N_18800,N_18373);
and U19345 (N_19345,N_18160,N_18284);
and U19346 (N_19346,N_18204,N_18501);
and U19347 (N_19347,N_18767,N_18938);
or U19348 (N_19348,N_18096,N_18185);
nor U19349 (N_19349,N_19038,N_19060);
xor U19350 (N_19350,N_19064,N_18858);
or U19351 (N_19351,N_19100,N_18399);
xnor U19352 (N_19352,N_18118,N_18394);
nand U19353 (N_19353,N_18921,N_19184);
xor U19354 (N_19354,N_18860,N_18289);
or U19355 (N_19355,N_19036,N_18961);
and U19356 (N_19356,N_18733,N_18843);
nand U19357 (N_19357,N_18320,N_18830);
xnor U19358 (N_19358,N_18016,N_18701);
or U19359 (N_19359,N_18209,N_18758);
or U19360 (N_19360,N_18856,N_18873);
and U19361 (N_19361,N_18230,N_19137);
and U19362 (N_19362,N_18005,N_18268);
xnor U19363 (N_19363,N_18604,N_19043);
or U19364 (N_19364,N_18153,N_18586);
nor U19365 (N_19365,N_18377,N_19126);
xnor U19366 (N_19366,N_18567,N_18940);
or U19367 (N_19367,N_18435,N_18510);
nand U19368 (N_19368,N_18280,N_18488);
nand U19369 (N_19369,N_18414,N_19047);
and U19370 (N_19370,N_18939,N_18912);
nor U19371 (N_19371,N_18606,N_18763);
or U19372 (N_19372,N_19133,N_18884);
or U19373 (N_19373,N_18423,N_18451);
nor U19374 (N_19374,N_18047,N_18352);
nand U19375 (N_19375,N_18673,N_18093);
nand U19376 (N_19376,N_18054,N_18443);
nand U19377 (N_19377,N_18454,N_18527);
and U19378 (N_19378,N_18235,N_18290);
nor U19379 (N_19379,N_19076,N_18405);
xnor U19380 (N_19380,N_18799,N_18065);
xor U19381 (N_19381,N_18937,N_18670);
and U19382 (N_19382,N_18711,N_18933);
and U19383 (N_19383,N_18136,N_18082);
nand U19384 (N_19384,N_18892,N_18696);
and U19385 (N_19385,N_19167,N_19173);
nor U19386 (N_19386,N_18123,N_18574);
nor U19387 (N_19387,N_18078,N_18911);
nand U19388 (N_19388,N_18041,N_18079);
nor U19389 (N_19389,N_18383,N_18879);
nand U19390 (N_19390,N_18764,N_18750);
xnor U19391 (N_19391,N_18159,N_18195);
and U19392 (N_19392,N_18844,N_18176);
xnor U19393 (N_19393,N_18270,N_19198);
nor U19394 (N_19394,N_18643,N_18647);
nand U19395 (N_19395,N_18636,N_18877);
xor U19396 (N_19396,N_18650,N_18142);
nor U19397 (N_19397,N_18171,N_18649);
nor U19398 (N_19398,N_19122,N_18406);
nor U19399 (N_19399,N_19128,N_18146);
or U19400 (N_19400,N_19174,N_19130);
nand U19401 (N_19401,N_18611,N_19028);
nor U19402 (N_19402,N_18869,N_18006);
xor U19403 (N_19403,N_18395,N_18101);
and U19404 (N_19404,N_18231,N_18919);
and U19405 (N_19405,N_18404,N_18663);
nor U19406 (N_19406,N_19101,N_18720);
nand U19407 (N_19407,N_18001,N_19096);
nand U19408 (N_19408,N_18515,N_18177);
or U19409 (N_19409,N_19055,N_18687);
xor U19410 (N_19410,N_18039,N_18319);
nand U19411 (N_19411,N_18903,N_18854);
xnor U19412 (N_19412,N_18476,N_19124);
or U19413 (N_19413,N_18987,N_18438);
or U19414 (N_19414,N_19151,N_19010);
nor U19415 (N_19415,N_18003,N_19039);
xnor U19416 (N_19416,N_18154,N_18379);
xor U19417 (N_19417,N_18427,N_18797);
xor U19418 (N_19418,N_18400,N_19062);
nor U19419 (N_19419,N_18552,N_18089);
nand U19420 (N_19420,N_18470,N_18975);
nand U19421 (N_19421,N_19048,N_19178);
xor U19422 (N_19422,N_18240,N_18493);
and U19423 (N_19423,N_19119,N_18949);
nand U19424 (N_19424,N_19144,N_18074);
nand U19425 (N_19425,N_18958,N_18703);
nand U19426 (N_19426,N_18348,N_18278);
xnor U19427 (N_19427,N_18943,N_18809);
and U19428 (N_19428,N_18298,N_18848);
nor U19429 (N_19429,N_18834,N_18492);
xor U19430 (N_19430,N_18186,N_19095);
xor U19431 (N_19431,N_18737,N_18697);
xor U19432 (N_19432,N_18090,N_18532);
nor U19433 (N_19433,N_18324,N_18539);
and U19434 (N_19434,N_19034,N_18429);
and U19435 (N_19435,N_18807,N_18666);
xnor U19436 (N_19436,N_18732,N_18715);
xor U19437 (N_19437,N_18803,N_18068);
xor U19438 (N_19438,N_18672,N_18336);
nand U19439 (N_19439,N_19069,N_18533);
xnor U19440 (N_19440,N_18572,N_18543);
nand U19441 (N_19441,N_18918,N_18009);
xor U19442 (N_19442,N_18467,N_18983);
nand U19443 (N_19443,N_18248,N_19149);
xnor U19444 (N_19444,N_18170,N_18999);
nand U19445 (N_19445,N_18648,N_18833);
xor U19446 (N_19446,N_18842,N_18354);
nor U19447 (N_19447,N_18836,N_18969);
nor U19448 (N_19448,N_18549,N_18486);
or U19449 (N_19449,N_18201,N_18207);
or U19450 (N_19450,N_19083,N_18753);
xnor U19451 (N_19451,N_19185,N_18031);
or U19452 (N_19452,N_18302,N_18024);
nor U19453 (N_19453,N_18683,N_18840);
or U19454 (N_19454,N_18317,N_18602);
nand U19455 (N_19455,N_18318,N_18658);
nand U19456 (N_19456,N_18128,N_18456);
xor U19457 (N_19457,N_18898,N_18148);
nor U19458 (N_19458,N_18942,N_18772);
xnor U19459 (N_19459,N_18895,N_18450);
and U19460 (N_19460,N_18747,N_18049);
and U19461 (N_19461,N_18688,N_18368);
or U19462 (N_19462,N_18013,N_18077);
xor U19463 (N_19463,N_18260,N_19006);
nor U19464 (N_19464,N_18452,N_18927);
and U19465 (N_19465,N_19183,N_18559);
nand U19466 (N_19466,N_18255,N_18010);
xor U19467 (N_19467,N_18085,N_19059);
or U19468 (N_19468,N_18917,N_19113);
nand U19469 (N_19469,N_18751,N_18783);
nor U19470 (N_19470,N_18876,N_18059);
nand U19471 (N_19471,N_18340,N_19041);
or U19472 (N_19472,N_19023,N_18613);
nor U19473 (N_19473,N_18308,N_18924);
or U19474 (N_19474,N_18823,N_19110);
or U19475 (N_19475,N_19152,N_18885);
and U19476 (N_19476,N_18865,N_18689);
nor U19477 (N_19477,N_18358,N_18622);
nand U19478 (N_19478,N_18200,N_18113);
and U19479 (N_19479,N_18222,N_18482);
or U19480 (N_19480,N_18162,N_18037);
xor U19481 (N_19481,N_18487,N_18430);
xnor U19482 (N_19482,N_18011,N_18223);
nor U19483 (N_19483,N_18050,N_19088);
nand U19484 (N_19484,N_18735,N_18237);
or U19485 (N_19485,N_18321,N_18208);
or U19486 (N_19486,N_18882,N_19134);
and U19487 (N_19487,N_18557,N_19007);
and U19488 (N_19488,N_18070,N_19024);
nand U19489 (N_19489,N_18306,N_18710);
and U19490 (N_19490,N_18812,N_18402);
xor U19491 (N_19491,N_18591,N_19044);
nand U19492 (N_19492,N_18788,N_18676);
and U19493 (N_19493,N_19074,N_18126);
xor U19494 (N_19494,N_18634,N_19075);
nand U19495 (N_19495,N_18568,N_18855);
and U19496 (N_19496,N_18002,N_19117);
and U19497 (N_19497,N_18657,N_18233);
nor U19498 (N_19498,N_18627,N_18794);
xor U19499 (N_19499,N_18517,N_18785);
nand U19500 (N_19500,N_18360,N_19106);
nand U19501 (N_19501,N_18722,N_18092);
and U19502 (N_19502,N_18684,N_18151);
xor U19503 (N_19503,N_18900,N_18471);
nand U19504 (N_19504,N_18172,N_18334);
xnor U19505 (N_19505,N_18875,N_18806);
or U19506 (N_19506,N_18391,N_19013);
nand U19507 (N_19507,N_19066,N_19156);
or U19508 (N_19508,N_18595,N_18828);
nor U19509 (N_19509,N_18386,N_18106);
and U19510 (N_19510,N_18274,N_18158);
nor U19511 (N_19511,N_19033,N_19032);
xor U19512 (N_19512,N_18707,N_19019);
nand U19513 (N_19513,N_18227,N_18769);
and U19514 (N_19514,N_18731,N_18069);
nor U19515 (N_19515,N_18372,N_18594);
or U19516 (N_19516,N_19163,N_18421);
nand U19517 (N_19517,N_18135,N_18793);
or U19518 (N_19518,N_18469,N_18562);
nand U19519 (N_19519,N_18531,N_18887);
nand U19520 (N_19520,N_19188,N_18294);
and U19521 (N_19521,N_19168,N_19132);
or U19522 (N_19522,N_18440,N_18546);
and U19523 (N_19523,N_18690,N_18712);
xor U19524 (N_19524,N_18149,N_18871);
nand U19525 (N_19525,N_19016,N_18174);
xnor U19526 (N_19526,N_18639,N_18365);
or U19527 (N_19527,N_19143,N_19046);
or U19528 (N_19528,N_18188,N_18433);
nand U19529 (N_19529,N_18313,N_19051);
and U19530 (N_19530,N_18651,N_18382);
and U19531 (N_19531,N_18385,N_18808);
or U19532 (N_19532,N_18581,N_18446);
xnor U19533 (N_19533,N_18555,N_18139);
and U19534 (N_19534,N_18163,N_18359);
xnor U19535 (N_19535,N_18014,N_18027);
nor U19536 (N_19536,N_18770,N_19147);
nand U19537 (N_19537,N_18315,N_18225);
and U19538 (N_19538,N_18759,N_18682);
nor U19539 (N_19539,N_18152,N_18872);
nand U19540 (N_19540,N_19099,N_18130);
or U19541 (N_19541,N_18109,N_18122);
nor U19542 (N_19542,N_18287,N_19080);
or U19543 (N_19543,N_18955,N_19004);
and U19544 (N_19544,N_18973,N_18121);
nor U19545 (N_19545,N_18455,N_18058);
and U19546 (N_19546,N_18893,N_19053);
xnor U19547 (N_19547,N_18214,N_18035);
and U19548 (N_19548,N_18277,N_18959);
or U19549 (N_19549,N_18616,N_18953);
nand U19550 (N_19550,N_18859,N_19021);
and U19551 (N_19551,N_18789,N_18717);
or U19552 (N_19552,N_18063,N_19093);
nand U19553 (N_19553,N_18513,N_18846);
nand U19554 (N_19554,N_18963,N_19140);
or U19555 (N_19555,N_18947,N_18708);
or U19556 (N_19556,N_18242,N_18584);
xor U19557 (N_19557,N_18017,N_18980);
nand U19558 (N_19558,N_19089,N_18700);
or U19559 (N_19559,N_18252,N_18357);
nor U19560 (N_19560,N_18580,N_18795);
or U19561 (N_19561,N_18787,N_18076);
nor U19562 (N_19562,N_18996,N_18083);
and U19563 (N_19563,N_18028,N_18642);
and U19564 (N_19564,N_19003,N_18761);
xnor U19565 (N_19565,N_18889,N_18038);
nand U19566 (N_19566,N_18662,N_19162);
or U19567 (N_19567,N_18550,N_19114);
nand U19568 (N_19568,N_18444,N_19177);
nand U19569 (N_19569,N_18468,N_18740);
nand U19570 (N_19570,N_18694,N_18951);
xor U19571 (N_19571,N_19090,N_18279);
and U19572 (N_19572,N_19077,N_18991);
nand U19573 (N_19573,N_18098,N_19150);
xnor U19574 (N_19574,N_18743,N_18810);
and U19575 (N_19575,N_18491,N_19104);
nand U19576 (N_19576,N_18590,N_18551);
or U19577 (N_19577,N_18219,N_18754);
nand U19578 (N_19578,N_18837,N_18520);
nor U19579 (N_19579,N_18349,N_18403);
and U19580 (N_19580,N_18623,N_18380);
nor U19581 (N_19581,N_19063,N_18202);
or U19582 (N_19582,N_18992,N_18905);
nor U19583 (N_19583,N_18292,N_18625);
nand U19584 (N_19584,N_18250,N_18588);
or U19585 (N_19585,N_18374,N_19139);
and U19586 (N_19586,N_18140,N_18322);
and U19587 (N_19587,N_18906,N_18044);
xor U19588 (N_19588,N_18111,N_18480);
nand U19589 (N_19589,N_18052,N_18345);
and U19590 (N_19590,N_18247,N_18952);
or U19591 (N_19591,N_19181,N_18529);
nand U19592 (N_19592,N_18351,N_18375);
and U19593 (N_19593,N_18966,N_18674);
nor U19594 (N_19594,N_18032,N_18704);
nand U19595 (N_19595,N_18053,N_18757);
nand U19596 (N_19596,N_18212,N_18282);
nand U19597 (N_19597,N_18516,N_18946);
xnor U19598 (N_19598,N_18021,N_18494);
nor U19599 (N_19599,N_18099,N_18691);
nand U19600 (N_19600,N_18587,N_18727);
nor U19601 (N_19601,N_18108,N_18781);
nor U19602 (N_19602,N_18630,N_18525);
xor U19603 (N_19603,N_18665,N_18653);
and U19604 (N_19604,N_18926,N_18695);
or U19605 (N_19605,N_18363,N_19040);
and U19606 (N_19606,N_18408,N_19002);
or U19607 (N_19607,N_18305,N_18948);
or U19608 (N_19608,N_18137,N_18178);
nand U19609 (N_19609,N_18620,N_18015);
and U19610 (N_19610,N_18742,N_18729);
nand U19611 (N_19611,N_18641,N_19078);
nor U19612 (N_19612,N_18447,N_18821);
and U19613 (N_19613,N_18441,N_19025);
nand U19614 (N_19614,N_18888,N_18928);
and U19615 (N_19615,N_19190,N_18156);
nand U19616 (N_19616,N_18271,N_18503);
and U19617 (N_19617,N_18234,N_18461);
xnor U19618 (N_19618,N_18300,N_18583);
or U19619 (N_19619,N_18291,N_18025);
nand U19620 (N_19620,N_19135,N_18018);
xnor U19621 (N_19621,N_18378,N_19070);
nor U19622 (N_19622,N_18734,N_18190);
and U19623 (N_19623,N_19169,N_18107);
nand U19624 (N_19624,N_18536,N_18936);
or U19625 (N_19625,N_18640,N_18495);
nand U19626 (N_19626,N_18901,N_18565);
xnor U19627 (N_19627,N_18519,N_18460);
nand U19628 (N_19628,N_18985,N_18561);
xor U19629 (N_19629,N_18745,N_18206);
or U19630 (N_19630,N_18288,N_19180);
or U19631 (N_19631,N_18422,N_18328);
or U19632 (N_19632,N_18332,N_18164);
or U19633 (N_19633,N_18095,N_18243);
and U19634 (N_19634,N_18576,N_19103);
nor U19635 (N_19635,N_18496,N_18479);
xnor U19636 (N_19636,N_19020,N_18297);
nor U19637 (N_19637,N_18205,N_18904);
and U19638 (N_19638,N_18197,N_18213);
xnor U19639 (N_19639,N_18390,N_18827);
nor U19640 (N_19640,N_19154,N_18605);
xor U19641 (N_19641,N_18582,N_18542);
nand U19642 (N_19642,N_18804,N_18593);
nor U19643 (N_19643,N_18442,N_18409);
nand U19644 (N_19644,N_18081,N_18629);
nand U19645 (N_19645,N_18048,N_18878);
nor U19646 (N_19646,N_18864,N_18376);
xor U19647 (N_19647,N_18124,N_18784);
nand U19648 (N_19648,N_18051,N_18786);
and U19649 (N_19649,N_18342,N_18624);
xor U19650 (N_19650,N_18654,N_18986);
and U19651 (N_19651,N_18415,N_19187);
nor U19652 (N_19652,N_18343,N_18338);
or U19653 (N_19653,N_18776,N_18432);
xor U19654 (N_19654,N_18272,N_18655);
nand U19655 (N_19655,N_18522,N_19105);
or U19656 (N_19656,N_19022,N_18210);
nor U19657 (N_19657,N_18180,N_19015);
and U19658 (N_19658,N_18072,N_18896);
nor U19659 (N_19659,N_18686,N_18239);
nor U19660 (N_19660,N_18042,N_18922);
xnor U19661 (N_19661,N_19026,N_19058);
and U19662 (N_19662,N_18412,N_18179);
or U19663 (N_19663,N_18431,N_18474);
and U19664 (N_19664,N_18333,N_19146);
and U19665 (N_19665,N_18218,N_19091);
nand U19666 (N_19666,N_18466,N_19087);
and U19667 (N_19667,N_18034,N_18579);
nand U19668 (N_19668,N_18245,N_18309);
or U19669 (N_19669,N_18908,N_18597);
and U19670 (N_19670,N_18796,N_18972);
nand U19671 (N_19671,N_19030,N_18886);
and U19672 (N_19672,N_19138,N_18782);
or U19673 (N_19673,N_18685,N_18500);
nor U19674 (N_19674,N_18608,N_18838);
and U19675 (N_19675,N_19193,N_18269);
xnor U19676 (N_19676,N_18850,N_18792);
nand U19677 (N_19677,N_18802,N_18392);
nand U19678 (N_19678,N_18066,N_18954);
and U19679 (N_19679,N_18897,N_18192);
xor U19680 (N_19680,N_18698,N_18692);
and U19681 (N_19681,N_18512,N_18547);
xor U19682 (N_19682,N_18478,N_18134);
xnor U19683 (N_19683,N_19191,N_18238);
nor U19684 (N_19684,N_18853,N_18671);
nand U19685 (N_19685,N_18416,N_18267);
and U19686 (N_19686,N_18607,N_18341);
nand U19687 (N_19687,N_18299,N_18563);
nand U19688 (N_19688,N_19009,N_18073);
and U19689 (N_19689,N_18988,N_18216);
or U19690 (N_19690,N_18762,N_19067);
or U19691 (N_19691,N_18490,N_18813);
nand U19692 (N_19692,N_18964,N_18890);
xnor U19693 (N_19693,N_18524,N_18229);
nand U19694 (N_19694,N_19194,N_18147);
nand U19695 (N_19695,N_18350,N_19142);
and U19696 (N_19696,N_19136,N_18483);
xor U19697 (N_19697,N_18119,N_18257);
nand U19698 (N_19698,N_18064,N_18424);
nor U19699 (N_19699,N_19012,N_18618);
nor U19700 (N_19700,N_18194,N_18022);
nand U19701 (N_19701,N_19035,N_18075);
xnor U19702 (N_19702,N_18993,N_18571);
xor U19703 (N_19703,N_18475,N_18220);
nand U19704 (N_19704,N_18445,N_18008);
and U19705 (N_19705,N_18805,N_19199);
nor U19706 (N_19706,N_18485,N_18719);
nand U19707 (N_19707,N_18420,N_18832);
or U19708 (N_19708,N_18981,N_18323);
xnor U19709 (N_19709,N_18849,N_18457);
xnor U19710 (N_19710,N_18203,N_18347);
or U19711 (N_19711,N_18449,N_18033);
or U19712 (N_19712,N_19175,N_18913);
and U19713 (N_19713,N_18633,N_18548);
nor U19714 (N_19714,N_18464,N_18867);
nand U19715 (N_19715,N_18244,N_18353);
or U19716 (N_19716,N_18709,N_18425);
or U19717 (N_19717,N_18296,N_18556);
and U19718 (N_19718,N_18866,N_19082);
nand U19719 (N_19719,N_18057,N_18756);
and U19720 (N_19720,N_18040,N_18071);
or U19721 (N_19721,N_18839,N_18950);
and U19722 (N_19722,N_18046,N_18396);
and U19723 (N_19723,N_19086,N_18314);
xnor U19724 (N_19724,N_18199,N_18765);
nor U19725 (N_19725,N_18251,N_19127);
nor U19726 (N_19726,N_18506,N_18091);
nand U19727 (N_19727,N_18702,N_18193);
and U19728 (N_19728,N_18191,N_18967);
and U19729 (N_19729,N_18398,N_18599);
nor U19730 (N_19730,N_18325,N_18554);
xor U19731 (N_19731,N_19145,N_18631);
or U19732 (N_19732,N_18741,N_19170);
nor U19733 (N_19733,N_18829,N_18411);
and U19734 (N_19734,N_19017,N_18381);
and U19735 (N_19735,N_18175,N_18167);
and U19736 (N_19736,N_18166,N_18677);
or U19737 (N_19737,N_18184,N_19109);
nand U19738 (N_19738,N_18521,N_18100);
xnor U19739 (N_19739,N_18659,N_19116);
nand U19740 (N_19740,N_18577,N_19186);
xnor U19741 (N_19741,N_18780,N_18728);
and U19742 (N_19742,N_18413,N_18744);
or U19743 (N_19743,N_19158,N_18371);
or U19744 (N_19744,N_19164,N_19042);
xor U19745 (N_19745,N_18998,N_18518);
nor U19746 (N_19746,N_18356,N_18266);
and U19747 (N_19747,N_18726,N_18637);
or U19748 (N_19748,N_18870,N_18979);
nand U19749 (N_19749,N_18635,N_19092);
and U19750 (N_19750,N_19102,N_18228);
nand U19751 (N_19751,N_18505,N_18097);
xnor U19752 (N_19752,N_19094,N_18127);
nor U19753 (N_19753,N_18984,N_18335);
and U19754 (N_19754,N_18462,N_18615);
nor U19755 (N_19755,N_18189,N_18056);
nand U19756 (N_19756,N_18570,N_18337);
nor U19757 (N_19757,N_19148,N_18752);
xnor U19758 (N_19758,N_18329,N_19018);
nor U19759 (N_19759,N_19008,N_18169);
and U19760 (N_19760,N_18165,N_18393);
and U19761 (N_19761,N_18661,N_18628);
xor U19762 (N_19762,N_19031,N_19056);
nand U19763 (N_19763,N_18407,N_18774);
and U19764 (N_19764,N_18960,N_18944);
nor U19765 (N_19765,N_18384,N_18327);
or U19766 (N_19766,N_19165,N_18932);
nand U19767 (N_19767,N_18120,N_18526);
nor U19768 (N_19768,N_18632,N_18112);
nand U19769 (N_19769,N_18133,N_19108);
nand U19770 (N_19770,N_18929,N_18934);
or U19771 (N_19771,N_18907,N_18935);
nand U19772 (N_19772,N_18779,N_18699);
and U19773 (N_19773,N_18232,N_18861);
nor U19774 (N_19774,N_18974,N_18801);
nor U19775 (N_19775,N_18771,N_19160);
or U19776 (N_19776,N_18370,N_18241);
nor U19777 (N_19777,N_18962,N_18217);
xor U19778 (N_19778,N_18925,N_18874);
nand U19779 (N_19779,N_18965,N_18990);
xnor U19780 (N_19780,N_18211,N_18881);
nand U19781 (N_19781,N_18739,N_18831);
nor U19782 (N_19782,N_18619,N_18534);
nor U19783 (N_19783,N_18249,N_19000);
xor U19784 (N_19784,N_18931,N_18553);
xnor U19785 (N_19785,N_18646,N_18263);
xor U19786 (N_19786,N_19014,N_18401);
and U19787 (N_19787,N_19054,N_18705);
xor U19788 (N_19788,N_18264,N_18458);
and U19789 (N_19789,N_18062,N_18060);
or U19790 (N_19790,N_18664,N_18566);
nand U19791 (N_19791,N_18226,N_18110);
nor U19792 (N_19792,N_18537,N_18236);
xnor U19793 (N_19793,N_18899,N_18326);
and U19794 (N_19794,N_18721,N_18814);
xor U19795 (N_19795,N_18144,N_18307);
nand U19796 (N_19796,N_18575,N_18410);
nor U19797 (N_19797,N_18977,N_18117);
or U19798 (N_19798,N_18498,N_18592);
xor U19799 (N_19799,N_18626,N_18645);
or U19800 (N_19800,N_18014,N_18162);
nor U19801 (N_19801,N_19091,N_18420);
and U19802 (N_19802,N_18864,N_18096);
or U19803 (N_19803,N_18491,N_18668);
nand U19804 (N_19804,N_18920,N_18848);
and U19805 (N_19805,N_18826,N_18457);
nand U19806 (N_19806,N_18991,N_18146);
or U19807 (N_19807,N_18854,N_18149);
and U19808 (N_19808,N_18743,N_18455);
or U19809 (N_19809,N_18184,N_18980);
xor U19810 (N_19810,N_18631,N_18600);
and U19811 (N_19811,N_18074,N_18958);
xnor U19812 (N_19812,N_18449,N_18940);
nor U19813 (N_19813,N_19142,N_18495);
and U19814 (N_19814,N_18168,N_18016);
nand U19815 (N_19815,N_19068,N_18265);
and U19816 (N_19816,N_19085,N_18269);
xnor U19817 (N_19817,N_18561,N_18630);
nor U19818 (N_19818,N_18519,N_18161);
xor U19819 (N_19819,N_18616,N_18096);
nor U19820 (N_19820,N_19155,N_18821);
xor U19821 (N_19821,N_18997,N_18208);
nor U19822 (N_19822,N_19164,N_18963);
nor U19823 (N_19823,N_18741,N_19196);
xor U19824 (N_19824,N_18227,N_18633);
xor U19825 (N_19825,N_18660,N_18348);
nor U19826 (N_19826,N_18799,N_18473);
nor U19827 (N_19827,N_18696,N_18482);
nor U19828 (N_19828,N_18119,N_18642);
xnor U19829 (N_19829,N_19026,N_18675);
and U19830 (N_19830,N_18447,N_18672);
nand U19831 (N_19831,N_18002,N_19074);
and U19832 (N_19832,N_18662,N_18659);
and U19833 (N_19833,N_18470,N_18962);
nand U19834 (N_19834,N_18059,N_18974);
nand U19835 (N_19835,N_18294,N_18139);
xor U19836 (N_19836,N_18143,N_18908);
nor U19837 (N_19837,N_18920,N_19097);
or U19838 (N_19838,N_18229,N_18384);
nand U19839 (N_19839,N_18363,N_18159);
nand U19840 (N_19840,N_19113,N_18926);
or U19841 (N_19841,N_18007,N_18733);
nand U19842 (N_19842,N_18964,N_18683);
nor U19843 (N_19843,N_19146,N_18196);
and U19844 (N_19844,N_18309,N_18083);
nand U19845 (N_19845,N_18168,N_19012);
xor U19846 (N_19846,N_18860,N_19193);
or U19847 (N_19847,N_18959,N_18331);
nand U19848 (N_19848,N_18712,N_19096);
xor U19849 (N_19849,N_18233,N_18688);
nor U19850 (N_19850,N_18727,N_19053);
nor U19851 (N_19851,N_18634,N_18148);
or U19852 (N_19852,N_18935,N_18752);
or U19853 (N_19853,N_19038,N_18347);
nor U19854 (N_19854,N_18752,N_18512);
and U19855 (N_19855,N_19077,N_18912);
xnor U19856 (N_19856,N_19153,N_18240);
or U19857 (N_19857,N_18384,N_18591);
xnor U19858 (N_19858,N_18541,N_18014);
nor U19859 (N_19859,N_18535,N_18703);
or U19860 (N_19860,N_18265,N_18632);
nor U19861 (N_19861,N_18484,N_19190);
nor U19862 (N_19862,N_18537,N_18156);
nor U19863 (N_19863,N_18966,N_18906);
or U19864 (N_19864,N_18550,N_19066);
nand U19865 (N_19865,N_19155,N_18548);
and U19866 (N_19866,N_19089,N_18074);
nor U19867 (N_19867,N_18780,N_18031);
nand U19868 (N_19868,N_18087,N_18877);
nor U19869 (N_19869,N_18833,N_18470);
and U19870 (N_19870,N_18872,N_18141);
nand U19871 (N_19871,N_19002,N_18366);
or U19872 (N_19872,N_18414,N_19100);
xnor U19873 (N_19873,N_18859,N_18235);
xnor U19874 (N_19874,N_18731,N_19021);
and U19875 (N_19875,N_18805,N_18170);
nor U19876 (N_19876,N_18863,N_18896);
nand U19877 (N_19877,N_18749,N_18930);
or U19878 (N_19878,N_18644,N_18515);
xor U19879 (N_19879,N_19145,N_18568);
or U19880 (N_19880,N_18711,N_18079);
nor U19881 (N_19881,N_18905,N_18397);
and U19882 (N_19882,N_18931,N_18732);
xor U19883 (N_19883,N_19090,N_18030);
nor U19884 (N_19884,N_19190,N_19052);
and U19885 (N_19885,N_19058,N_18532);
nor U19886 (N_19886,N_18568,N_19194);
nor U19887 (N_19887,N_18526,N_18685);
or U19888 (N_19888,N_18792,N_18705);
nor U19889 (N_19889,N_18246,N_18577);
xor U19890 (N_19890,N_19014,N_18830);
nor U19891 (N_19891,N_19164,N_18957);
nand U19892 (N_19892,N_18115,N_19135);
xnor U19893 (N_19893,N_18611,N_18252);
xnor U19894 (N_19894,N_18112,N_18178);
and U19895 (N_19895,N_18174,N_19010);
nand U19896 (N_19896,N_19125,N_18644);
nor U19897 (N_19897,N_18379,N_18092);
nor U19898 (N_19898,N_18678,N_18133);
and U19899 (N_19899,N_18782,N_18010);
nor U19900 (N_19900,N_18391,N_18803);
nand U19901 (N_19901,N_18998,N_18352);
xor U19902 (N_19902,N_18765,N_18007);
or U19903 (N_19903,N_18683,N_19026);
or U19904 (N_19904,N_19103,N_18684);
and U19905 (N_19905,N_18713,N_18196);
nor U19906 (N_19906,N_18488,N_18999);
and U19907 (N_19907,N_18254,N_18765);
xor U19908 (N_19908,N_19097,N_18697);
nand U19909 (N_19909,N_18069,N_18788);
xor U19910 (N_19910,N_18776,N_18640);
or U19911 (N_19911,N_19063,N_18164);
nor U19912 (N_19912,N_18905,N_18951);
nand U19913 (N_19913,N_18810,N_18444);
nand U19914 (N_19914,N_18470,N_19128);
xor U19915 (N_19915,N_18972,N_18775);
nand U19916 (N_19916,N_18686,N_18342);
or U19917 (N_19917,N_18076,N_19068);
nand U19918 (N_19918,N_18679,N_18286);
xor U19919 (N_19919,N_18223,N_18696);
nand U19920 (N_19920,N_19195,N_18152);
or U19921 (N_19921,N_18542,N_19152);
and U19922 (N_19922,N_18387,N_18299);
xnor U19923 (N_19923,N_18914,N_18556);
nor U19924 (N_19924,N_19150,N_18751);
nor U19925 (N_19925,N_18461,N_18512);
nand U19926 (N_19926,N_18389,N_19092);
xnor U19927 (N_19927,N_18330,N_18917);
nor U19928 (N_19928,N_19130,N_18017);
or U19929 (N_19929,N_19174,N_18560);
and U19930 (N_19930,N_19009,N_18788);
or U19931 (N_19931,N_18748,N_18769);
nand U19932 (N_19932,N_18403,N_18260);
or U19933 (N_19933,N_18655,N_18791);
xnor U19934 (N_19934,N_18319,N_19088);
and U19935 (N_19935,N_18712,N_18155);
or U19936 (N_19936,N_18536,N_18445);
nor U19937 (N_19937,N_18637,N_18914);
nand U19938 (N_19938,N_18922,N_18197);
nand U19939 (N_19939,N_18823,N_19066);
xnor U19940 (N_19940,N_18415,N_18177);
nand U19941 (N_19941,N_18320,N_18657);
or U19942 (N_19942,N_18949,N_19009);
or U19943 (N_19943,N_18134,N_19013);
and U19944 (N_19944,N_18670,N_18006);
xnor U19945 (N_19945,N_19095,N_18914);
nand U19946 (N_19946,N_18521,N_18372);
and U19947 (N_19947,N_18424,N_18832);
nand U19948 (N_19948,N_18714,N_18571);
xor U19949 (N_19949,N_19163,N_18672);
nor U19950 (N_19950,N_19091,N_18746);
nand U19951 (N_19951,N_19045,N_18505);
nand U19952 (N_19952,N_19120,N_18999);
nor U19953 (N_19953,N_18922,N_18686);
xnor U19954 (N_19954,N_18390,N_18703);
nor U19955 (N_19955,N_18552,N_18349);
and U19956 (N_19956,N_18414,N_18617);
nor U19957 (N_19957,N_18906,N_18510);
or U19958 (N_19958,N_18725,N_18046);
or U19959 (N_19959,N_18208,N_18011);
nand U19960 (N_19960,N_19157,N_18299);
nor U19961 (N_19961,N_19141,N_18077);
and U19962 (N_19962,N_19041,N_18116);
nand U19963 (N_19963,N_19026,N_18574);
or U19964 (N_19964,N_18368,N_18610);
and U19965 (N_19965,N_18042,N_18965);
nor U19966 (N_19966,N_18364,N_18625);
or U19967 (N_19967,N_19030,N_18729);
xor U19968 (N_19968,N_18809,N_18307);
nor U19969 (N_19969,N_18720,N_18459);
nand U19970 (N_19970,N_18123,N_18327);
nand U19971 (N_19971,N_18207,N_18196);
nand U19972 (N_19972,N_18475,N_18818);
nor U19973 (N_19973,N_18079,N_18135);
and U19974 (N_19974,N_18647,N_18519);
and U19975 (N_19975,N_19196,N_19065);
and U19976 (N_19976,N_18322,N_18811);
or U19977 (N_19977,N_18533,N_18528);
and U19978 (N_19978,N_18821,N_18126);
or U19979 (N_19979,N_18009,N_18644);
nand U19980 (N_19980,N_19189,N_18931);
nor U19981 (N_19981,N_18059,N_19045);
or U19982 (N_19982,N_18027,N_18743);
xnor U19983 (N_19983,N_18424,N_18778);
and U19984 (N_19984,N_18560,N_18582);
or U19985 (N_19985,N_18982,N_18269);
nand U19986 (N_19986,N_18314,N_18095);
and U19987 (N_19987,N_19034,N_18991);
nand U19988 (N_19988,N_18181,N_18355);
and U19989 (N_19989,N_18596,N_18139);
or U19990 (N_19990,N_18090,N_19081);
or U19991 (N_19991,N_18283,N_18736);
and U19992 (N_19992,N_18689,N_18694);
nor U19993 (N_19993,N_18716,N_18575);
nor U19994 (N_19994,N_18769,N_19018);
and U19995 (N_19995,N_18739,N_18261);
and U19996 (N_19996,N_19052,N_19142);
or U19997 (N_19997,N_18642,N_18546);
and U19998 (N_19998,N_18864,N_18545);
nor U19999 (N_19999,N_18695,N_18639);
nor U20000 (N_20000,N_18094,N_18905);
xnor U20001 (N_20001,N_18951,N_18631);
or U20002 (N_20002,N_18738,N_18405);
nor U20003 (N_20003,N_18766,N_18611);
and U20004 (N_20004,N_18197,N_18020);
nand U20005 (N_20005,N_18164,N_18287);
nand U20006 (N_20006,N_18963,N_18032);
nor U20007 (N_20007,N_18350,N_18913);
nand U20008 (N_20008,N_18267,N_18888);
nor U20009 (N_20009,N_19189,N_18282);
nand U20010 (N_20010,N_18104,N_18504);
and U20011 (N_20011,N_18460,N_18642);
or U20012 (N_20012,N_18501,N_18710);
nor U20013 (N_20013,N_19079,N_18169);
or U20014 (N_20014,N_19036,N_19013);
nor U20015 (N_20015,N_18662,N_18701);
nand U20016 (N_20016,N_18460,N_18205);
or U20017 (N_20017,N_18695,N_18541);
nor U20018 (N_20018,N_18552,N_18487);
or U20019 (N_20019,N_18772,N_18078);
or U20020 (N_20020,N_18198,N_18515);
xnor U20021 (N_20021,N_18313,N_18272);
nor U20022 (N_20022,N_18789,N_18376);
xnor U20023 (N_20023,N_18133,N_18138);
or U20024 (N_20024,N_18996,N_19079);
nor U20025 (N_20025,N_18152,N_18875);
and U20026 (N_20026,N_18339,N_19173);
nand U20027 (N_20027,N_18097,N_18826);
or U20028 (N_20028,N_18872,N_19018);
xor U20029 (N_20029,N_19055,N_18758);
nand U20030 (N_20030,N_18603,N_18780);
xor U20031 (N_20031,N_18912,N_19059);
nand U20032 (N_20032,N_18182,N_18660);
nor U20033 (N_20033,N_18608,N_18606);
or U20034 (N_20034,N_18414,N_18622);
or U20035 (N_20035,N_18293,N_18144);
nand U20036 (N_20036,N_18455,N_18318);
or U20037 (N_20037,N_18022,N_18161);
nand U20038 (N_20038,N_18378,N_18097);
or U20039 (N_20039,N_18429,N_18138);
nand U20040 (N_20040,N_18167,N_18308);
xnor U20041 (N_20041,N_18447,N_18906);
nor U20042 (N_20042,N_18725,N_18433);
nand U20043 (N_20043,N_19018,N_18756);
nor U20044 (N_20044,N_19180,N_18380);
and U20045 (N_20045,N_18904,N_18848);
nand U20046 (N_20046,N_18094,N_18486);
xnor U20047 (N_20047,N_19133,N_18846);
xnor U20048 (N_20048,N_18891,N_18064);
nor U20049 (N_20049,N_18292,N_18549);
nor U20050 (N_20050,N_18955,N_18059);
or U20051 (N_20051,N_19044,N_18873);
xnor U20052 (N_20052,N_18082,N_18937);
nor U20053 (N_20053,N_18970,N_18330);
or U20054 (N_20054,N_19020,N_19029);
xnor U20055 (N_20055,N_18111,N_18336);
nand U20056 (N_20056,N_19144,N_18981);
or U20057 (N_20057,N_18114,N_19082);
nor U20058 (N_20058,N_18303,N_18000);
xnor U20059 (N_20059,N_18633,N_18656);
or U20060 (N_20060,N_18322,N_18754);
and U20061 (N_20061,N_18746,N_18247);
xor U20062 (N_20062,N_18245,N_18105);
xor U20063 (N_20063,N_18899,N_18909);
nor U20064 (N_20064,N_18749,N_18048);
nor U20065 (N_20065,N_18768,N_18868);
and U20066 (N_20066,N_19177,N_19142);
and U20067 (N_20067,N_18503,N_18832);
xnor U20068 (N_20068,N_19032,N_18962);
nand U20069 (N_20069,N_18998,N_18923);
nand U20070 (N_20070,N_18928,N_18347);
and U20071 (N_20071,N_19097,N_18653);
nand U20072 (N_20072,N_18895,N_18959);
xor U20073 (N_20073,N_18567,N_18329);
or U20074 (N_20074,N_18104,N_18615);
nand U20075 (N_20075,N_19059,N_19146);
and U20076 (N_20076,N_18025,N_18372);
and U20077 (N_20077,N_18671,N_18246);
nand U20078 (N_20078,N_19086,N_18362);
nor U20079 (N_20079,N_18061,N_18308);
or U20080 (N_20080,N_18866,N_18537);
and U20081 (N_20081,N_18743,N_18996);
xor U20082 (N_20082,N_18699,N_19011);
and U20083 (N_20083,N_18303,N_19044);
xor U20084 (N_20084,N_18390,N_18874);
nand U20085 (N_20085,N_18064,N_18448);
xor U20086 (N_20086,N_18392,N_18649);
xor U20087 (N_20087,N_18991,N_18782);
or U20088 (N_20088,N_18563,N_18617);
or U20089 (N_20089,N_18230,N_18538);
nand U20090 (N_20090,N_18682,N_19051);
nor U20091 (N_20091,N_18883,N_18109);
or U20092 (N_20092,N_18446,N_18515);
or U20093 (N_20093,N_18057,N_19169);
nor U20094 (N_20094,N_18680,N_18817);
xnor U20095 (N_20095,N_18791,N_18685);
nor U20096 (N_20096,N_18104,N_18981);
nand U20097 (N_20097,N_19099,N_18009);
xor U20098 (N_20098,N_18714,N_18977);
nor U20099 (N_20099,N_18420,N_18399);
nand U20100 (N_20100,N_18922,N_18924);
nand U20101 (N_20101,N_19109,N_18773);
nor U20102 (N_20102,N_19160,N_19184);
xor U20103 (N_20103,N_19192,N_18369);
nand U20104 (N_20104,N_18905,N_19102);
or U20105 (N_20105,N_18776,N_18991);
or U20106 (N_20106,N_18230,N_18366);
or U20107 (N_20107,N_19178,N_18178);
nor U20108 (N_20108,N_18707,N_19137);
nor U20109 (N_20109,N_18093,N_18547);
or U20110 (N_20110,N_18822,N_19125);
or U20111 (N_20111,N_18084,N_18249);
nand U20112 (N_20112,N_18175,N_18555);
nand U20113 (N_20113,N_18448,N_19084);
xor U20114 (N_20114,N_18548,N_18464);
and U20115 (N_20115,N_18948,N_18558);
nand U20116 (N_20116,N_18187,N_18597);
nand U20117 (N_20117,N_18494,N_18787);
or U20118 (N_20118,N_18872,N_18090);
nor U20119 (N_20119,N_18841,N_18548);
nor U20120 (N_20120,N_18163,N_18200);
nand U20121 (N_20121,N_18271,N_18203);
xnor U20122 (N_20122,N_18429,N_18723);
nand U20123 (N_20123,N_19102,N_18836);
nand U20124 (N_20124,N_18324,N_18154);
and U20125 (N_20125,N_18618,N_18138);
nor U20126 (N_20126,N_18099,N_18981);
xor U20127 (N_20127,N_18296,N_18226);
nand U20128 (N_20128,N_19003,N_19105);
nand U20129 (N_20129,N_18323,N_18944);
nor U20130 (N_20130,N_18386,N_18959);
and U20131 (N_20131,N_18212,N_18202);
nand U20132 (N_20132,N_18366,N_18595);
nand U20133 (N_20133,N_18704,N_18315);
or U20134 (N_20134,N_18567,N_18424);
nand U20135 (N_20135,N_18056,N_18013);
xnor U20136 (N_20136,N_18061,N_18072);
and U20137 (N_20137,N_18777,N_18541);
or U20138 (N_20138,N_18941,N_19146);
xor U20139 (N_20139,N_18314,N_18887);
or U20140 (N_20140,N_18491,N_18966);
nand U20141 (N_20141,N_18834,N_19167);
nor U20142 (N_20142,N_18991,N_18592);
nand U20143 (N_20143,N_18057,N_18846);
or U20144 (N_20144,N_18756,N_18275);
and U20145 (N_20145,N_18922,N_18338);
xor U20146 (N_20146,N_18854,N_18807);
xor U20147 (N_20147,N_18623,N_18550);
nor U20148 (N_20148,N_18475,N_18362);
and U20149 (N_20149,N_18392,N_18011);
nand U20150 (N_20150,N_18836,N_18676);
nand U20151 (N_20151,N_18597,N_18792);
or U20152 (N_20152,N_18832,N_18233);
nor U20153 (N_20153,N_18102,N_18844);
nand U20154 (N_20154,N_19044,N_18974);
xor U20155 (N_20155,N_18875,N_18334);
and U20156 (N_20156,N_18419,N_19030);
xnor U20157 (N_20157,N_18554,N_18457);
and U20158 (N_20158,N_18263,N_18247);
or U20159 (N_20159,N_18665,N_18333);
nand U20160 (N_20160,N_18493,N_18749);
nand U20161 (N_20161,N_18567,N_18511);
and U20162 (N_20162,N_18438,N_18158);
and U20163 (N_20163,N_18628,N_18961);
xor U20164 (N_20164,N_18656,N_18829);
or U20165 (N_20165,N_18933,N_18372);
nand U20166 (N_20166,N_18193,N_18823);
nor U20167 (N_20167,N_18757,N_18862);
xnor U20168 (N_20168,N_18976,N_18219);
and U20169 (N_20169,N_18785,N_18679);
nor U20170 (N_20170,N_19090,N_18038);
or U20171 (N_20171,N_18624,N_18265);
xor U20172 (N_20172,N_18960,N_18760);
xor U20173 (N_20173,N_18827,N_18001);
nand U20174 (N_20174,N_18294,N_18350);
nor U20175 (N_20175,N_18527,N_18868);
or U20176 (N_20176,N_18351,N_18142);
nor U20177 (N_20177,N_19185,N_18243);
nor U20178 (N_20178,N_18644,N_18632);
xor U20179 (N_20179,N_18607,N_18305);
nor U20180 (N_20180,N_18608,N_19033);
nor U20181 (N_20181,N_18138,N_18640);
or U20182 (N_20182,N_18893,N_18619);
xnor U20183 (N_20183,N_18350,N_18663);
or U20184 (N_20184,N_18577,N_18997);
xnor U20185 (N_20185,N_18052,N_18739);
nand U20186 (N_20186,N_18462,N_18983);
nor U20187 (N_20187,N_18048,N_19182);
nand U20188 (N_20188,N_18208,N_18910);
nor U20189 (N_20189,N_18270,N_18681);
nand U20190 (N_20190,N_18980,N_18307);
or U20191 (N_20191,N_18649,N_18291);
nor U20192 (N_20192,N_18818,N_18235);
nand U20193 (N_20193,N_18922,N_18224);
xor U20194 (N_20194,N_18962,N_19142);
or U20195 (N_20195,N_18043,N_18227);
nand U20196 (N_20196,N_19007,N_18213);
or U20197 (N_20197,N_18112,N_18456);
nor U20198 (N_20198,N_18110,N_18569);
nor U20199 (N_20199,N_18043,N_18957);
nor U20200 (N_20200,N_18787,N_18664);
and U20201 (N_20201,N_18333,N_18144);
xnor U20202 (N_20202,N_18144,N_18415);
xnor U20203 (N_20203,N_18292,N_18515);
and U20204 (N_20204,N_18560,N_18641);
xnor U20205 (N_20205,N_18714,N_18609);
xor U20206 (N_20206,N_18850,N_18241);
and U20207 (N_20207,N_18637,N_18419);
xnor U20208 (N_20208,N_18681,N_18241);
nor U20209 (N_20209,N_18907,N_19197);
and U20210 (N_20210,N_18313,N_18490);
and U20211 (N_20211,N_18726,N_18254);
and U20212 (N_20212,N_18213,N_18558);
nand U20213 (N_20213,N_18324,N_18382);
or U20214 (N_20214,N_18133,N_18019);
nand U20215 (N_20215,N_19107,N_18022);
xnor U20216 (N_20216,N_18747,N_18973);
nand U20217 (N_20217,N_18014,N_18768);
or U20218 (N_20218,N_18917,N_18924);
nand U20219 (N_20219,N_19005,N_18409);
nor U20220 (N_20220,N_18375,N_18852);
and U20221 (N_20221,N_18032,N_18171);
nor U20222 (N_20222,N_19073,N_19125);
or U20223 (N_20223,N_18483,N_18666);
nand U20224 (N_20224,N_18251,N_18844);
xor U20225 (N_20225,N_18726,N_19088);
and U20226 (N_20226,N_18335,N_18763);
nor U20227 (N_20227,N_18330,N_18834);
xnor U20228 (N_20228,N_18285,N_18796);
nor U20229 (N_20229,N_18312,N_18695);
nor U20230 (N_20230,N_18593,N_18586);
nand U20231 (N_20231,N_19139,N_18298);
nor U20232 (N_20232,N_18066,N_19063);
xnor U20233 (N_20233,N_18794,N_18790);
nor U20234 (N_20234,N_19069,N_18052);
xor U20235 (N_20235,N_18396,N_19189);
or U20236 (N_20236,N_18229,N_18231);
nor U20237 (N_20237,N_18291,N_19038);
nor U20238 (N_20238,N_18856,N_18398);
or U20239 (N_20239,N_18318,N_18429);
xnor U20240 (N_20240,N_18892,N_18139);
nand U20241 (N_20241,N_18438,N_18181);
xor U20242 (N_20242,N_18473,N_18235);
and U20243 (N_20243,N_18116,N_19034);
and U20244 (N_20244,N_19198,N_18810);
xor U20245 (N_20245,N_18583,N_18401);
or U20246 (N_20246,N_18054,N_18491);
and U20247 (N_20247,N_18302,N_18175);
and U20248 (N_20248,N_18214,N_18516);
nor U20249 (N_20249,N_18614,N_18743);
or U20250 (N_20250,N_18232,N_18761);
xnor U20251 (N_20251,N_18574,N_18851);
xor U20252 (N_20252,N_18282,N_18839);
nand U20253 (N_20253,N_18965,N_18560);
nor U20254 (N_20254,N_18584,N_18686);
or U20255 (N_20255,N_19134,N_18738);
nand U20256 (N_20256,N_18032,N_18414);
xor U20257 (N_20257,N_18009,N_18464);
xnor U20258 (N_20258,N_18895,N_18909);
nor U20259 (N_20259,N_18305,N_18738);
nor U20260 (N_20260,N_18013,N_18573);
xor U20261 (N_20261,N_18986,N_18278);
xor U20262 (N_20262,N_18694,N_19179);
xor U20263 (N_20263,N_18091,N_19194);
or U20264 (N_20264,N_18666,N_18237);
nor U20265 (N_20265,N_18428,N_18047);
xor U20266 (N_20266,N_18730,N_18296);
or U20267 (N_20267,N_18798,N_18804);
nor U20268 (N_20268,N_18022,N_18824);
xnor U20269 (N_20269,N_18587,N_19009);
nand U20270 (N_20270,N_18899,N_18396);
or U20271 (N_20271,N_18072,N_18978);
and U20272 (N_20272,N_18388,N_19150);
nor U20273 (N_20273,N_18572,N_18141);
xor U20274 (N_20274,N_18646,N_18693);
nand U20275 (N_20275,N_18571,N_18328);
and U20276 (N_20276,N_18285,N_18928);
and U20277 (N_20277,N_18413,N_18925);
or U20278 (N_20278,N_18395,N_18939);
or U20279 (N_20279,N_18235,N_18862);
or U20280 (N_20280,N_18507,N_19022);
and U20281 (N_20281,N_18236,N_18147);
nor U20282 (N_20282,N_18254,N_18771);
xnor U20283 (N_20283,N_18208,N_18515);
and U20284 (N_20284,N_18614,N_18144);
or U20285 (N_20285,N_19045,N_18904);
nand U20286 (N_20286,N_18024,N_18456);
nand U20287 (N_20287,N_18882,N_18552);
nand U20288 (N_20288,N_19004,N_18726);
or U20289 (N_20289,N_18510,N_18577);
xor U20290 (N_20290,N_18252,N_18259);
nand U20291 (N_20291,N_18550,N_19038);
or U20292 (N_20292,N_19018,N_18548);
nand U20293 (N_20293,N_19108,N_18220);
or U20294 (N_20294,N_18916,N_18712);
and U20295 (N_20295,N_18776,N_18877);
nand U20296 (N_20296,N_18311,N_18462);
or U20297 (N_20297,N_18425,N_18904);
nor U20298 (N_20298,N_18783,N_18632);
nor U20299 (N_20299,N_18669,N_18828);
nand U20300 (N_20300,N_18333,N_18575);
xor U20301 (N_20301,N_18828,N_18100);
nor U20302 (N_20302,N_18719,N_18938);
nor U20303 (N_20303,N_18583,N_19172);
and U20304 (N_20304,N_18072,N_18105);
xnor U20305 (N_20305,N_18143,N_19124);
xor U20306 (N_20306,N_18684,N_18708);
xor U20307 (N_20307,N_18836,N_18960);
or U20308 (N_20308,N_19008,N_18566);
and U20309 (N_20309,N_18396,N_18217);
and U20310 (N_20310,N_19078,N_18669);
and U20311 (N_20311,N_18991,N_18382);
or U20312 (N_20312,N_19132,N_18367);
xnor U20313 (N_20313,N_18679,N_18255);
or U20314 (N_20314,N_18357,N_18598);
nand U20315 (N_20315,N_18072,N_18409);
nor U20316 (N_20316,N_18825,N_18621);
xor U20317 (N_20317,N_18916,N_18787);
or U20318 (N_20318,N_18025,N_18283);
nand U20319 (N_20319,N_18434,N_18325);
nor U20320 (N_20320,N_18817,N_18991);
nor U20321 (N_20321,N_18534,N_18464);
nor U20322 (N_20322,N_19000,N_18713);
xor U20323 (N_20323,N_18256,N_18425);
or U20324 (N_20324,N_19093,N_19197);
and U20325 (N_20325,N_18863,N_18054);
or U20326 (N_20326,N_19196,N_18111);
xnor U20327 (N_20327,N_18865,N_18177);
xor U20328 (N_20328,N_18012,N_18695);
nor U20329 (N_20329,N_18896,N_18322);
nor U20330 (N_20330,N_18735,N_18981);
or U20331 (N_20331,N_18671,N_18763);
nor U20332 (N_20332,N_18638,N_19143);
nand U20333 (N_20333,N_18633,N_18613);
nand U20334 (N_20334,N_18255,N_18369);
or U20335 (N_20335,N_18025,N_18695);
xor U20336 (N_20336,N_18991,N_18702);
nand U20337 (N_20337,N_18232,N_18310);
nor U20338 (N_20338,N_18759,N_18044);
and U20339 (N_20339,N_19036,N_18453);
xnor U20340 (N_20340,N_18549,N_18365);
and U20341 (N_20341,N_19133,N_18514);
xor U20342 (N_20342,N_19034,N_18392);
nor U20343 (N_20343,N_18793,N_18465);
and U20344 (N_20344,N_18958,N_18503);
nor U20345 (N_20345,N_18844,N_18694);
xor U20346 (N_20346,N_18834,N_18649);
or U20347 (N_20347,N_18226,N_18702);
or U20348 (N_20348,N_18282,N_18235);
xor U20349 (N_20349,N_18961,N_18682);
or U20350 (N_20350,N_19054,N_18640);
nor U20351 (N_20351,N_18528,N_18075);
nor U20352 (N_20352,N_19149,N_18284);
nand U20353 (N_20353,N_18222,N_19088);
nand U20354 (N_20354,N_18809,N_18317);
nand U20355 (N_20355,N_18858,N_18948);
or U20356 (N_20356,N_18789,N_18040);
nand U20357 (N_20357,N_18686,N_18638);
nand U20358 (N_20358,N_18185,N_18350);
xor U20359 (N_20359,N_18098,N_18682);
nor U20360 (N_20360,N_19060,N_18927);
nand U20361 (N_20361,N_18501,N_18183);
nand U20362 (N_20362,N_18843,N_19034);
nor U20363 (N_20363,N_18710,N_18086);
and U20364 (N_20364,N_18076,N_18288);
nand U20365 (N_20365,N_19154,N_18362);
nand U20366 (N_20366,N_18610,N_18848);
nand U20367 (N_20367,N_18367,N_18917);
xnor U20368 (N_20368,N_18773,N_18104);
nand U20369 (N_20369,N_18698,N_18405);
nand U20370 (N_20370,N_18278,N_18228);
xor U20371 (N_20371,N_18535,N_19050);
nor U20372 (N_20372,N_18212,N_18852);
and U20373 (N_20373,N_18079,N_18371);
and U20374 (N_20374,N_18431,N_18367);
or U20375 (N_20375,N_18938,N_18404);
nor U20376 (N_20376,N_18842,N_18529);
nand U20377 (N_20377,N_18264,N_19031);
xor U20378 (N_20378,N_18029,N_19050);
xor U20379 (N_20379,N_18120,N_18541);
xnor U20380 (N_20380,N_18915,N_18250);
nand U20381 (N_20381,N_19057,N_18389);
nor U20382 (N_20382,N_18391,N_18037);
or U20383 (N_20383,N_18673,N_18397);
nand U20384 (N_20384,N_18460,N_18129);
nand U20385 (N_20385,N_18702,N_18321);
xnor U20386 (N_20386,N_18637,N_18214);
or U20387 (N_20387,N_18423,N_18522);
nand U20388 (N_20388,N_19106,N_18775);
nand U20389 (N_20389,N_18890,N_18078);
nand U20390 (N_20390,N_18516,N_18825);
nand U20391 (N_20391,N_18846,N_19129);
xor U20392 (N_20392,N_18373,N_18096);
nor U20393 (N_20393,N_18832,N_18335);
or U20394 (N_20394,N_18793,N_18705);
nor U20395 (N_20395,N_19137,N_18619);
or U20396 (N_20396,N_18163,N_18248);
and U20397 (N_20397,N_19032,N_18288);
xnor U20398 (N_20398,N_18047,N_19105);
nor U20399 (N_20399,N_18425,N_18795);
or U20400 (N_20400,N_20018,N_20289);
nor U20401 (N_20401,N_19513,N_20262);
and U20402 (N_20402,N_19876,N_19431);
or U20403 (N_20403,N_20146,N_20391);
or U20404 (N_20404,N_19656,N_20252);
nor U20405 (N_20405,N_19556,N_20304);
nand U20406 (N_20406,N_19887,N_20075);
xnor U20407 (N_20407,N_19456,N_19952);
xor U20408 (N_20408,N_19633,N_20055);
nor U20409 (N_20409,N_19848,N_19672);
xor U20410 (N_20410,N_19951,N_19226);
xor U20411 (N_20411,N_19457,N_19806);
xor U20412 (N_20412,N_20179,N_20191);
and U20413 (N_20413,N_19590,N_19916);
nand U20414 (N_20414,N_20136,N_19717);
nand U20415 (N_20415,N_19896,N_20182);
xnor U20416 (N_20416,N_20323,N_20361);
nor U20417 (N_20417,N_19734,N_19446);
or U20418 (N_20418,N_20142,N_20219);
xor U20419 (N_20419,N_19266,N_19616);
nor U20420 (N_20420,N_19253,N_19571);
or U20421 (N_20421,N_19627,N_19336);
xnor U20422 (N_20422,N_19724,N_20054);
nor U20423 (N_20423,N_20270,N_20329);
and U20424 (N_20424,N_20254,N_20026);
xnor U20425 (N_20425,N_20390,N_20045);
nor U20426 (N_20426,N_19641,N_19706);
xor U20427 (N_20427,N_19488,N_19567);
xor U20428 (N_20428,N_20202,N_20171);
or U20429 (N_20429,N_20206,N_19500);
or U20430 (N_20430,N_19964,N_19747);
or U20431 (N_20431,N_19966,N_19882);
xor U20432 (N_20432,N_20068,N_19606);
or U20433 (N_20433,N_19455,N_19692);
or U20434 (N_20434,N_19603,N_20084);
nand U20435 (N_20435,N_20071,N_20389);
xnor U20436 (N_20436,N_19762,N_19698);
nand U20437 (N_20437,N_20152,N_19503);
nor U20438 (N_20438,N_20003,N_20034);
and U20439 (N_20439,N_20192,N_19945);
xnor U20440 (N_20440,N_19342,N_19995);
nor U20441 (N_20441,N_19785,N_20150);
nand U20442 (N_20442,N_19751,N_19398);
nor U20443 (N_20443,N_20324,N_19524);
xnor U20444 (N_20444,N_19244,N_19662);
nor U20445 (N_20445,N_20024,N_19671);
or U20446 (N_20446,N_19652,N_20157);
xor U20447 (N_20447,N_19333,N_20215);
nor U20448 (N_20448,N_19517,N_20271);
nor U20449 (N_20449,N_19468,N_19424);
nand U20450 (N_20450,N_19721,N_20246);
nand U20451 (N_20451,N_20067,N_19290);
nor U20452 (N_20452,N_19303,N_20053);
xor U20453 (N_20453,N_19328,N_19486);
nor U20454 (N_20454,N_20010,N_19286);
or U20455 (N_20455,N_20355,N_19217);
xor U20456 (N_20456,N_20030,N_19708);
nor U20457 (N_20457,N_19388,N_19920);
and U20458 (N_20458,N_20303,N_20106);
nand U20459 (N_20459,N_19994,N_19930);
or U20460 (N_20460,N_19400,N_19579);
nor U20461 (N_20461,N_19230,N_19666);
or U20462 (N_20462,N_19310,N_19414);
or U20463 (N_20463,N_20322,N_19643);
and U20464 (N_20464,N_20226,N_19704);
nor U20465 (N_20465,N_20048,N_19906);
nand U20466 (N_20466,N_19324,N_19454);
nand U20467 (N_20467,N_19955,N_19469);
xnor U20468 (N_20468,N_19772,N_19279);
and U20469 (N_20469,N_19776,N_19915);
and U20470 (N_20470,N_20032,N_19857);
nand U20471 (N_20471,N_19593,N_20284);
xor U20472 (N_20472,N_19936,N_19238);
and U20473 (N_20473,N_20058,N_19396);
nor U20474 (N_20474,N_20041,N_20300);
nand U20475 (N_20475,N_20044,N_19228);
and U20476 (N_20476,N_20096,N_20392);
nor U20477 (N_20477,N_20049,N_20004);
or U20478 (N_20478,N_19349,N_20159);
and U20479 (N_20479,N_19584,N_19744);
nand U20480 (N_20480,N_20187,N_19630);
and U20481 (N_20481,N_20188,N_20031);
or U20482 (N_20482,N_19550,N_20332);
xor U20483 (N_20483,N_20119,N_19783);
xor U20484 (N_20484,N_20275,N_19453);
nand U20485 (N_20485,N_19561,N_19805);
nand U20486 (N_20486,N_19629,N_19812);
and U20487 (N_20487,N_19752,N_19540);
and U20488 (N_20488,N_19673,N_19620);
or U20489 (N_20489,N_19216,N_20156);
xor U20490 (N_20490,N_20094,N_19528);
nor U20491 (N_20491,N_19270,N_19642);
and U20492 (N_20492,N_19760,N_19221);
nor U20493 (N_20493,N_19723,N_19660);
nand U20494 (N_20494,N_20394,N_19322);
xnor U20495 (N_20495,N_20302,N_19944);
xor U20496 (N_20496,N_19251,N_19663);
or U20497 (N_20497,N_20015,N_19722);
xor U20498 (N_20498,N_19378,N_19525);
nor U20499 (N_20499,N_19299,N_19465);
nor U20500 (N_20500,N_19413,N_19733);
nor U20501 (N_20501,N_19379,N_19852);
and U20502 (N_20502,N_20116,N_20241);
xor U20503 (N_20503,N_19731,N_19757);
nor U20504 (N_20504,N_19859,N_20100);
xor U20505 (N_20505,N_19452,N_19683);
nor U20506 (N_20506,N_19821,N_19509);
nor U20507 (N_20507,N_20133,N_19958);
nor U20508 (N_20508,N_19542,N_19773);
or U20509 (N_20509,N_20016,N_19287);
xor U20510 (N_20510,N_19613,N_20261);
and U20511 (N_20511,N_19931,N_19505);
nand U20512 (N_20512,N_19204,N_19661);
or U20513 (N_20513,N_20231,N_20283);
xnor U20514 (N_20514,N_19645,N_20139);
xor U20515 (N_20515,N_19419,N_19547);
nor U20516 (N_20516,N_19397,N_19969);
xnor U20517 (N_20517,N_20278,N_19913);
and U20518 (N_20518,N_20087,N_19485);
or U20519 (N_20519,N_20288,N_20277);
or U20520 (N_20520,N_19720,N_20359);
nand U20521 (N_20521,N_19972,N_20085);
or U20522 (N_20522,N_20124,N_19269);
nor U20523 (N_20523,N_20164,N_20235);
and U20524 (N_20524,N_19529,N_20110);
nor U20525 (N_20525,N_19306,N_20245);
nor U20526 (N_20526,N_19255,N_20145);
and U20527 (N_20527,N_20258,N_19715);
xnor U20528 (N_20528,N_19311,N_20073);
and U20529 (N_20529,N_20033,N_19410);
xor U20530 (N_20530,N_20040,N_20293);
and U20531 (N_20531,N_20263,N_19712);
nand U20532 (N_20532,N_19993,N_19364);
nor U20533 (N_20533,N_19243,N_19830);
and U20534 (N_20534,N_20372,N_20396);
xor U20535 (N_20535,N_20321,N_19834);
and U20536 (N_20536,N_19713,N_20209);
and U20537 (N_20537,N_19209,N_20169);
and U20538 (N_20538,N_19921,N_19572);
and U20539 (N_20539,N_19978,N_20057);
nand U20540 (N_20540,N_19585,N_19832);
nor U20541 (N_20541,N_19441,N_19604);
xnor U20542 (N_20542,N_19438,N_19746);
nor U20543 (N_20543,N_19638,N_20196);
or U20544 (N_20544,N_19440,N_19450);
or U20545 (N_20545,N_19300,N_19654);
xor U20546 (N_20546,N_20186,N_20248);
nand U20547 (N_20547,N_20217,N_19335);
xor U20548 (N_20548,N_19412,N_19735);
nand U20549 (N_20549,N_20028,N_19977);
and U20550 (N_20550,N_19777,N_19515);
xor U20551 (N_20551,N_19828,N_20341);
nor U20552 (N_20552,N_20297,N_19825);
nand U20553 (N_20553,N_19695,N_20266);
nand U20554 (N_20554,N_20222,N_19502);
or U20555 (N_20555,N_20077,N_19280);
nor U20556 (N_20556,N_20240,N_20279);
nor U20557 (N_20557,N_19658,N_19459);
nor U20558 (N_20558,N_19754,N_19587);
nand U20559 (N_20559,N_20051,N_20078);
xor U20560 (N_20560,N_19693,N_19490);
or U20561 (N_20561,N_19974,N_19808);
and U20562 (N_20562,N_19399,N_20346);
and U20563 (N_20563,N_19853,N_20313);
xor U20564 (N_20564,N_20162,N_19527);
nand U20565 (N_20565,N_19792,N_19725);
nand U20566 (N_20566,N_19258,N_20287);
and U20567 (N_20567,N_20072,N_19753);
and U20568 (N_20568,N_20325,N_19867);
nand U20569 (N_20569,N_19375,N_19614);
nand U20570 (N_20570,N_20035,N_19729);
or U20571 (N_20571,N_19790,N_19317);
nor U20572 (N_20572,N_20063,N_20330);
xnor U20573 (N_20573,N_19665,N_20269);
or U20574 (N_20574,N_20371,N_20345);
nor U20575 (N_20575,N_19411,N_19223);
nor U20576 (N_20576,N_20229,N_19910);
and U20577 (N_20577,N_20267,N_20099);
xor U20578 (N_20578,N_19981,N_19617);
or U20579 (N_20579,N_19248,N_19205);
nand U20580 (N_20580,N_19384,N_20397);
nand U20581 (N_20581,N_20247,N_19471);
nand U20582 (N_20582,N_20308,N_20023);
nand U20583 (N_20583,N_19222,N_19766);
xnor U20584 (N_20584,N_20036,N_19855);
nand U20585 (N_20585,N_19254,N_19647);
nor U20586 (N_20586,N_19596,N_19710);
and U20587 (N_20587,N_20008,N_19489);
nand U20588 (N_20588,N_20286,N_20234);
nor U20589 (N_20589,N_19391,N_19730);
xnor U20590 (N_20590,N_19566,N_19674);
or U20591 (N_20591,N_20006,N_20128);
xnor U20592 (N_20592,N_20014,N_19664);
or U20593 (N_20593,N_19940,N_20369);
nor U20594 (N_20594,N_19366,N_19804);
and U20595 (N_20595,N_20377,N_19680);
and U20596 (N_20596,N_20333,N_19236);
and U20597 (N_20597,N_19403,N_20052);
or U20598 (N_20598,N_19798,N_19481);
or U20599 (N_20599,N_19321,N_19780);
or U20600 (N_20600,N_20172,N_19743);
nor U20601 (N_20601,N_20280,N_19592);
xor U20602 (N_20602,N_19367,N_19778);
or U20603 (N_20603,N_19959,N_19562);
nor U20604 (N_20604,N_19430,N_20292);
nor U20605 (N_20605,N_20260,N_19339);
xor U20606 (N_20606,N_20257,N_20348);
nand U20607 (N_20607,N_19771,N_20367);
nand U20608 (N_20608,N_19554,N_20340);
nand U20609 (N_20609,N_20233,N_19582);
and U20610 (N_20610,N_20081,N_19467);
and U20611 (N_20611,N_19491,N_20170);
and U20612 (N_20612,N_20114,N_19395);
nand U20613 (N_20613,N_20368,N_20273);
xnor U20614 (N_20614,N_20294,N_20011);
or U20615 (N_20615,N_19738,N_20317);
nand U20616 (N_20616,N_19626,N_19847);
and U20617 (N_20617,N_19711,N_19507);
and U20618 (N_20618,N_19894,N_19901);
and U20619 (N_20619,N_19983,N_20210);
xnor U20620 (N_20620,N_20344,N_19681);
nand U20621 (N_20621,N_19911,N_19763);
xor U20622 (N_20622,N_20259,N_20125);
nor U20623 (N_20623,N_20319,N_20005);
xnor U20624 (N_20624,N_19595,N_19605);
or U20625 (N_20625,N_20109,N_20020);
xnor U20626 (N_20626,N_19831,N_20002);
nand U20627 (N_20627,N_19929,N_19536);
nand U20628 (N_20628,N_20199,N_20098);
xor U20629 (N_20629,N_19329,N_20339);
and U20630 (N_20630,N_20122,N_20358);
nor U20631 (N_20631,N_19922,N_19492);
and U20632 (N_20632,N_19219,N_19493);
nor U20633 (N_20633,N_19741,N_20129);
nand U20634 (N_20634,N_19954,N_20314);
nand U20635 (N_20635,N_20176,N_19863);
nor U20636 (N_20636,N_19420,N_19967);
or U20637 (N_20637,N_19416,N_19272);
xor U20638 (N_20638,N_19843,N_19569);
nand U20639 (N_20639,N_19979,N_19241);
or U20640 (N_20640,N_19239,N_19568);
nor U20641 (N_20641,N_19546,N_20197);
and U20642 (N_20642,N_20238,N_19774);
nand U20643 (N_20643,N_20046,N_20029);
nor U20644 (N_20644,N_20301,N_19232);
or U20645 (N_20645,N_19631,N_20079);
nand U20646 (N_20646,N_19314,N_20091);
nand U20647 (N_20647,N_19235,N_20165);
nor U20648 (N_20648,N_20306,N_19866);
xor U20649 (N_20649,N_19268,N_19895);
xnor U20650 (N_20650,N_19632,N_20112);
or U20651 (N_20651,N_20151,N_20126);
or U20652 (N_20652,N_19758,N_19991);
nand U20653 (N_20653,N_19845,N_19976);
nor U20654 (N_20654,N_20264,N_20092);
or U20655 (N_20655,N_19823,N_19942);
or U20656 (N_20656,N_19618,N_20174);
and U20657 (N_20657,N_19284,N_20309);
nand U20658 (N_20658,N_19338,N_20177);
nor U20659 (N_20659,N_19407,N_19415);
nor U20660 (N_20660,N_19427,N_19496);
xor U20661 (N_20661,N_19480,N_19477);
and U20662 (N_20662,N_19639,N_20042);
nor U20663 (N_20663,N_20378,N_20117);
nor U20664 (N_20664,N_20356,N_19353);
nand U20665 (N_20665,N_20000,N_19227);
nor U20666 (N_20666,N_19833,N_19409);
and U20667 (N_20667,N_19215,N_19343);
nor U20668 (N_20668,N_19689,N_19787);
and U20669 (N_20669,N_19878,N_19923);
and U20670 (N_20670,N_19522,N_19233);
nand U20671 (N_20671,N_20250,N_20127);
xnor U20672 (N_20672,N_19946,N_19668);
and U20673 (N_20673,N_19312,N_20061);
xnor U20674 (N_20674,N_20120,N_19838);
nand U20675 (N_20675,N_19225,N_20244);
nand U20676 (N_20676,N_19634,N_19950);
nand U20677 (N_20677,N_19301,N_19611);
and U20678 (N_20678,N_20101,N_19948);
nand U20679 (N_20679,N_19460,N_19851);
nor U20680 (N_20680,N_19897,N_19849);
nor U20681 (N_20681,N_19218,N_19256);
or U20682 (N_20682,N_20102,N_20331);
xor U20683 (N_20683,N_19799,N_19334);
and U20684 (N_20684,N_19612,N_20070);
and U20685 (N_20685,N_19240,N_19332);
nor U20686 (N_20686,N_20195,N_19581);
nand U20687 (N_20687,N_20347,N_20086);
or U20688 (N_20688,N_20316,N_19369);
nor U20689 (N_20689,N_19576,N_19383);
or U20690 (N_20690,N_19552,N_19348);
or U20691 (N_20691,N_19594,N_20059);
nand U20692 (N_20692,N_19992,N_19516);
or U20693 (N_20693,N_20335,N_19201);
or U20694 (N_20694,N_19323,N_19809);
and U20695 (N_20695,N_20296,N_19802);
nand U20696 (N_20696,N_20069,N_19473);
nor U20697 (N_20697,N_20350,N_19406);
xor U20698 (N_20698,N_19653,N_19390);
and U20699 (N_20699,N_19274,N_19675);
or U20700 (N_20700,N_20123,N_19260);
nand U20701 (N_20701,N_19417,N_19909);
nor U20702 (N_20702,N_19305,N_20342);
and U20703 (N_20703,N_19534,N_19445);
xnor U20704 (N_20704,N_19800,N_19242);
or U20705 (N_20705,N_19482,N_20365);
xor U20706 (N_20706,N_20290,N_20388);
and U20707 (N_20707,N_19423,N_19444);
nor U20708 (N_20708,N_20386,N_19988);
or U20709 (N_20709,N_19702,N_19302);
or U20710 (N_20710,N_19869,N_19868);
xor U20711 (N_20711,N_19487,N_19330);
nand U20712 (N_20712,N_19293,N_20095);
nand U20713 (N_20713,N_19376,N_19877);
and U20714 (N_20714,N_19926,N_20281);
nand U20715 (N_20715,N_19908,N_19862);
and U20716 (N_20716,N_19498,N_20009);
xor U20717 (N_20717,N_19354,N_19608);
nand U20718 (N_20718,N_20088,N_20194);
nand U20719 (N_20719,N_19893,N_20236);
or U20720 (N_20720,N_20375,N_19749);
or U20721 (N_20721,N_20334,N_19275);
and U20722 (N_20722,N_20097,N_19697);
and U20723 (N_20723,N_19237,N_19356);
xor U20724 (N_20724,N_19404,N_19841);
or U20725 (N_20725,N_19928,N_20083);
nor U20726 (N_20726,N_19484,N_20065);
and U20727 (N_20727,N_19870,N_19434);
nand U20728 (N_20728,N_20398,N_19659);
and U20729 (N_20729,N_20149,N_19361);
xnor U20730 (N_20730,N_19598,N_19351);
nor U20731 (N_20731,N_19933,N_20181);
nor U20732 (N_20732,N_19532,N_19728);
and U20733 (N_20733,N_19797,N_19288);
nand U20734 (N_20734,N_20265,N_19291);
and U20735 (N_20735,N_19984,N_19707);
or U20736 (N_20736,N_19884,N_19602);
nand U20737 (N_20737,N_20351,N_19919);
nand U20738 (N_20738,N_19885,N_19347);
nor U20739 (N_20739,N_19943,N_19432);
nand U20740 (N_20740,N_20017,N_19801);
or U20741 (N_20741,N_19925,N_19970);
xor U20742 (N_20742,N_20295,N_19835);
nand U20743 (N_20743,N_20221,N_19640);
and U20744 (N_20744,N_20320,N_19912);
and U20745 (N_20745,N_19837,N_19858);
nand U20746 (N_20746,N_19827,N_19705);
and U20747 (N_20747,N_19313,N_19553);
or U20748 (N_20748,N_19883,N_19817);
nor U20749 (N_20749,N_20216,N_19686);
and U20750 (N_20750,N_20074,N_19245);
and U20751 (N_20751,N_19402,N_20242);
or U20752 (N_20752,N_20107,N_19900);
nor U20753 (N_20753,N_19971,N_19861);
nor U20754 (N_20754,N_20366,N_19401);
or U20755 (N_20755,N_20349,N_19565);
and U20756 (N_20756,N_19296,N_20056);
and U20757 (N_20757,N_20019,N_20189);
nand U20758 (N_20758,N_19325,N_19985);
xnor U20759 (N_20759,N_19212,N_20311);
nor U20760 (N_20760,N_19609,N_19259);
xnor U20761 (N_20761,N_20025,N_20363);
nor U20762 (N_20762,N_19842,N_20080);
xnor U20763 (N_20763,N_19531,N_19365);
and U20764 (N_20764,N_20012,N_19651);
nor U20765 (N_20765,N_19815,N_20062);
nand U20766 (N_20766,N_20132,N_19650);
or U20767 (N_20767,N_19784,N_20038);
xnor U20768 (N_20768,N_20249,N_20180);
and U20769 (N_20769,N_20379,N_19386);
nor U20770 (N_20770,N_19224,N_19472);
or U20771 (N_20771,N_19782,N_19331);
or U20772 (N_20772,N_19263,N_19879);
nand U20773 (N_20773,N_19501,N_19850);
and U20774 (N_20774,N_19736,N_19687);
xor U20775 (N_20775,N_19676,N_19580);
nor U20776 (N_20776,N_19856,N_19368);
and U20777 (N_20777,N_19474,N_19816);
and U20778 (N_20778,N_19319,N_19914);
nand U20779 (N_20779,N_20001,N_19429);
or U20780 (N_20780,N_20239,N_19458);
or U20781 (N_20781,N_19437,N_20208);
nor U20782 (N_20782,N_19341,N_19678);
or U20783 (N_20783,N_19699,N_19257);
nor U20784 (N_20784,N_20364,N_19839);
nand U20785 (N_20785,N_20135,N_20113);
or U20786 (N_20786,N_19803,N_19271);
nor U20787 (N_20787,N_20305,N_19548);
nor U20788 (N_20788,N_19588,N_19352);
and U20789 (N_20789,N_19476,N_19961);
and U20790 (N_20790,N_20227,N_19514);
and U20791 (N_20791,N_19574,N_20118);
nand U20792 (N_20792,N_19479,N_19518);
nor U20793 (N_20793,N_20343,N_20121);
xnor U20794 (N_20794,N_20066,N_19889);
and U20795 (N_20795,N_19359,N_19449);
and U20796 (N_20796,N_19756,N_19563);
nand U20797 (N_20797,N_19504,N_19670);
nor U20798 (N_20798,N_19577,N_19220);
nand U20799 (N_20799,N_20357,N_19965);
and U20800 (N_20800,N_19211,N_19541);
nor U20801 (N_20801,N_20220,N_19903);
or U20802 (N_20802,N_20022,N_19628);
or U20803 (N_20803,N_19982,N_20093);
nor U20804 (N_20804,N_20212,N_19511);
or U20805 (N_20805,N_19559,N_19295);
or U20806 (N_20806,N_19905,N_20282);
or U20807 (N_20807,N_19573,N_19794);
xor U20808 (N_20808,N_19363,N_19558);
nand U20809 (N_20809,N_19874,N_20184);
nor U20810 (N_20810,N_20131,N_19506);
xor U20811 (N_20811,N_19973,N_19538);
nand U20812 (N_20812,N_19523,N_19382);
nand U20813 (N_20813,N_19648,N_20251);
nand U20814 (N_20814,N_19924,N_19261);
and U20815 (N_20815,N_19519,N_20173);
and U20816 (N_20816,N_19881,N_19826);
nor U20817 (N_20817,N_20076,N_19426);
and U20818 (N_20818,N_19764,N_19264);
nor U20819 (N_20819,N_19997,N_20168);
and U20820 (N_20820,N_20082,N_19583);
xnor U20821 (N_20821,N_19636,N_20362);
and U20822 (N_20822,N_19655,N_20115);
nor U20823 (N_20823,N_19769,N_19544);
and U20824 (N_20824,N_19937,N_19309);
xor U20825 (N_20825,N_19732,N_19880);
and U20826 (N_20826,N_19748,N_19273);
nand U20827 (N_20827,N_19907,N_19340);
nand U20828 (N_20828,N_19327,N_19987);
xor U20829 (N_20829,N_20272,N_19701);
xnor U20830 (N_20830,N_19557,N_20353);
and U20831 (N_20831,N_19840,N_20230);
xnor U20832 (N_20832,N_20013,N_20148);
or U20833 (N_20833,N_19962,N_20064);
nor U20834 (N_20834,N_19247,N_19387);
and U20835 (N_20835,N_19535,N_19370);
nor U20836 (N_20836,N_19750,N_19873);
nand U20837 (N_20837,N_20108,N_19865);
xor U20838 (N_20838,N_20089,N_19267);
or U20839 (N_20839,N_19439,N_20060);
nor U20840 (N_20840,N_19372,N_19373);
nor U20841 (N_20841,N_19854,N_19688);
nand U20842 (N_20842,N_19462,N_20318);
nor U20843 (N_20843,N_19591,N_19644);
and U20844 (N_20844,N_20143,N_20161);
nor U20845 (N_20845,N_20387,N_19278);
xor U20846 (N_20846,N_19408,N_19470);
nor U20847 (N_20847,N_19694,N_19307);
or U20848 (N_20848,N_19564,N_19326);
or U20849 (N_20849,N_19941,N_19345);
and U20850 (N_20850,N_19898,N_20370);
and U20851 (N_20851,N_19425,N_19872);
or U20852 (N_20852,N_20232,N_19765);
nand U20853 (N_20853,N_19207,N_19623);
nor U20854 (N_20854,N_20183,N_20207);
and U20855 (N_20855,N_20385,N_19234);
or U20856 (N_20856,N_20007,N_19788);
xor U20857 (N_20857,N_20198,N_19555);
or U20858 (N_20858,N_19599,N_19285);
nor U20859 (N_20859,N_19433,N_20352);
or U20860 (N_20860,N_19265,N_19545);
or U20861 (N_20861,N_19635,N_20047);
or U20862 (N_20862,N_20395,N_19814);
nand U20863 (N_20863,N_19451,N_19537);
or U20864 (N_20864,N_20228,N_19389);
and U20865 (N_20865,N_19813,N_20310);
and U20866 (N_20866,N_19520,N_20134);
and U20867 (N_20867,N_20163,N_19890);
nand U20868 (N_20868,N_19560,N_20328);
xor U20869 (N_20869,N_19727,N_19358);
and U20870 (N_20870,N_19975,N_19935);
nand U20871 (N_20871,N_20381,N_19461);
nor U20872 (N_20872,N_19394,N_19466);
nor U20873 (N_20873,N_19214,N_19298);
or U20874 (N_20874,N_19927,N_19277);
and U20875 (N_20875,N_20315,N_20382);
nor U20876 (N_20876,N_20336,N_19621);
nand U20877 (N_20877,N_19667,N_19996);
nor U20878 (N_20878,N_20383,N_19770);
nand U20879 (N_20879,N_19371,N_19475);
or U20880 (N_20880,N_19229,N_20050);
nand U20881 (N_20881,N_19337,N_19714);
nor U20882 (N_20882,N_20154,N_19289);
and U20883 (N_20883,N_19355,N_19478);
and U20884 (N_20884,N_19421,N_20155);
nand U20885 (N_20885,N_19779,N_19619);
xnor U20886 (N_20886,N_20255,N_20167);
nand U20887 (N_20887,N_19422,N_20160);
nand U20888 (N_20888,N_19249,N_20338);
and U20889 (N_20889,N_20312,N_19625);
nand U20890 (N_20890,N_19252,N_19202);
nand U20891 (N_20891,N_19691,N_19308);
and U20892 (N_20892,N_19939,N_20218);
and U20893 (N_20893,N_19539,N_19709);
or U20894 (N_20894,N_19957,N_19206);
nand U20895 (N_20895,N_20175,N_19622);
nand U20896 (N_20896,N_19807,N_20203);
xnor U20897 (N_20897,N_19350,N_19949);
nor U20898 (N_20898,N_19657,N_19677);
or U20899 (N_20899,N_19512,N_20268);
or U20900 (N_20900,N_19737,N_20021);
xor U20901 (N_20901,N_19637,N_19989);
and U20902 (N_20902,N_19294,N_20178);
and U20903 (N_20903,N_19447,N_19510);
and U20904 (N_20904,N_19904,N_19428);
or U20905 (N_20905,N_19947,N_20104);
xor U20906 (N_20906,N_19875,N_19768);
and U20907 (N_20907,N_19745,N_20037);
nand U20908 (N_20908,N_19963,N_19700);
nand U20909 (N_20909,N_19679,N_19418);
xnor U20910 (N_20910,N_20373,N_20224);
or U20911 (N_20911,N_19508,N_19682);
and U20912 (N_20912,N_19346,N_19597);
or U20913 (N_20913,N_19250,N_19917);
or U20914 (N_20914,N_19934,N_20130);
or U20915 (N_20915,N_19570,N_19886);
and U20916 (N_20916,N_19607,N_20299);
nand U20917 (N_20917,N_19615,N_19436);
and U20918 (N_20918,N_20326,N_19551);
xor U20919 (N_20919,N_19530,N_19385);
xor U20920 (N_20920,N_19980,N_19589);
nor U20921 (N_20921,N_19283,N_20166);
or U20922 (N_20922,N_19819,N_20360);
or U20923 (N_20923,N_19864,N_20185);
nor U20924 (N_20924,N_19786,N_19200);
and U20925 (N_20925,N_20298,N_20190);
and U20926 (N_20926,N_19740,N_19292);
and U20927 (N_20927,N_19393,N_19521);
nor U20928 (N_20928,N_19281,N_19775);
and U20929 (N_20929,N_19495,N_19276);
nor U20930 (N_20930,N_20201,N_20376);
nor U20931 (N_20931,N_19742,N_19795);
or U20932 (N_20932,N_19533,N_20043);
xor U20933 (N_20933,N_19381,N_19932);
xnor U20934 (N_20934,N_20354,N_19844);
or U20935 (N_20935,N_19836,N_20205);
xor U20936 (N_20936,N_20256,N_19231);
or U20937 (N_20937,N_19392,N_19820);
nand U20938 (N_20938,N_19318,N_20285);
xnor U20939 (N_20939,N_19448,N_19716);
xor U20940 (N_20940,N_19726,N_19210);
or U20941 (N_20941,N_19669,N_19953);
or U20942 (N_20942,N_20225,N_19986);
nand U20943 (N_20943,N_19781,N_20039);
or U20944 (N_20944,N_20204,N_19610);
or U20945 (N_20945,N_19968,N_19822);
nand U20946 (N_20946,N_19719,N_20393);
and U20947 (N_20947,N_19902,N_19767);
xor U20948 (N_20948,N_19601,N_19282);
nor U20949 (N_20949,N_19646,N_19297);
nand U20950 (N_20950,N_19499,N_19938);
or U20951 (N_20951,N_19549,N_19810);
xor U20952 (N_20952,N_20214,N_19600);
nand U20953 (N_20953,N_20237,N_19344);
nor U20954 (N_20954,N_19824,N_19320);
xnor U20955 (N_20955,N_19315,N_19755);
and U20956 (N_20956,N_19956,N_19871);
and U20957 (N_20957,N_19696,N_19442);
and U20958 (N_20958,N_20384,N_19435);
and U20959 (N_20959,N_20374,N_19860);
nor U20960 (N_20960,N_19960,N_19718);
or U20961 (N_20961,N_19796,N_19357);
xor U20962 (N_20962,N_19463,N_20213);
xnor U20963 (N_20963,N_19443,N_19526);
nor U20964 (N_20964,N_20253,N_19586);
or U20965 (N_20965,N_20337,N_20138);
xor U20966 (N_20966,N_19892,N_20103);
xor U20967 (N_20967,N_20200,N_19703);
xnor U20968 (N_20968,N_19793,N_20307);
or U20969 (N_20969,N_19759,N_19208);
xnor U20970 (N_20970,N_19203,N_19684);
nor U20971 (N_20971,N_19649,N_20223);
nor U20972 (N_20972,N_19829,N_19918);
nand U20973 (N_20973,N_19360,N_19899);
nand U20974 (N_20974,N_20291,N_20141);
xnor U20975 (N_20975,N_20380,N_19990);
nor U20976 (N_20976,N_19998,N_20193);
xnor U20977 (N_20977,N_19494,N_19213);
and U20978 (N_20978,N_20399,N_20105);
and U20979 (N_20979,N_19464,N_20243);
and U20980 (N_20980,N_20158,N_20276);
nor U20981 (N_20981,N_19789,N_19575);
or U20982 (N_20982,N_20090,N_19690);
xor U20983 (N_20983,N_19811,N_19791);
nand U20984 (N_20984,N_20140,N_19624);
nand U20985 (N_20985,N_20147,N_19761);
nand U20986 (N_20986,N_19685,N_19246);
or U20987 (N_20987,N_19483,N_19380);
and U20988 (N_20988,N_19739,N_19377);
xnor U20989 (N_20989,N_19578,N_20274);
and U20990 (N_20990,N_20327,N_19543);
or U20991 (N_20991,N_19362,N_19818);
xnor U20992 (N_20992,N_20211,N_19846);
and U20993 (N_20993,N_20153,N_19405);
and U20994 (N_20994,N_19888,N_20027);
nor U20995 (N_20995,N_19497,N_19999);
nor U20996 (N_20996,N_20137,N_19374);
nand U20997 (N_20997,N_20111,N_19316);
nand U20998 (N_20998,N_19304,N_19262);
nand U20999 (N_20999,N_19891,N_20144);
and U21000 (N_21000,N_19836,N_19818);
and U21001 (N_21001,N_20251,N_19986);
or U21002 (N_21002,N_20023,N_19575);
xor U21003 (N_21003,N_20284,N_20393);
xnor U21004 (N_21004,N_19605,N_19575);
or U21005 (N_21005,N_20038,N_20057);
xor U21006 (N_21006,N_19888,N_19450);
or U21007 (N_21007,N_19505,N_19644);
xor U21008 (N_21008,N_19342,N_19278);
and U21009 (N_21009,N_20146,N_19279);
or U21010 (N_21010,N_19471,N_19760);
nand U21011 (N_21011,N_19294,N_19634);
and U21012 (N_21012,N_19800,N_19816);
or U21013 (N_21013,N_19369,N_19925);
and U21014 (N_21014,N_19308,N_19795);
nand U21015 (N_21015,N_20332,N_19461);
nand U21016 (N_21016,N_19706,N_19386);
xnor U21017 (N_21017,N_20091,N_19734);
and U21018 (N_21018,N_19845,N_19400);
and U21019 (N_21019,N_19791,N_19511);
xnor U21020 (N_21020,N_20078,N_20219);
and U21021 (N_21021,N_20335,N_19639);
and U21022 (N_21022,N_19253,N_19629);
xor U21023 (N_21023,N_19965,N_20004);
nand U21024 (N_21024,N_20289,N_20209);
or U21025 (N_21025,N_19934,N_20232);
and U21026 (N_21026,N_19895,N_19380);
nand U21027 (N_21027,N_19374,N_20272);
nor U21028 (N_21028,N_20069,N_19596);
and U21029 (N_21029,N_19443,N_20035);
nand U21030 (N_21030,N_19644,N_19414);
or U21031 (N_21031,N_19207,N_19268);
nor U21032 (N_21032,N_19235,N_19610);
or U21033 (N_21033,N_20080,N_20192);
and U21034 (N_21034,N_20201,N_19454);
and U21035 (N_21035,N_19712,N_20189);
xnor U21036 (N_21036,N_19872,N_19245);
or U21037 (N_21037,N_19476,N_19956);
xnor U21038 (N_21038,N_19698,N_20370);
or U21039 (N_21039,N_20246,N_20010);
nor U21040 (N_21040,N_19616,N_19527);
nand U21041 (N_21041,N_19289,N_19715);
or U21042 (N_21042,N_19795,N_20091);
nor U21043 (N_21043,N_19796,N_19573);
or U21044 (N_21044,N_19681,N_19997);
and U21045 (N_21045,N_19651,N_19670);
xor U21046 (N_21046,N_20284,N_20008);
or U21047 (N_21047,N_20339,N_19208);
and U21048 (N_21048,N_19431,N_19808);
nand U21049 (N_21049,N_19674,N_19269);
or U21050 (N_21050,N_20135,N_20395);
xnor U21051 (N_21051,N_19667,N_19404);
nor U21052 (N_21052,N_20051,N_19289);
nand U21053 (N_21053,N_19642,N_19267);
nand U21054 (N_21054,N_20276,N_19384);
nor U21055 (N_21055,N_19917,N_20103);
and U21056 (N_21056,N_20089,N_20102);
xor U21057 (N_21057,N_19506,N_19516);
xnor U21058 (N_21058,N_19928,N_20179);
and U21059 (N_21059,N_19796,N_19503);
nor U21060 (N_21060,N_20241,N_19565);
and U21061 (N_21061,N_20251,N_19840);
nand U21062 (N_21062,N_19425,N_20130);
xor U21063 (N_21063,N_20034,N_20120);
nand U21064 (N_21064,N_20339,N_20051);
and U21065 (N_21065,N_19359,N_20144);
xor U21066 (N_21066,N_20225,N_19349);
nand U21067 (N_21067,N_19915,N_19549);
or U21068 (N_21068,N_20083,N_20169);
and U21069 (N_21069,N_20289,N_19771);
xor U21070 (N_21070,N_19265,N_19388);
or U21071 (N_21071,N_19986,N_19969);
nand U21072 (N_21072,N_20310,N_19856);
nand U21073 (N_21073,N_20199,N_19556);
or U21074 (N_21074,N_19301,N_19636);
xnor U21075 (N_21075,N_20091,N_20210);
or U21076 (N_21076,N_19953,N_19366);
xor U21077 (N_21077,N_19876,N_20367);
nor U21078 (N_21078,N_19608,N_19468);
xor U21079 (N_21079,N_19389,N_20024);
and U21080 (N_21080,N_20394,N_19204);
nand U21081 (N_21081,N_19710,N_20311);
nor U21082 (N_21082,N_19560,N_19993);
nand U21083 (N_21083,N_19851,N_19595);
nand U21084 (N_21084,N_19821,N_19835);
and U21085 (N_21085,N_19364,N_20036);
nand U21086 (N_21086,N_19566,N_20004);
nand U21087 (N_21087,N_19401,N_19463);
and U21088 (N_21088,N_19394,N_19794);
and U21089 (N_21089,N_20005,N_20073);
xnor U21090 (N_21090,N_20089,N_19704);
nor U21091 (N_21091,N_20209,N_19975);
nor U21092 (N_21092,N_19380,N_19515);
and U21093 (N_21093,N_20167,N_20047);
nor U21094 (N_21094,N_19395,N_19603);
or U21095 (N_21095,N_19968,N_20054);
nor U21096 (N_21096,N_20058,N_19682);
nor U21097 (N_21097,N_20192,N_20020);
xnor U21098 (N_21098,N_19212,N_20321);
nor U21099 (N_21099,N_19334,N_19233);
or U21100 (N_21100,N_20349,N_19575);
nand U21101 (N_21101,N_19519,N_19501);
and U21102 (N_21102,N_20316,N_20179);
nor U21103 (N_21103,N_19629,N_19289);
nor U21104 (N_21104,N_19676,N_20339);
and U21105 (N_21105,N_20088,N_19508);
and U21106 (N_21106,N_19927,N_19888);
xnor U21107 (N_21107,N_19445,N_19741);
or U21108 (N_21108,N_19976,N_19747);
xnor U21109 (N_21109,N_19819,N_19633);
xor U21110 (N_21110,N_19532,N_19283);
or U21111 (N_21111,N_19698,N_19694);
xnor U21112 (N_21112,N_19527,N_19751);
nor U21113 (N_21113,N_20080,N_20204);
nor U21114 (N_21114,N_20231,N_19659);
or U21115 (N_21115,N_19840,N_19906);
nand U21116 (N_21116,N_19656,N_20152);
and U21117 (N_21117,N_19401,N_19635);
and U21118 (N_21118,N_19318,N_20253);
nand U21119 (N_21119,N_19512,N_20175);
and U21120 (N_21120,N_20277,N_19352);
and U21121 (N_21121,N_19328,N_19832);
nor U21122 (N_21122,N_19271,N_19907);
and U21123 (N_21123,N_20102,N_19230);
or U21124 (N_21124,N_20197,N_19846);
nand U21125 (N_21125,N_20143,N_19314);
xnor U21126 (N_21126,N_20181,N_20029);
nor U21127 (N_21127,N_19680,N_19638);
nor U21128 (N_21128,N_19513,N_19261);
and U21129 (N_21129,N_19889,N_19937);
nand U21130 (N_21130,N_19468,N_19763);
and U21131 (N_21131,N_19985,N_19244);
or U21132 (N_21132,N_19635,N_19422);
nor U21133 (N_21133,N_19452,N_19444);
nor U21134 (N_21134,N_19661,N_19520);
nor U21135 (N_21135,N_20133,N_20298);
xnor U21136 (N_21136,N_19866,N_19586);
or U21137 (N_21137,N_20273,N_19976);
nor U21138 (N_21138,N_19205,N_19830);
nand U21139 (N_21139,N_19627,N_19912);
nor U21140 (N_21140,N_19517,N_19662);
and U21141 (N_21141,N_19376,N_19937);
xnor U21142 (N_21142,N_19983,N_19959);
and U21143 (N_21143,N_19490,N_20316);
nand U21144 (N_21144,N_19563,N_19327);
xnor U21145 (N_21145,N_19817,N_20398);
or U21146 (N_21146,N_19212,N_19982);
or U21147 (N_21147,N_19502,N_19456);
or U21148 (N_21148,N_19743,N_19661);
xor U21149 (N_21149,N_19261,N_20312);
nor U21150 (N_21150,N_19305,N_20129);
or U21151 (N_21151,N_19302,N_19551);
nand U21152 (N_21152,N_19207,N_20078);
nor U21153 (N_21153,N_19432,N_20102);
and U21154 (N_21154,N_20060,N_19580);
or U21155 (N_21155,N_19281,N_19627);
nor U21156 (N_21156,N_19214,N_20148);
nor U21157 (N_21157,N_19539,N_20373);
or U21158 (N_21158,N_19568,N_19339);
xor U21159 (N_21159,N_19286,N_19556);
or U21160 (N_21160,N_20397,N_20232);
and U21161 (N_21161,N_20208,N_20124);
nand U21162 (N_21162,N_20033,N_20387);
and U21163 (N_21163,N_19887,N_20377);
and U21164 (N_21164,N_20113,N_20246);
nor U21165 (N_21165,N_19523,N_19669);
nor U21166 (N_21166,N_19424,N_19324);
nor U21167 (N_21167,N_19894,N_19860);
nand U21168 (N_21168,N_19432,N_20065);
nand U21169 (N_21169,N_20256,N_19907);
xnor U21170 (N_21170,N_19900,N_20147);
nor U21171 (N_21171,N_19897,N_19956);
and U21172 (N_21172,N_19451,N_19771);
nand U21173 (N_21173,N_19373,N_19789);
and U21174 (N_21174,N_19935,N_20030);
nor U21175 (N_21175,N_20351,N_19941);
xnor U21176 (N_21176,N_19354,N_19661);
xnor U21177 (N_21177,N_19821,N_20203);
or U21178 (N_21178,N_19939,N_20046);
nor U21179 (N_21179,N_19830,N_20125);
or U21180 (N_21180,N_19841,N_20219);
and U21181 (N_21181,N_19634,N_19205);
nand U21182 (N_21182,N_19599,N_20199);
or U21183 (N_21183,N_19572,N_19723);
nand U21184 (N_21184,N_19790,N_19341);
nand U21185 (N_21185,N_20191,N_19671);
or U21186 (N_21186,N_19527,N_19671);
xnor U21187 (N_21187,N_19995,N_20171);
nand U21188 (N_21188,N_19265,N_19329);
nor U21189 (N_21189,N_19991,N_20161);
nand U21190 (N_21190,N_19415,N_19793);
nand U21191 (N_21191,N_19976,N_20093);
and U21192 (N_21192,N_20282,N_19756);
nand U21193 (N_21193,N_19606,N_19396);
and U21194 (N_21194,N_19967,N_19350);
or U21195 (N_21195,N_20035,N_19620);
or U21196 (N_21196,N_19988,N_19833);
or U21197 (N_21197,N_19465,N_19866);
nor U21198 (N_21198,N_19725,N_19297);
xor U21199 (N_21199,N_19315,N_20241);
xnor U21200 (N_21200,N_20226,N_20102);
or U21201 (N_21201,N_20011,N_20162);
or U21202 (N_21202,N_20215,N_19389);
xnor U21203 (N_21203,N_19351,N_19431);
nand U21204 (N_21204,N_20326,N_20282);
xor U21205 (N_21205,N_19234,N_19405);
xor U21206 (N_21206,N_19556,N_19253);
or U21207 (N_21207,N_19434,N_19678);
and U21208 (N_21208,N_19910,N_19334);
nor U21209 (N_21209,N_19880,N_19841);
nor U21210 (N_21210,N_19534,N_19246);
or U21211 (N_21211,N_19616,N_20022);
nand U21212 (N_21212,N_20180,N_20387);
and U21213 (N_21213,N_19672,N_19511);
nand U21214 (N_21214,N_19766,N_20269);
or U21215 (N_21215,N_19565,N_20245);
nor U21216 (N_21216,N_19521,N_20155);
and U21217 (N_21217,N_19220,N_20047);
or U21218 (N_21218,N_19899,N_20357);
or U21219 (N_21219,N_20005,N_19355);
or U21220 (N_21220,N_20147,N_20032);
and U21221 (N_21221,N_19244,N_19891);
nand U21222 (N_21222,N_19320,N_19281);
nand U21223 (N_21223,N_20181,N_19493);
xnor U21224 (N_21224,N_19700,N_19709);
or U21225 (N_21225,N_19240,N_19565);
xor U21226 (N_21226,N_19857,N_20003);
nor U21227 (N_21227,N_19721,N_19357);
xor U21228 (N_21228,N_20030,N_19261);
and U21229 (N_21229,N_20003,N_19812);
xor U21230 (N_21230,N_19465,N_20220);
nand U21231 (N_21231,N_20340,N_19593);
xor U21232 (N_21232,N_20007,N_19990);
nand U21233 (N_21233,N_19721,N_19450);
xor U21234 (N_21234,N_20398,N_20024);
xnor U21235 (N_21235,N_19603,N_19210);
and U21236 (N_21236,N_19298,N_20003);
xnor U21237 (N_21237,N_19404,N_19730);
xor U21238 (N_21238,N_19692,N_19925);
xor U21239 (N_21239,N_20121,N_20114);
xor U21240 (N_21240,N_20052,N_20328);
or U21241 (N_21241,N_20010,N_20087);
nand U21242 (N_21242,N_19273,N_19561);
nand U21243 (N_21243,N_20021,N_20398);
or U21244 (N_21244,N_19245,N_19798);
nor U21245 (N_21245,N_19706,N_19595);
or U21246 (N_21246,N_19901,N_19661);
xnor U21247 (N_21247,N_19247,N_19525);
and U21248 (N_21248,N_19471,N_20337);
nand U21249 (N_21249,N_19331,N_19421);
nor U21250 (N_21250,N_19301,N_19324);
or U21251 (N_21251,N_19945,N_20120);
and U21252 (N_21252,N_20220,N_20354);
xor U21253 (N_21253,N_19829,N_19766);
and U21254 (N_21254,N_19635,N_19560);
nor U21255 (N_21255,N_19821,N_19988);
xnor U21256 (N_21256,N_19724,N_19759);
nor U21257 (N_21257,N_20298,N_19443);
nand U21258 (N_21258,N_20155,N_19893);
or U21259 (N_21259,N_19905,N_19962);
and U21260 (N_21260,N_19960,N_20390);
nand U21261 (N_21261,N_19597,N_19329);
nand U21262 (N_21262,N_19769,N_19765);
nand U21263 (N_21263,N_20248,N_20300);
and U21264 (N_21264,N_19438,N_19545);
and U21265 (N_21265,N_19220,N_19460);
and U21266 (N_21266,N_20206,N_20203);
xor U21267 (N_21267,N_20230,N_19571);
xor U21268 (N_21268,N_19574,N_19469);
xnor U21269 (N_21269,N_19997,N_19737);
nand U21270 (N_21270,N_19714,N_20254);
or U21271 (N_21271,N_19231,N_19339);
nor U21272 (N_21272,N_19478,N_19357);
nor U21273 (N_21273,N_19328,N_19914);
nor U21274 (N_21274,N_19708,N_19927);
or U21275 (N_21275,N_19807,N_19230);
nand U21276 (N_21276,N_20215,N_20104);
or U21277 (N_21277,N_20115,N_19460);
or U21278 (N_21278,N_19250,N_19798);
and U21279 (N_21279,N_19961,N_20179);
nor U21280 (N_21280,N_19751,N_19367);
or U21281 (N_21281,N_19920,N_19366);
xnor U21282 (N_21282,N_19204,N_19897);
or U21283 (N_21283,N_20050,N_20099);
or U21284 (N_21284,N_19778,N_19572);
or U21285 (N_21285,N_19275,N_19407);
xor U21286 (N_21286,N_19484,N_20259);
nand U21287 (N_21287,N_19961,N_19689);
nor U21288 (N_21288,N_20142,N_19255);
and U21289 (N_21289,N_19773,N_19287);
and U21290 (N_21290,N_19349,N_19558);
xnor U21291 (N_21291,N_19611,N_19586);
nor U21292 (N_21292,N_20398,N_19871);
xnor U21293 (N_21293,N_19513,N_19467);
nor U21294 (N_21294,N_20042,N_20052);
nand U21295 (N_21295,N_19794,N_20377);
nor U21296 (N_21296,N_19796,N_19337);
nor U21297 (N_21297,N_19850,N_19545);
nor U21298 (N_21298,N_19568,N_19740);
or U21299 (N_21299,N_19681,N_20252);
and U21300 (N_21300,N_19935,N_19345);
or U21301 (N_21301,N_19952,N_19394);
nand U21302 (N_21302,N_20310,N_19872);
nor U21303 (N_21303,N_19842,N_19361);
and U21304 (N_21304,N_19982,N_19965);
xor U21305 (N_21305,N_19858,N_19890);
xor U21306 (N_21306,N_19491,N_19471);
nand U21307 (N_21307,N_19275,N_19843);
or U21308 (N_21308,N_20207,N_19368);
xnor U21309 (N_21309,N_19221,N_20096);
nor U21310 (N_21310,N_20270,N_19480);
or U21311 (N_21311,N_19877,N_19768);
xnor U21312 (N_21312,N_20212,N_19606);
or U21313 (N_21313,N_20026,N_19529);
nor U21314 (N_21314,N_19847,N_19986);
and U21315 (N_21315,N_20173,N_19730);
xnor U21316 (N_21316,N_19499,N_19952);
or U21317 (N_21317,N_19834,N_19872);
and U21318 (N_21318,N_20341,N_19346);
and U21319 (N_21319,N_19863,N_19595);
xor U21320 (N_21320,N_19679,N_20349);
or U21321 (N_21321,N_20027,N_19545);
or U21322 (N_21322,N_19755,N_20366);
and U21323 (N_21323,N_19785,N_20176);
nand U21324 (N_21324,N_19581,N_19968);
nor U21325 (N_21325,N_19463,N_19772);
xnor U21326 (N_21326,N_20362,N_19334);
xor U21327 (N_21327,N_20222,N_20137);
xnor U21328 (N_21328,N_19273,N_20382);
nand U21329 (N_21329,N_19317,N_19687);
xnor U21330 (N_21330,N_19698,N_19706);
or U21331 (N_21331,N_19963,N_19219);
or U21332 (N_21332,N_19798,N_19440);
xnor U21333 (N_21333,N_19311,N_19426);
nand U21334 (N_21334,N_19472,N_19946);
and U21335 (N_21335,N_19463,N_19273);
and U21336 (N_21336,N_19876,N_19621);
or U21337 (N_21337,N_19606,N_20272);
xor U21338 (N_21338,N_20208,N_20267);
and U21339 (N_21339,N_19807,N_20365);
xnor U21340 (N_21340,N_20083,N_19319);
nand U21341 (N_21341,N_20255,N_20333);
or U21342 (N_21342,N_20352,N_19861);
nor U21343 (N_21343,N_20385,N_20045);
xor U21344 (N_21344,N_20258,N_20092);
nor U21345 (N_21345,N_19897,N_19552);
or U21346 (N_21346,N_19225,N_20131);
nand U21347 (N_21347,N_19688,N_19866);
nand U21348 (N_21348,N_19493,N_20370);
nand U21349 (N_21349,N_19899,N_19988);
or U21350 (N_21350,N_19651,N_20302);
nand U21351 (N_21351,N_19314,N_19207);
xnor U21352 (N_21352,N_20215,N_20320);
and U21353 (N_21353,N_19641,N_19558);
nand U21354 (N_21354,N_19475,N_19313);
and U21355 (N_21355,N_20078,N_19534);
nand U21356 (N_21356,N_20324,N_19857);
nor U21357 (N_21357,N_19861,N_20069);
or U21358 (N_21358,N_19424,N_19217);
and U21359 (N_21359,N_19776,N_20358);
or U21360 (N_21360,N_20174,N_19996);
or U21361 (N_21361,N_20367,N_19932);
nor U21362 (N_21362,N_19626,N_19608);
nand U21363 (N_21363,N_19889,N_19469);
xor U21364 (N_21364,N_19520,N_19788);
or U21365 (N_21365,N_20357,N_19512);
nand U21366 (N_21366,N_20072,N_20076);
xnor U21367 (N_21367,N_19514,N_19283);
nand U21368 (N_21368,N_19337,N_19709);
nor U21369 (N_21369,N_19920,N_19434);
nand U21370 (N_21370,N_19322,N_20373);
xnor U21371 (N_21371,N_19650,N_19579);
and U21372 (N_21372,N_19730,N_20060);
xnor U21373 (N_21373,N_19516,N_19400);
nand U21374 (N_21374,N_19635,N_19602);
xor U21375 (N_21375,N_19473,N_19878);
and U21376 (N_21376,N_19918,N_19396);
nand U21377 (N_21377,N_19287,N_19226);
and U21378 (N_21378,N_19871,N_19546);
or U21379 (N_21379,N_19600,N_19213);
xnor U21380 (N_21380,N_19904,N_19954);
and U21381 (N_21381,N_20303,N_20193);
or U21382 (N_21382,N_19257,N_19595);
and U21383 (N_21383,N_20218,N_20180);
xnor U21384 (N_21384,N_19659,N_20174);
and U21385 (N_21385,N_19253,N_19962);
or U21386 (N_21386,N_19956,N_20305);
nor U21387 (N_21387,N_19887,N_20127);
nand U21388 (N_21388,N_19950,N_20146);
xor U21389 (N_21389,N_19328,N_19949);
nand U21390 (N_21390,N_19875,N_20394);
nor U21391 (N_21391,N_19249,N_20115);
xnor U21392 (N_21392,N_20169,N_19761);
xor U21393 (N_21393,N_20117,N_19676);
or U21394 (N_21394,N_19378,N_19573);
nor U21395 (N_21395,N_19216,N_19712);
xnor U21396 (N_21396,N_19909,N_19349);
and U21397 (N_21397,N_20283,N_20184);
or U21398 (N_21398,N_20081,N_19387);
or U21399 (N_21399,N_19726,N_20017);
xnor U21400 (N_21400,N_19840,N_19233);
or U21401 (N_21401,N_20228,N_19662);
nand U21402 (N_21402,N_19549,N_19574);
and U21403 (N_21403,N_20093,N_19458);
and U21404 (N_21404,N_19742,N_19448);
nor U21405 (N_21405,N_19804,N_19734);
nor U21406 (N_21406,N_19415,N_20089);
nor U21407 (N_21407,N_19742,N_19867);
nand U21408 (N_21408,N_19962,N_19246);
nor U21409 (N_21409,N_19847,N_19394);
or U21410 (N_21410,N_19306,N_19687);
or U21411 (N_21411,N_19227,N_19956);
nand U21412 (N_21412,N_20398,N_19688);
nand U21413 (N_21413,N_20181,N_19313);
and U21414 (N_21414,N_19884,N_19973);
or U21415 (N_21415,N_19408,N_20001);
xnor U21416 (N_21416,N_20081,N_19800);
nor U21417 (N_21417,N_19893,N_19794);
xnor U21418 (N_21418,N_19261,N_20075);
nor U21419 (N_21419,N_19474,N_20370);
or U21420 (N_21420,N_19727,N_20121);
xor U21421 (N_21421,N_19478,N_19627);
or U21422 (N_21422,N_19368,N_20079);
xor U21423 (N_21423,N_19598,N_19281);
and U21424 (N_21424,N_19340,N_20301);
and U21425 (N_21425,N_19641,N_19892);
or U21426 (N_21426,N_19700,N_19654);
or U21427 (N_21427,N_20249,N_20124);
nor U21428 (N_21428,N_19953,N_19525);
nor U21429 (N_21429,N_19348,N_20049);
and U21430 (N_21430,N_19219,N_19245);
xnor U21431 (N_21431,N_19624,N_19626);
nand U21432 (N_21432,N_19591,N_19277);
nor U21433 (N_21433,N_20053,N_20387);
or U21434 (N_21434,N_19201,N_20234);
nand U21435 (N_21435,N_19203,N_20147);
or U21436 (N_21436,N_19327,N_20327);
xor U21437 (N_21437,N_20339,N_19296);
xnor U21438 (N_21438,N_20046,N_20126);
and U21439 (N_21439,N_19590,N_20336);
nor U21440 (N_21440,N_20250,N_19334);
and U21441 (N_21441,N_20334,N_19785);
nor U21442 (N_21442,N_20131,N_20141);
or U21443 (N_21443,N_20208,N_19771);
or U21444 (N_21444,N_19480,N_19215);
nor U21445 (N_21445,N_19706,N_20123);
nand U21446 (N_21446,N_19523,N_19945);
and U21447 (N_21447,N_19832,N_19956);
nor U21448 (N_21448,N_19476,N_19634);
nor U21449 (N_21449,N_19224,N_20020);
and U21450 (N_21450,N_20215,N_20117);
and U21451 (N_21451,N_19567,N_20162);
and U21452 (N_21452,N_19627,N_20031);
xor U21453 (N_21453,N_19412,N_19349);
or U21454 (N_21454,N_19630,N_20191);
and U21455 (N_21455,N_20014,N_20089);
and U21456 (N_21456,N_20339,N_19308);
or U21457 (N_21457,N_20262,N_19552);
or U21458 (N_21458,N_19778,N_20086);
or U21459 (N_21459,N_19348,N_19216);
nand U21460 (N_21460,N_20277,N_19842);
nand U21461 (N_21461,N_19274,N_19983);
and U21462 (N_21462,N_20333,N_19425);
or U21463 (N_21463,N_20356,N_20084);
or U21464 (N_21464,N_19403,N_20344);
nor U21465 (N_21465,N_20124,N_19390);
nand U21466 (N_21466,N_19675,N_19972);
nor U21467 (N_21467,N_19751,N_19292);
nor U21468 (N_21468,N_19797,N_20182);
and U21469 (N_21469,N_19833,N_19355);
xor U21470 (N_21470,N_19332,N_19246);
nand U21471 (N_21471,N_19835,N_20255);
or U21472 (N_21472,N_19232,N_19535);
xor U21473 (N_21473,N_20281,N_19976);
and U21474 (N_21474,N_19829,N_19585);
xnor U21475 (N_21475,N_19619,N_19747);
and U21476 (N_21476,N_20386,N_20247);
nor U21477 (N_21477,N_20305,N_19483);
nand U21478 (N_21478,N_19669,N_19526);
or U21479 (N_21479,N_19751,N_19957);
nor U21480 (N_21480,N_20141,N_20050);
xor U21481 (N_21481,N_20268,N_20220);
and U21482 (N_21482,N_19635,N_19693);
xnor U21483 (N_21483,N_19316,N_20012);
and U21484 (N_21484,N_19612,N_19528);
nand U21485 (N_21485,N_20080,N_19281);
xor U21486 (N_21486,N_19610,N_20228);
nand U21487 (N_21487,N_19620,N_19888);
and U21488 (N_21488,N_19617,N_19635);
nor U21489 (N_21489,N_19397,N_19836);
xor U21490 (N_21490,N_19561,N_20110);
nand U21491 (N_21491,N_19416,N_19598);
xnor U21492 (N_21492,N_19923,N_20019);
xnor U21493 (N_21493,N_19749,N_19887);
xnor U21494 (N_21494,N_20197,N_19484);
or U21495 (N_21495,N_20069,N_20008);
and U21496 (N_21496,N_19528,N_20344);
or U21497 (N_21497,N_19942,N_19899);
nor U21498 (N_21498,N_19408,N_19602);
and U21499 (N_21499,N_20391,N_19647);
or U21500 (N_21500,N_19249,N_20227);
or U21501 (N_21501,N_19316,N_19571);
or U21502 (N_21502,N_19769,N_19916);
xor U21503 (N_21503,N_20250,N_19870);
nand U21504 (N_21504,N_20371,N_19591);
or U21505 (N_21505,N_20206,N_19212);
or U21506 (N_21506,N_19368,N_19909);
or U21507 (N_21507,N_19866,N_19917);
nor U21508 (N_21508,N_19580,N_19502);
and U21509 (N_21509,N_19812,N_19311);
xnor U21510 (N_21510,N_19450,N_19743);
and U21511 (N_21511,N_20296,N_20085);
and U21512 (N_21512,N_20102,N_19556);
and U21513 (N_21513,N_19483,N_19717);
xor U21514 (N_21514,N_19898,N_19670);
nand U21515 (N_21515,N_20378,N_19340);
nand U21516 (N_21516,N_19613,N_19417);
xor U21517 (N_21517,N_19572,N_20220);
and U21518 (N_21518,N_19615,N_19454);
xnor U21519 (N_21519,N_19780,N_19454);
nand U21520 (N_21520,N_19549,N_19360);
xor U21521 (N_21521,N_19390,N_19330);
xnor U21522 (N_21522,N_19351,N_19484);
and U21523 (N_21523,N_19560,N_19384);
and U21524 (N_21524,N_19551,N_19884);
and U21525 (N_21525,N_20115,N_19650);
xor U21526 (N_21526,N_19643,N_19591);
xnor U21527 (N_21527,N_19529,N_20170);
nor U21528 (N_21528,N_20103,N_19267);
nor U21529 (N_21529,N_19205,N_19660);
and U21530 (N_21530,N_20174,N_20168);
nor U21531 (N_21531,N_19388,N_19974);
and U21532 (N_21532,N_20067,N_19897);
xnor U21533 (N_21533,N_19286,N_19314);
or U21534 (N_21534,N_19628,N_19871);
xnor U21535 (N_21535,N_19884,N_20207);
and U21536 (N_21536,N_20103,N_19338);
and U21537 (N_21537,N_20353,N_19922);
nand U21538 (N_21538,N_20318,N_20037);
nor U21539 (N_21539,N_19254,N_19677);
nand U21540 (N_21540,N_20395,N_19255);
or U21541 (N_21541,N_19403,N_20322);
and U21542 (N_21542,N_19450,N_19409);
nand U21543 (N_21543,N_19889,N_19585);
xor U21544 (N_21544,N_19455,N_20177);
nand U21545 (N_21545,N_20112,N_19388);
nor U21546 (N_21546,N_19932,N_20278);
nand U21547 (N_21547,N_20372,N_19795);
xor U21548 (N_21548,N_19496,N_19673);
nor U21549 (N_21549,N_20382,N_20087);
nor U21550 (N_21550,N_19926,N_20150);
nor U21551 (N_21551,N_19632,N_19985);
xnor U21552 (N_21552,N_19349,N_20146);
and U21553 (N_21553,N_19503,N_19490);
xor U21554 (N_21554,N_20060,N_19480);
or U21555 (N_21555,N_19294,N_19989);
or U21556 (N_21556,N_19832,N_20262);
nor U21557 (N_21557,N_19731,N_20046);
nand U21558 (N_21558,N_20314,N_20210);
or U21559 (N_21559,N_19538,N_20352);
nor U21560 (N_21560,N_19251,N_19491);
xor U21561 (N_21561,N_19872,N_19433);
xor U21562 (N_21562,N_19388,N_20078);
and U21563 (N_21563,N_19343,N_19309);
or U21564 (N_21564,N_19339,N_19860);
nor U21565 (N_21565,N_19303,N_19348);
xor U21566 (N_21566,N_19756,N_19382);
and U21567 (N_21567,N_19205,N_20268);
xor U21568 (N_21568,N_19576,N_19571);
xor U21569 (N_21569,N_19578,N_19298);
nor U21570 (N_21570,N_19893,N_19346);
and U21571 (N_21571,N_19382,N_19431);
nand U21572 (N_21572,N_20043,N_19353);
xnor U21573 (N_21573,N_19249,N_19258);
and U21574 (N_21574,N_19707,N_19245);
nor U21575 (N_21575,N_19446,N_19486);
xor U21576 (N_21576,N_20132,N_20162);
nor U21577 (N_21577,N_20020,N_19916);
nand U21578 (N_21578,N_20057,N_20303);
or U21579 (N_21579,N_20139,N_19290);
nor U21580 (N_21580,N_20109,N_19688);
nor U21581 (N_21581,N_20170,N_20294);
xnor U21582 (N_21582,N_19236,N_20284);
nor U21583 (N_21583,N_19824,N_20289);
or U21584 (N_21584,N_20223,N_19583);
nand U21585 (N_21585,N_19501,N_19454);
nor U21586 (N_21586,N_19654,N_19929);
or U21587 (N_21587,N_19903,N_20228);
nor U21588 (N_21588,N_19625,N_19398);
nand U21589 (N_21589,N_19268,N_19985);
nand U21590 (N_21590,N_19421,N_19578);
and U21591 (N_21591,N_19497,N_19216);
nand U21592 (N_21592,N_20143,N_20323);
nor U21593 (N_21593,N_19356,N_19513);
xor U21594 (N_21594,N_19227,N_20039);
or U21595 (N_21595,N_20330,N_20126);
xor U21596 (N_21596,N_19487,N_20038);
nand U21597 (N_21597,N_19698,N_19926);
xnor U21598 (N_21598,N_19333,N_20213);
xnor U21599 (N_21599,N_20358,N_19853);
xor U21600 (N_21600,N_20628,N_21192);
or U21601 (N_21601,N_21266,N_21528);
and U21602 (N_21602,N_21015,N_21225);
nand U21603 (N_21603,N_20931,N_20783);
or U21604 (N_21604,N_20961,N_20774);
xor U21605 (N_21605,N_21345,N_21205);
and U21606 (N_21606,N_20549,N_21160);
xor U21607 (N_21607,N_20976,N_20901);
and U21608 (N_21608,N_20758,N_21170);
nor U21609 (N_21609,N_21348,N_21276);
xnor U21610 (N_21610,N_20874,N_21038);
nand U21611 (N_21611,N_21124,N_21508);
xnor U21612 (N_21612,N_20462,N_21434);
nand U21613 (N_21613,N_20975,N_21327);
or U21614 (N_21614,N_20969,N_21369);
and U21615 (N_21615,N_20442,N_20686);
nand U21616 (N_21616,N_21544,N_20737);
and U21617 (N_21617,N_21486,N_21041);
xor U21618 (N_21618,N_20814,N_21207);
or U21619 (N_21619,N_21010,N_20435);
or U21620 (N_21620,N_20721,N_20476);
and U21621 (N_21621,N_20830,N_20810);
nand U21622 (N_21622,N_20932,N_20775);
or U21623 (N_21623,N_20616,N_21495);
xnor U21624 (N_21624,N_20643,N_21011);
nand U21625 (N_21625,N_20727,N_21231);
and U21626 (N_21626,N_21248,N_20599);
nand U21627 (N_21627,N_21334,N_20589);
and U21628 (N_21628,N_21379,N_20834);
nor U21629 (N_21629,N_21338,N_20711);
nand U21630 (N_21630,N_20873,N_20920);
and U21631 (N_21631,N_21537,N_20909);
or U21632 (N_21632,N_20658,N_21412);
nand U21633 (N_21633,N_21573,N_21259);
and U21634 (N_21634,N_21216,N_20983);
nand U21635 (N_21635,N_21569,N_20576);
xnor U21636 (N_21636,N_20905,N_21430);
nor U21637 (N_21637,N_21553,N_21070);
nand U21638 (N_21638,N_21193,N_20743);
nand U21639 (N_21639,N_20703,N_21106);
and U21640 (N_21640,N_21415,N_21197);
xor U21641 (N_21641,N_21286,N_21488);
or U21642 (N_21642,N_20866,N_20937);
xor U21643 (N_21643,N_20844,N_21101);
nand U21644 (N_21644,N_20763,N_21213);
nor U21645 (N_21645,N_20620,N_21319);
or U21646 (N_21646,N_21526,N_20893);
nor U21647 (N_21647,N_21202,N_20872);
or U21648 (N_21648,N_20865,N_20537);
and U21649 (N_21649,N_21409,N_20451);
nor U21650 (N_21650,N_21318,N_21222);
and U21651 (N_21651,N_21543,N_20779);
nand U21652 (N_21652,N_20608,N_21227);
and U21653 (N_21653,N_21516,N_21463);
xnor U21654 (N_21654,N_20971,N_20887);
nor U21655 (N_21655,N_21159,N_21075);
nor U21656 (N_21656,N_20416,N_21140);
and U21657 (N_21657,N_20559,N_21191);
xor U21658 (N_21658,N_20452,N_20765);
or U21659 (N_21659,N_20815,N_21051);
xor U21660 (N_21660,N_21068,N_21313);
nand U21661 (N_21661,N_20696,N_20515);
and U21662 (N_21662,N_20657,N_20527);
nor U21663 (N_21663,N_21574,N_20835);
nor U21664 (N_21664,N_21314,N_21034);
nor U21665 (N_21665,N_20792,N_20558);
nor U21666 (N_21666,N_20430,N_21462);
nand U21667 (N_21667,N_21292,N_21400);
nand U21668 (N_21668,N_21432,N_21558);
nor U21669 (N_21669,N_21132,N_20736);
nor U21670 (N_21670,N_21477,N_20454);
and U21671 (N_21671,N_20767,N_21237);
or U21672 (N_21672,N_20544,N_20676);
nor U21673 (N_21673,N_21293,N_20572);
nand U21674 (N_21674,N_21572,N_20539);
xor U21675 (N_21675,N_21530,N_20456);
and U21676 (N_21676,N_20904,N_21211);
nand U21677 (N_21677,N_20738,N_21523);
nor U21678 (N_21678,N_20761,N_20922);
and U21679 (N_21679,N_21550,N_21282);
nand U21680 (N_21680,N_20974,N_20913);
or U21681 (N_21681,N_21448,N_20541);
or U21682 (N_21682,N_20751,N_21290);
nand U21683 (N_21683,N_21176,N_20916);
xor U21684 (N_21684,N_20784,N_20739);
and U21685 (N_21685,N_20970,N_21130);
and U21686 (N_21686,N_21531,N_21499);
nand U21687 (N_21687,N_21509,N_20843);
nand U21688 (N_21688,N_21308,N_21118);
xor U21689 (N_21689,N_20745,N_20989);
nor U21690 (N_21690,N_20998,N_21032);
nand U21691 (N_21691,N_21435,N_21552);
nand U21692 (N_21692,N_20687,N_21532);
nand U21693 (N_21693,N_20554,N_20584);
nand U21694 (N_21694,N_21316,N_21556);
or U21695 (N_21695,N_20595,N_21304);
or U21696 (N_21696,N_20458,N_21006);
and U21697 (N_21697,N_21299,N_20663);
or U21698 (N_21698,N_21458,N_20566);
nand U21699 (N_21699,N_21446,N_20809);
nand U21700 (N_21700,N_21263,N_20827);
nand U21701 (N_21701,N_21347,N_21000);
nand U21702 (N_21702,N_20940,N_21410);
and U21703 (N_21703,N_20871,N_21152);
nand U21704 (N_21704,N_21171,N_20440);
or U21705 (N_21705,N_21464,N_20591);
nor U21706 (N_21706,N_20886,N_21440);
xor U21707 (N_21707,N_21228,N_20606);
xnor U21708 (N_21708,N_20944,N_20627);
and U21709 (N_21709,N_20512,N_21284);
nor U21710 (N_21710,N_21009,N_21444);
nand U21711 (N_21711,N_20613,N_20517);
or U21712 (N_21712,N_21534,N_21538);
nand U21713 (N_21713,N_20694,N_21283);
or U21714 (N_21714,N_20744,N_20762);
and U21715 (N_21715,N_20542,N_20640);
xnor U21716 (N_21716,N_21247,N_21012);
or U21717 (N_21717,N_21058,N_21360);
and U21718 (N_21718,N_21264,N_21483);
and U21719 (N_21719,N_21023,N_21273);
xnor U21720 (N_21720,N_21503,N_20828);
and U21721 (N_21721,N_20609,N_20860);
nand U21722 (N_21722,N_20802,N_20884);
nor U21723 (N_21723,N_21529,N_20882);
and U21724 (N_21724,N_21461,N_21147);
nand U21725 (N_21725,N_21168,N_21076);
or U21726 (N_21726,N_20548,N_20641);
nor U21727 (N_21727,N_20956,N_20618);
and U21728 (N_21728,N_20417,N_21540);
nand U21729 (N_21729,N_20695,N_21235);
and U21730 (N_21730,N_21129,N_20593);
nand U21731 (N_21731,N_21351,N_21148);
or U21732 (N_21732,N_21405,N_21279);
xor U21733 (N_21733,N_21481,N_21172);
or U21734 (N_21734,N_21593,N_20723);
nand U21735 (N_21735,N_20497,N_20853);
nor U21736 (N_21736,N_20679,N_21219);
and U21737 (N_21737,N_21100,N_21524);
nand U21738 (N_21738,N_21494,N_20521);
and U21739 (N_21739,N_20448,N_21372);
nor U21740 (N_21740,N_20941,N_21115);
nor U21741 (N_21741,N_21303,N_21403);
or U21742 (N_21742,N_21019,N_20741);
nor U21743 (N_21743,N_20982,N_21332);
and U21744 (N_21744,N_21103,N_21389);
and U21745 (N_21745,N_21423,N_21510);
nand U21746 (N_21746,N_21598,N_21418);
nand U21747 (N_21747,N_21257,N_20449);
nor U21748 (N_21748,N_21567,N_21217);
xnor U21749 (N_21749,N_20413,N_21485);
nand U21750 (N_21750,N_20551,N_20499);
or U21751 (N_21751,N_20660,N_21088);
nor U21752 (N_21752,N_21066,N_21121);
nor U21753 (N_21753,N_20863,N_20612);
and U21754 (N_21754,N_20780,N_20807);
xor U21755 (N_21755,N_21554,N_20622);
xor U21756 (N_21756,N_21224,N_21595);
xnor U21757 (N_21757,N_20771,N_21511);
and U21758 (N_21758,N_20928,N_20670);
xor U21759 (N_21759,N_21295,N_21004);
and U21760 (N_21760,N_20796,N_20420);
xor U21761 (N_21761,N_21594,N_20691);
and U21762 (N_21762,N_20546,N_21375);
nand U21763 (N_21763,N_20564,N_21204);
xnor U21764 (N_21764,N_20474,N_20978);
and U21765 (N_21765,N_21230,N_21086);
or U21766 (N_21766,N_21186,N_21396);
nor U21767 (N_21767,N_21194,N_20858);
and U21768 (N_21768,N_20602,N_20519);
xnor U21769 (N_21769,N_21097,N_20506);
xnor U21770 (N_21770,N_21244,N_21126);
or U21771 (N_21771,N_20685,N_21465);
nor U21772 (N_21772,N_21312,N_21460);
xnor U21773 (N_21773,N_20649,N_21122);
or U21774 (N_21774,N_21081,N_20848);
or U21775 (N_21775,N_21320,N_20475);
and U21776 (N_21776,N_21575,N_21095);
xnor U21777 (N_21777,N_20678,N_21358);
xnor U21778 (N_21778,N_20414,N_21561);
or U21779 (N_21779,N_21035,N_21336);
or U21780 (N_21780,N_20650,N_21242);
nand U21781 (N_21781,N_20583,N_21424);
nor U21782 (N_21782,N_21031,N_21104);
nand U21783 (N_21783,N_21374,N_21245);
or U21784 (N_21784,N_20817,N_20428);
and U21785 (N_21785,N_21018,N_20592);
nand U21786 (N_21786,N_20733,N_21394);
and U21787 (N_21787,N_20625,N_20634);
and U21788 (N_21788,N_21373,N_20725);
and U21789 (N_21789,N_21519,N_20524);
nand U21790 (N_21790,N_20820,N_20750);
or U21791 (N_21791,N_20457,N_21107);
xnor U21792 (N_21792,N_21057,N_20411);
xor U21793 (N_21793,N_20522,N_21102);
nor U21794 (N_21794,N_20481,N_21089);
nand U21795 (N_21795,N_20494,N_20410);
or U21796 (N_21796,N_21028,N_21143);
nor U21797 (N_21797,N_20925,N_20405);
or U21798 (N_21798,N_21053,N_20438);
xor U21799 (N_21799,N_21493,N_20629);
xor U21800 (N_21800,N_20688,N_21046);
nand U21801 (N_21801,N_20590,N_20850);
nand U21802 (N_21802,N_20984,N_21223);
and U21803 (N_21803,N_20759,N_21069);
and U21804 (N_21804,N_20671,N_20423);
or U21805 (N_21805,N_20700,N_20735);
or U21806 (N_21806,N_21232,N_21220);
and U21807 (N_21807,N_20652,N_20706);
xor U21808 (N_21808,N_20536,N_20516);
and U21809 (N_21809,N_21149,N_20637);
xnor U21810 (N_21810,N_20776,N_20710);
nand U21811 (N_21811,N_20614,N_20578);
nand U21812 (N_21812,N_20406,N_20580);
nand U21813 (N_21813,N_21185,N_20885);
nand U21814 (N_21814,N_21215,N_20681);
or U21815 (N_21815,N_21047,N_20588);
xor U21816 (N_21816,N_20547,N_20868);
nand U21817 (N_21817,N_21001,N_20797);
or U21818 (N_21818,N_20846,N_21527);
and U21819 (N_21819,N_20579,N_21346);
and U21820 (N_21820,N_21354,N_20919);
or U21821 (N_21821,N_21475,N_20556);
nor U21822 (N_21822,N_21457,N_21470);
nand U21823 (N_21823,N_21431,N_21274);
or U21824 (N_21824,N_21560,N_21408);
nor U21825 (N_21825,N_21398,N_20917);
or U21826 (N_21826,N_20952,N_21178);
or U21827 (N_21827,N_21134,N_21388);
and U21828 (N_21828,N_21269,N_21512);
xnor U21829 (N_21829,N_21335,N_20450);
or U21830 (N_21830,N_20669,N_20824);
xor U21831 (N_21831,N_21184,N_21189);
nand U21832 (N_21832,N_21566,N_21155);
xor U21833 (N_21833,N_20740,N_20630);
or U21834 (N_21834,N_20540,N_20404);
and U21835 (N_21835,N_21326,N_21533);
xor U21836 (N_21836,N_20436,N_20415);
xor U21837 (N_21837,N_20714,N_20453);
or U21838 (N_21838,N_20907,N_21391);
xor U21839 (N_21839,N_21490,N_20503);
or U21840 (N_21840,N_21417,N_20673);
nand U21841 (N_21841,N_21449,N_20994);
xnor U21842 (N_21842,N_20662,N_20891);
or U21843 (N_21843,N_21513,N_20877);
xnor U21844 (N_21844,N_21551,N_21007);
and U21845 (N_21845,N_20471,N_21505);
nor U21846 (N_21846,N_20664,N_20626);
or U21847 (N_21847,N_20949,N_20756);
xor U21848 (N_21848,N_21061,N_20930);
xor U21849 (N_21849,N_20441,N_21381);
and U21850 (N_21850,N_21339,N_20400);
xnor U21851 (N_21851,N_21411,N_21386);
and U21852 (N_21852,N_21507,N_20666);
xor U21853 (N_21853,N_20926,N_21164);
nor U21854 (N_21854,N_20432,N_20621);
xnor U21855 (N_21855,N_21397,N_21447);
nand U21856 (N_21856,N_20644,N_21246);
and U21857 (N_21857,N_21071,N_21474);
and U21858 (N_21858,N_21166,N_20854);
nand U21859 (N_21859,N_20601,N_21317);
or U21860 (N_21860,N_21361,N_21144);
and U21861 (N_21861,N_21040,N_21281);
or U21862 (N_21862,N_21413,N_21298);
nand U21863 (N_21863,N_21514,N_20507);
nand U21864 (N_21864,N_21436,N_20942);
nor U21865 (N_21865,N_21310,N_20419);
nand U21866 (N_21866,N_21323,N_21277);
or U21867 (N_21867,N_21063,N_21250);
or U21868 (N_21868,N_21016,N_20842);
nor U21869 (N_21869,N_21506,N_20624);
and U21870 (N_21870,N_20734,N_20800);
and U21871 (N_21871,N_20480,N_20955);
and U21872 (N_21872,N_20560,N_21406);
or U21873 (N_21873,N_21401,N_21133);
nor U21874 (N_21874,N_20674,N_20680);
nor U21875 (N_21875,N_20794,N_20823);
nand U21876 (N_21876,N_20513,N_20829);
xnor U21877 (N_21877,N_21201,N_21022);
xnor U21878 (N_21878,N_21060,N_20742);
nand U21879 (N_21879,N_20996,N_20728);
nand U21880 (N_21880,N_20689,N_21173);
xnor U21881 (N_21881,N_20988,N_20408);
nor U21882 (N_21882,N_20668,N_21517);
xor U21883 (N_21883,N_21294,N_21128);
xor U21884 (N_21884,N_20492,N_20957);
xor U21885 (N_21885,N_20791,N_21082);
xor U21886 (N_21886,N_20833,N_20642);
nand U21887 (N_21887,N_20466,N_21175);
xor U21888 (N_21888,N_20782,N_21003);
and U21889 (N_21889,N_21330,N_21062);
or U21890 (N_21890,N_20712,N_20575);
nand U21891 (N_21891,N_21482,N_20532);
nor U21892 (N_21892,N_21542,N_21226);
nand U21893 (N_21893,N_20439,N_21065);
nor U21894 (N_21894,N_21145,N_21467);
xnor U21895 (N_21895,N_20838,N_21238);
nand U21896 (N_21896,N_21045,N_20656);
and U21897 (N_21897,N_21289,N_20550);
xor U21898 (N_21898,N_20585,N_20493);
nor U21899 (N_21899,N_20699,N_20973);
or U21900 (N_21900,N_21139,N_21562);
nand U21901 (N_21901,N_21450,N_20505);
or U21902 (N_21902,N_21218,N_20535);
nor U21903 (N_21903,N_21547,N_21402);
nand U21904 (N_21904,N_20409,N_20773);
and U21905 (N_21905,N_21301,N_21592);
nand U21906 (N_21906,N_21198,N_20708);
or U21907 (N_21907,N_20713,N_20489);
xor U21908 (N_21908,N_20953,N_20772);
and U21909 (N_21909,N_21029,N_20897);
or U21910 (N_21910,N_20748,N_20862);
xor U21911 (N_21911,N_20446,N_20443);
and U21912 (N_21912,N_20615,N_20808);
xnor U21913 (N_21913,N_20473,N_20752);
or U21914 (N_21914,N_21052,N_20651);
and U21915 (N_21915,N_21200,N_20943);
xor U21916 (N_21916,N_21137,N_20667);
nand U21917 (N_21917,N_21174,N_21548);
and U21918 (N_21918,N_21119,N_21331);
xnor U21919 (N_21919,N_20993,N_20757);
nor U21920 (N_21920,N_20875,N_20465);
or U21921 (N_21921,N_21492,N_20545);
xor U21922 (N_21922,N_20531,N_21253);
and U21923 (N_21923,N_21048,N_20935);
nor U21924 (N_21924,N_20718,N_20870);
and U21925 (N_21925,N_21067,N_21039);
xnor U21926 (N_21926,N_21262,N_21091);
nand U21927 (N_21927,N_20604,N_21305);
nor U21928 (N_21928,N_20484,N_21350);
and U21929 (N_21929,N_20571,N_21385);
nand U21930 (N_21930,N_20799,N_20929);
nor U21931 (N_21931,N_21181,N_20729);
and U21932 (N_21932,N_21559,N_21329);
nand U21933 (N_21933,N_20698,N_21570);
nand U21934 (N_21934,N_21555,N_20760);
and U21935 (N_21935,N_21116,N_20661);
xor U21936 (N_21936,N_21291,N_21296);
nor U21937 (N_21937,N_21251,N_20684);
or U21938 (N_21938,N_20888,N_20654);
nor U21939 (N_21939,N_21014,N_21399);
xor U21940 (N_21940,N_21362,N_20908);
or U21941 (N_21941,N_21545,N_21206);
or U21942 (N_21942,N_21437,N_21254);
xnor U21943 (N_21943,N_20407,N_21599);
or U21944 (N_21944,N_21501,N_21363);
nand U21945 (N_21945,N_20965,N_21280);
nand U21946 (N_21946,N_20495,N_20582);
nor U21947 (N_21947,N_21341,N_21328);
and U21948 (N_21948,N_21142,N_21229);
and U21949 (N_21949,N_21256,N_21117);
nand U21950 (N_21950,N_21110,N_21453);
or U21951 (N_21951,N_21025,N_21199);
nand U21952 (N_21952,N_21576,N_21487);
or U21953 (N_21953,N_20895,N_21210);
xnor U21954 (N_21954,N_20594,N_21300);
nand U21955 (N_21955,N_21468,N_20402);
nor U21956 (N_21956,N_21577,N_21151);
xor U21957 (N_21957,N_21195,N_20951);
or U21958 (N_21958,N_21187,N_20825);
nor U21959 (N_21959,N_21472,N_20704);
and U21960 (N_21960,N_21518,N_20999);
nand U21961 (N_21961,N_20979,N_20880);
and U21962 (N_21962,N_21473,N_20730);
nor U21963 (N_21963,N_21272,N_20847);
xor U21964 (N_21964,N_20501,N_21582);
nand U21965 (N_21965,N_20682,N_21212);
nand U21966 (N_21966,N_20665,N_20509);
or U21967 (N_21967,N_20529,N_20839);
nor U21968 (N_21968,N_21208,N_20574);
and U21969 (N_21969,N_20633,N_21271);
and U21970 (N_21970,N_21491,N_20869);
and U21971 (N_21971,N_21055,N_21416);
or U21972 (N_21972,N_21096,N_21368);
nand U21973 (N_21973,N_20502,N_20798);
and U21974 (N_21974,N_20990,N_21563);
xor U21975 (N_21975,N_21020,N_20992);
nand U21976 (N_21976,N_20938,N_20470);
xnor U21977 (N_21977,N_21017,N_20463);
nand U21978 (N_21978,N_20921,N_21270);
or U21979 (N_21979,N_20849,N_21169);
xor U21980 (N_21980,N_21469,N_20504);
xnor U21981 (N_21981,N_20597,N_20605);
xnor U21982 (N_21982,N_21322,N_21059);
nand U21983 (N_21983,N_20581,N_20732);
nand U21984 (N_21984,N_20500,N_20822);
nand U21985 (N_21985,N_21421,N_20459);
nor U21986 (N_21986,N_20861,N_20526);
nor U21987 (N_21987,N_20562,N_21158);
and U21988 (N_21988,N_20964,N_21021);
nor U21989 (N_21989,N_20892,N_20464);
nor U21990 (N_21990,N_21008,N_20431);
nor U21991 (N_21991,N_21258,N_20934);
nor U21992 (N_21992,N_20485,N_20461);
and U21993 (N_21993,N_20939,N_21236);
and U21994 (N_21994,N_21377,N_21383);
xor U21995 (N_21995,N_21180,N_21285);
or U21996 (N_21996,N_20918,N_21030);
or U21997 (N_21997,N_20879,N_21157);
xor U21998 (N_21998,N_20915,N_21382);
nand U21999 (N_21999,N_20722,N_20460);
nand U22000 (N_22000,N_21525,N_20444);
xnor U22001 (N_22001,N_20587,N_20675);
xor U22002 (N_22002,N_20716,N_20720);
or U22003 (N_22003,N_20900,N_20520);
or U22004 (N_22004,N_20813,N_21367);
and U22005 (N_22005,N_21590,N_21583);
xnor U22006 (N_22006,N_21392,N_21183);
nor U22007 (N_22007,N_21353,N_20472);
nand U22008 (N_22008,N_20561,N_21267);
xor U22009 (N_22009,N_21504,N_21585);
nor U22010 (N_22010,N_20777,N_21153);
and U22011 (N_22011,N_20577,N_20401);
and U22012 (N_22012,N_20960,N_21565);
xnor U22013 (N_22013,N_21596,N_20933);
nand U22014 (N_22014,N_20857,N_21203);
nor U22015 (N_22015,N_21209,N_20518);
or U22016 (N_22016,N_21427,N_21275);
nand U22017 (N_22017,N_20906,N_20841);
nor U22018 (N_22018,N_21161,N_20646);
and U22019 (N_22019,N_20778,N_20425);
xor U22020 (N_22020,N_21138,N_21050);
xor U22021 (N_22021,N_20672,N_21114);
or U22022 (N_22022,N_21179,N_20790);
or U22023 (N_22023,N_21278,N_20766);
and U22024 (N_22024,N_20795,N_21090);
and U22025 (N_22025,N_20856,N_21260);
nand U22026 (N_22026,N_21131,N_20523);
xnor U22027 (N_22027,N_21520,N_20586);
or U22028 (N_22028,N_21241,N_20533);
and U22029 (N_22029,N_20903,N_21234);
and U22030 (N_22030,N_20488,N_20543);
and U22031 (N_22031,N_21196,N_21455);
and U22032 (N_22032,N_21094,N_20985);
xor U22033 (N_22033,N_21591,N_20514);
and U22034 (N_22034,N_20852,N_20573);
xor U22035 (N_22035,N_20468,N_20803);
or U22036 (N_22036,N_21498,N_20655);
nor U22037 (N_22037,N_21074,N_21376);
nor U22038 (N_22038,N_21182,N_21221);
nand U22039 (N_22039,N_21549,N_20555);
and U22040 (N_22040,N_20487,N_21404);
or U22041 (N_22041,N_21165,N_21371);
or U22042 (N_22042,N_20552,N_21111);
xnor U22043 (N_22043,N_20692,N_20426);
and U22044 (N_22044,N_20902,N_20788);
nand U22045 (N_22045,N_21466,N_20890);
and U22046 (N_22046,N_20659,N_20832);
nor U22047 (N_22047,N_21249,N_20632);
xnor U22048 (N_22048,N_20418,N_21092);
xor U22049 (N_22049,N_20709,N_21536);
or U22050 (N_22050,N_21502,N_20491);
or U22051 (N_22051,N_21541,N_20851);
nor U22052 (N_22052,N_20769,N_21355);
nand U22053 (N_22053,N_20963,N_21087);
or U22054 (N_22054,N_21233,N_21044);
nand U22055 (N_22055,N_20496,N_20421);
or U22056 (N_22056,N_20805,N_21586);
nand U22057 (N_22057,N_20845,N_20433);
xor U22058 (N_22058,N_20968,N_20837);
and U22059 (N_22059,N_20479,N_21497);
or U22060 (N_22060,N_20977,N_21243);
or U22061 (N_22061,N_20567,N_20482);
and U22062 (N_22062,N_21108,N_21442);
xnor U22063 (N_22063,N_21079,N_20568);
and U22064 (N_22064,N_20483,N_21240);
or U22065 (N_22065,N_20565,N_21078);
nand U22066 (N_22066,N_20936,N_20639);
or U22067 (N_22067,N_20607,N_21557);
xnor U22068 (N_22068,N_20954,N_20883);
and U22069 (N_22069,N_20596,N_20927);
nand U22070 (N_22070,N_21357,N_20947);
nor U22071 (N_22071,N_21579,N_21307);
nor U22072 (N_22072,N_21167,N_21580);
and U22073 (N_22073,N_21588,N_21037);
nand U22074 (N_22074,N_21364,N_21120);
and U22075 (N_22075,N_20726,N_21324);
and U22076 (N_22076,N_20635,N_20836);
nor U22077 (N_22077,N_21177,N_20981);
nor U22078 (N_22078,N_21422,N_20950);
nor U22079 (N_22079,N_21571,N_20924);
nand U22080 (N_22080,N_21581,N_21584);
and U22081 (N_22081,N_20455,N_21325);
or U22082 (N_22082,N_21265,N_21135);
and U22083 (N_22083,N_21564,N_21333);
or U22084 (N_22084,N_20731,N_21042);
nand U22085 (N_22085,N_20962,N_21073);
nand U22086 (N_22086,N_20693,N_20553);
nand U22087 (N_22087,N_20986,N_20889);
nand U22088 (N_22088,N_21478,N_21005);
and U22089 (N_22089,N_20600,N_21064);
or U22090 (N_22090,N_21359,N_21429);
or U22091 (N_22091,N_20770,N_20945);
and U22092 (N_22092,N_21036,N_21378);
and U22093 (N_22093,N_21479,N_21489);
nor U22094 (N_22094,N_20701,N_21365);
and U22095 (N_22095,N_21033,N_20816);
nand U22096 (N_22096,N_20490,N_20991);
nor U22097 (N_22097,N_21099,N_20840);
nor U22098 (N_22098,N_20569,N_20911);
and U22099 (N_22099,N_21027,N_21451);
and U22100 (N_22100,N_21288,N_21049);
and U22101 (N_22101,N_20511,N_21546);
nor U22102 (N_22102,N_20966,N_20746);
or U22103 (N_22103,N_21136,N_21522);
or U22104 (N_22104,N_20528,N_20648);
xor U22105 (N_22105,N_21419,N_20987);
nor U22106 (N_22106,N_20534,N_21428);
nand U22107 (N_22107,N_20530,N_20914);
xnor U22108 (N_22108,N_20821,N_21085);
nand U22109 (N_22109,N_21443,N_21456);
xnor U22110 (N_22110,N_20719,N_21080);
nor U22111 (N_22111,N_21420,N_21261);
xnor U22112 (N_22112,N_20958,N_21002);
xnor U22113 (N_22113,N_21287,N_20538);
nor U22114 (N_22114,N_21093,N_20972);
nor U22115 (N_22115,N_20747,N_21337);
nand U22116 (N_22116,N_20598,N_21013);
and U22117 (N_22117,N_20638,N_21188);
and U22118 (N_22118,N_21539,N_21521);
xor U22119 (N_22119,N_20768,N_21163);
nor U22120 (N_22120,N_20923,N_20910);
and U22121 (N_22121,N_21380,N_21390);
xnor U22122 (N_22122,N_20437,N_20631);
nor U22123 (N_22123,N_20995,N_20894);
xnor U22124 (N_22124,N_21370,N_20793);
nor U22125 (N_22125,N_20647,N_21343);
and U22126 (N_22126,N_20610,N_20997);
and U22127 (N_22127,N_20617,N_21414);
or U22128 (N_22128,N_21356,N_21393);
nor U22129 (N_22129,N_20715,N_21190);
nor U22130 (N_22130,N_20789,N_21315);
xor U22131 (N_22131,N_20980,N_21146);
xor U22132 (N_22132,N_20755,N_20705);
and U22133 (N_22133,N_20427,N_21587);
nand U22134 (N_22134,N_21072,N_21496);
and U22135 (N_22135,N_20867,N_20781);
xor U22136 (N_22136,N_21349,N_21239);
or U22137 (N_22137,N_20785,N_20948);
xnor U22138 (N_22138,N_20946,N_20645);
or U22139 (N_22139,N_20486,N_20855);
nand U22140 (N_22140,N_21127,N_21395);
or U22141 (N_22141,N_20754,N_20570);
nor U22142 (N_22142,N_20403,N_20753);
nor U22143 (N_22143,N_20749,N_21306);
xnor U22144 (N_22144,N_20859,N_20445);
nand U22145 (N_22145,N_21454,N_21255);
nand U22146 (N_22146,N_21515,N_21098);
xnor U22147 (N_22147,N_20619,N_20702);
or U22148 (N_22148,N_20707,N_21407);
xnor U22149 (N_22149,N_21366,N_21056);
xnor U22150 (N_22150,N_20477,N_21026);
or U22151 (N_22151,N_21441,N_20818);
nand U22152 (N_22152,N_21568,N_21484);
nor U22153 (N_22153,N_20898,N_20434);
nor U22154 (N_22154,N_21054,N_20959);
or U22155 (N_22155,N_21113,N_20724);
nor U22156 (N_22156,N_20896,N_20424);
or U22157 (N_22157,N_21439,N_21297);
nand U22158 (N_22158,N_20881,N_20912);
or U22159 (N_22159,N_20717,N_21309);
and U22160 (N_22160,N_20653,N_21535);
xnor U22161 (N_22161,N_21125,N_20508);
and U22162 (N_22162,N_20697,N_20787);
nor U22163 (N_22163,N_20764,N_20563);
nor U22164 (N_22164,N_21578,N_21252);
xnor U22165 (N_22165,N_21445,N_20786);
or U22166 (N_22166,N_20611,N_21342);
and U22167 (N_22167,N_21112,N_20683);
nand U22168 (N_22168,N_21352,N_21214);
nor U22169 (N_22169,N_21154,N_20690);
and U22170 (N_22170,N_21387,N_20876);
nand U22171 (N_22171,N_20510,N_20498);
xnor U22172 (N_22172,N_21500,N_21083);
nor U22173 (N_22173,N_21156,N_21452);
or U22174 (N_22174,N_20677,N_20804);
and U22175 (N_22175,N_21162,N_21597);
or U22176 (N_22176,N_20636,N_21471);
or U22177 (N_22177,N_20422,N_21433);
or U22178 (N_22178,N_21077,N_21268);
and U22179 (N_22179,N_20819,N_20478);
nor U22180 (N_22180,N_21109,N_20603);
and U22181 (N_22181,N_20878,N_21480);
nor U22182 (N_22182,N_20812,N_21476);
xor U22183 (N_22183,N_21105,N_21123);
nor U22184 (N_22184,N_20467,N_20831);
nand U22185 (N_22185,N_21459,N_21426);
xor U22186 (N_22186,N_20525,N_20967);
and U22187 (N_22187,N_21043,N_21084);
xor U22188 (N_22188,N_20826,N_20864);
and U22189 (N_22189,N_21344,N_20469);
and U22190 (N_22190,N_20899,N_20412);
xor U22191 (N_22191,N_20801,N_20557);
nor U22192 (N_22192,N_21384,N_21024);
nor U22193 (N_22193,N_20429,N_20623);
nor U22194 (N_22194,N_21321,N_21311);
or U22195 (N_22195,N_21150,N_21425);
nor U22196 (N_22196,N_21302,N_20447);
or U22197 (N_22197,N_21589,N_21340);
and U22198 (N_22198,N_21438,N_20811);
nor U22199 (N_22199,N_20806,N_21141);
and U22200 (N_22200,N_21253,N_20437);
nand U22201 (N_22201,N_21150,N_20595);
and U22202 (N_22202,N_21492,N_20616);
or U22203 (N_22203,N_20812,N_21138);
and U22204 (N_22204,N_20504,N_20465);
xnor U22205 (N_22205,N_20774,N_21430);
or U22206 (N_22206,N_20444,N_20703);
and U22207 (N_22207,N_21254,N_21524);
nand U22208 (N_22208,N_20460,N_20708);
xor U22209 (N_22209,N_20507,N_21461);
nand U22210 (N_22210,N_20540,N_21026);
xor U22211 (N_22211,N_20889,N_20662);
nand U22212 (N_22212,N_21104,N_20706);
xnor U22213 (N_22213,N_20654,N_20665);
and U22214 (N_22214,N_20866,N_20869);
and U22215 (N_22215,N_21457,N_20936);
or U22216 (N_22216,N_21284,N_20603);
and U22217 (N_22217,N_20909,N_21252);
and U22218 (N_22218,N_20695,N_21163);
and U22219 (N_22219,N_20727,N_21037);
and U22220 (N_22220,N_21264,N_20871);
and U22221 (N_22221,N_20818,N_20894);
nand U22222 (N_22222,N_21112,N_20786);
nor U22223 (N_22223,N_20730,N_21308);
nand U22224 (N_22224,N_21336,N_20954);
and U22225 (N_22225,N_20758,N_20865);
xor U22226 (N_22226,N_20574,N_20822);
nor U22227 (N_22227,N_21228,N_20895);
or U22228 (N_22228,N_20519,N_20763);
nor U22229 (N_22229,N_21382,N_21085);
nand U22230 (N_22230,N_20935,N_21015);
nor U22231 (N_22231,N_20886,N_21357);
nand U22232 (N_22232,N_20477,N_20946);
or U22233 (N_22233,N_20539,N_20449);
nand U22234 (N_22234,N_20840,N_21590);
and U22235 (N_22235,N_20468,N_20569);
and U22236 (N_22236,N_21270,N_21080);
or U22237 (N_22237,N_20940,N_20821);
nand U22238 (N_22238,N_21015,N_20828);
xor U22239 (N_22239,N_20694,N_21162);
nor U22240 (N_22240,N_21021,N_20414);
xor U22241 (N_22241,N_20599,N_20570);
and U22242 (N_22242,N_20532,N_20822);
nand U22243 (N_22243,N_21595,N_21579);
nor U22244 (N_22244,N_20450,N_20465);
or U22245 (N_22245,N_20878,N_20492);
nor U22246 (N_22246,N_21223,N_20573);
nor U22247 (N_22247,N_21201,N_21108);
or U22248 (N_22248,N_20811,N_21350);
and U22249 (N_22249,N_20669,N_21131);
or U22250 (N_22250,N_20746,N_20967);
xnor U22251 (N_22251,N_20492,N_21059);
nor U22252 (N_22252,N_20689,N_21054);
nand U22253 (N_22253,N_21063,N_21532);
xor U22254 (N_22254,N_21227,N_20422);
or U22255 (N_22255,N_21447,N_20533);
nor U22256 (N_22256,N_20730,N_21139);
or U22257 (N_22257,N_21596,N_20716);
nand U22258 (N_22258,N_21306,N_20856);
and U22259 (N_22259,N_20906,N_20759);
nand U22260 (N_22260,N_20535,N_20959);
or U22261 (N_22261,N_21377,N_21187);
and U22262 (N_22262,N_20500,N_20672);
nor U22263 (N_22263,N_21523,N_20869);
nand U22264 (N_22264,N_21581,N_20711);
nor U22265 (N_22265,N_21367,N_20549);
or U22266 (N_22266,N_20843,N_20850);
nand U22267 (N_22267,N_20467,N_20828);
nor U22268 (N_22268,N_20567,N_21189);
xnor U22269 (N_22269,N_21484,N_20449);
xnor U22270 (N_22270,N_21449,N_20898);
or U22271 (N_22271,N_21035,N_21160);
xnor U22272 (N_22272,N_21043,N_20771);
nand U22273 (N_22273,N_21522,N_21546);
nor U22274 (N_22274,N_20880,N_21367);
or U22275 (N_22275,N_21297,N_20469);
or U22276 (N_22276,N_20794,N_20793);
nand U22277 (N_22277,N_21292,N_21504);
xor U22278 (N_22278,N_20797,N_20967);
and U22279 (N_22279,N_20781,N_20423);
nor U22280 (N_22280,N_20540,N_20927);
nand U22281 (N_22281,N_21041,N_20952);
xor U22282 (N_22282,N_21345,N_20780);
nand U22283 (N_22283,N_21089,N_20627);
or U22284 (N_22284,N_21292,N_20929);
xor U22285 (N_22285,N_21248,N_20504);
nor U22286 (N_22286,N_20437,N_20895);
and U22287 (N_22287,N_21073,N_21134);
nand U22288 (N_22288,N_20823,N_20445);
and U22289 (N_22289,N_21474,N_21463);
nor U22290 (N_22290,N_20602,N_21142);
and U22291 (N_22291,N_21489,N_20732);
nand U22292 (N_22292,N_20767,N_20735);
or U22293 (N_22293,N_21501,N_21112);
and U22294 (N_22294,N_21281,N_20551);
xnor U22295 (N_22295,N_21334,N_21516);
nand U22296 (N_22296,N_21261,N_20948);
xnor U22297 (N_22297,N_20801,N_21596);
and U22298 (N_22298,N_21063,N_21190);
and U22299 (N_22299,N_21496,N_20871);
and U22300 (N_22300,N_20733,N_21484);
nand U22301 (N_22301,N_21285,N_20643);
xnor U22302 (N_22302,N_20716,N_21587);
and U22303 (N_22303,N_20647,N_20697);
or U22304 (N_22304,N_20666,N_21585);
or U22305 (N_22305,N_21290,N_20690);
nand U22306 (N_22306,N_21086,N_20789);
or U22307 (N_22307,N_20661,N_21437);
and U22308 (N_22308,N_20487,N_20791);
nor U22309 (N_22309,N_20516,N_20914);
nor U22310 (N_22310,N_20957,N_20780);
xor U22311 (N_22311,N_21413,N_20768);
nor U22312 (N_22312,N_21505,N_20605);
xnor U22313 (N_22313,N_21044,N_21273);
nor U22314 (N_22314,N_20702,N_20507);
nor U22315 (N_22315,N_20816,N_20832);
nor U22316 (N_22316,N_21129,N_21285);
and U22317 (N_22317,N_21015,N_20614);
xnor U22318 (N_22318,N_20454,N_20411);
nand U22319 (N_22319,N_20512,N_20993);
xor U22320 (N_22320,N_21436,N_21089);
nand U22321 (N_22321,N_20706,N_21472);
nand U22322 (N_22322,N_21138,N_20698);
xnor U22323 (N_22323,N_21036,N_20978);
xnor U22324 (N_22324,N_21524,N_21412);
nor U22325 (N_22325,N_21479,N_20475);
nand U22326 (N_22326,N_20563,N_20925);
and U22327 (N_22327,N_21513,N_21311);
xor U22328 (N_22328,N_20783,N_20793);
or U22329 (N_22329,N_20508,N_21523);
nand U22330 (N_22330,N_21314,N_21350);
nand U22331 (N_22331,N_21402,N_20843);
nand U22332 (N_22332,N_21549,N_21106);
xor U22333 (N_22333,N_21419,N_21342);
xnor U22334 (N_22334,N_20757,N_20775);
nand U22335 (N_22335,N_21386,N_21312);
or U22336 (N_22336,N_20902,N_20876);
or U22337 (N_22337,N_20413,N_21140);
xnor U22338 (N_22338,N_21006,N_21249);
and U22339 (N_22339,N_21558,N_20469);
xnor U22340 (N_22340,N_20576,N_20799);
and U22341 (N_22341,N_21432,N_21148);
xor U22342 (N_22342,N_20877,N_20500);
nand U22343 (N_22343,N_21235,N_20788);
nand U22344 (N_22344,N_20768,N_20820);
nand U22345 (N_22345,N_20446,N_20701);
nand U22346 (N_22346,N_21477,N_20653);
or U22347 (N_22347,N_20728,N_21242);
nand U22348 (N_22348,N_21476,N_20845);
or U22349 (N_22349,N_21318,N_20935);
or U22350 (N_22350,N_21364,N_21076);
or U22351 (N_22351,N_21352,N_21190);
nor U22352 (N_22352,N_20558,N_21328);
xnor U22353 (N_22353,N_21333,N_20542);
or U22354 (N_22354,N_21260,N_21041);
nand U22355 (N_22355,N_20765,N_21340);
nor U22356 (N_22356,N_20401,N_20800);
or U22357 (N_22357,N_21560,N_20639);
xnor U22358 (N_22358,N_21450,N_21059);
or U22359 (N_22359,N_21505,N_21244);
xnor U22360 (N_22360,N_21514,N_20442);
or U22361 (N_22361,N_20856,N_21104);
or U22362 (N_22362,N_21453,N_20927);
or U22363 (N_22363,N_20680,N_21271);
xnor U22364 (N_22364,N_21255,N_20439);
or U22365 (N_22365,N_21439,N_21219);
xnor U22366 (N_22366,N_21098,N_21317);
xnor U22367 (N_22367,N_21138,N_20826);
nor U22368 (N_22368,N_21323,N_20664);
nor U22369 (N_22369,N_21297,N_21446);
xnor U22370 (N_22370,N_21174,N_21149);
nand U22371 (N_22371,N_20943,N_20496);
and U22372 (N_22372,N_21364,N_20449);
and U22373 (N_22373,N_20948,N_20771);
xor U22374 (N_22374,N_21572,N_20688);
nor U22375 (N_22375,N_21402,N_20831);
and U22376 (N_22376,N_21563,N_20852);
and U22377 (N_22377,N_20726,N_20909);
nand U22378 (N_22378,N_20645,N_20860);
xnor U22379 (N_22379,N_21589,N_20980);
xor U22380 (N_22380,N_20447,N_20943);
nor U22381 (N_22381,N_21234,N_21419);
nand U22382 (N_22382,N_20523,N_21271);
or U22383 (N_22383,N_20634,N_21167);
and U22384 (N_22384,N_20536,N_21491);
and U22385 (N_22385,N_21590,N_21535);
or U22386 (N_22386,N_20681,N_21233);
and U22387 (N_22387,N_20661,N_21452);
xnor U22388 (N_22388,N_21084,N_21579);
nand U22389 (N_22389,N_21435,N_20797);
or U22390 (N_22390,N_21021,N_20987);
or U22391 (N_22391,N_20833,N_20581);
and U22392 (N_22392,N_21483,N_21185);
or U22393 (N_22393,N_20648,N_20894);
nor U22394 (N_22394,N_21524,N_21115);
or U22395 (N_22395,N_20416,N_21468);
or U22396 (N_22396,N_21016,N_20799);
or U22397 (N_22397,N_20769,N_20580);
nand U22398 (N_22398,N_20762,N_20725);
nor U22399 (N_22399,N_21561,N_21504);
nor U22400 (N_22400,N_20852,N_21478);
nor U22401 (N_22401,N_20434,N_21504);
nand U22402 (N_22402,N_21450,N_21023);
nor U22403 (N_22403,N_20762,N_20482);
nor U22404 (N_22404,N_21035,N_21579);
nand U22405 (N_22405,N_21077,N_20989);
or U22406 (N_22406,N_21495,N_21064);
xnor U22407 (N_22407,N_20762,N_21400);
and U22408 (N_22408,N_20549,N_20627);
or U22409 (N_22409,N_20880,N_20425);
nand U22410 (N_22410,N_20585,N_20429);
nor U22411 (N_22411,N_21094,N_20882);
and U22412 (N_22412,N_21082,N_20830);
or U22413 (N_22413,N_21069,N_20878);
nor U22414 (N_22414,N_20526,N_21277);
nand U22415 (N_22415,N_20425,N_21580);
nand U22416 (N_22416,N_21036,N_21158);
nor U22417 (N_22417,N_21128,N_21083);
xor U22418 (N_22418,N_20577,N_20409);
or U22419 (N_22419,N_20599,N_21027);
and U22420 (N_22420,N_21239,N_21192);
nand U22421 (N_22421,N_20995,N_21421);
xor U22422 (N_22422,N_21422,N_21144);
xor U22423 (N_22423,N_20774,N_21551);
nand U22424 (N_22424,N_20790,N_20414);
nand U22425 (N_22425,N_21257,N_21118);
nor U22426 (N_22426,N_20554,N_20494);
xnor U22427 (N_22427,N_21318,N_20517);
nand U22428 (N_22428,N_20817,N_20660);
nand U22429 (N_22429,N_21482,N_20785);
nand U22430 (N_22430,N_21395,N_21463);
or U22431 (N_22431,N_21003,N_21391);
xor U22432 (N_22432,N_21150,N_21008);
or U22433 (N_22433,N_20896,N_20894);
nor U22434 (N_22434,N_21443,N_21032);
or U22435 (N_22435,N_21385,N_21511);
nor U22436 (N_22436,N_20998,N_20503);
or U22437 (N_22437,N_21237,N_20850);
nor U22438 (N_22438,N_21386,N_20693);
xnor U22439 (N_22439,N_21521,N_20658);
nand U22440 (N_22440,N_20505,N_21367);
or U22441 (N_22441,N_20761,N_21130);
or U22442 (N_22442,N_20677,N_20912);
or U22443 (N_22443,N_21445,N_21510);
or U22444 (N_22444,N_21508,N_20401);
and U22445 (N_22445,N_21027,N_20411);
and U22446 (N_22446,N_21031,N_21037);
nor U22447 (N_22447,N_21508,N_20748);
or U22448 (N_22448,N_21074,N_20579);
or U22449 (N_22449,N_21483,N_21226);
xnor U22450 (N_22450,N_20735,N_21420);
or U22451 (N_22451,N_20509,N_20608);
and U22452 (N_22452,N_20529,N_20736);
xor U22453 (N_22453,N_21440,N_21274);
and U22454 (N_22454,N_21176,N_20613);
nor U22455 (N_22455,N_21062,N_21502);
nand U22456 (N_22456,N_20857,N_21556);
or U22457 (N_22457,N_20827,N_20866);
nor U22458 (N_22458,N_20874,N_21521);
xnor U22459 (N_22459,N_21172,N_20930);
or U22460 (N_22460,N_20477,N_20626);
or U22461 (N_22461,N_21270,N_21239);
xor U22462 (N_22462,N_21263,N_21247);
xnor U22463 (N_22463,N_21311,N_21518);
nor U22464 (N_22464,N_20533,N_21100);
and U22465 (N_22465,N_20517,N_21587);
nand U22466 (N_22466,N_21030,N_21014);
xor U22467 (N_22467,N_21403,N_20888);
and U22468 (N_22468,N_20741,N_20962);
nor U22469 (N_22469,N_20806,N_20884);
and U22470 (N_22470,N_21456,N_21067);
and U22471 (N_22471,N_21267,N_21016);
and U22472 (N_22472,N_20808,N_20716);
or U22473 (N_22473,N_20649,N_20984);
nand U22474 (N_22474,N_20558,N_20451);
nand U22475 (N_22475,N_20508,N_20850);
nor U22476 (N_22476,N_21517,N_21170);
and U22477 (N_22477,N_20819,N_20550);
nor U22478 (N_22478,N_21249,N_21026);
nand U22479 (N_22479,N_21387,N_20991);
and U22480 (N_22480,N_21241,N_21323);
and U22481 (N_22481,N_20941,N_21217);
nor U22482 (N_22482,N_20552,N_21179);
nor U22483 (N_22483,N_21458,N_20630);
or U22484 (N_22484,N_20991,N_20844);
nand U22485 (N_22485,N_20400,N_21574);
or U22486 (N_22486,N_21506,N_21024);
nor U22487 (N_22487,N_21144,N_21221);
and U22488 (N_22488,N_20937,N_20992);
and U22489 (N_22489,N_20703,N_21281);
xnor U22490 (N_22490,N_20947,N_20638);
and U22491 (N_22491,N_21209,N_20874);
nor U22492 (N_22492,N_21190,N_21384);
nand U22493 (N_22493,N_21166,N_20492);
nand U22494 (N_22494,N_20708,N_20570);
and U22495 (N_22495,N_21299,N_20834);
nor U22496 (N_22496,N_21510,N_21528);
nor U22497 (N_22497,N_20919,N_21540);
nand U22498 (N_22498,N_20923,N_20721);
or U22499 (N_22499,N_21504,N_20897);
or U22500 (N_22500,N_20939,N_20427);
nor U22501 (N_22501,N_20901,N_20646);
xnor U22502 (N_22502,N_21151,N_21091);
nor U22503 (N_22503,N_21516,N_20744);
xor U22504 (N_22504,N_20967,N_20580);
and U22505 (N_22505,N_21331,N_20845);
and U22506 (N_22506,N_20511,N_21023);
nor U22507 (N_22507,N_21343,N_21010);
nor U22508 (N_22508,N_20662,N_21245);
nor U22509 (N_22509,N_20653,N_21101);
and U22510 (N_22510,N_21269,N_20863);
xor U22511 (N_22511,N_21289,N_21133);
or U22512 (N_22512,N_20948,N_20827);
and U22513 (N_22513,N_20623,N_20511);
xor U22514 (N_22514,N_21371,N_21014);
or U22515 (N_22515,N_21114,N_20558);
or U22516 (N_22516,N_20749,N_20910);
nand U22517 (N_22517,N_20715,N_21100);
nand U22518 (N_22518,N_21368,N_20627);
nor U22519 (N_22519,N_20602,N_20743);
or U22520 (N_22520,N_21453,N_21167);
nor U22521 (N_22521,N_20443,N_20733);
or U22522 (N_22522,N_20713,N_21173);
nor U22523 (N_22523,N_21191,N_21301);
or U22524 (N_22524,N_20830,N_21028);
nand U22525 (N_22525,N_20703,N_20454);
nand U22526 (N_22526,N_21442,N_20516);
nor U22527 (N_22527,N_20792,N_20495);
and U22528 (N_22528,N_20820,N_20418);
and U22529 (N_22529,N_20521,N_21518);
xor U22530 (N_22530,N_20794,N_21059);
and U22531 (N_22531,N_20648,N_21267);
or U22532 (N_22532,N_21251,N_20989);
xnor U22533 (N_22533,N_20615,N_20451);
or U22534 (N_22534,N_20650,N_21227);
nor U22535 (N_22535,N_20544,N_21073);
and U22536 (N_22536,N_20503,N_20669);
and U22537 (N_22537,N_21291,N_20447);
nand U22538 (N_22538,N_20788,N_20540);
and U22539 (N_22539,N_21239,N_20954);
or U22540 (N_22540,N_21162,N_20860);
and U22541 (N_22541,N_21438,N_20737);
xor U22542 (N_22542,N_21056,N_20711);
or U22543 (N_22543,N_20421,N_21278);
nand U22544 (N_22544,N_21283,N_20705);
xor U22545 (N_22545,N_21174,N_21212);
nor U22546 (N_22546,N_21423,N_20875);
and U22547 (N_22547,N_20958,N_20652);
or U22548 (N_22548,N_21590,N_21255);
and U22549 (N_22549,N_20878,N_20553);
or U22550 (N_22550,N_20840,N_21054);
and U22551 (N_22551,N_20601,N_20546);
and U22552 (N_22552,N_20728,N_21021);
and U22553 (N_22553,N_20556,N_21388);
or U22554 (N_22554,N_21548,N_20415);
and U22555 (N_22555,N_21411,N_21567);
or U22556 (N_22556,N_20400,N_21419);
xor U22557 (N_22557,N_21511,N_20495);
and U22558 (N_22558,N_21126,N_21170);
nand U22559 (N_22559,N_20987,N_21369);
and U22560 (N_22560,N_20917,N_20763);
xnor U22561 (N_22561,N_21153,N_21104);
or U22562 (N_22562,N_21254,N_20624);
nor U22563 (N_22563,N_20900,N_21477);
nor U22564 (N_22564,N_20645,N_20859);
nand U22565 (N_22565,N_20527,N_20462);
nand U22566 (N_22566,N_21399,N_21369);
or U22567 (N_22567,N_21380,N_20434);
or U22568 (N_22568,N_20932,N_20540);
or U22569 (N_22569,N_21076,N_21214);
and U22570 (N_22570,N_20430,N_20437);
nand U22571 (N_22571,N_20446,N_21591);
nand U22572 (N_22572,N_21443,N_20590);
nand U22573 (N_22573,N_20725,N_20555);
and U22574 (N_22574,N_20786,N_21053);
and U22575 (N_22575,N_20609,N_21367);
xnor U22576 (N_22576,N_20887,N_20834);
nor U22577 (N_22577,N_21353,N_20703);
and U22578 (N_22578,N_20540,N_21447);
nor U22579 (N_22579,N_21289,N_20665);
xnor U22580 (N_22580,N_21313,N_20609);
nand U22581 (N_22581,N_20454,N_20842);
or U22582 (N_22582,N_21183,N_21063);
nor U22583 (N_22583,N_21442,N_20413);
or U22584 (N_22584,N_20882,N_21229);
and U22585 (N_22585,N_21564,N_20858);
nor U22586 (N_22586,N_21287,N_21142);
nand U22587 (N_22587,N_21075,N_20474);
nand U22588 (N_22588,N_21147,N_20841);
xor U22589 (N_22589,N_21102,N_21391);
nand U22590 (N_22590,N_21134,N_21360);
nand U22591 (N_22591,N_20539,N_21165);
nand U22592 (N_22592,N_21318,N_21192);
xnor U22593 (N_22593,N_20571,N_21145);
nor U22594 (N_22594,N_21505,N_21021);
xnor U22595 (N_22595,N_20470,N_20757);
and U22596 (N_22596,N_21317,N_20969);
nor U22597 (N_22597,N_21227,N_21020);
or U22598 (N_22598,N_21388,N_20664);
xor U22599 (N_22599,N_21492,N_20486);
nand U22600 (N_22600,N_20596,N_20749);
nand U22601 (N_22601,N_21263,N_20662);
or U22602 (N_22602,N_21085,N_20853);
or U22603 (N_22603,N_21578,N_20759);
and U22604 (N_22604,N_21589,N_20951);
or U22605 (N_22605,N_21424,N_20751);
nand U22606 (N_22606,N_21250,N_21217);
nor U22607 (N_22607,N_20954,N_20637);
xnor U22608 (N_22608,N_20977,N_20431);
xnor U22609 (N_22609,N_20526,N_21034);
nand U22610 (N_22610,N_20730,N_21239);
nand U22611 (N_22611,N_21176,N_21375);
xor U22612 (N_22612,N_20798,N_20666);
and U22613 (N_22613,N_21201,N_21501);
nand U22614 (N_22614,N_20925,N_20467);
nor U22615 (N_22615,N_21461,N_21320);
or U22616 (N_22616,N_21176,N_21488);
xnor U22617 (N_22617,N_21121,N_20993);
nor U22618 (N_22618,N_21027,N_20623);
and U22619 (N_22619,N_20794,N_21300);
and U22620 (N_22620,N_21487,N_20462);
or U22621 (N_22621,N_21149,N_20572);
and U22622 (N_22622,N_20660,N_20951);
or U22623 (N_22623,N_20626,N_20761);
xor U22624 (N_22624,N_21414,N_20903);
and U22625 (N_22625,N_20537,N_20474);
or U22626 (N_22626,N_20480,N_20950);
and U22627 (N_22627,N_21387,N_20586);
nor U22628 (N_22628,N_20726,N_20718);
nor U22629 (N_22629,N_21077,N_20404);
nand U22630 (N_22630,N_20672,N_21038);
or U22631 (N_22631,N_20755,N_20734);
nand U22632 (N_22632,N_21169,N_20810);
nand U22633 (N_22633,N_21039,N_20874);
and U22634 (N_22634,N_20913,N_21037);
nor U22635 (N_22635,N_21299,N_21389);
nand U22636 (N_22636,N_21595,N_20545);
xnor U22637 (N_22637,N_21278,N_20739);
or U22638 (N_22638,N_20450,N_20539);
and U22639 (N_22639,N_20411,N_21483);
nand U22640 (N_22640,N_21204,N_20939);
nand U22641 (N_22641,N_21312,N_21522);
and U22642 (N_22642,N_20913,N_20436);
and U22643 (N_22643,N_20981,N_21137);
and U22644 (N_22644,N_20576,N_20574);
xor U22645 (N_22645,N_21364,N_20811);
nand U22646 (N_22646,N_20861,N_20903);
and U22647 (N_22647,N_21529,N_21361);
and U22648 (N_22648,N_21087,N_21351);
nor U22649 (N_22649,N_21023,N_20594);
nor U22650 (N_22650,N_20859,N_21547);
nand U22651 (N_22651,N_21027,N_21022);
or U22652 (N_22652,N_20625,N_21276);
xor U22653 (N_22653,N_20959,N_20506);
nor U22654 (N_22654,N_21195,N_20611);
xnor U22655 (N_22655,N_20938,N_20659);
nor U22656 (N_22656,N_21459,N_21391);
or U22657 (N_22657,N_21282,N_20430);
nor U22658 (N_22658,N_21038,N_20782);
or U22659 (N_22659,N_21540,N_21479);
nor U22660 (N_22660,N_20702,N_20889);
and U22661 (N_22661,N_20605,N_21347);
and U22662 (N_22662,N_20847,N_21457);
xor U22663 (N_22663,N_21354,N_21048);
or U22664 (N_22664,N_21437,N_20613);
nand U22665 (N_22665,N_20880,N_21214);
and U22666 (N_22666,N_20635,N_21579);
xnor U22667 (N_22667,N_20554,N_20743);
nand U22668 (N_22668,N_20700,N_21509);
nor U22669 (N_22669,N_21511,N_20895);
and U22670 (N_22670,N_21561,N_20689);
or U22671 (N_22671,N_21264,N_20564);
or U22672 (N_22672,N_21195,N_21572);
xnor U22673 (N_22673,N_20468,N_21503);
or U22674 (N_22674,N_21313,N_21276);
xor U22675 (N_22675,N_21268,N_21238);
or U22676 (N_22676,N_21563,N_21279);
or U22677 (N_22677,N_20645,N_21129);
xnor U22678 (N_22678,N_20416,N_21241);
xor U22679 (N_22679,N_21119,N_20516);
xor U22680 (N_22680,N_21287,N_21182);
or U22681 (N_22681,N_20813,N_21446);
and U22682 (N_22682,N_20803,N_21577);
or U22683 (N_22683,N_21290,N_20475);
xor U22684 (N_22684,N_20648,N_20770);
nand U22685 (N_22685,N_20465,N_20828);
and U22686 (N_22686,N_21449,N_20789);
nor U22687 (N_22687,N_20893,N_21384);
or U22688 (N_22688,N_21254,N_21028);
xor U22689 (N_22689,N_20819,N_20497);
nand U22690 (N_22690,N_20991,N_21395);
xnor U22691 (N_22691,N_21327,N_20606);
xor U22692 (N_22692,N_21184,N_21524);
and U22693 (N_22693,N_20470,N_21189);
nand U22694 (N_22694,N_20902,N_20508);
nor U22695 (N_22695,N_21392,N_21346);
and U22696 (N_22696,N_21013,N_21432);
nand U22697 (N_22697,N_21052,N_21186);
or U22698 (N_22698,N_20935,N_21064);
nand U22699 (N_22699,N_20677,N_21537);
xor U22700 (N_22700,N_20706,N_21229);
nand U22701 (N_22701,N_21379,N_20638);
nand U22702 (N_22702,N_20888,N_20879);
and U22703 (N_22703,N_20575,N_20416);
xor U22704 (N_22704,N_20516,N_21224);
xor U22705 (N_22705,N_21576,N_21586);
and U22706 (N_22706,N_21428,N_20872);
xor U22707 (N_22707,N_20985,N_20624);
and U22708 (N_22708,N_21107,N_20873);
xnor U22709 (N_22709,N_21537,N_20506);
xnor U22710 (N_22710,N_21462,N_21233);
xor U22711 (N_22711,N_21282,N_21229);
and U22712 (N_22712,N_20620,N_20834);
and U22713 (N_22713,N_21306,N_20716);
nor U22714 (N_22714,N_21072,N_20495);
nor U22715 (N_22715,N_21415,N_21591);
nand U22716 (N_22716,N_20574,N_20859);
or U22717 (N_22717,N_21190,N_21134);
and U22718 (N_22718,N_21218,N_20807);
or U22719 (N_22719,N_21347,N_21520);
nand U22720 (N_22720,N_20500,N_20605);
nand U22721 (N_22721,N_21319,N_20601);
xor U22722 (N_22722,N_21038,N_20475);
nor U22723 (N_22723,N_21419,N_21166);
nand U22724 (N_22724,N_20525,N_21031);
or U22725 (N_22725,N_21526,N_20970);
nand U22726 (N_22726,N_20850,N_20876);
xor U22727 (N_22727,N_21082,N_20493);
xnor U22728 (N_22728,N_20561,N_21467);
nor U22729 (N_22729,N_21236,N_21570);
nand U22730 (N_22730,N_21194,N_21577);
nor U22731 (N_22731,N_20951,N_21029);
or U22732 (N_22732,N_21097,N_20545);
or U22733 (N_22733,N_20902,N_20402);
nor U22734 (N_22734,N_20596,N_20416);
xor U22735 (N_22735,N_20871,N_21589);
nor U22736 (N_22736,N_20972,N_21125);
nor U22737 (N_22737,N_20841,N_20446);
nor U22738 (N_22738,N_21135,N_20783);
nor U22739 (N_22739,N_20480,N_21594);
and U22740 (N_22740,N_20552,N_20597);
nor U22741 (N_22741,N_20402,N_21024);
xor U22742 (N_22742,N_20696,N_21385);
and U22743 (N_22743,N_21458,N_21390);
and U22744 (N_22744,N_21124,N_21277);
and U22745 (N_22745,N_21530,N_20416);
nand U22746 (N_22746,N_21097,N_20557);
nor U22747 (N_22747,N_20546,N_21480);
or U22748 (N_22748,N_21502,N_20583);
or U22749 (N_22749,N_21373,N_20835);
and U22750 (N_22750,N_20847,N_20703);
nor U22751 (N_22751,N_21312,N_20901);
or U22752 (N_22752,N_20569,N_20679);
and U22753 (N_22753,N_21000,N_20618);
nand U22754 (N_22754,N_21175,N_21363);
nor U22755 (N_22755,N_21450,N_20719);
nand U22756 (N_22756,N_20990,N_20788);
xnor U22757 (N_22757,N_20967,N_20687);
or U22758 (N_22758,N_21112,N_21450);
and U22759 (N_22759,N_21222,N_20615);
nand U22760 (N_22760,N_21137,N_21552);
and U22761 (N_22761,N_20805,N_21345);
nor U22762 (N_22762,N_20435,N_20491);
nor U22763 (N_22763,N_21195,N_20987);
and U22764 (N_22764,N_20779,N_20453);
or U22765 (N_22765,N_20798,N_20717);
or U22766 (N_22766,N_20796,N_21150);
nor U22767 (N_22767,N_21004,N_21240);
and U22768 (N_22768,N_20533,N_21529);
and U22769 (N_22769,N_21464,N_20511);
nand U22770 (N_22770,N_21205,N_21583);
and U22771 (N_22771,N_21481,N_21279);
xor U22772 (N_22772,N_21251,N_20961);
nand U22773 (N_22773,N_20576,N_20817);
or U22774 (N_22774,N_21475,N_20562);
xor U22775 (N_22775,N_20798,N_20441);
and U22776 (N_22776,N_20916,N_21302);
xnor U22777 (N_22777,N_20502,N_21077);
xor U22778 (N_22778,N_21299,N_21095);
nor U22779 (N_22779,N_21280,N_20738);
nor U22780 (N_22780,N_21107,N_21311);
nand U22781 (N_22781,N_20672,N_21253);
and U22782 (N_22782,N_21544,N_21538);
or U22783 (N_22783,N_20550,N_20956);
and U22784 (N_22784,N_20572,N_20990);
nand U22785 (N_22785,N_21431,N_20819);
or U22786 (N_22786,N_20533,N_21176);
and U22787 (N_22787,N_21188,N_20578);
xnor U22788 (N_22788,N_20662,N_21025);
and U22789 (N_22789,N_21297,N_21405);
and U22790 (N_22790,N_20939,N_20416);
or U22791 (N_22791,N_21410,N_20708);
nor U22792 (N_22792,N_21492,N_21371);
and U22793 (N_22793,N_21074,N_20919);
nor U22794 (N_22794,N_20507,N_20844);
nand U22795 (N_22795,N_21539,N_21423);
nor U22796 (N_22796,N_20488,N_20523);
nor U22797 (N_22797,N_21441,N_20477);
and U22798 (N_22798,N_20516,N_20738);
nand U22799 (N_22799,N_20457,N_21590);
or U22800 (N_22800,N_21758,N_22228);
or U22801 (N_22801,N_22100,N_22741);
and U22802 (N_22802,N_21932,N_21750);
nor U22803 (N_22803,N_21687,N_21966);
nand U22804 (N_22804,N_22040,N_22568);
nand U22805 (N_22805,N_22452,N_22639);
and U22806 (N_22806,N_21792,N_22250);
or U22807 (N_22807,N_22764,N_22717);
nand U22808 (N_22808,N_22150,N_21752);
nor U22809 (N_22809,N_22059,N_22345);
nand U22810 (N_22810,N_22265,N_22533);
xor U22811 (N_22811,N_21741,N_21828);
nand U22812 (N_22812,N_22223,N_21835);
nor U22813 (N_22813,N_21808,N_22609);
nand U22814 (N_22814,N_21886,N_22414);
xor U22815 (N_22815,N_22474,N_22726);
or U22816 (N_22816,N_22762,N_21855);
nand U22817 (N_22817,N_21601,N_22161);
or U22818 (N_22818,N_21760,N_22237);
or U22819 (N_22819,N_22053,N_22661);
xor U22820 (N_22820,N_22542,N_22106);
or U22821 (N_22821,N_22417,N_22143);
nor U22822 (N_22822,N_22224,N_22523);
and U22823 (N_22823,N_22623,N_22740);
nor U22824 (N_22824,N_21662,N_21611);
nand U22825 (N_22825,N_21774,N_22373);
nand U22826 (N_22826,N_21685,N_22225);
xor U22827 (N_22827,N_22455,N_21634);
nand U22828 (N_22828,N_21674,N_22317);
and U22829 (N_22829,N_21749,N_22774);
or U22830 (N_22830,N_22030,N_21747);
or U22831 (N_22831,N_22567,N_22546);
and U22832 (N_22832,N_21751,N_22102);
nor U22833 (N_22833,N_22739,N_22320);
xor U22834 (N_22834,N_22140,N_22737);
or U22835 (N_22835,N_22169,N_21728);
nand U22836 (N_22836,N_22309,N_21690);
xor U22837 (N_22837,N_22627,N_22663);
xnor U22838 (N_22838,N_21904,N_21938);
xnor U22839 (N_22839,N_22486,N_22561);
nand U22840 (N_22840,N_21719,N_22798);
xor U22841 (N_22841,N_22460,N_21974);
nand U22842 (N_22842,N_22166,N_22752);
or U22843 (N_22843,N_21898,N_21646);
nor U22844 (N_22844,N_22278,N_22026);
xor U22845 (N_22845,N_22123,N_22778);
nand U22846 (N_22846,N_21629,N_21632);
nor U22847 (N_22847,N_21650,N_21665);
nor U22848 (N_22848,N_21794,N_22274);
xor U22849 (N_22849,N_22355,N_22553);
xnor U22850 (N_22850,N_21782,N_22200);
nor U22851 (N_22851,N_22687,N_21890);
and U22852 (N_22852,N_22372,N_21780);
and U22853 (N_22853,N_22594,N_22298);
nand U22854 (N_22854,N_22665,N_21891);
nor U22855 (N_22855,N_22066,N_21871);
or U22856 (N_22856,N_22360,N_22173);
xor U22857 (N_22857,N_22605,N_22338);
nor U22858 (N_22858,N_22674,N_22732);
nor U22859 (N_22859,N_22441,N_21820);
or U22860 (N_22860,N_22286,N_21988);
or U22861 (N_22861,N_21952,N_22773);
and U22862 (N_22862,N_22330,N_22733);
and U22863 (N_22863,N_22758,N_22093);
xor U22864 (N_22864,N_22349,N_22604);
xnor U22865 (N_22865,N_22648,N_22148);
nor U22866 (N_22866,N_21762,N_22128);
or U22867 (N_22867,N_22729,N_22755);
nor U22868 (N_22868,N_22033,N_22593);
or U22869 (N_22869,N_21743,N_21999);
nand U22870 (N_22870,N_21799,N_22199);
nor U22871 (N_22871,N_22451,N_22689);
or U22872 (N_22872,N_22396,N_22548);
and U22873 (N_22873,N_22696,N_22101);
nor U22874 (N_22874,N_21735,N_21893);
nand U22875 (N_22875,N_22704,N_21831);
or U22876 (N_22876,N_22555,N_22400);
nor U22877 (N_22877,N_22036,N_21681);
nor U22878 (N_22878,N_22052,N_22473);
and U22879 (N_22879,N_22531,N_22235);
xnor U22880 (N_22880,N_22493,N_22783);
nand U22881 (N_22881,N_22693,N_21708);
xor U22882 (N_22882,N_22666,N_21876);
and U22883 (N_22883,N_22406,N_21658);
xor U22884 (N_22884,N_22728,N_22233);
nand U22885 (N_22885,N_22552,N_22280);
or U22886 (N_22886,N_22769,N_22675);
and U22887 (N_22887,N_21888,N_21942);
nor U22888 (N_22888,N_22554,N_22112);
nor U22889 (N_22889,N_21963,N_21955);
nor U22890 (N_22890,N_22227,N_21703);
or U22891 (N_22891,N_22087,N_22343);
nor U22892 (N_22892,N_22480,N_22050);
nand U22893 (N_22893,N_21772,N_22727);
or U22894 (N_22894,N_22705,N_22057);
nor U22895 (N_22895,N_22526,N_21705);
xor U22896 (N_22896,N_22403,N_21935);
nor U22897 (N_22897,N_22181,N_22312);
nor U22898 (N_22898,N_21967,N_22212);
or U22899 (N_22899,N_22281,N_22346);
nand U22900 (N_22900,N_21956,N_22618);
or U22901 (N_22901,N_21713,N_21869);
and U22902 (N_22902,N_22263,N_22119);
nand U22903 (N_22903,N_21842,N_21931);
xnor U22904 (N_22904,N_22044,N_21720);
and U22905 (N_22905,N_21661,N_22768);
or U22906 (N_22906,N_22147,N_21788);
or U22907 (N_22907,N_22370,N_22209);
or U22908 (N_22908,N_22067,N_21996);
xnor U22909 (N_22909,N_21918,N_21639);
xnor U22910 (N_22910,N_22375,N_21982);
nor U22911 (N_22911,N_22624,N_22008);
nor U22912 (N_22912,N_22489,N_22725);
or U22913 (N_22913,N_22069,N_22013);
xnor U22914 (N_22914,N_22015,N_22364);
or U22915 (N_22915,N_22230,N_21771);
xnor U22916 (N_22916,N_22562,N_22469);
nor U22917 (N_22917,N_22384,N_22468);
or U22918 (N_22918,N_22239,N_22077);
and U22919 (N_22919,N_22405,N_22304);
nor U22920 (N_22920,N_21895,N_22642);
xor U22921 (N_22921,N_22242,N_22679);
and U22922 (N_22922,N_22167,N_22507);
nor U22923 (N_22923,N_21615,N_22793);
nand U22924 (N_22924,N_21882,N_22515);
xnor U22925 (N_22925,N_22660,N_22306);
or U22926 (N_22926,N_22014,N_22688);
nor U22927 (N_22927,N_22327,N_22433);
xnor U22928 (N_22928,N_22572,N_22638);
and U22929 (N_22929,N_21626,N_22075);
and U22930 (N_22930,N_22021,N_21666);
nand U22931 (N_22931,N_22471,N_22334);
nor U22932 (N_22932,N_21764,N_21654);
and U22933 (N_22933,N_21715,N_22607);
xor U22934 (N_22934,N_22600,N_22336);
and U22935 (N_22935,N_22766,N_21985);
nand U22936 (N_22936,N_22790,N_22530);
or U22937 (N_22937,N_22647,N_21770);
xor U22938 (N_22938,N_21810,N_21804);
xnor U22939 (N_22939,N_21976,N_21856);
xnor U22940 (N_22940,N_21864,N_22487);
xnor U22941 (N_22941,N_22264,N_22082);
and U22942 (N_22942,N_22423,N_22498);
nand U22943 (N_22943,N_22437,N_22363);
xor U22944 (N_22944,N_21987,N_22564);
nor U22945 (N_22945,N_22586,N_22415);
nor U22946 (N_22946,N_21644,N_21754);
nor U22947 (N_22947,N_21669,N_21817);
and U22948 (N_22948,N_21887,N_22585);
or U22949 (N_22949,N_22061,N_21722);
nor U22950 (N_22950,N_22756,N_21683);
xor U22951 (N_22951,N_22208,N_22601);
nor U22952 (N_22952,N_21973,N_21714);
or U22953 (N_22953,N_21691,N_22458);
nor U22954 (N_22954,N_22387,N_22528);
nand U22955 (N_22955,N_22436,N_22001);
and U22956 (N_22956,N_21672,N_22168);
nor U22957 (N_22957,N_21922,N_21655);
nor U22958 (N_22958,N_22096,N_21775);
xnor U22959 (N_22959,N_22152,N_21899);
xnor U22960 (N_22960,N_22643,N_22133);
and U22961 (N_22961,N_21930,N_22656);
nand U22962 (N_22962,N_22470,N_21700);
or U22963 (N_22963,N_21843,N_21923);
and U22964 (N_22964,N_22164,N_22522);
and U22965 (N_22965,N_22635,N_21628);
xnor U22966 (N_22966,N_21657,N_22310);
and U22967 (N_22967,N_22794,N_22730);
or U22968 (N_22968,N_21620,N_22767);
and U22969 (N_22969,N_22465,N_22534);
xnor U22970 (N_22970,N_21710,N_21619);
or U22971 (N_22971,N_22620,N_21746);
or U22972 (N_22972,N_22020,N_21627);
nand U22973 (N_22973,N_22284,N_22380);
or U22974 (N_22974,N_22277,N_21924);
xnor U22975 (N_22975,N_21643,N_22456);
nor U22976 (N_22976,N_22429,N_22625);
and U22977 (N_22977,N_22290,N_22784);
and U22978 (N_22978,N_21962,N_22457);
nand U22979 (N_22979,N_22357,N_22058);
nand U22980 (N_22980,N_22019,N_22422);
nand U22981 (N_22981,N_22395,N_22179);
xor U22982 (N_22982,N_22580,N_22525);
or U22983 (N_22983,N_22394,N_22719);
nand U22984 (N_22984,N_22344,N_21791);
nand U22985 (N_22985,N_22260,N_22207);
nor U22986 (N_22986,N_22645,N_21901);
and U22987 (N_22987,N_21850,N_21875);
nor U22988 (N_22988,N_22016,N_22248);
and U22989 (N_22989,N_22590,N_22464);
nor U22990 (N_22990,N_22269,N_22226);
nor U22991 (N_22991,N_21822,N_22131);
nand U22992 (N_22992,N_22113,N_22502);
nor U22993 (N_22993,N_22246,N_22398);
and U22994 (N_22994,N_22462,N_22293);
or U22995 (N_22995,N_22673,N_21902);
or U22996 (N_22996,N_22314,N_21933);
nand U22997 (N_22997,N_22434,N_22117);
xor U22998 (N_22998,N_21696,N_22723);
or U22999 (N_22999,N_22479,N_21797);
xor U23000 (N_23000,N_22583,N_21706);
or U23001 (N_23001,N_21675,N_22407);
nor U23002 (N_23002,N_22408,N_22089);
and U23003 (N_23003,N_22389,N_22628);
nand U23004 (N_23004,N_21784,N_22124);
nor U23005 (N_23005,N_21995,N_21981);
nor U23006 (N_23006,N_22362,N_22517);
xnor U23007 (N_23007,N_21604,N_22146);
nand U23008 (N_23008,N_21821,N_22105);
or U23009 (N_23009,N_22171,N_22114);
nand U23010 (N_23010,N_22511,N_21641);
xor U23011 (N_23011,N_22676,N_21844);
and U23012 (N_23012,N_22187,N_22132);
nand U23013 (N_23013,N_22744,N_21653);
nor U23014 (N_23014,N_21740,N_22027);
xnor U23015 (N_23015,N_22410,N_22401);
and U23016 (N_23016,N_22680,N_22599);
xor U23017 (N_23017,N_21965,N_21631);
or U23018 (N_23018,N_22738,N_21824);
or U23019 (N_23019,N_22291,N_22701);
or U23020 (N_23020,N_21786,N_22300);
nor U23021 (N_23021,N_22151,N_22356);
nand U23022 (N_23022,N_22413,N_21625);
nor U23023 (N_23023,N_22116,N_22512);
nand U23024 (N_23024,N_22614,N_21753);
xnor U23025 (N_23025,N_21921,N_22570);
nor U23026 (N_23026,N_21948,N_22043);
nand U23027 (N_23027,N_22107,N_21652);
and U23028 (N_23028,N_22220,N_22025);
nand U23029 (N_23029,N_22243,N_22651);
and U23030 (N_23030,N_22399,N_21768);
or U23031 (N_23031,N_22340,N_21636);
xnor U23032 (N_23032,N_22477,N_22289);
nor U23033 (N_23033,N_22497,N_22103);
xnor U23034 (N_23034,N_22777,N_21847);
xor U23035 (N_23035,N_22307,N_21676);
nor U23036 (N_23036,N_22598,N_22508);
or U23037 (N_23037,N_21711,N_22323);
xor U23038 (N_23038,N_21785,N_22404);
and U23039 (N_23039,N_21870,N_22039);
xor U23040 (N_23040,N_21633,N_22703);
xor U23041 (N_23041,N_22313,N_21756);
nand U23042 (N_23042,N_22708,N_22393);
nor U23043 (N_23043,N_22296,N_22445);
nand U23044 (N_23044,N_21868,N_21825);
or U23045 (N_23045,N_22251,N_22467);
or U23046 (N_23046,N_22383,N_22294);
nand U23047 (N_23047,N_21663,N_22084);
nor U23048 (N_23048,N_22022,N_22420);
nand U23049 (N_23049,N_22094,N_22359);
nand U23050 (N_23050,N_22641,N_22472);
or U23051 (N_23051,N_22198,N_21885);
and U23052 (N_23052,N_22495,N_22667);
and U23053 (N_23053,N_21867,N_21861);
nand U23054 (N_23054,N_21637,N_22134);
nor U23055 (N_23055,N_21829,N_22485);
nor U23056 (N_23056,N_21980,N_21697);
or U23057 (N_23057,N_22035,N_22587);
xnor U23058 (N_23058,N_21813,N_21896);
nand U23059 (N_23059,N_22615,N_21879);
or U23060 (N_23060,N_22158,N_22543);
or U23061 (N_23061,N_22484,N_22170);
nand U23062 (N_23062,N_22201,N_22379);
nand U23063 (N_23063,N_22700,N_22315);
xnor U23064 (N_23064,N_21977,N_22453);
nand U23065 (N_23065,N_22038,N_22210);
or U23066 (N_23066,N_21621,N_21939);
xnor U23067 (N_23067,N_21677,N_21695);
xor U23068 (N_23068,N_22073,N_22136);
nand U23069 (N_23069,N_22162,N_22521);
xnor U23070 (N_23070,N_22771,N_22063);
xor U23071 (N_23071,N_22613,N_21789);
xnor U23072 (N_23072,N_21698,N_22229);
and U23073 (N_23073,N_21991,N_22478);
nand U23074 (N_23074,N_21668,N_21769);
nor U23075 (N_23075,N_22789,N_22529);
xnor U23076 (N_23076,N_22750,N_22652);
nor U23077 (N_23077,N_21993,N_21727);
nand U23078 (N_23078,N_22367,N_22257);
and U23079 (N_23079,N_22621,N_21915);
xnor U23080 (N_23080,N_22139,N_22440);
nand U23081 (N_23081,N_22062,N_21881);
or U23082 (N_23082,N_22551,N_22442);
nand U23083 (N_23083,N_22516,N_22010);
and U23084 (N_23084,N_22731,N_21857);
and U23085 (N_23085,N_21910,N_22002);
or U23086 (N_23086,N_21927,N_22760);
and U23087 (N_23087,N_22347,N_22378);
xnor U23088 (N_23088,N_22549,N_21742);
and U23089 (N_23089,N_21717,N_22185);
and U23090 (N_23090,N_21950,N_21671);
nor U23091 (N_23091,N_21779,N_22361);
nand U23092 (N_23092,N_22716,N_22713);
xor U23093 (N_23093,N_22004,N_21622);
nor U23094 (N_23094,N_21841,N_21694);
xnor U23095 (N_23095,N_22799,N_21600);
nor U23096 (N_23096,N_22017,N_21994);
nor U23097 (N_23097,N_22626,N_22617);
nor U23098 (N_23098,N_22509,N_21680);
and U23099 (N_23099,N_22202,N_21865);
nand U23100 (N_23100,N_22056,N_22556);
or U23101 (N_23101,N_22326,N_22753);
xnor U23102 (N_23102,N_21640,N_21712);
nand U23103 (N_23103,N_22761,N_22046);
nor U23104 (N_23104,N_22098,N_22273);
or U23105 (N_23105,N_22097,N_22770);
or U23106 (N_23106,N_22520,N_22706);
nor U23107 (N_23107,N_22060,N_22707);
and U23108 (N_23108,N_22563,N_21725);
or U23109 (N_23109,N_21701,N_21718);
and U23110 (N_23110,N_22749,N_22686);
and U23111 (N_23111,N_22178,N_22135);
or U23112 (N_23112,N_22421,N_21866);
xnor U23113 (N_23113,N_22272,N_21819);
and U23114 (N_23114,N_22711,N_22782);
nor U23115 (N_23115,N_22154,N_22322);
and U23116 (N_23116,N_21607,N_22215);
and U23117 (N_23117,N_22329,N_22092);
nor U23118 (N_23118,N_22425,N_21787);
nand U23119 (N_23119,N_22637,N_22255);
nand U23120 (N_23120,N_22218,N_22256);
nor U23121 (N_23121,N_22541,N_22332);
xor U23122 (N_23122,N_22579,N_22644);
nor U23123 (N_23123,N_21907,N_21734);
or U23124 (N_23124,N_22566,N_22721);
nand U23125 (N_23125,N_21815,N_21909);
xnor U23126 (N_23126,N_22177,N_22258);
or U23127 (N_23127,N_22348,N_22757);
nor U23128 (N_23128,N_22654,N_21878);
or U23129 (N_23129,N_22204,N_21679);
xor U23130 (N_23130,N_22369,N_22217);
nand U23131 (N_23131,N_22055,N_22699);
nor U23132 (N_23132,N_22254,N_21998);
nand U23133 (N_23133,N_22341,N_22302);
or U23134 (N_23134,N_21726,N_22048);
nand U23135 (N_23135,N_21947,N_22611);
nand U23136 (N_23136,N_22715,N_21983);
xnor U23137 (N_23137,N_22668,N_22271);
xnor U23138 (N_23138,N_22702,N_22331);
xnor U23139 (N_23139,N_22144,N_21826);
and U23140 (N_23140,N_22710,N_21903);
xor U23141 (N_23141,N_21894,N_22439);
nor U23142 (N_23142,N_22023,N_22610);
xnor U23143 (N_23143,N_22589,N_22785);
nor U23144 (N_23144,N_21678,N_22714);
and U23145 (N_23145,N_22018,N_22482);
nand U23146 (N_23146,N_22476,N_22795);
xor U23147 (N_23147,N_21883,N_21997);
nand U23148 (N_23148,N_21961,N_22049);
or U23149 (N_23149,N_21840,N_22122);
nor U23150 (N_23150,N_22350,N_21807);
or U23151 (N_23151,N_21651,N_21862);
nand U23152 (N_23152,N_22427,N_21833);
xor U23153 (N_23153,N_22392,N_21709);
xnor U23154 (N_23154,N_21849,N_22672);
xnor U23155 (N_23155,N_22402,N_21755);
nor U23156 (N_23156,N_22619,N_21814);
and U23157 (N_23157,N_22698,N_22595);
or U23158 (N_23158,N_21759,N_22718);
nor U23159 (N_23159,N_22388,N_21897);
and U23160 (N_23160,N_22206,N_21941);
nand U23161 (N_23161,N_21623,N_21827);
nor U23162 (N_23162,N_22045,N_21839);
or U23163 (N_23163,N_21776,N_21964);
xnor U23164 (N_23164,N_21724,N_22537);
nand U23165 (N_23165,N_22104,N_21832);
nor U23166 (N_23166,N_22011,N_21739);
nand U23167 (N_23167,N_22694,N_21730);
nor U23168 (N_23168,N_21913,N_21630);
and U23169 (N_23169,N_22259,N_22252);
or U23170 (N_23170,N_21968,N_21610);
and U23171 (N_23171,N_22244,N_22214);
and U23172 (N_23172,N_22276,N_22308);
nor U23173 (N_23173,N_22682,N_22079);
and U23174 (N_23174,N_21649,N_22261);
nand U23175 (N_23175,N_21969,N_22371);
xnor U23176 (N_23176,N_21702,N_22126);
and U23177 (N_23177,N_21925,N_22792);
nand U23178 (N_23178,N_22622,N_21693);
nor U23179 (N_23179,N_22282,N_22000);
or U23180 (N_23180,N_21940,N_21790);
nand U23181 (N_23181,N_22754,N_22759);
nor U23182 (N_23182,N_22591,N_22390);
nor U23183 (N_23183,N_22031,N_21765);
xnor U23184 (N_23184,N_21837,N_21795);
or U23185 (N_23185,N_22496,N_22426);
xor U23186 (N_23186,N_22382,N_21806);
xnor U23187 (N_23187,N_22358,N_21616);
nand U23188 (N_23188,N_21834,N_22193);
and U23189 (N_23189,N_22629,N_22160);
or U23190 (N_23190,N_21684,N_22763);
nor U23191 (N_23191,N_22279,N_21818);
nor U23192 (N_23192,N_22649,N_22137);
xnor U23193 (N_23193,N_22746,N_22029);
xnor U23194 (N_23194,N_22505,N_21971);
nand U23195 (N_23195,N_21989,N_22443);
nand U23196 (N_23196,N_21953,N_22419);
or U23197 (N_23197,N_21816,N_21889);
nor U23198 (N_23198,N_22184,N_22028);
nor U23199 (N_23199,N_22483,N_22145);
xor U23200 (N_23200,N_22670,N_21944);
nor U23201 (N_23201,N_22109,N_21811);
and U23202 (N_23202,N_21892,N_22466);
nor U23203 (N_23203,N_22163,N_22747);
nor U23204 (N_23204,N_21738,N_21624);
nor U23205 (N_23205,N_22582,N_22070);
or U23206 (N_23206,N_22099,N_22270);
xor U23207 (N_23207,N_22127,N_22175);
nand U23208 (N_23208,N_22671,N_21608);
nor U23209 (N_23209,N_22032,N_21614);
and U23210 (N_23210,N_22397,N_21877);
nor U23211 (N_23211,N_21926,N_21914);
and U23212 (N_23212,N_22797,N_22129);
nor U23213 (N_23213,N_22065,N_22234);
nor U23214 (N_23214,N_21733,N_21686);
nor U23215 (N_23215,N_22337,N_21737);
nand U23216 (N_23216,N_21809,N_22368);
or U23217 (N_23217,N_21838,N_21958);
xor U23218 (N_23218,N_21929,N_22176);
and U23219 (N_23219,N_22034,N_22424);
nor U23220 (N_23220,N_22086,N_22321);
nor U23221 (N_23221,N_22159,N_22491);
xnor U23222 (N_23222,N_22742,N_22596);
nand U23223 (N_23223,N_21603,N_22157);
nor U23224 (N_23224,N_22188,N_22662);
or U23225 (N_23225,N_22412,N_22138);
and U23226 (N_23226,N_22558,N_22720);
nand U23227 (N_23227,N_22560,N_22547);
xor U23228 (N_23228,N_22779,N_22655);
nand U23229 (N_23229,N_22351,N_22374);
or U23230 (N_23230,N_22183,N_22475);
and U23231 (N_23231,N_22535,N_22203);
or U23232 (N_23232,N_22636,N_22448);
xor U23233 (N_23233,N_21781,N_22791);
nand U23234 (N_23234,N_21884,N_22325);
or U23235 (N_23235,N_21736,N_22051);
xnor U23236 (N_23236,N_21744,N_22630);
and U23237 (N_23237,N_21748,N_22612);
nor U23238 (N_23238,N_21602,N_21943);
xnor U23239 (N_23239,N_21642,N_21846);
nand U23240 (N_23240,N_22735,N_22565);
xor U23241 (N_23241,N_22444,N_21905);
xor U23242 (N_23242,N_21638,N_22054);
or U23243 (N_23243,N_21729,N_22411);
nand U23244 (N_23244,N_21970,N_21957);
nand U23245 (N_23245,N_21617,N_22712);
or U23246 (N_23246,N_22189,N_22303);
or U23247 (N_23247,N_22120,N_22697);
and U23248 (N_23248,N_22205,N_21802);
nand U23249 (N_23249,N_22125,N_22335);
xnor U23250 (N_23250,N_22090,N_22446);
nand U23251 (N_23251,N_22449,N_22299);
and U23252 (N_23252,N_22095,N_22581);
xnor U23253 (N_23253,N_22539,N_21812);
xnor U23254 (N_23254,N_22775,N_22301);
or U23255 (N_23255,N_22353,N_22165);
nand U23256 (N_23256,N_22447,N_22241);
nor U23257 (N_23257,N_22366,N_22236);
or U23258 (N_23258,N_21863,N_21801);
xor U23259 (N_23259,N_22354,N_22249);
xor U23260 (N_23260,N_22499,N_22385);
or U23261 (N_23261,N_21777,N_22544);
and U23262 (N_23262,N_22216,N_22432);
nor U23263 (N_23263,N_22080,N_22450);
xnor U23264 (N_23264,N_22182,N_22650);
nor U23265 (N_23265,N_22751,N_22194);
or U23266 (N_23266,N_21836,N_21648);
xor U23267 (N_23267,N_22664,N_22003);
nand U23268 (N_23268,N_22081,N_21766);
nor U23269 (N_23269,N_22435,N_22012);
nand U23270 (N_23270,N_22042,N_22071);
or U23271 (N_23271,N_21798,N_21908);
and U23272 (N_23272,N_22722,N_22695);
nand U23273 (N_23273,N_22640,N_21618);
or U23274 (N_23274,N_22213,N_22683);
xnor U23275 (N_23275,N_22780,N_22319);
nand U23276 (N_23276,N_22431,N_22037);
xnor U23277 (N_23277,N_22342,N_22550);
and U23278 (N_23278,N_22692,N_21860);
nand U23279 (N_23279,N_22527,N_21670);
or U23280 (N_23280,N_22083,N_22559);
xor U23281 (N_23281,N_22283,N_22574);
or U23282 (N_23282,N_21761,N_22153);
nor U23283 (N_23283,N_22454,N_22292);
and U23284 (N_23284,N_21906,N_21699);
nand U23285 (N_23285,N_21900,N_22634);
nor U23286 (N_23286,N_21704,N_22245);
or U23287 (N_23287,N_22268,N_21635);
nor U23288 (N_23288,N_22339,N_22219);
nor U23289 (N_23289,N_22041,N_22288);
xor U23290 (N_23290,N_22172,N_21972);
nand U23291 (N_23291,N_22633,N_21659);
nor U23292 (N_23292,N_21934,N_22240);
and U23293 (N_23293,N_21851,N_22118);
nor U23294 (N_23294,N_21745,N_21783);
xor U23295 (N_23295,N_22381,N_21979);
xnor U23296 (N_23296,N_22076,N_22736);
nand U23297 (N_23297,N_22510,N_22130);
nor U23298 (N_23298,N_22745,N_21853);
nor U23299 (N_23299,N_21796,N_21800);
nand U23300 (N_23300,N_22616,N_21664);
xor U23301 (N_23301,N_21605,N_22681);
and U23302 (N_23302,N_22592,N_21613);
nor U23303 (N_23303,N_22494,N_21949);
or U23304 (N_23304,N_22748,N_22438);
nor U23305 (N_23305,N_21990,N_22519);
xor U23306 (N_23306,N_22575,N_22518);
or U23307 (N_23307,N_22588,N_22232);
nand U23308 (N_23308,N_22631,N_22262);
and U23309 (N_23309,N_22238,N_22006);
or U23310 (N_23310,N_22155,N_21986);
xnor U23311 (N_23311,N_22333,N_21854);
nand U23312 (N_23312,N_22174,N_22538);
xor U23313 (N_23313,N_21805,N_22409);
and U23314 (N_23314,N_22386,N_21606);
nand U23315 (N_23315,N_22074,N_22141);
or U23316 (N_23316,N_22266,N_21612);
xor U23317 (N_23317,N_22197,N_22192);
and U23318 (N_23318,N_22186,N_22391);
xor U23319 (N_23319,N_22328,N_22787);
and U23320 (N_23320,N_22776,N_22602);
xor U23321 (N_23321,N_21848,N_22573);
nor U23322 (N_23322,N_22772,N_22690);
or U23323 (N_23323,N_22305,N_22490);
or U23324 (N_23324,N_22222,N_21936);
xor U23325 (N_23325,N_21823,N_22532);
and U23326 (N_23326,N_22142,N_22024);
or U23327 (N_23327,N_22488,N_21928);
nand U23328 (N_23328,N_22085,N_22653);
nand U23329 (N_23329,N_22691,N_21692);
and U23330 (N_23330,N_22734,N_22196);
or U23331 (N_23331,N_21937,N_21872);
or U23332 (N_23332,N_21660,N_21919);
and U23333 (N_23333,N_22578,N_21803);
nor U23334 (N_23334,N_21858,N_22513);
or U23335 (N_23335,N_21689,N_22608);
and U23336 (N_23336,N_22191,N_22318);
nand U23337 (N_23337,N_22603,N_22149);
and U23338 (N_23338,N_22285,N_22577);
xnor U23339 (N_23339,N_22416,N_21946);
and U23340 (N_23340,N_22658,N_22078);
or U23341 (N_23341,N_21945,N_22156);
and U23342 (N_23342,N_22418,N_22576);
xor U23343 (N_23343,N_22287,N_22743);
nor U23344 (N_23344,N_22669,N_21767);
nor U23345 (N_23345,N_21763,N_22091);
xor U23346 (N_23346,N_22503,N_22557);
nor U23347 (N_23347,N_22009,N_22068);
nand U23348 (N_23348,N_22481,N_22110);
and U23349 (N_23349,N_21656,N_21975);
or U23350 (N_23350,N_22765,N_22461);
or U23351 (N_23351,N_22463,N_21688);
and U23352 (N_23352,N_22545,N_22180);
xnor U23353 (N_23353,N_22247,N_22524);
or U23354 (N_23354,N_22064,N_21873);
or U23355 (N_23355,N_22428,N_22501);
or U23356 (N_23356,N_21992,N_21984);
nor U23357 (N_23357,N_22677,N_22504);
nand U23358 (N_23358,N_22500,N_22709);
nand U23359 (N_23359,N_22324,N_21880);
xnor U23360 (N_23360,N_22781,N_21960);
nor U23361 (N_23361,N_21954,N_21757);
nor U23362 (N_23362,N_22646,N_21830);
and U23363 (N_23363,N_21645,N_22571);
or U23364 (N_23364,N_21773,N_22685);
xor U23365 (N_23365,N_21721,N_21978);
nand U23366 (N_23366,N_22659,N_21845);
nor U23367 (N_23367,N_22606,N_22678);
nor U23368 (N_23368,N_22221,N_22788);
nor U23369 (N_23369,N_22365,N_21667);
nand U23370 (N_23370,N_22211,N_22724);
nand U23371 (N_23371,N_21793,N_22540);
nand U23372 (N_23372,N_22796,N_21647);
or U23373 (N_23373,N_22536,N_21917);
xnor U23374 (N_23374,N_21912,N_22459);
xor U23375 (N_23375,N_22007,N_21716);
and U23376 (N_23376,N_21859,N_22632);
nor U23377 (N_23377,N_22311,N_22108);
or U23378 (N_23378,N_22514,N_22088);
xor U23379 (N_23379,N_22352,N_22376);
nand U23380 (N_23380,N_22657,N_22195);
or U23381 (N_23381,N_22684,N_22190);
nand U23382 (N_23382,N_21852,N_21673);
xor U23383 (N_23383,N_22295,N_21609);
nand U23384 (N_23384,N_22072,N_21707);
nor U23385 (N_23385,N_22005,N_22597);
nor U23386 (N_23386,N_21778,N_22430);
nor U23387 (N_23387,N_22316,N_21732);
nor U23388 (N_23388,N_22569,N_22121);
xor U23389 (N_23389,N_21731,N_22253);
nor U23390 (N_23390,N_22111,N_21682);
xor U23391 (N_23391,N_21951,N_22267);
or U23392 (N_23392,N_22047,N_21723);
or U23393 (N_23393,N_21916,N_21874);
or U23394 (N_23394,N_22297,N_21911);
and U23395 (N_23395,N_22492,N_21920);
or U23396 (N_23396,N_22786,N_22231);
and U23397 (N_23397,N_22115,N_21959);
nor U23398 (N_23398,N_22584,N_22506);
or U23399 (N_23399,N_22275,N_22377);
or U23400 (N_23400,N_22186,N_21730);
nor U23401 (N_23401,N_22416,N_21774);
or U23402 (N_23402,N_21869,N_22343);
xnor U23403 (N_23403,N_22673,N_22749);
and U23404 (N_23404,N_21651,N_22528);
xor U23405 (N_23405,N_22744,N_22655);
or U23406 (N_23406,N_22686,N_21977);
nor U23407 (N_23407,N_22400,N_22624);
xor U23408 (N_23408,N_22069,N_21719);
and U23409 (N_23409,N_22393,N_21787);
and U23410 (N_23410,N_21919,N_21985);
or U23411 (N_23411,N_22018,N_22453);
nor U23412 (N_23412,N_22187,N_22000);
nand U23413 (N_23413,N_22340,N_22777);
xor U23414 (N_23414,N_22715,N_22624);
nand U23415 (N_23415,N_22481,N_22145);
nor U23416 (N_23416,N_22760,N_21783);
nor U23417 (N_23417,N_22357,N_21990);
nor U23418 (N_23418,N_21699,N_22283);
nand U23419 (N_23419,N_22242,N_21885);
nor U23420 (N_23420,N_22021,N_22127);
nand U23421 (N_23421,N_22666,N_22341);
nand U23422 (N_23422,N_22201,N_22073);
xor U23423 (N_23423,N_22384,N_22358);
nand U23424 (N_23424,N_21927,N_22173);
and U23425 (N_23425,N_22245,N_21699);
or U23426 (N_23426,N_22219,N_22047);
xor U23427 (N_23427,N_22611,N_21713);
and U23428 (N_23428,N_22146,N_21994);
xnor U23429 (N_23429,N_22631,N_22244);
nand U23430 (N_23430,N_22319,N_22240);
nand U23431 (N_23431,N_21800,N_22222);
nor U23432 (N_23432,N_22179,N_21620);
or U23433 (N_23433,N_22581,N_22260);
nor U23434 (N_23434,N_21887,N_22159);
and U23435 (N_23435,N_22687,N_22123);
nand U23436 (N_23436,N_22404,N_22699);
and U23437 (N_23437,N_21733,N_21956);
nor U23438 (N_23438,N_22352,N_22670);
nand U23439 (N_23439,N_21704,N_21945);
or U23440 (N_23440,N_22234,N_22551);
or U23441 (N_23441,N_22591,N_22206);
xor U23442 (N_23442,N_21696,N_22664);
nor U23443 (N_23443,N_22094,N_21811);
nor U23444 (N_23444,N_22541,N_21945);
or U23445 (N_23445,N_21751,N_22177);
nand U23446 (N_23446,N_21869,N_22792);
and U23447 (N_23447,N_22108,N_21972);
xnor U23448 (N_23448,N_22602,N_21875);
xnor U23449 (N_23449,N_21675,N_21826);
nand U23450 (N_23450,N_22646,N_22726);
nor U23451 (N_23451,N_21998,N_22496);
nand U23452 (N_23452,N_21714,N_22225);
nor U23453 (N_23453,N_21742,N_22131);
nor U23454 (N_23454,N_22767,N_22484);
and U23455 (N_23455,N_22463,N_21816);
or U23456 (N_23456,N_21616,N_22301);
nor U23457 (N_23457,N_22239,N_22590);
xnor U23458 (N_23458,N_21690,N_21861);
xor U23459 (N_23459,N_22361,N_21825);
nand U23460 (N_23460,N_21960,N_22694);
or U23461 (N_23461,N_22467,N_22771);
or U23462 (N_23462,N_22344,N_22356);
or U23463 (N_23463,N_21927,N_22499);
nand U23464 (N_23464,N_22348,N_21943);
nand U23465 (N_23465,N_22217,N_22597);
and U23466 (N_23466,N_22480,N_21888);
nand U23467 (N_23467,N_21753,N_22133);
xnor U23468 (N_23468,N_22036,N_22245);
or U23469 (N_23469,N_22682,N_22555);
xnor U23470 (N_23470,N_22662,N_22089);
and U23471 (N_23471,N_22426,N_22582);
nand U23472 (N_23472,N_22433,N_22447);
xor U23473 (N_23473,N_22746,N_22618);
or U23474 (N_23474,N_21890,N_21717);
xnor U23475 (N_23475,N_21923,N_21975);
xnor U23476 (N_23476,N_21808,N_22773);
nand U23477 (N_23477,N_22650,N_22286);
xor U23478 (N_23478,N_22743,N_21657);
xnor U23479 (N_23479,N_22014,N_22353);
and U23480 (N_23480,N_21911,N_22690);
nand U23481 (N_23481,N_21693,N_22233);
xnor U23482 (N_23482,N_21769,N_22228);
xnor U23483 (N_23483,N_22465,N_21711);
nand U23484 (N_23484,N_22375,N_21601);
xnor U23485 (N_23485,N_22338,N_22637);
and U23486 (N_23486,N_21979,N_22394);
or U23487 (N_23487,N_22057,N_22074);
nand U23488 (N_23488,N_22513,N_22533);
and U23489 (N_23489,N_21904,N_22494);
xor U23490 (N_23490,N_21822,N_21777);
nor U23491 (N_23491,N_22260,N_21766);
and U23492 (N_23492,N_22173,N_21911);
or U23493 (N_23493,N_21676,N_22695);
or U23494 (N_23494,N_21906,N_21662);
or U23495 (N_23495,N_22351,N_22179);
nor U23496 (N_23496,N_21621,N_22664);
nand U23497 (N_23497,N_22147,N_21976);
or U23498 (N_23498,N_22772,N_22696);
nor U23499 (N_23499,N_22317,N_22071);
nand U23500 (N_23500,N_21957,N_22257);
nor U23501 (N_23501,N_21618,N_21892);
or U23502 (N_23502,N_21883,N_22233);
nand U23503 (N_23503,N_21911,N_22431);
nand U23504 (N_23504,N_21856,N_22349);
and U23505 (N_23505,N_22062,N_22142);
nand U23506 (N_23506,N_22708,N_22183);
nand U23507 (N_23507,N_21869,N_21617);
and U23508 (N_23508,N_21979,N_22431);
xor U23509 (N_23509,N_22178,N_22252);
and U23510 (N_23510,N_22488,N_22108);
or U23511 (N_23511,N_22733,N_21872);
nand U23512 (N_23512,N_22756,N_22639);
nor U23513 (N_23513,N_21830,N_22106);
nand U23514 (N_23514,N_21922,N_22727);
nand U23515 (N_23515,N_22624,N_22072);
nand U23516 (N_23516,N_22112,N_21680);
or U23517 (N_23517,N_22103,N_21671);
or U23518 (N_23518,N_22334,N_22599);
nor U23519 (N_23519,N_22075,N_22716);
xnor U23520 (N_23520,N_22678,N_22604);
or U23521 (N_23521,N_21894,N_22763);
nor U23522 (N_23522,N_21653,N_22268);
and U23523 (N_23523,N_22633,N_22345);
nand U23524 (N_23524,N_22533,N_22109);
xor U23525 (N_23525,N_22770,N_21641);
or U23526 (N_23526,N_22095,N_22451);
nor U23527 (N_23527,N_21754,N_21852);
or U23528 (N_23528,N_21791,N_22696);
xor U23529 (N_23529,N_21710,N_21876);
xnor U23530 (N_23530,N_22151,N_21869);
nor U23531 (N_23531,N_21935,N_21756);
xor U23532 (N_23532,N_22394,N_21651);
nor U23533 (N_23533,N_22016,N_22311);
or U23534 (N_23534,N_22682,N_22598);
nand U23535 (N_23535,N_21789,N_22218);
nand U23536 (N_23536,N_22499,N_21784);
nor U23537 (N_23537,N_22313,N_22019);
or U23538 (N_23538,N_22343,N_21678);
nand U23539 (N_23539,N_21890,N_21885);
nand U23540 (N_23540,N_21764,N_22591);
and U23541 (N_23541,N_21829,N_22246);
or U23542 (N_23542,N_22542,N_21913);
xor U23543 (N_23543,N_22515,N_21707);
nor U23544 (N_23544,N_22536,N_22270);
nand U23545 (N_23545,N_21682,N_21817);
and U23546 (N_23546,N_22665,N_21866);
xnor U23547 (N_23547,N_22189,N_22324);
or U23548 (N_23548,N_22683,N_21810);
and U23549 (N_23549,N_21750,N_22713);
xnor U23550 (N_23550,N_22684,N_22359);
nand U23551 (N_23551,N_21870,N_22750);
and U23552 (N_23552,N_21608,N_22321);
nand U23553 (N_23553,N_22784,N_21818);
or U23554 (N_23554,N_21712,N_22392);
nand U23555 (N_23555,N_22579,N_21827);
or U23556 (N_23556,N_22676,N_22183);
nand U23557 (N_23557,N_21939,N_22012);
and U23558 (N_23558,N_21728,N_21925);
and U23559 (N_23559,N_21704,N_22609);
or U23560 (N_23560,N_22148,N_22611);
nand U23561 (N_23561,N_22421,N_22048);
nor U23562 (N_23562,N_22231,N_22547);
nand U23563 (N_23563,N_21978,N_22275);
nand U23564 (N_23564,N_22649,N_21977);
nand U23565 (N_23565,N_22051,N_22112);
nand U23566 (N_23566,N_22596,N_22156);
nand U23567 (N_23567,N_21846,N_22757);
or U23568 (N_23568,N_21634,N_22426);
nor U23569 (N_23569,N_22250,N_22240);
or U23570 (N_23570,N_22269,N_22706);
nand U23571 (N_23571,N_22768,N_22352);
nand U23572 (N_23572,N_22299,N_21900);
nor U23573 (N_23573,N_22228,N_22163);
or U23574 (N_23574,N_22210,N_22330);
or U23575 (N_23575,N_22704,N_22496);
xor U23576 (N_23576,N_22140,N_22722);
nand U23577 (N_23577,N_22171,N_22634);
nor U23578 (N_23578,N_22623,N_22280);
xor U23579 (N_23579,N_22203,N_22409);
nor U23580 (N_23580,N_22610,N_22468);
and U23581 (N_23581,N_22236,N_21845);
xnor U23582 (N_23582,N_22406,N_22589);
nor U23583 (N_23583,N_21835,N_21746);
or U23584 (N_23584,N_21772,N_21778);
xor U23585 (N_23585,N_22153,N_22486);
nand U23586 (N_23586,N_22765,N_21840);
nor U23587 (N_23587,N_21840,N_21654);
nor U23588 (N_23588,N_22792,N_22005);
nand U23589 (N_23589,N_22639,N_22202);
nor U23590 (N_23590,N_22628,N_21941);
nor U23591 (N_23591,N_22116,N_21899);
or U23592 (N_23592,N_21946,N_22718);
xnor U23593 (N_23593,N_22077,N_22485);
nand U23594 (N_23594,N_22613,N_22303);
or U23595 (N_23595,N_22135,N_21863);
xnor U23596 (N_23596,N_21602,N_22682);
xnor U23597 (N_23597,N_22580,N_22275);
nor U23598 (N_23598,N_22705,N_21928);
or U23599 (N_23599,N_21928,N_22595);
or U23600 (N_23600,N_22388,N_22699);
xor U23601 (N_23601,N_22001,N_22636);
nand U23602 (N_23602,N_22508,N_22087);
nand U23603 (N_23603,N_22181,N_22682);
and U23604 (N_23604,N_21760,N_21672);
and U23605 (N_23605,N_22652,N_22468);
nor U23606 (N_23606,N_22231,N_22446);
xnor U23607 (N_23607,N_21733,N_21711);
or U23608 (N_23608,N_21881,N_22539);
xnor U23609 (N_23609,N_21851,N_21922);
nor U23610 (N_23610,N_22125,N_22153);
xnor U23611 (N_23611,N_22678,N_22545);
nand U23612 (N_23612,N_22247,N_22602);
nand U23613 (N_23613,N_21747,N_22421);
nand U23614 (N_23614,N_22210,N_22041);
xnor U23615 (N_23615,N_21722,N_22602);
nor U23616 (N_23616,N_22081,N_22079);
xor U23617 (N_23617,N_22570,N_21737);
nand U23618 (N_23618,N_22198,N_22338);
nor U23619 (N_23619,N_22454,N_22463);
or U23620 (N_23620,N_22150,N_22171);
nand U23621 (N_23621,N_22463,N_22495);
nor U23622 (N_23622,N_21749,N_22227);
and U23623 (N_23623,N_22737,N_22777);
nor U23624 (N_23624,N_22380,N_21623);
and U23625 (N_23625,N_22550,N_22103);
or U23626 (N_23626,N_22503,N_21702);
nand U23627 (N_23627,N_21972,N_22191);
and U23628 (N_23628,N_21691,N_22439);
nand U23629 (N_23629,N_22508,N_22185);
xor U23630 (N_23630,N_22004,N_21605);
nand U23631 (N_23631,N_22324,N_22442);
nor U23632 (N_23632,N_22096,N_22574);
or U23633 (N_23633,N_21916,N_22438);
or U23634 (N_23634,N_22197,N_22774);
or U23635 (N_23635,N_22565,N_22417);
nor U23636 (N_23636,N_22790,N_21790);
or U23637 (N_23637,N_21796,N_22260);
and U23638 (N_23638,N_22573,N_22435);
nand U23639 (N_23639,N_21803,N_22094);
xnor U23640 (N_23640,N_22125,N_22749);
or U23641 (N_23641,N_21867,N_22677);
xnor U23642 (N_23642,N_22616,N_21921);
or U23643 (N_23643,N_21867,N_21688);
nand U23644 (N_23644,N_22089,N_22619);
nand U23645 (N_23645,N_22589,N_22640);
nor U23646 (N_23646,N_22642,N_22237);
nor U23647 (N_23647,N_22144,N_21778);
or U23648 (N_23648,N_21608,N_21735);
nor U23649 (N_23649,N_22796,N_21775);
and U23650 (N_23650,N_22702,N_21815);
nand U23651 (N_23651,N_22675,N_22425);
xor U23652 (N_23652,N_22007,N_21924);
nor U23653 (N_23653,N_22733,N_21782);
xor U23654 (N_23654,N_22542,N_22431);
nor U23655 (N_23655,N_22760,N_22088);
or U23656 (N_23656,N_22645,N_22021);
nor U23657 (N_23657,N_22078,N_21894);
nor U23658 (N_23658,N_21745,N_22103);
nand U23659 (N_23659,N_22408,N_22524);
or U23660 (N_23660,N_21949,N_21957);
and U23661 (N_23661,N_22162,N_22695);
nor U23662 (N_23662,N_21646,N_21862);
nor U23663 (N_23663,N_22285,N_22557);
or U23664 (N_23664,N_22289,N_21793);
and U23665 (N_23665,N_22727,N_21961);
xor U23666 (N_23666,N_22290,N_21927);
or U23667 (N_23667,N_21686,N_22372);
or U23668 (N_23668,N_22070,N_22704);
or U23669 (N_23669,N_21979,N_21833);
or U23670 (N_23670,N_22236,N_22011);
or U23671 (N_23671,N_21971,N_22436);
nor U23672 (N_23672,N_22633,N_22066);
or U23673 (N_23673,N_22079,N_21948);
nor U23674 (N_23674,N_22133,N_22141);
or U23675 (N_23675,N_22132,N_22346);
nor U23676 (N_23676,N_21610,N_22083);
xnor U23677 (N_23677,N_22084,N_21761);
and U23678 (N_23678,N_22466,N_22795);
xnor U23679 (N_23679,N_22357,N_21735);
xor U23680 (N_23680,N_22394,N_22168);
nand U23681 (N_23681,N_22687,N_21615);
and U23682 (N_23682,N_21903,N_22673);
and U23683 (N_23683,N_22068,N_21641);
nor U23684 (N_23684,N_21773,N_22052);
and U23685 (N_23685,N_22342,N_22795);
nor U23686 (N_23686,N_22322,N_22777);
xnor U23687 (N_23687,N_21807,N_22209);
nor U23688 (N_23688,N_22236,N_21779);
nand U23689 (N_23689,N_22456,N_21744);
and U23690 (N_23690,N_22772,N_22383);
nand U23691 (N_23691,N_22616,N_22730);
xnor U23692 (N_23692,N_21722,N_22230);
nand U23693 (N_23693,N_21823,N_22186);
nand U23694 (N_23694,N_21907,N_21902);
nand U23695 (N_23695,N_22079,N_22045);
and U23696 (N_23696,N_21902,N_22642);
and U23697 (N_23697,N_21700,N_22205);
nor U23698 (N_23698,N_21687,N_22528);
nand U23699 (N_23699,N_21624,N_22772);
and U23700 (N_23700,N_21752,N_22529);
and U23701 (N_23701,N_21737,N_22562);
and U23702 (N_23702,N_21955,N_21605);
xnor U23703 (N_23703,N_22797,N_21763);
xnor U23704 (N_23704,N_22712,N_21663);
and U23705 (N_23705,N_21854,N_22669);
nand U23706 (N_23706,N_22601,N_22011);
nor U23707 (N_23707,N_21897,N_21875);
xnor U23708 (N_23708,N_22292,N_21949);
or U23709 (N_23709,N_22534,N_22284);
or U23710 (N_23710,N_22757,N_22371);
nand U23711 (N_23711,N_21816,N_21639);
and U23712 (N_23712,N_21826,N_22453);
xnor U23713 (N_23713,N_22141,N_22455);
nand U23714 (N_23714,N_22334,N_21930);
and U23715 (N_23715,N_22741,N_21705);
nor U23716 (N_23716,N_21997,N_21904);
and U23717 (N_23717,N_22275,N_22171);
or U23718 (N_23718,N_21767,N_22689);
nor U23719 (N_23719,N_21786,N_22367);
nand U23720 (N_23720,N_22334,N_22081);
nand U23721 (N_23721,N_21697,N_22565);
nand U23722 (N_23722,N_21818,N_22422);
nand U23723 (N_23723,N_22200,N_22078);
nor U23724 (N_23724,N_21950,N_22583);
xnor U23725 (N_23725,N_22015,N_22592);
nor U23726 (N_23726,N_21785,N_22685);
nor U23727 (N_23727,N_22345,N_21601);
nor U23728 (N_23728,N_22424,N_22147);
nor U23729 (N_23729,N_22113,N_22154);
and U23730 (N_23730,N_22013,N_21973);
xnor U23731 (N_23731,N_22424,N_21988);
or U23732 (N_23732,N_21820,N_21977);
nor U23733 (N_23733,N_22007,N_22287);
and U23734 (N_23734,N_22631,N_22539);
xor U23735 (N_23735,N_22401,N_22465);
xor U23736 (N_23736,N_22168,N_21807);
or U23737 (N_23737,N_21783,N_22069);
and U23738 (N_23738,N_22453,N_22125);
nor U23739 (N_23739,N_22288,N_22325);
and U23740 (N_23740,N_22118,N_22136);
nor U23741 (N_23741,N_22701,N_22418);
nor U23742 (N_23742,N_22659,N_21636);
nor U23743 (N_23743,N_22153,N_22581);
nand U23744 (N_23744,N_21639,N_22033);
xnor U23745 (N_23745,N_21851,N_22796);
nor U23746 (N_23746,N_22229,N_22334);
and U23747 (N_23747,N_22353,N_22108);
xor U23748 (N_23748,N_22007,N_22256);
nor U23749 (N_23749,N_22038,N_22569);
and U23750 (N_23750,N_22778,N_21773);
nand U23751 (N_23751,N_22027,N_22471);
xnor U23752 (N_23752,N_22062,N_22280);
and U23753 (N_23753,N_21638,N_21822);
nand U23754 (N_23754,N_22626,N_22194);
nor U23755 (N_23755,N_22184,N_22003);
xor U23756 (N_23756,N_21910,N_22121);
and U23757 (N_23757,N_22160,N_21776);
nor U23758 (N_23758,N_21770,N_22089);
and U23759 (N_23759,N_22604,N_21700);
or U23760 (N_23760,N_22518,N_21726);
nor U23761 (N_23761,N_22428,N_22693);
nor U23762 (N_23762,N_22799,N_22730);
and U23763 (N_23763,N_21974,N_22389);
or U23764 (N_23764,N_22535,N_21918);
or U23765 (N_23765,N_22632,N_21760);
and U23766 (N_23766,N_22149,N_21740);
xnor U23767 (N_23767,N_22666,N_21741);
or U23768 (N_23768,N_21935,N_22349);
nor U23769 (N_23769,N_22577,N_22329);
xnor U23770 (N_23770,N_22068,N_21715);
xnor U23771 (N_23771,N_22521,N_22514);
and U23772 (N_23772,N_22420,N_22089);
and U23773 (N_23773,N_22002,N_21625);
or U23774 (N_23774,N_21614,N_22069);
nor U23775 (N_23775,N_21624,N_22177);
xnor U23776 (N_23776,N_21617,N_21998);
or U23777 (N_23777,N_22101,N_21942);
nor U23778 (N_23778,N_22285,N_22202);
or U23779 (N_23779,N_22628,N_21633);
nand U23780 (N_23780,N_22590,N_22150);
and U23781 (N_23781,N_22396,N_21985);
nor U23782 (N_23782,N_22028,N_22186);
xnor U23783 (N_23783,N_22262,N_21723);
nand U23784 (N_23784,N_21663,N_22065);
and U23785 (N_23785,N_21841,N_22685);
nand U23786 (N_23786,N_22515,N_21968);
or U23787 (N_23787,N_22243,N_22212);
or U23788 (N_23788,N_22049,N_22085);
or U23789 (N_23789,N_22638,N_22587);
nand U23790 (N_23790,N_22013,N_22024);
nand U23791 (N_23791,N_21979,N_21911);
and U23792 (N_23792,N_22470,N_22212);
or U23793 (N_23793,N_22704,N_21653);
nor U23794 (N_23794,N_21866,N_22141);
nor U23795 (N_23795,N_22656,N_21675);
nand U23796 (N_23796,N_21985,N_22403);
nor U23797 (N_23797,N_22796,N_22547);
or U23798 (N_23798,N_22335,N_22150);
or U23799 (N_23799,N_21771,N_21667);
or U23800 (N_23800,N_21602,N_22530);
nor U23801 (N_23801,N_21745,N_21696);
or U23802 (N_23802,N_22462,N_22199);
or U23803 (N_23803,N_21761,N_22392);
or U23804 (N_23804,N_22071,N_22316);
nor U23805 (N_23805,N_21655,N_21912);
nand U23806 (N_23806,N_22758,N_22209);
nor U23807 (N_23807,N_21855,N_22383);
and U23808 (N_23808,N_21959,N_22778);
nand U23809 (N_23809,N_22349,N_22038);
xor U23810 (N_23810,N_22699,N_21684);
or U23811 (N_23811,N_21981,N_22798);
nor U23812 (N_23812,N_22680,N_22544);
or U23813 (N_23813,N_22627,N_21863);
or U23814 (N_23814,N_22658,N_21688);
or U23815 (N_23815,N_21841,N_21711);
nand U23816 (N_23816,N_22301,N_22771);
nor U23817 (N_23817,N_22604,N_22719);
or U23818 (N_23818,N_21969,N_22255);
and U23819 (N_23819,N_21679,N_21735);
nor U23820 (N_23820,N_21930,N_21924);
and U23821 (N_23821,N_22700,N_21912);
or U23822 (N_23822,N_22667,N_21607);
nor U23823 (N_23823,N_22406,N_22620);
nor U23824 (N_23824,N_21915,N_22061);
xor U23825 (N_23825,N_22011,N_22128);
and U23826 (N_23826,N_22292,N_22799);
or U23827 (N_23827,N_22047,N_22036);
or U23828 (N_23828,N_21709,N_21804);
nor U23829 (N_23829,N_21804,N_22510);
nor U23830 (N_23830,N_22551,N_22437);
xor U23831 (N_23831,N_22490,N_22154);
xor U23832 (N_23832,N_22224,N_21787);
nor U23833 (N_23833,N_22177,N_22068);
or U23834 (N_23834,N_22637,N_22554);
nand U23835 (N_23835,N_21769,N_22139);
and U23836 (N_23836,N_22588,N_22693);
and U23837 (N_23837,N_22326,N_22583);
xnor U23838 (N_23838,N_21956,N_21978);
or U23839 (N_23839,N_22714,N_22024);
and U23840 (N_23840,N_21964,N_22017);
and U23841 (N_23841,N_22760,N_21650);
xnor U23842 (N_23842,N_22710,N_22749);
or U23843 (N_23843,N_22312,N_22689);
nand U23844 (N_23844,N_22547,N_22169);
or U23845 (N_23845,N_22245,N_22748);
xor U23846 (N_23846,N_22201,N_22411);
xor U23847 (N_23847,N_22015,N_22406);
nand U23848 (N_23848,N_21761,N_22295);
or U23849 (N_23849,N_22023,N_22164);
xnor U23850 (N_23850,N_21975,N_22700);
xor U23851 (N_23851,N_22523,N_22724);
nand U23852 (N_23852,N_22734,N_22461);
nand U23853 (N_23853,N_21637,N_21968);
and U23854 (N_23854,N_21860,N_22519);
xnor U23855 (N_23855,N_21987,N_21743);
and U23856 (N_23856,N_22697,N_22404);
xor U23857 (N_23857,N_21959,N_22323);
and U23858 (N_23858,N_22727,N_22184);
or U23859 (N_23859,N_22184,N_22461);
xnor U23860 (N_23860,N_22579,N_21991);
or U23861 (N_23861,N_22681,N_22463);
or U23862 (N_23862,N_22747,N_22377);
nor U23863 (N_23863,N_22065,N_22044);
and U23864 (N_23864,N_22148,N_22673);
or U23865 (N_23865,N_22198,N_22052);
xnor U23866 (N_23866,N_22506,N_22687);
nand U23867 (N_23867,N_22341,N_21724);
or U23868 (N_23868,N_22127,N_22289);
xor U23869 (N_23869,N_21846,N_22705);
xnor U23870 (N_23870,N_21647,N_22069);
or U23871 (N_23871,N_21728,N_21641);
nor U23872 (N_23872,N_22388,N_22533);
nand U23873 (N_23873,N_22101,N_22390);
nand U23874 (N_23874,N_22432,N_22267);
xor U23875 (N_23875,N_22165,N_22624);
nor U23876 (N_23876,N_22553,N_22521);
or U23877 (N_23877,N_21813,N_22636);
nor U23878 (N_23878,N_22784,N_22071);
nand U23879 (N_23879,N_21773,N_21863);
xor U23880 (N_23880,N_22503,N_22130);
nor U23881 (N_23881,N_22283,N_22541);
nand U23882 (N_23882,N_21698,N_21811);
and U23883 (N_23883,N_22678,N_22123);
nand U23884 (N_23884,N_22147,N_22374);
and U23885 (N_23885,N_22039,N_22080);
and U23886 (N_23886,N_22590,N_21894);
xor U23887 (N_23887,N_22052,N_22091);
and U23888 (N_23888,N_22268,N_22199);
and U23889 (N_23889,N_22255,N_22077);
or U23890 (N_23890,N_21972,N_22327);
nand U23891 (N_23891,N_21835,N_22526);
or U23892 (N_23892,N_22543,N_22060);
xor U23893 (N_23893,N_21811,N_22730);
or U23894 (N_23894,N_22245,N_21884);
nand U23895 (N_23895,N_21821,N_22135);
nor U23896 (N_23896,N_22495,N_22100);
xnor U23897 (N_23897,N_22453,N_22744);
or U23898 (N_23898,N_22766,N_21762);
or U23899 (N_23899,N_22133,N_21786);
xor U23900 (N_23900,N_22746,N_22154);
nor U23901 (N_23901,N_22103,N_22592);
xor U23902 (N_23902,N_22013,N_22605);
nand U23903 (N_23903,N_22781,N_22764);
nor U23904 (N_23904,N_21788,N_22046);
or U23905 (N_23905,N_22136,N_21620);
or U23906 (N_23906,N_22245,N_21793);
nor U23907 (N_23907,N_21978,N_22608);
nand U23908 (N_23908,N_22308,N_22067);
xnor U23909 (N_23909,N_22658,N_22493);
xnor U23910 (N_23910,N_21946,N_22070);
nor U23911 (N_23911,N_21695,N_21600);
or U23912 (N_23912,N_21601,N_22484);
or U23913 (N_23913,N_21941,N_22115);
xor U23914 (N_23914,N_22119,N_22073);
nand U23915 (N_23915,N_22081,N_22030);
nor U23916 (N_23916,N_22746,N_21650);
nor U23917 (N_23917,N_22781,N_22229);
nor U23918 (N_23918,N_21767,N_22174);
nand U23919 (N_23919,N_22121,N_22249);
and U23920 (N_23920,N_21868,N_22297);
and U23921 (N_23921,N_22109,N_21854);
and U23922 (N_23922,N_22355,N_22474);
or U23923 (N_23923,N_22258,N_21608);
nor U23924 (N_23924,N_22419,N_22282);
and U23925 (N_23925,N_22517,N_22475);
xnor U23926 (N_23926,N_22613,N_21680);
nand U23927 (N_23927,N_22431,N_21871);
nand U23928 (N_23928,N_21895,N_22252);
or U23929 (N_23929,N_22524,N_22551);
or U23930 (N_23930,N_21707,N_22229);
nor U23931 (N_23931,N_21745,N_21729);
and U23932 (N_23932,N_21999,N_22270);
xor U23933 (N_23933,N_22098,N_21914);
or U23934 (N_23934,N_22566,N_21955);
xnor U23935 (N_23935,N_22363,N_22450);
nor U23936 (N_23936,N_22508,N_21954);
xnor U23937 (N_23937,N_22773,N_22292);
or U23938 (N_23938,N_21639,N_22776);
nand U23939 (N_23939,N_21949,N_22010);
xnor U23940 (N_23940,N_22513,N_22078);
nand U23941 (N_23941,N_22577,N_21789);
or U23942 (N_23942,N_21809,N_22766);
and U23943 (N_23943,N_21679,N_22334);
xnor U23944 (N_23944,N_22733,N_22626);
xnor U23945 (N_23945,N_22074,N_22360);
nor U23946 (N_23946,N_22625,N_22305);
or U23947 (N_23947,N_22670,N_22564);
and U23948 (N_23948,N_22544,N_21969);
and U23949 (N_23949,N_21892,N_22772);
or U23950 (N_23950,N_22272,N_21859);
or U23951 (N_23951,N_21614,N_22638);
nor U23952 (N_23952,N_21813,N_22277);
xnor U23953 (N_23953,N_22565,N_22282);
xor U23954 (N_23954,N_22252,N_21723);
nor U23955 (N_23955,N_22058,N_22701);
xor U23956 (N_23956,N_22758,N_22426);
or U23957 (N_23957,N_22132,N_21958);
xor U23958 (N_23958,N_22069,N_22486);
and U23959 (N_23959,N_21976,N_21673);
or U23960 (N_23960,N_22159,N_22572);
and U23961 (N_23961,N_22619,N_22262);
nor U23962 (N_23962,N_22572,N_22506);
nand U23963 (N_23963,N_21773,N_22713);
or U23964 (N_23964,N_22081,N_21995);
xnor U23965 (N_23965,N_21840,N_21758);
nand U23966 (N_23966,N_21976,N_22237);
xor U23967 (N_23967,N_22117,N_22751);
or U23968 (N_23968,N_21945,N_21983);
xnor U23969 (N_23969,N_21745,N_22608);
or U23970 (N_23970,N_21646,N_22041);
nand U23971 (N_23971,N_22537,N_22247);
or U23972 (N_23972,N_22221,N_21970);
or U23973 (N_23973,N_21736,N_21884);
nor U23974 (N_23974,N_22079,N_21853);
nand U23975 (N_23975,N_22223,N_21722);
nor U23976 (N_23976,N_22761,N_22684);
and U23977 (N_23977,N_22352,N_22740);
and U23978 (N_23978,N_21765,N_22506);
xnor U23979 (N_23979,N_21755,N_21929);
and U23980 (N_23980,N_21724,N_22608);
xor U23981 (N_23981,N_21997,N_22773);
nor U23982 (N_23982,N_21636,N_22065);
and U23983 (N_23983,N_22435,N_21612);
nor U23984 (N_23984,N_22186,N_21935);
or U23985 (N_23985,N_22457,N_21658);
xor U23986 (N_23986,N_22396,N_21799);
and U23987 (N_23987,N_22205,N_22105);
nor U23988 (N_23988,N_21641,N_21984);
nor U23989 (N_23989,N_22081,N_22150);
xor U23990 (N_23990,N_22037,N_22289);
or U23991 (N_23991,N_21898,N_22634);
nand U23992 (N_23992,N_22111,N_21683);
and U23993 (N_23993,N_22119,N_22345);
nand U23994 (N_23994,N_22033,N_22198);
and U23995 (N_23995,N_22539,N_22325);
nor U23996 (N_23996,N_22489,N_22511);
and U23997 (N_23997,N_22682,N_21806);
nor U23998 (N_23998,N_22107,N_21659);
and U23999 (N_23999,N_22386,N_22729);
xnor U24000 (N_24000,N_23862,N_23275);
and U24001 (N_24001,N_23786,N_23751);
nor U24002 (N_24002,N_23288,N_23908);
nor U24003 (N_24003,N_23363,N_23007);
nor U24004 (N_24004,N_23216,N_23134);
nand U24005 (N_24005,N_23925,N_23434);
xnor U24006 (N_24006,N_23082,N_23579);
xnor U24007 (N_24007,N_22936,N_23924);
and U24008 (N_24008,N_23826,N_23109);
nand U24009 (N_24009,N_23457,N_23191);
and U24010 (N_24010,N_23237,N_22989);
nor U24011 (N_24011,N_23310,N_23565);
nor U24012 (N_24012,N_23196,N_22933);
nor U24013 (N_24013,N_23845,N_23651);
nor U24014 (N_24014,N_23367,N_22822);
or U24015 (N_24015,N_23108,N_23125);
xnor U24016 (N_24016,N_22973,N_23614);
or U24017 (N_24017,N_23485,N_23267);
or U24018 (N_24018,N_23951,N_23365);
nand U24019 (N_24019,N_22957,N_23509);
and U24020 (N_24020,N_23088,N_23936);
and U24021 (N_24021,N_23830,N_22921);
nand U24022 (N_24022,N_23374,N_23020);
or U24023 (N_24023,N_22984,N_23624);
xor U24024 (N_24024,N_22892,N_23915);
or U24025 (N_24025,N_22820,N_23793);
or U24026 (N_24026,N_23084,N_23206);
xnor U24027 (N_24027,N_23824,N_23145);
and U24028 (N_24028,N_23256,N_23211);
and U24029 (N_24029,N_23037,N_23320);
xnor U24030 (N_24030,N_23203,N_23343);
and U24031 (N_24031,N_23164,N_23791);
or U24032 (N_24032,N_23946,N_23055);
or U24033 (N_24033,N_23980,N_22879);
or U24034 (N_24034,N_22849,N_23159);
nor U24035 (N_24035,N_23494,N_23723);
or U24036 (N_24036,N_23212,N_23431);
or U24037 (N_24037,N_23883,N_23876);
or U24038 (N_24038,N_23905,N_23198);
nor U24039 (N_24039,N_23248,N_23810);
nand U24040 (N_24040,N_22859,N_22944);
and U24041 (N_24041,N_23694,N_23874);
and U24042 (N_24042,N_23429,N_23419);
nand U24043 (N_24043,N_23536,N_23776);
xnor U24044 (N_24044,N_23403,N_23263);
nor U24045 (N_24045,N_23653,N_23903);
and U24046 (N_24046,N_23843,N_23337);
nor U24047 (N_24047,N_23714,N_23075);
xnor U24048 (N_24048,N_22929,N_23650);
nand U24049 (N_24049,N_23846,N_23923);
xnor U24050 (N_24050,N_22874,N_23617);
or U24051 (N_24051,N_23993,N_23062);
xnor U24052 (N_24052,N_22922,N_23249);
nand U24053 (N_24053,N_23455,N_23024);
nand U24054 (N_24054,N_23604,N_23214);
nor U24055 (N_24055,N_23978,N_23551);
and U24056 (N_24056,N_22814,N_23478);
or U24057 (N_24057,N_23398,N_22997);
xor U24058 (N_24058,N_23931,N_22927);
or U24059 (N_24059,N_23736,N_22812);
nand U24060 (N_24060,N_23277,N_23641);
xor U24061 (N_24061,N_22888,N_23972);
and U24062 (N_24062,N_23576,N_22991);
nand U24063 (N_24063,N_23050,N_23748);
or U24064 (N_24064,N_23065,N_23852);
nand U24065 (N_24065,N_22924,N_22817);
and U24066 (N_24066,N_22899,N_23882);
nor U24067 (N_24067,N_23500,N_22966);
nor U24068 (N_24068,N_23526,N_23264);
or U24069 (N_24069,N_22914,N_23864);
xor U24070 (N_24070,N_23302,N_23807);
or U24071 (N_24071,N_23013,N_23195);
and U24072 (N_24072,N_23632,N_22951);
nand U24073 (N_24073,N_23290,N_23008);
xor U24074 (N_24074,N_23954,N_23785);
or U24075 (N_24075,N_23546,N_22902);
nor U24076 (N_24076,N_23016,N_23540);
or U24077 (N_24077,N_23691,N_22836);
xnor U24078 (N_24078,N_23352,N_23401);
or U24079 (N_24079,N_23067,N_23340);
and U24080 (N_24080,N_23459,N_23577);
nor U24081 (N_24081,N_23230,N_23667);
nor U24082 (N_24082,N_22808,N_23964);
xnor U24083 (N_24083,N_23628,N_22988);
and U24084 (N_24084,N_23996,N_23312);
nand U24085 (N_24085,N_23848,N_22915);
xor U24086 (N_24086,N_23440,N_22815);
or U24087 (N_24087,N_23180,N_23407);
and U24088 (N_24088,N_23507,N_23997);
nand U24089 (N_24089,N_23122,N_22947);
xnor U24090 (N_24090,N_23974,N_22945);
and U24091 (N_24091,N_22845,N_23814);
and U24092 (N_24092,N_22930,N_23520);
and U24093 (N_24093,N_23270,N_23127);
nor U24094 (N_24094,N_23589,N_23816);
nand U24095 (N_24095,N_23737,N_23408);
nor U24096 (N_24096,N_22940,N_23592);
or U24097 (N_24097,N_23866,N_23095);
nand U24098 (N_24098,N_23409,N_23378);
and U24099 (N_24099,N_22829,N_22956);
nor U24100 (N_24100,N_23101,N_23178);
and U24101 (N_24101,N_22979,N_23514);
nand U24102 (N_24102,N_23911,N_23770);
or U24103 (N_24103,N_23413,N_23734);
and U24104 (N_24104,N_23420,N_22962);
nand U24105 (N_24105,N_23949,N_22861);
or U24106 (N_24106,N_23029,N_22972);
and U24107 (N_24107,N_23053,N_23492);
xor U24108 (N_24108,N_23342,N_23451);
or U24109 (N_24109,N_23228,N_23059);
and U24110 (N_24110,N_23727,N_23498);
nand U24111 (N_24111,N_23435,N_23182);
or U24112 (N_24112,N_23747,N_23556);
nand U24113 (N_24113,N_23684,N_23966);
and U24114 (N_24114,N_23271,N_23390);
nor U24115 (N_24115,N_23875,N_22967);
nor U24116 (N_24116,N_23427,N_23539);
nor U24117 (N_24117,N_23806,N_23620);
or U24118 (N_24118,N_23855,N_23238);
and U24119 (N_24119,N_22865,N_23326);
and U24120 (N_24120,N_23932,N_23803);
xnor U24121 (N_24121,N_23040,N_23332);
nand U24122 (N_24122,N_22877,N_23857);
and U24123 (N_24123,N_22838,N_23150);
nor U24124 (N_24124,N_23917,N_23276);
or U24125 (N_24125,N_23169,N_23242);
or U24126 (N_24126,N_23510,N_23126);
and U24127 (N_24127,N_22863,N_22906);
or U24128 (N_24128,N_22913,N_23464);
or U24129 (N_24129,N_23496,N_23381);
nand U24130 (N_24130,N_23718,N_23710);
or U24131 (N_24131,N_23597,N_23475);
xnor U24132 (N_24132,N_23382,N_23143);
and U24133 (N_24133,N_23041,N_23690);
and U24134 (N_24134,N_23023,N_22975);
xnor U24135 (N_24135,N_22942,N_23517);
or U24136 (N_24136,N_23422,N_23662);
or U24137 (N_24137,N_23328,N_23295);
nor U24138 (N_24138,N_23351,N_23851);
xor U24139 (N_24139,N_23397,N_22918);
or U24140 (N_24140,N_22923,N_23490);
xor U24141 (N_24141,N_23686,N_23891);
nand U24142 (N_24142,N_23387,N_22847);
nor U24143 (N_24143,N_23591,N_23912);
nor U24144 (N_24144,N_23032,N_22883);
and U24145 (N_24145,N_23813,N_23133);
or U24146 (N_24146,N_23282,N_23977);
nand U24147 (N_24147,N_23140,N_23835);
or U24148 (N_24148,N_23713,N_23728);
xnor U24149 (N_24149,N_23942,N_22809);
and U24150 (N_24150,N_23116,N_23439);
and U24151 (N_24151,N_23399,N_23601);
and U24152 (N_24152,N_23889,N_23784);
nor U24153 (N_24153,N_23341,N_23179);
and U24154 (N_24154,N_22968,N_22981);
or U24155 (N_24155,N_23453,N_23112);
nor U24156 (N_24156,N_22810,N_23961);
nor U24157 (N_24157,N_23550,N_23354);
xor U24158 (N_24158,N_23504,N_23314);
or U24159 (N_24159,N_23028,N_23102);
or U24160 (N_24160,N_23789,N_23994);
or U24161 (N_24161,N_23202,N_23670);
nor U24162 (N_24162,N_23877,N_23898);
nand U24163 (N_24163,N_23637,N_23749);
and U24164 (N_24164,N_22803,N_22931);
or U24165 (N_24165,N_23247,N_23554);
nor U24166 (N_24166,N_23372,N_23036);
xor U24167 (N_24167,N_23255,N_23741);
or U24168 (N_24168,N_22807,N_22986);
or U24169 (N_24169,N_23658,N_23618);
nand U24170 (N_24170,N_23045,N_23769);
nor U24171 (N_24171,N_23516,N_22985);
nand U24172 (N_24172,N_23735,N_23965);
nand U24173 (N_24173,N_23787,N_23750);
nor U24174 (N_24174,N_23009,N_23957);
nand U24175 (N_24175,N_22959,N_23757);
or U24176 (N_24176,N_22909,N_23103);
xnor U24177 (N_24177,N_22891,N_23582);
or U24178 (N_24178,N_23183,N_22998);
or U24179 (N_24179,N_23406,N_23521);
and U24180 (N_24180,N_23031,N_23742);
or U24181 (N_24181,N_23569,N_23437);
xnor U24182 (N_24182,N_23677,N_23782);
xor U24183 (N_24183,N_22955,N_23347);
or U24184 (N_24184,N_22920,N_23501);
and U24185 (N_24185,N_23884,N_23473);
nor U24186 (N_24186,N_23623,N_23405);
or U24187 (N_24187,N_23168,N_23380);
or U24188 (N_24188,N_23330,N_22885);
xnor U24189 (N_24189,N_23357,N_23469);
nor U24190 (N_24190,N_23336,N_22905);
or U24191 (N_24191,N_23708,N_23812);
xor U24192 (N_24192,N_23064,N_23269);
or U24193 (N_24193,N_23232,N_23079);
or U24194 (N_24194,N_23881,N_22974);
xnor U24195 (N_24195,N_23926,N_23331);
nand U24196 (N_24196,N_22965,N_23960);
nand U24197 (N_24197,N_23615,N_23385);
nor U24198 (N_24198,N_23110,N_23892);
nand U24199 (N_24199,N_22848,N_23513);
nand U24200 (N_24200,N_23557,N_23066);
nor U24201 (N_24201,N_23467,N_23743);
nand U24202 (N_24202,N_23729,N_23304);
and U24203 (N_24203,N_23488,N_23430);
and U24204 (N_24204,N_23188,N_23524);
or U24205 (N_24205,N_23758,N_23364);
nand U24206 (N_24206,N_23493,N_23860);
and U24207 (N_24207,N_23480,N_23679);
nand U24208 (N_24208,N_23698,N_23976);
xnor U24209 (N_24209,N_23004,N_23091);
and U24210 (N_24210,N_23847,N_22987);
and U24211 (N_24211,N_23483,N_23224);
and U24212 (N_24212,N_22978,N_23362);
or U24213 (N_24213,N_23135,N_23764);
nand U24214 (N_24214,N_23703,N_22939);
xnor U24215 (N_24215,N_23280,N_23098);
xor U24216 (N_24216,N_23260,N_23265);
and U24217 (N_24217,N_23731,N_23808);
xnor U24218 (N_24218,N_23074,N_23804);
xor U24219 (N_24219,N_23291,N_23285);
and U24220 (N_24220,N_23619,N_23479);
and U24221 (N_24221,N_23610,N_23712);
and U24222 (N_24222,N_23542,N_23535);
and U24223 (N_24223,N_23210,N_23021);
xor U24224 (N_24224,N_23730,N_23940);
nor U24225 (N_24225,N_23121,N_23279);
nand U24226 (N_24226,N_22823,N_23571);
xor U24227 (N_24227,N_22977,N_23896);
nand U24228 (N_24228,N_23096,N_23201);
xnor U24229 (N_24229,N_23069,N_23695);
xor U24230 (N_24230,N_23154,N_23722);
and U24231 (N_24231,N_23689,N_23167);
nor U24232 (N_24232,N_23950,N_23828);
and U24233 (N_24233,N_22843,N_23715);
xnor U24234 (N_24234,N_22867,N_23880);
xnor U24235 (N_24235,N_23570,N_23990);
and U24236 (N_24236,N_23945,N_23692);
nor U24237 (N_24237,N_23660,N_23989);
nand U24238 (N_24238,N_23389,N_23057);
xnor U24239 (N_24239,N_22811,N_23600);
or U24240 (N_24240,N_23815,N_23350);
nand U24241 (N_24241,N_23172,N_23305);
xnor U24242 (N_24242,N_23035,N_23001);
nand U24243 (N_24243,N_23481,N_23308);
nor U24244 (N_24244,N_23158,N_23083);
nand U24245 (N_24245,N_23334,N_23811);
and U24246 (N_24246,N_23197,N_23837);
and U24247 (N_24247,N_23709,N_23893);
and U24248 (N_24248,N_22844,N_22887);
xor U24249 (N_24249,N_23596,N_23680);
nor U24250 (N_24250,N_23253,N_23243);
nand U24251 (N_24251,N_23717,N_23348);
and U24252 (N_24252,N_23186,N_23117);
nand U24253 (N_24253,N_23250,N_23400);
and U24254 (N_24254,N_23744,N_23929);
nor U24255 (N_24255,N_23258,N_22964);
and U24256 (N_24256,N_23138,N_23338);
xor U24257 (N_24257,N_23817,N_23652);
xor U24258 (N_24258,N_23583,N_23073);
and U24259 (N_24259,N_23773,N_23227);
nor U24260 (N_24260,N_23704,N_23987);
or U24261 (N_24261,N_22880,N_23026);
nand U24262 (N_24262,N_23732,N_22841);
xnor U24263 (N_24263,N_22871,N_22969);
or U24264 (N_24264,N_23199,N_22901);
nand U24265 (N_24265,N_23969,N_23752);
xnor U24266 (N_24266,N_23840,N_23044);
nor U24267 (N_24267,N_23598,N_23502);
nor U24268 (N_24268,N_23130,N_23661);
and U24269 (N_24269,N_23349,N_23106);
or U24270 (N_24270,N_23962,N_23913);
nand U24271 (N_24271,N_23886,N_23858);
and U24272 (N_24272,N_23878,N_22916);
or U24273 (N_24273,N_23656,N_22800);
or U24274 (N_24274,N_23933,N_23373);
xnor U24275 (N_24275,N_23834,N_23952);
nand U24276 (N_24276,N_23584,N_23417);
nand U24277 (N_24277,N_23992,N_23754);
nand U24278 (N_24278,N_23809,N_23111);
xor U24279 (N_24279,N_23200,N_23937);
nand U24280 (N_24280,N_23284,N_23297);
nor U24281 (N_24281,N_23534,N_23625);
and U24282 (N_24282,N_23027,N_22805);
nand U24283 (N_24283,N_23985,N_23982);
or U24284 (N_24284,N_23426,N_23772);
or U24285 (N_24285,N_23185,N_23823);
nor U24286 (N_24286,N_23124,N_23825);
or U24287 (N_24287,N_23162,N_23423);
xor U24288 (N_24288,N_23468,N_23450);
and U24289 (N_24289,N_23017,N_22903);
or U24290 (N_24290,N_23466,N_23697);
nor U24291 (N_24291,N_23240,N_23902);
xnor U24292 (N_24292,N_22819,N_23533);
and U24293 (N_24293,N_23085,N_23051);
or U24294 (N_24294,N_22853,N_23100);
or U24295 (N_24295,N_22864,N_22941);
xnor U24296 (N_24296,N_23543,N_23899);
or U24297 (N_24297,N_23165,N_23904);
xor U24298 (N_24298,N_23963,N_23801);
and U24299 (N_24299,N_23244,N_23463);
nor U24300 (N_24300,N_23089,N_23170);
nand U24301 (N_24301,N_23799,N_23246);
xnor U24302 (N_24302,N_23916,N_23360);
xnor U24303 (N_24303,N_22976,N_23425);
and U24304 (N_24304,N_23161,N_23292);
and U24305 (N_24305,N_23506,N_23668);
xnor U24306 (N_24306,N_22821,N_22983);
xnor U24307 (N_24307,N_23287,N_23000);
and U24308 (N_24308,N_23574,N_23943);
nand U24309 (N_24309,N_23766,N_23266);
or U24310 (N_24310,N_22850,N_23907);
and U24311 (N_24311,N_23011,N_23345);
nor U24312 (N_24312,N_22866,N_22961);
nand U24313 (N_24313,N_23975,N_23396);
nor U24314 (N_24314,N_23298,N_22881);
nor U24315 (N_24315,N_23118,N_23669);
nor U24316 (N_24316,N_23433,N_23633);
xnor U24317 (N_24317,N_23339,N_23208);
or U24318 (N_24318,N_23094,N_23671);
nor U24319 (N_24319,N_22872,N_23289);
and U24320 (N_24320,N_23887,N_22895);
nor U24321 (N_24321,N_23831,N_23317);
xor U24322 (N_24322,N_23410,N_23636);
and U24323 (N_24323,N_23645,N_23152);
nand U24324 (N_24324,N_22889,N_23300);
and U24325 (N_24325,N_23802,N_23225);
nor U24326 (N_24326,N_23261,N_23820);
or U24327 (N_24327,N_23080,N_23153);
and U24328 (N_24328,N_23113,N_23296);
xor U24329 (N_24329,N_23696,N_22862);
nor U24330 (N_24330,N_23315,N_23586);
nand U24331 (N_24331,N_23002,N_22897);
and U24332 (N_24332,N_23958,N_22952);
xor U24333 (N_24333,N_23092,N_23299);
and U24334 (N_24334,N_23181,N_23048);
nor U24335 (N_24335,N_23449,N_23622);
nand U24336 (N_24336,N_23254,N_23104);
and U24337 (N_24337,N_23497,N_23593);
nor U24338 (N_24338,N_22935,N_23909);
nor U24339 (N_24339,N_23528,N_23587);
nor U24340 (N_24340,N_23523,N_23190);
or U24341 (N_24341,N_23944,N_23647);
or U24342 (N_24342,N_23685,N_23272);
or U24343 (N_24343,N_23595,N_23724);
and U24344 (N_24344,N_22801,N_23303);
and U24345 (N_24345,N_23086,N_23829);
nand U24346 (N_24346,N_23719,N_23678);
and U24347 (N_24347,N_23664,N_22834);
and U24348 (N_24348,N_23914,N_23527);
and U24349 (N_24349,N_23355,N_23832);
nand U24350 (N_24350,N_22857,N_22953);
nand U24351 (N_24351,N_23640,N_23682);
xor U24352 (N_24352,N_23762,N_23229);
or U24353 (N_24353,N_23155,N_22831);
nor U24354 (N_24354,N_23885,N_23765);
and U24355 (N_24355,N_23935,N_23959);
or U24356 (N_24356,N_23967,N_23612);
and U24357 (N_24357,N_23683,N_23879);
nor U24358 (N_24358,N_23968,N_23755);
nand U24359 (N_24359,N_23491,N_23444);
nand U24360 (N_24360,N_23672,N_23953);
nor U24361 (N_24361,N_23115,N_23311);
xor U24362 (N_24362,N_23177,N_23646);
nor U24363 (N_24363,N_23033,N_22904);
nor U24364 (N_24364,N_23489,N_23499);
nand U24365 (N_24365,N_23821,N_23239);
nand U24366 (N_24366,N_23532,N_23827);
nor U24367 (N_24367,N_23090,N_23235);
and U24368 (N_24368,N_23128,N_23204);
nand U24369 (N_24369,N_23441,N_23505);
nor U24370 (N_24370,N_23215,N_23659);
nand U24371 (N_24371,N_23839,N_22900);
nand U24372 (N_24372,N_23983,N_22928);
nand U24373 (N_24373,N_23642,N_23148);
xnor U24374 (N_24374,N_23868,N_22886);
and U24375 (N_24375,N_23323,N_23301);
and U24376 (N_24376,N_23054,N_23262);
or U24377 (N_24377,N_23564,N_23870);
nor U24378 (N_24378,N_22934,N_23316);
or U24379 (N_24379,N_23166,N_23231);
xnor U24380 (N_24380,N_23687,N_23581);
and U24381 (N_24381,N_23973,N_23906);
or U24382 (N_24382,N_23460,N_23139);
nor U24383 (N_24383,N_23699,N_23721);
or U24384 (N_24384,N_23850,N_22893);
nor U24385 (N_24385,N_23395,N_23321);
or U24386 (N_24386,N_23105,N_23391);
and U24387 (N_24387,N_23495,N_23412);
nor U24388 (N_24388,N_22894,N_23344);
and U24389 (N_24389,N_23043,N_23222);
or U24390 (N_24390,N_23572,N_23512);
or U24391 (N_24391,N_23529,N_22898);
xnor U24392 (N_24392,N_22846,N_22937);
and U24393 (N_24393,N_23049,N_22832);
and U24394 (N_24394,N_23818,N_23606);
nor U24395 (N_24395,N_22996,N_23998);
nor U24396 (N_24396,N_23871,N_23761);
nand U24397 (N_24397,N_23218,N_23307);
xnor U24398 (N_24398,N_23800,N_23462);
nand U24399 (N_24399,N_22828,N_23482);
nand U24400 (N_24400,N_23654,N_23010);
and U24401 (N_24401,N_23281,N_22982);
nor U24402 (N_24402,N_23873,N_23187);
nand U24403 (N_24403,N_23627,N_23702);
nand U24404 (N_24404,N_23071,N_23418);
nand U24405 (N_24405,N_23955,N_23771);
xor U24406 (N_24406,N_23783,N_23038);
and U24407 (N_24407,N_23484,N_23384);
nor U24408 (N_24408,N_23921,N_23649);
nand U24409 (N_24409,N_23836,N_23798);
and U24410 (N_24410,N_23580,N_23184);
nand U24411 (N_24411,N_23077,N_23209);
nor U24412 (N_24412,N_23665,N_23366);
or U24413 (N_24413,N_23626,N_23558);
and U24414 (N_24414,N_23555,N_23644);
nand U24415 (N_24415,N_23402,N_23849);
nand U24416 (N_24416,N_22840,N_23676);
and U24417 (N_24417,N_23888,N_23538);
nor U24418 (N_24418,N_23566,N_23988);
xor U24419 (N_24419,N_23777,N_23778);
or U24420 (N_24420,N_23171,N_23854);
and U24421 (N_24421,N_23072,N_23356);
or U24422 (N_24422,N_22873,N_23971);
nor U24423 (N_24423,N_23192,N_23233);
or U24424 (N_24424,N_22908,N_23530);
xnor U24425 (N_24425,N_23445,N_23745);
nor U24426 (N_24426,N_23221,N_23226);
and U24427 (N_24427,N_23394,N_23869);
or U24428 (N_24428,N_23223,N_23438);
nor U24429 (N_24429,N_23099,N_23984);
or U24430 (N_24430,N_23213,N_23386);
nor U24431 (N_24431,N_23613,N_23369);
and U24432 (N_24432,N_22860,N_23779);
or U24433 (N_24433,N_22851,N_22912);
or U24434 (N_24434,N_23415,N_22995);
nand U24435 (N_24435,N_23609,N_23070);
or U24436 (N_24436,N_23286,N_23383);
and U24437 (N_24437,N_23442,N_23819);
nor U24438 (N_24438,N_23531,N_23544);
xnor U24439 (N_24439,N_23207,N_23022);
xnor U24440 (N_24440,N_23052,N_23910);
and U24441 (N_24441,N_23970,N_23432);
xor U24442 (N_24442,N_23194,N_23144);
or U24443 (N_24443,N_23093,N_23900);
and U24444 (N_24444,N_23327,N_23377);
xnor U24445 (N_24445,N_23930,N_23563);
or U24446 (N_24446,N_23081,N_23019);
nand U24447 (N_24447,N_23547,N_23018);
and U24448 (N_24448,N_23928,N_23657);
xnor U24449 (N_24449,N_22875,N_23567);
nor U24450 (N_24450,N_23278,N_23634);
xnor U24451 (N_24451,N_23309,N_23608);
or U24452 (N_24452,N_23322,N_23294);
or U24453 (N_24453,N_23141,N_23436);
nand U24454 (N_24454,N_23999,N_23794);
and U24455 (N_24455,N_23841,N_22950);
nand U24456 (N_24456,N_23795,N_23805);
xor U24457 (N_24457,N_23313,N_22833);
xor U24458 (N_24458,N_23947,N_23456);
xor U24459 (N_24459,N_23443,N_23060);
nand U24460 (N_24460,N_22806,N_23895);
or U24461 (N_24461,N_23346,N_23585);
nor U24462 (N_24462,N_23371,N_23424);
and U24463 (N_24463,N_23726,N_23941);
or U24464 (N_24464,N_23353,N_23447);
nand U24465 (N_24465,N_23867,N_23979);
nand U24466 (N_24466,N_23790,N_23068);
and U24467 (N_24467,N_23552,N_23607);
xor U24468 (N_24468,N_23701,N_23132);
or U24469 (N_24469,N_22946,N_22980);
nand U24470 (N_24470,N_23006,N_23861);
xor U24471 (N_24471,N_23087,N_23594);
and U24472 (N_24472,N_23919,N_23688);
and U24473 (N_24473,N_23123,N_23939);
xnor U24474 (N_24474,N_23251,N_23590);
nor U24475 (N_24475,N_23934,N_23446);
xnor U24476 (N_24476,N_22890,N_23545);
nor U24477 (N_24477,N_23205,N_23780);
xnor U24478 (N_24478,N_22839,N_23176);
xnor U24479 (N_24479,N_23030,N_23245);
nor U24480 (N_24480,N_23560,N_23525);
nand U24481 (N_24481,N_23515,N_23631);
nand U24482 (N_24482,N_23666,N_22990);
xor U24483 (N_24483,N_23897,N_23901);
or U24484 (N_24484,N_23421,N_23486);
xor U24485 (N_24485,N_22994,N_23120);
and U24486 (N_24486,N_23042,N_23872);
and U24487 (N_24487,N_23471,N_23306);
and U24488 (N_24488,N_22963,N_23760);
xor U24489 (N_24489,N_23781,N_23474);
nand U24490 (N_24490,N_23142,N_23217);
and U24491 (N_24491,N_22856,N_23706);
nand U24492 (N_24492,N_23890,N_23605);
nand U24493 (N_24493,N_23163,N_23548);
and U24494 (N_24494,N_23693,N_23853);
or U24495 (N_24495,N_23611,N_23711);
nand U24496 (N_24496,N_23241,N_22858);
nor U24497 (N_24497,N_23648,N_23157);
or U24498 (N_24498,N_22910,N_23136);
xor U24499 (N_24499,N_23325,N_23477);
or U24500 (N_24500,N_23005,N_22813);
and U24501 (N_24501,N_23918,N_23025);
nor U24502 (N_24502,N_23234,N_23573);
or U24503 (N_24503,N_23675,N_23274);
or U24504 (N_24504,N_23797,N_22917);
xor U24505 (N_24505,N_23324,N_23599);
xor U24506 (N_24506,N_23537,N_23511);
nor U24507 (N_24507,N_23461,N_23716);
nor U24508 (N_24508,N_23268,N_23920);
nor U24509 (N_24509,N_23114,N_22919);
nor U24510 (N_24510,N_23193,N_23635);
xor U24511 (N_24511,N_23151,N_23472);
nand U24512 (N_24512,N_23333,N_22884);
xnor U24513 (N_24513,N_23220,N_23404);
and U24514 (N_24514,N_23707,N_23519);
xnor U24515 (N_24515,N_23375,N_23379);
nor U24516 (N_24516,N_23061,N_23189);
and U24517 (N_24517,N_23173,N_23639);
and U24518 (N_24518,N_22868,N_22999);
or U24519 (N_24519,N_23470,N_23518);
or U24520 (N_24520,N_23562,N_23259);
nor U24521 (N_24521,N_22911,N_23725);
xnor U24522 (N_24522,N_23318,N_23131);
xor U24523 (N_24523,N_23047,N_23454);
and U24524 (N_24524,N_23012,N_23465);
or U24525 (N_24525,N_23014,N_23865);
and U24526 (N_24526,N_23575,N_23578);
xor U24527 (N_24527,N_23046,N_23856);
xnor U24528 (N_24528,N_23995,N_23863);
nor U24529 (N_24529,N_23938,N_23767);
and U24530 (N_24530,N_23549,N_23948);
nor U24531 (N_24531,N_23700,N_22971);
or U24532 (N_24532,N_23621,N_23522);
xor U24533 (N_24533,N_22855,N_23107);
and U24534 (N_24534,N_23559,N_22925);
xnor U24535 (N_24535,N_23759,N_23147);
nor U24536 (N_24536,N_23319,N_23361);
nor U24537 (N_24537,N_22835,N_23986);
xor U24538 (N_24538,N_22958,N_23753);
and U24539 (N_24539,N_23561,N_23137);
xor U24540 (N_24540,N_23359,N_23738);
nand U24541 (N_24541,N_23844,N_23015);
nand U24542 (N_24542,N_23388,N_23927);
nand U24543 (N_24543,N_23788,N_22954);
or U24544 (N_24544,N_23175,N_23894);
xor U24545 (N_24545,N_23775,N_23792);
or U24546 (N_24546,N_22878,N_23981);
and U24547 (N_24547,N_22992,N_23416);
nor U24548 (N_24548,N_23039,N_22960);
nand U24549 (N_24549,N_23156,N_23003);
and U24550 (N_24550,N_23842,N_23219);
nor U24551 (N_24551,N_23746,N_22818);
nor U24552 (N_24552,N_23655,N_23956);
nand U24553 (N_24553,N_22830,N_22938);
nor U24554 (N_24554,N_23739,N_23283);
nor U24555 (N_24555,N_23119,N_22825);
nand U24556 (N_24556,N_23063,N_23756);
xor U24557 (N_24557,N_22802,N_22852);
and U24558 (N_24558,N_22870,N_22816);
xor U24559 (N_24559,N_22907,N_23273);
xnor U24560 (N_24560,N_23673,N_23146);
nor U24561 (N_24561,N_23588,N_23740);
or U24562 (N_24562,N_23922,N_23160);
or U24563 (N_24563,N_22876,N_23058);
or U24564 (N_24564,N_23392,N_23293);
nor U24565 (N_24565,N_23733,N_23822);
nor U24566 (N_24566,N_23428,N_22842);
xnor U24567 (N_24567,N_23411,N_23838);
or U24568 (N_24568,N_23078,N_23638);
and U24569 (N_24569,N_23257,N_23768);
or U24570 (N_24570,N_23368,N_22943);
xnor U24571 (N_24571,N_22932,N_23663);
nor U24572 (N_24572,N_23376,N_23487);
nand U24573 (N_24573,N_23252,N_22869);
or U24574 (N_24574,N_23503,N_23174);
nor U24575 (N_24575,N_23358,N_23076);
and U24576 (N_24576,N_22949,N_22826);
and U24577 (N_24577,N_22970,N_23681);
xor U24578 (N_24578,N_23393,N_23458);
nor U24579 (N_24579,N_22993,N_23508);
xor U24580 (N_24580,N_23629,N_23603);
nor U24581 (N_24581,N_23452,N_23705);
and U24582 (N_24582,N_23859,N_23720);
nor U24583 (N_24583,N_22926,N_22824);
nand U24584 (N_24584,N_23149,N_22896);
xnor U24585 (N_24585,N_23476,N_23643);
xor U24586 (N_24586,N_22854,N_23414);
nor U24587 (N_24587,N_23034,N_23763);
nor U24588 (N_24588,N_23448,N_23991);
or U24589 (N_24589,N_23553,N_23630);
nor U24590 (N_24590,N_23370,N_23097);
and U24591 (N_24591,N_23236,N_22827);
nor U24592 (N_24592,N_22882,N_23056);
xnor U24593 (N_24593,N_23602,N_22804);
or U24594 (N_24594,N_22837,N_23774);
or U24595 (N_24595,N_23833,N_23335);
and U24596 (N_24596,N_23674,N_23568);
or U24597 (N_24597,N_23796,N_22948);
or U24598 (N_24598,N_23541,N_23129);
nor U24599 (N_24599,N_23329,N_23616);
or U24600 (N_24600,N_23209,N_23892);
nand U24601 (N_24601,N_22933,N_22890);
nor U24602 (N_24602,N_22927,N_22924);
or U24603 (N_24603,N_23957,N_23872);
or U24604 (N_24604,N_23999,N_23740);
and U24605 (N_24605,N_23282,N_23341);
and U24606 (N_24606,N_23307,N_23109);
nand U24607 (N_24607,N_22853,N_23363);
nor U24608 (N_24608,N_23053,N_23167);
and U24609 (N_24609,N_23103,N_23447);
xnor U24610 (N_24610,N_23961,N_23371);
and U24611 (N_24611,N_23306,N_22971);
nand U24612 (N_24612,N_22948,N_23970);
and U24613 (N_24613,N_23185,N_23954);
nor U24614 (N_24614,N_22961,N_23821);
xnor U24615 (N_24615,N_23234,N_23178);
or U24616 (N_24616,N_23985,N_22872);
xnor U24617 (N_24617,N_23474,N_23878);
xor U24618 (N_24618,N_23491,N_23929);
and U24619 (N_24619,N_23688,N_23343);
nand U24620 (N_24620,N_23205,N_23160);
or U24621 (N_24621,N_23919,N_22889);
or U24622 (N_24622,N_23290,N_23114);
xnor U24623 (N_24623,N_23600,N_23860);
or U24624 (N_24624,N_23767,N_23356);
or U24625 (N_24625,N_23489,N_23219);
nand U24626 (N_24626,N_22951,N_22963);
xor U24627 (N_24627,N_22850,N_23798);
or U24628 (N_24628,N_22885,N_23509);
and U24629 (N_24629,N_23449,N_23304);
xor U24630 (N_24630,N_22829,N_23131);
or U24631 (N_24631,N_23270,N_23833);
or U24632 (N_24632,N_23538,N_23972);
and U24633 (N_24633,N_23064,N_23173);
xor U24634 (N_24634,N_23652,N_22938);
nor U24635 (N_24635,N_23874,N_23612);
and U24636 (N_24636,N_22935,N_23016);
nor U24637 (N_24637,N_22945,N_23746);
nand U24638 (N_24638,N_23450,N_23563);
xnor U24639 (N_24639,N_23473,N_22814);
nor U24640 (N_24640,N_23295,N_23297);
xor U24641 (N_24641,N_23124,N_23834);
nor U24642 (N_24642,N_23665,N_23229);
and U24643 (N_24643,N_22864,N_23905);
and U24644 (N_24644,N_23173,N_23661);
nand U24645 (N_24645,N_23067,N_23037);
xnor U24646 (N_24646,N_23541,N_23328);
xor U24647 (N_24647,N_23193,N_23220);
nor U24648 (N_24648,N_23200,N_22965);
and U24649 (N_24649,N_23712,N_22819);
or U24650 (N_24650,N_23911,N_23690);
nor U24651 (N_24651,N_23952,N_23132);
xnor U24652 (N_24652,N_23886,N_23392);
nand U24653 (N_24653,N_23197,N_23410);
and U24654 (N_24654,N_23218,N_23691);
or U24655 (N_24655,N_23081,N_23283);
nor U24656 (N_24656,N_23316,N_23242);
and U24657 (N_24657,N_23867,N_23443);
nor U24658 (N_24658,N_23088,N_23804);
xor U24659 (N_24659,N_22807,N_23721);
nor U24660 (N_24660,N_23763,N_23153);
nor U24661 (N_24661,N_23408,N_23282);
nand U24662 (N_24662,N_23079,N_23829);
and U24663 (N_24663,N_23531,N_22827);
or U24664 (N_24664,N_23098,N_23360);
xor U24665 (N_24665,N_23595,N_23068);
xnor U24666 (N_24666,N_23229,N_23661);
or U24667 (N_24667,N_22850,N_23717);
and U24668 (N_24668,N_23235,N_23323);
nor U24669 (N_24669,N_22879,N_23185);
and U24670 (N_24670,N_23547,N_23796);
xor U24671 (N_24671,N_22822,N_23593);
and U24672 (N_24672,N_23509,N_23672);
nand U24673 (N_24673,N_23981,N_23931);
or U24674 (N_24674,N_22939,N_23915);
and U24675 (N_24675,N_23105,N_22810);
nand U24676 (N_24676,N_23152,N_23313);
nor U24677 (N_24677,N_23184,N_23441);
or U24678 (N_24678,N_23710,N_23870);
nor U24679 (N_24679,N_23010,N_23279);
or U24680 (N_24680,N_23535,N_23714);
xor U24681 (N_24681,N_22851,N_22897);
nor U24682 (N_24682,N_23894,N_23177);
or U24683 (N_24683,N_23313,N_22882);
or U24684 (N_24684,N_22950,N_23432);
nor U24685 (N_24685,N_23733,N_22885);
nor U24686 (N_24686,N_23184,N_23643);
or U24687 (N_24687,N_23253,N_22963);
xnor U24688 (N_24688,N_22945,N_23939);
nand U24689 (N_24689,N_23813,N_23778);
xnor U24690 (N_24690,N_23830,N_23407);
nor U24691 (N_24691,N_23985,N_23767);
nor U24692 (N_24692,N_23480,N_23813);
nand U24693 (N_24693,N_23625,N_22922);
nor U24694 (N_24694,N_22921,N_23044);
and U24695 (N_24695,N_23389,N_23452);
xor U24696 (N_24696,N_23689,N_23860);
nand U24697 (N_24697,N_22832,N_23410);
xor U24698 (N_24698,N_23046,N_23091);
xnor U24699 (N_24699,N_22930,N_23420);
nand U24700 (N_24700,N_23730,N_23471);
or U24701 (N_24701,N_22800,N_23891);
xnor U24702 (N_24702,N_23688,N_23169);
or U24703 (N_24703,N_23059,N_23092);
xnor U24704 (N_24704,N_23379,N_23586);
or U24705 (N_24705,N_23931,N_23365);
and U24706 (N_24706,N_23219,N_23788);
and U24707 (N_24707,N_23610,N_23356);
or U24708 (N_24708,N_23813,N_23431);
or U24709 (N_24709,N_23337,N_23619);
or U24710 (N_24710,N_23982,N_23798);
nand U24711 (N_24711,N_23365,N_23217);
nand U24712 (N_24712,N_22999,N_23805);
xor U24713 (N_24713,N_22963,N_23131);
or U24714 (N_24714,N_23142,N_23116);
nor U24715 (N_24715,N_23285,N_23753);
and U24716 (N_24716,N_23403,N_23594);
nand U24717 (N_24717,N_22939,N_23355);
nor U24718 (N_24718,N_23475,N_22815);
nor U24719 (N_24719,N_23591,N_22903);
or U24720 (N_24720,N_23393,N_23154);
or U24721 (N_24721,N_23051,N_23077);
xnor U24722 (N_24722,N_23154,N_22804);
and U24723 (N_24723,N_23622,N_23641);
nor U24724 (N_24724,N_23058,N_23669);
nor U24725 (N_24725,N_23448,N_23275);
or U24726 (N_24726,N_23218,N_23263);
nor U24727 (N_24727,N_23002,N_22906);
nand U24728 (N_24728,N_23815,N_23291);
and U24729 (N_24729,N_22931,N_23074);
and U24730 (N_24730,N_23516,N_23346);
nor U24731 (N_24731,N_23011,N_23674);
and U24732 (N_24732,N_23661,N_23235);
or U24733 (N_24733,N_23801,N_22966);
and U24734 (N_24734,N_23165,N_22935);
and U24735 (N_24735,N_23494,N_23639);
xnor U24736 (N_24736,N_23518,N_23236);
xor U24737 (N_24737,N_22847,N_23974);
nor U24738 (N_24738,N_23529,N_23155);
xnor U24739 (N_24739,N_23105,N_23493);
nand U24740 (N_24740,N_23568,N_23738);
xor U24741 (N_24741,N_23421,N_23480);
and U24742 (N_24742,N_23354,N_23511);
or U24743 (N_24743,N_23100,N_23709);
nor U24744 (N_24744,N_22944,N_23207);
and U24745 (N_24745,N_22908,N_23096);
and U24746 (N_24746,N_23558,N_23209);
or U24747 (N_24747,N_23664,N_22992);
and U24748 (N_24748,N_23894,N_23301);
nand U24749 (N_24749,N_23717,N_23127);
or U24750 (N_24750,N_23772,N_23817);
or U24751 (N_24751,N_23684,N_23282);
nand U24752 (N_24752,N_23701,N_23423);
and U24753 (N_24753,N_23518,N_22933);
xor U24754 (N_24754,N_23274,N_23909);
nor U24755 (N_24755,N_23532,N_23900);
nand U24756 (N_24756,N_22920,N_22874);
xnor U24757 (N_24757,N_23931,N_23881);
xnor U24758 (N_24758,N_23821,N_23581);
xor U24759 (N_24759,N_22845,N_22908);
nand U24760 (N_24760,N_23809,N_23852);
xnor U24761 (N_24761,N_22910,N_23573);
xnor U24762 (N_24762,N_23793,N_23224);
or U24763 (N_24763,N_22814,N_23181);
or U24764 (N_24764,N_22961,N_23800);
nand U24765 (N_24765,N_23222,N_23176);
xor U24766 (N_24766,N_23504,N_23136);
nand U24767 (N_24767,N_23308,N_23517);
nor U24768 (N_24768,N_23380,N_23395);
nor U24769 (N_24769,N_23221,N_23384);
nand U24770 (N_24770,N_23428,N_23054);
nand U24771 (N_24771,N_23424,N_23014);
nand U24772 (N_24772,N_23714,N_23485);
nor U24773 (N_24773,N_23192,N_23361);
and U24774 (N_24774,N_22896,N_22905);
or U24775 (N_24775,N_22963,N_22803);
xor U24776 (N_24776,N_23431,N_22885);
nor U24777 (N_24777,N_23968,N_23854);
or U24778 (N_24778,N_23930,N_22861);
or U24779 (N_24779,N_23668,N_23990);
nand U24780 (N_24780,N_23101,N_23107);
or U24781 (N_24781,N_23488,N_23056);
nand U24782 (N_24782,N_23875,N_23789);
or U24783 (N_24783,N_23085,N_23421);
nor U24784 (N_24784,N_23756,N_23369);
nor U24785 (N_24785,N_23530,N_23598);
or U24786 (N_24786,N_23953,N_22853);
nor U24787 (N_24787,N_23778,N_23259);
nand U24788 (N_24788,N_23129,N_23945);
and U24789 (N_24789,N_22851,N_23394);
nor U24790 (N_24790,N_23632,N_23279);
xor U24791 (N_24791,N_23931,N_23926);
and U24792 (N_24792,N_23542,N_23125);
nand U24793 (N_24793,N_23391,N_22868);
nor U24794 (N_24794,N_22908,N_23669);
or U24795 (N_24795,N_23005,N_23587);
or U24796 (N_24796,N_23714,N_23024);
nor U24797 (N_24797,N_23237,N_22983);
nand U24798 (N_24798,N_23226,N_23198);
nand U24799 (N_24799,N_23131,N_23962);
nand U24800 (N_24800,N_23967,N_23201);
nor U24801 (N_24801,N_23056,N_23425);
or U24802 (N_24802,N_23341,N_23266);
and U24803 (N_24803,N_22897,N_23048);
nor U24804 (N_24804,N_22851,N_23038);
xor U24805 (N_24805,N_23235,N_23969);
nor U24806 (N_24806,N_23184,N_22897);
or U24807 (N_24807,N_23858,N_23755);
nand U24808 (N_24808,N_23240,N_23583);
nand U24809 (N_24809,N_22930,N_23480);
or U24810 (N_24810,N_23704,N_22888);
nor U24811 (N_24811,N_23019,N_23135);
and U24812 (N_24812,N_23039,N_23641);
or U24813 (N_24813,N_22939,N_23638);
and U24814 (N_24814,N_23974,N_23635);
nor U24815 (N_24815,N_23691,N_23853);
or U24816 (N_24816,N_23915,N_22923);
nor U24817 (N_24817,N_23768,N_23762);
nand U24818 (N_24818,N_23469,N_23405);
or U24819 (N_24819,N_23846,N_23739);
nand U24820 (N_24820,N_23540,N_23212);
nand U24821 (N_24821,N_23097,N_23273);
nand U24822 (N_24822,N_22942,N_23000);
or U24823 (N_24823,N_23257,N_22823);
and U24824 (N_24824,N_23693,N_23609);
nor U24825 (N_24825,N_23618,N_22980);
or U24826 (N_24826,N_23905,N_22857);
nor U24827 (N_24827,N_23341,N_23577);
or U24828 (N_24828,N_23445,N_22837);
xnor U24829 (N_24829,N_23888,N_23142);
xnor U24830 (N_24830,N_23635,N_23300);
xor U24831 (N_24831,N_23561,N_23396);
or U24832 (N_24832,N_23422,N_23016);
or U24833 (N_24833,N_23822,N_23891);
or U24834 (N_24834,N_22818,N_23213);
nand U24835 (N_24835,N_23553,N_23192);
xnor U24836 (N_24836,N_23066,N_23753);
nand U24837 (N_24837,N_23016,N_23454);
nor U24838 (N_24838,N_23662,N_23489);
or U24839 (N_24839,N_23784,N_23042);
nand U24840 (N_24840,N_23736,N_23616);
xor U24841 (N_24841,N_23980,N_22848);
nand U24842 (N_24842,N_23661,N_22918);
nand U24843 (N_24843,N_23614,N_23434);
or U24844 (N_24844,N_23575,N_22882);
xnor U24845 (N_24845,N_22941,N_23198);
xor U24846 (N_24846,N_23206,N_23619);
or U24847 (N_24847,N_23385,N_23741);
or U24848 (N_24848,N_23843,N_23100);
nor U24849 (N_24849,N_23702,N_23607);
xnor U24850 (N_24850,N_23090,N_23808);
or U24851 (N_24851,N_23998,N_23281);
and U24852 (N_24852,N_23756,N_23619);
nand U24853 (N_24853,N_23288,N_23831);
nor U24854 (N_24854,N_22871,N_23287);
nor U24855 (N_24855,N_23728,N_22949);
or U24856 (N_24856,N_22845,N_23020);
nor U24857 (N_24857,N_23609,N_23117);
or U24858 (N_24858,N_23688,N_23678);
or U24859 (N_24859,N_23896,N_22880);
or U24860 (N_24860,N_22845,N_23628);
nand U24861 (N_24861,N_23505,N_23589);
nand U24862 (N_24862,N_23557,N_23718);
nor U24863 (N_24863,N_23463,N_23803);
nand U24864 (N_24864,N_23964,N_23898);
xor U24865 (N_24865,N_23971,N_23822);
xor U24866 (N_24866,N_23322,N_23976);
xor U24867 (N_24867,N_23507,N_23898);
and U24868 (N_24868,N_23784,N_23823);
and U24869 (N_24869,N_23389,N_23299);
or U24870 (N_24870,N_23494,N_23921);
and U24871 (N_24871,N_22993,N_23232);
nand U24872 (N_24872,N_23078,N_23323);
nand U24873 (N_24873,N_23669,N_23358);
nand U24874 (N_24874,N_23857,N_22951);
or U24875 (N_24875,N_23701,N_23760);
nor U24876 (N_24876,N_23067,N_23586);
xor U24877 (N_24877,N_23714,N_23523);
nand U24878 (N_24878,N_23449,N_22969);
and U24879 (N_24879,N_23602,N_22870);
or U24880 (N_24880,N_23086,N_23052);
and U24881 (N_24881,N_22829,N_23403);
or U24882 (N_24882,N_23170,N_23533);
xnor U24883 (N_24883,N_22984,N_23676);
nor U24884 (N_24884,N_23485,N_23110);
nand U24885 (N_24885,N_23693,N_23975);
nor U24886 (N_24886,N_23655,N_23980);
or U24887 (N_24887,N_23239,N_23027);
and U24888 (N_24888,N_23918,N_22823);
nand U24889 (N_24889,N_23614,N_22891);
nand U24890 (N_24890,N_23375,N_23378);
nor U24891 (N_24891,N_23796,N_23248);
and U24892 (N_24892,N_22914,N_23211);
or U24893 (N_24893,N_23838,N_22880);
xnor U24894 (N_24894,N_22888,N_23858);
and U24895 (N_24895,N_23345,N_23065);
and U24896 (N_24896,N_23808,N_23263);
xor U24897 (N_24897,N_23624,N_22801);
nor U24898 (N_24898,N_23899,N_23869);
nand U24899 (N_24899,N_22962,N_23077);
and U24900 (N_24900,N_23756,N_23346);
and U24901 (N_24901,N_22802,N_23045);
xor U24902 (N_24902,N_23146,N_23896);
nand U24903 (N_24903,N_23244,N_23978);
nor U24904 (N_24904,N_23768,N_23838);
xnor U24905 (N_24905,N_22869,N_23283);
nor U24906 (N_24906,N_23368,N_23085);
and U24907 (N_24907,N_23642,N_23777);
and U24908 (N_24908,N_23082,N_23997);
nor U24909 (N_24909,N_23730,N_22893);
nor U24910 (N_24910,N_23573,N_23686);
nor U24911 (N_24911,N_23296,N_23954);
and U24912 (N_24912,N_23254,N_23600);
or U24913 (N_24913,N_23797,N_23205);
nand U24914 (N_24914,N_23871,N_23523);
nand U24915 (N_24915,N_23048,N_23136);
nand U24916 (N_24916,N_23238,N_22848);
xnor U24917 (N_24917,N_23350,N_23100);
xor U24918 (N_24918,N_23977,N_23163);
xor U24919 (N_24919,N_23232,N_22943);
or U24920 (N_24920,N_23024,N_23150);
and U24921 (N_24921,N_23211,N_23264);
nand U24922 (N_24922,N_23016,N_23411);
nor U24923 (N_24923,N_23970,N_23052);
nand U24924 (N_24924,N_23098,N_23537);
nor U24925 (N_24925,N_23944,N_23792);
nor U24926 (N_24926,N_23788,N_23440);
nand U24927 (N_24927,N_23922,N_22989);
nor U24928 (N_24928,N_23788,N_23561);
or U24929 (N_24929,N_23885,N_23509);
nand U24930 (N_24930,N_22926,N_23243);
nor U24931 (N_24931,N_23950,N_23372);
nand U24932 (N_24932,N_23098,N_23566);
or U24933 (N_24933,N_23698,N_23475);
or U24934 (N_24934,N_23142,N_22953);
nor U24935 (N_24935,N_23314,N_22842);
nand U24936 (N_24936,N_23840,N_23121);
and U24937 (N_24937,N_23767,N_22832);
nand U24938 (N_24938,N_23810,N_23942);
or U24939 (N_24939,N_23301,N_23244);
xor U24940 (N_24940,N_22915,N_23521);
nor U24941 (N_24941,N_23246,N_23886);
xor U24942 (N_24942,N_23336,N_23277);
xor U24943 (N_24943,N_23708,N_23298);
and U24944 (N_24944,N_23356,N_23587);
xnor U24945 (N_24945,N_22860,N_23416);
xnor U24946 (N_24946,N_23579,N_23622);
nand U24947 (N_24947,N_23213,N_23415);
nand U24948 (N_24948,N_23308,N_23518);
xnor U24949 (N_24949,N_23887,N_22912);
and U24950 (N_24950,N_22878,N_23626);
nor U24951 (N_24951,N_23291,N_23427);
or U24952 (N_24952,N_23103,N_23327);
and U24953 (N_24953,N_23167,N_23313);
nor U24954 (N_24954,N_22977,N_22940);
nor U24955 (N_24955,N_23049,N_23969);
or U24956 (N_24956,N_23890,N_23285);
nand U24957 (N_24957,N_23009,N_23879);
xor U24958 (N_24958,N_23580,N_23814);
nand U24959 (N_24959,N_22858,N_23728);
xnor U24960 (N_24960,N_23108,N_22866);
nor U24961 (N_24961,N_23515,N_23106);
nor U24962 (N_24962,N_23308,N_23600);
or U24963 (N_24963,N_23608,N_22958);
or U24964 (N_24964,N_23311,N_22960);
nand U24965 (N_24965,N_23791,N_23368);
or U24966 (N_24966,N_23634,N_23387);
nor U24967 (N_24967,N_23304,N_23006);
xnor U24968 (N_24968,N_23708,N_23052);
or U24969 (N_24969,N_23063,N_23708);
and U24970 (N_24970,N_22843,N_22834);
nand U24971 (N_24971,N_23906,N_22930);
nor U24972 (N_24972,N_23278,N_23176);
xnor U24973 (N_24973,N_23858,N_23074);
and U24974 (N_24974,N_23706,N_23390);
nand U24975 (N_24975,N_23896,N_23291);
nor U24976 (N_24976,N_23431,N_22895);
xnor U24977 (N_24977,N_23172,N_23997);
nand U24978 (N_24978,N_23496,N_23621);
nor U24979 (N_24979,N_23496,N_23986);
xor U24980 (N_24980,N_23793,N_23902);
nand U24981 (N_24981,N_23762,N_22947);
nand U24982 (N_24982,N_23212,N_23215);
nor U24983 (N_24983,N_23798,N_22835);
nand U24984 (N_24984,N_23101,N_23306);
or U24985 (N_24985,N_23537,N_23279);
nor U24986 (N_24986,N_23266,N_22909);
or U24987 (N_24987,N_23687,N_23355);
nand U24988 (N_24988,N_23375,N_23958);
nand U24989 (N_24989,N_23065,N_23988);
nor U24990 (N_24990,N_23833,N_23171);
and U24991 (N_24991,N_23029,N_23710);
xor U24992 (N_24992,N_23897,N_22944);
or U24993 (N_24993,N_23403,N_23110);
nor U24994 (N_24994,N_23748,N_23494);
nand U24995 (N_24995,N_23107,N_23699);
nand U24996 (N_24996,N_23441,N_23466);
and U24997 (N_24997,N_23285,N_23497);
or U24998 (N_24998,N_23727,N_22834);
and U24999 (N_24999,N_23724,N_23966);
and U25000 (N_25000,N_23149,N_23022);
nand U25001 (N_25001,N_23767,N_22918);
and U25002 (N_25002,N_23819,N_23527);
and U25003 (N_25003,N_23180,N_23237);
xor U25004 (N_25004,N_23743,N_23551);
nand U25005 (N_25005,N_23001,N_23056);
nor U25006 (N_25006,N_23758,N_23844);
xnor U25007 (N_25007,N_23980,N_22985);
nor U25008 (N_25008,N_23603,N_23383);
nand U25009 (N_25009,N_23699,N_23960);
nor U25010 (N_25010,N_23488,N_23752);
and U25011 (N_25011,N_23755,N_23444);
and U25012 (N_25012,N_23408,N_23864);
nor U25013 (N_25013,N_23449,N_23834);
nor U25014 (N_25014,N_23614,N_23003);
and U25015 (N_25015,N_23638,N_23232);
or U25016 (N_25016,N_23789,N_23227);
and U25017 (N_25017,N_23286,N_23260);
xnor U25018 (N_25018,N_23907,N_23674);
nor U25019 (N_25019,N_23260,N_23898);
nand U25020 (N_25020,N_23664,N_23715);
and U25021 (N_25021,N_23155,N_23402);
nand U25022 (N_25022,N_23663,N_23864);
xor U25023 (N_25023,N_23853,N_23782);
or U25024 (N_25024,N_23139,N_22888);
nand U25025 (N_25025,N_23318,N_23092);
and U25026 (N_25026,N_23653,N_23770);
and U25027 (N_25027,N_23425,N_22817);
nor U25028 (N_25028,N_23033,N_23816);
nor U25029 (N_25029,N_23527,N_23890);
nand U25030 (N_25030,N_23049,N_23439);
xnor U25031 (N_25031,N_23575,N_22890);
nor U25032 (N_25032,N_23772,N_23082);
nor U25033 (N_25033,N_23237,N_23113);
or U25034 (N_25034,N_23545,N_23812);
and U25035 (N_25035,N_23403,N_23341);
xor U25036 (N_25036,N_23498,N_23258);
xnor U25037 (N_25037,N_23404,N_23079);
nand U25038 (N_25038,N_23456,N_23502);
nand U25039 (N_25039,N_22820,N_23347);
xnor U25040 (N_25040,N_22979,N_23178);
nor U25041 (N_25041,N_23814,N_22856);
or U25042 (N_25042,N_23330,N_22888);
nor U25043 (N_25043,N_22835,N_23056);
xnor U25044 (N_25044,N_23565,N_23281);
nand U25045 (N_25045,N_23499,N_23946);
and U25046 (N_25046,N_23374,N_23462);
or U25047 (N_25047,N_23561,N_23417);
and U25048 (N_25048,N_23007,N_23752);
or U25049 (N_25049,N_23559,N_23474);
and U25050 (N_25050,N_23857,N_23488);
and U25051 (N_25051,N_23203,N_22814);
xor U25052 (N_25052,N_23056,N_23253);
and U25053 (N_25053,N_23345,N_22874);
and U25054 (N_25054,N_23629,N_23218);
nand U25055 (N_25055,N_23199,N_22978);
nand U25056 (N_25056,N_23807,N_23621);
xor U25057 (N_25057,N_23798,N_23130);
nand U25058 (N_25058,N_23113,N_23815);
or U25059 (N_25059,N_23587,N_23481);
nand U25060 (N_25060,N_23895,N_23685);
or U25061 (N_25061,N_23643,N_22937);
nor U25062 (N_25062,N_22813,N_23233);
nand U25063 (N_25063,N_23971,N_23714);
nor U25064 (N_25064,N_22988,N_23965);
xnor U25065 (N_25065,N_23218,N_23782);
xor U25066 (N_25066,N_23652,N_23297);
nand U25067 (N_25067,N_23591,N_23621);
or U25068 (N_25068,N_23830,N_22970);
and U25069 (N_25069,N_23440,N_22956);
nand U25070 (N_25070,N_22802,N_23517);
nor U25071 (N_25071,N_23876,N_23433);
nor U25072 (N_25072,N_23177,N_22844);
nor U25073 (N_25073,N_23216,N_23273);
and U25074 (N_25074,N_22966,N_23684);
and U25075 (N_25075,N_23718,N_23808);
nor U25076 (N_25076,N_22966,N_23946);
nand U25077 (N_25077,N_23194,N_23140);
and U25078 (N_25078,N_23095,N_23361);
nand U25079 (N_25079,N_23842,N_23640);
or U25080 (N_25080,N_23040,N_23597);
xor U25081 (N_25081,N_23740,N_23755);
or U25082 (N_25082,N_23494,N_23858);
and U25083 (N_25083,N_23321,N_23157);
and U25084 (N_25084,N_23976,N_23046);
and U25085 (N_25085,N_23562,N_23082);
or U25086 (N_25086,N_23583,N_23276);
nor U25087 (N_25087,N_23127,N_23883);
nand U25088 (N_25088,N_22832,N_23455);
nand U25089 (N_25089,N_23024,N_23132);
xor U25090 (N_25090,N_23153,N_23432);
nor U25091 (N_25091,N_23486,N_22982);
or U25092 (N_25092,N_23404,N_23147);
and U25093 (N_25093,N_23643,N_23543);
and U25094 (N_25094,N_22939,N_23651);
nand U25095 (N_25095,N_23795,N_23529);
xor U25096 (N_25096,N_23318,N_23548);
xnor U25097 (N_25097,N_22883,N_23894);
and U25098 (N_25098,N_23167,N_23341);
nand U25099 (N_25099,N_23637,N_23351);
nor U25100 (N_25100,N_23589,N_23259);
nor U25101 (N_25101,N_23893,N_23384);
or U25102 (N_25102,N_23193,N_23680);
or U25103 (N_25103,N_23120,N_23132);
and U25104 (N_25104,N_23905,N_23223);
xnor U25105 (N_25105,N_23354,N_23098);
nand U25106 (N_25106,N_23064,N_22887);
nor U25107 (N_25107,N_23501,N_23637);
nor U25108 (N_25108,N_23964,N_23078);
nor U25109 (N_25109,N_23215,N_23654);
xnor U25110 (N_25110,N_23566,N_23071);
nor U25111 (N_25111,N_23923,N_23790);
and U25112 (N_25112,N_23686,N_22969);
and U25113 (N_25113,N_23499,N_22893);
nand U25114 (N_25114,N_23719,N_23261);
nor U25115 (N_25115,N_22984,N_23368);
or U25116 (N_25116,N_23176,N_23820);
xor U25117 (N_25117,N_22989,N_23105);
and U25118 (N_25118,N_22989,N_23308);
nand U25119 (N_25119,N_22979,N_22953);
nor U25120 (N_25120,N_23932,N_23322);
nor U25121 (N_25121,N_22923,N_23935);
and U25122 (N_25122,N_23649,N_23797);
and U25123 (N_25123,N_22836,N_23228);
nor U25124 (N_25124,N_22985,N_23866);
nand U25125 (N_25125,N_23544,N_23649);
xor U25126 (N_25126,N_23776,N_23404);
or U25127 (N_25127,N_23450,N_23781);
and U25128 (N_25128,N_23304,N_23723);
nor U25129 (N_25129,N_23253,N_23099);
xnor U25130 (N_25130,N_23799,N_23280);
nand U25131 (N_25131,N_22805,N_23759);
nand U25132 (N_25132,N_23969,N_23050);
and U25133 (N_25133,N_23963,N_23941);
xor U25134 (N_25134,N_23832,N_23897);
xnor U25135 (N_25135,N_23629,N_23712);
xor U25136 (N_25136,N_23717,N_23438);
nor U25137 (N_25137,N_22971,N_23663);
and U25138 (N_25138,N_23938,N_23687);
and U25139 (N_25139,N_22954,N_23592);
or U25140 (N_25140,N_23538,N_23950);
and U25141 (N_25141,N_23090,N_23993);
or U25142 (N_25142,N_23230,N_22905);
xnor U25143 (N_25143,N_22835,N_23557);
or U25144 (N_25144,N_23301,N_23398);
nand U25145 (N_25145,N_23627,N_23441);
nor U25146 (N_25146,N_23972,N_23581);
xor U25147 (N_25147,N_22926,N_23345);
nor U25148 (N_25148,N_22847,N_23391);
xor U25149 (N_25149,N_23408,N_23670);
and U25150 (N_25150,N_23042,N_23401);
and U25151 (N_25151,N_23487,N_22813);
or U25152 (N_25152,N_23647,N_23917);
nand U25153 (N_25153,N_23012,N_22956);
nand U25154 (N_25154,N_23388,N_23726);
xnor U25155 (N_25155,N_23285,N_23450);
and U25156 (N_25156,N_23411,N_23819);
xor U25157 (N_25157,N_23183,N_23358);
nor U25158 (N_25158,N_23149,N_23117);
nor U25159 (N_25159,N_23872,N_22982);
or U25160 (N_25160,N_23460,N_23386);
nor U25161 (N_25161,N_23897,N_23725);
xor U25162 (N_25162,N_23596,N_23793);
nand U25163 (N_25163,N_23349,N_23337);
xor U25164 (N_25164,N_23110,N_23829);
xor U25165 (N_25165,N_23978,N_23156);
xnor U25166 (N_25166,N_23402,N_23902);
or U25167 (N_25167,N_22901,N_22917);
nor U25168 (N_25168,N_22886,N_23856);
or U25169 (N_25169,N_23842,N_23651);
nor U25170 (N_25170,N_23616,N_23965);
and U25171 (N_25171,N_23902,N_23647);
nand U25172 (N_25172,N_23958,N_23384);
xnor U25173 (N_25173,N_22822,N_23664);
and U25174 (N_25174,N_23525,N_23896);
xnor U25175 (N_25175,N_22922,N_23467);
and U25176 (N_25176,N_22866,N_23256);
nor U25177 (N_25177,N_23329,N_23220);
nand U25178 (N_25178,N_23071,N_23249);
nand U25179 (N_25179,N_23808,N_23201);
and U25180 (N_25180,N_23270,N_23781);
nand U25181 (N_25181,N_23053,N_23814);
and U25182 (N_25182,N_23720,N_22836);
xnor U25183 (N_25183,N_23523,N_23152);
nor U25184 (N_25184,N_22927,N_23804);
or U25185 (N_25185,N_23902,N_22911);
xnor U25186 (N_25186,N_23400,N_23190);
xor U25187 (N_25187,N_23241,N_23957);
xor U25188 (N_25188,N_22974,N_23586);
and U25189 (N_25189,N_23172,N_23384);
xnor U25190 (N_25190,N_23424,N_23604);
nor U25191 (N_25191,N_23853,N_23001);
nor U25192 (N_25192,N_23003,N_23714);
or U25193 (N_25193,N_23584,N_23984);
nand U25194 (N_25194,N_23407,N_23161);
xor U25195 (N_25195,N_23132,N_23931);
or U25196 (N_25196,N_23820,N_22967);
xor U25197 (N_25197,N_23020,N_23137);
and U25198 (N_25198,N_23515,N_23386);
or U25199 (N_25199,N_23318,N_23827);
and U25200 (N_25200,N_24093,N_24861);
and U25201 (N_25201,N_24050,N_24577);
and U25202 (N_25202,N_24470,N_24844);
or U25203 (N_25203,N_24984,N_24647);
or U25204 (N_25204,N_24010,N_24567);
and U25205 (N_25205,N_24664,N_25108);
and U25206 (N_25206,N_24157,N_25188);
nor U25207 (N_25207,N_24649,N_24877);
xor U25208 (N_25208,N_24570,N_24156);
nand U25209 (N_25209,N_24055,N_24442);
xnor U25210 (N_25210,N_24252,N_24441);
xnor U25211 (N_25211,N_24428,N_25152);
nor U25212 (N_25212,N_24163,N_24932);
xor U25213 (N_25213,N_24939,N_24888);
and U25214 (N_25214,N_24316,N_24020);
xnor U25215 (N_25215,N_25055,N_24119);
nor U25216 (N_25216,N_24762,N_25088);
and U25217 (N_25217,N_24137,N_24746);
nor U25218 (N_25218,N_24096,N_25021);
nand U25219 (N_25219,N_24601,N_25130);
or U25220 (N_25220,N_24091,N_24735);
xor U25221 (N_25221,N_24634,N_24065);
nor U25222 (N_25222,N_24941,N_24794);
nor U25223 (N_25223,N_24040,N_24685);
nand U25224 (N_25224,N_24711,N_24381);
or U25225 (N_25225,N_25120,N_24704);
xnor U25226 (N_25226,N_24788,N_24307);
xor U25227 (N_25227,N_24856,N_24404);
and U25228 (N_25228,N_24004,N_24727);
nor U25229 (N_25229,N_24658,N_24573);
or U25230 (N_25230,N_24579,N_24412);
xor U25231 (N_25231,N_25114,N_25176);
nand U25232 (N_25232,N_24668,N_24853);
nor U25233 (N_25233,N_24125,N_24189);
nor U25234 (N_25234,N_24029,N_24009);
and U25235 (N_25235,N_24437,N_25047);
or U25236 (N_25236,N_24945,N_24636);
and U25237 (N_25237,N_24838,N_24966);
nand U25238 (N_25238,N_24011,N_24980);
nor U25239 (N_25239,N_24348,N_24660);
nand U25240 (N_25240,N_24247,N_24534);
xor U25241 (N_25241,N_24253,N_24198);
and U25242 (N_25242,N_24070,N_24708);
xor U25243 (N_25243,N_25184,N_24349);
or U25244 (N_25244,N_24483,N_24041);
xnor U25245 (N_25245,N_24633,N_24213);
nor U25246 (N_25246,N_24960,N_24002);
nor U25247 (N_25247,N_24904,N_24695);
and U25248 (N_25248,N_25058,N_24515);
and U25249 (N_25249,N_25041,N_24149);
or U25250 (N_25250,N_24518,N_25175);
nand U25251 (N_25251,N_24243,N_24582);
or U25252 (N_25252,N_25039,N_25071);
and U25253 (N_25253,N_24763,N_24774);
nand U25254 (N_25254,N_24802,N_24384);
or U25255 (N_25255,N_24211,N_24488);
nand U25256 (N_25256,N_25013,N_24118);
or U25257 (N_25257,N_24288,N_24102);
xor U25258 (N_25258,N_24106,N_24602);
nor U25259 (N_25259,N_25089,N_24342);
xor U25260 (N_25260,N_24075,N_24265);
and U25261 (N_25261,N_24885,N_24849);
xnor U25262 (N_25262,N_25032,N_24204);
and U25263 (N_25263,N_24353,N_25099);
xnor U25264 (N_25264,N_25098,N_24425);
xnor U25265 (N_25265,N_24789,N_24955);
and U25266 (N_25266,N_24071,N_25082);
and U25267 (N_25267,N_24741,N_24187);
or U25268 (N_25268,N_25036,N_24300);
xnor U25269 (N_25269,N_24299,N_24394);
and U25270 (N_25270,N_24832,N_24988);
nor U25271 (N_25271,N_24476,N_24031);
or U25272 (N_25272,N_25040,N_24268);
nor U25273 (N_25273,N_24641,N_24646);
nand U25274 (N_25274,N_24403,N_24094);
and U25275 (N_25275,N_24599,N_25094);
nor U25276 (N_25276,N_24245,N_24327);
xor U25277 (N_25277,N_24703,N_25111);
xnor U25278 (N_25278,N_24712,N_24807);
and U25279 (N_25279,N_25006,N_24795);
nor U25280 (N_25280,N_24555,N_24090);
nand U25281 (N_25281,N_24781,N_24206);
nor U25282 (N_25282,N_24554,N_24336);
and U25283 (N_25283,N_24016,N_24655);
nand U25284 (N_25284,N_24144,N_24449);
and U25285 (N_25285,N_24236,N_25012);
xnor U25286 (N_25286,N_24957,N_25074);
nand U25287 (N_25287,N_25155,N_24550);
or U25288 (N_25288,N_24473,N_25007);
xor U25289 (N_25289,N_24419,N_24337);
and U25290 (N_25290,N_24858,N_24026);
nand U25291 (N_25291,N_25044,N_25078);
xor U25292 (N_25292,N_24768,N_24507);
nor U25293 (N_25293,N_25056,N_24148);
nand U25294 (N_25294,N_24521,N_24220);
nor U25295 (N_25295,N_24495,N_24811);
and U25296 (N_25296,N_24973,N_24304);
or U25297 (N_25297,N_24350,N_24538);
xnor U25298 (N_25298,N_24716,N_25001);
xnor U25299 (N_25299,N_24669,N_25080);
nor U25300 (N_25300,N_24110,N_24295);
and U25301 (N_25301,N_24701,N_25073);
nand U25302 (N_25302,N_24458,N_24522);
nand U25303 (N_25303,N_24101,N_24235);
nor U25304 (N_25304,N_24535,N_24017);
or U25305 (N_25305,N_24146,N_24320);
or U25306 (N_25306,N_25186,N_25196);
or U25307 (N_25307,N_24635,N_24631);
or U25308 (N_25308,N_24971,N_24462);
nand U25309 (N_25309,N_24183,N_25023);
and U25310 (N_25310,N_25124,N_24175);
nor U25311 (N_25311,N_24386,N_24439);
and U25312 (N_25312,N_24938,N_24045);
and U25313 (N_25313,N_24876,N_24451);
nand U25314 (N_25314,N_24315,N_24200);
nor U25315 (N_25315,N_24296,N_24594);
or U25316 (N_25316,N_24022,N_24563);
nor U25317 (N_25317,N_24623,N_24410);
and U25318 (N_25318,N_24291,N_25125);
nand U25319 (N_25319,N_24747,N_24651);
and U25320 (N_25320,N_24810,N_24078);
or U25321 (N_25321,N_24355,N_24466);
or U25322 (N_25322,N_24924,N_24943);
and U25323 (N_25323,N_24151,N_24277);
and U25324 (N_25324,N_25109,N_24196);
or U25325 (N_25325,N_24835,N_24834);
and U25326 (N_25326,N_24696,N_24529);
nor U25327 (N_25327,N_25000,N_25171);
xor U25328 (N_25328,N_24620,N_24383);
nor U25329 (N_25329,N_24608,N_24082);
xnor U25330 (N_25330,N_24049,N_24132);
nand U25331 (N_25331,N_24598,N_24457);
nor U25332 (N_25332,N_24025,N_24749);
or U25333 (N_25333,N_24677,N_24580);
nor U25334 (N_25334,N_24186,N_24697);
xor U25335 (N_25335,N_24516,N_24848);
nand U25336 (N_25336,N_24285,N_24143);
nand U25337 (N_25337,N_24940,N_24318);
xor U25338 (N_25338,N_25095,N_24072);
and U25339 (N_25339,N_24409,N_24073);
nand U25340 (N_25340,N_24926,N_25031);
or U25341 (N_25341,N_24339,N_24038);
or U25342 (N_25342,N_24389,N_24818);
and U25343 (N_25343,N_25028,N_24417);
or U25344 (N_25344,N_24165,N_24205);
nor U25345 (N_25345,N_24622,N_25057);
or U25346 (N_25346,N_24364,N_24923);
nor U25347 (N_25347,N_25160,N_24278);
nor U25348 (N_25348,N_24574,N_24797);
nand U25349 (N_25349,N_24482,N_25113);
and U25350 (N_25350,N_24153,N_24314);
nand U25351 (N_25351,N_24237,N_24341);
nand U25352 (N_25352,N_24572,N_24970);
and U25353 (N_25353,N_24232,N_24880);
or U25354 (N_25354,N_24357,N_24775);
xnor U25355 (N_25355,N_25133,N_24748);
or U25356 (N_25356,N_24657,N_24780);
xor U25357 (N_25357,N_25167,N_24257);
or U25358 (N_25358,N_24497,N_24120);
nand U25359 (N_25359,N_25198,N_24290);
or U25360 (N_25360,N_24855,N_24498);
or U25361 (N_25361,N_24991,N_24737);
and U25362 (N_25362,N_24714,N_24413);
xnor U25363 (N_25363,N_24281,N_24546);
and U25364 (N_25364,N_24124,N_25003);
nand U25365 (N_25365,N_24385,N_24105);
nand U25366 (N_25366,N_24760,N_24445);
xnor U25367 (N_25367,N_24282,N_24432);
or U25368 (N_25368,N_24951,N_24393);
nor U25369 (N_25369,N_24373,N_24301);
xnor U25370 (N_25370,N_25153,N_24905);
xnor U25371 (N_25371,N_24773,N_24562);
nand U25372 (N_25372,N_24347,N_24167);
or U25373 (N_25373,N_24533,N_24638);
xnor U25374 (N_25374,N_24551,N_24370);
nand U25375 (N_25375,N_24830,N_24944);
nor U25376 (N_25376,N_25024,N_24074);
or U25377 (N_25377,N_24424,N_24345);
or U25378 (N_25378,N_24934,N_24799);
nor U25379 (N_25379,N_24680,N_24193);
xor U25380 (N_25380,N_24272,N_24911);
and U25381 (N_25381,N_24374,N_24308);
and U25382 (N_25382,N_24251,N_24850);
xor U25383 (N_25383,N_25178,N_25187);
or U25384 (N_25384,N_25164,N_25062);
or U25385 (N_25385,N_24821,N_24012);
xor U25386 (N_25386,N_24879,N_24242);
nand U25387 (N_25387,N_25191,N_25180);
or U25388 (N_25388,N_24293,N_24104);
nor U25389 (N_25389,N_24994,N_24450);
nand U25390 (N_25390,N_24600,N_24197);
xnor U25391 (N_25391,N_24999,N_24116);
or U25392 (N_25392,N_24590,N_24454);
nor U25393 (N_25393,N_24258,N_24099);
or U25394 (N_25394,N_24979,N_24881);
nand U25395 (N_25395,N_24732,N_24214);
or U25396 (N_25396,N_24210,N_24612);
nand U25397 (N_25397,N_24079,N_24378);
or U25398 (N_25398,N_24887,N_24405);
xor U25399 (N_25399,N_24867,N_24048);
nor U25400 (N_25400,N_24279,N_24665);
and U25401 (N_25401,N_24241,N_24765);
or U25402 (N_25402,N_24037,N_24962);
nor U25403 (N_25403,N_24840,N_24808);
nand U25404 (N_25404,N_24618,N_24134);
or U25405 (N_25405,N_25190,N_24207);
nand U25406 (N_25406,N_24063,N_24418);
or U25407 (N_25407,N_24560,N_25179);
xnor U25408 (N_25408,N_24069,N_25137);
nor U25409 (N_25409,N_24202,N_24001);
xnor U25410 (N_25410,N_24035,N_24319);
nor U25411 (N_25411,N_25157,N_24606);
or U25412 (N_25412,N_24178,N_24740);
and U25413 (N_25413,N_24162,N_24261);
nor U25414 (N_25414,N_24224,N_24369);
nor U25415 (N_25415,N_24733,N_24414);
nor U25416 (N_25416,N_24985,N_25106);
or U25417 (N_25417,N_24216,N_24731);
nand U25418 (N_25418,N_24603,N_25090);
or U25419 (N_25419,N_24547,N_24054);
xnor U25420 (N_25420,N_24201,N_24524);
and U25421 (N_25421,N_24890,N_24906);
or U25422 (N_25422,N_24557,N_24707);
and U25423 (N_25423,N_24356,N_24313);
and U25424 (N_25424,N_24455,N_24123);
xnor U25425 (N_25425,N_24682,N_25129);
or U25426 (N_25426,N_24109,N_24897);
xor U25427 (N_25427,N_24303,N_24138);
xnor U25428 (N_25428,N_24064,N_24929);
nor U25429 (N_25429,N_24791,N_24586);
nand U25430 (N_25430,N_25034,N_24761);
xnor U25431 (N_25431,N_24292,N_24159);
and U25432 (N_25432,N_24294,N_24523);
nor U25433 (N_25433,N_24346,N_24916);
or U25434 (N_25434,N_24368,N_24478);
and U25435 (N_25435,N_24751,N_25181);
xnor U25436 (N_25436,N_24479,N_24539);
and U25437 (N_25437,N_24467,N_24103);
nor U25438 (N_25438,N_24352,N_24757);
xnor U25439 (N_25439,N_24689,N_25189);
nor U25440 (N_25440,N_24726,N_24782);
or U25441 (N_25441,N_24267,N_24325);
or U25442 (N_25442,N_24833,N_24796);
or U25443 (N_25443,N_24305,N_24397);
or U25444 (N_25444,N_24542,N_24800);
or U25445 (N_25445,N_24433,N_24812);
nand U25446 (N_25446,N_24902,N_24392);
nor U25447 (N_25447,N_24095,N_25117);
nor U25448 (N_25448,N_24687,N_25151);
nand U25449 (N_25449,N_24710,N_25022);
or U25450 (N_25450,N_25037,N_24042);
or U25451 (N_25451,N_24464,N_24842);
or U25452 (N_25452,N_24720,N_25146);
nand U25453 (N_25453,N_24785,N_25011);
and U25454 (N_25454,N_24475,N_24884);
nand U25455 (N_25455,N_25059,N_24387);
nor U25456 (N_25456,N_25101,N_24047);
xor U25457 (N_25457,N_24229,N_24508);
and U25458 (N_25458,N_24899,N_24595);
or U25459 (N_25459,N_24003,N_24452);
nand U25460 (N_25460,N_24209,N_25045);
nand U25461 (N_25461,N_24000,N_24164);
or U25462 (N_25462,N_24158,N_24772);
or U25463 (N_25463,N_24868,N_25173);
xnor U25464 (N_25464,N_24058,N_24171);
nor U25465 (N_25465,N_24321,N_24597);
or U25466 (N_25466,N_24836,N_24656);
nor U25467 (N_25467,N_25131,N_24400);
nand U25468 (N_25468,N_24130,N_24051);
or U25469 (N_25469,N_24783,N_24401);
and U25470 (N_25470,N_24262,N_25030);
and U25471 (N_25471,N_24920,N_24552);
and U25472 (N_25472,N_24827,N_25107);
xor U25473 (N_25473,N_24630,N_24584);
nand U25474 (N_25474,N_24334,N_24415);
nor U25475 (N_25475,N_24972,N_24933);
nor U25476 (N_25476,N_24825,N_25063);
nor U25477 (N_25477,N_24676,N_24605);
xor U25478 (N_25478,N_25132,N_24406);
nor U25479 (N_25479,N_25068,N_24375);
nor U25480 (N_25480,N_25118,N_24922);
or U25481 (N_25481,N_24632,N_24208);
or U25482 (N_25482,N_24983,N_25069);
nand U25483 (N_25483,N_24203,N_24097);
or U25484 (N_25484,N_24264,N_24581);
or U25485 (N_25485,N_24489,N_24244);
or U25486 (N_25486,N_24390,N_24246);
and U25487 (N_25487,N_24826,N_24005);
nor U25488 (N_25488,N_24684,N_24107);
xor U25489 (N_25489,N_24564,N_24512);
nand U25490 (N_25490,N_25075,N_24553);
or U25491 (N_25491,N_24233,N_24841);
nand U25492 (N_25492,N_24989,N_25064);
xor U25493 (N_25493,N_24587,N_24952);
nand U25494 (N_25494,N_25136,N_24862);
xnor U25495 (N_25495,N_24184,N_24487);
nor U25496 (N_25496,N_25084,N_24959);
nand U25497 (N_25497,N_25104,N_24459);
nor U25498 (N_25498,N_24366,N_24526);
nand U25499 (N_25499,N_24700,N_24066);
xor U25500 (N_25500,N_24947,N_24930);
and U25501 (N_25501,N_24444,N_24869);
nor U25502 (N_25502,N_24886,N_24613);
xnor U25503 (N_25503,N_24472,N_25017);
or U25504 (N_25504,N_24578,N_24817);
nand U25505 (N_25505,N_25083,N_24191);
nand U25506 (N_25506,N_24873,N_24532);
and U25507 (N_25507,N_24662,N_24477);
and U25508 (N_25508,N_24344,N_24212);
and U25509 (N_25509,N_24592,N_24126);
nor U25510 (N_25510,N_24297,N_24667);
nor U25511 (N_25511,N_24510,N_24083);
nor U25512 (N_25512,N_24129,N_24845);
nor U25513 (N_25513,N_24117,N_24798);
or U25514 (N_25514,N_24898,N_24484);
xor U25515 (N_25515,N_24982,N_25154);
nand U25516 (N_25516,N_24639,N_24872);
nor U25517 (N_25517,N_24958,N_24621);
or U25518 (N_25518,N_24976,N_25072);
or U25519 (N_25519,N_24494,N_25066);
xnor U25520 (N_25520,N_25170,N_24195);
xnor U25521 (N_25521,N_24504,N_25004);
and U25522 (N_25522,N_25018,N_24006);
nand U25523 (N_25523,N_24576,N_24756);
or U25524 (N_25524,N_24217,N_24030);
nor U25525 (N_25525,N_24739,N_24806);
nand U25526 (N_25526,N_25014,N_24372);
nand U25527 (N_25527,N_24227,N_24367);
xor U25528 (N_25528,N_25195,N_24527);
and U25529 (N_25529,N_24683,N_24371);
nor U25530 (N_25530,N_24505,N_25135);
and U25531 (N_25531,N_24447,N_24702);
or U25532 (N_25532,N_24270,N_24098);
and U25533 (N_25533,N_25065,N_25070);
nand U25534 (N_25534,N_24430,N_25161);
nand U25535 (N_25535,N_24274,N_24287);
nand U25536 (N_25536,N_24531,N_24892);
xnor U25537 (N_25537,N_24626,N_24147);
and U25538 (N_25538,N_24928,N_24427);
and U25539 (N_25539,N_24420,N_24990);
xor U25540 (N_25540,N_24617,N_24263);
nand U25541 (N_25541,N_24921,N_24583);
nor U25542 (N_25542,N_24998,N_25100);
nor U25543 (N_25543,N_24034,N_24610);
xor U25544 (N_25544,N_24736,N_24615);
or U25545 (N_25545,N_24276,N_24435);
and U25546 (N_25546,N_24250,N_24771);
nor U25547 (N_25547,N_24672,N_24331);
nor U25548 (N_25548,N_24218,N_24568);
and U25549 (N_25549,N_24721,N_24745);
xnor U25550 (N_25550,N_24330,N_25122);
or U25551 (N_25551,N_24152,N_24561);
nor U25552 (N_25552,N_24269,N_24831);
xnor U25553 (N_25553,N_24306,N_25144);
xor U25554 (N_25554,N_24062,N_25015);
or U25555 (N_25555,N_24688,N_24589);
nand U25556 (N_25556,N_24540,N_24174);
or U25557 (N_25557,N_24650,N_25081);
nand U25558 (N_25558,N_24543,N_24335);
nand U25559 (N_25559,N_24486,N_24659);
and U25560 (N_25560,N_25019,N_24429);
or U25561 (N_25561,N_24057,N_25020);
and U25562 (N_25562,N_24717,N_24490);
and U25563 (N_25563,N_24226,N_24919);
nand U25564 (N_25564,N_25005,N_24170);
nor U25565 (N_25565,N_25172,N_24365);
xor U25566 (N_25566,N_24565,N_24338);
xor U25567 (N_25567,N_24675,N_24804);
nor U25568 (N_25568,N_24160,N_25029);
or U25569 (N_25569,N_24502,N_24734);
xnor U25570 (N_25570,N_24333,N_24814);
and U25571 (N_25571,N_25141,N_24456);
xnor U25572 (N_25572,N_24240,N_24076);
and U25573 (N_25573,N_25116,N_24190);
xor U25574 (N_25574,N_24380,N_24377);
nor U25575 (N_25575,N_24993,N_24640);
or U25576 (N_25576,N_25199,N_24360);
and U25577 (N_25577,N_25166,N_24931);
and U25578 (N_25578,N_24624,N_24828);
nor U25579 (N_25579,N_24286,N_24870);
and U25580 (N_25580,N_24769,N_24100);
nor U25581 (N_25581,N_24113,N_24021);
xnor U25582 (N_25582,N_24758,N_24018);
or U25583 (N_25583,N_24019,N_24222);
or U25584 (N_25584,N_24837,N_25182);
nor U25585 (N_25585,N_24081,N_25105);
nor U25586 (N_25586,N_24997,N_24750);
and U25587 (N_25587,N_24426,N_24629);
and U25588 (N_25588,N_24228,N_24396);
and U25589 (N_25589,N_24503,N_24815);
and U25590 (N_25590,N_24092,N_24864);
or U25591 (N_25591,N_24436,N_24086);
xnor U25592 (N_25592,N_24168,N_24225);
nor U25593 (N_25593,N_24046,N_24754);
xnor U25594 (N_25594,N_24637,N_24465);
and U25595 (N_25595,N_24248,N_24914);
nand U25596 (N_25596,N_24219,N_25016);
nand U25597 (N_25597,N_24391,N_24537);
or U25598 (N_25598,N_24752,N_24181);
nand U25599 (N_25599,N_24779,N_24363);
or U25600 (N_25600,N_24678,N_25147);
nor U25601 (N_25601,N_24154,N_25127);
xnor U25602 (N_25602,N_24014,N_24878);
nand U25603 (N_25603,N_25138,N_24525);
and U25604 (N_25604,N_24585,N_24961);
nand U25605 (N_25605,N_24852,N_24974);
and U25606 (N_25606,N_24423,N_24388);
or U25607 (N_25607,N_24801,N_24645);
nand U25608 (N_25608,N_24199,N_24298);
nand U25609 (N_25609,N_24694,N_24491);
nor U25610 (N_25610,N_24142,N_25126);
or U25611 (N_25611,N_24709,N_24896);
nor U25612 (N_25612,N_24544,N_24813);
xnor U25613 (N_25613,N_25183,N_24273);
nand U25614 (N_25614,N_24770,N_24173);
nand U25615 (N_25615,N_24965,N_24936);
xnor U25616 (N_25616,N_25010,N_24468);
and U25617 (N_25617,N_24949,N_24463);
xor U25618 (N_25618,N_25162,N_24903);
nor U25619 (N_25619,N_24056,N_24013);
nand U25620 (N_25620,N_24492,N_24416);
nand U25621 (N_25621,N_25163,N_24963);
xor U25622 (N_25622,N_24786,N_24343);
nor U25623 (N_25623,N_24275,N_24948);
or U25624 (N_25624,N_24609,N_24362);
and U25625 (N_25625,N_24431,N_24398);
or U25626 (N_25626,N_24742,N_24023);
nor U25627 (N_25627,N_25159,N_24556);
xnor U25628 (N_25628,N_24900,N_24625);
or U25629 (N_25629,N_24642,N_24511);
nand U25630 (N_25630,N_24713,N_24942);
or U25631 (N_25631,N_24145,N_24935);
nand U25632 (N_25632,N_24514,N_24666);
and U25633 (N_25633,N_24180,N_24628);
and U25634 (N_25634,N_24176,N_24569);
xnor U25635 (N_25635,N_24728,N_24112);
or U25636 (N_25636,N_24499,N_24824);
or U25637 (N_25637,N_24692,N_24161);
and U25638 (N_25638,N_24820,N_24172);
nand U25639 (N_25639,N_24854,N_24975);
nand U25640 (N_25640,N_25165,N_24596);
or U25641 (N_25641,N_25121,N_24359);
nor U25642 (N_25642,N_25026,N_24255);
xor U25643 (N_25643,N_24964,N_24706);
or U25644 (N_25644,N_25145,N_24496);
nand U25645 (N_25645,N_24185,N_24604);
nand U25646 (N_25646,N_24715,N_24528);
nor U25647 (N_25647,N_25123,N_24559);
and U25648 (N_25648,N_24925,N_24913);
and U25649 (N_25649,N_24188,N_24328);
xnor U25650 (N_25650,N_25093,N_24857);
or U25651 (N_25651,N_24619,N_24908);
and U25652 (N_25652,N_24968,N_24249);
and U25653 (N_25653,N_24670,N_24422);
nand U25654 (N_25654,N_24223,N_24088);
or U25655 (N_25655,N_24611,N_24215);
or U25656 (N_25656,N_24446,N_25158);
and U25657 (N_25657,N_24068,N_24067);
or U25658 (N_25658,N_24027,N_24329);
nor U25659 (N_25659,N_24653,N_24509);
nor U25660 (N_25660,N_24558,N_24591);
or U25661 (N_25661,N_24956,N_24260);
nor U25662 (N_25662,N_25148,N_24053);
nand U25663 (N_25663,N_24399,N_24408);
xor U25664 (N_25664,N_24875,N_24889);
nor U25665 (N_25665,N_24823,N_25128);
nand U25666 (N_25666,N_24860,N_24309);
nor U25667 (N_25667,N_24015,N_24805);
nand U25668 (N_25668,N_24150,N_24052);
xnor U25669 (N_25669,N_24310,N_24407);
or U25670 (N_25670,N_24266,N_24661);
xnor U25671 (N_25671,N_25096,N_24133);
and U25672 (N_25672,N_24139,N_24480);
nand U25673 (N_25673,N_24777,N_24461);
or U25674 (N_25674,N_24089,N_24673);
and U25675 (N_25675,N_24778,N_24493);
nor U25676 (N_25676,N_24460,N_24859);
nand U25677 (N_25677,N_25050,N_24691);
xor U25678 (N_25678,N_24995,N_24326);
nor U25679 (N_25679,N_25150,N_24738);
nand U25680 (N_25680,N_24520,N_24108);
nand U25681 (N_25681,N_24722,N_24231);
or U25682 (N_25682,N_25052,N_24753);
or U25683 (N_25683,N_25008,N_24182);
or U25684 (N_25684,N_24743,N_24954);
or U25685 (N_25685,N_25038,N_24256);
xor U25686 (N_25686,N_24787,N_24500);
xor U25687 (N_25687,N_24032,N_24893);
nand U25688 (N_25688,N_24969,N_24283);
nor U25689 (N_25689,N_25002,N_25142);
nand U25690 (N_25690,N_24977,N_24767);
nand U25691 (N_25691,N_25097,N_24663);
xor U25692 (N_25692,N_24114,N_24978);
and U25693 (N_25693,N_24474,N_24485);
and U25694 (N_25694,N_25087,N_24725);
xnor U25695 (N_25695,N_24155,N_24322);
nand U25696 (N_25696,N_24803,N_24891);
and U25697 (N_25697,N_24847,N_24085);
nand U25698 (N_25698,N_24239,N_24084);
and U25699 (N_25699,N_24448,N_25102);
xnor U25700 (N_25700,N_24593,N_24127);
nor U25701 (N_25701,N_25025,N_24059);
nor U25702 (N_25702,N_24894,N_24588);
and U25703 (N_25703,N_24843,N_24043);
or U25704 (N_25704,N_24332,N_24271);
and U25705 (N_25705,N_25168,N_24519);
or U25706 (N_25706,N_25067,N_24744);
or U25707 (N_25707,N_24351,N_24866);
nor U25708 (N_25708,N_24967,N_24379);
or U25709 (N_25709,N_24627,N_24421);
xnor U25710 (N_25710,N_25134,N_25143);
or U25711 (N_25711,N_25009,N_24901);
and U25712 (N_25712,N_25043,N_24179);
and U25713 (N_25713,N_24044,N_24471);
nand U25714 (N_25714,N_24776,N_24536);
nor U25715 (N_25715,N_24324,N_24996);
nand U25716 (N_25716,N_24284,N_24469);
or U25717 (N_25717,N_24259,N_24729);
and U25718 (N_25718,N_24221,N_24946);
nand U25719 (N_25719,N_24131,N_24140);
nor U25720 (N_25720,N_24912,N_24614);
nor U25721 (N_25721,N_24575,N_24871);
or U25722 (N_25722,N_25054,N_25053);
nor U25723 (N_25723,N_24289,N_24863);
or U25724 (N_25724,N_24644,N_24135);
nor U25725 (N_25725,N_25177,N_24616);
or U25726 (N_25726,N_24166,N_25033);
nor U25727 (N_25727,N_24809,N_24513);
xor U25728 (N_25728,N_24671,N_24438);
or U25729 (N_25729,N_24302,N_24033);
and U25730 (N_25730,N_25086,N_24953);
nor U25731 (N_25731,N_24443,N_24061);
nor U25732 (N_25732,N_24312,N_24506);
and U25733 (N_25733,N_24907,N_25076);
nand U25734 (N_25734,N_24723,N_25110);
nand U25735 (N_25735,N_24177,N_25049);
or U25736 (N_25736,N_25085,N_24501);
and U25737 (N_25737,N_24764,N_24937);
nand U25738 (N_25738,N_24883,N_24453);
and U25739 (N_25739,N_24829,N_24238);
or U25740 (N_25740,N_24910,N_24987);
nor U25741 (N_25741,N_24643,N_25042);
nand U25742 (N_25742,N_24517,N_24755);
nand U25743 (N_25743,N_24822,N_24909);
nand U25744 (N_25744,N_24674,N_24950);
and U25745 (N_25745,N_24784,N_25091);
nor U25746 (N_25746,N_24060,N_25139);
nand U25747 (N_25747,N_24693,N_24541);
nand U25748 (N_25748,N_25194,N_24816);
and U25749 (N_25749,N_24411,N_24234);
and U25750 (N_25750,N_24915,N_24354);
nor U25751 (N_25751,N_24918,N_24402);
nand U25752 (N_25752,N_25193,N_24549);
xor U25753 (N_25753,N_24992,N_24361);
nor U25754 (N_25754,N_25192,N_24169);
and U25755 (N_25755,N_24607,N_24254);
nand U25756 (N_25756,N_24686,N_24759);
and U25757 (N_25757,N_24340,N_24730);
and U25758 (N_25758,N_24882,N_24927);
nand U25759 (N_25759,N_24548,N_24652);
and U25760 (N_25760,N_25197,N_24481);
xnor U25761 (N_25761,N_24376,N_24382);
xnor U25762 (N_25762,N_24039,N_24395);
nand U25763 (N_25763,N_24895,N_24981);
and U25764 (N_25764,N_25060,N_24036);
nand U25765 (N_25765,N_24566,N_24545);
and U25766 (N_25766,N_25092,N_24192);
or U25767 (N_25767,N_24280,N_24317);
nand U25768 (N_25768,N_25035,N_24681);
xnor U25769 (N_25769,N_25061,N_24194);
or U25770 (N_25770,N_24986,N_24115);
nand U25771 (N_25771,N_24440,N_24128);
nand U25772 (N_25772,N_24699,N_25119);
and U25773 (N_25773,N_25149,N_24679);
nor U25774 (N_25774,N_25169,N_24024);
or U25775 (N_25775,N_24851,N_24724);
xnor U25776 (N_25776,N_24122,N_25077);
nor U25777 (N_25777,N_24874,N_25140);
nand U25778 (N_25778,N_24917,N_24121);
and U25779 (N_25779,N_24434,N_25079);
xor U25780 (N_25780,N_24028,N_24077);
nand U25781 (N_25781,N_24323,N_24571);
or U25782 (N_25782,N_24087,N_24719);
nor U25783 (N_25783,N_24698,N_24080);
xnor U25784 (N_25784,N_24839,N_24111);
nor U25785 (N_25785,N_24358,N_24865);
nand U25786 (N_25786,N_24230,N_25156);
and U25787 (N_25787,N_24846,N_24648);
and U25788 (N_25788,N_24790,N_24690);
or U25789 (N_25789,N_24141,N_24718);
and U25790 (N_25790,N_24793,N_24792);
or U25791 (N_25791,N_25174,N_25051);
xor U25792 (N_25792,N_25046,N_24530);
or U25793 (N_25793,N_24136,N_24819);
and U25794 (N_25794,N_25048,N_25027);
or U25795 (N_25795,N_24705,N_25103);
and U25796 (N_25796,N_25112,N_24007);
nand U25797 (N_25797,N_24008,N_24766);
nand U25798 (N_25798,N_24311,N_25115);
and U25799 (N_25799,N_25185,N_24654);
nand U25800 (N_25800,N_24631,N_24222);
nand U25801 (N_25801,N_24322,N_24409);
nand U25802 (N_25802,N_24769,N_24396);
and U25803 (N_25803,N_25162,N_24866);
and U25804 (N_25804,N_24809,N_24742);
nor U25805 (N_25805,N_25180,N_24606);
and U25806 (N_25806,N_24991,N_24620);
xor U25807 (N_25807,N_24099,N_24935);
nand U25808 (N_25808,N_24796,N_24578);
nor U25809 (N_25809,N_24279,N_24384);
and U25810 (N_25810,N_25094,N_24346);
nor U25811 (N_25811,N_24079,N_24403);
nor U25812 (N_25812,N_24733,N_24570);
nand U25813 (N_25813,N_24996,N_24302);
xor U25814 (N_25814,N_25032,N_25031);
or U25815 (N_25815,N_24579,N_24192);
nor U25816 (N_25816,N_24159,N_24536);
nor U25817 (N_25817,N_25112,N_25181);
xor U25818 (N_25818,N_24318,N_24307);
nor U25819 (N_25819,N_24429,N_24040);
or U25820 (N_25820,N_24071,N_25003);
or U25821 (N_25821,N_25068,N_24475);
and U25822 (N_25822,N_24786,N_24566);
and U25823 (N_25823,N_24978,N_24802);
nand U25824 (N_25824,N_24590,N_24860);
nor U25825 (N_25825,N_24402,N_24397);
nand U25826 (N_25826,N_24435,N_24907);
or U25827 (N_25827,N_25063,N_24540);
and U25828 (N_25828,N_24996,N_24958);
nor U25829 (N_25829,N_24243,N_24497);
nand U25830 (N_25830,N_24883,N_25000);
nor U25831 (N_25831,N_24294,N_24328);
or U25832 (N_25832,N_25110,N_24742);
xor U25833 (N_25833,N_24537,N_24270);
and U25834 (N_25834,N_24386,N_24170);
nor U25835 (N_25835,N_24405,N_24513);
xor U25836 (N_25836,N_24854,N_24179);
and U25837 (N_25837,N_24611,N_24832);
and U25838 (N_25838,N_24009,N_24998);
xnor U25839 (N_25839,N_25083,N_24790);
or U25840 (N_25840,N_24518,N_24428);
xor U25841 (N_25841,N_24147,N_24860);
nor U25842 (N_25842,N_25062,N_24393);
nand U25843 (N_25843,N_24718,N_24859);
nor U25844 (N_25844,N_24891,N_25011);
nand U25845 (N_25845,N_25107,N_24882);
nand U25846 (N_25846,N_24369,N_24438);
nand U25847 (N_25847,N_24705,N_24723);
nor U25848 (N_25848,N_24127,N_24300);
xor U25849 (N_25849,N_24067,N_24456);
nor U25850 (N_25850,N_24100,N_24514);
nor U25851 (N_25851,N_24503,N_24044);
and U25852 (N_25852,N_25191,N_24913);
nand U25853 (N_25853,N_24150,N_24740);
and U25854 (N_25854,N_24230,N_25107);
and U25855 (N_25855,N_24273,N_24788);
nor U25856 (N_25856,N_24244,N_24875);
xnor U25857 (N_25857,N_24171,N_24061);
or U25858 (N_25858,N_24299,N_24061);
and U25859 (N_25859,N_24172,N_24131);
or U25860 (N_25860,N_24349,N_24631);
xnor U25861 (N_25861,N_24370,N_25159);
or U25862 (N_25862,N_24485,N_25099);
xor U25863 (N_25863,N_24323,N_24054);
or U25864 (N_25864,N_24065,N_24796);
nand U25865 (N_25865,N_24230,N_24674);
nand U25866 (N_25866,N_25184,N_24839);
or U25867 (N_25867,N_24157,N_24091);
xor U25868 (N_25868,N_24272,N_24447);
nand U25869 (N_25869,N_24717,N_24227);
nand U25870 (N_25870,N_24855,N_24101);
nor U25871 (N_25871,N_24680,N_24412);
xor U25872 (N_25872,N_24644,N_24660);
nor U25873 (N_25873,N_24752,N_24211);
xnor U25874 (N_25874,N_24859,N_24409);
nand U25875 (N_25875,N_24207,N_24587);
nand U25876 (N_25876,N_24567,N_24318);
and U25877 (N_25877,N_24856,N_24918);
nor U25878 (N_25878,N_24972,N_25117);
nor U25879 (N_25879,N_24339,N_24147);
and U25880 (N_25880,N_24650,N_25088);
or U25881 (N_25881,N_24353,N_24025);
xnor U25882 (N_25882,N_24126,N_24357);
nand U25883 (N_25883,N_24660,N_24205);
nor U25884 (N_25884,N_25165,N_24161);
nor U25885 (N_25885,N_24003,N_24011);
nand U25886 (N_25886,N_24820,N_24046);
nor U25887 (N_25887,N_24327,N_24254);
nand U25888 (N_25888,N_24760,N_24806);
nor U25889 (N_25889,N_25116,N_24272);
nand U25890 (N_25890,N_24996,N_24797);
nand U25891 (N_25891,N_24174,N_25100);
nand U25892 (N_25892,N_24259,N_25075);
nor U25893 (N_25893,N_25093,N_25028);
nor U25894 (N_25894,N_24510,N_24577);
nand U25895 (N_25895,N_24308,N_24201);
nand U25896 (N_25896,N_24967,N_24495);
nor U25897 (N_25897,N_24171,N_24292);
xor U25898 (N_25898,N_25092,N_24315);
nand U25899 (N_25899,N_24170,N_24455);
xnor U25900 (N_25900,N_24659,N_24127);
nand U25901 (N_25901,N_24500,N_24247);
and U25902 (N_25902,N_24287,N_24364);
or U25903 (N_25903,N_24944,N_24120);
xor U25904 (N_25904,N_25098,N_24073);
and U25905 (N_25905,N_24637,N_24113);
nor U25906 (N_25906,N_25147,N_24499);
nor U25907 (N_25907,N_24377,N_24544);
nor U25908 (N_25908,N_25176,N_24832);
and U25909 (N_25909,N_24838,N_24980);
nor U25910 (N_25910,N_24432,N_24083);
nor U25911 (N_25911,N_24756,N_24063);
nand U25912 (N_25912,N_25003,N_24589);
and U25913 (N_25913,N_24760,N_24591);
nor U25914 (N_25914,N_24773,N_24081);
and U25915 (N_25915,N_24697,N_24788);
nand U25916 (N_25916,N_24560,N_24244);
and U25917 (N_25917,N_24286,N_24967);
and U25918 (N_25918,N_24456,N_24020);
xnor U25919 (N_25919,N_24993,N_24179);
or U25920 (N_25920,N_24695,N_24512);
nand U25921 (N_25921,N_24776,N_25027);
nor U25922 (N_25922,N_24392,N_24144);
and U25923 (N_25923,N_24892,N_24376);
and U25924 (N_25924,N_24345,N_24204);
or U25925 (N_25925,N_24819,N_24931);
nand U25926 (N_25926,N_25043,N_24335);
nor U25927 (N_25927,N_24087,N_25197);
nor U25928 (N_25928,N_24847,N_24257);
and U25929 (N_25929,N_24138,N_24624);
nand U25930 (N_25930,N_24695,N_24700);
or U25931 (N_25931,N_25137,N_24488);
and U25932 (N_25932,N_24967,N_24859);
or U25933 (N_25933,N_24931,N_24871);
or U25934 (N_25934,N_24156,N_24419);
xnor U25935 (N_25935,N_24096,N_24495);
nand U25936 (N_25936,N_24987,N_24259);
xor U25937 (N_25937,N_24184,N_24697);
nand U25938 (N_25938,N_25166,N_24598);
nand U25939 (N_25939,N_24696,N_24813);
xnor U25940 (N_25940,N_24223,N_24316);
or U25941 (N_25941,N_24764,N_25025);
and U25942 (N_25942,N_24196,N_24652);
or U25943 (N_25943,N_24941,N_25191);
or U25944 (N_25944,N_24287,N_24670);
or U25945 (N_25945,N_24433,N_24173);
nand U25946 (N_25946,N_24859,N_24165);
and U25947 (N_25947,N_24384,N_24096);
nor U25948 (N_25948,N_24271,N_24142);
and U25949 (N_25949,N_24337,N_24140);
nand U25950 (N_25950,N_24616,N_25135);
nand U25951 (N_25951,N_24988,N_24006);
nor U25952 (N_25952,N_24462,N_24913);
nor U25953 (N_25953,N_24967,N_24370);
xnor U25954 (N_25954,N_24556,N_24400);
nand U25955 (N_25955,N_24135,N_25049);
nor U25956 (N_25956,N_24405,N_24577);
xnor U25957 (N_25957,N_25126,N_24360);
nand U25958 (N_25958,N_24459,N_24177);
and U25959 (N_25959,N_25190,N_24813);
and U25960 (N_25960,N_24014,N_24364);
nand U25961 (N_25961,N_25002,N_24730);
or U25962 (N_25962,N_24888,N_24918);
and U25963 (N_25963,N_24389,N_24854);
nor U25964 (N_25964,N_24247,N_24205);
nand U25965 (N_25965,N_24605,N_24616);
xnor U25966 (N_25966,N_24037,N_24702);
nor U25967 (N_25967,N_24730,N_24613);
or U25968 (N_25968,N_24162,N_24978);
and U25969 (N_25969,N_24495,N_24663);
and U25970 (N_25970,N_24980,N_24214);
xor U25971 (N_25971,N_24029,N_24160);
nor U25972 (N_25972,N_24402,N_24027);
and U25973 (N_25973,N_24994,N_24415);
nand U25974 (N_25974,N_24381,N_25079);
nand U25975 (N_25975,N_24011,N_24290);
xor U25976 (N_25976,N_24698,N_24458);
nand U25977 (N_25977,N_24005,N_24683);
xor U25978 (N_25978,N_24457,N_24218);
nand U25979 (N_25979,N_24053,N_24159);
xnor U25980 (N_25980,N_24009,N_24751);
xnor U25981 (N_25981,N_24374,N_24608);
and U25982 (N_25982,N_24423,N_24506);
or U25983 (N_25983,N_24454,N_24425);
xnor U25984 (N_25984,N_25025,N_24102);
and U25985 (N_25985,N_24555,N_24549);
nand U25986 (N_25986,N_24252,N_24079);
or U25987 (N_25987,N_24268,N_24887);
nand U25988 (N_25988,N_25039,N_25106);
nor U25989 (N_25989,N_24190,N_24484);
nand U25990 (N_25990,N_24392,N_24053);
xnor U25991 (N_25991,N_24705,N_24579);
or U25992 (N_25992,N_24184,N_24274);
nor U25993 (N_25993,N_25114,N_24189);
or U25994 (N_25994,N_24328,N_24585);
and U25995 (N_25995,N_24973,N_24389);
and U25996 (N_25996,N_24140,N_24791);
xnor U25997 (N_25997,N_24954,N_24226);
nor U25998 (N_25998,N_24688,N_25128);
nor U25999 (N_25999,N_24464,N_24467);
nor U26000 (N_26000,N_24637,N_25168);
nand U26001 (N_26001,N_24240,N_24766);
or U26002 (N_26002,N_24356,N_25125);
nand U26003 (N_26003,N_24513,N_24508);
nor U26004 (N_26004,N_24261,N_24943);
or U26005 (N_26005,N_24256,N_24110);
nor U26006 (N_26006,N_25015,N_25027);
nor U26007 (N_26007,N_24125,N_25076);
nand U26008 (N_26008,N_24064,N_24026);
or U26009 (N_26009,N_24497,N_25072);
xor U26010 (N_26010,N_24996,N_24474);
or U26011 (N_26011,N_24604,N_24380);
nand U26012 (N_26012,N_24236,N_24473);
or U26013 (N_26013,N_24549,N_24353);
or U26014 (N_26014,N_24785,N_24845);
nor U26015 (N_26015,N_24695,N_24187);
nand U26016 (N_26016,N_24369,N_24687);
nor U26017 (N_26017,N_24079,N_24331);
xor U26018 (N_26018,N_24580,N_24427);
xnor U26019 (N_26019,N_24076,N_25058);
xor U26020 (N_26020,N_24875,N_25003);
and U26021 (N_26021,N_25087,N_24336);
and U26022 (N_26022,N_24913,N_25031);
xnor U26023 (N_26023,N_24731,N_24732);
nor U26024 (N_26024,N_24464,N_24421);
nor U26025 (N_26025,N_24070,N_24506);
nand U26026 (N_26026,N_25175,N_24089);
and U26027 (N_26027,N_24343,N_24513);
nand U26028 (N_26028,N_24748,N_24668);
and U26029 (N_26029,N_24249,N_24736);
and U26030 (N_26030,N_24278,N_24949);
nor U26031 (N_26031,N_24872,N_25088);
nand U26032 (N_26032,N_24411,N_24521);
xnor U26033 (N_26033,N_25025,N_24319);
xnor U26034 (N_26034,N_24982,N_24608);
xor U26035 (N_26035,N_25006,N_24991);
nand U26036 (N_26036,N_24313,N_24525);
nor U26037 (N_26037,N_24676,N_24536);
nand U26038 (N_26038,N_24376,N_24783);
nand U26039 (N_26039,N_24889,N_24809);
xor U26040 (N_26040,N_24957,N_25030);
or U26041 (N_26041,N_24751,N_25053);
and U26042 (N_26042,N_24540,N_24740);
and U26043 (N_26043,N_24080,N_25171);
or U26044 (N_26044,N_24439,N_24609);
or U26045 (N_26045,N_24335,N_24595);
and U26046 (N_26046,N_24007,N_24116);
xor U26047 (N_26047,N_25000,N_24888);
and U26048 (N_26048,N_24149,N_24290);
nor U26049 (N_26049,N_25106,N_24263);
nor U26050 (N_26050,N_24150,N_24287);
or U26051 (N_26051,N_24170,N_25040);
and U26052 (N_26052,N_25105,N_24438);
and U26053 (N_26053,N_24654,N_25150);
or U26054 (N_26054,N_24745,N_24160);
and U26055 (N_26055,N_24753,N_24684);
xnor U26056 (N_26056,N_24731,N_24809);
or U26057 (N_26057,N_24850,N_24057);
nor U26058 (N_26058,N_24138,N_25094);
nor U26059 (N_26059,N_24282,N_24292);
and U26060 (N_26060,N_24345,N_25019);
or U26061 (N_26061,N_24917,N_24783);
nand U26062 (N_26062,N_24372,N_24857);
nand U26063 (N_26063,N_24151,N_25001);
xor U26064 (N_26064,N_25032,N_25158);
nand U26065 (N_26065,N_24345,N_24961);
or U26066 (N_26066,N_24076,N_24237);
and U26067 (N_26067,N_24649,N_24356);
nand U26068 (N_26068,N_24240,N_24946);
or U26069 (N_26069,N_25193,N_25186);
and U26070 (N_26070,N_24560,N_24624);
xnor U26071 (N_26071,N_25021,N_24057);
and U26072 (N_26072,N_24068,N_24525);
xor U26073 (N_26073,N_24699,N_24437);
and U26074 (N_26074,N_24253,N_24489);
or U26075 (N_26075,N_24028,N_24337);
nor U26076 (N_26076,N_24342,N_24486);
or U26077 (N_26077,N_24416,N_24986);
or U26078 (N_26078,N_25024,N_24515);
nand U26079 (N_26079,N_25022,N_24491);
xor U26080 (N_26080,N_24270,N_25044);
xor U26081 (N_26081,N_25097,N_24614);
nand U26082 (N_26082,N_24938,N_24828);
and U26083 (N_26083,N_24507,N_24518);
xnor U26084 (N_26084,N_24217,N_24463);
nand U26085 (N_26085,N_24824,N_24560);
nand U26086 (N_26086,N_24383,N_24680);
or U26087 (N_26087,N_24799,N_24514);
and U26088 (N_26088,N_24301,N_24026);
xnor U26089 (N_26089,N_24519,N_24882);
xor U26090 (N_26090,N_24936,N_24165);
xor U26091 (N_26091,N_24574,N_24146);
nand U26092 (N_26092,N_25067,N_24432);
and U26093 (N_26093,N_24031,N_24463);
and U26094 (N_26094,N_25149,N_24515);
xor U26095 (N_26095,N_24926,N_25117);
or U26096 (N_26096,N_24824,N_25023);
or U26097 (N_26097,N_24395,N_24604);
and U26098 (N_26098,N_25180,N_25020);
and U26099 (N_26099,N_24600,N_24168);
or U26100 (N_26100,N_24467,N_24183);
and U26101 (N_26101,N_24829,N_24706);
xor U26102 (N_26102,N_25180,N_24911);
nor U26103 (N_26103,N_25076,N_25136);
xor U26104 (N_26104,N_24417,N_24732);
and U26105 (N_26105,N_24758,N_24388);
nand U26106 (N_26106,N_24018,N_24474);
or U26107 (N_26107,N_24209,N_25048);
nand U26108 (N_26108,N_24541,N_24859);
xor U26109 (N_26109,N_25036,N_24071);
or U26110 (N_26110,N_24438,N_24308);
xor U26111 (N_26111,N_24372,N_24701);
and U26112 (N_26112,N_24153,N_24112);
xor U26113 (N_26113,N_24512,N_24989);
or U26114 (N_26114,N_24491,N_24104);
or U26115 (N_26115,N_25063,N_24582);
and U26116 (N_26116,N_24909,N_24091);
and U26117 (N_26117,N_24587,N_24569);
xor U26118 (N_26118,N_24667,N_24556);
or U26119 (N_26119,N_24765,N_24317);
or U26120 (N_26120,N_24304,N_24863);
xnor U26121 (N_26121,N_24459,N_24568);
and U26122 (N_26122,N_24576,N_24395);
or U26123 (N_26123,N_24912,N_24360);
nor U26124 (N_26124,N_24426,N_24979);
xnor U26125 (N_26125,N_24966,N_24753);
nand U26126 (N_26126,N_25039,N_24911);
nand U26127 (N_26127,N_24091,N_24015);
xnor U26128 (N_26128,N_24658,N_24694);
nor U26129 (N_26129,N_24568,N_24343);
or U26130 (N_26130,N_24292,N_24039);
or U26131 (N_26131,N_24136,N_24124);
nor U26132 (N_26132,N_24441,N_25081);
and U26133 (N_26133,N_24798,N_25020);
nand U26134 (N_26134,N_24783,N_24645);
nand U26135 (N_26135,N_24239,N_25114);
or U26136 (N_26136,N_24240,N_24649);
xnor U26137 (N_26137,N_24660,N_24118);
or U26138 (N_26138,N_24871,N_24973);
nand U26139 (N_26139,N_24764,N_24824);
nor U26140 (N_26140,N_24891,N_24646);
xor U26141 (N_26141,N_25035,N_25081);
and U26142 (N_26142,N_24528,N_24705);
and U26143 (N_26143,N_25107,N_24904);
nor U26144 (N_26144,N_24329,N_24425);
and U26145 (N_26145,N_24640,N_24397);
nand U26146 (N_26146,N_24975,N_24266);
and U26147 (N_26147,N_24230,N_24752);
xnor U26148 (N_26148,N_24480,N_24742);
nand U26149 (N_26149,N_24346,N_24055);
and U26150 (N_26150,N_25173,N_24860);
xor U26151 (N_26151,N_24870,N_25038);
nand U26152 (N_26152,N_25038,N_24451);
and U26153 (N_26153,N_24508,N_24992);
and U26154 (N_26154,N_24981,N_24739);
or U26155 (N_26155,N_24378,N_24374);
or U26156 (N_26156,N_24285,N_24923);
nand U26157 (N_26157,N_24173,N_24335);
xor U26158 (N_26158,N_24196,N_24282);
xor U26159 (N_26159,N_25152,N_24582);
or U26160 (N_26160,N_25119,N_24356);
xor U26161 (N_26161,N_25114,N_24961);
nand U26162 (N_26162,N_24314,N_25092);
nor U26163 (N_26163,N_24381,N_25026);
xnor U26164 (N_26164,N_24743,N_24426);
or U26165 (N_26165,N_24826,N_24425);
or U26166 (N_26166,N_24520,N_24469);
and U26167 (N_26167,N_24765,N_24154);
and U26168 (N_26168,N_24965,N_24155);
xnor U26169 (N_26169,N_25036,N_24029);
nor U26170 (N_26170,N_24923,N_24034);
and U26171 (N_26171,N_24670,N_24564);
nor U26172 (N_26172,N_24767,N_24381);
nor U26173 (N_26173,N_24064,N_24417);
and U26174 (N_26174,N_24067,N_24085);
or U26175 (N_26175,N_24369,N_24810);
xor U26176 (N_26176,N_24646,N_24474);
nand U26177 (N_26177,N_24930,N_25116);
nand U26178 (N_26178,N_24975,N_24478);
and U26179 (N_26179,N_25011,N_24004);
nand U26180 (N_26180,N_24621,N_24420);
or U26181 (N_26181,N_24714,N_24419);
nor U26182 (N_26182,N_24509,N_24193);
xor U26183 (N_26183,N_25139,N_24687);
nor U26184 (N_26184,N_25169,N_24983);
or U26185 (N_26185,N_24427,N_25062);
xor U26186 (N_26186,N_24380,N_25063);
nor U26187 (N_26187,N_24824,N_24095);
or U26188 (N_26188,N_24364,N_24767);
and U26189 (N_26189,N_24119,N_24344);
xnor U26190 (N_26190,N_24556,N_24919);
or U26191 (N_26191,N_24840,N_24362);
or U26192 (N_26192,N_24239,N_24601);
nand U26193 (N_26193,N_24560,N_24901);
nor U26194 (N_26194,N_24234,N_24987);
xor U26195 (N_26195,N_24597,N_24249);
and U26196 (N_26196,N_25184,N_24680);
and U26197 (N_26197,N_24623,N_24955);
nand U26198 (N_26198,N_24555,N_24270);
nor U26199 (N_26199,N_24006,N_25127);
xor U26200 (N_26200,N_24809,N_24535);
nor U26201 (N_26201,N_24538,N_24497);
xnor U26202 (N_26202,N_24760,N_24922);
or U26203 (N_26203,N_24850,N_24453);
nor U26204 (N_26204,N_24904,N_24014);
or U26205 (N_26205,N_24798,N_24247);
nand U26206 (N_26206,N_24114,N_24004);
and U26207 (N_26207,N_25121,N_24205);
xnor U26208 (N_26208,N_24184,N_24405);
nor U26209 (N_26209,N_25113,N_24261);
nor U26210 (N_26210,N_24687,N_24459);
xnor U26211 (N_26211,N_24935,N_24452);
nor U26212 (N_26212,N_24343,N_25029);
and U26213 (N_26213,N_25129,N_25099);
nor U26214 (N_26214,N_24228,N_24293);
or U26215 (N_26215,N_24160,N_24996);
nor U26216 (N_26216,N_24041,N_24099);
nand U26217 (N_26217,N_24983,N_24230);
nor U26218 (N_26218,N_25130,N_24341);
and U26219 (N_26219,N_24637,N_24377);
and U26220 (N_26220,N_24884,N_24932);
xor U26221 (N_26221,N_24367,N_24659);
and U26222 (N_26222,N_24127,N_24428);
nor U26223 (N_26223,N_24740,N_24028);
nor U26224 (N_26224,N_24221,N_24861);
nand U26225 (N_26225,N_24407,N_24488);
and U26226 (N_26226,N_24990,N_24635);
nor U26227 (N_26227,N_24575,N_24306);
or U26228 (N_26228,N_25019,N_24302);
or U26229 (N_26229,N_24377,N_24463);
nor U26230 (N_26230,N_24471,N_25100);
xor U26231 (N_26231,N_24631,N_24264);
or U26232 (N_26232,N_24889,N_25078);
or U26233 (N_26233,N_25153,N_24960);
nand U26234 (N_26234,N_24388,N_24947);
xnor U26235 (N_26235,N_24866,N_24672);
nor U26236 (N_26236,N_24150,N_24717);
nand U26237 (N_26237,N_24976,N_25164);
nand U26238 (N_26238,N_24292,N_24831);
and U26239 (N_26239,N_24025,N_24922);
nor U26240 (N_26240,N_24073,N_24378);
or U26241 (N_26241,N_24417,N_24967);
nor U26242 (N_26242,N_24533,N_25173);
xnor U26243 (N_26243,N_24056,N_24491);
nand U26244 (N_26244,N_24900,N_24141);
and U26245 (N_26245,N_24736,N_25115);
xor U26246 (N_26246,N_25020,N_24421);
xnor U26247 (N_26247,N_24578,N_24063);
or U26248 (N_26248,N_24023,N_24743);
or U26249 (N_26249,N_24034,N_24161);
or U26250 (N_26250,N_24431,N_25071);
xnor U26251 (N_26251,N_24750,N_24920);
nand U26252 (N_26252,N_25117,N_24683);
and U26253 (N_26253,N_25041,N_25148);
or U26254 (N_26254,N_24048,N_25098);
nor U26255 (N_26255,N_24189,N_24170);
or U26256 (N_26256,N_24133,N_24326);
and U26257 (N_26257,N_24970,N_24026);
nand U26258 (N_26258,N_24080,N_25140);
xor U26259 (N_26259,N_24281,N_24873);
nand U26260 (N_26260,N_24491,N_25171);
nand U26261 (N_26261,N_24832,N_24051);
or U26262 (N_26262,N_24201,N_24331);
or U26263 (N_26263,N_24833,N_24782);
xor U26264 (N_26264,N_25047,N_24516);
and U26265 (N_26265,N_24518,N_24670);
nor U26266 (N_26266,N_24723,N_24262);
xnor U26267 (N_26267,N_24983,N_24034);
or U26268 (N_26268,N_24606,N_24535);
xnor U26269 (N_26269,N_25037,N_24153);
xor U26270 (N_26270,N_24185,N_24638);
nand U26271 (N_26271,N_24094,N_24340);
nand U26272 (N_26272,N_24492,N_24930);
or U26273 (N_26273,N_25149,N_24325);
xor U26274 (N_26274,N_24397,N_24240);
xnor U26275 (N_26275,N_25063,N_24713);
or U26276 (N_26276,N_24990,N_24085);
xnor U26277 (N_26277,N_24473,N_24965);
and U26278 (N_26278,N_24685,N_25073);
xor U26279 (N_26279,N_24867,N_24979);
nand U26280 (N_26280,N_24713,N_24259);
or U26281 (N_26281,N_25036,N_24612);
nand U26282 (N_26282,N_24697,N_24428);
and U26283 (N_26283,N_24612,N_25052);
nand U26284 (N_26284,N_24412,N_24728);
nand U26285 (N_26285,N_24871,N_25104);
and U26286 (N_26286,N_25118,N_24155);
nand U26287 (N_26287,N_24838,N_24297);
and U26288 (N_26288,N_25174,N_24898);
nand U26289 (N_26289,N_25008,N_24819);
and U26290 (N_26290,N_25187,N_24063);
or U26291 (N_26291,N_24259,N_24180);
nand U26292 (N_26292,N_24047,N_24540);
or U26293 (N_26293,N_24139,N_24733);
nand U26294 (N_26294,N_24502,N_24421);
xor U26295 (N_26295,N_24729,N_25115);
or U26296 (N_26296,N_24231,N_24447);
and U26297 (N_26297,N_24248,N_24823);
nor U26298 (N_26298,N_24494,N_24760);
and U26299 (N_26299,N_25107,N_24284);
nor U26300 (N_26300,N_24105,N_24877);
nand U26301 (N_26301,N_24404,N_24068);
nor U26302 (N_26302,N_25055,N_25161);
and U26303 (N_26303,N_25015,N_24530);
and U26304 (N_26304,N_24542,N_24921);
or U26305 (N_26305,N_24825,N_25053);
or U26306 (N_26306,N_25179,N_24583);
nand U26307 (N_26307,N_24193,N_24296);
nand U26308 (N_26308,N_25026,N_24195);
xor U26309 (N_26309,N_24152,N_24806);
nand U26310 (N_26310,N_24081,N_24847);
nor U26311 (N_26311,N_24746,N_25088);
or U26312 (N_26312,N_24774,N_24894);
or U26313 (N_26313,N_25177,N_24309);
or U26314 (N_26314,N_24749,N_24486);
and U26315 (N_26315,N_24785,N_24064);
xor U26316 (N_26316,N_24348,N_24538);
or U26317 (N_26317,N_25120,N_24622);
nor U26318 (N_26318,N_24802,N_24762);
nor U26319 (N_26319,N_24548,N_24312);
or U26320 (N_26320,N_24088,N_24940);
and U26321 (N_26321,N_24357,N_25190);
xor U26322 (N_26322,N_24626,N_24506);
nor U26323 (N_26323,N_25115,N_24152);
nor U26324 (N_26324,N_24867,N_24053);
nand U26325 (N_26325,N_25088,N_24859);
or U26326 (N_26326,N_24274,N_24424);
xnor U26327 (N_26327,N_24527,N_25166);
xor U26328 (N_26328,N_24425,N_24209);
and U26329 (N_26329,N_24517,N_24506);
or U26330 (N_26330,N_24245,N_24504);
nand U26331 (N_26331,N_24214,N_24102);
nand U26332 (N_26332,N_24620,N_24117);
and U26333 (N_26333,N_24269,N_24707);
or U26334 (N_26334,N_24616,N_24413);
nand U26335 (N_26335,N_24429,N_24101);
or U26336 (N_26336,N_24415,N_24413);
or U26337 (N_26337,N_24057,N_24349);
and U26338 (N_26338,N_25150,N_24559);
xnor U26339 (N_26339,N_24745,N_24775);
nor U26340 (N_26340,N_24015,N_24747);
xnor U26341 (N_26341,N_25169,N_24356);
nand U26342 (N_26342,N_24253,N_24767);
xor U26343 (N_26343,N_24167,N_24851);
nor U26344 (N_26344,N_24703,N_24294);
nor U26345 (N_26345,N_24897,N_24851);
nor U26346 (N_26346,N_24053,N_24245);
nand U26347 (N_26347,N_24421,N_24259);
and U26348 (N_26348,N_24288,N_24893);
or U26349 (N_26349,N_24661,N_25137);
or U26350 (N_26350,N_25133,N_24044);
xnor U26351 (N_26351,N_25123,N_24319);
or U26352 (N_26352,N_24323,N_24942);
xor U26353 (N_26353,N_24786,N_25069);
and U26354 (N_26354,N_25138,N_24858);
and U26355 (N_26355,N_24884,N_24648);
xnor U26356 (N_26356,N_24654,N_24806);
nand U26357 (N_26357,N_25111,N_25105);
and U26358 (N_26358,N_24944,N_24598);
or U26359 (N_26359,N_25186,N_24573);
and U26360 (N_26360,N_24822,N_24990);
xor U26361 (N_26361,N_24470,N_25063);
or U26362 (N_26362,N_24800,N_24162);
nor U26363 (N_26363,N_24815,N_24945);
nand U26364 (N_26364,N_24483,N_24325);
nor U26365 (N_26365,N_24587,N_24951);
xor U26366 (N_26366,N_24079,N_24569);
nand U26367 (N_26367,N_24167,N_24760);
or U26368 (N_26368,N_24333,N_25084);
and U26369 (N_26369,N_24529,N_24425);
nand U26370 (N_26370,N_24564,N_25172);
and U26371 (N_26371,N_25109,N_25193);
or U26372 (N_26372,N_24062,N_25002);
nand U26373 (N_26373,N_24133,N_24187);
or U26374 (N_26374,N_25044,N_24104);
or U26375 (N_26375,N_25038,N_25184);
nand U26376 (N_26376,N_24052,N_25093);
nand U26377 (N_26377,N_24616,N_24994);
xor U26378 (N_26378,N_25187,N_24335);
or U26379 (N_26379,N_24604,N_24283);
nand U26380 (N_26380,N_24729,N_24958);
xnor U26381 (N_26381,N_24459,N_25129);
nand U26382 (N_26382,N_24019,N_25178);
xnor U26383 (N_26383,N_24126,N_24244);
or U26384 (N_26384,N_24368,N_24462);
and U26385 (N_26385,N_24188,N_25181);
and U26386 (N_26386,N_24050,N_24591);
xor U26387 (N_26387,N_25096,N_24255);
or U26388 (N_26388,N_24241,N_24000);
xnor U26389 (N_26389,N_24338,N_24066);
and U26390 (N_26390,N_24067,N_24715);
or U26391 (N_26391,N_24801,N_24093);
xnor U26392 (N_26392,N_24436,N_24279);
and U26393 (N_26393,N_24750,N_24092);
nor U26394 (N_26394,N_24145,N_24091);
xnor U26395 (N_26395,N_25023,N_24099);
and U26396 (N_26396,N_24968,N_25155);
and U26397 (N_26397,N_24199,N_24335);
or U26398 (N_26398,N_24786,N_24356);
nand U26399 (N_26399,N_25011,N_24685);
and U26400 (N_26400,N_25529,N_25656);
xor U26401 (N_26401,N_25997,N_26080);
nor U26402 (N_26402,N_26215,N_25821);
or U26403 (N_26403,N_26246,N_26355);
nand U26404 (N_26404,N_25991,N_26257);
nand U26405 (N_26405,N_25905,N_26082);
and U26406 (N_26406,N_25744,N_26216);
xor U26407 (N_26407,N_25210,N_25893);
or U26408 (N_26408,N_25830,N_25449);
or U26409 (N_26409,N_25450,N_25583);
and U26410 (N_26410,N_25874,N_25316);
xnor U26411 (N_26411,N_25347,N_26230);
nor U26412 (N_26412,N_25851,N_26190);
nor U26413 (N_26413,N_25668,N_25589);
or U26414 (N_26414,N_26389,N_26092);
and U26415 (N_26415,N_26101,N_25435);
nand U26416 (N_26416,N_25405,N_25452);
xnor U26417 (N_26417,N_25585,N_25681);
and U26418 (N_26418,N_26179,N_25341);
or U26419 (N_26419,N_25766,N_26142);
nand U26420 (N_26420,N_25776,N_25535);
nor U26421 (N_26421,N_25528,N_25361);
xor U26422 (N_26422,N_25500,N_26383);
xnor U26423 (N_26423,N_25643,N_25454);
nor U26424 (N_26424,N_25732,N_25843);
and U26425 (N_26425,N_25556,N_25423);
or U26426 (N_26426,N_25741,N_26020);
and U26427 (N_26427,N_25721,N_25385);
xnor U26428 (N_26428,N_26288,N_26342);
nand U26429 (N_26429,N_25456,N_25909);
xor U26430 (N_26430,N_26391,N_25531);
nor U26431 (N_26431,N_26211,N_25526);
and U26432 (N_26432,N_25394,N_25389);
xor U26433 (N_26433,N_26398,N_26220);
and U26434 (N_26434,N_26185,N_25639);
and U26435 (N_26435,N_25919,N_26160);
nor U26436 (N_26436,N_25504,N_25969);
nand U26437 (N_26437,N_25574,N_25952);
xnor U26438 (N_26438,N_26366,N_26236);
xor U26439 (N_26439,N_26223,N_25687);
xnor U26440 (N_26440,N_25773,N_25860);
nor U26441 (N_26441,N_26194,N_25641);
nand U26442 (N_26442,N_25957,N_25671);
xnor U26443 (N_26443,N_26325,N_25376);
xor U26444 (N_26444,N_26197,N_25395);
xor U26445 (N_26445,N_25428,N_25418);
and U26446 (N_26446,N_26386,N_25259);
xnor U26447 (N_26447,N_25939,N_25425);
and U26448 (N_26448,N_26137,N_25820);
or U26449 (N_26449,N_26121,N_26356);
nand U26450 (N_26450,N_26273,N_25416);
and U26451 (N_26451,N_26169,N_25896);
nor U26452 (N_26452,N_25749,N_25448);
and U26453 (N_26453,N_26295,N_25949);
nand U26454 (N_26454,N_25495,N_25914);
nand U26455 (N_26455,N_25768,N_25755);
and U26456 (N_26456,N_25541,N_25483);
or U26457 (N_26457,N_25211,N_25699);
nand U26458 (N_26458,N_25387,N_25831);
nor U26459 (N_26459,N_26077,N_25616);
xor U26460 (N_26460,N_26345,N_25795);
and U26461 (N_26461,N_26265,N_25291);
nand U26462 (N_26462,N_25217,N_26312);
nand U26463 (N_26463,N_25417,N_25520);
nand U26464 (N_26464,N_25993,N_25840);
nor U26465 (N_26465,N_26291,N_25335);
and U26466 (N_26466,N_26118,N_25212);
xnor U26467 (N_26467,N_26244,N_25748);
nor U26468 (N_26468,N_25824,N_25223);
xnor U26469 (N_26469,N_25963,N_26243);
and U26470 (N_26470,N_26192,N_26340);
nor U26471 (N_26471,N_25973,N_25492);
or U26472 (N_26472,N_26298,N_26181);
or U26473 (N_26473,N_25443,N_25578);
xnor U26474 (N_26474,N_25678,N_25360);
nor U26475 (N_26475,N_25393,N_25754);
nand U26476 (N_26476,N_25459,N_26313);
and U26477 (N_26477,N_26394,N_26175);
and U26478 (N_26478,N_25396,N_25612);
or U26479 (N_26479,N_25277,N_25723);
and U26480 (N_26480,N_25779,N_25884);
or U26481 (N_26481,N_25868,N_25793);
and U26482 (N_26482,N_25299,N_26155);
and U26483 (N_26483,N_25968,N_25314);
or U26484 (N_26484,N_25622,N_25995);
or U26485 (N_26485,N_26209,N_25994);
xnor U26486 (N_26486,N_25850,N_25225);
or U26487 (N_26487,N_25849,N_25606);
or U26488 (N_26488,N_26059,N_25265);
or U26489 (N_26489,N_25724,N_25374);
xnor U26490 (N_26490,N_26364,N_25427);
or U26491 (N_26491,N_26350,N_26287);
nor U26492 (N_26492,N_25352,N_25215);
nor U26493 (N_26493,N_25813,N_26128);
and U26494 (N_26494,N_25708,N_26173);
or U26495 (N_26495,N_26286,N_25826);
nor U26496 (N_26496,N_25561,N_26060);
xnor U26497 (N_26497,N_25981,N_26005);
and U26498 (N_26498,N_25653,N_25305);
nor U26499 (N_26499,N_25750,N_25859);
xnor U26500 (N_26500,N_26114,N_26013);
xnor U26501 (N_26501,N_26382,N_25486);
nor U26502 (N_26502,N_26262,N_25301);
xnor U26503 (N_26503,N_26213,N_25260);
or U26504 (N_26504,N_26148,N_25588);
or U26505 (N_26505,N_26285,N_25867);
nand U26506 (N_26506,N_25604,N_26311);
or U26507 (N_26507,N_26376,N_25224);
nor U26508 (N_26508,N_26308,N_25367);
nor U26509 (N_26509,N_25739,N_26097);
or U26510 (N_26510,N_25282,N_25392);
and U26511 (N_26511,N_25864,N_25657);
or U26512 (N_26512,N_25717,N_26307);
nand U26513 (N_26513,N_26384,N_25664);
nand U26514 (N_26514,N_25207,N_25828);
nor U26515 (N_26515,N_25298,N_25818);
and U26516 (N_26516,N_26122,N_25244);
or U26517 (N_26517,N_26078,N_25659);
xor U26518 (N_26518,N_25373,N_25789);
or U26519 (N_26519,N_25325,N_25380);
xor U26520 (N_26520,N_25594,N_25953);
nor U26521 (N_26521,N_25987,N_26015);
nor U26522 (N_26522,N_26163,N_25303);
or U26523 (N_26523,N_26075,N_26214);
or U26524 (N_26524,N_26202,N_25990);
xnor U26525 (N_26525,N_25431,N_25798);
and U26526 (N_26526,N_26027,N_25568);
xnor U26527 (N_26527,N_25227,N_26306);
nor U26528 (N_26528,N_25565,N_25257);
and U26529 (N_26529,N_25557,N_26079);
and U26530 (N_26530,N_25734,N_25623);
or U26531 (N_26531,N_25845,N_26167);
and U26532 (N_26532,N_26309,N_25965);
nor U26533 (N_26533,N_25407,N_25488);
nand U26534 (N_26534,N_26222,N_25652);
or U26535 (N_26535,N_25371,N_25894);
or U26536 (N_26536,N_25327,N_26186);
nor U26537 (N_26537,N_26344,N_25958);
or U26538 (N_26538,N_26260,N_25365);
xor U26539 (N_26539,N_25966,N_25572);
and U26540 (N_26540,N_25937,N_26043);
nand U26541 (N_26541,N_25581,N_25400);
and U26542 (N_26542,N_25890,N_26224);
and U26543 (N_26543,N_26371,N_25285);
xor U26544 (N_26544,N_25209,N_26041);
nor U26545 (N_26545,N_25555,N_25735);
and U26546 (N_26546,N_25985,N_26333);
xor U26547 (N_26547,N_25370,N_26226);
or U26548 (N_26548,N_25662,N_25803);
and U26549 (N_26549,N_25988,N_25899);
and U26550 (N_26550,N_26094,N_25917);
nand U26551 (N_26551,N_25543,N_26237);
nor U26552 (N_26552,N_25892,N_26293);
nor U26553 (N_26553,N_26289,N_26045);
and U26554 (N_26554,N_25745,N_25722);
nor U26555 (N_26555,N_26145,N_26305);
xnor U26556 (N_26556,N_25762,N_26251);
nor U26557 (N_26557,N_25839,N_26357);
nor U26558 (N_26558,N_25916,N_25362);
or U26559 (N_26559,N_26178,N_26234);
and U26560 (N_26560,N_26087,N_25608);
nor U26561 (N_26561,N_25644,N_25240);
nor U26562 (N_26562,N_25466,N_26008);
and U26563 (N_26563,N_26009,N_25689);
and U26564 (N_26564,N_26256,N_25221);
nor U26565 (N_26565,N_25494,N_25967);
nand U26566 (N_26566,N_25458,N_25978);
or U26567 (N_26567,N_25636,N_26314);
xor U26568 (N_26568,N_25465,N_26136);
nand U26569 (N_26569,N_26171,N_25709);
xor U26570 (N_26570,N_25251,N_25710);
or U26571 (N_26571,N_26166,N_25880);
nor U26572 (N_26572,N_25794,N_25551);
and U26573 (N_26573,N_26055,N_25386);
or U26574 (N_26574,N_25312,N_26347);
xnor U26575 (N_26575,N_25942,N_25307);
nand U26576 (N_26576,N_25467,N_26238);
or U26577 (N_26577,N_25955,N_25539);
and U26578 (N_26578,N_26058,N_25442);
nor U26579 (N_26579,N_26107,N_26248);
or U26580 (N_26580,N_25796,N_26219);
nor U26581 (N_26581,N_26116,N_25777);
xnor U26582 (N_26582,N_26396,N_26139);
nand U26583 (N_26583,N_26200,N_26143);
xor U26584 (N_26584,N_25889,N_25271);
nor U26585 (N_26585,N_26051,N_25629);
xor U26586 (N_26586,N_25640,N_25879);
and U26587 (N_26587,N_26172,N_25747);
nand U26588 (N_26588,N_26032,N_25614);
nand U26589 (N_26589,N_25328,N_26000);
nand U26590 (N_26590,N_25476,N_25638);
nor U26591 (N_26591,N_25252,N_26241);
or U26592 (N_26592,N_25261,N_25357);
nor U26593 (N_26593,N_26146,N_26199);
xor U26594 (N_26594,N_25847,N_25489);
and U26595 (N_26595,N_26084,N_25219);
xnor U26596 (N_26596,N_25999,N_25584);
nand U26597 (N_26597,N_26004,N_25502);
nor U26598 (N_26598,N_25478,N_26258);
xor U26599 (N_26599,N_25404,N_25402);
and U26600 (N_26600,N_25497,N_26110);
or U26601 (N_26601,N_25961,N_26158);
and U26602 (N_26602,N_25704,N_26064);
nor U26603 (N_26603,N_26062,N_25635);
nor U26604 (N_26604,N_26050,N_26123);
xnor U26605 (N_26605,N_26296,N_25712);
nand U26606 (N_26606,N_26281,N_25355);
nor U26607 (N_26607,N_26096,N_25401);
or U26608 (N_26608,N_25984,N_25740);
nor U26609 (N_26609,N_26099,N_25288);
nor U26610 (N_26610,N_26011,N_25536);
and U26611 (N_26611,N_26204,N_25731);
nand U26612 (N_26612,N_25615,N_25356);
and U26613 (N_26613,N_26358,N_25586);
nand U26614 (N_26614,N_25715,N_25888);
xor U26615 (N_26615,N_26003,N_25493);
nor U26616 (N_26616,N_25924,N_25617);
nand U26617 (N_26617,N_25992,N_25974);
xor U26618 (N_26618,N_26182,N_26034);
xnor U26619 (N_26619,N_25941,N_26029);
and U26620 (N_26620,N_26030,N_26337);
or U26621 (N_26621,N_26271,N_25487);
nand U26622 (N_26622,N_26381,N_25628);
and U26623 (N_26623,N_25945,N_25881);
xnor U26624 (N_26624,N_25757,N_25563);
and U26625 (N_26625,N_25655,N_26367);
xnor U26626 (N_26626,N_26001,N_26205);
xnor U26627 (N_26627,N_25782,N_25982);
or U26628 (N_26628,N_25245,N_26072);
nand U26629 (N_26629,N_26069,N_26152);
nand U26630 (N_26630,N_25420,N_26090);
xnor U26631 (N_26631,N_26022,N_26250);
xnor U26632 (N_26632,N_26012,N_26073);
or U26633 (N_26633,N_25481,N_25844);
nand U26634 (N_26634,N_25775,N_26089);
nand U26635 (N_26635,N_25948,N_25296);
xor U26636 (N_26636,N_26259,N_25759);
nand U26637 (N_26637,N_26195,N_26377);
nand U26638 (N_26638,N_25691,N_25203);
nor U26639 (N_26639,N_25354,N_26033);
and U26640 (N_26640,N_25885,N_25564);
nor U26641 (N_26641,N_26112,N_25419);
or U26642 (N_26642,N_26188,N_25672);
nor U26643 (N_26643,N_25650,N_25313);
and U26644 (N_26644,N_25625,N_25562);
xnor U26645 (N_26645,N_26266,N_25339);
or U26646 (N_26646,N_25243,N_25742);
nand U26647 (N_26647,N_25771,N_25887);
nand U26648 (N_26648,N_25372,N_25797);
nand U26649 (N_26649,N_25802,N_25979);
and U26650 (N_26650,N_25727,N_25334);
xor U26651 (N_26651,N_25876,N_26363);
nor U26652 (N_26652,N_25455,N_26331);
nand U26653 (N_26653,N_25247,N_25573);
xnor U26654 (N_26654,N_25838,N_26274);
xor U26655 (N_26655,N_25897,N_26379);
or U26656 (N_26656,N_25514,N_26385);
and U26657 (N_26657,N_25451,N_25345);
and U26658 (N_26658,N_25571,N_26362);
nor U26659 (N_26659,N_25854,N_25834);
nor U26660 (N_26660,N_25342,N_25618);
xnor U26661 (N_26661,N_26231,N_25507);
nor U26662 (N_26662,N_25553,N_25554);
xnor U26663 (N_26663,N_25809,N_26267);
xnor U26664 (N_26664,N_25324,N_25829);
xnor U26665 (N_26665,N_25284,N_25413);
and U26666 (N_26666,N_26397,N_25511);
or U26667 (N_26667,N_25343,N_25841);
nand U26668 (N_26668,N_25415,N_26046);
and U26669 (N_26669,N_26300,N_26225);
or U26670 (N_26670,N_25645,N_25311);
or U26671 (N_26671,N_26310,N_25944);
nand U26672 (N_26672,N_25411,N_25632);
nand U26673 (N_26673,N_25522,N_25457);
nand U26674 (N_26674,N_26252,N_25403);
xor U26675 (N_26675,N_25234,N_25501);
nand U26676 (N_26676,N_26091,N_26157);
nand U26677 (N_26677,N_25787,N_25853);
xor U26678 (N_26678,N_25607,N_25577);
and U26679 (N_26679,N_26242,N_25218);
nor U26680 (N_26680,N_25906,N_26024);
and U26681 (N_26681,N_25432,N_25464);
xnor U26682 (N_26682,N_25214,N_25280);
and U26683 (N_26683,N_25231,N_25290);
nand U26684 (N_26684,N_26232,N_25575);
or U26685 (N_26685,N_25682,N_25900);
nor U26686 (N_26686,N_25254,N_25326);
and U26687 (N_26687,N_25769,N_25238);
or U26688 (N_26688,N_26028,N_26361);
or U26689 (N_26689,N_25695,N_25471);
xnor U26690 (N_26690,N_25950,N_25509);
xnor U26691 (N_26691,N_25579,N_25624);
nor U26692 (N_26692,N_26352,N_26221);
or U26693 (N_26693,N_26254,N_25790);
xor U26694 (N_26694,N_25667,N_26125);
nand U26695 (N_26695,N_25286,N_25477);
or U26696 (N_26696,N_25814,N_26002);
nor U26697 (N_26697,N_25409,N_26061);
or U26698 (N_26698,N_25576,N_25752);
xor U26699 (N_26699,N_25513,N_25700);
or U26700 (N_26700,N_25649,N_25346);
nor U26701 (N_26701,N_26294,N_25846);
nand U26702 (N_26702,N_25725,N_26135);
or U26703 (N_26703,N_26218,N_26161);
and U26704 (N_26704,N_25527,N_25698);
or U26705 (N_26705,N_25533,N_26320);
nand U26706 (N_26706,N_25980,N_25783);
or U26707 (N_26707,N_25515,N_26301);
nand U26708 (N_26708,N_26187,N_26323);
and U26709 (N_26709,N_25878,N_25737);
nor U26710 (N_26710,N_25518,N_25460);
nor U26711 (N_26711,N_26113,N_25743);
or U26712 (N_26712,N_26159,N_25570);
and U26713 (N_26713,N_25758,N_25619);
and U26714 (N_26714,N_25304,N_25414);
or U26715 (N_26715,N_25801,N_25300);
xnor U26716 (N_26716,N_25631,N_26303);
nand U26717 (N_26717,N_25626,N_26374);
xor U26718 (N_26718,N_26368,N_26280);
nand U26719 (N_26719,N_25852,N_26006);
or U26720 (N_26720,N_26268,N_26353);
nor U26721 (N_26721,N_25877,N_26229);
xnor U26722 (N_26722,N_26036,N_25947);
and U26723 (N_26723,N_25837,N_26130);
nand U26724 (N_26724,N_25201,N_25253);
or U26725 (N_26725,N_25268,N_26201);
or U26726 (N_26726,N_25318,N_25634);
xnor U26727 (N_26727,N_25600,N_26191);
or U26728 (N_26728,N_25669,N_25901);
xor U26729 (N_26729,N_25907,N_26279);
or U26730 (N_26730,N_25331,N_25598);
and U26731 (N_26731,N_25677,N_25788);
or U26732 (N_26732,N_25491,N_25663);
and U26733 (N_26733,N_25596,N_25283);
and U26734 (N_26734,N_25805,N_25437);
or U26735 (N_26735,N_25666,N_25951);
xor U26736 (N_26736,N_25525,N_25292);
or U26737 (N_26737,N_26047,N_26054);
xnor U26738 (N_26738,N_25825,N_26359);
or U26739 (N_26739,N_26304,N_25774);
xnor U26740 (N_26740,N_25320,N_26212);
and U26741 (N_26741,N_26007,N_25366);
nand U26742 (N_26742,N_26315,N_26253);
and U26743 (N_26743,N_25422,N_25383);
nor U26744 (N_26744,N_26198,N_25397);
xnor U26745 (N_26745,N_25791,N_25381);
nand U26746 (N_26746,N_25751,N_25646);
or U26747 (N_26747,N_25249,N_25675);
or U26748 (N_26748,N_26144,N_26245);
xor U26749 (N_26749,N_26035,N_26162);
nor U26750 (N_26750,N_25351,N_25302);
or U26751 (N_26751,N_25858,N_26247);
nor U26752 (N_26752,N_25654,N_25236);
xor U26753 (N_26753,N_25902,N_25239);
and U26754 (N_26754,N_25591,N_26120);
nand U26755 (N_26755,N_25424,N_25545);
nand U26756 (N_26756,N_25279,N_26138);
or U26757 (N_26757,N_25819,N_26210);
nor U26758 (N_26758,N_25960,N_25815);
nand U26759 (N_26759,N_26275,N_25621);
nor U26760 (N_26760,N_25637,N_25983);
and U26761 (N_26761,N_25333,N_25222);
nor U26762 (N_26762,N_25547,N_25806);
and U26763 (N_26763,N_25627,N_26151);
nand U26764 (N_26764,N_25287,N_25883);
and U26765 (N_26765,N_26105,N_25266);
nor U26766 (N_26766,N_26348,N_25613);
xor U26767 (N_26767,N_25378,N_26102);
or U26768 (N_26768,N_25270,N_25886);
or U26769 (N_26769,N_25469,N_26039);
nand U26770 (N_26770,N_25359,N_26351);
nand U26771 (N_26771,N_26154,N_26193);
nor U26772 (N_26772,N_26129,N_26322);
and U26773 (N_26773,N_25683,N_25857);
nand U26774 (N_26774,N_25546,N_25760);
or U26775 (N_26775,N_25697,N_25692);
or U26776 (N_26776,N_26233,N_25463);
nor U26777 (N_26777,N_26392,N_26184);
nand U26778 (N_26778,N_26086,N_26127);
nand U26779 (N_26779,N_26149,N_25242);
nor U26780 (N_26780,N_26170,N_26206);
or U26781 (N_26781,N_25706,N_25205);
nand U26782 (N_26782,N_25363,N_26263);
or U26783 (N_26783,N_26018,N_25332);
nand U26784 (N_26784,N_26071,N_25926);
nor U26785 (N_26785,N_25676,N_25792);
xnor U26786 (N_26786,N_26264,N_26180);
nand U26787 (N_26787,N_26053,N_25317);
nand U26788 (N_26788,N_25559,N_25808);
nand U26789 (N_26789,N_25696,N_26334);
or U26790 (N_26790,N_25473,N_25693);
and U26791 (N_26791,N_26319,N_25915);
nor U26792 (N_26792,N_26066,N_25611);
nor U26793 (N_26793,N_25707,N_25764);
and U26794 (N_26794,N_25927,N_25329);
xnor U26795 (N_26795,N_25321,N_25264);
nand U26796 (N_26796,N_26276,N_26065);
and U26797 (N_26797,N_26038,N_25661);
xnor U26798 (N_26798,N_25338,N_25785);
and U26799 (N_26799,N_26168,N_26056);
or U26800 (N_26800,N_26228,N_25728);
xnor U26801 (N_26801,N_25865,N_25936);
xor U26802 (N_26802,N_25904,N_26019);
nor U26803 (N_26803,N_25538,N_26150);
nand U26804 (N_26804,N_25817,N_25323);
nor U26805 (N_26805,N_25781,N_25421);
xor U26806 (N_26806,N_25954,N_26057);
nor U26807 (N_26807,N_26302,N_26278);
xnor U26808 (N_26808,N_26131,N_25255);
and U26809 (N_26809,N_25548,N_25694);
nor U26810 (N_26810,N_25964,N_25350);
xor U26811 (N_26811,N_25484,N_26284);
and U26812 (N_26812,N_26100,N_26330);
xor U26813 (N_26813,N_25756,N_25680);
and U26814 (N_26814,N_25800,N_25315);
nand U26815 (N_26815,N_25972,N_25610);
xor U26816 (N_26816,N_26126,N_25462);
nand U26817 (N_26817,N_25256,N_25595);
xor U26818 (N_26818,N_26387,N_25508);
and U26819 (N_26819,N_25412,N_26372);
or U26820 (N_26820,N_25474,N_25701);
or U26821 (N_26821,N_25807,N_25989);
and U26822 (N_26822,N_26140,N_26141);
or U26823 (N_26823,N_25827,N_26378);
or U26824 (N_26824,N_25399,N_26388);
and U26825 (N_26825,N_26085,N_25872);
xor U26826 (N_26826,N_25934,N_25358);
or U26827 (N_26827,N_25241,N_26156);
nor U26828 (N_26828,N_25832,N_25230);
nand U26829 (N_26829,N_25461,N_25716);
nor U26830 (N_26830,N_25761,N_25479);
or U26831 (N_26831,N_25862,N_26134);
nand U26832 (N_26832,N_26365,N_26067);
xnor U26833 (N_26833,N_25620,N_25534);
nor U26834 (N_26834,N_25597,N_25337);
xor U26835 (N_26835,N_26189,N_25517);
nand U26836 (N_26836,N_26349,N_25882);
nand U26837 (N_26837,N_25869,N_25673);
and U26838 (N_26838,N_26346,N_26026);
nor U26839 (N_26839,N_26063,N_25811);
nor U26840 (N_26840,N_25379,N_26176);
and U26841 (N_26841,N_26341,N_26052);
and U26842 (N_26842,N_26360,N_25943);
or U26843 (N_26843,N_26239,N_25833);
and U26844 (N_26844,N_26153,N_26261);
or U26845 (N_26845,N_25935,N_25580);
xor U26846 (N_26846,N_25861,N_25702);
nand U26847 (N_26847,N_26023,N_26321);
or U26848 (N_26848,N_25310,N_25956);
nor U26849 (N_26849,N_25532,N_26017);
and U26850 (N_26850,N_25524,N_25684);
nor U26851 (N_26851,N_25922,N_26070);
xnor U26852 (N_26852,N_25590,N_25660);
and U26853 (N_26853,N_26031,N_26328);
nor U26854 (N_26854,N_25810,N_25946);
and U26855 (N_26855,N_26088,N_26272);
or U26856 (N_26856,N_25705,N_26164);
and U26857 (N_26857,N_25962,N_25587);
and U26858 (N_26858,N_25521,N_25891);
xnor U26859 (N_26859,N_25920,N_26016);
xor U26860 (N_26860,N_25592,N_25267);
or U26861 (N_26861,N_25903,N_26240);
and U26862 (N_26862,N_25938,N_26332);
xnor U26863 (N_26863,N_26021,N_25364);
xnor U26864 (N_26864,N_25933,N_25248);
nand U26865 (N_26865,N_25530,N_25925);
xnor U26866 (N_26866,N_25932,N_25633);
or U26867 (N_26867,N_25281,N_25278);
nand U26868 (N_26868,N_25237,N_25912);
nor U26869 (N_26869,N_25308,N_25599);
and U26870 (N_26870,N_26196,N_25384);
xnor U26871 (N_26871,N_25447,N_25275);
nor U26872 (N_26872,N_25648,N_26025);
and U26873 (N_26873,N_25388,N_26203);
xor U26874 (N_26874,N_25433,N_26044);
nor U26875 (N_26875,N_25510,N_25552);
nand U26876 (N_26876,N_25382,N_25200);
or U26877 (N_26877,N_26336,N_25498);
nand U26878 (N_26878,N_25786,N_25330);
and U26879 (N_26879,N_25601,N_26249);
and U26880 (N_26880,N_25647,N_25746);
and U26881 (N_26881,N_26338,N_26335);
or U26882 (N_26882,N_26297,N_25726);
or U26883 (N_26883,N_25738,N_25229);
nor U26884 (N_26884,N_25665,N_25441);
nor U26885 (N_26885,N_26369,N_25918);
or U26886 (N_26886,N_25765,N_26068);
xor U26887 (N_26887,N_25630,N_25928);
and U26888 (N_26888,N_26399,N_26010);
nand U26889 (N_26889,N_25519,N_26370);
and U26890 (N_26890,N_26040,N_25703);
xnor U26891 (N_26891,N_25674,N_25713);
and U26892 (N_26892,N_25603,N_25921);
nand U26893 (N_26893,N_25569,N_25506);
and U26894 (N_26894,N_25499,N_25246);
xnor U26895 (N_26895,N_25322,N_26174);
or U26896 (N_26896,N_25986,N_25540);
xor U26897 (N_26897,N_25472,N_25799);
xor U26898 (N_26898,N_25439,N_25228);
xor U26899 (N_26899,N_25642,N_25276);
and U26900 (N_26900,N_26208,N_25567);
xor U26901 (N_26901,N_25816,N_25767);
nor U26902 (N_26902,N_25537,N_25480);
and U26903 (N_26903,N_25468,N_25289);
nor U26904 (N_26904,N_25679,N_25866);
and U26905 (N_26905,N_25812,N_26083);
or U26906 (N_26906,N_25959,N_26292);
and U26907 (N_26907,N_25998,N_26014);
xnor U26908 (N_26908,N_25542,N_26317);
or U26909 (N_26909,N_25485,N_25375);
xnor U26910 (N_26910,N_25319,N_25658);
xor U26911 (N_26911,N_26109,N_25670);
xnor U26912 (N_26912,N_25344,N_25688);
or U26913 (N_26913,N_25871,N_26277);
nand U26914 (N_26914,N_25975,N_25368);
nand U26915 (N_26915,N_25309,N_25898);
nand U26916 (N_26916,N_26282,N_25377);
nand U26917 (N_26917,N_26049,N_25855);
xnor U26918 (N_26918,N_26177,N_25895);
xnor U26919 (N_26919,N_25482,N_25685);
nand U26920 (N_26920,N_25202,N_25390);
nor U26921 (N_26921,N_25971,N_25490);
xor U26922 (N_26922,N_25408,N_26119);
nand U26923 (N_26923,N_25908,N_25923);
nor U26924 (N_26924,N_25250,N_25720);
xnor U26925 (N_26925,N_25269,N_25566);
or U26926 (N_26926,N_25516,N_26108);
or U26927 (N_26927,N_25446,N_25274);
nand U26928 (N_26928,N_26390,N_25842);
and U26929 (N_26929,N_25582,N_25729);
nor U26930 (N_26930,N_25505,N_25391);
xor U26931 (N_26931,N_26098,N_25856);
or U26932 (N_26932,N_25306,N_25398);
and U26933 (N_26933,N_26133,N_25445);
nor U26934 (N_26934,N_25208,N_26299);
nand U26935 (N_26935,N_25550,N_26147);
xnor U26936 (N_26936,N_26111,N_25730);
nor U26937 (N_26937,N_25426,N_25910);
nor U26938 (N_26938,N_25733,N_26103);
nor U26939 (N_26939,N_25863,N_25503);
nand U26940 (N_26940,N_25258,N_25353);
xnor U26941 (N_26941,N_25686,N_25213);
nand U26942 (N_26942,N_26207,N_26048);
nor U26943 (N_26943,N_26115,N_25470);
xor U26944 (N_26944,N_25204,N_25602);
or U26945 (N_26945,N_25930,N_25848);
xnor U26946 (N_26946,N_26269,N_26037);
nor U26947 (N_26947,N_25605,N_25349);
nor U26948 (N_26948,N_25206,N_26093);
nor U26949 (N_26949,N_25233,N_25336);
or U26950 (N_26950,N_25294,N_26326);
and U26951 (N_26951,N_26327,N_26235);
xor U26952 (N_26952,N_26343,N_26329);
nor U26953 (N_26953,N_25453,N_26324);
and U26954 (N_26954,N_25835,N_25544);
and U26955 (N_26955,N_26255,N_26318);
xor U26956 (N_26956,N_25875,N_25976);
nor U26957 (N_26957,N_25690,N_26339);
nand U26958 (N_26958,N_25753,N_26290);
nand U26959 (N_26959,N_25444,N_25711);
xor U26960 (N_26960,N_25438,N_25340);
nor U26961 (N_26961,N_26393,N_26165);
xnor U26962 (N_26962,N_25295,N_25931);
xnor U26963 (N_26963,N_26095,N_25558);
and U26964 (N_26964,N_25929,N_25496);
nor U26965 (N_26965,N_25410,N_25778);
nand U26966 (N_26966,N_25823,N_25436);
and U26967 (N_26967,N_26375,N_25429);
nand U26968 (N_26968,N_25836,N_25780);
nand U26969 (N_26969,N_25235,N_25736);
nand U26970 (N_26970,N_25273,N_25772);
nand U26971 (N_26971,N_26354,N_25609);
xnor U26972 (N_26972,N_25714,N_25977);
nand U26973 (N_26973,N_25549,N_25770);
and U26974 (N_26974,N_25406,N_26217);
nand U26975 (N_26975,N_26316,N_25512);
nor U26976 (N_26976,N_25369,N_25348);
xor U26977 (N_26977,N_25996,N_25475);
nor U26978 (N_26978,N_25263,N_25870);
nor U26979 (N_26979,N_26183,N_26380);
xnor U26980 (N_26980,N_25430,N_25719);
xor U26981 (N_26981,N_25822,N_26042);
xor U26982 (N_26982,N_26104,N_25784);
xnor U26983 (N_26983,N_26227,N_26106);
xor U26984 (N_26984,N_25262,N_26117);
xnor U26985 (N_26985,N_25560,N_26132);
and U26986 (N_26986,N_26283,N_25216);
xnor U26987 (N_26987,N_25272,N_26081);
or U26988 (N_26988,N_25913,N_26076);
or U26989 (N_26989,N_25940,N_25523);
xor U26990 (N_26990,N_25226,N_26074);
nand U26991 (N_26991,N_25220,N_25593);
xnor U26992 (N_26992,N_25651,N_26270);
and U26993 (N_26993,N_25970,N_26124);
xor U26994 (N_26994,N_26373,N_25718);
nor U26995 (N_26995,N_25440,N_25911);
and U26996 (N_26996,N_25804,N_26395);
xnor U26997 (N_26997,N_25232,N_25293);
and U26998 (N_26998,N_25763,N_25297);
or U26999 (N_26999,N_25873,N_25434);
and U27000 (N_27000,N_26247,N_26124);
xor U27001 (N_27001,N_25792,N_26158);
and U27002 (N_27002,N_25884,N_25486);
or U27003 (N_27003,N_25917,N_25736);
nand U27004 (N_27004,N_26069,N_25856);
xnor U27005 (N_27005,N_25253,N_25779);
nand U27006 (N_27006,N_25742,N_26122);
and U27007 (N_27007,N_25522,N_25948);
xor U27008 (N_27008,N_25809,N_25237);
nor U27009 (N_27009,N_25991,N_26122);
nor U27010 (N_27010,N_25744,N_26030);
and U27011 (N_27011,N_25827,N_25559);
nand U27012 (N_27012,N_25442,N_25981);
xor U27013 (N_27013,N_25545,N_25936);
nand U27014 (N_27014,N_25229,N_26003);
or U27015 (N_27015,N_25946,N_25410);
or U27016 (N_27016,N_26073,N_25927);
nor U27017 (N_27017,N_25280,N_26083);
or U27018 (N_27018,N_25404,N_25499);
or U27019 (N_27019,N_26136,N_26274);
nor U27020 (N_27020,N_26201,N_26129);
nand U27021 (N_27021,N_25506,N_26166);
or U27022 (N_27022,N_25447,N_26069);
nand U27023 (N_27023,N_25738,N_26075);
nand U27024 (N_27024,N_26333,N_25350);
xnor U27025 (N_27025,N_25841,N_26287);
nor U27026 (N_27026,N_25994,N_26121);
nand U27027 (N_27027,N_25349,N_25583);
or U27028 (N_27028,N_25650,N_25639);
nor U27029 (N_27029,N_26070,N_26071);
or U27030 (N_27030,N_26306,N_26346);
nor U27031 (N_27031,N_26324,N_26068);
nor U27032 (N_27032,N_25586,N_25539);
xnor U27033 (N_27033,N_25814,N_26092);
nor U27034 (N_27034,N_25456,N_25992);
and U27035 (N_27035,N_25770,N_25610);
and U27036 (N_27036,N_26315,N_25288);
nor U27037 (N_27037,N_26349,N_25736);
or U27038 (N_27038,N_25754,N_25721);
xor U27039 (N_27039,N_25554,N_25573);
or U27040 (N_27040,N_25974,N_25710);
nand U27041 (N_27041,N_25226,N_26353);
xnor U27042 (N_27042,N_25783,N_25899);
xnor U27043 (N_27043,N_25367,N_25858);
and U27044 (N_27044,N_26083,N_25468);
and U27045 (N_27045,N_25497,N_25226);
or U27046 (N_27046,N_25263,N_26228);
or U27047 (N_27047,N_25527,N_25289);
nand U27048 (N_27048,N_26161,N_25336);
xnor U27049 (N_27049,N_26078,N_25605);
nor U27050 (N_27050,N_25583,N_25517);
nand U27051 (N_27051,N_25859,N_25960);
nor U27052 (N_27052,N_25680,N_25494);
nor U27053 (N_27053,N_25694,N_25966);
nor U27054 (N_27054,N_25604,N_26350);
and U27055 (N_27055,N_26067,N_25222);
and U27056 (N_27056,N_26081,N_25271);
nand U27057 (N_27057,N_25850,N_25564);
nand U27058 (N_27058,N_25741,N_26220);
nor U27059 (N_27059,N_25330,N_25829);
xnor U27060 (N_27060,N_25471,N_25630);
nand U27061 (N_27061,N_25925,N_25313);
nand U27062 (N_27062,N_25425,N_26023);
xor U27063 (N_27063,N_25274,N_25651);
or U27064 (N_27064,N_26267,N_26076);
nor U27065 (N_27065,N_25873,N_26000);
xor U27066 (N_27066,N_25358,N_26292);
xnor U27067 (N_27067,N_25872,N_25543);
and U27068 (N_27068,N_25976,N_25905);
xnor U27069 (N_27069,N_25536,N_25819);
nand U27070 (N_27070,N_25764,N_25885);
or U27071 (N_27071,N_26303,N_25798);
or U27072 (N_27072,N_25861,N_25672);
nor U27073 (N_27073,N_25598,N_26105);
or U27074 (N_27074,N_26162,N_26215);
nor U27075 (N_27075,N_26011,N_26316);
or U27076 (N_27076,N_25831,N_26195);
and U27077 (N_27077,N_25490,N_26387);
nand U27078 (N_27078,N_26383,N_25578);
nor U27079 (N_27079,N_26252,N_25598);
nand U27080 (N_27080,N_25930,N_25259);
or U27081 (N_27081,N_26185,N_26124);
nand U27082 (N_27082,N_26321,N_25913);
and U27083 (N_27083,N_25634,N_25633);
nand U27084 (N_27084,N_25926,N_25269);
nor U27085 (N_27085,N_25698,N_26004);
or U27086 (N_27086,N_26148,N_25415);
xnor U27087 (N_27087,N_25284,N_25504);
nor U27088 (N_27088,N_25384,N_25841);
or U27089 (N_27089,N_25496,N_26217);
nor U27090 (N_27090,N_26013,N_25391);
and U27091 (N_27091,N_25736,N_26134);
xnor U27092 (N_27092,N_25411,N_26349);
nand U27093 (N_27093,N_25448,N_25453);
and U27094 (N_27094,N_25342,N_26117);
nor U27095 (N_27095,N_25273,N_25604);
nand U27096 (N_27096,N_25454,N_25962);
xnor U27097 (N_27097,N_26333,N_25967);
xor U27098 (N_27098,N_25240,N_25385);
or U27099 (N_27099,N_25948,N_25428);
or U27100 (N_27100,N_25915,N_26264);
nand U27101 (N_27101,N_25943,N_25376);
or U27102 (N_27102,N_25534,N_25536);
or U27103 (N_27103,N_26304,N_26177);
or U27104 (N_27104,N_26123,N_25285);
or U27105 (N_27105,N_25474,N_25727);
and U27106 (N_27106,N_25605,N_25401);
nand U27107 (N_27107,N_25613,N_25883);
nand U27108 (N_27108,N_25671,N_25806);
or U27109 (N_27109,N_25986,N_25701);
nand U27110 (N_27110,N_25954,N_25780);
and U27111 (N_27111,N_25442,N_25731);
nand U27112 (N_27112,N_26247,N_25696);
or U27113 (N_27113,N_25488,N_25805);
nor U27114 (N_27114,N_25640,N_25755);
nand U27115 (N_27115,N_25511,N_25969);
or U27116 (N_27116,N_25564,N_26117);
and U27117 (N_27117,N_25643,N_25372);
nand U27118 (N_27118,N_25802,N_26093);
nand U27119 (N_27119,N_26100,N_25517);
xnor U27120 (N_27120,N_26273,N_25308);
and U27121 (N_27121,N_25967,N_25770);
nor U27122 (N_27122,N_25311,N_26044);
nor U27123 (N_27123,N_25531,N_25478);
nor U27124 (N_27124,N_26124,N_25915);
xnor U27125 (N_27125,N_25361,N_26004);
nand U27126 (N_27126,N_25281,N_25994);
nor U27127 (N_27127,N_25264,N_26347);
and U27128 (N_27128,N_26010,N_26364);
nand U27129 (N_27129,N_26358,N_25840);
xnor U27130 (N_27130,N_26247,N_25953);
nand U27131 (N_27131,N_25495,N_25295);
or U27132 (N_27132,N_26085,N_25748);
nand U27133 (N_27133,N_26278,N_25570);
nor U27134 (N_27134,N_25514,N_26277);
nor U27135 (N_27135,N_26031,N_26134);
or U27136 (N_27136,N_25950,N_25213);
xor U27137 (N_27137,N_26091,N_26329);
xor U27138 (N_27138,N_26202,N_26312);
or U27139 (N_27139,N_25689,N_25292);
or U27140 (N_27140,N_25811,N_25250);
and U27141 (N_27141,N_26089,N_25700);
xor U27142 (N_27142,N_26184,N_25379);
nand U27143 (N_27143,N_25847,N_25836);
or U27144 (N_27144,N_25535,N_25861);
xnor U27145 (N_27145,N_26335,N_25632);
xnor U27146 (N_27146,N_26021,N_25931);
and U27147 (N_27147,N_25987,N_25507);
xnor U27148 (N_27148,N_25334,N_25318);
xnor U27149 (N_27149,N_25692,N_25715);
xnor U27150 (N_27150,N_25780,N_26365);
xor U27151 (N_27151,N_26360,N_25465);
nor U27152 (N_27152,N_25278,N_26395);
nand U27153 (N_27153,N_25572,N_26258);
or U27154 (N_27154,N_25388,N_25328);
nor U27155 (N_27155,N_26077,N_26275);
xor U27156 (N_27156,N_25709,N_25230);
nand U27157 (N_27157,N_25860,N_25909);
and U27158 (N_27158,N_25554,N_25597);
or U27159 (N_27159,N_25740,N_25225);
nand U27160 (N_27160,N_26313,N_25523);
nand U27161 (N_27161,N_25450,N_25548);
or U27162 (N_27162,N_26162,N_25530);
xnor U27163 (N_27163,N_25904,N_25721);
or U27164 (N_27164,N_26018,N_25960);
or U27165 (N_27165,N_25312,N_26357);
xor U27166 (N_27166,N_25836,N_26251);
and U27167 (N_27167,N_25441,N_26028);
xnor U27168 (N_27168,N_26171,N_26190);
and U27169 (N_27169,N_26287,N_26244);
or U27170 (N_27170,N_26089,N_25320);
and U27171 (N_27171,N_26115,N_25871);
nand U27172 (N_27172,N_26219,N_25891);
nor U27173 (N_27173,N_26091,N_26018);
or U27174 (N_27174,N_26209,N_25576);
nand U27175 (N_27175,N_25731,N_25857);
nand U27176 (N_27176,N_25566,N_26135);
or U27177 (N_27177,N_26050,N_26164);
or U27178 (N_27178,N_25340,N_25625);
xnor U27179 (N_27179,N_25367,N_26322);
nor U27180 (N_27180,N_25554,N_25634);
and U27181 (N_27181,N_25861,N_25569);
nand U27182 (N_27182,N_25260,N_25308);
and U27183 (N_27183,N_25764,N_25719);
or U27184 (N_27184,N_25956,N_25217);
and U27185 (N_27185,N_26175,N_26022);
or U27186 (N_27186,N_26126,N_26076);
nor U27187 (N_27187,N_25797,N_25993);
xor U27188 (N_27188,N_25511,N_25592);
and U27189 (N_27189,N_25564,N_25997);
or U27190 (N_27190,N_25682,N_25754);
xnor U27191 (N_27191,N_26213,N_25620);
xor U27192 (N_27192,N_26394,N_25784);
or U27193 (N_27193,N_25924,N_25791);
and U27194 (N_27194,N_26197,N_25891);
nor U27195 (N_27195,N_25643,N_25452);
or U27196 (N_27196,N_25230,N_26088);
xnor U27197 (N_27197,N_25666,N_26231);
or U27198 (N_27198,N_25589,N_25648);
and U27199 (N_27199,N_25584,N_25818);
or U27200 (N_27200,N_25877,N_25613);
xor U27201 (N_27201,N_26228,N_26120);
or U27202 (N_27202,N_25550,N_25275);
or U27203 (N_27203,N_26268,N_26107);
nand U27204 (N_27204,N_25773,N_25346);
xnor U27205 (N_27205,N_25956,N_25201);
nor U27206 (N_27206,N_26367,N_25711);
nor U27207 (N_27207,N_26131,N_25346);
and U27208 (N_27208,N_25511,N_25679);
or U27209 (N_27209,N_25793,N_25780);
nor U27210 (N_27210,N_26267,N_25632);
and U27211 (N_27211,N_25935,N_25819);
nor U27212 (N_27212,N_25274,N_25937);
and U27213 (N_27213,N_25791,N_25377);
and U27214 (N_27214,N_25595,N_25923);
xnor U27215 (N_27215,N_25822,N_25642);
xor U27216 (N_27216,N_25410,N_25466);
or U27217 (N_27217,N_25826,N_25930);
and U27218 (N_27218,N_26233,N_26188);
or U27219 (N_27219,N_26328,N_25772);
nor U27220 (N_27220,N_25748,N_25890);
and U27221 (N_27221,N_26366,N_25412);
nor U27222 (N_27222,N_25794,N_25923);
nor U27223 (N_27223,N_26350,N_25546);
nor U27224 (N_27224,N_25973,N_26132);
or U27225 (N_27225,N_25243,N_26279);
and U27226 (N_27226,N_25530,N_25535);
nand U27227 (N_27227,N_25920,N_26356);
or U27228 (N_27228,N_26140,N_26094);
or U27229 (N_27229,N_25537,N_26319);
or U27230 (N_27230,N_26046,N_25245);
xnor U27231 (N_27231,N_25790,N_25388);
nand U27232 (N_27232,N_25840,N_26322);
or U27233 (N_27233,N_25929,N_25913);
nand U27234 (N_27234,N_26097,N_25549);
nor U27235 (N_27235,N_26192,N_26194);
nor U27236 (N_27236,N_26053,N_26358);
and U27237 (N_27237,N_25314,N_26037);
nand U27238 (N_27238,N_26075,N_26159);
nand U27239 (N_27239,N_26133,N_25959);
xor U27240 (N_27240,N_25600,N_25462);
nand U27241 (N_27241,N_25225,N_25476);
or U27242 (N_27242,N_25334,N_26249);
xor U27243 (N_27243,N_25303,N_25501);
nor U27244 (N_27244,N_25864,N_25326);
and U27245 (N_27245,N_25753,N_25969);
xnor U27246 (N_27246,N_25296,N_26108);
nor U27247 (N_27247,N_26003,N_25573);
nand U27248 (N_27248,N_25782,N_26240);
and U27249 (N_27249,N_26347,N_26292);
nor U27250 (N_27250,N_25751,N_25575);
nor U27251 (N_27251,N_25282,N_26297);
xor U27252 (N_27252,N_25904,N_26295);
xor U27253 (N_27253,N_26262,N_26003);
and U27254 (N_27254,N_25261,N_25228);
and U27255 (N_27255,N_25226,N_25326);
or U27256 (N_27256,N_25924,N_26245);
nand U27257 (N_27257,N_26020,N_25544);
xor U27258 (N_27258,N_25441,N_26190);
and U27259 (N_27259,N_26303,N_25930);
or U27260 (N_27260,N_26058,N_25786);
and U27261 (N_27261,N_25384,N_26366);
or U27262 (N_27262,N_25518,N_25502);
and U27263 (N_27263,N_25575,N_26005);
and U27264 (N_27264,N_25490,N_26147);
nor U27265 (N_27265,N_26128,N_26197);
nand U27266 (N_27266,N_25896,N_25417);
nand U27267 (N_27267,N_26272,N_25640);
nand U27268 (N_27268,N_26266,N_25411);
xnor U27269 (N_27269,N_25903,N_25823);
nor U27270 (N_27270,N_25516,N_26192);
xor U27271 (N_27271,N_25881,N_25693);
nand U27272 (N_27272,N_25594,N_25691);
nand U27273 (N_27273,N_25879,N_26249);
xor U27274 (N_27274,N_25386,N_25383);
and U27275 (N_27275,N_25843,N_25587);
and U27276 (N_27276,N_25329,N_26195);
nand U27277 (N_27277,N_25989,N_25200);
or U27278 (N_27278,N_26213,N_26208);
nor U27279 (N_27279,N_25296,N_25289);
nor U27280 (N_27280,N_25325,N_25577);
nand U27281 (N_27281,N_25398,N_25485);
or U27282 (N_27282,N_26367,N_26238);
and U27283 (N_27283,N_26194,N_25233);
and U27284 (N_27284,N_25653,N_26004);
nand U27285 (N_27285,N_26062,N_25728);
nand U27286 (N_27286,N_26302,N_26146);
nand U27287 (N_27287,N_25631,N_25228);
nor U27288 (N_27288,N_26015,N_26146);
xnor U27289 (N_27289,N_26356,N_25288);
nand U27290 (N_27290,N_25795,N_25242);
and U27291 (N_27291,N_25648,N_25564);
and U27292 (N_27292,N_26090,N_26086);
nand U27293 (N_27293,N_25973,N_25257);
nand U27294 (N_27294,N_25764,N_25808);
nor U27295 (N_27295,N_26216,N_25729);
nor U27296 (N_27296,N_25943,N_25851);
nand U27297 (N_27297,N_26034,N_26246);
and U27298 (N_27298,N_25324,N_25407);
or U27299 (N_27299,N_25923,N_25208);
nand U27300 (N_27300,N_26021,N_26108);
or U27301 (N_27301,N_26046,N_25724);
nand U27302 (N_27302,N_26350,N_25247);
nand U27303 (N_27303,N_26363,N_25502);
nor U27304 (N_27304,N_26313,N_25610);
nor U27305 (N_27305,N_25906,N_26114);
and U27306 (N_27306,N_25237,N_26315);
xnor U27307 (N_27307,N_25711,N_26219);
nor U27308 (N_27308,N_26188,N_26054);
xor U27309 (N_27309,N_25208,N_26328);
nor U27310 (N_27310,N_25689,N_26137);
nor U27311 (N_27311,N_25508,N_25873);
nor U27312 (N_27312,N_26145,N_26155);
and U27313 (N_27313,N_26038,N_26350);
nor U27314 (N_27314,N_25557,N_26021);
nand U27315 (N_27315,N_26181,N_25927);
or U27316 (N_27316,N_25584,N_25350);
nor U27317 (N_27317,N_25737,N_25267);
nand U27318 (N_27318,N_25416,N_25769);
or U27319 (N_27319,N_25694,N_25503);
nor U27320 (N_27320,N_26114,N_26397);
and U27321 (N_27321,N_25803,N_25308);
nand U27322 (N_27322,N_25595,N_25873);
xor U27323 (N_27323,N_26087,N_26066);
xnor U27324 (N_27324,N_25481,N_26213);
xnor U27325 (N_27325,N_25702,N_25812);
nand U27326 (N_27326,N_26352,N_26116);
and U27327 (N_27327,N_26310,N_26308);
xnor U27328 (N_27328,N_25631,N_26329);
xnor U27329 (N_27329,N_25708,N_25713);
nor U27330 (N_27330,N_26280,N_25995);
or U27331 (N_27331,N_25621,N_26287);
nor U27332 (N_27332,N_25612,N_26080);
and U27333 (N_27333,N_25788,N_25296);
and U27334 (N_27334,N_26297,N_26115);
nor U27335 (N_27335,N_25627,N_25430);
and U27336 (N_27336,N_25476,N_25775);
or U27337 (N_27337,N_25490,N_25704);
or U27338 (N_27338,N_26396,N_26266);
nand U27339 (N_27339,N_25389,N_25444);
or U27340 (N_27340,N_25220,N_25250);
nand U27341 (N_27341,N_26084,N_25484);
nor U27342 (N_27342,N_26215,N_26271);
nand U27343 (N_27343,N_25679,N_26231);
nor U27344 (N_27344,N_25567,N_25638);
or U27345 (N_27345,N_25419,N_25462);
nor U27346 (N_27346,N_25774,N_25796);
nand U27347 (N_27347,N_26029,N_25615);
or U27348 (N_27348,N_26133,N_25563);
and U27349 (N_27349,N_26220,N_25872);
xor U27350 (N_27350,N_25945,N_26269);
nand U27351 (N_27351,N_25729,N_25602);
or U27352 (N_27352,N_25802,N_25485);
nor U27353 (N_27353,N_25708,N_26079);
xor U27354 (N_27354,N_25952,N_25210);
nand U27355 (N_27355,N_25294,N_25637);
and U27356 (N_27356,N_26120,N_25220);
and U27357 (N_27357,N_25328,N_25914);
xnor U27358 (N_27358,N_26280,N_26379);
and U27359 (N_27359,N_26228,N_25750);
xor U27360 (N_27360,N_25243,N_25347);
and U27361 (N_27361,N_25397,N_26303);
nor U27362 (N_27362,N_25281,N_25678);
and U27363 (N_27363,N_25786,N_25316);
and U27364 (N_27364,N_25883,N_26023);
and U27365 (N_27365,N_26371,N_25260);
nor U27366 (N_27366,N_26352,N_25244);
xnor U27367 (N_27367,N_25282,N_26033);
nand U27368 (N_27368,N_25985,N_25742);
or U27369 (N_27369,N_25691,N_25491);
nand U27370 (N_27370,N_26374,N_25792);
nand U27371 (N_27371,N_25275,N_25584);
xnor U27372 (N_27372,N_26279,N_25671);
xor U27373 (N_27373,N_26021,N_25727);
or U27374 (N_27374,N_25536,N_26300);
xnor U27375 (N_27375,N_25375,N_25250);
and U27376 (N_27376,N_25496,N_25574);
and U27377 (N_27377,N_25794,N_25683);
and U27378 (N_27378,N_25448,N_25295);
nand U27379 (N_27379,N_26106,N_26326);
nand U27380 (N_27380,N_25814,N_25689);
and U27381 (N_27381,N_26108,N_25529);
and U27382 (N_27382,N_26315,N_26125);
xnor U27383 (N_27383,N_26265,N_25515);
xnor U27384 (N_27384,N_25602,N_25521);
and U27385 (N_27385,N_26369,N_25602);
xnor U27386 (N_27386,N_25817,N_26347);
or U27387 (N_27387,N_25466,N_25882);
nand U27388 (N_27388,N_25735,N_26225);
nand U27389 (N_27389,N_26085,N_25809);
and U27390 (N_27390,N_25888,N_26197);
xor U27391 (N_27391,N_26063,N_25297);
and U27392 (N_27392,N_26198,N_26324);
xor U27393 (N_27393,N_25811,N_25679);
or U27394 (N_27394,N_26052,N_25766);
or U27395 (N_27395,N_26327,N_25991);
and U27396 (N_27396,N_25351,N_25750);
nor U27397 (N_27397,N_25270,N_25818);
and U27398 (N_27398,N_25251,N_25594);
xor U27399 (N_27399,N_25362,N_26210);
nor U27400 (N_27400,N_26038,N_26193);
nor U27401 (N_27401,N_25770,N_26036);
xor U27402 (N_27402,N_26266,N_25291);
and U27403 (N_27403,N_26054,N_26162);
and U27404 (N_27404,N_25579,N_25799);
and U27405 (N_27405,N_25396,N_25843);
or U27406 (N_27406,N_25694,N_26329);
xor U27407 (N_27407,N_25716,N_26375);
xor U27408 (N_27408,N_25502,N_25530);
nor U27409 (N_27409,N_26000,N_25677);
and U27410 (N_27410,N_26269,N_25890);
nand U27411 (N_27411,N_25200,N_25246);
nand U27412 (N_27412,N_25833,N_25332);
and U27413 (N_27413,N_25450,N_26011);
or U27414 (N_27414,N_25479,N_25685);
nor U27415 (N_27415,N_26230,N_25825);
nand U27416 (N_27416,N_26124,N_25586);
and U27417 (N_27417,N_25345,N_25560);
xor U27418 (N_27418,N_25746,N_26231);
nor U27419 (N_27419,N_25996,N_25312);
nand U27420 (N_27420,N_26340,N_26136);
nor U27421 (N_27421,N_25268,N_25975);
or U27422 (N_27422,N_25289,N_25449);
xnor U27423 (N_27423,N_25348,N_25995);
nand U27424 (N_27424,N_25885,N_25451);
xor U27425 (N_27425,N_25350,N_26374);
nand U27426 (N_27426,N_25284,N_26144);
nand U27427 (N_27427,N_25456,N_25214);
or U27428 (N_27428,N_25573,N_25729);
and U27429 (N_27429,N_25855,N_25377);
and U27430 (N_27430,N_26131,N_26044);
and U27431 (N_27431,N_26318,N_26045);
nor U27432 (N_27432,N_26227,N_26300);
nand U27433 (N_27433,N_25454,N_26092);
nand U27434 (N_27434,N_25938,N_25895);
nor U27435 (N_27435,N_25373,N_25277);
or U27436 (N_27436,N_26158,N_26230);
nand U27437 (N_27437,N_26365,N_25717);
and U27438 (N_27438,N_25446,N_25911);
and U27439 (N_27439,N_25886,N_25285);
nand U27440 (N_27440,N_25578,N_25625);
and U27441 (N_27441,N_25466,N_26349);
nor U27442 (N_27442,N_26080,N_25254);
or U27443 (N_27443,N_25986,N_25267);
xnor U27444 (N_27444,N_25840,N_26386);
xor U27445 (N_27445,N_26367,N_26320);
or U27446 (N_27446,N_25957,N_26127);
xor U27447 (N_27447,N_25426,N_26368);
nand U27448 (N_27448,N_26071,N_26389);
nor U27449 (N_27449,N_25563,N_25281);
or U27450 (N_27450,N_25823,N_25557);
xnor U27451 (N_27451,N_25699,N_26261);
xnor U27452 (N_27452,N_26197,N_25956);
nor U27453 (N_27453,N_25966,N_25646);
or U27454 (N_27454,N_25438,N_25679);
and U27455 (N_27455,N_26117,N_25608);
nor U27456 (N_27456,N_25572,N_26220);
nand U27457 (N_27457,N_25336,N_25472);
xnor U27458 (N_27458,N_26282,N_25617);
xnor U27459 (N_27459,N_25379,N_25646);
nand U27460 (N_27460,N_25466,N_25656);
nand U27461 (N_27461,N_25932,N_25704);
and U27462 (N_27462,N_25322,N_25641);
nand U27463 (N_27463,N_25516,N_25226);
nand U27464 (N_27464,N_25982,N_25428);
or U27465 (N_27465,N_25869,N_26381);
nand U27466 (N_27466,N_26026,N_25759);
nand U27467 (N_27467,N_25314,N_25542);
or U27468 (N_27468,N_25768,N_25483);
nor U27469 (N_27469,N_26045,N_26007);
and U27470 (N_27470,N_26095,N_25447);
xnor U27471 (N_27471,N_25917,N_26100);
xor U27472 (N_27472,N_25741,N_25381);
and U27473 (N_27473,N_25934,N_26008);
nor U27474 (N_27474,N_26374,N_25397);
nor U27475 (N_27475,N_25999,N_25956);
xor U27476 (N_27476,N_25836,N_26258);
and U27477 (N_27477,N_25703,N_26081);
or U27478 (N_27478,N_25659,N_26200);
or U27479 (N_27479,N_25746,N_26024);
xnor U27480 (N_27480,N_25834,N_26290);
and U27481 (N_27481,N_26317,N_25215);
nor U27482 (N_27482,N_25977,N_25282);
or U27483 (N_27483,N_25389,N_25858);
nor U27484 (N_27484,N_25445,N_25935);
and U27485 (N_27485,N_25539,N_25689);
nand U27486 (N_27486,N_25427,N_25488);
xor U27487 (N_27487,N_25294,N_26306);
nor U27488 (N_27488,N_25478,N_25947);
and U27489 (N_27489,N_25209,N_25671);
xor U27490 (N_27490,N_25857,N_25781);
or U27491 (N_27491,N_25984,N_26346);
nand U27492 (N_27492,N_25448,N_26294);
nor U27493 (N_27493,N_26187,N_26217);
nand U27494 (N_27494,N_25647,N_26321);
nand U27495 (N_27495,N_25741,N_26375);
nor U27496 (N_27496,N_25625,N_26024);
xor U27497 (N_27497,N_25916,N_26357);
nor U27498 (N_27498,N_25803,N_25419);
nand U27499 (N_27499,N_25387,N_26194);
and U27500 (N_27500,N_25547,N_25607);
xor U27501 (N_27501,N_25953,N_25504);
and U27502 (N_27502,N_25233,N_25933);
or U27503 (N_27503,N_26132,N_25466);
xnor U27504 (N_27504,N_25604,N_25539);
or U27505 (N_27505,N_25928,N_25263);
and U27506 (N_27506,N_26344,N_25308);
nor U27507 (N_27507,N_26244,N_26340);
nor U27508 (N_27508,N_26164,N_25389);
or U27509 (N_27509,N_25377,N_26293);
xor U27510 (N_27510,N_26142,N_25956);
or U27511 (N_27511,N_26379,N_25377);
or U27512 (N_27512,N_26265,N_26050);
nand U27513 (N_27513,N_26193,N_25272);
nand U27514 (N_27514,N_25497,N_25920);
xnor U27515 (N_27515,N_25781,N_26329);
nand U27516 (N_27516,N_25858,N_25211);
nand U27517 (N_27517,N_25393,N_25839);
nor U27518 (N_27518,N_25925,N_26171);
nand U27519 (N_27519,N_25859,N_25525);
and U27520 (N_27520,N_26206,N_26394);
xnor U27521 (N_27521,N_26048,N_25419);
xnor U27522 (N_27522,N_25360,N_26290);
nor U27523 (N_27523,N_26108,N_25418);
and U27524 (N_27524,N_26310,N_25713);
and U27525 (N_27525,N_25549,N_25448);
nand U27526 (N_27526,N_26049,N_25536);
nand U27527 (N_27527,N_25208,N_26225);
nor U27528 (N_27528,N_26243,N_25879);
or U27529 (N_27529,N_26153,N_26248);
nand U27530 (N_27530,N_25566,N_26246);
and U27531 (N_27531,N_25661,N_25726);
nor U27532 (N_27532,N_25491,N_25334);
and U27533 (N_27533,N_25705,N_25311);
or U27534 (N_27534,N_26256,N_25937);
nor U27535 (N_27535,N_25592,N_25814);
or U27536 (N_27536,N_25480,N_25364);
xnor U27537 (N_27537,N_25598,N_26187);
nor U27538 (N_27538,N_26357,N_25690);
xor U27539 (N_27539,N_25688,N_25858);
or U27540 (N_27540,N_26259,N_26084);
xor U27541 (N_27541,N_26009,N_25940);
xor U27542 (N_27542,N_25687,N_25645);
nand U27543 (N_27543,N_26065,N_25755);
nand U27544 (N_27544,N_26262,N_25210);
xnor U27545 (N_27545,N_25362,N_25636);
xor U27546 (N_27546,N_25208,N_26273);
nor U27547 (N_27547,N_26249,N_25611);
and U27548 (N_27548,N_25833,N_25411);
xnor U27549 (N_27549,N_25852,N_25222);
or U27550 (N_27550,N_25617,N_26118);
and U27551 (N_27551,N_25610,N_26341);
nand U27552 (N_27552,N_25354,N_26150);
and U27553 (N_27553,N_25961,N_25643);
nand U27554 (N_27554,N_26171,N_25400);
xor U27555 (N_27555,N_25640,N_25464);
nand U27556 (N_27556,N_25283,N_25464);
and U27557 (N_27557,N_25607,N_25213);
nor U27558 (N_27558,N_26058,N_26372);
xnor U27559 (N_27559,N_25969,N_26308);
nor U27560 (N_27560,N_25222,N_25392);
nor U27561 (N_27561,N_25758,N_25802);
nor U27562 (N_27562,N_25381,N_26034);
and U27563 (N_27563,N_25885,N_25822);
nand U27564 (N_27564,N_26306,N_25841);
nor U27565 (N_27565,N_25475,N_25959);
and U27566 (N_27566,N_25647,N_25319);
and U27567 (N_27567,N_25526,N_25988);
nand U27568 (N_27568,N_26380,N_25453);
xor U27569 (N_27569,N_26017,N_25735);
or U27570 (N_27570,N_25296,N_26011);
nor U27571 (N_27571,N_25501,N_26176);
and U27572 (N_27572,N_25491,N_26297);
xor U27573 (N_27573,N_25526,N_26201);
and U27574 (N_27574,N_25731,N_25335);
xnor U27575 (N_27575,N_25794,N_25906);
xnor U27576 (N_27576,N_25557,N_25479);
xnor U27577 (N_27577,N_26235,N_25422);
nand U27578 (N_27578,N_25724,N_25499);
xor U27579 (N_27579,N_25265,N_25377);
and U27580 (N_27580,N_25814,N_25507);
nand U27581 (N_27581,N_26029,N_25729);
and U27582 (N_27582,N_26326,N_26041);
xnor U27583 (N_27583,N_26226,N_25592);
and U27584 (N_27584,N_25395,N_25752);
xnor U27585 (N_27585,N_25721,N_25563);
or U27586 (N_27586,N_26210,N_25208);
nor U27587 (N_27587,N_25985,N_26153);
nand U27588 (N_27588,N_25803,N_25804);
and U27589 (N_27589,N_25890,N_25953);
or U27590 (N_27590,N_25919,N_26008);
xnor U27591 (N_27591,N_25474,N_26108);
nor U27592 (N_27592,N_25974,N_26281);
and U27593 (N_27593,N_25862,N_25928);
or U27594 (N_27594,N_25586,N_25756);
nand U27595 (N_27595,N_25679,N_25695);
or U27596 (N_27596,N_26373,N_25264);
or U27597 (N_27597,N_25962,N_26044);
nand U27598 (N_27598,N_26224,N_25899);
and U27599 (N_27599,N_25652,N_26084);
or U27600 (N_27600,N_26557,N_26595);
nor U27601 (N_27601,N_27005,N_27043);
xnor U27602 (N_27602,N_27328,N_27022);
nor U27603 (N_27603,N_26427,N_27322);
xor U27604 (N_27604,N_27369,N_26946);
or U27605 (N_27605,N_26588,N_26492);
and U27606 (N_27606,N_27024,N_26716);
xor U27607 (N_27607,N_27231,N_27408);
and U27608 (N_27608,N_27078,N_26610);
nand U27609 (N_27609,N_27352,N_26520);
nor U27610 (N_27610,N_27407,N_26835);
and U27611 (N_27611,N_26795,N_26552);
nand U27612 (N_27612,N_26685,N_27382);
xnor U27613 (N_27613,N_27004,N_26504);
xor U27614 (N_27614,N_27112,N_26819);
nand U27615 (N_27615,N_26505,N_26511);
and U27616 (N_27616,N_26777,N_27470);
nand U27617 (N_27617,N_26961,N_26831);
or U27618 (N_27618,N_27472,N_27528);
nand U27619 (N_27619,N_26626,N_26986);
xor U27620 (N_27620,N_27038,N_26900);
nand U27621 (N_27621,N_26995,N_27154);
xor U27622 (N_27622,N_27228,N_26927);
xnor U27623 (N_27623,N_27145,N_27313);
nand U27624 (N_27624,N_27340,N_27456);
xor U27625 (N_27625,N_26928,N_26600);
and U27626 (N_27626,N_27416,N_27594);
nand U27627 (N_27627,N_27214,N_26516);
nand U27628 (N_27628,N_26471,N_27324);
nor U27629 (N_27629,N_26637,N_26838);
or U27630 (N_27630,N_27204,N_27089);
nor U27631 (N_27631,N_27372,N_27277);
xnor U27632 (N_27632,N_27373,N_26810);
nor U27633 (N_27633,N_27557,N_27297);
xnor U27634 (N_27634,N_26655,N_26765);
nor U27635 (N_27635,N_26878,N_26875);
xnor U27636 (N_27636,N_26815,N_27220);
and U27637 (N_27637,N_27240,N_27578);
nand U27638 (N_27638,N_26867,N_27377);
and U27639 (N_27639,N_26828,N_27044);
nor U27640 (N_27640,N_27325,N_27545);
xor U27641 (N_27641,N_26524,N_27099);
nor U27642 (N_27642,N_26638,N_27055);
and U27643 (N_27643,N_27344,N_26873);
nor U27644 (N_27644,N_26969,N_27567);
or U27645 (N_27645,N_26847,N_26434);
or U27646 (N_27646,N_26973,N_26899);
and U27647 (N_27647,N_27579,N_27315);
or U27648 (N_27648,N_26688,N_27410);
nand U27649 (N_27649,N_27386,N_27589);
or U27650 (N_27650,N_27559,N_26984);
nor U27651 (N_27651,N_26431,N_26517);
nand U27652 (N_27652,N_26958,N_27433);
nor U27653 (N_27653,N_26842,N_26786);
and U27654 (N_27654,N_26743,N_26449);
nor U27655 (N_27655,N_27029,N_26499);
nor U27656 (N_27656,N_27124,N_26792);
xor U27657 (N_27657,N_27212,N_26910);
or U27658 (N_27658,N_27039,N_26893);
xor U27659 (N_27659,N_27343,N_26465);
or U27660 (N_27660,N_26660,N_26843);
or U27661 (N_27661,N_26923,N_27292);
nand U27662 (N_27662,N_26543,N_26953);
nand U27663 (N_27663,N_26938,N_26460);
or U27664 (N_27664,N_26715,N_26426);
nand U27665 (N_27665,N_26955,N_26904);
and U27666 (N_27666,N_26436,N_27356);
nand U27667 (N_27667,N_26531,N_26745);
nor U27668 (N_27668,N_27013,N_26635);
xnor U27669 (N_27669,N_27139,N_26523);
nor U27670 (N_27670,N_27573,N_26456);
xnor U27671 (N_27671,N_26494,N_27192);
nand U27672 (N_27672,N_26420,N_27244);
and U27673 (N_27673,N_26732,N_27429);
and U27674 (N_27674,N_26664,N_27002);
nand U27675 (N_27675,N_27025,N_27412);
or U27676 (N_27676,N_26858,N_27235);
or U27677 (N_27677,N_27580,N_27184);
nand U27678 (N_27678,N_27418,N_26539);
nor U27679 (N_27679,N_26982,N_26445);
nor U27680 (N_27680,N_27193,N_27367);
xor U27681 (N_27681,N_27040,N_26981);
nor U27682 (N_27682,N_27009,N_26924);
or U27683 (N_27683,N_27018,N_26856);
nand U27684 (N_27684,N_26992,N_26763);
or U27685 (N_27685,N_26750,N_26797);
or U27686 (N_27686,N_26443,N_27522);
nand U27687 (N_27687,N_26562,N_27434);
or U27688 (N_27688,N_26439,N_26423);
or U27689 (N_27689,N_27052,N_26599);
or U27690 (N_27690,N_27444,N_26811);
and U27691 (N_27691,N_27469,N_27098);
nor U27692 (N_27692,N_27525,N_27458);
nand U27693 (N_27693,N_26921,N_26729);
nor U27694 (N_27694,N_26941,N_26617);
xnor U27695 (N_27695,N_26816,N_27249);
nor U27696 (N_27696,N_27065,N_27069);
xnor U27697 (N_27697,N_27405,N_27076);
nand U27698 (N_27698,N_26653,N_27530);
nor U27699 (N_27699,N_27426,N_26753);
or U27700 (N_27700,N_26530,N_26448);
nor U27701 (N_27701,N_27033,N_26922);
nand U27702 (N_27702,N_26556,N_27534);
or U27703 (N_27703,N_27218,N_27385);
xnor U27704 (N_27704,N_26911,N_26880);
nor U27705 (N_27705,N_27394,N_26441);
nor U27706 (N_27706,N_27122,N_26738);
nand U27707 (N_27707,N_26812,N_27587);
and U27708 (N_27708,N_27132,N_26592);
and U27709 (N_27709,N_27540,N_26979);
xnor U27710 (N_27710,N_27135,N_26891);
nor U27711 (N_27711,N_27273,N_27019);
or U27712 (N_27712,N_26467,N_27404);
and U27713 (N_27713,N_26693,N_26883);
xnor U27714 (N_27714,N_27310,N_26806);
or U27715 (N_27715,N_26951,N_27552);
and U27716 (N_27716,N_27420,N_27115);
nand U27717 (N_27717,N_27493,N_27028);
and U27718 (N_27718,N_27261,N_27541);
and U27719 (N_27719,N_27161,N_27391);
nor U27720 (N_27720,N_26846,N_27143);
nor U27721 (N_27721,N_27358,N_26598);
nor U27722 (N_27722,N_26771,N_27357);
and U27723 (N_27723,N_26578,N_27320);
or U27724 (N_27724,N_27498,N_26702);
and U27725 (N_27725,N_27383,N_27542);
and U27726 (N_27726,N_27409,N_27048);
or U27727 (N_27727,N_26490,N_26721);
and U27728 (N_27728,N_27437,N_27129);
and U27729 (N_27729,N_26485,N_26968);
nor U27730 (N_27730,N_27021,N_27269);
nand U27731 (N_27731,N_26521,N_27349);
and U27732 (N_27732,N_27275,N_27413);
xor U27733 (N_27733,N_26746,N_26773);
or U27734 (N_27734,N_27387,N_27338);
or U27735 (N_27735,N_27150,N_26590);
nand U27736 (N_27736,N_27570,N_27224);
nor U27737 (N_27737,N_26542,N_27219);
and U27738 (N_27738,N_26895,N_26491);
or U27739 (N_27739,N_27347,N_27422);
and U27740 (N_27740,N_27398,N_26890);
nor U27741 (N_27741,N_26737,N_26886);
nor U27742 (N_27742,N_26468,N_26458);
and U27743 (N_27743,N_27564,N_27482);
nor U27744 (N_27744,N_26768,N_27531);
xnor U27745 (N_27745,N_26534,N_27399);
xnor U27746 (N_27746,N_26413,N_26674);
nand U27747 (N_27747,N_26778,N_26671);
xor U27748 (N_27748,N_27465,N_27524);
or U27749 (N_27749,N_26594,N_27074);
and U27750 (N_27750,N_26967,N_27484);
nand U27751 (N_27751,N_27179,N_27223);
nor U27752 (N_27752,N_27478,N_26647);
and U27753 (N_27753,N_26579,N_27480);
nand U27754 (N_27754,N_27554,N_27274);
xor U27755 (N_27755,N_27206,N_27189);
nand U27756 (N_27756,N_27263,N_27226);
or U27757 (N_27757,N_26774,N_27473);
nor U27758 (N_27758,N_26990,N_27451);
nand U27759 (N_27759,N_27014,N_27242);
or U27760 (N_27760,N_27003,N_26506);
nor U27761 (N_27761,N_27363,N_26735);
nor U27762 (N_27762,N_26412,N_27543);
and U27763 (N_27763,N_27067,N_27421);
nand U27764 (N_27764,N_27503,N_26945);
xnor U27765 (N_27765,N_27533,N_26462);
nor U27766 (N_27766,N_26428,N_27331);
or U27767 (N_27767,N_27509,N_26430);
or U27768 (N_27768,N_26493,N_27280);
nor U27769 (N_27769,N_26759,N_27237);
xnor U27770 (N_27770,N_26963,N_27481);
or U27771 (N_27771,N_26642,N_26697);
nor U27772 (N_27772,N_26994,N_27158);
nor U27773 (N_27773,N_26453,N_27515);
or U27774 (N_27774,N_26554,N_27510);
xor U27775 (N_27775,N_27359,N_27474);
nor U27776 (N_27776,N_27215,N_26495);
and U27777 (N_27777,N_26615,N_27319);
and U27778 (N_27778,N_26636,N_27448);
and U27779 (N_27779,N_26618,N_27351);
nor U27780 (N_27780,N_27217,N_26619);
nand U27781 (N_27781,N_26849,N_27303);
and U27782 (N_27782,N_27031,N_27479);
xnor U27783 (N_27783,N_27051,N_27428);
nand U27784 (N_27784,N_27137,N_27070);
or U27785 (N_27785,N_26587,N_27186);
or U27786 (N_27786,N_26553,N_26489);
nand U27787 (N_27787,N_27468,N_26708);
nand U27788 (N_27788,N_26459,N_26421);
xnor U27789 (N_27789,N_26711,N_27467);
or U27790 (N_27790,N_26871,N_27599);
nor U27791 (N_27791,N_26563,N_26570);
or U27792 (N_27792,N_27430,N_26832);
nand U27793 (N_27793,N_26474,N_26903);
and U27794 (N_27794,N_27294,N_27544);
xnor U27795 (N_27795,N_27252,N_26976);
xor U27796 (N_27796,N_27027,N_27536);
and U27797 (N_27797,N_26998,N_26977);
or U27798 (N_27798,N_27107,N_26853);
and U27799 (N_27799,N_27000,N_27317);
nand U27800 (N_27800,N_27301,N_26607);
nor U27801 (N_27801,N_27379,N_27314);
xor U27802 (N_27802,N_26947,N_26498);
xnor U27803 (N_27803,N_26438,N_27400);
xnor U27804 (N_27804,N_27160,N_27288);
nor U27805 (N_27805,N_26507,N_27134);
nand U27806 (N_27806,N_27131,N_26809);
or U27807 (N_27807,N_26596,N_27284);
nand U27808 (N_27808,N_27095,N_26703);
and U27809 (N_27809,N_26544,N_27165);
and U27810 (N_27810,N_27417,N_26681);
and U27811 (N_27811,N_26827,N_27266);
and U27812 (N_27812,N_26589,N_27300);
nand U27813 (N_27813,N_27374,N_27056);
nand U27814 (N_27814,N_27485,N_27058);
and U27815 (N_27815,N_26793,N_26783);
nand U27816 (N_27816,N_27336,N_26622);
and U27817 (N_27817,N_27327,N_27339);
nor U27818 (N_27818,N_27380,N_26678);
nand U27819 (N_27819,N_26571,N_27091);
nor U27820 (N_27820,N_26665,N_26502);
and U27821 (N_27821,N_26403,N_27576);
or U27822 (N_27822,N_26555,N_26720);
xnor U27823 (N_27823,N_26881,N_26576);
nor U27824 (N_27824,N_26402,N_26789);
nand U27825 (N_27825,N_27305,N_26912);
or U27826 (N_27826,N_27201,N_26608);
and U27827 (N_27827,N_27415,N_27198);
xor U27828 (N_27828,N_27360,N_26796);
and U27829 (N_27829,N_26957,N_26645);
nor U27830 (N_27830,N_26799,N_26509);
and U27831 (N_27831,N_26444,N_27549);
nand U27832 (N_27832,N_26864,N_27167);
nor U27833 (N_27833,N_26609,N_26582);
xnor U27834 (N_27834,N_26548,N_26541);
or U27835 (N_27835,N_26794,N_26758);
nor U27836 (N_27836,N_26829,N_27243);
xor U27837 (N_27837,N_26861,N_26457);
nand U27838 (N_27838,N_27087,N_27030);
nor U27839 (N_27839,N_27105,N_26836);
nand U27840 (N_27840,N_26987,N_26902);
xnor U27841 (N_27841,N_26700,N_26725);
xor U27842 (N_27842,N_27155,N_27560);
and U27843 (N_27843,N_27532,N_26602);
or U27844 (N_27844,N_27225,N_26942);
xnor U27845 (N_27845,N_27411,N_27568);
xnor U27846 (N_27846,N_27401,N_26776);
and U27847 (N_27847,N_27289,N_26476);
and U27848 (N_27848,N_27246,N_27488);
xnor U27849 (N_27849,N_27395,N_26915);
and U27850 (N_27850,N_27156,N_26687);
or U27851 (N_27851,N_27034,N_26632);
or U27852 (N_27852,N_26802,N_27211);
or U27853 (N_27853,N_26522,N_26868);
xor U27854 (N_27854,N_26442,N_26888);
and U27855 (N_27855,N_27236,N_26862);
and U27856 (N_27856,N_26744,N_26480);
nor U27857 (N_27857,N_27248,N_26717);
or U27858 (N_27858,N_27290,N_27439);
xor U27859 (N_27859,N_26850,N_26762);
or U27860 (N_27860,N_27123,N_27085);
xnor U27861 (N_27861,N_26934,N_27092);
and U27862 (N_27862,N_26780,N_27450);
nand U27863 (N_27863,N_27169,N_26549);
and U27864 (N_27864,N_27362,N_26892);
xor U27865 (N_27865,N_27517,N_27334);
nand U27866 (N_27866,N_27210,N_27550);
nor U27867 (N_27867,N_27523,N_26401);
xnor U27868 (N_27868,N_27453,N_26897);
nor U27869 (N_27869,N_27538,N_26482);
or U27870 (N_27870,N_27403,N_26821);
nor U27871 (N_27871,N_26907,N_27208);
xor U27872 (N_27872,N_26691,N_27016);
and U27873 (N_27873,N_27520,N_27487);
nor U27874 (N_27874,N_26630,N_26787);
and U27875 (N_27875,N_26701,N_26497);
xor U27876 (N_27876,N_26918,N_26527);
nor U27877 (N_27877,N_26845,N_27494);
xor U27878 (N_27878,N_26848,N_27307);
nor U27879 (N_27879,N_26705,N_26734);
nand U27880 (N_27880,N_26488,N_27256);
or U27881 (N_27881,N_27348,N_27513);
nand U27882 (N_27882,N_26761,N_27558);
and U27883 (N_27883,N_26882,N_26477);
and U27884 (N_27884,N_26695,N_26991);
nor U27885 (N_27885,N_26677,N_27010);
nor U27886 (N_27886,N_27504,N_27311);
and U27887 (N_27887,N_27125,N_26755);
and U27888 (N_27888,N_27518,N_26501);
nand U27889 (N_27889,N_27229,N_26978);
or U27890 (N_27890,N_27203,N_27177);
xor U27891 (N_27891,N_27397,N_26616);
xnor U27892 (N_27892,N_27326,N_27191);
xor U27893 (N_27893,N_27323,N_26686);
and U27894 (N_27894,N_26639,N_27370);
nor U27895 (N_27895,N_26624,N_26852);
nand U27896 (N_27896,N_27088,N_26860);
nand U27897 (N_27897,N_26770,N_26601);
xor U27898 (N_27898,N_27262,N_27440);
nor U27899 (N_27899,N_26575,N_27133);
nand U27900 (N_27900,N_26574,N_27381);
xnor U27901 (N_27901,N_26651,N_26649);
nor U27902 (N_27902,N_26840,N_27388);
or U27903 (N_27903,N_26633,N_27232);
nand U27904 (N_27904,N_26964,N_27454);
and U27905 (N_27905,N_26989,N_27152);
xor U27906 (N_27906,N_26971,N_27227);
nor U27907 (N_27907,N_26533,N_26584);
and U27908 (N_27908,N_27234,N_26839);
nor U27909 (N_27909,N_26803,N_26820);
xnor U27910 (N_27910,N_27384,N_26739);
nor U27911 (N_27911,N_27572,N_26914);
xnor U27912 (N_27912,N_26440,N_27283);
nand U27913 (N_27913,N_27597,N_27071);
nand U27914 (N_27914,N_27306,N_26707);
nor U27915 (N_27915,N_26784,N_26411);
nand U27916 (N_27916,N_27535,N_26675);
and U27917 (N_27917,N_26932,N_27060);
nor U27918 (N_27918,N_26631,N_26673);
and U27919 (N_27919,N_27431,N_26560);
and U27920 (N_27920,N_27445,N_27304);
and U27921 (N_27921,N_27268,N_26805);
nand U27922 (N_27922,N_27166,N_27516);
nand U27923 (N_27923,N_27146,N_26733);
or U27924 (N_27924,N_26996,N_27569);
xnor U27925 (N_27925,N_27299,N_27508);
xor U27926 (N_27926,N_27142,N_27527);
nor U27927 (N_27927,N_27278,N_27461);
nand U27928 (N_27928,N_27287,N_26625);
nor U27929 (N_27929,N_27455,N_26514);
or U27930 (N_27930,N_26405,N_26785);
or U27931 (N_27931,N_26919,N_26668);
nor U27932 (N_27932,N_26433,N_27015);
nand U27933 (N_27933,N_27462,N_27207);
or U27934 (N_27934,N_26407,N_27062);
or U27935 (N_27935,N_27355,N_26817);
nor U27936 (N_27936,N_26450,N_27118);
and U27937 (N_27937,N_27180,N_27079);
nor U27938 (N_27938,N_26825,N_26525);
and U27939 (N_27939,N_27017,N_27205);
nand U27940 (N_27940,N_26690,N_26908);
nand U27941 (N_27941,N_26604,N_27393);
xnor U27942 (N_27942,N_27157,N_26680);
xnor U27943 (N_27943,N_27457,N_27130);
and U27944 (N_27944,N_27563,N_26567);
nor U27945 (N_27945,N_27368,N_26551);
or U27946 (N_27946,N_27586,N_26545);
xor U27947 (N_27947,N_27257,N_26807);
nor U27948 (N_27948,N_26779,N_26916);
or U27949 (N_27949,N_27001,N_26767);
or U27950 (N_27950,N_27419,N_27584);
or U27951 (N_27951,N_26920,N_27332);
or U27952 (N_27952,N_26463,N_26538);
or U27953 (N_27953,N_26515,N_27061);
nand U27954 (N_27954,N_26764,N_26727);
xnor U27955 (N_27955,N_26826,N_26558);
and U27956 (N_27956,N_27276,N_26939);
nand U27957 (N_27957,N_27562,N_26801);
nor U27958 (N_27958,N_27222,N_27459);
xnor U27959 (N_27959,N_27501,N_27011);
nor U27960 (N_27960,N_27593,N_26855);
nor U27961 (N_27961,N_27298,N_26841);
or U27962 (N_27962,N_26757,N_27113);
and U27963 (N_27963,N_26999,N_27209);
or U27964 (N_27964,N_27068,N_27392);
or U27965 (N_27965,N_27047,N_26469);
xor U27966 (N_27966,N_26550,N_27486);
or U27967 (N_27967,N_27312,N_27553);
and U27968 (N_27968,N_26756,N_26454);
and U27969 (N_27969,N_27106,N_26722);
or U27970 (N_27970,N_26791,N_27221);
and U27971 (N_27971,N_26901,N_27446);
or U27972 (N_27972,N_27499,N_27309);
nor U27973 (N_27973,N_27565,N_26896);
xor U27974 (N_27974,N_27502,N_27436);
or U27975 (N_27975,N_27505,N_27471);
nand U27976 (N_27976,N_26749,N_26972);
nor U27977 (N_27977,N_27286,N_26935);
xnor U27978 (N_27978,N_27185,N_26419);
nor U27979 (N_27979,N_26648,N_27447);
xor U27980 (N_27980,N_27571,N_27053);
xor U27981 (N_27981,N_26754,N_26415);
nor U27982 (N_27982,N_26593,N_27110);
or U27983 (N_27983,N_26870,N_26585);
xor U27984 (N_27984,N_26662,N_27080);
and U27985 (N_27985,N_27495,N_26466);
and U27986 (N_27986,N_27316,N_27476);
or U27987 (N_27987,N_27006,N_26698);
xnor U27988 (N_27988,N_27136,N_26414);
nand U27989 (N_27989,N_27199,N_26966);
and U27990 (N_27990,N_26742,N_26682);
xnor U27991 (N_27991,N_27500,N_26547);
nor U27992 (N_27992,N_27396,N_27159);
nand U27993 (N_27993,N_27581,N_26718);
nor U27994 (N_27994,N_26859,N_27036);
xor U27995 (N_27995,N_26656,N_27475);
and U27996 (N_27996,N_27296,N_26940);
nor U27997 (N_27997,N_27466,N_27342);
xnor U27998 (N_27998,N_26503,N_27585);
or U27999 (N_27999,N_26887,N_26537);
nand U28000 (N_28000,N_26620,N_27353);
nand U28001 (N_28001,N_26731,N_26913);
xor U28002 (N_28002,N_26834,N_27141);
xor U28003 (N_28003,N_26813,N_27041);
nor U28004 (N_28004,N_27114,N_26930);
and U28005 (N_28005,N_27574,N_26962);
nand U28006 (N_28006,N_27188,N_27270);
nand U28007 (N_28007,N_27032,N_27216);
nor U28008 (N_28008,N_27081,N_27254);
xnor U28009 (N_28009,N_26659,N_26461);
xnor U28010 (N_28010,N_27045,N_27170);
and U28011 (N_28011,N_26435,N_27483);
xor U28012 (N_28012,N_26993,N_27337);
nand U28013 (N_28013,N_26566,N_27057);
and U28014 (N_28014,N_27230,N_26606);
nand U28015 (N_28015,N_26980,N_26905);
and U28016 (N_28016,N_26464,N_26726);
or U28017 (N_28017,N_26706,N_26676);
and U28018 (N_28018,N_27054,N_27120);
or U28019 (N_28019,N_27364,N_27064);
xor U28020 (N_28020,N_27202,N_26565);
or U28021 (N_28021,N_26564,N_26451);
xnor U28022 (N_28022,N_27595,N_26960);
nor U28023 (N_28023,N_27341,N_26741);
nor U28024 (N_28024,N_26432,N_27424);
or U28025 (N_28025,N_26874,N_26876);
nand U28026 (N_28026,N_26894,N_26470);
nand U28027 (N_28027,N_26577,N_26483);
or U28028 (N_28028,N_27555,N_26614);
nor U28029 (N_28029,N_26472,N_26728);
nor U28030 (N_28030,N_27138,N_27583);
xnor U28031 (N_28031,N_26748,N_26869);
or U28032 (N_28032,N_26724,N_26657);
or U28033 (N_28033,N_27102,N_27402);
nand U28034 (N_28034,N_27194,N_27260);
or U28035 (N_28035,N_26487,N_26719);
nor U28036 (N_28036,N_26486,N_27514);
nor U28037 (N_28037,N_27598,N_26959);
nor U28038 (N_28038,N_27111,N_26628);
xnor U28039 (N_28039,N_27238,N_27490);
xor U28040 (N_28040,N_27477,N_27007);
xnor U28041 (N_28041,N_27255,N_26824);
or U28042 (N_28042,N_27196,N_27176);
or U28043 (N_28043,N_26723,N_27163);
and U28044 (N_28044,N_27376,N_27241);
or U28045 (N_28045,N_27077,N_26404);
nand U28046 (N_28046,N_27406,N_26591);
nand U28047 (N_28047,N_26672,N_26879);
and U28048 (N_28048,N_27008,N_26546);
xnor U28049 (N_28049,N_27366,N_26536);
nor U28050 (N_28050,N_26410,N_26623);
and U28051 (N_28051,N_27464,N_27090);
xor U28052 (N_28052,N_27049,N_26823);
and U28053 (N_28053,N_27174,N_27097);
xor U28054 (N_28054,N_26667,N_26400);
nand U28055 (N_28055,N_26933,N_27452);
nor U28056 (N_28056,N_26736,N_27121);
xnor U28057 (N_28057,N_26709,N_27104);
xor U28058 (N_28058,N_26712,N_26713);
xnor U28059 (N_28059,N_27588,N_27259);
xor U28060 (N_28060,N_26475,N_26772);
and U28061 (N_28061,N_27126,N_26478);
nand U28062 (N_28062,N_27330,N_26561);
xnor U28063 (N_28063,N_26699,N_27190);
and U28064 (N_28064,N_27020,N_26949);
nor U28065 (N_28065,N_26814,N_26455);
xnor U28066 (N_28066,N_27195,N_27213);
xor U28067 (N_28067,N_26526,N_27042);
nand U28068 (N_28068,N_26621,N_27258);
or U28069 (N_28069,N_27247,N_27548);
nand U28070 (N_28070,N_27577,N_26936);
xnor U28071 (N_28071,N_27390,N_27361);
xor U28072 (N_28072,N_27172,N_26409);
xor U28073 (N_28073,N_27059,N_27103);
and U28074 (N_28074,N_26528,N_27521);
or U28075 (N_28075,N_27108,N_27519);
nor U28076 (N_28076,N_26679,N_27183);
or U28077 (N_28077,N_26997,N_27489);
nor U28078 (N_28078,N_26611,N_27181);
nor U28079 (N_28079,N_27200,N_26535);
nand U28080 (N_28080,N_26429,N_27119);
or U28081 (N_28081,N_26529,N_26417);
nand U28082 (N_28082,N_26865,N_26666);
xnor U28083 (N_28083,N_27389,N_26884);
nor U28084 (N_28084,N_26714,N_26909);
nor U28085 (N_28085,N_26760,N_27438);
and U28086 (N_28086,N_27365,N_27425);
or U28087 (N_28087,N_26583,N_26866);
nor U28088 (N_28088,N_27037,N_27094);
or U28089 (N_28089,N_27023,N_27046);
nor U28090 (N_28090,N_27318,N_26692);
nor U28091 (N_28091,N_27147,N_26766);
or U28092 (N_28092,N_27511,N_27295);
nor U28093 (N_28093,N_26661,N_27267);
nor U28094 (N_28094,N_26654,N_27427);
or U28095 (N_28095,N_27302,N_27281);
nand U28096 (N_28096,N_27093,N_27497);
nor U28097 (N_28097,N_26446,N_26447);
xor U28098 (N_28098,N_26710,N_27075);
xnor U28099 (N_28099,N_26670,N_26694);
or U28100 (N_28100,N_27162,N_27293);
nor U28101 (N_28101,N_27148,N_27083);
xnor U28102 (N_28102,N_27149,N_27175);
nand U28103 (N_28103,N_26818,N_26627);
xnor U28104 (N_28104,N_26518,N_27251);
or U28105 (N_28105,N_27590,N_27250);
or U28106 (N_28106,N_27566,N_26950);
and U28107 (N_28107,N_26650,N_27371);
or U28108 (N_28108,N_26985,N_26956);
nor U28109 (N_28109,N_26603,N_27432);
xor U28110 (N_28110,N_27116,N_26872);
xor U28111 (N_28111,N_26572,N_26798);
nor U28112 (N_28112,N_27128,N_26641);
nor U28113 (N_28113,N_26500,N_26775);
xnor U28114 (N_28114,N_27443,N_26481);
nand U28115 (N_28115,N_26747,N_27378);
nor U28116 (N_28116,N_26974,N_26408);
xor U28117 (N_28117,N_26658,N_27096);
or U28118 (N_28118,N_27329,N_26644);
nor U28119 (N_28119,N_27086,N_26704);
and U28120 (N_28120,N_26863,N_26808);
or U28121 (N_28121,N_26629,N_26800);
nand U28122 (N_28122,N_26512,N_27308);
nand U28123 (N_28123,N_26437,N_27272);
nand U28124 (N_28124,N_27239,N_27012);
and U28125 (N_28125,N_26983,N_27512);
nand U28126 (N_28126,N_26790,N_26422);
nor U28127 (N_28127,N_26643,N_26751);
nor U28128 (N_28128,N_26669,N_26822);
xor U28129 (N_28129,N_26926,N_26851);
or U28130 (N_28130,N_26683,N_26944);
nand U28131 (N_28131,N_27491,N_26837);
or U28132 (N_28132,N_26513,N_27050);
and U28133 (N_28133,N_27345,N_27460);
nor U28134 (N_28134,N_26929,N_27556);
and U28135 (N_28135,N_27333,N_27350);
xor U28136 (N_28136,N_27233,N_27375);
and U28137 (N_28137,N_26769,N_26597);
or U28138 (N_28138,N_26479,N_27546);
nor U28139 (N_28139,N_26568,N_26740);
xnor U28140 (N_28140,N_26612,N_26418);
nor U28141 (N_28141,N_27354,N_27182);
xnor U28142 (N_28142,N_26540,N_27507);
nand U28143 (N_28143,N_27171,N_26857);
nand U28144 (N_28144,N_26586,N_26559);
xor U28145 (N_28145,N_27151,N_27264);
nand U28146 (N_28146,N_27526,N_26854);
nand U28147 (N_28147,N_26684,N_27321);
and U28148 (N_28148,N_27109,N_26943);
xor U28149 (N_28149,N_27082,N_26925);
or U28150 (N_28150,N_26646,N_27117);
nor U28151 (N_28151,N_26452,N_26508);
xnor U28152 (N_28152,N_27492,N_26532);
xor U28153 (N_28153,N_26425,N_26752);
and U28154 (N_28154,N_26965,N_27253);
nand U28155 (N_28155,N_26484,N_27063);
or U28156 (N_28156,N_27285,N_27414);
and U28157 (N_28157,N_26696,N_27072);
and U28158 (N_28158,N_26605,N_27271);
xnor U28159 (N_28159,N_27144,N_26937);
xor U28160 (N_28160,N_27127,N_27496);
or U28161 (N_28161,N_26906,N_27100);
nor U28162 (N_28162,N_26663,N_26952);
or U28163 (N_28163,N_27435,N_26970);
and U28164 (N_28164,N_27423,N_27547);
xnor U28165 (N_28165,N_26496,N_27506);
xor U28166 (N_28166,N_26804,N_26830);
or U28167 (N_28167,N_27291,N_27592);
or U28168 (N_28168,N_27539,N_27463);
nor U28169 (N_28169,N_27596,N_27582);
xor U28170 (N_28170,N_27187,N_26975);
nand U28171 (N_28171,N_27026,N_27265);
nand U28172 (N_28172,N_27066,N_26954);
nor U28173 (N_28173,N_26782,N_26573);
nor U28174 (N_28174,N_26416,N_26877);
and U28175 (N_28175,N_26833,N_27575);
xor U28176 (N_28176,N_26640,N_26889);
xor U28177 (N_28177,N_26781,N_26689);
or U28178 (N_28178,N_27551,N_26613);
nor U28179 (N_28179,N_26898,N_26510);
or U28180 (N_28180,N_26988,N_26634);
xnor U28181 (N_28181,N_27442,N_27449);
or U28182 (N_28182,N_26885,N_27153);
and U28183 (N_28183,N_26652,N_27164);
or U28184 (N_28184,N_26406,N_27140);
nand U28185 (N_28185,N_26424,N_27245);
or U28186 (N_28186,N_27529,N_27168);
and U28187 (N_28187,N_26580,N_27084);
xnor U28188 (N_28188,N_27537,N_27073);
nor U28189 (N_28189,N_26788,N_27035);
or U28190 (N_28190,N_26948,N_26844);
and U28191 (N_28191,N_26473,N_27279);
or U28192 (N_28192,N_26519,N_26581);
or U28193 (N_28193,N_27282,N_27335);
or U28194 (N_28194,N_26730,N_27591);
nor U28195 (N_28195,N_27178,N_27101);
nand U28196 (N_28196,N_27173,N_26917);
nand U28197 (N_28197,N_26569,N_26931);
and U28198 (N_28198,N_27346,N_27561);
nor U28199 (N_28199,N_27441,N_27197);
nand U28200 (N_28200,N_26433,N_26592);
xnor U28201 (N_28201,N_27240,N_27137);
nand U28202 (N_28202,N_27537,N_26890);
or U28203 (N_28203,N_26913,N_27370);
or U28204 (N_28204,N_27066,N_27503);
nor U28205 (N_28205,N_27008,N_27131);
and U28206 (N_28206,N_27451,N_27055);
nor U28207 (N_28207,N_27352,N_26748);
nand U28208 (N_28208,N_27128,N_27405);
and U28209 (N_28209,N_26655,N_27270);
nand U28210 (N_28210,N_26927,N_27550);
nor U28211 (N_28211,N_26822,N_27088);
and U28212 (N_28212,N_26909,N_27038);
nand U28213 (N_28213,N_27418,N_27532);
xor U28214 (N_28214,N_26424,N_27469);
or U28215 (N_28215,N_26815,N_27093);
xor U28216 (N_28216,N_27553,N_26930);
xnor U28217 (N_28217,N_27141,N_27387);
nand U28218 (N_28218,N_27001,N_26495);
xor U28219 (N_28219,N_26478,N_26919);
and U28220 (N_28220,N_27392,N_26479);
xnor U28221 (N_28221,N_26808,N_27595);
xnor U28222 (N_28222,N_26995,N_27584);
nand U28223 (N_28223,N_27256,N_27420);
nand U28224 (N_28224,N_26992,N_26506);
nor U28225 (N_28225,N_26545,N_27472);
nor U28226 (N_28226,N_26814,N_26641);
and U28227 (N_28227,N_26888,N_27230);
nor U28228 (N_28228,N_26866,N_26572);
xor U28229 (N_28229,N_27443,N_27046);
xnor U28230 (N_28230,N_27018,N_27183);
and U28231 (N_28231,N_27160,N_26526);
nor U28232 (N_28232,N_27203,N_27183);
xnor U28233 (N_28233,N_27104,N_26963);
and U28234 (N_28234,N_26626,N_27472);
or U28235 (N_28235,N_26868,N_27438);
nor U28236 (N_28236,N_26798,N_26503);
xor U28237 (N_28237,N_26808,N_26697);
and U28238 (N_28238,N_27356,N_27255);
and U28239 (N_28239,N_26851,N_26750);
or U28240 (N_28240,N_26695,N_27263);
nor U28241 (N_28241,N_26911,N_26648);
nand U28242 (N_28242,N_26642,N_26971);
xnor U28243 (N_28243,N_26845,N_26805);
nor U28244 (N_28244,N_27463,N_27587);
and U28245 (N_28245,N_26446,N_26677);
xor U28246 (N_28246,N_26848,N_27506);
or U28247 (N_28247,N_27350,N_26724);
and U28248 (N_28248,N_27525,N_27574);
nand U28249 (N_28249,N_27597,N_27246);
nor U28250 (N_28250,N_26982,N_27251);
nor U28251 (N_28251,N_27315,N_27456);
xnor U28252 (N_28252,N_26443,N_26431);
nor U28253 (N_28253,N_27442,N_27010);
or U28254 (N_28254,N_26504,N_26884);
xnor U28255 (N_28255,N_27482,N_27010);
xor U28256 (N_28256,N_26533,N_27125);
xor U28257 (N_28257,N_26727,N_26431);
nand U28258 (N_28258,N_26621,N_27270);
and U28259 (N_28259,N_27157,N_26898);
nand U28260 (N_28260,N_27243,N_26642);
nand U28261 (N_28261,N_26891,N_27461);
nor U28262 (N_28262,N_27268,N_27405);
nand U28263 (N_28263,N_26457,N_26992);
or U28264 (N_28264,N_26620,N_26945);
nand U28265 (N_28265,N_27009,N_27322);
or U28266 (N_28266,N_27438,N_26484);
xnor U28267 (N_28267,N_27411,N_26820);
or U28268 (N_28268,N_26784,N_26780);
nor U28269 (N_28269,N_26996,N_26559);
nor U28270 (N_28270,N_27276,N_27568);
nor U28271 (N_28271,N_27480,N_27097);
or U28272 (N_28272,N_27079,N_27413);
nand U28273 (N_28273,N_27138,N_27495);
or U28274 (N_28274,N_26997,N_26501);
nor U28275 (N_28275,N_27022,N_26495);
xnor U28276 (N_28276,N_26775,N_27255);
or U28277 (N_28277,N_26966,N_27528);
or U28278 (N_28278,N_27374,N_27407);
and U28279 (N_28279,N_26805,N_27456);
xnor U28280 (N_28280,N_27101,N_27017);
and U28281 (N_28281,N_26894,N_27281);
or U28282 (N_28282,N_26845,N_27120);
nor U28283 (N_28283,N_27507,N_27262);
nand U28284 (N_28284,N_26845,N_26590);
nor U28285 (N_28285,N_27368,N_27562);
nor U28286 (N_28286,N_26745,N_27378);
or U28287 (N_28287,N_26672,N_27429);
nand U28288 (N_28288,N_27305,N_26969);
xor U28289 (N_28289,N_26609,N_26636);
xnor U28290 (N_28290,N_27176,N_27276);
nand U28291 (N_28291,N_27534,N_27543);
nor U28292 (N_28292,N_26798,N_27259);
and U28293 (N_28293,N_26684,N_26423);
xor U28294 (N_28294,N_26720,N_27259);
xor U28295 (N_28295,N_26473,N_26781);
nor U28296 (N_28296,N_26639,N_26633);
xor U28297 (N_28297,N_26801,N_27199);
and U28298 (N_28298,N_26455,N_27113);
xor U28299 (N_28299,N_26725,N_27172);
or U28300 (N_28300,N_26772,N_27103);
or U28301 (N_28301,N_27303,N_27349);
or U28302 (N_28302,N_27033,N_27246);
and U28303 (N_28303,N_27009,N_27073);
nor U28304 (N_28304,N_27178,N_27405);
nor U28305 (N_28305,N_26907,N_26952);
nand U28306 (N_28306,N_27104,N_26553);
nand U28307 (N_28307,N_26609,N_26480);
xnor U28308 (N_28308,N_26989,N_27305);
nor U28309 (N_28309,N_26626,N_26602);
xor U28310 (N_28310,N_27204,N_26940);
or U28311 (N_28311,N_27208,N_26428);
and U28312 (N_28312,N_26599,N_26903);
and U28313 (N_28313,N_27512,N_27398);
nand U28314 (N_28314,N_27484,N_27075);
and U28315 (N_28315,N_26722,N_26725);
nor U28316 (N_28316,N_27156,N_26680);
and U28317 (N_28317,N_27424,N_27238);
nor U28318 (N_28318,N_27235,N_27232);
xor U28319 (N_28319,N_27411,N_26566);
nand U28320 (N_28320,N_26832,N_26838);
nand U28321 (N_28321,N_26652,N_27233);
xor U28322 (N_28322,N_26429,N_26716);
xor U28323 (N_28323,N_27555,N_27508);
nand U28324 (N_28324,N_26512,N_27569);
and U28325 (N_28325,N_26622,N_26866);
and U28326 (N_28326,N_27510,N_27065);
nor U28327 (N_28327,N_27010,N_26443);
nor U28328 (N_28328,N_26895,N_26673);
nand U28329 (N_28329,N_27253,N_27563);
nand U28330 (N_28330,N_26515,N_27424);
nand U28331 (N_28331,N_26883,N_26447);
xor U28332 (N_28332,N_27311,N_27521);
xnor U28333 (N_28333,N_27501,N_26721);
nor U28334 (N_28334,N_27330,N_27269);
and U28335 (N_28335,N_27105,N_27275);
nor U28336 (N_28336,N_27273,N_27534);
or U28337 (N_28337,N_27199,N_26695);
nand U28338 (N_28338,N_26985,N_27319);
nor U28339 (N_28339,N_26710,N_26585);
or U28340 (N_28340,N_26804,N_26808);
xnor U28341 (N_28341,N_27504,N_27276);
xnor U28342 (N_28342,N_26422,N_27550);
or U28343 (N_28343,N_26906,N_27031);
nor U28344 (N_28344,N_26613,N_27128);
nand U28345 (N_28345,N_26800,N_27372);
and U28346 (N_28346,N_27179,N_27057);
and U28347 (N_28347,N_27009,N_27163);
nor U28348 (N_28348,N_27198,N_27509);
and U28349 (N_28349,N_26943,N_27395);
xnor U28350 (N_28350,N_27416,N_26900);
and U28351 (N_28351,N_26456,N_27369);
nor U28352 (N_28352,N_26877,N_26563);
and U28353 (N_28353,N_27101,N_27053);
nand U28354 (N_28354,N_26963,N_27471);
nor U28355 (N_28355,N_26604,N_26534);
or U28356 (N_28356,N_26749,N_27003);
and U28357 (N_28357,N_27393,N_26895);
nand U28358 (N_28358,N_27044,N_27155);
nor U28359 (N_28359,N_27287,N_27495);
xnor U28360 (N_28360,N_26612,N_27377);
or U28361 (N_28361,N_26538,N_27026);
nand U28362 (N_28362,N_27454,N_27263);
nand U28363 (N_28363,N_27125,N_27025);
or U28364 (N_28364,N_26998,N_27251);
nand U28365 (N_28365,N_26741,N_26591);
or U28366 (N_28366,N_27223,N_26842);
nand U28367 (N_28367,N_26908,N_27287);
or U28368 (N_28368,N_26620,N_27310);
xnor U28369 (N_28369,N_26450,N_26609);
or U28370 (N_28370,N_27461,N_26515);
or U28371 (N_28371,N_27415,N_27406);
nor U28372 (N_28372,N_26724,N_26628);
nand U28373 (N_28373,N_26662,N_26794);
and U28374 (N_28374,N_27527,N_27195);
nand U28375 (N_28375,N_26641,N_26988);
xnor U28376 (N_28376,N_26779,N_26539);
xnor U28377 (N_28377,N_27125,N_26930);
nand U28378 (N_28378,N_27143,N_26971);
xor U28379 (N_28379,N_26959,N_26494);
nand U28380 (N_28380,N_26653,N_26900);
xor U28381 (N_28381,N_26531,N_27088);
or U28382 (N_28382,N_26768,N_27066);
and U28383 (N_28383,N_26961,N_27171);
and U28384 (N_28384,N_27496,N_26452);
nor U28385 (N_28385,N_27443,N_27114);
and U28386 (N_28386,N_27406,N_26484);
xor U28387 (N_28387,N_27142,N_26597);
nand U28388 (N_28388,N_27267,N_26883);
nand U28389 (N_28389,N_26406,N_27082);
and U28390 (N_28390,N_27509,N_26756);
or U28391 (N_28391,N_26851,N_27580);
or U28392 (N_28392,N_27447,N_26522);
nor U28393 (N_28393,N_27333,N_26462);
or U28394 (N_28394,N_27032,N_26805);
nand U28395 (N_28395,N_27100,N_26676);
nand U28396 (N_28396,N_27466,N_27213);
or U28397 (N_28397,N_27515,N_26577);
nor U28398 (N_28398,N_26702,N_26879);
and U28399 (N_28399,N_26494,N_26473);
nor U28400 (N_28400,N_27043,N_27040);
nor U28401 (N_28401,N_26984,N_26434);
nand U28402 (N_28402,N_27538,N_27428);
and U28403 (N_28403,N_26781,N_27040);
nor U28404 (N_28404,N_26823,N_26793);
nand U28405 (N_28405,N_27360,N_26798);
or U28406 (N_28406,N_27164,N_27550);
nand U28407 (N_28407,N_26772,N_27566);
nand U28408 (N_28408,N_27226,N_26484);
and U28409 (N_28409,N_26527,N_26816);
or U28410 (N_28410,N_27431,N_26527);
xnor U28411 (N_28411,N_26911,N_27250);
xnor U28412 (N_28412,N_27362,N_27335);
or U28413 (N_28413,N_26425,N_27355);
xor U28414 (N_28414,N_27545,N_26791);
and U28415 (N_28415,N_26636,N_26947);
nand U28416 (N_28416,N_27082,N_26945);
and U28417 (N_28417,N_26986,N_27478);
nor U28418 (N_28418,N_26749,N_26714);
and U28419 (N_28419,N_27018,N_27378);
nand U28420 (N_28420,N_26926,N_27002);
nand U28421 (N_28421,N_27162,N_27051);
or U28422 (N_28422,N_26520,N_26910);
xnor U28423 (N_28423,N_26557,N_26972);
nand U28424 (N_28424,N_27441,N_27274);
or U28425 (N_28425,N_26873,N_26606);
nand U28426 (N_28426,N_26826,N_27004);
nor U28427 (N_28427,N_27446,N_27251);
or U28428 (N_28428,N_26664,N_26877);
or U28429 (N_28429,N_26567,N_27027);
nand U28430 (N_28430,N_27158,N_26453);
nand U28431 (N_28431,N_27407,N_27452);
nor U28432 (N_28432,N_27589,N_26909);
xor U28433 (N_28433,N_26984,N_27005);
nor U28434 (N_28434,N_27237,N_27045);
nand U28435 (N_28435,N_27280,N_27585);
xnor U28436 (N_28436,N_26990,N_26992);
nand U28437 (N_28437,N_27142,N_26773);
nor U28438 (N_28438,N_26412,N_26446);
xnor U28439 (N_28439,N_26512,N_26699);
xor U28440 (N_28440,N_26656,N_26979);
nor U28441 (N_28441,N_26840,N_27124);
and U28442 (N_28442,N_26990,N_27044);
and U28443 (N_28443,N_26424,N_26763);
nor U28444 (N_28444,N_26716,N_26607);
or U28445 (N_28445,N_26696,N_27351);
or U28446 (N_28446,N_27314,N_27214);
nand U28447 (N_28447,N_27152,N_27492);
and U28448 (N_28448,N_27573,N_27163);
xor U28449 (N_28449,N_27146,N_27020);
or U28450 (N_28450,N_27379,N_27570);
xnor U28451 (N_28451,N_27583,N_26537);
nand U28452 (N_28452,N_27377,N_27409);
or U28453 (N_28453,N_27200,N_26642);
xnor U28454 (N_28454,N_27219,N_27581);
nand U28455 (N_28455,N_26837,N_26865);
and U28456 (N_28456,N_26717,N_27414);
xor U28457 (N_28457,N_27194,N_27230);
and U28458 (N_28458,N_26405,N_27413);
xor U28459 (N_28459,N_27418,N_27000);
and U28460 (N_28460,N_26459,N_27554);
xor U28461 (N_28461,N_27083,N_26790);
xor U28462 (N_28462,N_27366,N_27116);
and U28463 (N_28463,N_26868,N_27509);
and U28464 (N_28464,N_27599,N_27117);
or U28465 (N_28465,N_27093,N_26949);
and U28466 (N_28466,N_26807,N_26782);
nand U28467 (N_28467,N_26587,N_26835);
and U28468 (N_28468,N_27469,N_26937);
or U28469 (N_28469,N_27067,N_26733);
and U28470 (N_28470,N_27215,N_26931);
or U28471 (N_28471,N_27048,N_27455);
and U28472 (N_28472,N_26977,N_26792);
nor U28473 (N_28473,N_26502,N_27494);
nand U28474 (N_28474,N_27291,N_26873);
nand U28475 (N_28475,N_26484,N_27139);
and U28476 (N_28476,N_27595,N_27164);
xnor U28477 (N_28477,N_27474,N_26538);
xor U28478 (N_28478,N_26529,N_26525);
xor U28479 (N_28479,N_26971,N_26533);
nand U28480 (N_28480,N_26520,N_27410);
xor U28481 (N_28481,N_26876,N_26922);
and U28482 (N_28482,N_27497,N_27000);
or U28483 (N_28483,N_26697,N_26856);
and U28484 (N_28484,N_26803,N_27397);
nand U28485 (N_28485,N_26782,N_26883);
nor U28486 (N_28486,N_26906,N_26444);
xnor U28487 (N_28487,N_27476,N_26583);
nor U28488 (N_28488,N_27399,N_26480);
nand U28489 (N_28489,N_27463,N_26420);
nand U28490 (N_28490,N_26675,N_27490);
or U28491 (N_28491,N_27082,N_26702);
nor U28492 (N_28492,N_26879,N_26550);
and U28493 (N_28493,N_26978,N_26521);
and U28494 (N_28494,N_26741,N_27414);
xnor U28495 (N_28495,N_26838,N_27085);
and U28496 (N_28496,N_26943,N_27435);
and U28497 (N_28497,N_27399,N_27344);
nor U28498 (N_28498,N_27138,N_26549);
nor U28499 (N_28499,N_27393,N_27399);
nand U28500 (N_28500,N_27168,N_26937);
nand U28501 (N_28501,N_26617,N_27517);
nand U28502 (N_28502,N_26738,N_26852);
xor U28503 (N_28503,N_27151,N_26580);
and U28504 (N_28504,N_26860,N_27399);
nand U28505 (N_28505,N_27393,N_26446);
nor U28506 (N_28506,N_26622,N_27006);
xor U28507 (N_28507,N_26572,N_26545);
nor U28508 (N_28508,N_26521,N_26941);
nor U28509 (N_28509,N_26616,N_26406);
or U28510 (N_28510,N_27309,N_26926);
xor U28511 (N_28511,N_27527,N_27061);
and U28512 (N_28512,N_27048,N_26546);
and U28513 (N_28513,N_27382,N_27096);
and U28514 (N_28514,N_26559,N_27414);
nor U28515 (N_28515,N_26607,N_27579);
xnor U28516 (N_28516,N_26801,N_27433);
or U28517 (N_28517,N_26435,N_27570);
or U28518 (N_28518,N_27249,N_27541);
and U28519 (N_28519,N_26531,N_27141);
and U28520 (N_28520,N_26592,N_27041);
nor U28521 (N_28521,N_26583,N_26861);
xnor U28522 (N_28522,N_26480,N_27185);
or U28523 (N_28523,N_26658,N_26858);
nor U28524 (N_28524,N_27287,N_27016);
nand U28525 (N_28525,N_27163,N_26463);
and U28526 (N_28526,N_27379,N_26535);
and U28527 (N_28527,N_27068,N_27497);
nor U28528 (N_28528,N_27393,N_26415);
and U28529 (N_28529,N_26980,N_27429);
xor U28530 (N_28530,N_27462,N_26681);
or U28531 (N_28531,N_27019,N_27255);
and U28532 (N_28532,N_27577,N_27345);
nor U28533 (N_28533,N_27492,N_26638);
and U28534 (N_28534,N_26623,N_27161);
or U28535 (N_28535,N_27347,N_27242);
nand U28536 (N_28536,N_26707,N_27545);
and U28537 (N_28537,N_27271,N_26546);
nor U28538 (N_28538,N_27177,N_27195);
nand U28539 (N_28539,N_27387,N_27563);
xor U28540 (N_28540,N_27440,N_26651);
xnor U28541 (N_28541,N_27542,N_26969);
xor U28542 (N_28542,N_27204,N_27159);
nand U28543 (N_28543,N_27391,N_27131);
xnor U28544 (N_28544,N_27382,N_27400);
or U28545 (N_28545,N_27207,N_27047);
and U28546 (N_28546,N_26887,N_27558);
xor U28547 (N_28547,N_26955,N_27190);
nand U28548 (N_28548,N_26639,N_27247);
xnor U28549 (N_28549,N_27196,N_27487);
and U28550 (N_28550,N_27413,N_26830);
nor U28551 (N_28551,N_27497,N_27014);
nand U28552 (N_28552,N_27503,N_27377);
nor U28553 (N_28553,N_27319,N_27437);
xnor U28554 (N_28554,N_26476,N_27348);
nor U28555 (N_28555,N_27565,N_26909);
xnor U28556 (N_28556,N_27155,N_27394);
and U28557 (N_28557,N_26871,N_27117);
xnor U28558 (N_28558,N_27573,N_26662);
and U28559 (N_28559,N_27558,N_26549);
nand U28560 (N_28560,N_27550,N_27090);
nor U28561 (N_28561,N_26546,N_27295);
or U28562 (N_28562,N_26684,N_27093);
or U28563 (N_28563,N_27385,N_26916);
or U28564 (N_28564,N_26972,N_27153);
xnor U28565 (N_28565,N_27321,N_26891);
or U28566 (N_28566,N_27245,N_26951);
nor U28567 (N_28567,N_26467,N_27215);
or U28568 (N_28568,N_27176,N_27415);
nor U28569 (N_28569,N_27059,N_26448);
and U28570 (N_28570,N_26565,N_26973);
and U28571 (N_28571,N_26707,N_26564);
xor U28572 (N_28572,N_26605,N_26548);
xor U28573 (N_28573,N_27518,N_26577);
or U28574 (N_28574,N_26610,N_26885);
nor U28575 (N_28575,N_27196,N_27337);
nor U28576 (N_28576,N_26647,N_26724);
or U28577 (N_28577,N_27151,N_26486);
nor U28578 (N_28578,N_26561,N_27410);
nand U28579 (N_28579,N_26579,N_27364);
and U28580 (N_28580,N_27517,N_26690);
nor U28581 (N_28581,N_26511,N_27104);
or U28582 (N_28582,N_26640,N_27348);
nand U28583 (N_28583,N_26688,N_27057);
nor U28584 (N_28584,N_27000,N_26457);
xnor U28585 (N_28585,N_26845,N_27038);
or U28586 (N_28586,N_26513,N_26686);
xor U28587 (N_28587,N_26517,N_27316);
nand U28588 (N_28588,N_27550,N_27499);
nand U28589 (N_28589,N_26891,N_26787);
xnor U28590 (N_28590,N_27194,N_27295);
and U28591 (N_28591,N_26711,N_26417);
nor U28592 (N_28592,N_27515,N_26603);
or U28593 (N_28593,N_27208,N_27545);
nor U28594 (N_28594,N_27269,N_26516);
xnor U28595 (N_28595,N_27508,N_26975);
nand U28596 (N_28596,N_27037,N_27090);
xnor U28597 (N_28597,N_26545,N_26998);
nand U28598 (N_28598,N_26667,N_27368);
xnor U28599 (N_28599,N_26453,N_27302);
nand U28600 (N_28600,N_27568,N_27450);
xor U28601 (N_28601,N_27303,N_27283);
and U28602 (N_28602,N_26863,N_26744);
and U28603 (N_28603,N_26460,N_27237);
nor U28604 (N_28604,N_27447,N_26548);
and U28605 (N_28605,N_27311,N_27332);
or U28606 (N_28606,N_27448,N_27259);
nand U28607 (N_28607,N_27043,N_26762);
and U28608 (N_28608,N_26725,N_26833);
or U28609 (N_28609,N_26504,N_26593);
nand U28610 (N_28610,N_26411,N_26525);
and U28611 (N_28611,N_27113,N_26470);
xnor U28612 (N_28612,N_26897,N_26777);
nand U28613 (N_28613,N_27518,N_26995);
or U28614 (N_28614,N_27074,N_27179);
nor U28615 (N_28615,N_26934,N_26631);
and U28616 (N_28616,N_26930,N_26601);
and U28617 (N_28617,N_27371,N_26902);
xor U28618 (N_28618,N_26934,N_27265);
and U28619 (N_28619,N_27276,N_26479);
and U28620 (N_28620,N_27474,N_27458);
xnor U28621 (N_28621,N_26606,N_27216);
or U28622 (N_28622,N_26792,N_26417);
nand U28623 (N_28623,N_26413,N_27188);
xnor U28624 (N_28624,N_27059,N_27406);
xor U28625 (N_28625,N_27468,N_27510);
xnor U28626 (N_28626,N_26624,N_26400);
xnor U28627 (N_28627,N_26656,N_27301);
xor U28628 (N_28628,N_27527,N_26574);
xor U28629 (N_28629,N_27346,N_26715);
nand U28630 (N_28630,N_26509,N_26516);
and U28631 (N_28631,N_26785,N_27421);
or U28632 (N_28632,N_27456,N_27035);
xor U28633 (N_28633,N_27168,N_26532);
nand U28634 (N_28634,N_26453,N_27050);
nand U28635 (N_28635,N_27472,N_26638);
nand U28636 (N_28636,N_27595,N_27323);
and U28637 (N_28637,N_26605,N_26416);
nand U28638 (N_28638,N_27335,N_27507);
xnor U28639 (N_28639,N_26443,N_26516);
nand U28640 (N_28640,N_27561,N_26802);
or U28641 (N_28641,N_26620,N_26663);
nand U28642 (N_28642,N_26788,N_27041);
or U28643 (N_28643,N_27389,N_26588);
and U28644 (N_28644,N_27504,N_27438);
xor U28645 (N_28645,N_27297,N_26986);
and U28646 (N_28646,N_27416,N_27192);
and U28647 (N_28647,N_26790,N_26453);
or U28648 (N_28648,N_27488,N_26803);
xor U28649 (N_28649,N_27268,N_27450);
or U28650 (N_28650,N_26403,N_26839);
xor U28651 (N_28651,N_26932,N_26572);
and U28652 (N_28652,N_27060,N_26510);
or U28653 (N_28653,N_27133,N_27023);
nor U28654 (N_28654,N_26502,N_26980);
nand U28655 (N_28655,N_27527,N_26496);
or U28656 (N_28656,N_27501,N_27573);
xor U28657 (N_28657,N_27049,N_27079);
xor U28658 (N_28658,N_27017,N_27360);
xnor U28659 (N_28659,N_27203,N_26824);
nor U28660 (N_28660,N_26828,N_26863);
xnor U28661 (N_28661,N_27543,N_26852);
and U28662 (N_28662,N_27079,N_26581);
nand U28663 (N_28663,N_26867,N_26476);
nor U28664 (N_28664,N_27450,N_26992);
xor U28665 (N_28665,N_27024,N_27123);
nand U28666 (N_28666,N_27363,N_26854);
xor U28667 (N_28667,N_26715,N_27320);
or U28668 (N_28668,N_26865,N_26504);
xnor U28669 (N_28669,N_27379,N_27408);
nor U28670 (N_28670,N_27569,N_26486);
nand U28671 (N_28671,N_27484,N_27269);
nor U28672 (N_28672,N_27096,N_26499);
or U28673 (N_28673,N_26488,N_27378);
or U28674 (N_28674,N_26962,N_26443);
xor U28675 (N_28675,N_27001,N_26916);
xnor U28676 (N_28676,N_27566,N_26580);
nor U28677 (N_28677,N_27469,N_26567);
and U28678 (N_28678,N_26515,N_26732);
nand U28679 (N_28679,N_26600,N_26668);
nand U28680 (N_28680,N_27072,N_27195);
xor U28681 (N_28681,N_27395,N_26608);
or U28682 (N_28682,N_27445,N_26565);
nand U28683 (N_28683,N_27252,N_27568);
xor U28684 (N_28684,N_26493,N_26885);
or U28685 (N_28685,N_26792,N_26966);
or U28686 (N_28686,N_26464,N_26828);
xor U28687 (N_28687,N_26653,N_26651);
or U28688 (N_28688,N_26722,N_27441);
and U28689 (N_28689,N_26764,N_27487);
nor U28690 (N_28690,N_26782,N_26922);
and U28691 (N_28691,N_27548,N_26999);
nor U28692 (N_28692,N_26723,N_26687);
nand U28693 (N_28693,N_27104,N_27505);
nand U28694 (N_28694,N_26967,N_26899);
nor U28695 (N_28695,N_26529,N_26903);
xor U28696 (N_28696,N_27116,N_26883);
nor U28697 (N_28697,N_26643,N_26647);
nand U28698 (N_28698,N_26637,N_27557);
and U28699 (N_28699,N_27479,N_27549);
and U28700 (N_28700,N_27452,N_27317);
nand U28701 (N_28701,N_27231,N_27371);
nor U28702 (N_28702,N_27293,N_26646);
nor U28703 (N_28703,N_27591,N_26690);
nand U28704 (N_28704,N_27443,N_27421);
or U28705 (N_28705,N_26733,N_26913);
xnor U28706 (N_28706,N_27089,N_26803);
nand U28707 (N_28707,N_26487,N_27259);
nand U28708 (N_28708,N_27249,N_27444);
or U28709 (N_28709,N_26589,N_26810);
or U28710 (N_28710,N_26747,N_26476);
and U28711 (N_28711,N_27150,N_26922);
nor U28712 (N_28712,N_27519,N_27159);
nand U28713 (N_28713,N_26606,N_27355);
and U28714 (N_28714,N_27386,N_27192);
and U28715 (N_28715,N_26929,N_27259);
and U28716 (N_28716,N_26440,N_26532);
xor U28717 (N_28717,N_27008,N_26801);
xnor U28718 (N_28718,N_27268,N_27094);
and U28719 (N_28719,N_27507,N_26967);
nor U28720 (N_28720,N_26939,N_27434);
xnor U28721 (N_28721,N_27543,N_26887);
xnor U28722 (N_28722,N_27460,N_27281);
nor U28723 (N_28723,N_27577,N_26683);
nand U28724 (N_28724,N_26712,N_26559);
or U28725 (N_28725,N_27141,N_27290);
and U28726 (N_28726,N_27460,N_26494);
xor U28727 (N_28727,N_27082,N_27555);
nand U28728 (N_28728,N_26651,N_26609);
xor U28729 (N_28729,N_27473,N_27511);
xnor U28730 (N_28730,N_26403,N_27007);
and U28731 (N_28731,N_27506,N_27462);
or U28732 (N_28732,N_26729,N_26539);
nand U28733 (N_28733,N_26801,N_27000);
nor U28734 (N_28734,N_27452,N_26425);
or U28735 (N_28735,N_26759,N_27520);
or U28736 (N_28736,N_27283,N_26409);
nor U28737 (N_28737,N_26592,N_27385);
nand U28738 (N_28738,N_26536,N_26624);
and U28739 (N_28739,N_27045,N_26914);
nor U28740 (N_28740,N_26934,N_26865);
nor U28741 (N_28741,N_27044,N_26758);
nand U28742 (N_28742,N_26408,N_26697);
or U28743 (N_28743,N_27111,N_26549);
xor U28744 (N_28744,N_26866,N_26434);
xor U28745 (N_28745,N_27071,N_26684);
and U28746 (N_28746,N_26518,N_26957);
xnor U28747 (N_28747,N_27331,N_27021);
nand U28748 (N_28748,N_27346,N_27513);
xnor U28749 (N_28749,N_27129,N_26967);
or U28750 (N_28750,N_27161,N_27164);
xor U28751 (N_28751,N_27137,N_26536);
and U28752 (N_28752,N_27470,N_27467);
xor U28753 (N_28753,N_26835,N_27183);
nor U28754 (N_28754,N_27494,N_27296);
and U28755 (N_28755,N_27420,N_26904);
and U28756 (N_28756,N_26743,N_27576);
and U28757 (N_28757,N_26594,N_26520);
or U28758 (N_28758,N_26567,N_27262);
nor U28759 (N_28759,N_26882,N_27315);
xnor U28760 (N_28760,N_26826,N_26444);
nand U28761 (N_28761,N_27169,N_26776);
nor U28762 (N_28762,N_26824,N_27393);
and U28763 (N_28763,N_27008,N_26576);
and U28764 (N_28764,N_26779,N_27070);
xor U28765 (N_28765,N_26441,N_26420);
or U28766 (N_28766,N_26418,N_26532);
nand U28767 (N_28767,N_26779,N_26744);
xor U28768 (N_28768,N_27422,N_27334);
nor U28769 (N_28769,N_26806,N_27086);
or U28770 (N_28770,N_27579,N_27216);
xor U28771 (N_28771,N_26428,N_26988);
and U28772 (N_28772,N_26463,N_27269);
nand U28773 (N_28773,N_26436,N_26648);
nand U28774 (N_28774,N_27167,N_27426);
or U28775 (N_28775,N_27440,N_27186);
xnor U28776 (N_28776,N_26991,N_26682);
and U28777 (N_28777,N_27450,N_26643);
nand U28778 (N_28778,N_26856,N_26814);
or U28779 (N_28779,N_27475,N_27476);
or U28780 (N_28780,N_27001,N_27003);
nor U28781 (N_28781,N_27369,N_27325);
or U28782 (N_28782,N_26874,N_27488);
nand U28783 (N_28783,N_26533,N_26431);
xnor U28784 (N_28784,N_27106,N_27584);
xor U28785 (N_28785,N_27382,N_26498);
and U28786 (N_28786,N_27090,N_26993);
and U28787 (N_28787,N_26650,N_26957);
and U28788 (N_28788,N_27425,N_26751);
xnor U28789 (N_28789,N_26834,N_26488);
nor U28790 (N_28790,N_26958,N_26431);
and U28791 (N_28791,N_27514,N_27091);
nand U28792 (N_28792,N_26978,N_27343);
or U28793 (N_28793,N_27510,N_27014);
nand U28794 (N_28794,N_26683,N_26956);
xnor U28795 (N_28795,N_26593,N_27525);
nand U28796 (N_28796,N_26645,N_26654);
and U28797 (N_28797,N_26974,N_26817);
nor U28798 (N_28798,N_26882,N_26755);
nand U28799 (N_28799,N_26735,N_26599);
nand U28800 (N_28800,N_28505,N_28547);
and U28801 (N_28801,N_27653,N_28630);
or U28802 (N_28802,N_28738,N_27781);
xnor U28803 (N_28803,N_28464,N_27835);
nand U28804 (N_28804,N_28302,N_27971);
nand U28805 (N_28805,N_28152,N_27896);
nand U28806 (N_28806,N_28461,N_28694);
and U28807 (N_28807,N_28089,N_28028);
nor U28808 (N_28808,N_28600,N_28787);
nor U28809 (N_28809,N_28478,N_28115);
nand U28810 (N_28810,N_27820,N_27759);
or U28811 (N_28811,N_28242,N_28445);
xnor U28812 (N_28812,N_28003,N_28327);
and U28813 (N_28813,N_28253,N_27868);
nand U28814 (N_28814,N_28382,N_28648);
nand U28815 (N_28815,N_27733,N_28351);
nand U28816 (N_28816,N_28013,N_28424);
xnor U28817 (N_28817,N_28365,N_28226);
nor U28818 (N_28818,N_28333,N_27834);
or U28819 (N_28819,N_28294,N_28356);
and U28820 (N_28820,N_27840,N_27703);
or U28821 (N_28821,N_28504,N_27916);
nor U28822 (N_28822,N_28580,N_28598);
or U28823 (N_28823,N_27708,N_28133);
or U28824 (N_28824,N_27743,N_27659);
or U28825 (N_28825,N_28128,N_28777);
nor U28826 (N_28826,N_28679,N_27687);
and U28827 (N_28827,N_28293,N_27706);
nand U28828 (N_28828,N_27692,N_28651);
or U28829 (N_28829,N_28716,N_28262);
nand U28830 (N_28830,N_28350,N_27824);
or U28831 (N_28831,N_27668,N_27787);
and U28832 (N_28832,N_28267,N_28565);
nor U28833 (N_28833,N_28397,N_27823);
nand U28834 (N_28834,N_28289,N_28779);
or U28835 (N_28835,N_27927,N_27673);
nand U28836 (N_28836,N_28724,N_28368);
nand U28837 (N_28837,N_27772,N_27911);
and U28838 (N_28838,N_28774,N_27764);
and U28839 (N_28839,N_28196,N_28221);
nor U28840 (N_28840,N_27860,N_27749);
or U28841 (N_28841,N_27757,N_28174);
nand U28842 (N_28842,N_28366,N_28576);
or U28843 (N_28843,N_28216,N_28195);
xor U28844 (N_28844,N_27890,N_28674);
or U28845 (N_28845,N_27917,N_27934);
and U28846 (N_28846,N_28538,N_28561);
and U28847 (N_28847,N_27893,N_28096);
nand U28848 (N_28848,N_28312,N_28307);
and U28849 (N_28849,N_27880,N_27650);
nand U28850 (N_28850,N_27850,N_28522);
nor U28851 (N_28851,N_28243,N_28258);
nor U28852 (N_28852,N_28180,N_28126);
nand U28853 (N_28853,N_28783,N_28415);
nand U28854 (N_28854,N_28446,N_28497);
and U28855 (N_28855,N_28410,N_28256);
and U28856 (N_28856,N_28029,N_28465);
nor U28857 (N_28857,N_27672,N_27995);
nand U28858 (N_28858,N_28392,N_27740);
or U28859 (N_28859,N_28755,N_28532);
xnor U28860 (N_28860,N_28427,N_28177);
or U28861 (N_28861,N_28662,N_28291);
and U28862 (N_28862,N_27907,N_27931);
nor U28863 (N_28863,N_28166,N_27935);
and U28864 (N_28864,N_28147,N_27973);
and U28865 (N_28865,N_27997,N_28124);
and U28866 (N_28866,N_27685,N_28157);
nor U28867 (N_28867,N_28117,N_27908);
nand U28868 (N_28868,N_28414,N_27679);
and U28869 (N_28869,N_28572,N_28438);
nor U28870 (N_28870,N_28406,N_27681);
and U28871 (N_28871,N_27807,N_27613);
or U28872 (N_28872,N_27878,N_28757);
or U28873 (N_28873,N_28090,N_27720);
xor U28874 (N_28874,N_27904,N_28223);
or U28875 (N_28875,N_27830,N_28103);
and U28876 (N_28876,N_27925,N_28364);
nand U28877 (N_28877,N_28190,N_27991);
nand U28878 (N_28878,N_28502,N_28635);
nor U28879 (N_28879,N_28586,N_28619);
nand U28880 (N_28880,N_28006,N_27951);
or U28881 (N_28881,N_27751,N_28620);
nor U28882 (N_28882,N_28151,N_28672);
or U28883 (N_28883,N_28788,N_28409);
nor U28884 (N_28884,N_27755,N_28769);
or U28885 (N_28885,N_28764,N_28313);
nand U28886 (N_28886,N_28765,N_28568);
and U28887 (N_28887,N_27667,N_28661);
nand U28888 (N_28888,N_28105,N_28563);
nor U28889 (N_28889,N_28112,N_27760);
and U28890 (N_28890,N_27622,N_27870);
nand U28891 (N_28891,N_27876,N_27848);
or U28892 (N_28892,N_27885,N_28012);
nor U28893 (N_28893,N_27956,N_28400);
xor U28894 (N_28894,N_28344,N_28439);
nor U28895 (N_28895,N_28039,N_27822);
and U28896 (N_28896,N_28069,N_27905);
xnor U28897 (N_28897,N_28376,N_27739);
or U28898 (N_28898,N_28317,N_28318);
nand U28899 (N_28899,N_27981,N_28125);
nand U28900 (N_28900,N_27637,N_27865);
and U28901 (N_28901,N_28271,N_28049);
or U28902 (N_28902,N_28078,N_28160);
nor U28903 (N_28903,N_28621,N_28129);
nand U28904 (N_28904,N_28573,N_28199);
and U28905 (N_28905,N_27621,N_28489);
or U28906 (N_28906,N_28099,N_28536);
and U28907 (N_28907,N_28466,N_28544);
or U28908 (N_28908,N_28791,N_28419);
nor U28909 (N_28909,N_27871,N_28211);
and U28910 (N_28910,N_28785,N_28746);
and U28911 (N_28911,N_28299,N_28136);
xor U28912 (N_28912,N_28132,N_28664);
or U28913 (N_28913,N_28653,N_28668);
and U28914 (N_28914,N_28706,N_27984);
and U28915 (N_28915,N_28388,N_28389);
nand U28916 (N_28916,N_28119,N_28411);
nor U28917 (N_28917,N_28331,N_27634);
or U28918 (N_28918,N_28754,N_27800);
and U28919 (N_28919,N_28176,N_28794);
nor U28920 (N_28920,N_28035,N_28690);
and U28921 (N_28921,N_27906,N_28405);
nor U28922 (N_28922,N_28259,N_27627);
nor U28923 (N_28923,N_28321,N_28705);
and U28924 (N_28924,N_28276,N_27922);
or U28925 (N_28925,N_28748,N_27736);
xnor U28926 (N_28926,N_28628,N_28760);
xor U28927 (N_28927,N_28562,N_27992);
nand U28928 (N_28928,N_28094,N_28110);
and U28929 (N_28929,N_28556,N_28245);
nor U28930 (N_28930,N_28220,N_28440);
nor U28931 (N_28931,N_28383,N_27811);
nand U28932 (N_28932,N_27620,N_27709);
and U28933 (N_28933,N_27888,N_27980);
or U28934 (N_28934,N_28062,N_28075);
or U28935 (N_28935,N_28676,N_28283);
and U28936 (N_28936,N_28772,N_28091);
or U28937 (N_28937,N_27617,N_27698);
nor U28938 (N_28938,N_28338,N_27901);
xnor U28939 (N_28939,N_28444,N_28675);
nor U28940 (N_28940,N_28191,N_28542);
nand U28941 (N_28941,N_28369,N_28009);
nor U28942 (N_28942,N_28182,N_28287);
or U28943 (N_28943,N_28083,N_27633);
nand U28944 (N_28944,N_27797,N_28740);
nor U28945 (N_28945,N_28448,N_27854);
and U28946 (N_28946,N_28387,N_27766);
or U28947 (N_28947,N_27898,N_28689);
and U28948 (N_28948,N_27961,N_28325);
nor U28949 (N_28949,N_28683,N_28487);
xnor U28950 (N_28950,N_28493,N_28343);
nand U28951 (N_28951,N_27604,N_28541);
nor U28952 (N_28952,N_27891,N_28380);
and U28953 (N_28953,N_28064,N_28044);
or U28954 (N_28954,N_28107,N_28145);
xnor U28955 (N_28955,N_27831,N_28719);
xnor U28956 (N_28956,N_27623,N_28530);
or U28957 (N_28957,N_28797,N_28649);
nand U28958 (N_28958,N_27929,N_28247);
and U28959 (N_28959,N_28559,N_28534);
xnor U28960 (N_28960,N_27808,N_28314);
or U28961 (N_28961,N_27689,N_28637);
nor U28962 (N_28962,N_28763,N_27962);
or U28963 (N_28963,N_28452,N_28781);
nor U28964 (N_28964,N_27939,N_28474);
xor U28965 (N_28965,N_28052,N_28703);
xnor U28966 (N_28966,N_28412,N_27600);
xor U28967 (N_28967,N_28713,N_28591);
xnor U28968 (N_28968,N_27690,N_28730);
or U28969 (N_28969,N_28686,N_27899);
xnor U28970 (N_28970,N_28347,N_28458);
nor U28971 (N_28971,N_27982,N_28552);
and U28972 (N_28972,N_28656,N_28775);
xor U28973 (N_28973,N_28531,N_28490);
or U28974 (N_28974,N_28193,N_28071);
nand U28975 (N_28975,N_28610,N_27863);
xor U28976 (N_28976,N_27978,N_28034);
nand U28977 (N_28977,N_28222,N_27866);
or U28978 (N_28978,N_28139,N_28639);
or U28979 (N_28979,N_28334,N_27853);
nor U28980 (N_28980,N_28155,N_27771);
nor U28981 (N_28981,N_28025,N_28214);
xor U28982 (N_28982,N_27928,N_28286);
xnor U28983 (N_28983,N_28413,N_27955);
xor U28984 (N_28984,N_28026,N_28123);
or U28985 (N_28985,N_28798,N_28575);
and U28986 (N_28986,N_27846,N_27624);
xor U28987 (N_28987,N_28043,N_28279);
nand U28988 (N_28988,N_28352,N_28607);
and U28989 (N_28989,N_28646,N_27785);
and U28990 (N_28990,N_27809,N_28260);
nor U28991 (N_28991,N_28718,N_27915);
and U28992 (N_28992,N_27861,N_27729);
nor U28993 (N_28993,N_28605,N_28033);
or U28994 (N_28994,N_28304,N_28692);
xor U28995 (N_28995,N_28184,N_27847);
or U28996 (N_28996,N_28254,N_28500);
xor U28997 (N_28997,N_28642,N_28138);
or U28998 (N_28998,N_28345,N_27684);
and U28999 (N_28999,N_27676,N_28583);
and U29000 (N_29000,N_27645,N_28205);
or U29001 (N_29001,N_27782,N_27651);
nand U29002 (N_29002,N_27776,N_28192);
nor U29003 (N_29003,N_28167,N_27680);
and U29004 (N_29004,N_28460,N_28697);
or U29005 (N_29005,N_28215,N_27874);
or U29006 (N_29006,N_28077,N_27707);
or U29007 (N_29007,N_28002,N_28015);
nor U29008 (N_29008,N_27762,N_27943);
nor U29009 (N_29009,N_28523,N_28643);
xnor U29010 (N_29010,N_28442,N_28000);
and U29011 (N_29011,N_28582,N_27819);
xnor U29012 (N_29012,N_28564,N_28353);
nand U29013 (N_29013,N_28153,N_28178);
xnor U29014 (N_29014,N_28525,N_28599);
nand U29015 (N_29015,N_28782,N_28189);
or U29016 (N_29016,N_28161,N_27608);
nand U29017 (N_29017,N_28244,N_28611);
xnor U29018 (N_29018,N_27833,N_27926);
xor U29019 (N_29019,N_27881,N_28421);
nor U29020 (N_29020,N_28756,N_27695);
nor U29021 (N_29021,N_28722,N_27769);
or U29022 (N_29022,N_27836,N_27789);
and U29023 (N_29023,N_28473,N_27867);
or U29024 (N_29024,N_27738,N_28209);
xor U29025 (N_29025,N_28162,N_28357);
xnor U29026 (N_29026,N_28527,N_28073);
or U29027 (N_29027,N_28156,N_27758);
xnor U29028 (N_29028,N_27849,N_27859);
nand U29029 (N_29029,N_28456,N_28081);
or U29030 (N_29030,N_27938,N_28758);
nor U29031 (N_29031,N_27986,N_28394);
and U29032 (N_29032,N_28227,N_28492);
or U29033 (N_29033,N_28308,N_27662);
nor U29034 (N_29034,N_28434,N_27711);
nor U29035 (N_29035,N_28305,N_27998);
nor U29036 (N_29036,N_28736,N_27775);
nor U29037 (N_29037,N_27948,N_27941);
and U29038 (N_29038,N_27828,N_28766);
or U29039 (N_29039,N_28455,N_27696);
xnor U29040 (N_29040,N_28375,N_27697);
nand U29041 (N_29041,N_27748,N_27829);
nand U29042 (N_29042,N_28249,N_27952);
or U29043 (N_29043,N_28018,N_27994);
or U29044 (N_29044,N_27855,N_28097);
and U29045 (N_29045,N_27747,N_28631);
xor U29046 (N_29046,N_28059,N_27875);
or U29047 (N_29047,N_28263,N_27644);
nand U29048 (N_29048,N_28606,N_28274);
nor U29049 (N_29049,N_27727,N_28390);
nand U29050 (N_29050,N_27784,N_28471);
and U29051 (N_29051,N_28589,N_28592);
nor U29052 (N_29052,N_28560,N_28799);
xor U29053 (N_29053,N_28200,N_27841);
nand U29054 (N_29054,N_27805,N_28596);
and U29055 (N_29055,N_28217,N_28399);
or U29056 (N_29056,N_28319,N_28720);
nand U29057 (N_29057,N_27942,N_28609);
nor U29058 (N_29058,N_27910,N_28503);
or U29059 (N_29059,N_28443,N_27741);
xnor U29060 (N_29060,N_28688,N_27832);
nand U29061 (N_29061,N_27856,N_28159);
or U29062 (N_29062,N_27826,N_27605);
nor U29063 (N_29063,N_28617,N_28238);
nor U29064 (N_29064,N_27798,N_28007);
or U29065 (N_29065,N_28601,N_28031);
xor U29066 (N_29066,N_28173,N_28426);
and U29067 (N_29067,N_27806,N_27777);
nand U29068 (N_29068,N_27852,N_28252);
or U29069 (N_29069,N_27753,N_28204);
xor U29070 (N_29070,N_28535,N_28048);
and U29071 (N_29071,N_27628,N_27933);
or U29072 (N_29072,N_28185,N_27658);
nor U29073 (N_29073,N_27641,N_28771);
and U29074 (N_29074,N_28201,N_28727);
and U29075 (N_29075,N_27682,N_27654);
and U29076 (N_29076,N_28257,N_27730);
and U29077 (N_29077,N_27958,N_28528);
nor U29078 (N_29078,N_28644,N_28454);
nor U29079 (N_29079,N_28498,N_28301);
xor U29080 (N_29080,N_28717,N_28225);
and U29081 (N_29081,N_27843,N_27718);
nor U29082 (N_29082,N_28432,N_28374);
nor U29083 (N_29083,N_28168,N_27635);
or U29084 (N_29084,N_28494,N_27724);
xor U29085 (N_29085,N_28587,N_28425);
and U29086 (N_29086,N_27655,N_28793);
nand U29087 (N_29087,N_28197,N_28100);
or U29088 (N_29088,N_28054,N_27990);
or U29089 (N_29089,N_27701,N_28051);
xor U29090 (N_29090,N_27677,N_28549);
nor U29091 (N_29091,N_28303,N_28170);
or U29092 (N_29092,N_27702,N_27970);
and U29093 (N_29093,N_28430,N_28558);
xor U29094 (N_29094,N_28417,N_28768);
nor U29095 (N_29095,N_27606,N_28261);
and U29096 (N_29096,N_28708,N_28543);
nand U29097 (N_29097,N_27774,N_28594);
nand U29098 (N_29098,N_28285,N_28017);
and U29099 (N_29099,N_28418,N_28508);
and U29100 (N_29100,N_27746,N_28459);
nand U29101 (N_29101,N_27723,N_28248);
nor U29102 (N_29102,N_27919,N_28087);
xnor U29103 (N_29103,N_27979,N_27669);
or U29104 (N_29104,N_28457,N_28593);
and U29105 (N_29105,N_28737,N_27872);
or U29106 (N_29106,N_28084,N_28614);
xor U29107 (N_29107,N_28761,N_28602);
nand U29108 (N_29108,N_28297,N_28691);
xnor U29109 (N_29109,N_28513,N_27814);
xor U29110 (N_29110,N_28346,N_28624);
nor U29111 (N_29111,N_28194,N_27683);
xnor U29112 (N_29112,N_28208,N_27710);
nand U29113 (N_29113,N_28336,N_28358);
or U29114 (N_29114,N_28067,N_28171);
and U29115 (N_29115,N_28010,N_28056);
and U29116 (N_29116,N_28349,N_27914);
nand U29117 (N_29117,N_28362,N_28086);
xor U29118 (N_29118,N_28379,N_27857);
and U29119 (N_29119,N_28751,N_28695);
nor U29120 (N_29120,N_28612,N_28577);
xnor U29121 (N_29121,N_27884,N_28550);
xor U29122 (N_29122,N_28516,N_27946);
or U29123 (N_29123,N_28235,N_28265);
or U29124 (N_29124,N_27873,N_28554);
and U29125 (N_29125,N_28407,N_27794);
or U29126 (N_29126,N_27629,N_28792);
xor U29127 (N_29127,N_28330,N_27618);
nor U29128 (N_29128,N_27968,N_27699);
xnor U29129 (N_29129,N_28468,N_28704);
nand U29130 (N_29130,N_27799,N_28743);
nor U29131 (N_29131,N_28423,N_27949);
and U29132 (N_29132,N_28210,N_28158);
and U29133 (N_29133,N_28436,N_27993);
nor U29134 (N_29134,N_28712,N_28450);
and U29135 (N_29135,N_27879,N_27900);
nand U29136 (N_29136,N_28645,N_28507);
and U29137 (N_29137,N_28753,N_28290);
xor U29138 (N_29138,N_28739,N_27964);
or U29139 (N_29139,N_27902,N_28680);
xnor U29140 (N_29140,N_28469,N_28711);
and U29141 (N_29141,N_28036,N_28479);
and U29142 (N_29142,N_28481,N_27924);
or U29143 (N_29143,N_28747,N_27999);
or U29144 (N_29144,N_27851,N_27607);
and U29145 (N_29145,N_28234,N_28732);
or U29146 (N_29146,N_28266,N_27649);
and U29147 (N_29147,N_27754,N_27639);
and U29148 (N_29148,N_28485,N_28641);
and U29149 (N_29149,N_27788,N_28361);
xnor U29150 (N_29150,N_28574,N_28323);
and U29151 (N_29151,N_28186,N_28332);
xnor U29152 (N_29152,N_28790,N_28623);
xor U29153 (N_29153,N_27657,N_28172);
nor U29154 (N_29154,N_28268,N_28693);
or U29155 (N_29155,N_28627,N_28187);
xor U29156 (N_29156,N_28367,N_27609);
nand U29157 (N_29157,N_27947,N_27715);
and U29158 (N_29158,N_28433,N_27612);
nand U29159 (N_29159,N_28475,N_28696);
nor U29160 (N_29160,N_27671,N_28275);
nor U29161 (N_29161,N_27967,N_27603);
or U29162 (N_29162,N_28510,N_28288);
nand U29163 (N_29163,N_28633,N_28578);
nor U29164 (N_29164,N_28373,N_27909);
and U29165 (N_29165,N_28058,N_28429);
nor U29166 (N_29166,N_28678,N_28109);
or U29167 (N_29167,N_27957,N_28306);
or U29168 (N_29168,N_28219,N_28618);
xnor U29169 (N_29169,N_27803,N_28684);
nand U29170 (N_29170,N_27678,N_28038);
nor U29171 (N_29171,N_28328,N_27988);
nor U29172 (N_29172,N_28041,N_28472);
xnor U29173 (N_29173,N_27818,N_28229);
xnor U29174 (N_29174,N_27717,N_28169);
nand U29175 (N_29175,N_28045,N_28340);
xor U29176 (N_29176,N_28435,N_27940);
nand U29177 (N_29177,N_28278,N_27773);
and U29178 (N_29178,N_28453,N_27742);
nand U29179 (N_29179,N_27725,N_28309);
or U29180 (N_29180,N_27732,N_28557);
and U29181 (N_29181,N_28773,N_28240);
and U29182 (N_29182,N_28707,N_28470);
xor U29183 (N_29183,N_28506,N_27937);
nor U29184 (N_29184,N_28251,N_27792);
or U29185 (N_29185,N_28311,N_27691);
nor U29186 (N_29186,N_28114,N_28681);
xnor U29187 (N_29187,N_28236,N_28329);
nor U29188 (N_29188,N_27768,N_28008);
xor U29189 (N_29189,N_27625,N_28032);
nand U29190 (N_29190,N_27704,N_28207);
nand U29191 (N_29191,N_28422,N_28517);
nor U29192 (N_29192,N_28659,N_28188);
nand U29193 (N_29193,N_28246,N_27661);
or U29194 (N_29194,N_27821,N_28514);
and U29195 (N_29195,N_27960,N_28230);
xnor U29196 (N_29196,N_27844,N_28698);
nand U29197 (N_29197,N_27883,N_28480);
and U29198 (N_29198,N_28298,N_27705);
nand U29199 (N_29199,N_28181,N_28237);
nand U29200 (N_29200,N_27770,N_28142);
or U29201 (N_29201,N_28408,N_28141);
xnor U29202 (N_29202,N_28685,N_28320);
and U29203 (N_29203,N_28284,N_28250);
or U29204 (N_29204,N_28626,N_27714);
nor U29205 (N_29205,N_28677,N_28673);
and U29206 (N_29206,N_28687,N_28163);
nand U29207 (N_29207,N_28515,N_28046);
and U29208 (N_29208,N_28377,N_28776);
and U29209 (N_29209,N_28604,N_28076);
nand U29210 (N_29210,N_27903,N_28721);
nor U29211 (N_29211,N_27974,N_28786);
nor U29212 (N_29212,N_27965,N_27780);
and U29213 (N_29213,N_28355,N_28057);
xor U29214 (N_29214,N_27675,N_27886);
or U29215 (N_29215,N_28540,N_27932);
and U29216 (N_29216,N_27894,N_28228);
xor U29217 (N_29217,N_28569,N_28735);
and U29218 (N_29218,N_27642,N_27745);
nor U29219 (N_29219,N_28654,N_27839);
nor U29220 (N_29220,N_28616,N_28005);
xor U29221 (N_29221,N_28122,N_28518);
and U29222 (N_29222,N_27666,N_28016);
xor U29223 (N_29223,N_28079,N_28710);
nand U29224 (N_29224,N_27663,N_28482);
nand U29225 (N_29225,N_28665,N_28566);
and U29226 (N_29226,N_27801,N_28037);
xor U29227 (N_29227,N_28613,N_28486);
and U29228 (N_29228,N_28396,N_28337);
and U29229 (N_29229,N_27977,N_28270);
or U29230 (N_29230,N_28121,N_28496);
or U29231 (N_29231,N_28526,N_27616);
or U29232 (N_29232,N_28416,N_27779);
nand U29233 (N_29233,N_28636,N_27923);
or U29234 (N_29234,N_28092,N_28512);
nand U29235 (N_29235,N_28371,N_28233);
and U29236 (N_29236,N_28767,N_28324);
nor U29237 (N_29237,N_27793,N_28019);
nor U29238 (N_29238,N_28657,N_27640);
or U29239 (N_29239,N_27626,N_28060);
nor U29240 (N_29240,N_27631,N_27636);
or U29241 (N_29241,N_28590,N_28632);
nor U29242 (N_29242,N_27877,N_28101);
or U29243 (N_29243,N_28402,N_28795);
or U29244 (N_29244,N_28011,N_28175);
nand U29245 (N_29245,N_28137,N_27945);
or U29246 (N_29246,N_28666,N_28702);
and U29247 (N_29247,N_28539,N_28529);
and U29248 (N_29248,N_28477,N_28488);
and U29249 (N_29249,N_27987,N_27638);
xnor U29250 (N_29250,N_28491,N_28239);
nand U29251 (N_29251,N_28206,N_28022);
nor U29252 (N_29252,N_28608,N_27944);
xor U29253 (N_29253,N_27744,N_27795);
and U29254 (N_29254,N_27750,N_28341);
and U29255 (N_29255,N_28729,N_28629);
nor U29256 (N_29256,N_28749,N_27752);
and U29257 (N_29257,N_28537,N_28570);
nor U29258 (N_29258,N_27756,N_28074);
and U29259 (N_29259,N_28533,N_28131);
nand U29260 (N_29260,N_28752,N_27765);
xor U29261 (N_29261,N_27869,N_28447);
nor U29262 (N_29262,N_28555,N_28140);
and U29263 (N_29263,N_28551,N_28495);
and U29264 (N_29264,N_28118,N_27632);
xnor U29265 (N_29265,N_28398,N_28296);
and U29266 (N_29266,N_27619,N_27670);
nor U29267 (N_29267,N_28682,N_28667);
xor U29268 (N_29268,N_27665,N_27812);
and U29269 (N_29269,N_27686,N_28431);
xor U29270 (N_29270,N_28203,N_27716);
nand U29271 (N_29271,N_28106,N_27726);
and U29272 (N_29272,N_28581,N_28733);
nor U29273 (N_29273,N_28709,N_27786);
nor U29274 (N_29274,N_27763,N_28269);
nor U29275 (N_29275,N_28295,N_28650);
xor U29276 (N_29276,N_28784,N_27989);
nor U29277 (N_29277,N_27862,N_27817);
xor U29278 (N_29278,N_27660,N_28483);
and U29279 (N_29279,N_27647,N_28640);
nand U29280 (N_29280,N_27950,N_27913);
or U29281 (N_29281,N_27737,N_27731);
nor U29282 (N_29282,N_28545,N_28378);
and U29283 (N_29283,N_28053,N_28403);
nand U29284 (N_29284,N_28381,N_28622);
xnor U29285 (N_29285,N_28030,N_28437);
nand U29286 (N_29286,N_28714,N_28047);
or U29287 (N_29287,N_28770,N_28744);
and U29288 (N_29288,N_28134,N_28386);
nor U29289 (N_29289,N_28104,N_27897);
and U29290 (N_29290,N_28521,N_28088);
nor U29291 (N_29291,N_28135,N_28055);
xor U29292 (N_29292,N_28042,N_28660);
nand U29293 (N_29293,N_28070,N_27796);
nand U29294 (N_29294,N_28360,N_28553);
and U29295 (N_29295,N_27953,N_28342);
and U29296 (N_29296,N_27827,N_28462);
or U29297 (N_29297,N_27721,N_28441);
xor U29298 (N_29298,N_27611,N_28241);
or U29299 (N_29299,N_27996,N_27966);
or U29300 (N_29300,N_28164,N_27674);
or U29301 (N_29301,N_28699,N_27802);
nor U29302 (N_29302,N_28428,N_28584);
nor U29303 (N_29303,N_27652,N_28255);
xor U29304 (N_29304,N_27845,N_28102);
xnor U29305 (N_29305,N_28120,N_28264);
or U29306 (N_29306,N_27778,N_27610);
nand U29307 (N_29307,N_27889,N_28728);
nand U29308 (N_29308,N_28232,N_27804);
nor U29309 (N_29309,N_28499,N_27972);
nand U29310 (N_29310,N_28395,N_27864);
nand U29311 (N_29311,N_28647,N_28014);
nor U29312 (N_29312,N_27921,N_28050);
nand U29313 (N_29313,N_28401,N_28218);
and U29314 (N_29314,N_28310,N_27954);
or U29315 (N_29315,N_28780,N_28146);
xor U29316 (N_29316,N_27664,N_28082);
xor U29317 (N_29317,N_28280,N_28315);
nand U29318 (N_29318,N_27646,N_28509);
nor U29319 (N_29319,N_27918,N_27892);
nor U29320 (N_29320,N_27630,N_27936);
and U29321 (N_29321,N_28597,N_27761);
xor U29322 (N_29322,N_27783,N_28595);
nand U29323 (N_29323,N_27656,N_27734);
and U29324 (N_29324,N_28655,N_27688);
nand U29325 (N_29325,N_28080,N_28085);
nor U29326 (N_29326,N_28322,N_28700);
nand U29327 (N_29327,N_28198,N_28404);
nor U29328 (N_29328,N_28212,N_27816);
nand U29329 (N_29329,N_28476,N_28548);
nor U29330 (N_29330,N_28148,N_27813);
nor U29331 (N_29331,N_27825,N_27694);
and U29332 (N_29332,N_28634,N_27791);
xnor U29333 (N_29333,N_28484,N_27643);
or U29334 (N_29334,N_27614,N_28670);
or U29335 (N_29335,N_28023,N_28282);
and U29336 (N_29336,N_27735,N_27887);
or U29337 (N_29337,N_28734,N_27963);
xor U29338 (N_29338,N_27882,N_28385);
nand U29339 (N_29339,N_27648,N_28359);
nand U29340 (N_29340,N_28546,N_27858);
or U29341 (N_29341,N_28715,N_27722);
or U29342 (N_29342,N_28393,N_28669);
nand U29343 (N_29343,N_27601,N_27983);
nand U29344 (N_29344,N_27713,N_28281);
or U29345 (N_29345,N_28027,N_28063);
xor U29346 (N_29346,N_28567,N_28093);
or U29347 (N_29347,N_28143,N_27700);
nand U29348 (N_29348,N_28762,N_28759);
or U29349 (N_29349,N_28796,N_28272);
and U29350 (N_29350,N_27842,N_28149);
or U29351 (N_29351,N_28348,N_28384);
xnor U29352 (N_29352,N_28001,N_28391);
nor U29353 (N_29353,N_27959,N_28130);
nor U29354 (N_29354,N_28335,N_27712);
and U29355 (N_29355,N_28098,N_28095);
xor U29356 (N_29356,N_28588,N_28066);
nor U29357 (N_29357,N_28004,N_27969);
and U29358 (N_29358,N_27790,N_28020);
and U29359 (N_29359,N_28778,N_28021);
nor U29360 (N_29360,N_28467,N_28511);
nor U29361 (N_29361,N_28370,N_28520);
xor U29362 (N_29362,N_28524,N_28108);
nand U29363 (N_29363,N_28316,N_28231);
xnor U29364 (N_29364,N_27728,N_28671);
nor U29365 (N_29365,N_28463,N_28065);
or U29366 (N_29366,N_28701,N_28113);
and U29367 (N_29367,N_28726,N_27976);
nor U29368 (N_29368,N_28061,N_27920);
or U29369 (N_29369,N_28585,N_27602);
or U29370 (N_29370,N_28354,N_28731);
nand U29371 (N_29371,N_28451,N_28277);
xor U29372 (N_29372,N_28741,N_28638);
xor U29373 (N_29373,N_28040,N_27985);
and U29374 (N_29374,N_28449,N_28024);
and U29375 (N_29375,N_28625,N_28116);
xnor U29376 (N_29376,N_28420,N_27810);
and U29377 (N_29377,N_28658,N_28750);
xnor U29378 (N_29378,N_28292,N_28144);
nor U29379 (N_29379,N_27912,N_28789);
xnor U29380 (N_29380,N_28111,N_28224);
nand U29381 (N_29381,N_27838,N_28501);
or U29382 (N_29382,N_28127,N_28723);
xor U29383 (N_29383,N_28579,N_27767);
nor U29384 (N_29384,N_28652,N_28519);
or U29385 (N_29385,N_28154,N_28150);
xnor U29386 (N_29386,N_28603,N_27895);
nand U29387 (N_29387,N_28663,N_28179);
and U29388 (N_29388,N_27975,N_28068);
or U29389 (N_29389,N_28165,N_28072);
nor U29390 (N_29390,N_28571,N_27837);
and U29391 (N_29391,N_28183,N_28615);
nand U29392 (N_29392,N_27719,N_28372);
nand U29393 (N_29393,N_28326,N_28745);
xor U29394 (N_29394,N_28363,N_27693);
xnor U29395 (N_29395,N_28742,N_27615);
or U29396 (N_29396,N_28273,N_27930);
nor U29397 (N_29397,N_28202,N_28725);
xnor U29398 (N_29398,N_28300,N_27815);
nand U29399 (N_29399,N_28339,N_28213);
and U29400 (N_29400,N_28178,N_28536);
xor U29401 (N_29401,N_28536,N_27929);
nand U29402 (N_29402,N_28428,N_27711);
nand U29403 (N_29403,N_28513,N_28132);
and U29404 (N_29404,N_28157,N_27954);
xnor U29405 (N_29405,N_28397,N_27737);
or U29406 (N_29406,N_27939,N_28231);
nor U29407 (N_29407,N_27722,N_28547);
nor U29408 (N_29408,N_28685,N_28660);
or U29409 (N_29409,N_28770,N_27975);
nand U29410 (N_29410,N_28065,N_28167);
xnor U29411 (N_29411,N_28339,N_28016);
and U29412 (N_29412,N_27686,N_27754);
or U29413 (N_29413,N_27707,N_27965);
nor U29414 (N_29414,N_28436,N_27911);
nor U29415 (N_29415,N_28760,N_28599);
nand U29416 (N_29416,N_27791,N_28069);
nand U29417 (N_29417,N_27632,N_28338);
nand U29418 (N_29418,N_28012,N_27745);
nor U29419 (N_29419,N_28554,N_27882);
nand U29420 (N_29420,N_28626,N_27644);
and U29421 (N_29421,N_27829,N_28368);
nor U29422 (N_29422,N_28651,N_27882);
or U29423 (N_29423,N_27724,N_28689);
and U29424 (N_29424,N_28120,N_27643);
nor U29425 (N_29425,N_28383,N_28111);
or U29426 (N_29426,N_27612,N_28005);
nor U29427 (N_29427,N_28574,N_28380);
and U29428 (N_29428,N_27986,N_28367);
and U29429 (N_29429,N_28480,N_28745);
nand U29430 (N_29430,N_27877,N_28421);
and U29431 (N_29431,N_27733,N_28163);
and U29432 (N_29432,N_28314,N_28396);
and U29433 (N_29433,N_28458,N_28183);
and U29434 (N_29434,N_28470,N_28682);
nand U29435 (N_29435,N_28055,N_27652);
or U29436 (N_29436,N_28548,N_28096);
xnor U29437 (N_29437,N_27666,N_27659);
nor U29438 (N_29438,N_28498,N_28086);
nor U29439 (N_29439,N_28691,N_27968);
and U29440 (N_29440,N_28735,N_28154);
and U29441 (N_29441,N_28499,N_28368);
xnor U29442 (N_29442,N_27874,N_28151);
and U29443 (N_29443,N_28366,N_27615);
or U29444 (N_29444,N_28762,N_28534);
xor U29445 (N_29445,N_28536,N_28151);
xnor U29446 (N_29446,N_27885,N_28160);
or U29447 (N_29447,N_28764,N_28258);
and U29448 (N_29448,N_28449,N_28191);
or U29449 (N_29449,N_28547,N_28101);
and U29450 (N_29450,N_28662,N_27834);
and U29451 (N_29451,N_27783,N_28733);
xnor U29452 (N_29452,N_27815,N_27842);
nand U29453 (N_29453,N_28531,N_27853);
xnor U29454 (N_29454,N_28755,N_28307);
nor U29455 (N_29455,N_27602,N_27824);
nand U29456 (N_29456,N_28695,N_28717);
nor U29457 (N_29457,N_28736,N_28534);
nor U29458 (N_29458,N_28712,N_28769);
nand U29459 (N_29459,N_28403,N_28340);
xor U29460 (N_29460,N_28385,N_27927);
and U29461 (N_29461,N_28085,N_28426);
xor U29462 (N_29462,N_28761,N_28208);
and U29463 (N_29463,N_28354,N_27692);
and U29464 (N_29464,N_27808,N_28412);
or U29465 (N_29465,N_27984,N_27708);
nor U29466 (N_29466,N_28665,N_28764);
or U29467 (N_29467,N_28337,N_28399);
xnor U29468 (N_29468,N_27942,N_28700);
or U29469 (N_29469,N_28538,N_27687);
nand U29470 (N_29470,N_28059,N_28703);
xnor U29471 (N_29471,N_28121,N_28718);
or U29472 (N_29472,N_27810,N_27742);
xor U29473 (N_29473,N_28070,N_27659);
nand U29474 (N_29474,N_28759,N_27887);
xor U29475 (N_29475,N_28388,N_28739);
nand U29476 (N_29476,N_28721,N_28048);
xnor U29477 (N_29477,N_28107,N_28582);
or U29478 (N_29478,N_28327,N_27944);
and U29479 (N_29479,N_28779,N_27914);
nor U29480 (N_29480,N_28229,N_28480);
nor U29481 (N_29481,N_28728,N_28022);
or U29482 (N_29482,N_27832,N_28312);
or U29483 (N_29483,N_28079,N_28049);
nand U29484 (N_29484,N_28197,N_27826);
and U29485 (N_29485,N_27985,N_28297);
or U29486 (N_29486,N_27786,N_28518);
or U29487 (N_29487,N_28709,N_27773);
nor U29488 (N_29488,N_28165,N_28211);
nor U29489 (N_29489,N_28032,N_27846);
nand U29490 (N_29490,N_28699,N_28105);
and U29491 (N_29491,N_28648,N_28429);
nand U29492 (N_29492,N_28335,N_28242);
nand U29493 (N_29493,N_27846,N_28087);
and U29494 (N_29494,N_28607,N_27977);
and U29495 (N_29495,N_27936,N_28169);
and U29496 (N_29496,N_28361,N_27910);
xor U29497 (N_29497,N_28679,N_27709);
or U29498 (N_29498,N_27804,N_28263);
nor U29499 (N_29499,N_28516,N_28469);
xor U29500 (N_29500,N_28581,N_28732);
or U29501 (N_29501,N_28539,N_27810);
nor U29502 (N_29502,N_28424,N_27609);
nor U29503 (N_29503,N_27952,N_27734);
and U29504 (N_29504,N_27876,N_27652);
nor U29505 (N_29505,N_28130,N_28237);
nor U29506 (N_29506,N_28487,N_28621);
and U29507 (N_29507,N_27898,N_28667);
xor U29508 (N_29508,N_28291,N_27968);
nor U29509 (N_29509,N_28322,N_28794);
or U29510 (N_29510,N_28191,N_27831);
and U29511 (N_29511,N_28459,N_28134);
nor U29512 (N_29512,N_28101,N_27605);
and U29513 (N_29513,N_28099,N_28787);
xnor U29514 (N_29514,N_28326,N_28612);
xor U29515 (N_29515,N_28403,N_28319);
and U29516 (N_29516,N_28581,N_28528);
nor U29517 (N_29517,N_27960,N_28748);
or U29518 (N_29518,N_27828,N_27822);
xnor U29519 (N_29519,N_28223,N_27957);
or U29520 (N_29520,N_27947,N_27974);
or U29521 (N_29521,N_28111,N_27753);
nand U29522 (N_29522,N_28594,N_28470);
and U29523 (N_29523,N_27981,N_28022);
or U29524 (N_29524,N_27928,N_27944);
and U29525 (N_29525,N_28013,N_27917);
nor U29526 (N_29526,N_27761,N_27654);
and U29527 (N_29527,N_27622,N_28548);
nor U29528 (N_29528,N_28783,N_28534);
nand U29529 (N_29529,N_27953,N_27629);
nor U29530 (N_29530,N_28553,N_27733);
xor U29531 (N_29531,N_27977,N_27781);
or U29532 (N_29532,N_27846,N_27766);
xor U29533 (N_29533,N_28655,N_27860);
nor U29534 (N_29534,N_28503,N_28784);
and U29535 (N_29535,N_28313,N_28657);
and U29536 (N_29536,N_28384,N_28297);
nand U29537 (N_29537,N_28346,N_28317);
xor U29538 (N_29538,N_28394,N_28560);
and U29539 (N_29539,N_27900,N_27730);
or U29540 (N_29540,N_27709,N_27677);
xnor U29541 (N_29541,N_28623,N_27769);
and U29542 (N_29542,N_28679,N_28293);
nor U29543 (N_29543,N_28215,N_28545);
or U29544 (N_29544,N_27826,N_27768);
and U29545 (N_29545,N_28343,N_28183);
and U29546 (N_29546,N_27774,N_27959);
nand U29547 (N_29547,N_27816,N_28797);
or U29548 (N_29548,N_27968,N_28612);
and U29549 (N_29549,N_27976,N_27652);
or U29550 (N_29550,N_27932,N_27699);
and U29551 (N_29551,N_28564,N_27878);
nand U29552 (N_29552,N_27785,N_28773);
and U29553 (N_29553,N_27655,N_28643);
or U29554 (N_29554,N_28426,N_27619);
xor U29555 (N_29555,N_28502,N_28185);
nor U29556 (N_29556,N_28443,N_27963);
or U29557 (N_29557,N_28421,N_28706);
nor U29558 (N_29558,N_28663,N_28782);
nand U29559 (N_29559,N_27919,N_28118);
and U29560 (N_29560,N_27830,N_28619);
xor U29561 (N_29561,N_28790,N_28229);
nor U29562 (N_29562,N_28425,N_28504);
xnor U29563 (N_29563,N_28327,N_27905);
nand U29564 (N_29564,N_28228,N_27732);
xnor U29565 (N_29565,N_28716,N_28259);
nand U29566 (N_29566,N_27657,N_28288);
or U29567 (N_29567,N_27761,N_28245);
and U29568 (N_29568,N_27995,N_28393);
and U29569 (N_29569,N_28261,N_28600);
and U29570 (N_29570,N_28364,N_27612);
or U29571 (N_29571,N_27826,N_27843);
nor U29572 (N_29572,N_28082,N_28351);
xnor U29573 (N_29573,N_28731,N_27860);
nand U29574 (N_29574,N_28232,N_28636);
and U29575 (N_29575,N_28191,N_28528);
or U29576 (N_29576,N_28352,N_28393);
nor U29577 (N_29577,N_28621,N_28391);
and U29578 (N_29578,N_28645,N_28261);
nand U29579 (N_29579,N_27841,N_28337);
or U29580 (N_29580,N_28763,N_28597);
nand U29581 (N_29581,N_28175,N_28113);
nand U29582 (N_29582,N_27930,N_28503);
or U29583 (N_29583,N_28004,N_28610);
nand U29584 (N_29584,N_27632,N_28545);
and U29585 (N_29585,N_28156,N_28488);
nand U29586 (N_29586,N_28047,N_28130);
nor U29587 (N_29587,N_28614,N_27806);
and U29588 (N_29588,N_28173,N_27690);
nand U29589 (N_29589,N_27995,N_28195);
nand U29590 (N_29590,N_28439,N_28124);
and U29591 (N_29591,N_28402,N_27917);
or U29592 (N_29592,N_28625,N_27956);
nor U29593 (N_29593,N_28663,N_28495);
nor U29594 (N_29594,N_28656,N_28203);
xnor U29595 (N_29595,N_28751,N_28055);
and U29596 (N_29596,N_27602,N_27822);
and U29597 (N_29597,N_28031,N_27685);
or U29598 (N_29598,N_28204,N_27897);
or U29599 (N_29599,N_28501,N_27604);
or U29600 (N_29600,N_28286,N_28409);
and U29601 (N_29601,N_28370,N_27936);
nor U29602 (N_29602,N_28437,N_28584);
and U29603 (N_29603,N_28752,N_28053);
nand U29604 (N_29604,N_28130,N_28051);
or U29605 (N_29605,N_27715,N_28050);
and U29606 (N_29606,N_28266,N_28522);
nor U29607 (N_29607,N_28672,N_27668);
xnor U29608 (N_29608,N_27824,N_28198);
and U29609 (N_29609,N_28391,N_28422);
and U29610 (N_29610,N_28256,N_28335);
xnor U29611 (N_29611,N_28259,N_27736);
nand U29612 (N_29612,N_28728,N_28581);
xnor U29613 (N_29613,N_28397,N_27923);
xor U29614 (N_29614,N_28095,N_27860);
nor U29615 (N_29615,N_28168,N_27765);
or U29616 (N_29616,N_28125,N_28715);
xor U29617 (N_29617,N_28731,N_28582);
nor U29618 (N_29618,N_28353,N_28379);
and U29619 (N_29619,N_28717,N_27696);
nand U29620 (N_29620,N_28754,N_28110);
and U29621 (N_29621,N_28097,N_28201);
or U29622 (N_29622,N_28033,N_28601);
nand U29623 (N_29623,N_28421,N_28251);
nand U29624 (N_29624,N_27610,N_28051);
and U29625 (N_29625,N_27714,N_27920);
xnor U29626 (N_29626,N_27761,N_28375);
xor U29627 (N_29627,N_27843,N_27896);
xor U29628 (N_29628,N_28435,N_28543);
nand U29629 (N_29629,N_27825,N_27806);
or U29630 (N_29630,N_28194,N_28374);
nand U29631 (N_29631,N_27671,N_28502);
nor U29632 (N_29632,N_28109,N_28577);
nor U29633 (N_29633,N_27971,N_28735);
nand U29634 (N_29634,N_28158,N_28034);
nand U29635 (N_29635,N_28643,N_28453);
and U29636 (N_29636,N_28045,N_28589);
nand U29637 (N_29637,N_28730,N_28772);
and U29638 (N_29638,N_28475,N_28431);
and U29639 (N_29639,N_28373,N_27667);
xnor U29640 (N_29640,N_28427,N_28034);
xor U29641 (N_29641,N_28543,N_27835);
and U29642 (N_29642,N_28195,N_28059);
xnor U29643 (N_29643,N_28791,N_28706);
or U29644 (N_29644,N_27873,N_27816);
xnor U29645 (N_29645,N_28479,N_27878);
nand U29646 (N_29646,N_28248,N_28309);
nand U29647 (N_29647,N_27971,N_28782);
nor U29648 (N_29648,N_28520,N_28505);
nand U29649 (N_29649,N_28061,N_28439);
nand U29650 (N_29650,N_28157,N_28348);
and U29651 (N_29651,N_27781,N_28454);
xor U29652 (N_29652,N_28414,N_28035);
nor U29653 (N_29653,N_28458,N_28110);
and U29654 (N_29654,N_28287,N_27839);
xnor U29655 (N_29655,N_28393,N_28161);
nor U29656 (N_29656,N_28780,N_28601);
or U29657 (N_29657,N_28026,N_28691);
nor U29658 (N_29658,N_28097,N_28230);
and U29659 (N_29659,N_27624,N_28372);
nand U29660 (N_29660,N_27985,N_28783);
or U29661 (N_29661,N_27680,N_28383);
and U29662 (N_29662,N_27736,N_27862);
nand U29663 (N_29663,N_28234,N_27889);
nand U29664 (N_29664,N_28646,N_27790);
nand U29665 (N_29665,N_27674,N_28644);
and U29666 (N_29666,N_27980,N_28649);
nor U29667 (N_29667,N_28677,N_28312);
nand U29668 (N_29668,N_28180,N_27722);
xnor U29669 (N_29669,N_28237,N_28123);
nor U29670 (N_29670,N_28608,N_27919);
nor U29671 (N_29671,N_28271,N_28444);
or U29672 (N_29672,N_28408,N_28737);
xor U29673 (N_29673,N_28587,N_27890);
nand U29674 (N_29674,N_28580,N_27651);
nor U29675 (N_29675,N_28197,N_27662);
and U29676 (N_29676,N_27894,N_28067);
xor U29677 (N_29677,N_28720,N_27672);
or U29678 (N_29678,N_28694,N_28695);
nand U29679 (N_29679,N_28706,N_27952);
xnor U29680 (N_29680,N_27865,N_28017);
or U29681 (N_29681,N_27847,N_27927);
nand U29682 (N_29682,N_28081,N_27978);
nor U29683 (N_29683,N_28177,N_28566);
or U29684 (N_29684,N_28633,N_28789);
and U29685 (N_29685,N_27993,N_28097);
nor U29686 (N_29686,N_28181,N_27705);
and U29687 (N_29687,N_27706,N_28324);
and U29688 (N_29688,N_27938,N_28287);
or U29689 (N_29689,N_28747,N_27756);
and U29690 (N_29690,N_27630,N_27906);
xnor U29691 (N_29691,N_27899,N_27701);
and U29692 (N_29692,N_27633,N_28445);
xnor U29693 (N_29693,N_27697,N_28595);
nand U29694 (N_29694,N_28379,N_27808);
and U29695 (N_29695,N_28671,N_27936);
nor U29696 (N_29696,N_28183,N_27808);
nand U29697 (N_29697,N_28580,N_28134);
xnor U29698 (N_29698,N_27953,N_28749);
or U29699 (N_29699,N_27802,N_27811);
nand U29700 (N_29700,N_28190,N_28150);
and U29701 (N_29701,N_27738,N_28436);
or U29702 (N_29702,N_28597,N_28369);
and U29703 (N_29703,N_27795,N_28652);
xor U29704 (N_29704,N_28336,N_28137);
or U29705 (N_29705,N_28060,N_27700);
and U29706 (N_29706,N_27792,N_28034);
nor U29707 (N_29707,N_28173,N_28675);
nand U29708 (N_29708,N_27844,N_28560);
xnor U29709 (N_29709,N_28506,N_28323);
xor U29710 (N_29710,N_28464,N_28733);
and U29711 (N_29711,N_28590,N_28516);
xnor U29712 (N_29712,N_28098,N_27744);
nand U29713 (N_29713,N_28192,N_27764);
xor U29714 (N_29714,N_27834,N_28434);
and U29715 (N_29715,N_28734,N_27643);
xnor U29716 (N_29716,N_28346,N_28666);
nand U29717 (N_29717,N_28309,N_27958);
or U29718 (N_29718,N_28423,N_27887);
or U29719 (N_29719,N_28556,N_28740);
nand U29720 (N_29720,N_28618,N_28614);
and U29721 (N_29721,N_28539,N_28006);
nor U29722 (N_29722,N_27689,N_28596);
and U29723 (N_29723,N_27825,N_27975);
nand U29724 (N_29724,N_28028,N_28718);
or U29725 (N_29725,N_28182,N_28565);
nor U29726 (N_29726,N_28172,N_28298);
or U29727 (N_29727,N_27757,N_27716);
xnor U29728 (N_29728,N_28637,N_28652);
and U29729 (N_29729,N_27872,N_28101);
nor U29730 (N_29730,N_28195,N_28539);
nor U29731 (N_29731,N_27777,N_28059);
nor U29732 (N_29732,N_27977,N_27693);
and U29733 (N_29733,N_27880,N_28400);
nor U29734 (N_29734,N_28341,N_28095);
or U29735 (N_29735,N_28026,N_27679);
and U29736 (N_29736,N_27989,N_28294);
or U29737 (N_29737,N_28143,N_27885);
nand U29738 (N_29738,N_28081,N_27721);
xor U29739 (N_29739,N_28095,N_27630);
nor U29740 (N_29740,N_28786,N_27648);
nand U29741 (N_29741,N_27931,N_28285);
nor U29742 (N_29742,N_28551,N_27709);
and U29743 (N_29743,N_28387,N_28233);
or U29744 (N_29744,N_28216,N_28717);
xnor U29745 (N_29745,N_27918,N_28246);
and U29746 (N_29746,N_28652,N_28131);
nor U29747 (N_29747,N_27961,N_28138);
or U29748 (N_29748,N_28132,N_27649);
xnor U29749 (N_29749,N_27872,N_27624);
nand U29750 (N_29750,N_28374,N_28269);
or U29751 (N_29751,N_28339,N_27906);
xor U29752 (N_29752,N_28493,N_27967);
nand U29753 (N_29753,N_27893,N_27678);
and U29754 (N_29754,N_27742,N_27683);
or U29755 (N_29755,N_28156,N_27612);
and U29756 (N_29756,N_27819,N_27711);
and U29757 (N_29757,N_27942,N_28372);
or U29758 (N_29758,N_28233,N_28491);
xnor U29759 (N_29759,N_27940,N_27626);
nor U29760 (N_29760,N_27854,N_28781);
and U29761 (N_29761,N_28458,N_28506);
nand U29762 (N_29762,N_28298,N_27972);
and U29763 (N_29763,N_28044,N_28340);
and U29764 (N_29764,N_27792,N_27850);
nor U29765 (N_29765,N_28734,N_28132);
nor U29766 (N_29766,N_28473,N_28359);
nor U29767 (N_29767,N_27612,N_27777);
nor U29768 (N_29768,N_28612,N_28506);
nand U29769 (N_29769,N_28484,N_27783);
nand U29770 (N_29770,N_28272,N_27940);
nand U29771 (N_29771,N_27757,N_28764);
nor U29772 (N_29772,N_28129,N_28521);
nor U29773 (N_29773,N_28012,N_28356);
or U29774 (N_29774,N_28598,N_27943);
nor U29775 (N_29775,N_28654,N_27651);
nor U29776 (N_29776,N_28090,N_27754);
nor U29777 (N_29777,N_28496,N_27607);
or U29778 (N_29778,N_27851,N_27693);
and U29779 (N_29779,N_28189,N_27881);
nor U29780 (N_29780,N_27620,N_28570);
nand U29781 (N_29781,N_27618,N_27977);
nand U29782 (N_29782,N_28065,N_28731);
xnor U29783 (N_29783,N_28391,N_27936);
nor U29784 (N_29784,N_27976,N_27939);
nor U29785 (N_29785,N_28323,N_27975);
xnor U29786 (N_29786,N_28282,N_28776);
and U29787 (N_29787,N_28308,N_28417);
nand U29788 (N_29788,N_28509,N_28487);
and U29789 (N_29789,N_28686,N_28359);
nand U29790 (N_29790,N_28523,N_27619);
or U29791 (N_29791,N_27695,N_27860);
or U29792 (N_29792,N_27733,N_28079);
or U29793 (N_29793,N_28294,N_27666);
xor U29794 (N_29794,N_28777,N_27649);
xnor U29795 (N_29795,N_28781,N_27944);
or U29796 (N_29796,N_28219,N_28666);
nor U29797 (N_29797,N_27662,N_28520);
or U29798 (N_29798,N_28732,N_28682);
nor U29799 (N_29799,N_28603,N_28483);
or U29800 (N_29800,N_28386,N_28796);
xnor U29801 (N_29801,N_28394,N_28314);
and U29802 (N_29802,N_27690,N_28703);
or U29803 (N_29803,N_28543,N_27693);
and U29804 (N_29804,N_28250,N_28222);
or U29805 (N_29805,N_28509,N_27669);
and U29806 (N_29806,N_28353,N_28641);
and U29807 (N_29807,N_28227,N_28594);
and U29808 (N_29808,N_28737,N_28150);
xnor U29809 (N_29809,N_28010,N_27698);
nor U29810 (N_29810,N_28539,N_27943);
and U29811 (N_29811,N_27778,N_27857);
nor U29812 (N_29812,N_28327,N_27711);
nor U29813 (N_29813,N_28794,N_28770);
nand U29814 (N_29814,N_28599,N_27890);
nand U29815 (N_29815,N_28527,N_27792);
nor U29816 (N_29816,N_27854,N_27954);
nand U29817 (N_29817,N_27989,N_28449);
or U29818 (N_29818,N_28580,N_28384);
xor U29819 (N_29819,N_27771,N_27993);
nand U29820 (N_29820,N_28407,N_28647);
nand U29821 (N_29821,N_27755,N_28731);
nor U29822 (N_29822,N_28659,N_27749);
and U29823 (N_29823,N_28516,N_28445);
xor U29824 (N_29824,N_28134,N_28036);
nor U29825 (N_29825,N_28189,N_27726);
nand U29826 (N_29826,N_27634,N_27826);
nor U29827 (N_29827,N_28018,N_28221);
nor U29828 (N_29828,N_28276,N_28384);
and U29829 (N_29829,N_28570,N_28151);
and U29830 (N_29830,N_27813,N_27999);
or U29831 (N_29831,N_28583,N_28617);
and U29832 (N_29832,N_27925,N_27678);
and U29833 (N_29833,N_28106,N_28325);
nand U29834 (N_29834,N_28250,N_27711);
and U29835 (N_29835,N_28686,N_28774);
xor U29836 (N_29836,N_27906,N_28177);
and U29837 (N_29837,N_28374,N_28650);
nand U29838 (N_29838,N_28651,N_27854);
nand U29839 (N_29839,N_28082,N_28048);
nand U29840 (N_29840,N_28788,N_28285);
nand U29841 (N_29841,N_27930,N_28407);
nor U29842 (N_29842,N_28686,N_27867);
xnor U29843 (N_29843,N_27922,N_28305);
nor U29844 (N_29844,N_28770,N_28566);
and U29845 (N_29845,N_28772,N_28189);
nand U29846 (N_29846,N_28294,N_28340);
or U29847 (N_29847,N_27855,N_28576);
nor U29848 (N_29848,N_28111,N_28411);
xor U29849 (N_29849,N_28645,N_28569);
xnor U29850 (N_29850,N_28497,N_28711);
nor U29851 (N_29851,N_27947,N_27732);
nor U29852 (N_29852,N_28759,N_27648);
nand U29853 (N_29853,N_28752,N_28005);
and U29854 (N_29854,N_28111,N_28604);
or U29855 (N_29855,N_27684,N_27834);
or U29856 (N_29856,N_28726,N_28237);
and U29857 (N_29857,N_27640,N_28410);
and U29858 (N_29858,N_27878,N_27639);
and U29859 (N_29859,N_28016,N_28678);
nor U29860 (N_29860,N_28193,N_28680);
and U29861 (N_29861,N_28552,N_28493);
nor U29862 (N_29862,N_28391,N_27652);
nand U29863 (N_29863,N_28613,N_28775);
nand U29864 (N_29864,N_27813,N_27739);
or U29865 (N_29865,N_27859,N_28119);
and U29866 (N_29866,N_28199,N_28113);
nand U29867 (N_29867,N_27769,N_28148);
and U29868 (N_29868,N_28145,N_27768);
and U29869 (N_29869,N_28737,N_28362);
nand U29870 (N_29870,N_28075,N_27881);
xnor U29871 (N_29871,N_28459,N_28763);
and U29872 (N_29872,N_28718,N_28261);
nor U29873 (N_29873,N_27833,N_28219);
or U29874 (N_29874,N_28707,N_28416);
xor U29875 (N_29875,N_27809,N_28588);
and U29876 (N_29876,N_28182,N_28568);
and U29877 (N_29877,N_28617,N_27921);
nand U29878 (N_29878,N_28515,N_27863);
or U29879 (N_29879,N_28349,N_28152);
and U29880 (N_29880,N_28385,N_28522);
xnor U29881 (N_29881,N_27679,N_28145);
nand U29882 (N_29882,N_28531,N_27684);
or U29883 (N_29883,N_28302,N_28349);
or U29884 (N_29884,N_28408,N_27636);
nand U29885 (N_29885,N_28102,N_27965);
or U29886 (N_29886,N_28599,N_28139);
and U29887 (N_29887,N_28701,N_27896);
or U29888 (N_29888,N_27910,N_28737);
or U29889 (N_29889,N_28323,N_27877);
nand U29890 (N_29890,N_27621,N_27626);
and U29891 (N_29891,N_27617,N_28486);
nor U29892 (N_29892,N_28115,N_28364);
and U29893 (N_29893,N_27641,N_28239);
and U29894 (N_29894,N_28664,N_27808);
or U29895 (N_29895,N_27798,N_28226);
nand U29896 (N_29896,N_28514,N_27755);
nand U29897 (N_29897,N_27894,N_28158);
nand U29898 (N_29898,N_28278,N_28286);
and U29899 (N_29899,N_28169,N_28188);
xor U29900 (N_29900,N_28234,N_27731);
nor U29901 (N_29901,N_27935,N_27754);
nor U29902 (N_29902,N_27747,N_27978);
xnor U29903 (N_29903,N_28003,N_28168);
or U29904 (N_29904,N_27727,N_28455);
nor U29905 (N_29905,N_28359,N_28287);
and U29906 (N_29906,N_27705,N_28196);
and U29907 (N_29907,N_27633,N_28109);
or U29908 (N_29908,N_28008,N_27870);
xnor U29909 (N_29909,N_27906,N_28198);
nor U29910 (N_29910,N_27970,N_28752);
nand U29911 (N_29911,N_28382,N_28571);
or U29912 (N_29912,N_28764,N_28732);
nor U29913 (N_29913,N_28658,N_28243);
and U29914 (N_29914,N_27827,N_27800);
nand U29915 (N_29915,N_28140,N_27740);
nor U29916 (N_29916,N_28738,N_28189);
nand U29917 (N_29917,N_28289,N_28171);
xor U29918 (N_29918,N_28753,N_28379);
and U29919 (N_29919,N_27682,N_28385);
or U29920 (N_29920,N_28742,N_28288);
nor U29921 (N_29921,N_28505,N_28006);
or U29922 (N_29922,N_28147,N_27865);
and U29923 (N_29923,N_28782,N_28740);
xor U29924 (N_29924,N_28161,N_28174);
nor U29925 (N_29925,N_28599,N_28282);
nand U29926 (N_29926,N_27950,N_28181);
nor U29927 (N_29927,N_28565,N_28783);
or U29928 (N_29928,N_27939,N_28290);
nand U29929 (N_29929,N_28598,N_27918);
and U29930 (N_29930,N_28687,N_28136);
nand U29931 (N_29931,N_28501,N_28340);
or U29932 (N_29932,N_28060,N_27749);
and U29933 (N_29933,N_28166,N_28328);
nand U29934 (N_29934,N_28747,N_28067);
xnor U29935 (N_29935,N_28321,N_28213);
xor U29936 (N_29936,N_28096,N_28254);
nand U29937 (N_29937,N_28456,N_28249);
or U29938 (N_29938,N_28115,N_28321);
nand U29939 (N_29939,N_28448,N_28174);
and U29940 (N_29940,N_27871,N_28316);
nor U29941 (N_29941,N_27665,N_27656);
or U29942 (N_29942,N_28755,N_28219);
nand U29943 (N_29943,N_28079,N_28697);
or U29944 (N_29944,N_28267,N_28098);
or U29945 (N_29945,N_28036,N_28245);
or U29946 (N_29946,N_28626,N_28291);
or U29947 (N_29947,N_28517,N_28239);
xor U29948 (N_29948,N_28001,N_28294);
nor U29949 (N_29949,N_27740,N_28449);
nor U29950 (N_29950,N_27918,N_28334);
xor U29951 (N_29951,N_28054,N_27984);
nor U29952 (N_29952,N_28056,N_28421);
nor U29953 (N_29953,N_28743,N_28101);
xnor U29954 (N_29954,N_28482,N_28328);
nand U29955 (N_29955,N_28391,N_28768);
nor U29956 (N_29956,N_27887,N_28219);
xor U29957 (N_29957,N_28737,N_27902);
or U29958 (N_29958,N_28463,N_28041);
xnor U29959 (N_29959,N_28302,N_27932);
nor U29960 (N_29960,N_27988,N_28379);
xnor U29961 (N_29961,N_28029,N_28225);
or U29962 (N_29962,N_27719,N_28676);
xor U29963 (N_29963,N_28421,N_28201);
and U29964 (N_29964,N_28246,N_27795);
xor U29965 (N_29965,N_27806,N_28694);
and U29966 (N_29966,N_28796,N_27902);
and U29967 (N_29967,N_27696,N_28676);
nor U29968 (N_29968,N_28535,N_28313);
and U29969 (N_29969,N_28707,N_28606);
and U29970 (N_29970,N_28095,N_28115);
nand U29971 (N_29971,N_27876,N_27862);
nor U29972 (N_29972,N_28427,N_27985);
nand U29973 (N_29973,N_28153,N_27991);
xnor U29974 (N_29974,N_28514,N_27655);
nor U29975 (N_29975,N_27872,N_27911);
or U29976 (N_29976,N_27946,N_28477);
xor U29977 (N_29977,N_27827,N_28301);
and U29978 (N_29978,N_28776,N_28257);
xnor U29979 (N_29979,N_27826,N_27948);
xor U29980 (N_29980,N_28071,N_28650);
nor U29981 (N_29981,N_28633,N_28675);
and U29982 (N_29982,N_28424,N_27847);
or U29983 (N_29983,N_28222,N_28005);
and U29984 (N_29984,N_28352,N_28491);
and U29985 (N_29985,N_28118,N_28246);
or U29986 (N_29986,N_27695,N_28763);
nand U29987 (N_29987,N_28231,N_28182);
nor U29988 (N_29988,N_28262,N_27942);
nand U29989 (N_29989,N_28415,N_28711);
xor U29990 (N_29990,N_27654,N_28140);
nand U29991 (N_29991,N_28609,N_27866);
or U29992 (N_29992,N_28285,N_28680);
xnor U29993 (N_29993,N_28030,N_28069);
xor U29994 (N_29994,N_28675,N_28375);
or U29995 (N_29995,N_27943,N_27738);
nor U29996 (N_29996,N_28446,N_27700);
or U29997 (N_29997,N_28199,N_27952);
or U29998 (N_29998,N_27662,N_28485);
or U29999 (N_29999,N_27788,N_28229);
nand UO_0 (O_0,N_29680,N_29099);
xnor UO_1 (O_1,N_29624,N_29421);
and UO_2 (O_2,N_28936,N_29644);
and UO_3 (O_3,N_28824,N_29242);
and UO_4 (O_4,N_28973,N_29512);
nor UO_5 (O_5,N_29326,N_29703);
xnor UO_6 (O_6,N_29258,N_29031);
or UO_7 (O_7,N_29652,N_29145);
nand UO_8 (O_8,N_29581,N_29197);
and UO_9 (O_9,N_29759,N_29308);
nor UO_10 (O_10,N_29494,N_29231);
xor UO_11 (O_11,N_28888,N_29007);
nor UO_12 (O_12,N_29393,N_29929);
or UO_13 (O_13,N_29996,N_29428);
nor UO_14 (O_14,N_28903,N_29232);
nor UO_15 (O_15,N_28800,N_29317);
or UO_16 (O_16,N_29061,N_29685);
nor UO_17 (O_17,N_29637,N_29123);
nand UO_18 (O_18,N_29977,N_29737);
xnor UO_19 (O_19,N_28807,N_29122);
or UO_20 (O_20,N_29464,N_28943);
and UO_21 (O_21,N_29631,N_29873);
nand UO_22 (O_22,N_29828,N_29447);
nand UO_23 (O_23,N_29905,N_29141);
and UO_24 (O_24,N_28933,N_29520);
nor UO_25 (O_25,N_29654,N_29064);
and UO_26 (O_26,N_28978,N_29405);
or UO_27 (O_27,N_28905,N_29869);
and UO_28 (O_28,N_29279,N_28853);
nand UO_29 (O_29,N_29395,N_29057);
xnor UO_30 (O_30,N_29062,N_29424);
nor UO_31 (O_31,N_29843,N_29283);
nor UO_32 (O_32,N_29356,N_29620);
xnor UO_33 (O_33,N_28842,N_29738);
or UO_34 (O_34,N_29128,N_29388);
nand UO_35 (O_35,N_29327,N_29149);
nand UO_36 (O_36,N_29842,N_29855);
xnor UO_37 (O_37,N_28884,N_29210);
nand UO_38 (O_38,N_29343,N_28965);
nand UO_39 (O_39,N_29780,N_29935);
and UO_40 (O_40,N_29697,N_28935);
or UO_41 (O_41,N_29275,N_29962);
or UO_42 (O_42,N_29406,N_29720);
and UO_43 (O_43,N_29303,N_29413);
and UO_44 (O_44,N_29067,N_29300);
xor UO_45 (O_45,N_28873,N_29604);
nor UO_46 (O_46,N_29095,N_28822);
nor UO_47 (O_47,N_29221,N_29993);
and UO_48 (O_48,N_29950,N_28855);
nor UO_49 (O_49,N_28830,N_28963);
nand UO_50 (O_50,N_29609,N_29556);
nor UO_51 (O_51,N_29881,N_29490);
or UO_52 (O_52,N_28945,N_29107);
or UO_53 (O_53,N_29757,N_29941);
nor UO_54 (O_54,N_29389,N_29382);
or UO_55 (O_55,N_29055,N_29955);
nand UO_56 (O_56,N_29176,N_29365);
nand UO_57 (O_57,N_29074,N_29169);
nor UO_58 (O_58,N_29953,N_29079);
xor UO_59 (O_59,N_29900,N_29345);
or UO_60 (O_60,N_29882,N_28849);
xor UO_61 (O_61,N_29222,N_29758);
xor UO_62 (O_62,N_28840,N_29046);
or UO_63 (O_63,N_29845,N_29196);
or UO_64 (O_64,N_28901,N_29323);
nor UO_65 (O_65,N_29133,N_29948);
nor UO_66 (O_66,N_29593,N_29786);
nand UO_67 (O_67,N_28990,N_29366);
nor UO_68 (O_68,N_29618,N_28871);
or UO_69 (O_69,N_29466,N_28832);
or UO_70 (O_70,N_29807,N_29493);
nor UO_71 (O_71,N_29238,N_28815);
nand UO_72 (O_72,N_29336,N_28804);
or UO_73 (O_73,N_28836,N_29188);
nor UO_74 (O_74,N_29653,N_29982);
or UO_75 (O_75,N_29250,N_29126);
xor UO_76 (O_76,N_29130,N_29816);
or UO_77 (O_77,N_29983,N_29723);
and UO_78 (O_78,N_29529,N_29476);
nand UO_79 (O_79,N_29316,N_29741);
and UO_80 (O_80,N_29420,N_28860);
nand UO_81 (O_81,N_29853,N_29314);
xor UO_82 (O_82,N_29156,N_28899);
or UO_83 (O_83,N_28808,N_29949);
and UO_84 (O_84,N_28874,N_28916);
and UO_85 (O_85,N_29722,N_29290);
and UO_86 (O_86,N_29607,N_28861);
xor UO_87 (O_87,N_28959,N_29147);
nor UO_88 (O_88,N_29091,N_29098);
or UO_89 (O_89,N_28881,N_29375);
nand UO_90 (O_90,N_29230,N_29818);
and UO_91 (O_91,N_29416,N_29093);
nand UO_92 (O_92,N_28908,N_29785);
or UO_93 (O_93,N_29744,N_29553);
xor UO_94 (O_94,N_29665,N_28927);
or UO_95 (O_95,N_29177,N_29331);
and UO_96 (O_96,N_29641,N_29585);
or UO_97 (O_97,N_29349,N_29837);
or UO_98 (O_98,N_28955,N_29158);
and UO_99 (O_99,N_29047,N_29391);
nand UO_100 (O_100,N_29752,N_29746);
or UO_101 (O_101,N_29655,N_29364);
nor UO_102 (O_102,N_29782,N_29440);
nor UO_103 (O_103,N_29472,N_29599);
or UO_104 (O_104,N_29932,N_28917);
or UO_105 (O_105,N_29204,N_29632);
nand UO_106 (O_106,N_29352,N_29633);
or UO_107 (O_107,N_29713,N_29059);
nand UO_108 (O_108,N_29338,N_29183);
nor UO_109 (O_109,N_28866,N_29658);
or UO_110 (O_110,N_29749,N_29508);
nand UO_111 (O_111,N_29090,N_29358);
and UO_112 (O_112,N_29524,N_29400);
and UO_113 (O_113,N_28940,N_29261);
or UO_114 (O_114,N_28895,N_29274);
and UO_115 (O_115,N_28829,N_29245);
nor UO_116 (O_116,N_29501,N_29425);
nand UO_117 (O_117,N_29306,N_29159);
nor UO_118 (O_118,N_29913,N_29004);
nor UO_119 (O_119,N_29468,N_29333);
xnor UO_120 (O_120,N_29198,N_29127);
or UO_121 (O_121,N_29482,N_28988);
or UO_122 (O_122,N_29050,N_29346);
and UO_123 (O_123,N_29502,N_29080);
or UO_124 (O_124,N_29259,N_28872);
or UO_125 (O_125,N_29495,N_29761);
or UO_126 (O_126,N_29342,N_29286);
nor UO_127 (O_127,N_28954,N_28956);
xor UO_128 (O_128,N_28854,N_29084);
or UO_129 (O_129,N_28809,N_29817);
nand UO_130 (O_130,N_29419,N_29864);
or UO_131 (O_131,N_29619,N_29826);
and UO_132 (O_132,N_29042,N_29203);
and UO_133 (O_133,N_28968,N_28801);
xnor UO_134 (O_134,N_29426,N_29536);
xnor UO_135 (O_135,N_29399,N_29148);
and UO_136 (O_136,N_28983,N_29726);
or UO_137 (O_137,N_29835,N_28883);
xor UO_138 (O_138,N_28930,N_29574);
nand UO_139 (O_139,N_28868,N_29034);
nand UO_140 (O_140,N_29000,N_28987);
or UO_141 (O_141,N_29721,N_29243);
or UO_142 (O_142,N_29220,N_29473);
or UO_143 (O_143,N_29480,N_29020);
xor UO_144 (O_144,N_28948,N_29712);
and UO_145 (O_145,N_29857,N_29293);
nor UO_146 (O_146,N_29288,N_29899);
nor UO_147 (O_147,N_29871,N_29554);
nand UO_148 (O_148,N_29862,N_29821);
or UO_149 (O_149,N_29995,N_29487);
or UO_150 (O_150,N_28896,N_29990);
xor UO_151 (O_151,N_29451,N_29454);
xor UO_152 (O_152,N_29477,N_29299);
nor UO_153 (O_153,N_29374,N_28915);
and UO_154 (O_154,N_29304,N_29372);
or UO_155 (O_155,N_29182,N_29954);
nor UO_156 (O_156,N_29827,N_29465);
nand UO_157 (O_157,N_29439,N_29320);
nand UO_158 (O_158,N_29269,N_29268);
nand UO_159 (O_159,N_29796,N_29280);
nor UO_160 (O_160,N_28957,N_29498);
nand UO_161 (O_161,N_28938,N_29992);
nand UO_162 (O_162,N_29262,N_28816);
or UO_163 (O_163,N_29690,N_29265);
or UO_164 (O_164,N_29709,N_28929);
nand UO_165 (O_165,N_29435,N_28827);
xnor UO_166 (O_166,N_29150,N_29162);
nand UO_167 (O_167,N_29952,N_29001);
and UO_168 (O_168,N_29040,N_29016);
xor UO_169 (O_169,N_29926,N_29939);
and UO_170 (O_170,N_29676,N_29925);
xor UO_171 (O_171,N_29525,N_29707);
nand UO_172 (O_172,N_29861,N_29630);
nor UO_173 (O_173,N_29589,N_29890);
and UO_174 (O_174,N_29777,N_29436);
nor UO_175 (O_175,N_29448,N_29339);
and UO_176 (O_176,N_29915,N_29155);
or UO_177 (O_177,N_29887,N_28985);
xor UO_178 (O_178,N_29392,N_29402);
xor UO_179 (O_179,N_29089,N_28900);
nor UO_180 (O_180,N_28946,N_29313);
nand UO_181 (O_181,N_28879,N_29533);
nand UO_182 (O_182,N_29594,N_29963);
nor UO_183 (O_183,N_29643,N_29063);
nor UO_184 (O_184,N_29657,N_29276);
nand UO_185 (O_185,N_29174,N_29052);
nor UO_186 (O_186,N_29234,N_29792);
xor UO_187 (O_187,N_29385,N_29394);
nand UO_188 (O_188,N_28970,N_29663);
and UO_189 (O_189,N_29892,N_29783);
xnor UO_190 (O_190,N_28865,N_29297);
and UO_191 (O_191,N_29809,N_29615);
and UO_192 (O_192,N_29635,N_29408);
nand UO_193 (O_193,N_29808,N_29559);
nand UO_194 (O_194,N_28918,N_29852);
nor UO_195 (O_195,N_29705,N_29613);
nand UO_196 (O_196,N_29056,N_29820);
xnor UO_197 (O_197,N_29612,N_28996);
nor UO_198 (O_198,N_29073,N_29626);
and UO_199 (O_199,N_29832,N_29354);
xnor UO_200 (O_200,N_29218,N_28810);
nand UO_201 (O_201,N_29499,N_29701);
nor UO_202 (O_202,N_29934,N_29166);
and UO_203 (O_203,N_28835,N_29544);
and UO_204 (O_204,N_29891,N_29740);
or UO_205 (O_205,N_29679,N_29614);
xnor UO_206 (O_206,N_29695,N_28999);
and UO_207 (O_207,N_29824,N_29788);
nand UO_208 (O_208,N_29180,N_29083);
nor UO_209 (O_209,N_29884,N_29797);
nand UO_210 (O_210,N_29538,N_29754);
or UO_211 (O_211,N_29129,N_29458);
nor UO_212 (O_212,N_29442,N_29627);
nor UO_213 (O_213,N_29557,N_29551);
or UO_214 (O_214,N_29994,N_29805);
and UO_215 (O_215,N_28833,N_29718);
and UO_216 (O_216,N_29284,N_28890);
nor UO_217 (O_217,N_29906,N_29886);
nand UO_218 (O_218,N_29003,N_29489);
nor UO_219 (O_219,N_29138,N_29309);
and UO_220 (O_220,N_29178,N_28831);
or UO_221 (O_221,N_29927,N_29373);
nor UO_222 (O_222,N_29583,N_29564);
nor UO_223 (O_223,N_29651,N_28875);
or UO_224 (O_224,N_29312,N_29694);
nand UO_225 (O_225,N_28837,N_29662);
nor UO_226 (O_226,N_29812,N_29603);
nor UO_227 (O_227,N_29751,N_29264);
nor UO_228 (O_228,N_29931,N_29998);
and UO_229 (O_229,N_29347,N_29770);
xnor UO_230 (O_230,N_28806,N_29674);
nor UO_231 (O_231,N_29344,N_29191);
xnor UO_232 (O_232,N_29521,N_28931);
xnor UO_233 (O_233,N_29682,N_29254);
nand UO_234 (O_234,N_29933,N_29163);
nand UO_235 (O_235,N_29140,N_28911);
or UO_236 (O_236,N_28969,N_29119);
nand UO_237 (O_237,N_29164,N_29113);
and UO_238 (O_238,N_29103,N_28864);
nand UO_239 (O_239,N_29256,N_29184);
nand UO_240 (O_240,N_29763,N_29917);
nand UO_241 (O_241,N_29239,N_29266);
or UO_242 (O_242,N_28897,N_29516);
or UO_243 (O_243,N_28960,N_29810);
nor UO_244 (O_244,N_28993,N_28974);
or UO_245 (O_245,N_29901,N_29880);
xnor UO_246 (O_246,N_29431,N_29340);
nor UO_247 (O_247,N_29224,N_29137);
xor UO_248 (O_248,N_29659,N_29207);
xor UO_249 (O_249,N_29195,N_29171);
nor UO_250 (O_250,N_29959,N_29277);
or UO_251 (O_251,N_28820,N_29241);
or UO_252 (O_252,N_28975,N_29175);
or UO_253 (O_253,N_29865,N_29208);
or UO_254 (O_254,N_29018,N_29296);
nor UO_255 (O_255,N_29838,N_29965);
xor UO_256 (O_256,N_29729,N_29444);
nor UO_257 (O_257,N_28859,N_29823);
or UO_258 (O_258,N_29371,N_29360);
and UO_259 (O_259,N_29211,N_29748);
and UO_260 (O_260,N_29443,N_29687);
xnor UO_261 (O_261,N_29033,N_29830);
xnor UO_262 (O_262,N_29492,N_28907);
or UO_263 (O_263,N_29131,N_29606);
nor UO_264 (O_264,N_28921,N_29453);
nand UO_265 (O_265,N_28949,N_29475);
xor UO_266 (O_266,N_29844,N_28850);
or UO_267 (O_267,N_29839,N_29681);
nand UO_268 (O_268,N_29692,N_29152);
nand UO_269 (O_269,N_29968,N_28906);
or UO_270 (O_270,N_29505,N_29597);
xnor UO_271 (O_271,N_29854,N_29700);
nor UO_272 (O_272,N_29135,N_29247);
xnor UO_273 (O_273,N_29918,N_29904);
nand UO_274 (O_274,N_29936,N_29908);
xor UO_275 (O_275,N_28997,N_29579);
xnor UO_276 (O_276,N_29071,N_29571);
or UO_277 (O_277,N_29429,N_29656);
xnor UO_278 (O_278,N_28847,N_29106);
or UO_279 (O_279,N_29217,N_29455);
xor UO_280 (O_280,N_29251,N_29206);
nor UO_281 (O_281,N_28821,N_28998);
nor UO_282 (O_282,N_29878,N_29628);
nor UO_283 (O_283,N_29575,N_29157);
xor UO_284 (O_284,N_29975,N_29021);
and UO_285 (O_285,N_29831,N_29380);
nand UO_286 (O_286,N_29947,N_29212);
nor UO_287 (O_287,N_29822,N_29229);
xnor UO_288 (O_288,N_29923,N_29847);
and UO_289 (O_289,N_29005,N_29181);
nand UO_290 (O_290,N_28803,N_29072);
or UO_291 (O_291,N_29910,N_29577);
xor UO_292 (O_292,N_28814,N_29856);
nand UO_293 (O_293,N_28889,N_28986);
nand UO_294 (O_294,N_29790,N_29417);
or UO_295 (O_295,N_29795,N_29096);
nand UO_296 (O_296,N_29699,N_28932);
xnor UO_297 (O_297,N_29036,N_29094);
xnor UO_298 (O_298,N_29240,N_29298);
nor UO_299 (O_299,N_29228,N_29573);
and UO_300 (O_300,N_29236,N_29872);
and UO_301 (O_301,N_29580,N_29986);
and UO_302 (O_302,N_29885,N_28919);
nor UO_303 (O_303,N_29045,N_29528);
xor UO_304 (O_304,N_29909,N_29545);
nand UO_305 (O_305,N_28852,N_28839);
or UO_306 (O_306,N_29111,N_29200);
or UO_307 (O_307,N_28898,N_29441);
and UO_308 (O_308,N_29903,N_28811);
and UO_309 (O_309,N_29307,N_29038);
nand UO_310 (O_310,N_29246,N_29534);
xor UO_311 (O_311,N_29060,N_28812);
nor UO_312 (O_312,N_29984,N_29086);
nor UO_313 (O_313,N_29483,N_29840);
or UO_314 (O_314,N_29134,N_29562);
xnor UO_315 (O_315,N_29860,N_29226);
and UO_316 (O_316,N_29957,N_29139);
xnor UO_317 (O_317,N_29289,N_29849);
or UO_318 (O_318,N_29081,N_28980);
and UO_319 (O_319,N_29278,N_29112);
nor UO_320 (O_320,N_29146,N_29069);
or UO_321 (O_321,N_29076,N_29459);
nor UO_322 (O_322,N_29814,N_29077);
and UO_323 (O_323,N_29486,N_29334);
and UO_324 (O_324,N_29698,N_29725);
and UO_325 (O_325,N_29396,N_29542);
nor UO_326 (O_326,N_29980,N_29370);
or UO_327 (O_327,N_29944,N_28976);
xor UO_328 (O_328,N_29558,N_29561);
nand UO_329 (O_329,N_29760,N_29418);
nor UO_330 (O_330,N_29255,N_29315);
xor UO_331 (O_331,N_29012,N_29017);
xor UO_332 (O_332,N_29404,N_29478);
nand UO_333 (O_333,N_29895,N_28834);
nand UO_334 (O_334,N_28991,N_29517);
xor UO_335 (O_335,N_29118,N_29876);
nand UO_336 (O_336,N_29078,N_29590);
and UO_337 (O_337,N_29252,N_29467);
xnor UO_338 (O_338,N_29781,N_29715);
xnor UO_339 (O_339,N_29514,N_28951);
and UO_340 (O_340,N_29154,N_28813);
nand UO_341 (O_341,N_29006,N_29249);
nor UO_342 (O_342,N_29319,N_28924);
or UO_343 (O_343,N_29728,N_29811);
or UO_344 (O_344,N_29430,N_29622);
or UO_345 (O_345,N_29523,N_28902);
xnor UO_346 (O_346,N_29011,N_29522);
nand UO_347 (O_347,N_29548,N_29225);
and UO_348 (O_348,N_29964,N_29543);
or UO_349 (O_349,N_29834,N_29945);
and UO_350 (O_350,N_29087,N_28862);
xnor UO_351 (O_351,N_29105,N_29648);
xor UO_352 (O_352,N_29967,N_29030);
nand UO_353 (O_353,N_29914,N_28802);
nand UO_354 (O_354,N_29019,N_29570);
or UO_355 (O_355,N_29800,N_29706);
and UO_356 (O_356,N_29969,N_29341);
and UO_357 (O_357,N_28870,N_29693);
nand UO_358 (O_358,N_28942,N_29190);
and UO_359 (O_359,N_29065,N_28926);
xor UO_360 (O_360,N_28920,N_29647);
nor UO_361 (O_361,N_29841,N_29732);
or UO_362 (O_362,N_28972,N_28967);
or UO_363 (O_363,N_29337,N_29291);
xnor UO_364 (O_364,N_28982,N_28856);
or UO_365 (O_365,N_28989,N_29686);
nand UO_366 (O_366,N_29025,N_29970);
and UO_367 (O_367,N_29661,N_29068);
and UO_368 (O_368,N_29775,N_29422);
nor UO_369 (O_369,N_28909,N_28863);
nand UO_370 (O_370,N_28844,N_29547);
xnor UO_371 (O_371,N_29114,N_29646);
or UO_372 (O_372,N_29048,N_29791);
xnor UO_373 (O_373,N_29649,N_29889);
and UO_374 (O_374,N_29024,N_29414);
nand UO_375 (O_375,N_29596,N_29032);
or UO_376 (O_376,N_29121,N_29956);
and UO_377 (O_377,N_29769,N_29383);
or UO_378 (O_378,N_29285,N_29668);
nand UO_379 (O_379,N_29481,N_28923);
nor UO_380 (O_380,N_29958,N_28848);
nor UO_381 (O_381,N_29167,N_29946);
xor UO_382 (O_382,N_29199,N_29988);
nand UO_383 (O_383,N_29683,N_29407);
nor UO_384 (O_384,N_28979,N_29287);
nand UO_385 (O_385,N_29485,N_29474);
nor UO_386 (O_386,N_28886,N_29381);
nor UO_387 (O_387,N_29940,N_29888);
nand UO_388 (O_388,N_28817,N_29518);
or UO_389 (O_389,N_29051,N_29971);
and UO_390 (O_390,N_29896,N_29634);
or UO_391 (O_391,N_29640,N_29292);
and UO_392 (O_392,N_29507,N_28966);
xnor UO_393 (O_393,N_29773,N_29202);
and UO_394 (O_394,N_29423,N_29102);
nor UO_395 (O_395,N_29066,N_29829);
nor UO_396 (O_396,N_29710,N_29922);
nand UO_397 (O_397,N_29546,N_29803);
or UO_398 (O_398,N_29273,N_29696);
or UO_399 (O_399,N_29456,N_29858);
or UO_400 (O_400,N_29919,N_29353);
or UO_401 (O_401,N_29527,N_28869);
or UO_402 (O_402,N_29912,N_29041);
or UO_403 (O_403,N_29433,N_28995);
and UO_404 (O_404,N_29552,N_29201);
nor UO_405 (O_405,N_29739,N_29144);
xnor UO_406 (O_406,N_29755,N_29531);
and UO_407 (O_407,N_29010,N_29670);
nor UO_408 (O_408,N_29043,N_28878);
nor UO_409 (O_409,N_28838,N_29742);
xnor UO_410 (O_410,N_29153,N_29611);
xor UO_411 (O_411,N_29966,N_28941);
and UO_412 (O_412,N_29160,N_29974);
xnor UO_413 (O_413,N_29410,N_29802);
or UO_414 (O_414,N_29461,N_29578);
and UO_415 (O_415,N_28977,N_29743);
nand UO_416 (O_416,N_29263,N_29943);
xor UO_417 (O_417,N_29403,N_28992);
and UO_418 (O_418,N_29026,N_29774);
xnor UO_419 (O_419,N_29916,N_29675);
nor UO_420 (O_420,N_29348,N_29223);
xnor UO_421 (O_421,N_28858,N_29446);
nor UO_422 (O_422,N_29582,N_29397);
or UO_423 (O_423,N_29833,N_29961);
or UO_424 (O_424,N_28928,N_29125);
or UO_425 (O_425,N_28876,N_29766);
xor UO_426 (O_426,N_29376,N_29667);
xor UO_427 (O_427,N_29227,N_29727);
or UO_428 (O_428,N_29677,N_29806);
and UO_429 (O_429,N_29463,N_29415);
and UO_430 (O_430,N_29151,N_29897);
xor UO_431 (O_431,N_29669,N_29576);
and UO_432 (O_432,N_29870,N_29355);
nand UO_433 (O_433,N_29765,N_29330);
or UO_434 (O_434,N_28846,N_28934);
or UO_435 (O_435,N_29629,N_29716);
or UO_436 (O_436,N_29815,N_29555);
nand UO_437 (O_437,N_29951,N_29793);
xor UO_438 (O_438,N_29022,N_29506);
or UO_439 (O_439,N_28828,N_29617);
or UO_440 (O_440,N_29412,N_28912);
or UO_441 (O_441,N_28893,N_29602);
nor UO_442 (O_442,N_29318,N_29601);
or UO_443 (O_443,N_29539,N_29846);
xor UO_444 (O_444,N_29504,N_29733);
nor UO_445 (O_445,N_29438,N_29039);
or UO_446 (O_446,N_29650,N_29161);
nor UO_447 (O_447,N_28826,N_29271);
nor UO_448 (O_448,N_28922,N_29708);
and UO_449 (O_449,N_29002,N_29013);
nand UO_450 (O_450,N_29471,N_29704);
or UO_451 (O_451,N_29401,N_29978);
nor UO_452 (O_452,N_29328,N_28851);
nor UO_453 (O_453,N_29192,N_29101);
nor UO_454 (O_454,N_28818,N_29666);
or UO_455 (O_455,N_28981,N_29526);
xnor UO_456 (O_456,N_29115,N_29866);
or UO_457 (O_457,N_29605,N_29282);
or UO_458 (O_458,N_29563,N_29863);
or UO_459 (O_459,N_29058,N_29771);
nor UO_460 (O_460,N_29462,N_29497);
nor UO_461 (O_461,N_28882,N_28885);
xor UO_462 (O_462,N_29270,N_28962);
nor UO_463 (O_463,N_29764,N_29642);
nor UO_464 (O_464,N_29351,N_29928);
nand UO_465 (O_465,N_29515,N_29660);
or UO_466 (O_466,N_29350,N_29689);
nand UO_467 (O_467,N_29215,N_29363);
nor UO_468 (O_468,N_29819,N_29859);
xnor UO_469 (O_469,N_28819,N_28937);
or UO_470 (O_470,N_29684,N_29898);
and UO_471 (O_471,N_29608,N_29049);
or UO_472 (O_472,N_29734,N_29789);
and UO_473 (O_473,N_29804,N_29850);
or UO_474 (O_474,N_29029,N_28984);
and UO_475 (O_475,N_29550,N_29836);
nand UO_476 (O_476,N_29037,N_29999);
xor UO_477 (O_477,N_29310,N_29623);
xnor UO_478 (O_478,N_29437,N_28877);
nand UO_479 (O_479,N_29193,N_28950);
or UO_480 (O_480,N_29894,N_29997);
xnor UO_481 (O_481,N_29027,N_29621);
nor UO_482 (O_482,N_28891,N_29569);
or UO_483 (O_483,N_28894,N_29092);
nor UO_484 (O_484,N_29257,N_29768);
and UO_485 (O_485,N_28958,N_29595);
or UO_486 (O_486,N_29717,N_29496);
xnor UO_487 (O_487,N_29588,N_29108);
xor UO_488 (O_488,N_29452,N_29636);
xnor UO_489 (O_489,N_29902,N_29981);
nand UO_490 (O_490,N_29235,N_29124);
or UO_491 (O_491,N_29479,N_28892);
nor UO_492 (O_492,N_29302,N_29750);
nor UO_493 (O_493,N_29519,N_29924);
xnor UO_494 (O_494,N_29053,N_29205);
and UO_495 (O_495,N_29384,N_29168);
nor UO_496 (O_496,N_29100,N_29600);
or UO_497 (O_497,N_29879,N_29530);
xor UO_498 (O_498,N_29719,N_29549);
xnor UO_499 (O_499,N_29491,N_29591);
and UO_500 (O_500,N_29672,N_29387);
or UO_501 (O_501,N_29378,N_28823);
and UO_502 (O_502,N_29398,N_29784);
xor UO_503 (O_503,N_29120,N_28947);
or UO_504 (O_504,N_29295,N_29104);
nand UO_505 (O_505,N_28880,N_28952);
xor UO_506 (O_506,N_29813,N_29484);
or UO_507 (O_507,N_29979,N_29972);
or UO_508 (O_508,N_29116,N_29173);
xnor UO_509 (O_509,N_29592,N_28825);
and UO_510 (O_510,N_29976,N_29678);
xnor UO_511 (O_511,N_29253,N_29367);
xnor UO_512 (O_512,N_29893,N_28914);
and UO_513 (O_513,N_29469,N_29445);
and UO_514 (O_514,N_29434,N_29851);
and UO_515 (O_515,N_29085,N_29321);
xor UO_516 (O_516,N_29427,N_29960);
nand UO_517 (O_517,N_29762,N_29794);
and UO_518 (O_518,N_29500,N_29097);
or UO_519 (O_519,N_29987,N_28913);
xor UO_520 (O_520,N_29610,N_29142);
nor UO_521 (O_521,N_29023,N_29332);
and UO_522 (O_522,N_29921,N_29799);
and UO_523 (O_523,N_29260,N_29187);
and UO_524 (O_524,N_29432,N_29008);
nor UO_525 (O_525,N_29711,N_29324);
or UO_526 (O_526,N_29368,N_29179);
nand UO_527 (O_527,N_29883,N_29054);
or UO_528 (O_528,N_29671,N_29237);
nor UO_529 (O_529,N_29014,N_29736);
and UO_530 (O_530,N_28994,N_29511);
nand UO_531 (O_531,N_29189,N_28961);
nor UO_532 (O_532,N_29165,N_29625);
nand UO_533 (O_533,N_29568,N_29244);
xor UO_534 (O_534,N_29688,N_29329);
xnor UO_535 (O_535,N_29572,N_29362);
nand UO_536 (O_536,N_29170,N_29532);
nand UO_537 (O_537,N_29503,N_29216);
or UO_538 (O_538,N_29776,N_29567);
or UO_539 (O_539,N_29136,N_29015);
nand UO_540 (O_540,N_29028,N_29541);
nand UO_541 (O_541,N_28944,N_29616);
and UO_542 (O_542,N_29639,N_29848);
or UO_543 (O_543,N_29537,N_29778);
nor UO_544 (O_544,N_29488,N_29335);
nand UO_545 (O_545,N_29673,N_29450);
xnor UO_546 (O_546,N_28857,N_29143);
xnor UO_547 (O_547,N_29787,N_29691);
and UO_548 (O_548,N_29877,N_29379);
nor UO_549 (O_549,N_29513,N_28845);
nor UO_550 (O_550,N_29219,N_29117);
nor UO_551 (O_551,N_29540,N_29991);
nor UO_552 (O_552,N_29359,N_28964);
and UO_553 (O_553,N_29664,N_29801);
nand UO_554 (O_554,N_29560,N_29294);
nand UO_555 (O_555,N_28805,N_29460);
and UO_556 (O_556,N_29645,N_29305);
nand UO_557 (O_557,N_29584,N_29989);
or UO_558 (O_558,N_29301,N_29756);
nand UO_559 (O_559,N_29724,N_29779);
nor UO_560 (O_560,N_29772,N_29386);
and UO_561 (O_561,N_29369,N_29920);
xor UO_562 (O_562,N_29361,N_29044);
or UO_563 (O_563,N_29874,N_29937);
xor UO_564 (O_564,N_29911,N_29390);
nor UO_565 (O_565,N_28867,N_29248);
and UO_566 (O_566,N_29132,N_28910);
or UO_567 (O_567,N_29449,N_29233);
nand UO_568 (O_568,N_29868,N_29867);
xor UO_569 (O_569,N_29075,N_29272);
nand UO_570 (O_570,N_29745,N_29942);
xnor UO_571 (O_571,N_29907,N_29930);
or UO_572 (O_572,N_29035,N_29875);
nand UO_573 (O_573,N_29587,N_29510);
or UO_574 (O_574,N_29377,N_29731);
or UO_575 (O_575,N_29325,N_29586);
or UO_576 (O_576,N_29172,N_29214);
nor UO_577 (O_577,N_28841,N_28953);
or UO_578 (O_578,N_29565,N_29753);
xnor UO_579 (O_579,N_29825,N_29185);
nand UO_580 (O_580,N_29535,N_29973);
xor UO_581 (O_581,N_29186,N_29457);
or UO_582 (O_582,N_29411,N_29470);
nand UO_583 (O_583,N_28887,N_29194);
or UO_584 (O_584,N_29702,N_29714);
and UO_585 (O_585,N_28925,N_29088);
and UO_586 (O_586,N_29322,N_29509);
or UO_587 (O_587,N_28904,N_29598);
xor UO_588 (O_588,N_29070,N_29281);
and UO_589 (O_589,N_29082,N_29747);
xor UO_590 (O_590,N_29985,N_29209);
xnor UO_591 (O_591,N_29566,N_29109);
xnor UO_592 (O_592,N_29767,N_29638);
nand UO_593 (O_593,N_29735,N_29798);
nand UO_594 (O_594,N_29357,N_29213);
or UO_595 (O_595,N_28843,N_29311);
nor UO_596 (O_596,N_29730,N_29110);
nor UO_597 (O_597,N_28939,N_29009);
or UO_598 (O_598,N_28971,N_29938);
nand UO_599 (O_599,N_29267,N_29409);
nand UO_600 (O_600,N_28806,N_29952);
or UO_601 (O_601,N_29842,N_29838);
nand UO_602 (O_602,N_29388,N_29229);
nand UO_603 (O_603,N_29878,N_28945);
and UO_604 (O_604,N_29179,N_29552);
or UO_605 (O_605,N_29266,N_29911);
xnor UO_606 (O_606,N_29965,N_29464);
or UO_607 (O_607,N_29733,N_29854);
and UO_608 (O_608,N_29875,N_28971);
nand UO_609 (O_609,N_29699,N_28906);
nand UO_610 (O_610,N_29149,N_29247);
nor UO_611 (O_611,N_29553,N_28883);
or UO_612 (O_612,N_29450,N_29651);
nor UO_613 (O_613,N_29988,N_28819);
or UO_614 (O_614,N_29965,N_28865);
xnor UO_615 (O_615,N_28852,N_29408);
or UO_616 (O_616,N_28801,N_29970);
nor UO_617 (O_617,N_29736,N_29849);
xor UO_618 (O_618,N_29461,N_29625);
nor UO_619 (O_619,N_29446,N_29589);
nor UO_620 (O_620,N_29417,N_29263);
nand UO_621 (O_621,N_29618,N_29034);
nand UO_622 (O_622,N_29056,N_29747);
nor UO_623 (O_623,N_29692,N_29382);
and UO_624 (O_624,N_29334,N_29833);
nand UO_625 (O_625,N_29982,N_29689);
or UO_626 (O_626,N_29555,N_28826);
nand UO_627 (O_627,N_29367,N_29782);
nand UO_628 (O_628,N_29916,N_28933);
and UO_629 (O_629,N_29477,N_29516);
nor UO_630 (O_630,N_28943,N_29046);
nand UO_631 (O_631,N_29422,N_29902);
xor UO_632 (O_632,N_28888,N_29731);
and UO_633 (O_633,N_28982,N_29533);
or UO_634 (O_634,N_29972,N_29905);
or UO_635 (O_635,N_28931,N_28924);
nor UO_636 (O_636,N_29951,N_29359);
or UO_637 (O_637,N_29696,N_29145);
xnor UO_638 (O_638,N_29351,N_29627);
and UO_639 (O_639,N_29203,N_29730);
nor UO_640 (O_640,N_29241,N_29839);
or UO_641 (O_641,N_29156,N_28932);
nand UO_642 (O_642,N_29024,N_29030);
or UO_643 (O_643,N_29994,N_29183);
xnor UO_644 (O_644,N_29229,N_29755);
nor UO_645 (O_645,N_29156,N_29406);
nand UO_646 (O_646,N_29306,N_29882);
nand UO_647 (O_647,N_29652,N_29439);
nand UO_648 (O_648,N_29214,N_29372);
nand UO_649 (O_649,N_29955,N_29913);
nand UO_650 (O_650,N_29768,N_29101);
nand UO_651 (O_651,N_28872,N_28928);
xnor UO_652 (O_652,N_29423,N_29579);
nor UO_653 (O_653,N_29186,N_29547);
xor UO_654 (O_654,N_29638,N_29963);
and UO_655 (O_655,N_29367,N_28818);
xor UO_656 (O_656,N_29707,N_29063);
and UO_657 (O_657,N_29149,N_29974);
and UO_658 (O_658,N_29384,N_29154);
nand UO_659 (O_659,N_29145,N_29509);
xnor UO_660 (O_660,N_29845,N_29626);
nand UO_661 (O_661,N_28954,N_29199);
and UO_662 (O_662,N_28807,N_29656);
or UO_663 (O_663,N_29781,N_29940);
nand UO_664 (O_664,N_29134,N_29136);
nand UO_665 (O_665,N_29127,N_29206);
and UO_666 (O_666,N_29397,N_29216);
and UO_667 (O_667,N_29563,N_29697);
and UO_668 (O_668,N_28896,N_28905);
and UO_669 (O_669,N_29882,N_29632);
xor UO_670 (O_670,N_29091,N_29960);
or UO_671 (O_671,N_29979,N_29540);
nand UO_672 (O_672,N_29088,N_29966);
nor UO_673 (O_673,N_29114,N_29457);
or UO_674 (O_674,N_29828,N_29958);
xor UO_675 (O_675,N_29430,N_29955);
or UO_676 (O_676,N_29958,N_29377);
and UO_677 (O_677,N_29274,N_28986);
or UO_678 (O_678,N_29407,N_29465);
xnor UO_679 (O_679,N_28812,N_29091);
nand UO_680 (O_680,N_29075,N_28922);
or UO_681 (O_681,N_29989,N_29115);
and UO_682 (O_682,N_29526,N_29616);
nor UO_683 (O_683,N_29070,N_29825);
and UO_684 (O_684,N_29370,N_29621);
and UO_685 (O_685,N_29347,N_29532);
nand UO_686 (O_686,N_29874,N_29725);
or UO_687 (O_687,N_29455,N_29240);
and UO_688 (O_688,N_29442,N_28981);
and UO_689 (O_689,N_29867,N_28822);
nand UO_690 (O_690,N_29365,N_29820);
nor UO_691 (O_691,N_29967,N_29849);
nand UO_692 (O_692,N_28815,N_29753);
and UO_693 (O_693,N_28811,N_29051);
and UO_694 (O_694,N_29927,N_29046);
or UO_695 (O_695,N_29469,N_28827);
nand UO_696 (O_696,N_29548,N_29372);
nor UO_697 (O_697,N_28851,N_29786);
and UO_698 (O_698,N_29166,N_28874);
and UO_699 (O_699,N_29097,N_29124);
or UO_700 (O_700,N_28951,N_29774);
xor UO_701 (O_701,N_29506,N_29694);
and UO_702 (O_702,N_29632,N_28918);
and UO_703 (O_703,N_29098,N_29448);
or UO_704 (O_704,N_29595,N_29883);
nand UO_705 (O_705,N_29862,N_29053);
xor UO_706 (O_706,N_29628,N_29135);
or UO_707 (O_707,N_29182,N_29025);
xnor UO_708 (O_708,N_29297,N_29727);
xnor UO_709 (O_709,N_29036,N_29084);
nor UO_710 (O_710,N_29939,N_29457);
nand UO_711 (O_711,N_28886,N_29831);
nor UO_712 (O_712,N_29538,N_28861);
nand UO_713 (O_713,N_29669,N_29157);
or UO_714 (O_714,N_29185,N_28911);
nand UO_715 (O_715,N_29683,N_29111);
or UO_716 (O_716,N_28896,N_28957);
nor UO_717 (O_717,N_29472,N_29146);
nor UO_718 (O_718,N_29318,N_29308);
nand UO_719 (O_719,N_29484,N_28991);
and UO_720 (O_720,N_29246,N_29962);
xor UO_721 (O_721,N_29711,N_29671);
nor UO_722 (O_722,N_29153,N_29628);
and UO_723 (O_723,N_29256,N_28961);
nor UO_724 (O_724,N_29783,N_29753);
nand UO_725 (O_725,N_29153,N_29418);
nand UO_726 (O_726,N_29150,N_29586);
or UO_727 (O_727,N_29175,N_29632);
or UO_728 (O_728,N_29612,N_29438);
xor UO_729 (O_729,N_29633,N_29177);
and UO_730 (O_730,N_29575,N_29491);
xor UO_731 (O_731,N_29566,N_28968);
and UO_732 (O_732,N_29794,N_29555);
nand UO_733 (O_733,N_29809,N_29999);
or UO_734 (O_734,N_29635,N_28843);
nor UO_735 (O_735,N_29042,N_29497);
nand UO_736 (O_736,N_29418,N_28824);
or UO_737 (O_737,N_29663,N_29555);
or UO_738 (O_738,N_29257,N_29642);
nand UO_739 (O_739,N_28881,N_29058);
nand UO_740 (O_740,N_29211,N_29709);
nand UO_741 (O_741,N_29268,N_29234);
nor UO_742 (O_742,N_29555,N_29173);
and UO_743 (O_743,N_29192,N_29990);
and UO_744 (O_744,N_29394,N_29581);
nor UO_745 (O_745,N_29051,N_29774);
xnor UO_746 (O_746,N_29388,N_29302);
nand UO_747 (O_747,N_29559,N_29880);
and UO_748 (O_748,N_29146,N_29217);
nand UO_749 (O_749,N_29862,N_28975);
xnor UO_750 (O_750,N_29651,N_29508);
or UO_751 (O_751,N_28955,N_29245);
xor UO_752 (O_752,N_29463,N_29459);
or UO_753 (O_753,N_29826,N_29746);
xor UO_754 (O_754,N_29521,N_29630);
and UO_755 (O_755,N_29408,N_29751);
nand UO_756 (O_756,N_29009,N_29974);
and UO_757 (O_757,N_29974,N_28957);
nor UO_758 (O_758,N_29342,N_29078);
and UO_759 (O_759,N_29638,N_29219);
nand UO_760 (O_760,N_29063,N_29356);
nand UO_761 (O_761,N_28909,N_29458);
xor UO_762 (O_762,N_29353,N_29555);
xnor UO_763 (O_763,N_29160,N_29701);
nor UO_764 (O_764,N_29408,N_29055);
or UO_765 (O_765,N_29204,N_29095);
and UO_766 (O_766,N_29099,N_29000);
or UO_767 (O_767,N_29059,N_29453);
xor UO_768 (O_768,N_29159,N_29664);
nor UO_769 (O_769,N_29592,N_29701);
and UO_770 (O_770,N_29302,N_28806);
and UO_771 (O_771,N_29176,N_29010);
and UO_772 (O_772,N_29633,N_29407);
xnor UO_773 (O_773,N_29633,N_29944);
nor UO_774 (O_774,N_29753,N_28918);
xnor UO_775 (O_775,N_28994,N_29966);
xor UO_776 (O_776,N_29283,N_29439);
or UO_777 (O_777,N_29608,N_29442);
or UO_778 (O_778,N_29580,N_29809);
xor UO_779 (O_779,N_29789,N_29837);
nand UO_780 (O_780,N_28870,N_29984);
xnor UO_781 (O_781,N_28929,N_29559);
nor UO_782 (O_782,N_29486,N_29393);
xor UO_783 (O_783,N_29483,N_29993);
nor UO_784 (O_784,N_29817,N_29403);
or UO_785 (O_785,N_29199,N_29440);
nor UO_786 (O_786,N_28841,N_29356);
nand UO_787 (O_787,N_29519,N_29773);
nor UO_788 (O_788,N_29225,N_29514);
nor UO_789 (O_789,N_29791,N_29174);
and UO_790 (O_790,N_29080,N_29153);
or UO_791 (O_791,N_29643,N_29768);
nor UO_792 (O_792,N_29551,N_29398);
nor UO_793 (O_793,N_29557,N_29031);
and UO_794 (O_794,N_29656,N_29728);
and UO_795 (O_795,N_28889,N_29157);
nand UO_796 (O_796,N_29792,N_29909);
nor UO_797 (O_797,N_29223,N_29118);
xor UO_798 (O_798,N_29181,N_29340);
nor UO_799 (O_799,N_28821,N_28971);
nor UO_800 (O_800,N_29121,N_29243);
and UO_801 (O_801,N_29632,N_29358);
or UO_802 (O_802,N_28817,N_29974);
xor UO_803 (O_803,N_29043,N_29101);
xor UO_804 (O_804,N_29367,N_29810);
or UO_805 (O_805,N_29292,N_29612);
or UO_806 (O_806,N_29349,N_29211);
nand UO_807 (O_807,N_29794,N_28842);
or UO_808 (O_808,N_28819,N_29860);
nor UO_809 (O_809,N_29668,N_29743);
nor UO_810 (O_810,N_28992,N_29813);
nand UO_811 (O_811,N_29108,N_28902);
nand UO_812 (O_812,N_29020,N_28988);
or UO_813 (O_813,N_29406,N_29480);
nor UO_814 (O_814,N_29546,N_29722);
xor UO_815 (O_815,N_29901,N_28868);
nor UO_816 (O_816,N_29493,N_29509);
nand UO_817 (O_817,N_29458,N_28940);
or UO_818 (O_818,N_29921,N_29961);
xnor UO_819 (O_819,N_29993,N_28915);
nand UO_820 (O_820,N_29263,N_28826);
nor UO_821 (O_821,N_29153,N_29598);
xor UO_822 (O_822,N_29803,N_28999);
nor UO_823 (O_823,N_29138,N_29944);
and UO_824 (O_824,N_29783,N_29891);
nor UO_825 (O_825,N_29255,N_29532);
or UO_826 (O_826,N_29429,N_29621);
nand UO_827 (O_827,N_28824,N_28845);
or UO_828 (O_828,N_29532,N_29977);
and UO_829 (O_829,N_29255,N_29893);
and UO_830 (O_830,N_28868,N_29928);
xor UO_831 (O_831,N_29470,N_29929);
or UO_832 (O_832,N_29285,N_28894);
nand UO_833 (O_833,N_29140,N_28910);
xor UO_834 (O_834,N_29568,N_29404);
and UO_835 (O_835,N_29812,N_29521);
and UO_836 (O_836,N_29519,N_29371);
and UO_837 (O_837,N_28846,N_29782);
nor UO_838 (O_838,N_28990,N_29416);
nor UO_839 (O_839,N_29536,N_28805);
and UO_840 (O_840,N_29280,N_29621);
or UO_841 (O_841,N_28845,N_28814);
or UO_842 (O_842,N_28845,N_29209);
nand UO_843 (O_843,N_29140,N_29177);
or UO_844 (O_844,N_29237,N_29889);
and UO_845 (O_845,N_29332,N_29899);
or UO_846 (O_846,N_29724,N_28952);
or UO_847 (O_847,N_29035,N_29637);
nand UO_848 (O_848,N_29571,N_29224);
nand UO_849 (O_849,N_29653,N_29892);
nand UO_850 (O_850,N_29336,N_29129);
xnor UO_851 (O_851,N_29482,N_28937);
nand UO_852 (O_852,N_29049,N_29510);
and UO_853 (O_853,N_29165,N_29762);
xnor UO_854 (O_854,N_29756,N_29528);
and UO_855 (O_855,N_29041,N_29793);
nor UO_856 (O_856,N_29326,N_29505);
xor UO_857 (O_857,N_29677,N_28831);
xor UO_858 (O_858,N_29883,N_29483);
nand UO_859 (O_859,N_28823,N_29398);
or UO_860 (O_860,N_29915,N_29640);
nor UO_861 (O_861,N_29053,N_29793);
nand UO_862 (O_862,N_29821,N_29306);
xor UO_863 (O_863,N_29794,N_28858);
and UO_864 (O_864,N_29335,N_28982);
xor UO_865 (O_865,N_29502,N_28986);
nand UO_866 (O_866,N_28883,N_29586);
or UO_867 (O_867,N_29772,N_29114);
nor UO_868 (O_868,N_29777,N_29321);
xor UO_869 (O_869,N_28802,N_29059);
xnor UO_870 (O_870,N_29949,N_29557);
xor UO_871 (O_871,N_29509,N_29403);
nand UO_872 (O_872,N_29299,N_29506);
xnor UO_873 (O_873,N_29063,N_29670);
and UO_874 (O_874,N_28978,N_29458);
or UO_875 (O_875,N_29992,N_29501);
nor UO_876 (O_876,N_28885,N_29806);
nor UO_877 (O_877,N_29634,N_29012);
and UO_878 (O_878,N_29313,N_29203);
nor UO_879 (O_879,N_29763,N_29180);
or UO_880 (O_880,N_29704,N_29507);
xor UO_881 (O_881,N_29147,N_29261);
and UO_882 (O_882,N_29644,N_29885);
nand UO_883 (O_883,N_29431,N_29524);
nand UO_884 (O_884,N_29787,N_28998);
nor UO_885 (O_885,N_29666,N_29336);
or UO_886 (O_886,N_29473,N_29229);
nand UO_887 (O_887,N_29700,N_29094);
xor UO_888 (O_888,N_29841,N_28976);
and UO_889 (O_889,N_29013,N_29198);
xnor UO_890 (O_890,N_29317,N_29784);
xnor UO_891 (O_891,N_28821,N_29722);
and UO_892 (O_892,N_29433,N_28890);
xnor UO_893 (O_893,N_28939,N_29981);
nor UO_894 (O_894,N_29787,N_29933);
and UO_895 (O_895,N_29248,N_29708);
nor UO_896 (O_896,N_29845,N_29682);
xnor UO_897 (O_897,N_29585,N_28862);
xnor UO_898 (O_898,N_29745,N_29573);
nor UO_899 (O_899,N_29440,N_29895);
xnor UO_900 (O_900,N_29091,N_29875);
or UO_901 (O_901,N_29049,N_29566);
nand UO_902 (O_902,N_29585,N_29442);
xnor UO_903 (O_903,N_29880,N_29228);
xor UO_904 (O_904,N_29927,N_29155);
nand UO_905 (O_905,N_29475,N_29592);
or UO_906 (O_906,N_29695,N_29043);
nand UO_907 (O_907,N_29461,N_29278);
nor UO_908 (O_908,N_29884,N_29136);
and UO_909 (O_909,N_29190,N_28921);
nand UO_910 (O_910,N_28890,N_29895);
xor UO_911 (O_911,N_29331,N_29729);
xnor UO_912 (O_912,N_29718,N_28834);
nand UO_913 (O_913,N_29479,N_29843);
xor UO_914 (O_914,N_28842,N_29324);
xnor UO_915 (O_915,N_29206,N_29974);
or UO_916 (O_916,N_29047,N_28966);
nor UO_917 (O_917,N_29362,N_29232);
nor UO_918 (O_918,N_29828,N_29088);
or UO_919 (O_919,N_29556,N_29258);
xnor UO_920 (O_920,N_29293,N_29834);
xnor UO_921 (O_921,N_29485,N_28843);
xnor UO_922 (O_922,N_29700,N_29678);
or UO_923 (O_923,N_29778,N_29419);
nor UO_924 (O_924,N_29685,N_29921);
and UO_925 (O_925,N_29455,N_29277);
or UO_926 (O_926,N_29074,N_29044);
or UO_927 (O_927,N_29696,N_28812);
or UO_928 (O_928,N_28917,N_29547);
xnor UO_929 (O_929,N_29263,N_29111);
nand UO_930 (O_930,N_29544,N_29627);
or UO_931 (O_931,N_28944,N_29798);
or UO_932 (O_932,N_29573,N_28867);
or UO_933 (O_933,N_29960,N_29962);
nor UO_934 (O_934,N_29876,N_29041);
nand UO_935 (O_935,N_28896,N_28827);
nor UO_936 (O_936,N_29396,N_29704);
and UO_937 (O_937,N_29878,N_29988);
nor UO_938 (O_938,N_29264,N_29682);
xor UO_939 (O_939,N_29080,N_29117);
and UO_940 (O_940,N_29309,N_29044);
nor UO_941 (O_941,N_29890,N_29672);
and UO_942 (O_942,N_28804,N_29559);
and UO_943 (O_943,N_29203,N_29748);
nor UO_944 (O_944,N_29206,N_29953);
nand UO_945 (O_945,N_29386,N_29675);
nand UO_946 (O_946,N_28812,N_29159);
or UO_947 (O_947,N_29202,N_29879);
xor UO_948 (O_948,N_29023,N_28874);
nor UO_949 (O_949,N_28849,N_29320);
or UO_950 (O_950,N_28892,N_28971);
nor UO_951 (O_951,N_29551,N_29485);
xor UO_952 (O_952,N_29872,N_28853);
nor UO_953 (O_953,N_28831,N_29079);
or UO_954 (O_954,N_29879,N_29421);
xor UO_955 (O_955,N_29058,N_29310);
and UO_956 (O_956,N_29767,N_29864);
nor UO_957 (O_957,N_29901,N_29834);
nor UO_958 (O_958,N_29532,N_29467);
or UO_959 (O_959,N_29118,N_29983);
nand UO_960 (O_960,N_29332,N_29498);
or UO_961 (O_961,N_29040,N_29724);
nor UO_962 (O_962,N_29999,N_28909);
nand UO_963 (O_963,N_29962,N_28801);
nand UO_964 (O_964,N_29888,N_29329);
and UO_965 (O_965,N_29450,N_29864);
and UO_966 (O_966,N_29918,N_29657);
or UO_967 (O_967,N_29075,N_29798);
xor UO_968 (O_968,N_29714,N_28863);
nor UO_969 (O_969,N_29010,N_28977);
nand UO_970 (O_970,N_29227,N_29046);
xnor UO_971 (O_971,N_29398,N_29955);
xnor UO_972 (O_972,N_29677,N_29873);
xnor UO_973 (O_973,N_29292,N_29754);
and UO_974 (O_974,N_28898,N_29127);
and UO_975 (O_975,N_29619,N_29284);
and UO_976 (O_976,N_29173,N_29130);
and UO_977 (O_977,N_29785,N_29614);
nand UO_978 (O_978,N_29618,N_29852);
nand UO_979 (O_979,N_28896,N_29977);
and UO_980 (O_980,N_29847,N_29845);
xnor UO_981 (O_981,N_29927,N_29899);
and UO_982 (O_982,N_28912,N_29222);
nand UO_983 (O_983,N_29597,N_29767);
nand UO_984 (O_984,N_29915,N_29964);
and UO_985 (O_985,N_29347,N_29671);
or UO_986 (O_986,N_29073,N_29705);
or UO_987 (O_987,N_29871,N_29539);
nor UO_988 (O_988,N_29021,N_29629);
nor UO_989 (O_989,N_29754,N_29923);
nor UO_990 (O_990,N_29551,N_28951);
and UO_991 (O_991,N_29675,N_29266);
nor UO_992 (O_992,N_28896,N_29613);
xor UO_993 (O_993,N_29454,N_29637);
or UO_994 (O_994,N_28947,N_29956);
nand UO_995 (O_995,N_29022,N_29542);
nor UO_996 (O_996,N_29880,N_29077);
and UO_997 (O_997,N_29526,N_29393);
and UO_998 (O_998,N_29663,N_29839);
nor UO_999 (O_999,N_29257,N_28914);
and UO_1000 (O_1000,N_29812,N_29070);
xnor UO_1001 (O_1001,N_29670,N_29219);
nor UO_1002 (O_1002,N_29238,N_28853);
nand UO_1003 (O_1003,N_29705,N_29774);
and UO_1004 (O_1004,N_28912,N_29878);
and UO_1005 (O_1005,N_29122,N_29161);
xor UO_1006 (O_1006,N_29778,N_29079);
or UO_1007 (O_1007,N_28961,N_29395);
xor UO_1008 (O_1008,N_29950,N_28876);
xor UO_1009 (O_1009,N_29122,N_29834);
xnor UO_1010 (O_1010,N_28888,N_29400);
nand UO_1011 (O_1011,N_29247,N_28812);
nor UO_1012 (O_1012,N_29186,N_29624);
or UO_1013 (O_1013,N_29173,N_29689);
and UO_1014 (O_1014,N_29387,N_29880);
and UO_1015 (O_1015,N_29287,N_29028);
xor UO_1016 (O_1016,N_29883,N_29321);
xor UO_1017 (O_1017,N_29122,N_28895);
and UO_1018 (O_1018,N_29953,N_28952);
nand UO_1019 (O_1019,N_29173,N_29094);
xnor UO_1020 (O_1020,N_29984,N_29451);
nand UO_1021 (O_1021,N_29144,N_29498);
nand UO_1022 (O_1022,N_29420,N_29134);
and UO_1023 (O_1023,N_29560,N_29360);
nor UO_1024 (O_1024,N_29521,N_29744);
or UO_1025 (O_1025,N_29037,N_29549);
xor UO_1026 (O_1026,N_29165,N_29927);
and UO_1027 (O_1027,N_29879,N_29888);
nor UO_1028 (O_1028,N_29150,N_29064);
nor UO_1029 (O_1029,N_29873,N_29867);
and UO_1030 (O_1030,N_28984,N_29032);
and UO_1031 (O_1031,N_29203,N_29222);
or UO_1032 (O_1032,N_29966,N_29669);
or UO_1033 (O_1033,N_29254,N_29143);
xnor UO_1034 (O_1034,N_29309,N_29032);
nand UO_1035 (O_1035,N_29920,N_29687);
nor UO_1036 (O_1036,N_29794,N_29947);
nor UO_1037 (O_1037,N_29507,N_29461);
or UO_1038 (O_1038,N_28981,N_29360);
nor UO_1039 (O_1039,N_29537,N_29199);
and UO_1040 (O_1040,N_29224,N_29360);
nand UO_1041 (O_1041,N_29280,N_29096);
or UO_1042 (O_1042,N_28869,N_28826);
and UO_1043 (O_1043,N_28953,N_28901);
nor UO_1044 (O_1044,N_29518,N_29532);
nand UO_1045 (O_1045,N_29414,N_28888);
or UO_1046 (O_1046,N_29321,N_29638);
and UO_1047 (O_1047,N_29725,N_29512);
nor UO_1048 (O_1048,N_29211,N_29587);
nand UO_1049 (O_1049,N_29983,N_29579);
xnor UO_1050 (O_1050,N_29262,N_29517);
or UO_1051 (O_1051,N_29449,N_29912);
xor UO_1052 (O_1052,N_28873,N_29845);
nand UO_1053 (O_1053,N_29925,N_29078);
nand UO_1054 (O_1054,N_28807,N_29940);
nor UO_1055 (O_1055,N_29781,N_29680);
nand UO_1056 (O_1056,N_29491,N_29782);
xnor UO_1057 (O_1057,N_29631,N_29067);
xnor UO_1058 (O_1058,N_29528,N_29615);
nand UO_1059 (O_1059,N_29010,N_29707);
nand UO_1060 (O_1060,N_28805,N_29195);
nand UO_1061 (O_1061,N_29990,N_29570);
nor UO_1062 (O_1062,N_29715,N_29788);
xor UO_1063 (O_1063,N_29044,N_29623);
nor UO_1064 (O_1064,N_29468,N_28875);
xnor UO_1065 (O_1065,N_29988,N_28969);
xnor UO_1066 (O_1066,N_29973,N_29873);
and UO_1067 (O_1067,N_29211,N_29512);
and UO_1068 (O_1068,N_29662,N_29799);
and UO_1069 (O_1069,N_29380,N_28844);
and UO_1070 (O_1070,N_28979,N_29059);
and UO_1071 (O_1071,N_28939,N_28870);
nand UO_1072 (O_1072,N_28856,N_29832);
nand UO_1073 (O_1073,N_29617,N_29953);
nor UO_1074 (O_1074,N_29154,N_29901);
nand UO_1075 (O_1075,N_29908,N_29684);
or UO_1076 (O_1076,N_29112,N_29982);
nor UO_1077 (O_1077,N_29214,N_29330);
nor UO_1078 (O_1078,N_29638,N_29703);
xnor UO_1079 (O_1079,N_29161,N_29969);
nand UO_1080 (O_1080,N_29284,N_29491);
nand UO_1081 (O_1081,N_29402,N_29479);
or UO_1082 (O_1082,N_29059,N_29487);
and UO_1083 (O_1083,N_29944,N_28869);
or UO_1084 (O_1084,N_28993,N_28844);
xnor UO_1085 (O_1085,N_29518,N_29341);
xor UO_1086 (O_1086,N_29702,N_29537);
xnor UO_1087 (O_1087,N_28923,N_29266);
or UO_1088 (O_1088,N_29157,N_29509);
nor UO_1089 (O_1089,N_29970,N_29690);
xor UO_1090 (O_1090,N_29730,N_29534);
and UO_1091 (O_1091,N_29998,N_29790);
or UO_1092 (O_1092,N_29719,N_29442);
or UO_1093 (O_1093,N_28995,N_29264);
nand UO_1094 (O_1094,N_29414,N_28960);
nand UO_1095 (O_1095,N_29978,N_28976);
or UO_1096 (O_1096,N_29536,N_29911);
and UO_1097 (O_1097,N_29116,N_29472);
nor UO_1098 (O_1098,N_29336,N_29159);
xor UO_1099 (O_1099,N_29524,N_28842);
nor UO_1100 (O_1100,N_28896,N_29904);
xnor UO_1101 (O_1101,N_29612,N_29958);
nor UO_1102 (O_1102,N_29234,N_29297);
nand UO_1103 (O_1103,N_29683,N_29298);
nor UO_1104 (O_1104,N_28846,N_29946);
or UO_1105 (O_1105,N_29877,N_29372);
xor UO_1106 (O_1106,N_29878,N_29331);
nand UO_1107 (O_1107,N_29874,N_28972);
nand UO_1108 (O_1108,N_29295,N_28932);
or UO_1109 (O_1109,N_28990,N_29604);
nand UO_1110 (O_1110,N_29698,N_29280);
or UO_1111 (O_1111,N_29017,N_29992);
and UO_1112 (O_1112,N_29784,N_28847);
xnor UO_1113 (O_1113,N_29739,N_29641);
xor UO_1114 (O_1114,N_29790,N_29668);
nor UO_1115 (O_1115,N_29147,N_29626);
and UO_1116 (O_1116,N_29223,N_28886);
nor UO_1117 (O_1117,N_29193,N_29464);
nand UO_1118 (O_1118,N_29947,N_29672);
and UO_1119 (O_1119,N_28810,N_29401);
nor UO_1120 (O_1120,N_28938,N_29478);
xor UO_1121 (O_1121,N_28867,N_29665);
or UO_1122 (O_1122,N_29478,N_29508);
xor UO_1123 (O_1123,N_29073,N_29404);
nor UO_1124 (O_1124,N_28889,N_29246);
or UO_1125 (O_1125,N_29431,N_29542);
nor UO_1126 (O_1126,N_29136,N_29624);
nand UO_1127 (O_1127,N_29624,N_29685);
or UO_1128 (O_1128,N_29028,N_28893);
or UO_1129 (O_1129,N_29660,N_29149);
xnor UO_1130 (O_1130,N_29395,N_29284);
xnor UO_1131 (O_1131,N_29040,N_29655);
nand UO_1132 (O_1132,N_29518,N_29732);
nor UO_1133 (O_1133,N_29329,N_29183);
nand UO_1134 (O_1134,N_29224,N_28961);
nor UO_1135 (O_1135,N_29656,N_29605);
nand UO_1136 (O_1136,N_29439,N_29173);
xnor UO_1137 (O_1137,N_28876,N_29241);
or UO_1138 (O_1138,N_29357,N_29480);
nor UO_1139 (O_1139,N_29296,N_29587);
nand UO_1140 (O_1140,N_29194,N_29708);
nand UO_1141 (O_1141,N_28912,N_29494);
or UO_1142 (O_1142,N_29911,N_29959);
nor UO_1143 (O_1143,N_29847,N_28932);
and UO_1144 (O_1144,N_29902,N_29197);
nand UO_1145 (O_1145,N_29282,N_29179);
nor UO_1146 (O_1146,N_29881,N_28889);
xor UO_1147 (O_1147,N_29950,N_29511);
or UO_1148 (O_1148,N_29065,N_29825);
xnor UO_1149 (O_1149,N_29222,N_28869);
and UO_1150 (O_1150,N_28846,N_29789);
xnor UO_1151 (O_1151,N_29039,N_28862);
nand UO_1152 (O_1152,N_29473,N_29556);
nand UO_1153 (O_1153,N_29815,N_29896);
or UO_1154 (O_1154,N_29466,N_29896);
xnor UO_1155 (O_1155,N_29220,N_29346);
or UO_1156 (O_1156,N_29163,N_29155);
nand UO_1157 (O_1157,N_28966,N_29198);
and UO_1158 (O_1158,N_29556,N_28887);
xnor UO_1159 (O_1159,N_29943,N_29775);
or UO_1160 (O_1160,N_28851,N_29312);
or UO_1161 (O_1161,N_28829,N_29069);
nor UO_1162 (O_1162,N_29895,N_28810);
nand UO_1163 (O_1163,N_29639,N_29538);
nand UO_1164 (O_1164,N_29136,N_29785);
and UO_1165 (O_1165,N_29700,N_29924);
or UO_1166 (O_1166,N_28972,N_29861);
nand UO_1167 (O_1167,N_29448,N_29320);
nor UO_1168 (O_1168,N_29077,N_29608);
nand UO_1169 (O_1169,N_29937,N_29911);
or UO_1170 (O_1170,N_28925,N_29219);
xnor UO_1171 (O_1171,N_29791,N_29434);
nand UO_1172 (O_1172,N_29691,N_29114);
or UO_1173 (O_1173,N_29897,N_29429);
or UO_1174 (O_1174,N_29076,N_29034);
or UO_1175 (O_1175,N_29643,N_28873);
nor UO_1176 (O_1176,N_29390,N_29772);
or UO_1177 (O_1177,N_29707,N_29104);
or UO_1178 (O_1178,N_29738,N_29476);
nand UO_1179 (O_1179,N_28967,N_29110);
nand UO_1180 (O_1180,N_29611,N_28841);
and UO_1181 (O_1181,N_29992,N_29573);
or UO_1182 (O_1182,N_29587,N_29907);
nor UO_1183 (O_1183,N_29035,N_29213);
nand UO_1184 (O_1184,N_29339,N_29697);
and UO_1185 (O_1185,N_29382,N_29799);
and UO_1186 (O_1186,N_29031,N_29805);
xnor UO_1187 (O_1187,N_29260,N_29631);
and UO_1188 (O_1188,N_29127,N_29202);
xnor UO_1189 (O_1189,N_29286,N_29255);
xnor UO_1190 (O_1190,N_29546,N_28900);
and UO_1191 (O_1191,N_28999,N_29513);
and UO_1192 (O_1192,N_28914,N_29309);
xor UO_1193 (O_1193,N_29004,N_29806);
nor UO_1194 (O_1194,N_29418,N_29794);
xnor UO_1195 (O_1195,N_29474,N_29607);
or UO_1196 (O_1196,N_29487,N_29081);
or UO_1197 (O_1197,N_29393,N_28808);
xor UO_1198 (O_1198,N_29761,N_29064);
nor UO_1199 (O_1199,N_29468,N_29932);
nand UO_1200 (O_1200,N_28829,N_28942);
and UO_1201 (O_1201,N_29809,N_29893);
xor UO_1202 (O_1202,N_29268,N_29847);
nand UO_1203 (O_1203,N_28878,N_29383);
nand UO_1204 (O_1204,N_29779,N_29236);
nor UO_1205 (O_1205,N_29678,N_29093);
xor UO_1206 (O_1206,N_29514,N_28929);
or UO_1207 (O_1207,N_29182,N_29609);
nor UO_1208 (O_1208,N_28842,N_28861);
or UO_1209 (O_1209,N_29650,N_29725);
and UO_1210 (O_1210,N_28842,N_28844);
xor UO_1211 (O_1211,N_29838,N_29789);
xor UO_1212 (O_1212,N_29677,N_29216);
nor UO_1213 (O_1213,N_29295,N_29335);
nand UO_1214 (O_1214,N_28850,N_29239);
or UO_1215 (O_1215,N_29306,N_29284);
or UO_1216 (O_1216,N_29618,N_29517);
and UO_1217 (O_1217,N_29913,N_29777);
nor UO_1218 (O_1218,N_29205,N_29222);
nor UO_1219 (O_1219,N_29553,N_29528);
or UO_1220 (O_1220,N_29974,N_29113);
or UO_1221 (O_1221,N_29364,N_29588);
nand UO_1222 (O_1222,N_29375,N_29430);
or UO_1223 (O_1223,N_29956,N_29302);
nand UO_1224 (O_1224,N_29631,N_29170);
nand UO_1225 (O_1225,N_29311,N_28877);
xnor UO_1226 (O_1226,N_29665,N_29123);
or UO_1227 (O_1227,N_28932,N_29089);
nand UO_1228 (O_1228,N_29445,N_29832);
nand UO_1229 (O_1229,N_29133,N_29333);
and UO_1230 (O_1230,N_29663,N_29580);
nand UO_1231 (O_1231,N_29445,N_29768);
and UO_1232 (O_1232,N_29357,N_29294);
nor UO_1233 (O_1233,N_28836,N_29022);
and UO_1234 (O_1234,N_29837,N_29259);
or UO_1235 (O_1235,N_29731,N_29943);
nand UO_1236 (O_1236,N_29243,N_29945);
nand UO_1237 (O_1237,N_29183,N_29908);
xnor UO_1238 (O_1238,N_29709,N_29060);
xor UO_1239 (O_1239,N_28810,N_29648);
nand UO_1240 (O_1240,N_29716,N_29575);
and UO_1241 (O_1241,N_29897,N_29631);
or UO_1242 (O_1242,N_29335,N_28908);
nor UO_1243 (O_1243,N_29145,N_29244);
and UO_1244 (O_1244,N_29312,N_29487);
and UO_1245 (O_1245,N_29637,N_29157);
and UO_1246 (O_1246,N_29338,N_29232);
nor UO_1247 (O_1247,N_28935,N_29843);
or UO_1248 (O_1248,N_29968,N_28962);
xnor UO_1249 (O_1249,N_29903,N_29350);
or UO_1250 (O_1250,N_29403,N_28953);
or UO_1251 (O_1251,N_29631,N_29866);
xnor UO_1252 (O_1252,N_29620,N_29208);
nor UO_1253 (O_1253,N_28818,N_29039);
or UO_1254 (O_1254,N_29029,N_29612);
and UO_1255 (O_1255,N_29459,N_29938);
and UO_1256 (O_1256,N_29197,N_29136);
nor UO_1257 (O_1257,N_29652,N_29228);
nor UO_1258 (O_1258,N_28936,N_28921);
nor UO_1259 (O_1259,N_29295,N_28914);
or UO_1260 (O_1260,N_28978,N_29654);
nand UO_1261 (O_1261,N_29949,N_29617);
nor UO_1262 (O_1262,N_29728,N_29066);
nor UO_1263 (O_1263,N_29827,N_29260);
nor UO_1264 (O_1264,N_29699,N_29123);
nor UO_1265 (O_1265,N_29789,N_29519);
or UO_1266 (O_1266,N_29859,N_29268);
nor UO_1267 (O_1267,N_29511,N_29790);
or UO_1268 (O_1268,N_29079,N_29207);
nor UO_1269 (O_1269,N_29896,N_29337);
nand UO_1270 (O_1270,N_29685,N_29534);
nor UO_1271 (O_1271,N_29741,N_29687);
nand UO_1272 (O_1272,N_29456,N_29077);
or UO_1273 (O_1273,N_29186,N_28954);
or UO_1274 (O_1274,N_29988,N_29054);
nor UO_1275 (O_1275,N_29795,N_29388);
or UO_1276 (O_1276,N_29802,N_29043);
or UO_1277 (O_1277,N_29748,N_29563);
nand UO_1278 (O_1278,N_29022,N_29418);
nor UO_1279 (O_1279,N_29712,N_29373);
xnor UO_1280 (O_1280,N_29041,N_29507);
and UO_1281 (O_1281,N_29093,N_29643);
and UO_1282 (O_1282,N_29189,N_29778);
or UO_1283 (O_1283,N_29082,N_29223);
or UO_1284 (O_1284,N_29846,N_29784);
xnor UO_1285 (O_1285,N_29065,N_28853);
nand UO_1286 (O_1286,N_29482,N_29071);
nor UO_1287 (O_1287,N_29070,N_29820);
nor UO_1288 (O_1288,N_29251,N_29941);
or UO_1289 (O_1289,N_29018,N_29097);
and UO_1290 (O_1290,N_29356,N_29234);
or UO_1291 (O_1291,N_29382,N_28980);
xnor UO_1292 (O_1292,N_29236,N_29844);
and UO_1293 (O_1293,N_29781,N_29793);
nand UO_1294 (O_1294,N_29394,N_29261);
and UO_1295 (O_1295,N_29117,N_28968);
nand UO_1296 (O_1296,N_29175,N_29481);
xnor UO_1297 (O_1297,N_29626,N_29703);
or UO_1298 (O_1298,N_29227,N_29102);
nand UO_1299 (O_1299,N_29163,N_29065);
xnor UO_1300 (O_1300,N_28907,N_29372);
or UO_1301 (O_1301,N_28822,N_28887);
xnor UO_1302 (O_1302,N_29832,N_29913);
xor UO_1303 (O_1303,N_29823,N_29332);
and UO_1304 (O_1304,N_29294,N_29227);
xnor UO_1305 (O_1305,N_29920,N_29561);
nand UO_1306 (O_1306,N_28809,N_29082);
nor UO_1307 (O_1307,N_29005,N_29637);
and UO_1308 (O_1308,N_28991,N_29182);
nor UO_1309 (O_1309,N_29302,N_29350);
nand UO_1310 (O_1310,N_29493,N_28810);
xnor UO_1311 (O_1311,N_29614,N_29899);
nand UO_1312 (O_1312,N_29671,N_28925);
nor UO_1313 (O_1313,N_29145,N_28935);
nor UO_1314 (O_1314,N_29166,N_29428);
or UO_1315 (O_1315,N_29416,N_29297);
xor UO_1316 (O_1316,N_28926,N_29130);
nand UO_1317 (O_1317,N_29717,N_28875);
nand UO_1318 (O_1318,N_29420,N_29212);
xor UO_1319 (O_1319,N_28825,N_28852);
nand UO_1320 (O_1320,N_29010,N_29816);
and UO_1321 (O_1321,N_29755,N_29167);
xnor UO_1322 (O_1322,N_29337,N_29394);
or UO_1323 (O_1323,N_29508,N_29976);
xor UO_1324 (O_1324,N_29809,N_29956);
and UO_1325 (O_1325,N_29544,N_29382);
nor UO_1326 (O_1326,N_29309,N_29027);
nor UO_1327 (O_1327,N_29995,N_29580);
nand UO_1328 (O_1328,N_29958,N_29733);
nor UO_1329 (O_1329,N_28892,N_28843);
and UO_1330 (O_1330,N_29069,N_29143);
and UO_1331 (O_1331,N_29637,N_29881);
and UO_1332 (O_1332,N_29542,N_29158);
and UO_1333 (O_1333,N_29546,N_29105);
nor UO_1334 (O_1334,N_29416,N_29964);
nand UO_1335 (O_1335,N_29296,N_29781);
nand UO_1336 (O_1336,N_29740,N_29073);
and UO_1337 (O_1337,N_29924,N_29073);
nand UO_1338 (O_1338,N_28990,N_28831);
xnor UO_1339 (O_1339,N_29066,N_29643);
or UO_1340 (O_1340,N_29785,N_28962);
and UO_1341 (O_1341,N_29157,N_29854);
nand UO_1342 (O_1342,N_29973,N_29827);
xnor UO_1343 (O_1343,N_29286,N_28918);
nand UO_1344 (O_1344,N_29308,N_29032);
and UO_1345 (O_1345,N_29548,N_29833);
nor UO_1346 (O_1346,N_29264,N_29496);
nor UO_1347 (O_1347,N_29329,N_29278);
nand UO_1348 (O_1348,N_29893,N_28942);
nor UO_1349 (O_1349,N_29075,N_29320);
and UO_1350 (O_1350,N_29768,N_28812);
and UO_1351 (O_1351,N_28824,N_29464);
and UO_1352 (O_1352,N_28818,N_29546);
xor UO_1353 (O_1353,N_29110,N_29461);
xor UO_1354 (O_1354,N_29313,N_29902);
and UO_1355 (O_1355,N_29698,N_29917);
or UO_1356 (O_1356,N_29051,N_29066);
and UO_1357 (O_1357,N_28866,N_29788);
nor UO_1358 (O_1358,N_29196,N_29999);
or UO_1359 (O_1359,N_29914,N_29500);
nor UO_1360 (O_1360,N_29048,N_28867);
and UO_1361 (O_1361,N_29541,N_29284);
nand UO_1362 (O_1362,N_29776,N_29910);
or UO_1363 (O_1363,N_29702,N_29921);
and UO_1364 (O_1364,N_28899,N_29406);
or UO_1365 (O_1365,N_29277,N_28967);
xor UO_1366 (O_1366,N_28914,N_29702);
or UO_1367 (O_1367,N_28859,N_29055);
xor UO_1368 (O_1368,N_29050,N_29224);
and UO_1369 (O_1369,N_28995,N_29187);
xor UO_1370 (O_1370,N_29930,N_29784);
nor UO_1371 (O_1371,N_29368,N_29720);
xnor UO_1372 (O_1372,N_29905,N_29322);
xor UO_1373 (O_1373,N_28949,N_29783);
xnor UO_1374 (O_1374,N_28809,N_29726);
nand UO_1375 (O_1375,N_29380,N_29622);
and UO_1376 (O_1376,N_29758,N_28955);
and UO_1377 (O_1377,N_29373,N_29749);
xnor UO_1378 (O_1378,N_29431,N_29674);
and UO_1379 (O_1379,N_29468,N_29092);
nand UO_1380 (O_1380,N_29977,N_29976);
and UO_1381 (O_1381,N_29332,N_29789);
xor UO_1382 (O_1382,N_29376,N_29787);
nand UO_1383 (O_1383,N_29887,N_29319);
xor UO_1384 (O_1384,N_29301,N_28963);
or UO_1385 (O_1385,N_29517,N_29202);
and UO_1386 (O_1386,N_29108,N_29531);
nand UO_1387 (O_1387,N_29770,N_29120);
nand UO_1388 (O_1388,N_29710,N_29814);
or UO_1389 (O_1389,N_29036,N_29627);
nand UO_1390 (O_1390,N_29388,N_29723);
xnor UO_1391 (O_1391,N_29775,N_29477);
and UO_1392 (O_1392,N_28993,N_29070);
nand UO_1393 (O_1393,N_29476,N_29642);
nand UO_1394 (O_1394,N_28804,N_29316);
xnor UO_1395 (O_1395,N_28801,N_29688);
and UO_1396 (O_1396,N_29299,N_29452);
and UO_1397 (O_1397,N_29327,N_29509);
and UO_1398 (O_1398,N_29899,N_28951);
nand UO_1399 (O_1399,N_29106,N_29159);
and UO_1400 (O_1400,N_29685,N_28816);
nand UO_1401 (O_1401,N_29818,N_29549);
nor UO_1402 (O_1402,N_29766,N_28901);
or UO_1403 (O_1403,N_29718,N_29522);
or UO_1404 (O_1404,N_29680,N_29182);
and UO_1405 (O_1405,N_29511,N_29827);
or UO_1406 (O_1406,N_29965,N_29506);
nor UO_1407 (O_1407,N_29241,N_29202);
or UO_1408 (O_1408,N_29480,N_29143);
xor UO_1409 (O_1409,N_28863,N_29207);
or UO_1410 (O_1410,N_29148,N_29437);
and UO_1411 (O_1411,N_29936,N_29449);
and UO_1412 (O_1412,N_28931,N_29291);
or UO_1413 (O_1413,N_29574,N_29637);
nor UO_1414 (O_1414,N_29242,N_29195);
nand UO_1415 (O_1415,N_29531,N_29824);
and UO_1416 (O_1416,N_29494,N_29937);
nand UO_1417 (O_1417,N_28908,N_29938);
nor UO_1418 (O_1418,N_29625,N_29758);
or UO_1419 (O_1419,N_29083,N_29915);
or UO_1420 (O_1420,N_29371,N_28869);
nor UO_1421 (O_1421,N_28811,N_29402);
nand UO_1422 (O_1422,N_29340,N_28902);
nor UO_1423 (O_1423,N_29505,N_29774);
xnor UO_1424 (O_1424,N_29499,N_29400);
xor UO_1425 (O_1425,N_29659,N_29693);
or UO_1426 (O_1426,N_29182,N_29816);
nor UO_1427 (O_1427,N_29372,N_29349);
and UO_1428 (O_1428,N_29930,N_29708);
or UO_1429 (O_1429,N_29388,N_28906);
and UO_1430 (O_1430,N_29834,N_29453);
nand UO_1431 (O_1431,N_29967,N_28999);
or UO_1432 (O_1432,N_29272,N_29507);
and UO_1433 (O_1433,N_29155,N_28811);
xnor UO_1434 (O_1434,N_29621,N_29117);
and UO_1435 (O_1435,N_29242,N_29619);
nand UO_1436 (O_1436,N_28844,N_29201);
or UO_1437 (O_1437,N_29549,N_29517);
or UO_1438 (O_1438,N_28923,N_29054);
nor UO_1439 (O_1439,N_29656,N_29957);
and UO_1440 (O_1440,N_29255,N_29011);
xor UO_1441 (O_1441,N_29372,N_29723);
xnor UO_1442 (O_1442,N_29587,N_29692);
or UO_1443 (O_1443,N_29668,N_29949);
nor UO_1444 (O_1444,N_29446,N_29557);
nor UO_1445 (O_1445,N_29910,N_29071);
xor UO_1446 (O_1446,N_29676,N_29400);
and UO_1447 (O_1447,N_29275,N_29892);
or UO_1448 (O_1448,N_29611,N_29237);
xnor UO_1449 (O_1449,N_29512,N_28827);
and UO_1450 (O_1450,N_29493,N_28966);
nand UO_1451 (O_1451,N_29738,N_29576);
nor UO_1452 (O_1452,N_29362,N_29824);
or UO_1453 (O_1453,N_29528,N_29602);
or UO_1454 (O_1454,N_29417,N_29502);
or UO_1455 (O_1455,N_28979,N_29369);
and UO_1456 (O_1456,N_29749,N_29216);
or UO_1457 (O_1457,N_28864,N_29588);
nor UO_1458 (O_1458,N_29911,N_29291);
or UO_1459 (O_1459,N_29904,N_29798);
and UO_1460 (O_1460,N_28963,N_28860);
nand UO_1461 (O_1461,N_29655,N_29785);
xnor UO_1462 (O_1462,N_29655,N_28889);
or UO_1463 (O_1463,N_29189,N_29828);
xnor UO_1464 (O_1464,N_28842,N_29604);
xnor UO_1465 (O_1465,N_29528,N_28934);
or UO_1466 (O_1466,N_28818,N_29805);
xnor UO_1467 (O_1467,N_29665,N_29994);
or UO_1468 (O_1468,N_29165,N_29848);
nand UO_1469 (O_1469,N_29916,N_28969);
xnor UO_1470 (O_1470,N_29394,N_29947);
nand UO_1471 (O_1471,N_28901,N_28939);
nand UO_1472 (O_1472,N_28945,N_29559);
and UO_1473 (O_1473,N_28848,N_29007);
or UO_1474 (O_1474,N_29439,N_29433);
xnor UO_1475 (O_1475,N_29031,N_29409);
nand UO_1476 (O_1476,N_29652,N_28961);
nor UO_1477 (O_1477,N_29636,N_28896);
nor UO_1478 (O_1478,N_29421,N_29782);
or UO_1479 (O_1479,N_29513,N_29376);
and UO_1480 (O_1480,N_29712,N_29967);
and UO_1481 (O_1481,N_29667,N_29974);
nor UO_1482 (O_1482,N_29583,N_28976);
or UO_1483 (O_1483,N_29855,N_28858);
nand UO_1484 (O_1484,N_28886,N_28842);
xnor UO_1485 (O_1485,N_28878,N_29872);
nand UO_1486 (O_1486,N_29458,N_29672);
xor UO_1487 (O_1487,N_29932,N_29608);
and UO_1488 (O_1488,N_29246,N_28955);
or UO_1489 (O_1489,N_29215,N_29521);
xnor UO_1490 (O_1490,N_29351,N_29496);
nor UO_1491 (O_1491,N_28868,N_29900);
and UO_1492 (O_1492,N_29770,N_29714);
xor UO_1493 (O_1493,N_29056,N_29183);
xor UO_1494 (O_1494,N_28965,N_29143);
nand UO_1495 (O_1495,N_29897,N_29438);
or UO_1496 (O_1496,N_29150,N_29355);
or UO_1497 (O_1497,N_29537,N_29374);
and UO_1498 (O_1498,N_29308,N_29902);
nor UO_1499 (O_1499,N_29239,N_28955);
or UO_1500 (O_1500,N_29803,N_29122);
and UO_1501 (O_1501,N_29139,N_29707);
or UO_1502 (O_1502,N_28934,N_29415);
nand UO_1503 (O_1503,N_28870,N_29378);
nand UO_1504 (O_1504,N_29912,N_29151);
nand UO_1505 (O_1505,N_29923,N_29915);
xnor UO_1506 (O_1506,N_29851,N_29734);
xnor UO_1507 (O_1507,N_29150,N_29547);
nor UO_1508 (O_1508,N_29064,N_29687);
nand UO_1509 (O_1509,N_29648,N_29327);
or UO_1510 (O_1510,N_29562,N_29168);
or UO_1511 (O_1511,N_29007,N_29400);
and UO_1512 (O_1512,N_29356,N_28930);
and UO_1513 (O_1513,N_29962,N_29295);
or UO_1514 (O_1514,N_28996,N_29730);
and UO_1515 (O_1515,N_29464,N_29789);
or UO_1516 (O_1516,N_29016,N_29391);
or UO_1517 (O_1517,N_29723,N_29277);
nor UO_1518 (O_1518,N_29849,N_29361);
nand UO_1519 (O_1519,N_28843,N_29545);
and UO_1520 (O_1520,N_28830,N_29418);
nand UO_1521 (O_1521,N_29378,N_28893);
or UO_1522 (O_1522,N_29397,N_29464);
nor UO_1523 (O_1523,N_29979,N_29387);
and UO_1524 (O_1524,N_29214,N_28966);
or UO_1525 (O_1525,N_29176,N_29810);
or UO_1526 (O_1526,N_29075,N_29392);
xnor UO_1527 (O_1527,N_28966,N_29715);
and UO_1528 (O_1528,N_29236,N_29885);
or UO_1529 (O_1529,N_28843,N_28936);
nand UO_1530 (O_1530,N_29720,N_29599);
nand UO_1531 (O_1531,N_29135,N_29456);
or UO_1532 (O_1532,N_29538,N_29106);
xor UO_1533 (O_1533,N_29764,N_29236);
nor UO_1534 (O_1534,N_28826,N_29113);
and UO_1535 (O_1535,N_29605,N_29331);
nand UO_1536 (O_1536,N_29069,N_28821);
nor UO_1537 (O_1537,N_28949,N_29426);
nor UO_1538 (O_1538,N_29375,N_28818);
xnor UO_1539 (O_1539,N_29558,N_29035);
or UO_1540 (O_1540,N_29228,N_29916);
nor UO_1541 (O_1541,N_29783,N_29690);
nor UO_1542 (O_1542,N_28953,N_29864);
or UO_1543 (O_1543,N_29598,N_29135);
and UO_1544 (O_1544,N_29518,N_29543);
nor UO_1545 (O_1545,N_29064,N_29564);
nor UO_1546 (O_1546,N_29089,N_29251);
nand UO_1547 (O_1547,N_29412,N_29017);
nand UO_1548 (O_1548,N_29175,N_29619);
or UO_1549 (O_1549,N_28880,N_29264);
nand UO_1550 (O_1550,N_29300,N_28865);
xnor UO_1551 (O_1551,N_29606,N_29088);
and UO_1552 (O_1552,N_29779,N_29935);
or UO_1553 (O_1553,N_28835,N_29135);
and UO_1554 (O_1554,N_29379,N_29886);
xnor UO_1555 (O_1555,N_29956,N_29111);
nand UO_1556 (O_1556,N_29087,N_29546);
or UO_1557 (O_1557,N_29102,N_29916);
nor UO_1558 (O_1558,N_29758,N_29321);
and UO_1559 (O_1559,N_29082,N_28825);
nor UO_1560 (O_1560,N_29976,N_28962);
nand UO_1561 (O_1561,N_29613,N_29334);
and UO_1562 (O_1562,N_28852,N_28873);
nor UO_1563 (O_1563,N_29341,N_28834);
or UO_1564 (O_1564,N_29417,N_29115);
and UO_1565 (O_1565,N_29570,N_29411);
and UO_1566 (O_1566,N_29856,N_29236);
and UO_1567 (O_1567,N_28836,N_29523);
nand UO_1568 (O_1568,N_29610,N_29350);
nand UO_1569 (O_1569,N_29218,N_29869);
xor UO_1570 (O_1570,N_29966,N_29235);
nand UO_1571 (O_1571,N_28984,N_29199);
nor UO_1572 (O_1572,N_29792,N_28822);
or UO_1573 (O_1573,N_29201,N_29969);
xnor UO_1574 (O_1574,N_29737,N_29147);
xor UO_1575 (O_1575,N_29177,N_29653);
xnor UO_1576 (O_1576,N_28865,N_29375);
nor UO_1577 (O_1577,N_29072,N_28853);
nand UO_1578 (O_1578,N_29144,N_28967);
nor UO_1579 (O_1579,N_29908,N_29490);
or UO_1580 (O_1580,N_29127,N_28988);
and UO_1581 (O_1581,N_29442,N_29778);
and UO_1582 (O_1582,N_29500,N_28933);
nor UO_1583 (O_1583,N_29448,N_29558);
nor UO_1584 (O_1584,N_29870,N_29531);
xor UO_1585 (O_1585,N_29358,N_29494);
xnor UO_1586 (O_1586,N_29067,N_29132);
nor UO_1587 (O_1587,N_29211,N_29037);
or UO_1588 (O_1588,N_29107,N_29647);
nand UO_1589 (O_1589,N_29934,N_29397);
xnor UO_1590 (O_1590,N_29742,N_29886);
or UO_1591 (O_1591,N_29990,N_29478);
and UO_1592 (O_1592,N_29585,N_29266);
and UO_1593 (O_1593,N_29530,N_28818);
xnor UO_1594 (O_1594,N_29384,N_29802);
xnor UO_1595 (O_1595,N_29237,N_29988);
nand UO_1596 (O_1596,N_29952,N_29520);
or UO_1597 (O_1597,N_29804,N_29617);
or UO_1598 (O_1598,N_29434,N_29413);
or UO_1599 (O_1599,N_29265,N_29979);
and UO_1600 (O_1600,N_29383,N_28984);
and UO_1601 (O_1601,N_29299,N_29891);
or UO_1602 (O_1602,N_29492,N_29183);
nand UO_1603 (O_1603,N_28879,N_29256);
nand UO_1604 (O_1604,N_29396,N_29058);
nand UO_1605 (O_1605,N_29433,N_29871);
and UO_1606 (O_1606,N_29522,N_29616);
nor UO_1607 (O_1607,N_29989,N_28992);
or UO_1608 (O_1608,N_28973,N_29267);
nor UO_1609 (O_1609,N_29255,N_28881);
nor UO_1610 (O_1610,N_29929,N_29108);
nor UO_1611 (O_1611,N_29458,N_29104);
xor UO_1612 (O_1612,N_29318,N_29088);
or UO_1613 (O_1613,N_28886,N_29396);
nand UO_1614 (O_1614,N_28892,N_29426);
nand UO_1615 (O_1615,N_29647,N_29885);
nand UO_1616 (O_1616,N_28927,N_28929);
nand UO_1617 (O_1617,N_29321,N_29028);
or UO_1618 (O_1618,N_29671,N_28998);
and UO_1619 (O_1619,N_29698,N_29910);
nor UO_1620 (O_1620,N_28851,N_29778);
and UO_1621 (O_1621,N_29088,N_28948);
xor UO_1622 (O_1622,N_29939,N_29730);
xnor UO_1623 (O_1623,N_29857,N_29184);
or UO_1624 (O_1624,N_29339,N_29628);
nor UO_1625 (O_1625,N_29818,N_29053);
or UO_1626 (O_1626,N_29539,N_29683);
and UO_1627 (O_1627,N_28836,N_29300);
xor UO_1628 (O_1628,N_29469,N_28923);
nand UO_1629 (O_1629,N_29029,N_29493);
nand UO_1630 (O_1630,N_28860,N_29418);
and UO_1631 (O_1631,N_29700,N_29190);
and UO_1632 (O_1632,N_29145,N_29855);
or UO_1633 (O_1633,N_29314,N_29180);
nor UO_1634 (O_1634,N_29607,N_29790);
or UO_1635 (O_1635,N_28906,N_29956);
nor UO_1636 (O_1636,N_29829,N_29025);
nor UO_1637 (O_1637,N_28980,N_29562);
xnor UO_1638 (O_1638,N_29118,N_29277);
or UO_1639 (O_1639,N_29518,N_29101);
xnor UO_1640 (O_1640,N_29809,N_29456);
or UO_1641 (O_1641,N_29392,N_29669);
or UO_1642 (O_1642,N_29290,N_28971);
and UO_1643 (O_1643,N_28933,N_29113);
and UO_1644 (O_1644,N_28860,N_29977);
and UO_1645 (O_1645,N_29702,N_29299);
nor UO_1646 (O_1646,N_29594,N_28965);
or UO_1647 (O_1647,N_29461,N_29838);
xor UO_1648 (O_1648,N_29062,N_29856);
nor UO_1649 (O_1649,N_28935,N_28836);
nand UO_1650 (O_1650,N_29116,N_29695);
xor UO_1651 (O_1651,N_28922,N_29861);
nand UO_1652 (O_1652,N_28887,N_29768);
xor UO_1653 (O_1653,N_29376,N_29382);
nand UO_1654 (O_1654,N_28825,N_29067);
and UO_1655 (O_1655,N_28807,N_29515);
nand UO_1656 (O_1656,N_29146,N_29825);
nor UO_1657 (O_1657,N_29245,N_28899);
xnor UO_1658 (O_1658,N_29394,N_29949);
xnor UO_1659 (O_1659,N_29014,N_29941);
or UO_1660 (O_1660,N_29747,N_29172);
xor UO_1661 (O_1661,N_29901,N_29209);
or UO_1662 (O_1662,N_29838,N_29228);
xor UO_1663 (O_1663,N_28994,N_29670);
xor UO_1664 (O_1664,N_29133,N_29126);
xor UO_1665 (O_1665,N_29514,N_28927);
and UO_1666 (O_1666,N_29927,N_29573);
xnor UO_1667 (O_1667,N_29224,N_29532);
nand UO_1668 (O_1668,N_29609,N_29617);
or UO_1669 (O_1669,N_29186,N_29248);
and UO_1670 (O_1670,N_28813,N_29852);
or UO_1671 (O_1671,N_29232,N_29443);
nand UO_1672 (O_1672,N_29325,N_29729);
nor UO_1673 (O_1673,N_29281,N_29213);
and UO_1674 (O_1674,N_29559,N_28839);
or UO_1675 (O_1675,N_29818,N_29522);
nand UO_1676 (O_1676,N_29714,N_29917);
nand UO_1677 (O_1677,N_29213,N_29461);
nor UO_1678 (O_1678,N_29783,N_28896);
xnor UO_1679 (O_1679,N_29004,N_29950);
and UO_1680 (O_1680,N_29868,N_29291);
nor UO_1681 (O_1681,N_28813,N_29229);
and UO_1682 (O_1682,N_29405,N_29518);
nor UO_1683 (O_1683,N_29116,N_29750);
and UO_1684 (O_1684,N_29445,N_29814);
xor UO_1685 (O_1685,N_28983,N_28965);
xnor UO_1686 (O_1686,N_29325,N_29174);
and UO_1687 (O_1687,N_29573,N_28882);
or UO_1688 (O_1688,N_29304,N_29523);
nand UO_1689 (O_1689,N_29418,N_29143);
and UO_1690 (O_1690,N_29818,N_29099);
or UO_1691 (O_1691,N_29784,N_29534);
or UO_1692 (O_1692,N_29773,N_29851);
or UO_1693 (O_1693,N_29901,N_28860);
and UO_1694 (O_1694,N_29961,N_29689);
or UO_1695 (O_1695,N_29669,N_29461);
and UO_1696 (O_1696,N_29645,N_29847);
and UO_1697 (O_1697,N_29145,N_29033);
xnor UO_1698 (O_1698,N_29444,N_29284);
nor UO_1699 (O_1699,N_29121,N_29524);
nand UO_1700 (O_1700,N_29126,N_29472);
nand UO_1701 (O_1701,N_28914,N_29556);
or UO_1702 (O_1702,N_29803,N_28911);
or UO_1703 (O_1703,N_29070,N_29635);
nand UO_1704 (O_1704,N_29005,N_28988);
xnor UO_1705 (O_1705,N_28974,N_29566);
nor UO_1706 (O_1706,N_29218,N_29913);
xnor UO_1707 (O_1707,N_29493,N_29448);
nor UO_1708 (O_1708,N_29123,N_28861);
xor UO_1709 (O_1709,N_28988,N_29870);
or UO_1710 (O_1710,N_29976,N_29233);
nand UO_1711 (O_1711,N_29570,N_29714);
or UO_1712 (O_1712,N_29684,N_29139);
nor UO_1713 (O_1713,N_29898,N_29503);
nor UO_1714 (O_1714,N_29354,N_28804);
nand UO_1715 (O_1715,N_29835,N_28942);
nand UO_1716 (O_1716,N_28849,N_29558);
xnor UO_1717 (O_1717,N_29563,N_29842);
or UO_1718 (O_1718,N_29200,N_29441);
or UO_1719 (O_1719,N_29968,N_29005);
nor UO_1720 (O_1720,N_29492,N_29969);
or UO_1721 (O_1721,N_29490,N_29401);
and UO_1722 (O_1722,N_29971,N_29758);
nor UO_1723 (O_1723,N_29614,N_29228);
nand UO_1724 (O_1724,N_29740,N_29788);
and UO_1725 (O_1725,N_29356,N_29027);
nor UO_1726 (O_1726,N_29081,N_29773);
nand UO_1727 (O_1727,N_29055,N_29932);
xor UO_1728 (O_1728,N_29000,N_29396);
and UO_1729 (O_1729,N_29141,N_29235);
or UO_1730 (O_1730,N_29027,N_29538);
nand UO_1731 (O_1731,N_29009,N_29573);
or UO_1732 (O_1732,N_29728,N_29752);
or UO_1733 (O_1733,N_29726,N_28808);
nor UO_1734 (O_1734,N_28886,N_29863);
xor UO_1735 (O_1735,N_29428,N_29918);
and UO_1736 (O_1736,N_29865,N_29549);
nor UO_1737 (O_1737,N_28910,N_29139);
xor UO_1738 (O_1738,N_29597,N_29280);
and UO_1739 (O_1739,N_29441,N_29714);
nand UO_1740 (O_1740,N_29333,N_29515);
and UO_1741 (O_1741,N_29595,N_29309);
nor UO_1742 (O_1742,N_28959,N_29025);
nand UO_1743 (O_1743,N_29203,N_29443);
or UO_1744 (O_1744,N_29150,N_29484);
nor UO_1745 (O_1745,N_29787,N_29210);
or UO_1746 (O_1746,N_29986,N_29067);
nor UO_1747 (O_1747,N_29291,N_29558);
or UO_1748 (O_1748,N_29710,N_29439);
nand UO_1749 (O_1749,N_29045,N_28833);
nand UO_1750 (O_1750,N_29411,N_29888);
or UO_1751 (O_1751,N_29016,N_29144);
xor UO_1752 (O_1752,N_29397,N_29275);
nand UO_1753 (O_1753,N_29687,N_29586);
and UO_1754 (O_1754,N_29358,N_29473);
and UO_1755 (O_1755,N_29406,N_29547);
xnor UO_1756 (O_1756,N_29124,N_29988);
nor UO_1757 (O_1757,N_29452,N_29252);
nor UO_1758 (O_1758,N_28968,N_29919);
or UO_1759 (O_1759,N_29514,N_29079);
nor UO_1760 (O_1760,N_29957,N_29834);
nand UO_1761 (O_1761,N_28835,N_29339);
and UO_1762 (O_1762,N_29352,N_29250);
and UO_1763 (O_1763,N_29520,N_29369);
xor UO_1764 (O_1764,N_29796,N_29414);
nand UO_1765 (O_1765,N_28883,N_28885);
nor UO_1766 (O_1766,N_29617,N_28934);
xor UO_1767 (O_1767,N_29023,N_29185);
nand UO_1768 (O_1768,N_29893,N_28890);
or UO_1769 (O_1769,N_29948,N_29331);
nand UO_1770 (O_1770,N_28894,N_29343);
xor UO_1771 (O_1771,N_28961,N_29894);
nor UO_1772 (O_1772,N_28921,N_29847);
and UO_1773 (O_1773,N_29845,N_29065);
xor UO_1774 (O_1774,N_29908,N_29530);
nand UO_1775 (O_1775,N_29969,N_29913);
and UO_1776 (O_1776,N_29611,N_29931);
xor UO_1777 (O_1777,N_29205,N_29413);
nand UO_1778 (O_1778,N_29851,N_29639);
nand UO_1779 (O_1779,N_29093,N_29400);
and UO_1780 (O_1780,N_29590,N_29612);
xnor UO_1781 (O_1781,N_28830,N_28824);
or UO_1782 (O_1782,N_29502,N_29872);
nor UO_1783 (O_1783,N_29487,N_29592);
or UO_1784 (O_1784,N_29778,N_29559);
nor UO_1785 (O_1785,N_29573,N_29289);
xor UO_1786 (O_1786,N_29591,N_29187);
xnor UO_1787 (O_1787,N_28803,N_29019);
nor UO_1788 (O_1788,N_29691,N_29374);
nand UO_1789 (O_1789,N_28822,N_29084);
xor UO_1790 (O_1790,N_29663,N_29856);
xnor UO_1791 (O_1791,N_29183,N_29897);
xor UO_1792 (O_1792,N_29972,N_29937);
xor UO_1793 (O_1793,N_29161,N_29780);
xnor UO_1794 (O_1794,N_28888,N_29071);
nor UO_1795 (O_1795,N_29804,N_29153);
nor UO_1796 (O_1796,N_29624,N_28992);
nor UO_1797 (O_1797,N_28882,N_29927);
nand UO_1798 (O_1798,N_29515,N_29546);
xor UO_1799 (O_1799,N_29656,N_28842);
or UO_1800 (O_1800,N_28895,N_29732);
nor UO_1801 (O_1801,N_29269,N_29343);
or UO_1802 (O_1802,N_29256,N_29659);
nor UO_1803 (O_1803,N_29026,N_29723);
nand UO_1804 (O_1804,N_29167,N_29111);
xor UO_1805 (O_1805,N_28923,N_29556);
nand UO_1806 (O_1806,N_29720,N_29752);
xnor UO_1807 (O_1807,N_29189,N_29388);
nor UO_1808 (O_1808,N_29749,N_29879);
or UO_1809 (O_1809,N_29232,N_28912);
nor UO_1810 (O_1810,N_29200,N_29608);
nor UO_1811 (O_1811,N_29562,N_29815);
xor UO_1812 (O_1812,N_29979,N_28967);
and UO_1813 (O_1813,N_28894,N_29769);
nand UO_1814 (O_1814,N_29685,N_29946);
or UO_1815 (O_1815,N_29663,N_28980);
xor UO_1816 (O_1816,N_29357,N_29121);
or UO_1817 (O_1817,N_29269,N_29597);
nor UO_1818 (O_1818,N_29653,N_29758);
nand UO_1819 (O_1819,N_29145,N_29714);
nor UO_1820 (O_1820,N_29575,N_28909);
nor UO_1821 (O_1821,N_29723,N_28947);
and UO_1822 (O_1822,N_28926,N_28966);
nand UO_1823 (O_1823,N_29120,N_29640);
nand UO_1824 (O_1824,N_29715,N_29701);
and UO_1825 (O_1825,N_29564,N_29806);
nand UO_1826 (O_1826,N_29416,N_29568);
nand UO_1827 (O_1827,N_28943,N_29934);
nor UO_1828 (O_1828,N_29207,N_29433);
nor UO_1829 (O_1829,N_29239,N_28846);
and UO_1830 (O_1830,N_28972,N_29517);
xnor UO_1831 (O_1831,N_29745,N_29280);
and UO_1832 (O_1832,N_29114,N_29167);
nand UO_1833 (O_1833,N_29330,N_29360);
or UO_1834 (O_1834,N_29248,N_29552);
xor UO_1835 (O_1835,N_29765,N_29997);
and UO_1836 (O_1836,N_28893,N_28814);
nor UO_1837 (O_1837,N_29251,N_29579);
nand UO_1838 (O_1838,N_29708,N_29776);
nand UO_1839 (O_1839,N_29319,N_29333);
or UO_1840 (O_1840,N_29031,N_28952);
nand UO_1841 (O_1841,N_29670,N_28962);
xnor UO_1842 (O_1842,N_29906,N_29200);
xnor UO_1843 (O_1843,N_29839,N_28867);
or UO_1844 (O_1844,N_29437,N_29780);
nand UO_1845 (O_1845,N_29837,N_29372);
xor UO_1846 (O_1846,N_29127,N_29985);
or UO_1847 (O_1847,N_29109,N_29582);
xor UO_1848 (O_1848,N_28871,N_29592);
nand UO_1849 (O_1849,N_29864,N_29636);
nor UO_1850 (O_1850,N_29789,N_29834);
or UO_1851 (O_1851,N_29925,N_29865);
and UO_1852 (O_1852,N_29328,N_29893);
and UO_1853 (O_1853,N_29646,N_29243);
nor UO_1854 (O_1854,N_29188,N_29371);
or UO_1855 (O_1855,N_29930,N_29923);
nand UO_1856 (O_1856,N_29878,N_29372);
nor UO_1857 (O_1857,N_28929,N_28860);
nand UO_1858 (O_1858,N_29559,N_29372);
or UO_1859 (O_1859,N_29882,N_29010);
and UO_1860 (O_1860,N_29950,N_29912);
or UO_1861 (O_1861,N_29515,N_28924);
nor UO_1862 (O_1862,N_29073,N_29463);
and UO_1863 (O_1863,N_28996,N_28901);
xor UO_1864 (O_1864,N_29564,N_29396);
or UO_1865 (O_1865,N_29824,N_29092);
nand UO_1866 (O_1866,N_29163,N_29649);
nand UO_1867 (O_1867,N_28994,N_29675);
or UO_1868 (O_1868,N_29081,N_29855);
and UO_1869 (O_1869,N_29597,N_29318);
and UO_1870 (O_1870,N_29316,N_29177);
and UO_1871 (O_1871,N_29519,N_29551);
nor UO_1872 (O_1872,N_29842,N_29368);
xnor UO_1873 (O_1873,N_29589,N_29940);
and UO_1874 (O_1874,N_29313,N_29973);
and UO_1875 (O_1875,N_29116,N_29100);
xnor UO_1876 (O_1876,N_29731,N_29479);
nor UO_1877 (O_1877,N_29450,N_28904);
or UO_1878 (O_1878,N_29233,N_29106);
nand UO_1879 (O_1879,N_29513,N_29873);
nand UO_1880 (O_1880,N_28901,N_29603);
and UO_1881 (O_1881,N_29977,N_28917);
nand UO_1882 (O_1882,N_29909,N_29076);
nand UO_1883 (O_1883,N_29692,N_29643);
and UO_1884 (O_1884,N_29415,N_29814);
or UO_1885 (O_1885,N_29054,N_29731);
nor UO_1886 (O_1886,N_29726,N_29221);
or UO_1887 (O_1887,N_29999,N_29770);
nand UO_1888 (O_1888,N_29693,N_28868);
and UO_1889 (O_1889,N_28944,N_29435);
nor UO_1890 (O_1890,N_29180,N_29254);
nor UO_1891 (O_1891,N_29848,N_29025);
xnor UO_1892 (O_1892,N_29510,N_29720);
nor UO_1893 (O_1893,N_29696,N_29456);
nand UO_1894 (O_1894,N_29914,N_29016);
nand UO_1895 (O_1895,N_29451,N_29247);
nor UO_1896 (O_1896,N_29413,N_29451);
nand UO_1897 (O_1897,N_29219,N_29955);
or UO_1898 (O_1898,N_29544,N_28978);
and UO_1899 (O_1899,N_29595,N_29467);
nand UO_1900 (O_1900,N_29524,N_29243);
nor UO_1901 (O_1901,N_28817,N_29929);
nor UO_1902 (O_1902,N_28996,N_29842);
or UO_1903 (O_1903,N_29077,N_29791);
nor UO_1904 (O_1904,N_29943,N_29104);
nor UO_1905 (O_1905,N_28972,N_29476);
xor UO_1906 (O_1906,N_29730,N_29083);
nor UO_1907 (O_1907,N_29991,N_29872);
nand UO_1908 (O_1908,N_29288,N_28952);
nor UO_1909 (O_1909,N_29143,N_29552);
xor UO_1910 (O_1910,N_28905,N_29857);
nor UO_1911 (O_1911,N_29048,N_29479);
or UO_1912 (O_1912,N_28831,N_29826);
xnor UO_1913 (O_1913,N_29141,N_29758);
or UO_1914 (O_1914,N_29598,N_28800);
or UO_1915 (O_1915,N_29335,N_29926);
xor UO_1916 (O_1916,N_29087,N_28804);
nand UO_1917 (O_1917,N_29621,N_29740);
and UO_1918 (O_1918,N_29939,N_28907);
nor UO_1919 (O_1919,N_28888,N_29472);
and UO_1920 (O_1920,N_28991,N_29003);
xor UO_1921 (O_1921,N_29182,N_29657);
nor UO_1922 (O_1922,N_28901,N_29495);
and UO_1923 (O_1923,N_29657,N_29990);
or UO_1924 (O_1924,N_29648,N_28889);
nor UO_1925 (O_1925,N_29066,N_29846);
and UO_1926 (O_1926,N_29361,N_29078);
and UO_1927 (O_1927,N_29513,N_29743);
nor UO_1928 (O_1928,N_28933,N_29810);
xnor UO_1929 (O_1929,N_28842,N_29950);
nand UO_1930 (O_1930,N_29112,N_29971);
or UO_1931 (O_1931,N_29451,N_29721);
nor UO_1932 (O_1932,N_29089,N_29799);
nor UO_1933 (O_1933,N_29436,N_29081);
xor UO_1934 (O_1934,N_29845,N_29310);
or UO_1935 (O_1935,N_29187,N_29946);
and UO_1936 (O_1936,N_29815,N_28850);
and UO_1937 (O_1937,N_29940,N_29468);
xor UO_1938 (O_1938,N_29096,N_29810);
and UO_1939 (O_1939,N_29670,N_28801);
xor UO_1940 (O_1940,N_29421,N_29201);
or UO_1941 (O_1941,N_28825,N_29018);
xor UO_1942 (O_1942,N_29162,N_29582);
or UO_1943 (O_1943,N_28855,N_29758);
and UO_1944 (O_1944,N_29850,N_29891);
nand UO_1945 (O_1945,N_29895,N_29233);
or UO_1946 (O_1946,N_29316,N_29360);
or UO_1947 (O_1947,N_29810,N_29634);
nand UO_1948 (O_1948,N_29599,N_29561);
and UO_1949 (O_1949,N_29156,N_29704);
or UO_1950 (O_1950,N_29575,N_29840);
and UO_1951 (O_1951,N_29875,N_29791);
or UO_1952 (O_1952,N_29111,N_29593);
nor UO_1953 (O_1953,N_29074,N_29884);
nor UO_1954 (O_1954,N_29195,N_28927);
or UO_1955 (O_1955,N_29833,N_29347);
or UO_1956 (O_1956,N_29976,N_29943);
or UO_1957 (O_1957,N_29114,N_29132);
or UO_1958 (O_1958,N_29333,N_29974);
nor UO_1959 (O_1959,N_28940,N_29031);
nor UO_1960 (O_1960,N_29457,N_29090);
nor UO_1961 (O_1961,N_29063,N_29994);
and UO_1962 (O_1962,N_29773,N_29230);
xor UO_1963 (O_1963,N_28979,N_29432);
nand UO_1964 (O_1964,N_29723,N_28839);
or UO_1965 (O_1965,N_29893,N_29251);
nor UO_1966 (O_1966,N_29640,N_29571);
nor UO_1967 (O_1967,N_28959,N_29845);
and UO_1968 (O_1968,N_29317,N_29238);
and UO_1969 (O_1969,N_29107,N_29901);
nor UO_1970 (O_1970,N_29791,N_29232);
nor UO_1971 (O_1971,N_29489,N_29591);
nor UO_1972 (O_1972,N_29854,N_29406);
nor UO_1973 (O_1973,N_29669,N_29309);
and UO_1974 (O_1974,N_29271,N_29610);
or UO_1975 (O_1975,N_29509,N_29362);
nand UO_1976 (O_1976,N_29911,N_29677);
nor UO_1977 (O_1977,N_29969,N_28880);
or UO_1978 (O_1978,N_29684,N_29453);
or UO_1979 (O_1979,N_29680,N_29205);
and UO_1980 (O_1980,N_29007,N_29368);
and UO_1981 (O_1981,N_29396,N_29198);
or UO_1982 (O_1982,N_29236,N_29138);
or UO_1983 (O_1983,N_29083,N_29412);
nor UO_1984 (O_1984,N_28876,N_29698);
nor UO_1985 (O_1985,N_29331,N_29365);
and UO_1986 (O_1986,N_29349,N_29988);
and UO_1987 (O_1987,N_29675,N_29364);
and UO_1988 (O_1988,N_29560,N_29366);
nor UO_1989 (O_1989,N_29808,N_29432);
nand UO_1990 (O_1990,N_29359,N_29428);
nand UO_1991 (O_1991,N_29727,N_29316);
and UO_1992 (O_1992,N_29157,N_29249);
and UO_1993 (O_1993,N_28935,N_29034);
xnor UO_1994 (O_1994,N_29687,N_29177);
nand UO_1995 (O_1995,N_29935,N_29893);
and UO_1996 (O_1996,N_29469,N_29394);
and UO_1997 (O_1997,N_29347,N_29866);
or UO_1998 (O_1998,N_29284,N_29161);
nand UO_1999 (O_1999,N_29927,N_28867);
or UO_2000 (O_2000,N_29359,N_29287);
nor UO_2001 (O_2001,N_29325,N_28866);
and UO_2002 (O_2002,N_29935,N_28942);
nor UO_2003 (O_2003,N_29072,N_28868);
nor UO_2004 (O_2004,N_29295,N_29450);
and UO_2005 (O_2005,N_29059,N_29872);
and UO_2006 (O_2006,N_28978,N_29708);
nor UO_2007 (O_2007,N_28819,N_29823);
nand UO_2008 (O_2008,N_29490,N_29935);
xnor UO_2009 (O_2009,N_29368,N_29780);
and UO_2010 (O_2010,N_29955,N_28919);
nand UO_2011 (O_2011,N_29332,N_29234);
nor UO_2012 (O_2012,N_28815,N_29084);
and UO_2013 (O_2013,N_29743,N_29616);
and UO_2014 (O_2014,N_29473,N_28879);
xnor UO_2015 (O_2015,N_28946,N_29369);
nor UO_2016 (O_2016,N_29917,N_29383);
xor UO_2017 (O_2017,N_29792,N_28835);
nor UO_2018 (O_2018,N_29516,N_29633);
nor UO_2019 (O_2019,N_29048,N_28855);
nor UO_2020 (O_2020,N_29836,N_29049);
nor UO_2021 (O_2021,N_29955,N_28907);
nor UO_2022 (O_2022,N_29470,N_29987);
nor UO_2023 (O_2023,N_29191,N_29187);
nor UO_2024 (O_2024,N_29024,N_29086);
nand UO_2025 (O_2025,N_28813,N_28862);
nor UO_2026 (O_2026,N_28900,N_29780);
and UO_2027 (O_2027,N_29804,N_29142);
nand UO_2028 (O_2028,N_29470,N_28882);
and UO_2029 (O_2029,N_29172,N_29151);
or UO_2030 (O_2030,N_29190,N_29794);
xnor UO_2031 (O_2031,N_29090,N_29882);
and UO_2032 (O_2032,N_29616,N_29378);
nand UO_2033 (O_2033,N_29294,N_29605);
xnor UO_2034 (O_2034,N_29285,N_28851);
nor UO_2035 (O_2035,N_29885,N_29486);
xor UO_2036 (O_2036,N_28929,N_29108);
xor UO_2037 (O_2037,N_29139,N_29648);
xnor UO_2038 (O_2038,N_29342,N_29298);
nor UO_2039 (O_2039,N_29116,N_29182);
nand UO_2040 (O_2040,N_28897,N_29433);
nor UO_2041 (O_2041,N_29109,N_29776);
or UO_2042 (O_2042,N_29917,N_29394);
and UO_2043 (O_2043,N_28809,N_29156);
and UO_2044 (O_2044,N_29384,N_29749);
nand UO_2045 (O_2045,N_29816,N_29688);
or UO_2046 (O_2046,N_28850,N_29689);
and UO_2047 (O_2047,N_29028,N_28970);
and UO_2048 (O_2048,N_29393,N_29957);
xnor UO_2049 (O_2049,N_29603,N_29684);
or UO_2050 (O_2050,N_29947,N_29397);
or UO_2051 (O_2051,N_29156,N_29018);
or UO_2052 (O_2052,N_29420,N_29934);
xor UO_2053 (O_2053,N_29160,N_29271);
nor UO_2054 (O_2054,N_29938,N_29795);
nand UO_2055 (O_2055,N_29074,N_29984);
xor UO_2056 (O_2056,N_28982,N_29213);
nor UO_2057 (O_2057,N_29825,N_29844);
and UO_2058 (O_2058,N_29219,N_28818);
xor UO_2059 (O_2059,N_29790,N_29463);
xnor UO_2060 (O_2060,N_29514,N_29159);
nand UO_2061 (O_2061,N_29789,N_28804);
or UO_2062 (O_2062,N_29797,N_29364);
nor UO_2063 (O_2063,N_29165,N_28822);
nor UO_2064 (O_2064,N_29018,N_29012);
xnor UO_2065 (O_2065,N_29456,N_29582);
or UO_2066 (O_2066,N_29153,N_29879);
nand UO_2067 (O_2067,N_28867,N_29031);
or UO_2068 (O_2068,N_29506,N_29773);
xor UO_2069 (O_2069,N_29686,N_29827);
and UO_2070 (O_2070,N_29347,N_29238);
and UO_2071 (O_2071,N_29534,N_29311);
and UO_2072 (O_2072,N_29691,N_29491);
nor UO_2073 (O_2073,N_28815,N_29755);
xor UO_2074 (O_2074,N_29473,N_29858);
and UO_2075 (O_2075,N_29147,N_29162);
and UO_2076 (O_2076,N_29793,N_28877);
and UO_2077 (O_2077,N_28971,N_29785);
and UO_2078 (O_2078,N_29526,N_28871);
nor UO_2079 (O_2079,N_29721,N_29916);
nor UO_2080 (O_2080,N_29379,N_29096);
nand UO_2081 (O_2081,N_29546,N_28909);
xnor UO_2082 (O_2082,N_29678,N_29100);
nor UO_2083 (O_2083,N_28965,N_29757);
nand UO_2084 (O_2084,N_29185,N_28980);
or UO_2085 (O_2085,N_29496,N_29673);
nand UO_2086 (O_2086,N_29104,N_29433);
xor UO_2087 (O_2087,N_29726,N_29526);
xnor UO_2088 (O_2088,N_29571,N_29405);
nand UO_2089 (O_2089,N_29675,N_29234);
or UO_2090 (O_2090,N_29622,N_29328);
nand UO_2091 (O_2091,N_29904,N_28908);
and UO_2092 (O_2092,N_29658,N_28979);
nand UO_2093 (O_2093,N_29977,N_29595);
nand UO_2094 (O_2094,N_28983,N_29126);
nand UO_2095 (O_2095,N_28844,N_29600);
and UO_2096 (O_2096,N_29271,N_29773);
nor UO_2097 (O_2097,N_28982,N_28989);
xnor UO_2098 (O_2098,N_29915,N_29939);
nor UO_2099 (O_2099,N_29057,N_29661);
nand UO_2100 (O_2100,N_29144,N_29664);
nand UO_2101 (O_2101,N_29505,N_29491);
and UO_2102 (O_2102,N_29701,N_29116);
and UO_2103 (O_2103,N_29500,N_28940);
or UO_2104 (O_2104,N_29804,N_29636);
or UO_2105 (O_2105,N_29130,N_29085);
and UO_2106 (O_2106,N_29455,N_29548);
and UO_2107 (O_2107,N_28899,N_29285);
nand UO_2108 (O_2108,N_29636,N_28869);
nand UO_2109 (O_2109,N_28924,N_29194);
nand UO_2110 (O_2110,N_29058,N_29685);
or UO_2111 (O_2111,N_28859,N_28963);
nor UO_2112 (O_2112,N_28842,N_29767);
nand UO_2113 (O_2113,N_29749,N_29363);
nand UO_2114 (O_2114,N_29235,N_29436);
and UO_2115 (O_2115,N_29446,N_29738);
or UO_2116 (O_2116,N_29290,N_29021);
nand UO_2117 (O_2117,N_29080,N_29711);
nor UO_2118 (O_2118,N_28923,N_29138);
and UO_2119 (O_2119,N_29144,N_29709);
nand UO_2120 (O_2120,N_28881,N_28880);
nand UO_2121 (O_2121,N_29695,N_29664);
and UO_2122 (O_2122,N_28918,N_28855);
or UO_2123 (O_2123,N_29214,N_29095);
and UO_2124 (O_2124,N_29337,N_29597);
nor UO_2125 (O_2125,N_29475,N_29753);
nor UO_2126 (O_2126,N_28906,N_29237);
or UO_2127 (O_2127,N_29726,N_29689);
nor UO_2128 (O_2128,N_29326,N_29910);
or UO_2129 (O_2129,N_29191,N_29161);
nand UO_2130 (O_2130,N_29198,N_29559);
xor UO_2131 (O_2131,N_29488,N_29746);
or UO_2132 (O_2132,N_29542,N_28934);
or UO_2133 (O_2133,N_29077,N_29684);
nor UO_2134 (O_2134,N_29651,N_29740);
or UO_2135 (O_2135,N_29686,N_29365);
nand UO_2136 (O_2136,N_29872,N_29189);
and UO_2137 (O_2137,N_29465,N_29331);
or UO_2138 (O_2138,N_28940,N_29601);
and UO_2139 (O_2139,N_28854,N_29484);
nand UO_2140 (O_2140,N_28888,N_28886);
and UO_2141 (O_2141,N_29650,N_29281);
xnor UO_2142 (O_2142,N_29927,N_29226);
nor UO_2143 (O_2143,N_28870,N_28994);
and UO_2144 (O_2144,N_29135,N_29644);
or UO_2145 (O_2145,N_29449,N_28967);
nor UO_2146 (O_2146,N_29315,N_29575);
nand UO_2147 (O_2147,N_29504,N_29581);
or UO_2148 (O_2148,N_29081,N_29234);
xor UO_2149 (O_2149,N_29459,N_29989);
nand UO_2150 (O_2150,N_29600,N_29382);
or UO_2151 (O_2151,N_29930,N_28864);
nor UO_2152 (O_2152,N_29701,N_29074);
nand UO_2153 (O_2153,N_29468,N_29151);
or UO_2154 (O_2154,N_29865,N_28876);
and UO_2155 (O_2155,N_29112,N_29509);
or UO_2156 (O_2156,N_29493,N_28840);
nand UO_2157 (O_2157,N_29482,N_29599);
xnor UO_2158 (O_2158,N_29274,N_29894);
or UO_2159 (O_2159,N_29435,N_29718);
or UO_2160 (O_2160,N_28932,N_29880);
nor UO_2161 (O_2161,N_29700,N_29441);
xnor UO_2162 (O_2162,N_28995,N_29261);
nand UO_2163 (O_2163,N_29888,N_28871);
and UO_2164 (O_2164,N_29604,N_29285);
xor UO_2165 (O_2165,N_29962,N_29829);
xor UO_2166 (O_2166,N_28944,N_28835);
nor UO_2167 (O_2167,N_29889,N_29301);
xnor UO_2168 (O_2168,N_29495,N_28980);
nor UO_2169 (O_2169,N_29889,N_29931);
or UO_2170 (O_2170,N_28814,N_29476);
nand UO_2171 (O_2171,N_29179,N_28985);
nand UO_2172 (O_2172,N_28888,N_29106);
nor UO_2173 (O_2173,N_29086,N_29255);
nand UO_2174 (O_2174,N_29168,N_29808);
or UO_2175 (O_2175,N_29695,N_29469);
or UO_2176 (O_2176,N_29517,N_28804);
or UO_2177 (O_2177,N_29750,N_29754);
xor UO_2178 (O_2178,N_29315,N_29420);
nor UO_2179 (O_2179,N_29536,N_29249);
and UO_2180 (O_2180,N_29141,N_29171);
xor UO_2181 (O_2181,N_29884,N_29494);
nand UO_2182 (O_2182,N_29879,N_28830);
nand UO_2183 (O_2183,N_29865,N_29688);
nor UO_2184 (O_2184,N_29963,N_29927);
xnor UO_2185 (O_2185,N_29290,N_29273);
nand UO_2186 (O_2186,N_29713,N_29096);
or UO_2187 (O_2187,N_29175,N_29591);
nor UO_2188 (O_2188,N_29497,N_29784);
xnor UO_2189 (O_2189,N_29167,N_29890);
nand UO_2190 (O_2190,N_29452,N_29075);
nand UO_2191 (O_2191,N_29144,N_29752);
nand UO_2192 (O_2192,N_29596,N_29047);
and UO_2193 (O_2193,N_29108,N_29460);
nand UO_2194 (O_2194,N_29271,N_29466);
and UO_2195 (O_2195,N_29644,N_29759);
nor UO_2196 (O_2196,N_29259,N_29218);
nand UO_2197 (O_2197,N_29351,N_29993);
nand UO_2198 (O_2198,N_29288,N_29692);
or UO_2199 (O_2199,N_29215,N_29332);
or UO_2200 (O_2200,N_29578,N_29693);
nand UO_2201 (O_2201,N_29321,N_29867);
xor UO_2202 (O_2202,N_29168,N_28819);
nor UO_2203 (O_2203,N_29804,N_29599);
or UO_2204 (O_2204,N_29044,N_29620);
nand UO_2205 (O_2205,N_29647,N_29705);
nand UO_2206 (O_2206,N_29320,N_29488);
and UO_2207 (O_2207,N_29932,N_29800);
xor UO_2208 (O_2208,N_29781,N_29185);
xor UO_2209 (O_2209,N_29463,N_29120);
or UO_2210 (O_2210,N_29258,N_29236);
nor UO_2211 (O_2211,N_29205,N_29559);
xor UO_2212 (O_2212,N_29370,N_29347);
nand UO_2213 (O_2213,N_29851,N_28864);
and UO_2214 (O_2214,N_29680,N_29487);
xnor UO_2215 (O_2215,N_29346,N_29048);
or UO_2216 (O_2216,N_29271,N_29220);
and UO_2217 (O_2217,N_29808,N_29787);
nand UO_2218 (O_2218,N_28924,N_28920);
xnor UO_2219 (O_2219,N_29953,N_29128);
and UO_2220 (O_2220,N_29618,N_29292);
nor UO_2221 (O_2221,N_29455,N_28829);
or UO_2222 (O_2222,N_29476,N_29972);
nand UO_2223 (O_2223,N_29437,N_29870);
xor UO_2224 (O_2224,N_29868,N_28932);
nor UO_2225 (O_2225,N_29165,N_29637);
and UO_2226 (O_2226,N_29895,N_29741);
nand UO_2227 (O_2227,N_29808,N_29541);
nor UO_2228 (O_2228,N_29903,N_29347);
nor UO_2229 (O_2229,N_29790,N_29392);
nor UO_2230 (O_2230,N_28806,N_29055);
and UO_2231 (O_2231,N_29279,N_29532);
nor UO_2232 (O_2232,N_28945,N_29899);
xnor UO_2233 (O_2233,N_29654,N_29336);
nand UO_2234 (O_2234,N_29410,N_29493);
or UO_2235 (O_2235,N_29473,N_29351);
and UO_2236 (O_2236,N_29295,N_29921);
or UO_2237 (O_2237,N_29686,N_29188);
nand UO_2238 (O_2238,N_28819,N_29325);
xnor UO_2239 (O_2239,N_29762,N_28864);
nor UO_2240 (O_2240,N_29336,N_29509);
nor UO_2241 (O_2241,N_29254,N_29240);
and UO_2242 (O_2242,N_29799,N_29021);
nand UO_2243 (O_2243,N_29715,N_29666);
xnor UO_2244 (O_2244,N_28981,N_29334);
nand UO_2245 (O_2245,N_29830,N_29859);
or UO_2246 (O_2246,N_29319,N_28998);
nor UO_2247 (O_2247,N_29212,N_29627);
and UO_2248 (O_2248,N_29104,N_29676);
xor UO_2249 (O_2249,N_29769,N_29627);
and UO_2250 (O_2250,N_29861,N_29889);
xnor UO_2251 (O_2251,N_29369,N_29481);
and UO_2252 (O_2252,N_29206,N_29441);
or UO_2253 (O_2253,N_29249,N_29853);
nand UO_2254 (O_2254,N_29290,N_29677);
nand UO_2255 (O_2255,N_29455,N_29725);
or UO_2256 (O_2256,N_29653,N_29126);
xnor UO_2257 (O_2257,N_28987,N_29565);
and UO_2258 (O_2258,N_29777,N_29882);
nor UO_2259 (O_2259,N_29284,N_29984);
xnor UO_2260 (O_2260,N_28932,N_29217);
nor UO_2261 (O_2261,N_29285,N_29218);
nand UO_2262 (O_2262,N_28964,N_29731);
nor UO_2263 (O_2263,N_29248,N_28924);
nor UO_2264 (O_2264,N_28894,N_28813);
nor UO_2265 (O_2265,N_28827,N_29373);
xor UO_2266 (O_2266,N_29180,N_29125);
nand UO_2267 (O_2267,N_29690,N_29644);
or UO_2268 (O_2268,N_29225,N_28869);
xor UO_2269 (O_2269,N_28899,N_29161);
xor UO_2270 (O_2270,N_29137,N_29750);
or UO_2271 (O_2271,N_29374,N_29013);
xnor UO_2272 (O_2272,N_29535,N_29432);
xor UO_2273 (O_2273,N_29875,N_29723);
nand UO_2274 (O_2274,N_29037,N_29343);
nor UO_2275 (O_2275,N_29284,N_29589);
nand UO_2276 (O_2276,N_29810,N_28937);
xor UO_2277 (O_2277,N_28827,N_29257);
xor UO_2278 (O_2278,N_29072,N_28890);
xnor UO_2279 (O_2279,N_29633,N_29249);
nor UO_2280 (O_2280,N_29193,N_29133);
xnor UO_2281 (O_2281,N_28867,N_29161);
xnor UO_2282 (O_2282,N_28969,N_29608);
nand UO_2283 (O_2283,N_29505,N_29801);
or UO_2284 (O_2284,N_29319,N_29157);
and UO_2285 (O_2285,N_28919,N_28946);
nand UO_2286 (O_2286,N_29295,N_29770);
nor UO_2287 (O_2287,N_29361,N_29915);
or UO_2288 (O_2288,N_29725,N_29733);
and UO_2289 (O_2289,N_28801,N_29710);
xnor UO_2290 (O_2290,N_29099,N_29794);
or UO_2291 (O_2291,N_28944,N_29948);
xnor UO_2292 (O_2292,N_29631,N_29335);
or UO_2293 (O_2293,N_28919,N_29795);
and UO_2294 (O_2294,N_29740,N_29085);
nand UO_2295 (O_2295,N_29532,N_29588);
nand UO_2296 (O_2296,N_28866,N_28903);
xor UO_2297 (O_2297,N_28830,N_28945);
xor UO_2298 (O_2298,N_28972,N_29418);
xnor UO_2299 (O_2299,N_29655,N_29943);
nor UO_2300 (O_2300,N_28983,N_29563);
nand UO_2301 (O_2301,N_29822,N_29745);
and UO_2302 (O_2302,N_29948,N_28923);
nand UO_2303 (O_2303,N_29642,N_29425);
nand UO_2304 (O_2304,N_28939,N_29452);
or UO_2305 (O_2305,N_28821,N_28823);
xnor UO_2306 (O_2306,N_29074,N_28958);
and UO_2307 (O_2307,N_29256,N_29348);
xnor UO_2308 (O_2308,N_29094,N_29517);
and UO_2309 (O_2309,N_29482,N_29478);
nor UO_2310 (O_2310,N_29938,N_28841);
nor UO_2311 (O_2311,N_29645,N_29011);
nor UO_2312 (O_2312,N_29598,N_29560);
and UO_2313 (O_2313,N_29712,N_29958);
and UO_2314 (O_2314,N_29800,N_29597);
xnor UO_2315 (O_2315,N_29781,N_29079);
xnor UO_2316 (O_2316,N_29333,N_29240);
xnor UO_2317 (O_2317,N_29864,N_29862);
nand UO_2318 (O_2318,N_29591,N_29359);
xnor UO_2319 (O_2319,N_29620,N_29903);
and UO_2320 (O_2320,N_29588,N_29150);
or UO_2321 (O_2321,N_29437,N_29183);
nor UO_2322 (O_2322,N_28986,N_29815);
and UO_2323 (O_2323,N_29413,N_29845);
nor UO_2324 (O_2324,N_29035,N_29236);
nor UO_2325 (O_2325,N_29635,N_29654);
xor UO_2326 (O_2326,N_28866,N_29279);
xor UO_2327 (O_2327,N_29752,N_29938);
nand UO_2328 (O_2328,N_29130,N_29485);
nand UO_2329 (O_2329,N_29384,N_29860);
nor UO_2330 (O_2330,N_29575,N_29463);
xnor UO_2331 (O_2331,N_29284,N_29998);
xnor UO_2332 (O_2332,N_29048,N_29363);
nor UO_2333 (O_2333,N_29799,N_29623);
or UO_2334 (O_2334,N_29893,N_29153);
nor UO_2335 (O_2335,N_29419,N_29268);
or UO_2336 (O_2336,N_29475,N_29807);
nand UO_2337 (O_2337,N_29244,N_29853);
or UO_2338 (O_2338,N_29184,N_29142);
xnor UO_2339 (O_2339,N_29572,N_28920);
or UO_2340 (O_2340,N_29031,N_29608);
nand UO_2341 (O_2341,N_29916,N_28840);
or UO_2342 (O_2342,N_29191,N_28826);
nand UO_2343 (O_2343,N_29656,N_29133);
nand UO_2344 (O_2344,N_29741,N_28962);
or UO_2345 (O_2345,N_29187,N_29644);
nor UO_2346 (O_2346,N_28972,N_28867);
and UO_2347 (O_2347,N_28821,N_29769);
nor UO_2348 (O_2348,N_29028,N_29852);
nand UO_2349 (O_2349,N_29458,N_29526);
and UO_2350 (O_2350,N_28908,N_29050);
xnor UO_2351 (O_2351,N_29597,N_29130);
nand UO_2352 (O_2352,N_29663,N_29657);
xnor UO_2353 (O_2353,N_29389,N_29788);
nor UO_2354 (O_2354,N_29650,N_29955);
or UO_2355 (O_2355,N_29855,N_29316);
xnor UO_2356 (O_2356,N_28827,N_29262);
or UO_2357 (O_2357,N_29819,N_29403);
nand UO_2358 (O_2358,N_29309,N_29788);
nand UO_2359 (O_2359,N_29164,N_29834);
or UO_2360 (O_2360,N_28905,N_29586);
xor UO_2361 (O_2361,N_29264,N_29657);
nand UO_2362 (O_2362,N_29701,N_28932);
and UO_2363 (O_2363,N_29316,N_29108);
and UO_2364 (O_2364,N_28822,N_29259);
or UO_2365 (O_2365,N_29684,N_28937);
nand UO_2366 (O_2366,N_29505,N_29758);
nand UO_2367 (O_2367,N_29573,N_29940);
xnor UO_2368 (O_2368,N_28849,N_29076);
and UO_2369 (O_2369,N_29876,N_29435);
xor UO_2370 (O_2370,N_29372,N_28881);
and UO_2371 (O_2371,N_28981,N_28872);
or UO_2372 (O_2372,N_29243,N_29209);
nand UO_2373 (O_2373,N_29975,N_29034);
xor UO_2374 (O_2374,N_29742,N_29635);
nor UO_2375 (O_2375,N_28827,N_29510);
and UO_2376 (O_2376,N_29042,N_28889);
nor UO_2377 (O_2377,N_29398,N_29817);
or UO_2378 (O_2378,N_29493,N_29777);
or UO_2379 (O_2379,N_29401,N_29967);
and UO_2380 (O_2380,N_29637,N_29301);
xnor UO_2381 (O_2381,N_29838,N_29834);
nand UO_2382 (O_2382,N_28903,N_29575);
nor UO_2383 (O_2383,N_29883,N_29763);
nand UO_2384 (O_2384,N_29840,N_28936);
or UO_2385 (O_2385,N_29713,N_29233);
nand UO_2386 (O_2386,N_29279,N_28934);
or UO_2387 (O_2387,N_29529,N_29378);
nor UO_2388 (O_2388,N_29314,N_28852);
or UO_2389 (O_2389,N_29366,N_29630);
nor UO_2390 (O_2390,N_29673,N_29789);
and UO_2391 (O_2391,N_29471,N_29974);
or UO_2392 (O_2392,N_29261,N_29167);
nand UO_2393 (O_2393,N_29379,N_29246);
and UO_2394 (O_2394,N_28890,N_29813);
and UO_2395 (O_2395,N_29937,N_29387);
nor UO_2396 (O_2396,N_29730,N_28861);
and UO_2397 (O_2397,N_28886,N_29644);
nor UO_2398 (O_2398,N_29183,N_29069);
nor UO_2399 (O_2399,N_29406,N_29358);
or UO_2400 (O_2400,N_28958,N_29694);
nor UO_2401 (O_2401,N_29784,N_29235);
xor UO_2402 (O_2402,N_29415,N_29050);
or UO_2403 (O_2403,N_28869,N_29858);
nor UO_2404 (O_2404,N_29907,N_28959);
nor UO_2405 (O_2405,N_29051,N_29225);
and UO_2406 (O_2406,N_29496,N_29294);
nor UO_2407 (O_2407,N_29597,N_29929);
nand UO_2408 (O_2408,N_29936,N_29482);
xnor UO_2409 (O_2409,N_28956,N_29777);
nand UO_2410 (O_2410,N_28887,N_28852);
nor UO_2411 (O_2411,N_29567,N_29832);
nand UO_2412 (O_2412,N_29523,N_29283);
or UO_2413 (O_2413,N_29328,N_28935);
or UO_2414 (O_2414,N_29290,N_29702);
or UO_2415 (O_2415,N_29936,N_29939);
nand UO_2416 (O_2416,N_29345,N_29599);
nor UO_2417 (O_2417,N_29136,N_28876);
xnor UO_2418 (O_2418,N_29789,N_29264);
nor UO_2419 (O_2419,N_28972,N_29735);
nand UO_2420 (O_2420,N_29022,N_29784);
and UO_2421 (O_2421,N_29522,N_29966);
xnor UO_2422 (O_2422,N_28881,N_29726);
xor UO_2423 (O_2423,N_29663,N_29003);
nor UO_2424 (O_2424,N_29681,N_28954);
and UO_2425 (O_2425,N_29592,N_29542);
xnor UO_2426 (O_2426,N_29193,N_29219);
xnor UO_2427 (O_2427,N_28820,N_29344);
or UO_2428 (O_2428,N_29470,N_29919);
or UO_2429 (O_2429,N_29692,N_28850);
xor UO_2430 (O_2430,N_29101,N_29757);
or UO_2431 (O_2431,N_29077,N_29716);
xor UO_2432 (O_2432,N_29601,N_29691);
nand UO_2433 (O_2433,N_29399,N_29893);
nor UO_2434 (O_2434,N_29399,N_28833);
nand UO_2435 (O_2435,N_29276,N_29429);
and UO_2436 (O_2436,N_29846,N_29654);
nor UO_2437 (O_2437,N_29810,N_29105);
nand UO_2438 (O_2438,N_28802,N_28908);
or UO_2439 (O_2439,N_29187,N_29046);
or UO_2440 (O_2440,N_29726,N_29147);
nor UO_2441 (O_2441,N_29897,N_29373);
nor UO_2442 (O_2442,N_29204,N_29684);
and UO_2443 (O_2443,N_28856,N_29126);
nand UO_2444 (O_2444,N_29071,N_29133);
and UO_2445 (O_2445,N_29431,N_29378);
xor UO_2446 (O_2446,N_29325,N_29134);
nor UO_2447 (O_2447,N_28994,N_29645);
nand UO_2448 (O_2448,N_29884,N_29441);
or UO_2449 (O_2449,N_29753,N_29169);
and UO_2450 (O_2450,N_29055,N_28822);
nand UO_2451 (O_2451,N_29449,N_29146);
xnor UO_2452 (O_2452,N_29262,N_29327);
nand UO_2453 (O_2453,N_29909,N_29002);
and UO_2454 (O_2454,N_29663,N_29317);
nand UO_2455 (O_2455,N_29038,N_29883);
or UO_2456 (O_2456,N_29299,N_29677);
and UO_2457 (O_2457,N_29221,N_29673);
nor UO_2458 (O_2458,N_29344,N_29172);
nor UO_2459 (O_2459,N_28905,N_29993);
nor UO_2460 (O_2460,N_29841,N_29833);
xor UO_2461 (O_2461,N_29749,N_29103);
nor UO_2462 (O_2462,N_28993,N_29033);
nor UO_2463 (O_2463,N_29257,N_29340);
and UO_2464 (O_2464,N_29629,N_29878);
and UO_2465 (O_2465,N_28968,N_29775);
nand UO_2466 (O_2466,N_28933,N_29714);
nand UO_2467 (O_2467,N_28888,N_29074);
xor UO_2468 (O_2468,N_29830,N_28872);
or UO_2469 (O_2469,N_29497,N_29005);
and UO_2470 (O_2470,N_29948,N_29837);
or UO_2471 (O_2471,N_29563,N_29621);
xnor UO_2472 (O_2472,N_29852,N_29502);
nor UO_2473 (O_2473,N_29097,N_29854);
nor UO_2474 (O_2474,N_29119,N_29130);
xnor UO_2475 (O_2475,N_29600,N_28838);
or UO_2476 (O_2476,N_28840,N_29355);
nor UO_2477 (O_2477,N_29504,N_29489);
xnor UO_2478 (O_2478,N_28879,N_29077);
or UO_2479 (O_2479,N_28853,N_29964);
nand UO_2480 (O_2480,N_29598,N_29046);
or UO_2481 (O_2481,N_28817,N_29484);
nor UO_2482 (O_2482,N_29816,N_29619);
and UO_2483 (O_2483,N_29389,N_29764);
xor UO_2484 (O_2484,N_29233,N_29611);
nor UO_2485 (O_2485,N_29997,N_29985);
and UO_2486 (O_2486,N_28928,N_28938);
nor UO_2487 (O_2487,N_28872,N_29717);
nand UO_2488 (O_2488,N_29695,N_29822);
nor UO_2489 (O_2489,N_29539,N_29481);
and UO_2490 (O_2490,N_29409,N_29139);
nor UO_2491 (O_2491,N_29483,N_29500);
xnor UO_2492 (O_2492,N_29760,N_29233);
or UO_2493 (O_2493,N_28806,N_29233);
xor UO_2494 (O_2494,N_29142,N_29843);
and UO_2495 (O_2495,N_29488,N_29003);
nand UO_2496 (O_2496,N_28883,N_29324);
and UO_2497 (O_2497,N_29901,N_29557);
xnor UO_2498 (O_2498,N_28902,N_29109);
and UO_2499 (O_2499,N_28992,N_29246);
xnor UO_2500 (O_2500,N_29575,N_29753);
nor UO_2501 (O_2501,N_29015,N_29753);
nand UO_2502 (O_2502,N_28865,N_29583);
nor UO_2503 (O_2503,N_29656,N_29658);
nand UO_2504 (O_2504,N_29291,N_29644);
nand UO_2505 (O_2505,N_29595,N_29379);
and UO_2506 (O_2506,N_28965,N_29559);
or UO_2507 (O_2507,N_28898,N_29233);
and UO_2508 (O_2508,N_28859,N_29889);
nor UO_2509 (O_2509,N_29910,N_29980);
and UO_2510 (O_2510,N_29723,N_29250);
xnor UO_2511 (O_2511,N_29392,N_29535);
xor UO_2512 (O_2512,N_29530,N_28942);
nand UO_2513 (O_2513,N_29778,N_29520);
and UO_2514 (O_2514,N_29850,N_29199);
nand UO_2515 (O_2515,N_29525,N_29745);
nor UO_2516 (O_2516,N_29284,N_29069);
and UO_2517 (O_2517,N_29776,N_29967);
nor UO_2518 (O_2518,N_29546,N_29723);
xnor UO_2519 (O_2519,N_29734,N_29968);
nor UO_2520 (O_2520,N_29775,N_29459);
and UO_2521 (O_2521,N_29587,N_29292);
xnor UO_2522 (O_2522,N_28895,N_29150);
nor UO_2523 (O_2523,N_29630,N_28984);
nand UO_2524 (O_2524,N_28935,N_29007);
or UO_2525 (O_2525,N_29711,N_29776);
or UO_2526 (O_2526,N_28875,N_29273);
nand UO_2527 (O_2527,N_29993,N_29120);
xor UO_2528 (O_2528,N_29663,N_29435);
and UO_2529 (O_2529,N_29925,N_29093);
or UO_2530 (O_2530,N_29814,N_29400);
nor UO_2531 (O_2531,N_29767,N_29240);
or UO_2532 (O_2532,N_28840,N_29936);
and UO_2533 (O_2533,N_29731,N_29433);
nand UO_2534 (O_2534,N_29083,N_29239);
xor UO_2535 (O_2535,N_29022,N_29788);
and UO_2536 (O_2536,N_29842,N_29666);
or UO_2537 (O_2537,N_29699,N_29078);
nor UO_2538 (O_2538,N_29396,N_29681);
or UO_2539 (O_2539,N_29968,N_29608);
nand UO_2540 (O_2540,N_29207,N_29817);
or UO_2541 (O_2541,N_29714,N_29334);
nand UO_2542 (O_2542,N_29931,N_29554);
nand UO_2543 (O_2543,N_29639,N_29832);
or UO_2544 (O_2544,N_29154,N_29601);
and UO_2545 (O_2545,N_29509,N_29765);
nand UO_2546 (O_2546,N_29132,N_29589);
or UO_2547 (O_2547,N_29204,N_29340);
or UO_2548 (O_2548,N_29441,N_29289);
nor UO_2549 (O_2549,N_29257,N_29476);
nand UO_2550 (O_2550,N_29807,N_28815);
xor UO_2551 (O_2551,N_29053,N_29816);
and UO_2552 (O_2552,N_29433,N_28987);
xor UO_2553 (O_2553,N_29524,N_29816);
or UO_2554 (O_2554,N_29274,N_29714);
nor UO_2555 (O_2555,N_29328,N_29027);
and UO_2556 (O_2556,N_28825,N_29692);
or UO_2557 (O_2557,N_28955,N_29706);
or UO_2558 (O_2558,N_29132,N_29034);
nor UO_2559 (O_2559,N_29670,N_28904);
and UO_2560 (O_2560,N_29687,N_29778);
nor UO_2561 (O_2561,N_29151,N_29945);
xor UO_2562 (O_2562,N_29670,N_29255);
xor UO_2563 (O_2563,N_28979,N_28862);
and UO_2564 (O_2564,N_29669,N_29332);
nand UO_2565 (O_2565,N_29081,N_29935);
and UO_2566 (O_2566,N_29048,N_29009);
or UO_2567 (O_2567,N_29000,N_29721);
nor UO_2568 (O_2568,N_29718,N_29679);
or UO_2569 (O_2569,N_29022,N_29070);
and UO_2570 (O_2570,N_29094,N_29959);
and UO_2571 (O_2571,N_29747,N_29974);
nand UO_2572 (O_2572,N_29496,N_29105);
nor UO_2573 (O_2573,N_29759,N_29097);
nand UO_2574 (O_2574,N_29155,N_29073);
nand UO_2575 (O_2575,N_29242,N_29288);
nor UO_2576 (O_2576,N_29508,N_29875);
nand UO_2577 (O_2577,N_29964,N_29833);
and UO_2578 (O_2578,N_29830,N_29155);
and UO_2579 (O_2579,N_29407,N_29202);
nand UO_2580 (O_2580,N_29795,N_29674);
and UO_2581 (O_2581,N_29738,N_29261);
or UO_2582 (O_2582,N_29402,N_29028);
nor UO_2583 (O_2583,N_29968,N_29589);
and UO_2584 (O_2584,N_29827,N_29780);
or UO_2585 (O_2585,N_28962,N_28945);
or UO_2586 (O_2586,N_29954,N_29500);
or UO_2587 (O_2587,N_29512,N_28967);
or UO_2588 (O_2588,N_29951,N_29545);
xnor UO_2589 (O_2589,N_29024,N_29335);
xor UO_2590 (O_2590,N_29661,N_29301);
nand UO_2591 (O_2591,N_29289,N_29001);
or UO_2592 (O_2592,N_29661,N_29458);
and UO_2593 (O_2593,N_29510,N_28960);
and UO_2594 (O_2594,N_29740,N_29543);
and UO_2595 (O_2595,N_29102,N_28886);
and UO_2596 (O_2596,N_29345,N_29372);
or UO_2597 (O_2597,N_29947,N_29085);
and UO_2598 (O_2598,N_29775,N_29521);
and UO_2599 (O_2599,N_28924,N_29353);
nor UO_2600 (O_2600,N_28838,N_29877);
nor UO_2601 (O_2601,N_29401,N_29878);
nor UO_2602 (O_2602,N_29161,N_29913);
nor UO_2603 (O_2603,N_28808,N_29296);
or UO_2604 (O_2604,N_29852,N_29547);
nor UO_2605 (O_2605,N_28825,N_29734);
and UO_2606 (O_2606,N_29741,N_29265);
nand UO_2607 (O_2607,N_28950,N_29954);
or UO_2608 (O_2608,N_29590,N_29449);
nor UO_2609 (O_2609,N_29394,N_28998);
nand UO_2610 (O_2610,N_29717,N_29062);
or UO_2611 (O_2611,N_29457,N_29262);
nor UO_2612 (O_2612,N_28883,N_29500);
and UO_2613 (O_2613,N_29997,N_29299);
or UO_2614 (O_2614,N_29843,N_29375);
and UO_2615 (O_2615,N_29968,N_29281);
xor UO_2616 (O_2616,N_29751,N_29295);
and UO_2617 (O_2617,N_29609,N_29362);
nand UO_2618 (O_2618,N_29528,N_28963);
xor UO_2619 (O_2619,N_28942,N_29817);
or UO_2620 (O_2620,N_29500,N_29448);
or UO_2621 (O_2621,N_29311,N_29908);
nand UO_2622 (O_2622,N_29678,N_29313);
nor UO_2623 (O_2623,N_29091,N_29715);
and UO_2624 (O_2624,N_29361,N_29145);
nand UO_2625 (O_2625,N_29254,N_29148);
nand UO_2626 (O_2626,N_29454,N_28880);
nor UO_2627 (O_2627,N_28970,N_29163);
nor UO_2628 (O_2628,N_29958,N_29533);
nand UO_2629 (O_2629,N_29134,N_29686);
nor UO_2630 (O_2630,N_29488,N_29862);
xnor UO_2631 (O_2631,N_29569,N_29056);
or UO_2632 (O_2632,N_28997,N_29399);
nand UO_2633 (O_2633,N_29662,N_28919);
and UO_2634 (O_2634,N_29208,N_28857);
nor UO_2635 (O_2635,N_29780,N_28913);
nand UO_2636 (O_2636,N_29422,N_29071);
or UO_2637 (O_2637,N_29640,N_29728);
nor UO_2638 (O_2638,N_29025,N_28848);
nor UO_2639 (O_2639,N_29686,N_29731);
and UO_2640 (O_2640,N_28824,N_29173);
nor UO_2641 (O_2641,N_29048,N_29554);
and UO_2642 (O_2642,N_29200,N_29709);
nor UO_2643 (O_2643,N_28825,N_29072);
xnor UO_2644 (O_2644,N_28900,N_29472);
nand UO_2645 (O_2645,N_29527,N_29799);
xnor UO_2646 (O_2646,N_28866,N_29669);
and UO_2647 (O_2647,N_29893,N_29105);
xor UO_2648 (O_2648,N_29365,N_29716);
and UO_2649 (O_2649,N_29547,N_28938);
nor UO_2650 (O_2650,N_29003,N_29125);
and UO_2651 (O_2651,N_29147,N_29225);
nor UO_2652 (O_2652,N_29354,N_29159);
xor UO_2653 (O_2653,N_29496,N_29221);
and UO_2654 (O_2654,N_29102,N_29764);
nand UO_2655 (O_2655,N_29148,N_29352);
xor UO_2656 (O_2656,N_29432,N_29730);
nand UO_2657 (O_2657,N_29811,N_29947);
nor UO_2658 (O_2658,N_29333,N_28826);
xnor UO_2659 (O_2659,N_29392,N_29521);
xnor UO_2660 (O_2660,N_29771,N_29912);
and UO_2661 (O_2661,N_28957,N_28900);
nor UO_2662 (O_2662,N_29839,N_29524);
and UO_2663 (O_2663,N_28861,N_29621);
nor UO_2664 (O_2664,N_28985,N_29630);
and UO_2665 (O_2665,N_29640,N_29109);
nor UO_2666 (O_2666,N_29055,N_28838);
or UO_2667 (O_2667,N_29944,N_29491);
nor UO_2668 (O_2668,N_29314,N_29110);
and UO_2669 (O_2669,N_29810,N_29314);
or UO_2670 (O_2670,N_29991,N_29026);
and UO_2671 (O_2671,N_29975,N_29818);
or UO_2672 (O_2672,N_29912,N_29456);
and UO_2673 (O_2673,N_28811,N_29450);
nor UO_2674 (O_2674,N_29795,N_29152);
nand UO_2675 (O_2675,N_29602,N_29643);
nor UO_2676 (O_2676,N_28854,N_29922);
xor UO_2677 (O_2677,N_29481,N_29632);
xor UO_2678 (O_2678,N_29906,N_29945);
and UO_2679 (O_2679,N_29608,N_28992);
xor UO_2680 (O_2680,N_28887,N_29594);
and UO_2681 (O_2681,N_28846,N_29775);
and UO_2682 (O_2682,N_29815,N_29484);
nand UO_2683 (O_2683,N_29516,N_28907);
xnor UO_2684 (O_2684,N_29900,N_29665);
nor UO_2685 (O_2685,N_29893,N_29718);
nor UO_2686 (O_2686,N_29506,N_29950);
or UO_2687 (O_2687,N_29258,N_29799);
xnor UO_2688 (O_2688,N_29413,N_29637);
nor UO_2689 (O_2689,N_29359,N_29181);
and UO_2690 (O_2690,N_28921,N_29671);
nor UO_2691 (O_2691,N_29516,N_29470);
nand UO_2692 (O_2692,N_29307,N_29867);
or UO_2693 (O_2693,N_29786,N_28932);
and UO_2694 (O_2694,N_29776,N_29236);
xnor UO_2695 (O_2695,N_29366,N_29370);
and UO_2696 (O_2696,N_29711,N_29725);
nor UO_2697 (O_2697,N_29629,N_29800);
nor UO_2698 (O_2698,N_28859,N_28965);
or UO_2699 (O_2699,N_29903,N_29616);
or UO_2700 (O_2700,N_29757,N_28993);
xor UO_2701 (O_2701,N_29268,N_28928);
nand UO_2702 (O_2702,N_29247,N_28957);
nand UO_2703 (O_2703,N_29002,N_29682);
or UO_2704 (O_2704,N_29679,N_29962);
and UO_2705 (O_2705,N_29599,N_28830);
nor UO_2706 (O_2706,N_29575,N_29831);
xor UO_2707 (O_2707,N_29505,N_28992);
and UO_2708 (O_2708,N_29187,N_28890);
xnor UO_2709 (O_2709,N_29992,N_29373);
nand UO_2710 (O_2710,N_29378,N_28973);
or UO_2711 (O_2711,N_29932,N_29863);
or UO_2712 (O_2712,N_29588,N_29273);
nand UO_2713 (O_2713,N_29509,N_29432);
nand UO_2714 (O_2714,N_29732,N_29959);
and UO_2715 (O_2715,N_29601,N_29843);
nand UO_2716 (O_2716,N_29419,N_29942);
or UO_2717 (O_2717,N_28914,N_29190);
nor UO_2718 (O_2718,N_29531,N_29184);
nor UO_2719 (O_2719,N_29842,N_29641);
xor UO_2720 (O_2720,N_29146,N_29949);
and UO_2721 (O_2721,N_29449,N_29132);
nand UO_2722 (O_2722,N_29437,N_29600);
xnor UO_2723 (O_2723,N_29878,N_28812);
and UO_2724 (O_2724,N_29236,N_28992);
or UO_2725 (O_2725,N_28915,N_29961);
and UO_2726 (O_2726,N_29358,N_29750);
and UO_2727 (O_2727,N_29807,N_29077);
or UO_2728 (O_2728,N_29690,N_29653);
and UO_2729 (O_2729,N_29825,N_29565);
or UO_2730 (O_2730,N_29966,N_29677);
nor UO_2731 (O_2731,N_28827,N_29679);
nor UO_2732 (O_2732,N_29887,N_29415);
nand UO_2733 (O_2733,N_29999,N_28958);
and UO_2734 (O_2734,N_29864,N_29133);
or UO_2735 (O_2735,N_29382,N_28878);
or UO_2736 (O_2736,N_28996,N_29136);
nand UO_2737 (O_2737,N_29771,N_29975);
and UO_2738 (O_2738,N_29469,N_29053);
nor UO_2739 (O_2739,N_29696,N_29533);
and UO_2740 (O_2740,N_28803,N_29113);
nor UO_2741 (O_2741,N_29418,N_28810);
nand UO_2742 (O_2742,N_29192,N_29894);
or UO_2743 (O_2743,N_29364,N_28860);
nor UO_2744 (O_2744,N_29759,N_29512);
nand UO_2745 (O_2745,N_28826,N_29536);
nor UO_2746 (O_2746,N_29558,N_28816);
and UO_2747 (O_2747,N_29653,N_29364);
nor UO_2748 (O_2748,N_29332,N_29320);
or UO_2749 (O_2749,N_29894,N_29690);
and UO_2750 (O_2750,N_29676,N_29381);
nor UO_2751 (O_2751,N_29364,N_28886);
and UO_2752 (O_2752,N_29271,N_29438);
nor UO_2753 (O_2753,N_29158,N_29554);
nand UO_2754 (O_2754,N_29668,N_29645);
nand UO_2755 (O_2755,N_29344,N_29193);
and UO_2756 (O_2756,N_29904,N_29832);
nand UO_2757 (O_2757,N_29542,N_28917);
or UO_2758 (O_2758,N_28947,N_29094);
xor UO_2759 (O_2759,N_29694,N_29873);
or UO_2760 (O_2760,N_29353,N_29737);
and UO_2761 (O_2761,N_29810,N_29053);
or UO_2762 (O_2762,N_29283,N_29902);
or UO_2763 (O_2763,N_29929,N_29449);
xnor UO_2764 (O_2764,N_29155,N_29338);
nand UO_2765 (O_2765,N_29875,N_29475);
xor UO_2766 (O_2766,N_29938,N_29807);
or UO_2767 (O_2767,N_29766,N_28973);
xor UO_2768 (O_2768,N_29998,N_29639);
xor UO_2769 (O_2769,N_29595,N_29397);
and UO_2770 (O_2770,N_29333,N_29053);
or UO_2771 (O_2771,N_29999,N_29685);
nand UO_2772 (O_2772,N_29006,N_29839);
nor UO_2773 (O_2773,N_29374,N_29670);
nor UO_2774 (O_2774,N_29997,N_29613);
and UO_2775 (O_2775,N_29335,N_29340);
xor UO_2776 (O_2776,N_29074,N_29962);
xnor UO_2777 (O_2777,N_28975,N_29628);
xnor UO_2778 (O_2778,N_29023,N_29669);
and UO_2779 (O_2779,N_29834,N_29506);
and UO_2780 (O_2780,N_29929,N_28842);
nor UO_2781 (O_2781,N_29858,N_28895);
nor UO_2782 (O_2782,N_29085,N_29146);
nand UO_2783 (O_2783,N_29164,N_29695);
nor UO_2784 (O_2784,N_29209,N_29623);
nor UO_2785 (O_2785,N_29002,N_29104);
nor UO_2786 (O_2786,N_29591,N_29192);
or UO_2787 (O_2787,N_29278,N_29421);
and UO_2788 (O_2788,N_29782,N_29738);
nor UO_2789 (O_2789,N_29757,N_29524);
or UO_2790 (O_2790,N_29064,N_29217);
and UO_2791 (O_2791,N_28935,N_29861);
xnor UO_2792 (O_2792,N_28907,N_29785);
xor UO_2793 (O_2793,N_29418,N_29274);
and UO_2794 (O_2794,N_29368,N_28962);
and UO_2795 (O_2795,N_29328,N_29947);
and UO_2796 (O_2796,N_29525,N_29885);
or UO_2797 (O_2797,N_29362,N_29188);
and UO_2798 (O_2798,N_29552,N_28816);
or UO_2799 (O_2799,N_29987,N_29188);
nor UO_2800 (O_2800,N_28800,N_29638);
xnor UO_2801 (O_2801,N_29181,N_29868);
nor UO_2802 (O_2802,N_29250,N_29454);
nor UO_2803 (O_2803,N_29407,N_29739);
xnor UO_2804 (O_2804,N_28875,N_29064);
and UO_2805 (O_2805,N_29417,N_28804);
or UO_2806 (O_2806,N_28836,N_29568);
and UO_2807 (O_2807,N_29335,N_28893);
xnor UO_2808 (O_2808,N_28862,N_29537);
xor UO_2809 (O_2809,N_29555,N_29793);
and UO_2810 (O_2810,N_29215,N_29789);
xor UO_2811 (O_2811,N_29098,N_29417);
nand UO_2812 (O_2812,N_29500,N_29233);
or UO_2813 (O_2813,N_29727,N_29670);
xnor UO_2814 (O_2814,N_29405,N_29412);
nor UO_2815 (O_2815,N_29102,N_29792);
or UO_2816 (O_2816,N_29875,N_29004);
or UO_2817 (O_2817,N_29421,N_29312);
nor UO_2818 (O_2818,N_29896,N_29835);
or UO_2819 (O_2819,N_29794,N_29307);
or UO_2820 (O_2820,N_29795,N_29333);
nor UO_2821 (O_2821,N_29518,N_29884);
and UO_2822 (O_2822,N_29463,N_29948);
and UO_2823 (O_2823,N_29062,N_29415);
and UO_2824 (O_2824,N_29838,N_29569);
or UO_2825 (O_2825,N_28844,N_29088);
nor UO_2826 (O_2826,N_29957,N_29041);
xor UO_2827 (O_2827,N_28892,N_29789);
nand UO_2828 (O_2828,N_29058,N_29927);
and UO_2829 (O_2829,N_29293,N_29479);
and UO_2830 (O_2830,N_29441,N_29636);
or UO_2831 (O_2831,N_29496,N_29769);
nor UO_2832 (O_2832,N_29948,N_29597);
or UO_2833 (O_2833,N_29148,N_29773);
nand UO_2834 (O_2834,N_29246,N_28910);
xnor UO_2835 (O_2835,N_29628,N_28899);
xnor UO_2836 (O_2836,N_29430,N_29245);
and UO_2837 (O_2837,N_29104,N_29276);
nor UO_2838 (O_2838,N_29208,N_29675);
and UO_2839 (O_2839,N_29085,N_29375);
xor UO_2840 (O_2840,N_28983,N_29037);
nor UO_2841 (O_2841,N_29468,N_29083);
and UO_2842 (O_2842,N_29484,N_29202);
nor UO_2843 (O_2843,N_29362,N_29138);
xor UO_2844 (O_2844,N_29462,N_29053);
xnor UO_2845 (O_2845,N_29476,N_29871);
nor UO_2846 (O_2846,N_29877,N_29604);
nor UO_2847 (O_2847,N_29099,N_29498);
xnor UO_2848 (O_2848,N_29375,N_28858);
xor UO_2849 (O_2849,N_29693,N_29223);
and UO_2850 (O_2850,N_29805,N_29160);
nor UO_2851 (O_2851,N_29685,N_29333);
or UO_2852 (O_2852,N_28933,N_29246);
nor UO_2853 (O_2853,N_29240,N_29544);
or UO_2854 (O_2854,N_29045,N_28893);
nand UO_2855 (O_2855,N_29092,N_29839);
nand UO_2856 (O_2856,N_28972,N_28821);
nor UO_2857 (O_2857,N_29654,N_29533);
nand UO_2858 (O_2858,N_29105,N_28866);
and UO_2859 (O_2859,N_28877,N_29758);
or UO_2860 (O_2860,N_29942,N_29167);
nand UO_2861 (O_2861,N_29900,N_29526);
nand UO_2862 (O_2862,N_28843,N_29935);
nor UO_2863 (O_2863,N_29108,N_29430);
xnor UO_2864 (O_2864,N_29108,N_29840);
xnor UO_2865 (O_2865,N_29795,N_29187);
and UO_2866 (O_2866,N_29138,N_29365);
or UO_2867 (O_2867,N_28928,N_29731);
or UO_2868 (O_2868,N_29006,N_29032);
or UO_2869 (O_2869,N_29906,N_28927);
xnor UO_2870 (O_2870,N_29996,N_29156);
or UO_2871 (O_2871,N_29955,N_29006);
or UO_2872 (O_2872,N_29516,N_29464);
and UO_2873 (O_2873,N_29759,N_28990);
nand UO_2874 (O_2874,N_29546,N_28985);
xor UO_2875 (O_2875,N_29234,N_29394);
nand UO_2876 (O_2876,N_28984,N_28849);
or UO_2877 (O_2877,N_29990,N_29605);
nor UO_2878 (O_2878,N_29866,N_28993);
or UO_2879 (O_2879,N_28952,N_28917);
nand UO_2880 (O_2880,N_29709,N_29847);
nor UO_2881 (O_2881,N_29957,N_29057);
nand UO_2882 (O_2882,N_29720,N_29519);
and UO_2883 (O_2883,N_29875,N_29914);
and UO_2884 (O_2884,N_29005,N_29317);
and UO_2885 (O_2885,N_28983,N_29877);
nand UO_2886 (O_2886,N_29539,N_29353);
xor UO_2887 (O_2887,N_29743,N_29236);
nor UO_2888 (O_2888,N_29092,N_29736);
nand UO_2889 (O_2889,N_29581,N_28958);
nand UO_2890 (O_2890,N_29902,N_29349);
and UO_2891 (O_2891,N_29778,N_29596);
or UO_2892 (O_2892,N_29963,N_29772);
xor UO_2893 (O_2893,N_29521,N_29746);
xor UO_2894 (O_2894,N_29876,N_29855);
nor UO_2895 (O_2895,N_29019,N_29580);
and UO_2896 (O_2896,N_28894,N_29816);
nor UO_2897 (O_2897,N_29232,N_29202);
nand UO_2898 (O_2898,N_29678,N_29058);
or UO_2899 (O_2899,N_28800,N_29795);
and UO_2900 (O_2900,N_28841,N_28892);
or UO_2901 (O_2901,N_29235,N_29189);
nand UO_2902 (O_2902,N_29523,N_29154);
xnor UO_2903 (O_2903,N_29312,N_29099);
and UO_2904 (O_2904,N_29693,N_29248);
or UO_2905 (O_2905,N_29091,N_29494);
nand UO_2906 (O_2906,N_29727,N_29811);
xor UO_2907 (O_2907,N_28901,N_28980);
and UO_2908 (O_2908,N_29214,N_29615);
and UO_2909 (O_2909,N_29756,N_29415);
xnor UO_2910 (O_2910,N_29607,N_28944);
xnor UO_2911 (O_2911,N_28851,N_29051);
xor UO_2912 (O_2912,N_29505,N_29009);
nand UO_2913 (O_2913,N_29974,N_29814);
xnor UO_2914 (O_2914,N_29543,N_29200);
and UO_2915 (O_2915,N_29811,N_28985);
xor UO_2916 (O_2916,N_29440,N_29692);
and UO_2917 (O_2917,N_28839,N_29506);
or UO_2918 (O_2918,N_28866,N_28856);
nand UO_2919 (O_2919,N_29444,N_29552);
and UO_2920 (O_2920,N_29092,N_29903);
nor UO_2921 (O_2921,N_29947,N_29366);
or UO_2922 (O_2922,N_29749,N_28986);
nor UO_2923 (O_2923,N_29038,N_29216);
xnor UO_2924 (O_2924,N_29492,N_29445);
nand UO_2925 (O_2925,N_29804,N_29891);
xnor UO_2926 (O_2926,N_29154,N_29441);
or UO_2927 (O_2927,N_29291,N_28937);
nand UO_2928 (O_2928,N_29080,N_29007);
or UO_2929 (O_2929,N_29137,N_28897);
nand UO_2930 (O_2930,N_29896,N_29051);
nand UO_2931 (O_2931,N_29119,N_29866);
nor UO_2932 (O_2932,N_29457,N_29950);
nor UO_2933 (O_2933,N_29403,N_29933);
nor UO_2934 (O_2934,N_29924,N_28884);
xor UO_2935 (O_2935,N_29862,N_29598);
nand UO_2936 (O_2936,N_29203,N_29876);
nand UO_2937 (O_2937,N_29902,N_29838);
or UO_2938 (O_2938,N_28810,N_29247);
nand UO_2939 (O_2939,N_29787,N_29927);
nand UO_2940 (O_2940,N_28956,N_28990);
nor UO_2941 (O_2941,N_29834,N_29473);
nand UO_2942 (O_2942,N_29193,N_29702);
nand UO_2943 (O_2943,N_29598,N_28925);
and UO_2944 (O_2944,N_29417,N_29844);
nand UO_2945 (O_2945,N_29990,N_29568);
or UO_2946 (O_2946,N_29851,N_29801);
nor UO_2947 (O_2947,N_29656,N_29789);
nor UO_2948 (O_2948,N_28895,N_29742);
nand UO_2949 (O_2949,N_29131,N_29551);
nor UO_2950 (O_2950,N_29103,N_29026);
or UO_2951 (O_2951,N_29324,N_29566);
and UO_2952 (O_2952,N_28950,N_29931);
or UO_2953 (O_2953,N_29213,N_29517);
and UO_2954 (O_2954,N_29973,N_29305);
and UO_2955 (O_2955,N_29413,N_29262);
nand UO_2956 (O_2956,N_29298,N_29585);
and UO_2957 (O_2957,N_29154,N_29449);
xor UO_2958 (O_2958,N_29524,N_29351);
or UO_2959 (O_2959,N_29954,N_29927);
or UO_2960 (O_2960,N_28827,N_29736);
nor UO_2961 (O_2961,N_29555,N_29755);
xnor UO_2962 (O_2962,N_29488,N_29376);
and UO_2963 (O_2963,N_29892,N_29493);
nand UO_2964 (O_2964,N_29742,N_29216);
xor UO_2965 (O_2965,N_28847,N_29175);
or UO_2966 (O_2966,N_28835,N_29517);
nand UO_2967 (O_2967,N_29511,N_28873);
or UO_2968 (O_2968,N_29553,N_29996);
nand UO_2969 (O_2969,N_29114,N_29354);
nor UO_2970 (O_2970,N_29205,N_29557);
nand UO_2971 (O_2971,N_29267,N_29316);
and UO_2972 (O_2972,N_29708,N_28832);
and UO_2973 (O_2973,N_28979,N_29367);
nor UO_2974 (O_2974,N_29558,N_29615);
nor UO_2975 (O_2975,N_29150,N_29122);
xor UO_2976 (O_2976,N_28859,N_29607);
xnor UO_2977 (O_2977,N_29885,N_28802);
and UO_2978 (O_2978,N_28952,N_28920);
and UO_2979 (O_2979,N_29717,N_29442);
nand UO_2980 (O_2980,N_29668,N_29529);
xnor UO_2981 (O_2981,N_29087,N_29349);
xnor UO_2982 (O_2982,N_29494,N_29638);
nor UO_2983 (O_2983,N_29801,N_29427);
or UO_2984 (O_2984,N_29714,N_28917);
nand UO_2985 (O_2985,N_29610,N_29947);
or UO_2986 (O_2986,N_29025,N_29027);
or UO_2987 (O_2987,N_28995,N_28925);
and UO_2988 (O_2988,N_29531,N_29133);
xnor UO_2989 (O_2989,N_29126,N_29965);
and UO_2990 (O_2990,N_28931,N_29942);
xor UO_2991 (O_2991,N_29522,N_28934);
xnor UO_2992 (O_2992,N_28819,N_29047);
nand UO_2993 (O_2993,N_29457,N_29024);
and UO_2994 (O_2994,N_29441,N_29826);
or UO_2995 (O_2995,N_29545,N_28812);
nor UO_2996 (O_2996,N_29426,N_28815);
and UO_2997 (O_2997,N_29642,N_29682);
and UO_2998 (O_2998,N_28816,N_29091);
nor UO_2999 (O_2999,N_29092,N_29384);
xnor UO_3000 (O_3000,N_28907,N_29378);
or UO_3001 (O_3001,N_29370,N_29280);
and UO_3002 (O_3002,N_28940,N_29657);
or UO_3003 (O_3003,N_29422,N_28917);
nand UO_3004 (O_3004,N_29737,N_28913);
nand UO_3005 (O_3005,N_29261,N_28856);
and UO_3006 (O_3006,N_28863,N_29020);
xnor UO_3007 (O_3007,N_29177,N_29754);
nand UO_3008 (O_3008,N_29045,N_29199);
nand UO_3009 (O_3009,N_29988,N_29178);
and UO_3010 (O_3010,N_29461,N_29376);
and UO_3011 (O_3011,N_29190,N_28847);
or UO_3012 (O_3012,N_29605,N_29194);
nor UO_3013 (O_3013,N_29304,N_29351);
nand UO_3014 (O_3014,N_29957,N_29380);
nor UO_3015 (O_3015,N_29426,N_29900);
nand UO_3016 (O_3016,N_29601,N_29217);
nor UO_3017 (O_3017,N_29385,N_29695);
xnor UO_3018 (O_3018,N_29102,N_28975);
and UO_3019 (O_3019,N_29728,N_28805);
or UO_3020 (O_3020,N_29333,N_29809);
and UO_3021 (O_3021,N_29375,N_29555);
and UO_3022 (O_3022,N_29613,N_29304);
or UO_3023 (O_3023,N_29419,N_29132);
xnor UO_3024 (O_3024,N_29632,N_29191);
nand UO_3025 (O_3025,N_29530,N_29280);
xor UO_3026 (O_3026,N_29551,N_29231);
and UO_3027 (O_3027,N_29157,N_29615);
and UO_3028 (O_3028,N_29503,N_29353);
xnor UO_3029 (O_3029,N_28924,N_29983);
nor UO_3030 (O_3030,N_29358,N_29244);
nor UO_3031 (O_3031,N_29005,N_29484);
xor UO_3032 (O_3032,N_29901,N_29543);
or UO_3033 (O_3033,N_29079,N_29677);
or UO_3034 (O_3034,N_29651,N_29928);
and UO_3035 (O_3035,N_29689,N_29903);
or UO_3036 (O_3036,N_29884,N_28869);
nor UO_3037 (O_3037,N_29354,N_29043);
xnor UO_3038 (O_3038,N_29096,N_29324);
nor UO_3039 (O_3039,N_29020,N_28859);
nand UO_3040 (O_3040,N_29132,N_29284);
or UO_3041 (O_3041,N_28863,N_28901);
nor UO_3042 (O_3042,N_29532,N_29658);
nand UO_3043 (O_3043,N_29941,N_28953);
nand UO_3044 (O_3044,N_29007,N_29396);
xor UO_3045 (O_3045,N_29953,N_29949);
xor UO_3046 (O_3046,N_29013,N_29375);
nand UO_3047 (O_3047,N_29669,N_29054);
nand UO_3048 (O_3048,N_29276,N_28861);
nor UO_3049 (O_3049,N_29488,N_28913);
nand UO_3050 (O_3050,N_29330,N_29708);
nor UO_3051 (O_3051,N_29786,N_29962);
and UO_3052 (O_3052,N_29947,N_29483);
nand UO_3053 (O_3053,N_29886,N_29690);
nand UO_3054 (O_3054,N_28852,N_29234);
nor UO_3055 (O_3055,N_29846,N_29485);
nor UO_3056 (O_3056,N_29367,N_29911);
nor UO_3057 (O_3057,N_28984,N_29107);
or UO_3058 (O_3058,N_29945,N_29055);
nor UO_3059 (O_3059,N_29273,N_29302);
nor UO_3060 (O_3060,N_29636,N_28979);
nand UO_3061 (O_3061,N_29765,N_29665);
nor UO_3062 (O_3062,N_29404,N_29193);
and UO_3063 (O_3063,N_29481,N_28987);
nor UO_3064 (O_3064,N_29397,N_29407);
nor UO_3065 (O_3065,N_28872,N_29536);
nor UO_3066 (O_3066,N_28873,N_29958);
or UO_3067 (O_3067,N_29365,N_29264);
nand UO_3068 (O_3068,N_29449,N_29578);
nand UO_3069 (O_3069,N_29125,N_29234);
or UO_3070 (O_3070,N_28980,N_29564);
and UO_3071 (O_3071,N_28940,N_29468);
or UO_3072 (O_3072,N_29112,N_29191);
and UO_3073 (O_3073,N_29074,N_28918);
nand UO_3074 (O_3074,N_29019,N_29149);
nor UO_3075 (O_3075,N_29599,N_28836);
nor UO_3076 (O_3076,N_29241,N_29805);
nor UO_3077 (O_3077,N_29811,N_29983);
and UO_3078 (O_3078,N_29718,N_29358);
or UO_3079 (O_3079,N_28882,N_29835);
nor UO_3080 (O_3080,N_29686,N_29276);
or UO_3081 (O_3081,N_29366,N_29687);
nand UO_3082 (O_3082,N_29462,N_29307);
nand UO_3083 (O_3083,N_29230,N_29434);
or UO_3084 (O_3084,N_29899,N_29705);
nor UO_3085 (O_3085,N_29437,N_29508);
and UO_3086 (O_3086,N_28970,N_29785);
nor UO_3087 (O_3087,N_29777,N_29774);
nor UO_3088 (O_3088,N_29529,N_28827);
xor UO_3089 (O_3089,N_29050,N_29621);
nor UO_3090 (O_3090,N_29758,N_29406);
or UO_3091 (O_3091,N_29295,N_29516);
xor UO_3092 (O_3092,N_29504,N_29780);
nand UO_3093 (O_3093,N_29069,N_29234);
and UO_3094 (O_3094,N_29573,N_28801);
and UO_3095 (O_3095,N_29720,N_29948);
nor UO_3096 (O_3096,N_29416,N_29134);
or UO_3097 (O_3097,N_29967,N_29150);
and UO_3098 (O_3098,N_29383,N_29150);
nor UO_3099 (O_3099,N_29369,N_29770);
or UO_3100 (O_3100,N_29500,N_29206);
and UO_3101 (O_3101,N_29317,N_29274);
and UO_3102 (O_3102,N_29581,N_29014);
or UO_3103 (O_3103,N_29980,N_29547);
and UO_3104 (O_3104,N_29356,N_29954);
nand UO_3105 (O_3105,N_29533,N_29483);
or UO_3106 (O_3106,N_29691,N_29397);
or UO_3107 (O_3107,N_29929,N_28860);
nand UO_3108 (O_3108,N_29578,N_29816);
xnor UO_3109 (O_3109,N_29712,N_28998);
nand UO_3110 (O_3110,N_29999,N_28819);
or UO_3111 (O_3111,N_29164,N_29524);
or UO_3112 (O_3112,N_29261,N_29237);
and UO_3113 (O_3113,N_29384,N_29793);
or UO_3114 (O_3114,N_29026,N_29055);
xor UO_3115 (O_3115,N_29602,N_29961);
nand UO_3116 (O_3116,N_29197,N_29102);
and UO_3117 (O_3117,N_29629,N_29405);
or UO_3118 (O_3118,N_29319,N_29212);
nand UO_3119 (O_3119,N_28924,N_29365);
and UO_3120 (O_3120,N_28831,N_29416);
nor UO_3121 (O_3121,N_29338,N_29589);
xnor UO_3122 (O_3122,N_29697,N_29902);
and UO_3123 (O_3123,N_29359,N_29907);
xnor UO_3124 (O_3124,N_28945,N_29126);
xor UO_3125 (O_3125,N_29183,N_28917);
nand UO_3126 (O_3126,N_29666,N_29862);
nor UO_3127 (O_3127,N_29689,N_29527);
and UO_3128 (O_3128,N_29637,N_29718);
xnor UO_3129 (O_3129,N_29711,N_29982);
nand UO_3130 (O_3130,N_29229,N_29410);
nand UO_3131 (O_3131,N_29597,N_28851);
or UO_3132 (O_3132,N_28841,N_28921);
nor UO_3133 (O_3133,N_29948,N_29933);
xor UO_3134 (O_3134,N_28955,N_28992);
and UO_3135 (O_3135,N_29268,N_29278);
nor UO_3136 (O_3136,N_28981,N_28969);
xor UO_3137 (O_3137,N_28882,N_29219);
and UO_3138 (O_3138,N_29592,N_29458);
nand UO_3139 (O_3139,N_29597,N_29885);
nand UO_3140 (O_3140,N_28928,N_28836);
xnor UO_3141 (O_3141,N_29890,N_28978);
nand UO_3142 (O_3142,N_29388,N_28907);
and UO_3143 (O_3143,N_29459,N_29603);
xor UO_3144 (O_3144,N_29697,N_29743);
xnor UO_3145 (O_3145,N_29967,N_29189);
nor UO_3146 (O_3146,N_29753,N_28931);
nor UO_3147 (O_3147,N_29802,N_28992);
or UO_3148 (O_3148,N_29952,N_29824);
or UO_3149 (O_3149,N_29419,N_29312);
or UO_3150 (O_3150,N_28828,N_29112);
xor UO_3151 (O_3151,N_29183,N_29850);
xor UO_3152 (O_3152,N_29932,N_29477);
and UO_3153 (O_3153,N_29826,N_29474);
xnor UO_3154 (O_3154,N_28970,N_29334);
xor UO_3155 (O_3155,N_28875,N_28849);
or UO_3156 (O_3156,N_29366,N_29685);
xor UO_3157 (O_3157,N_29899,N_29116);
nand UO_3158 (O_3158,N_29038,N_29219);
nor UO_3159 (O_3159,N_29150,N_29897);
xnor UO_3160 (O_3160,N_29435,N_29672);
xnor UO_3161 (O_3161,N_29206,N_29210);
and UO_3162 (O_3162,N_28935,N_29931);
or UO_3163 (O_3163,N_29239,N_29138);
nor UO_3164 (O_3164,N_29206,N_29333);
or UO_3165 (O_3165,N_29110,N_29691);
nor UO_3166 (O_3166,N_28985,N_28818);
and UO_3167 (O_3167,N_29776,N_29865);
and UO_3168 (O_3168,N_29985,N_29880);
and UO_3169 (O_3169,N_28806,N_29788);
and UO_3170 (O_3170,N_29646,N_29592);
or UO_3171 (O_3171,N_29818,N_29258);
and UO_3172 (O_3172,N_29749,N_29104);
xor UO_3173 (O_3173,N_29249,N_29362);
and UO_3174 (O_3174,N_29658,N_29700);
nor UO_3175 (O_3175,N_29929,N_28851);
nor UO_3176 (O_3176,N_28888,N_29651);
nand UO_3177 (O_3177,N_29291,N_29493);
xnor UO_3178 (O_3178,N_29881,N_29663);
nand UO_3179 (O_3179,N_29182,N_29719);
and UO_3180 (O_3180,N_28865,N_29001);
and UO_3181 (O_3181,N_29391,N_29988);
nor UO_3182 (O_3182,N_29197,N_29623);
xor UO_3183 (O_3183,N_29068,N_28866);
xnor UO_3184 (O_3184,N_29972,N_28984);
and UO_3185 (O_3185,N_29742,N_29866);
xnor UO_3186 (O_3186,N_29081,N_29213);
or UO_3187 (O_3187,N_29432,N_29409);
nor UO_3188 (O_3188,N_29697,N_29374);
xor UO_3189 (O_3189,N_29702,N_29848);
xnor UO_3190 (O_3190,N_29069,N_28972);
or UO_3191 (O_3191,N_29128,N_29028);
or UO_3192 (O_3192,N_28973,N_29859);
or UO_3193 (O_3193,N_28958,N_29386);
nand UO_3194 (O_3194,N_29032,N_29961);
and UO_3195 (O_3195,N_28845,N_29316);
nor UO_3196 (O_3196,N_29938,N_29292);
nor UO_3197 (O_3197,N_29933,N_29020);
nand UO_3198 (O_3198,N_28821,N_29928);
or UO_3199 (O_3199,N_28842,N_29877);
xnor UO_3200 (O_3200,N_28857,N_29563);
and UO_3201 (O_3201,N_29841,N_29867);
xor UO_3202 (O_3202,N_29930,N_29002);
and UO_3203 (O_3203,N_28830,N_28969);
or UO_3204 (O_3204,N_29026,N_29583);
nor UO_3205 (O_3205,N_29625,N_29802);
nor UO_3206 (O_3206,N_29757,N_29129);
and UO_3207 (O_3207,N_29147,N_29643);
xor UO_3208 (O_3208,N_29005,N_29618);
nand UO_3209 (O_3209,N_29022,N_29055);
nor UO_3210 (O_3210,N_29398,N_29620);
nand UO_3211 (O_3211,N_29320,N_28916);
xnor UO_3212 (O_3212,N_29597,N_28832);
or UO_3213 (O_3213,N_29616,N_28891);
nor UO_3214 (O_3214,N_29965,N_29801);
nand UO_3215 (O_3215,N_28816,N_29991);
or UO_3216 (O_3216,N_29466,N_28800);
and UO_3217 (O_3217,N_28987,N_29954);
xor UO_3218 (O_3218,N_29487,N_28863);
or UO_3219 (O_3219,N_29565,N_29078);
xnor UO_3220 (O_3220,N_29143,N_29801);
nor UO_3221 (O_3221,N_29734,N_29511);
xor UO_3222 (O_3222,N_29849,N_29825);
xor UO_3223 (O_3223,N_29169,N_29024);
and UO_3224 (O_3224,N_29284,N_28906);
and UO_3225 (O_3225,N_29954,N_29799);
and UO_3226 (O_3226,N_29619,N_28875);
nor UO_3227 (O_3227,N_28952,N_28869);
nand UO_3228 (O_3228,N_29406,N_29448);
and UO_3229 (O_3229,N_29692,N_29488);
or UO_3230 (O_3230,N_29640,N_29264);
nor UO_3231 (O_3231,N_29470,N_29057);
nand UO_3232 (O_3232,N_29603,N_29460);
or UO_3233 (O_3233,N_28972,N_29216);
xnor UO_3234 (O_3234,N_29737,N_29514);
or UO_3235 (O_3235,N_29005,N_29983);
nand UO_3236 (O_3236,N_28834,N_29182);
nor UO_3237 (O_3237,N_29620,N_28948);
nand UO_3238 (O_3238,N_28838,N_29402);
nor UO_3239 (O_3239,N_29365,N_29578);
nand UO_3240 (O_3240,N_28923,N_29746);
and UO_3241 (O_3241,N_29408,N_29009);
and UO_3242 (O_3242,N_29242,N_29952);
or UO_3243 (O_3243,N_28979,N_28905);
xnor UO_3244 (O_3244,N_28841,N_29407);
and UO_3245 (O_3245,N_29132,N_29748);
and UO_3246 (O_3246,N_29237,N_28986);
and UO_3247 (O_3247,N_29973,N_29237);
or UO_3248 (O_3248,N_29240,N_29774);
nor UO_3249 (O_3249,N_29211,N_29137);
and UO_3250 (O_3250,N_29921,N_29806);
nand UO_3251 (O_3251,N_29728,N_29264);
nand UO_3252 (O_3252,N_28940,N_28841);
or UO_3253 (O_3253,N_29006,N_29045);
and UO_3254 (O_3254,N_29303,N_29619);
nor UO_3255 (O_3255,N_29977,N_29998);
or UO_3256 (O_3256,N_29412,N_29086);
and UO_3257 (O_3257,N_29102,N_29121);
or UO_3258 (O_3258,N_28903,N_29854);
or UO_3259 (O_3259,N_29575,N_29863);
nand UO_3260 (O_3260,N_29968,N_29196);
xor UO_3261 (O_3261,N_28855,N_29142);
nand UO_3262 (O_3262,N_29751,N_29249);
xnor UO_3263 (O_3263,N_29226,N_29318);
nor UO_3264 (O_3264,N_28806,N_29427);
nand UO_3265 (O_3265,N_28951,N_28901);
xnor UO_3266 (O_3266,N_29653,N_28959);
xnor UO_3267 (O_3267,N_29728,N_29497);
and UO_3268 (O_3268,N_29665,N_28886);
or UO_3269 (O_3269,N_29096,N_29809);
nor UO_3270 (O_3270,N_29784,N_29866);
xnor UO_3271 (O_3271,N_29034,N_28802);
nand UO_3272 (O_3272,N_29652,N_28890);
xnor UO_3273 (O_3273,N_28812,N_29337);
nor UO_3274 (O_3274,N_29340,N_29155);
nor UO_3275 (O_3275,N_28956,N_28808);
nor UO_3276 (O_3276,N_29479,N_29328);
nor UO_3277 (O_3277,N_29777,N_29566);
nor UO_3278 (O_3278,N_28999,N_29696);
and UO_3279 (O_3279,N_28845,N_29501);
nand UO_3280 (O_3280,N_29259,N_29529);
nand UO_3281 (O_3281,N_29777,N_29888);
nor UO_3282 (O_3282,N_29273,N_29611);
nand UO_3283 (O_3283,N_29648,N_29697);
nor UO_3284 (O_3284,N_29969,N_29173);
xor UO_3285 (O_3285,N_29041,N_29673);
xor UO_3286 (O_3286,N_28899,N_29611);
xnor UO_3287 (O_3287,N_29139,N_28946);
xor UO_3288 (O_3288,N_29782,N_29406);
and UO_3289 (O_3289,N_29581,N_29989);
xor UO_3290 (O_3290,N_29335,N_29580);
nand UO_3291 (O_3291,N_28923,N_29949);
or UO_3292 (O_3292,N_29135,N_29536);
xor UO_3293 (O_3293,N_28892,N_29124);
nor UO_3294 (O_3294,N_29437,N_29642);
and UO_3295 (O_3295,N_29736,N_29390);
and UO_3296 (O_3296,N_29496,N_29603);
xor UO_3297 (O_3297,N_28854,N_29069);
and UO_3298 (O_3298,N_29004,N_29548);
or UO_3299 (O_3299,N_29587,N_29329);
or UO_3300 (O_3300,N_29042,N_29188);
and UO_3301 (O_3301,N_28897,N_29184);
nor UO_3302 (O_3302,N_29513,N_29762);
nand UO_3303 (O_3303,N_29650,N_29777);
nor UO_3304 (O_3304,N_29861,N_29460);
xor UO_3305 (O_3305,N_29281,N_29599);
nand UO_3306 (O_3306,N_29815,N_29681);
xnor UO_3307 (O_3307,N_29956,N_28956);
and UO_3308 (O_3308,N_29647,N_29967);
xor UO_3309 (O_3309,N_29382,N_28922);
xnor UO_3310 (O_3310,N_29723,N_29812);
nor UO_3311 (O_3311,N_29569,N_29432);
nand UO_3312 (O_3312,N_29078,N_29304);
nor UO_3313 (O_3313,N_28803,N_29873);
nand UO_3314 (O_3314,N_28870,N_29305);
xor UO_3315 (O_3315,N_29025,N_28956);
and UO_3316 (O_3316,N_28869,N_29976);
nand UO_3317 (O_3317,N_29926,N_28827);
nand UO_3318 (O_3318,N_29019,N_29485);
nor UO_3319 (O_3319,N_29154,N_29579);
or UO_3320 (O_3320,N_29662,N_29650);
nor UO_3321 (O_3321,N_29291,N_28896);
nand UO_3322 (O_3322,N_29872,N_29909);
or UO_3323 (O_3323,N_29641,N_29028);
nor UO_3324 (O_3324,N_28826,N_29075);
and UO_3325 (O_3325,N_29760,N_29855);
nand UO_3326 (O_3326,N_29196,N_29407);
xor UO_3327 (O_3327,N_29445,N_28939);
nor UO_3328 (O_3328,N_29466,N_29504);
and UO_3329 (O_3329,N_29798,N_29755);
and UO_3330 (O_3330,N_29387,N_29356);
nor UO_3331 (O_3331,N_29140,N_28969);
or UO_3332 (O_3332,N_29173,N_29398);
nor UO_3333 (O_3333,N_29857,N_29211);
or UO_3334 (O_3334,N_29475,N_29047);
nand UO_3335 (O_3335,N_28828,N_29829);
and UO_3336 (O_3336,N_28910,N_28948);
xnor UO_3337 (O_3337,N_29001,N_29626);
and UO_3338 (O_3338,N_29061,N_29114);
or UO_3339 (O_3339,N_28953,N_29516);
or UO_3340 (O_3340,N_29196,N_29690);
xor UO_3341 (O_3341,N_29740,N_29976);
and UO_3342 (O_3342,N_29295,N_28832);
nor UO_3343 (O_3343,N_29013,N_29861);
and UO_3344 (O_3344,N_29923,N_29881);
nor UO_3345 (O_3345,N_28948,N_29830);
xor UO_3346 (O_3346,N_29910,N_29472);
nand UO_3347 (O_3347,N_29911,N_29859);
xor UO_3348 (O_3348,N_29445,N_29571);
or UO_3349 (O_3349,N_29751,N_28949);
and UO_3350 (O_3350,N_29871,N_29891);
nand UO_3351 (O_3351,N_29170,N_29708);
nor UO_3352 (O_3352,N_29155,N_29825);
and UO_3353 (O_3353,N_29811,N_29497);
or UO_3354 (O_3354,N_29362,N_29038);
nand UO_3355 (O_3355,N_29315,N_29253);
nand UO_3356 (O_3356,N_29373,N_28830);
nor UO_3357 (O_3357,N_29118,N_29229);
nand UO_3358 (O_3358,N_29871,N_29485);
xor UO_3359 (O_3359,N_29383,N_29035);
nand UO_3360 (O_3360,N_28905,N_28972);
nor UO_3361 (O_3361,N_29355,N_29806);
or UO_3362 (O_3362,N_29593,N_29255);
and UO_3363 (O_3363,N_29951,N_29061);
xnor UO_3364 (O_3364,N_29576,N_28831);
nor UO_3365 (O_3365,N_28977,N_29238);
nor UO_3366 (O_3366,N_29591,N_29462);
xnor UO_3367 (O_3367,N_29134,N_29754);
xnor UO_3368 (O_3368,N_29852,N_29486);
xor UO_3369 (O_3369,N_28842,N_28878);
or UO_3370 (O_3370,N_29081,N_29419);
nand UO_3371 (O_3371,N_29853,N_29820);
xnor UO_3372 (O_3372,N_29868,N_29774);
and UO_3373 (O_3373,N_29021,N_29543);
or UO_3374 (O_3374,N_29971,N_29009);
nand UO_3375 (O_3375,N_29984,N_29351);
and UO_3376 (O_3376,N_28845,N_29471);
xnor UO_3377 (O_3377,N_29940,N_29691);
xor UO_3378 (O_3378,N_29139,N_29986);
and UO_3379 (O_3379,N_29473,N_29431);
or UO_3380 (O_3380,N_28927,N_29342);
xnor UO_3381 (O_3381,N_28807,N_28875);
xor UO_3382 (O_3382,N_29880,N_29707);
xor UO_3383 (O_3383,N_29352,N_29601);
or UO_3384 (O_3384,N_29849,N_28865);
xor UO_3385 (O_3385,N_29199,N_28887);
nand UO_3386 (O_3386,N_29887,N_29339);
nor UO_3387 (O_3387,N_29193,N_29490);
nand UO_3388 (O_3388,N_29133,N_29484);
xnor UO_3389 (O_3389,N_29716,N_29128);
xnor UO_3390 (O_3390,N_29806,N_28840);
nand UO_3391 (O_3391,N_29329,N_29790);
and UO_3392 (O_3392,N_29528,N_29415);
and UO_3393 (O_3393,N_29018,N_29560);
or UO_3394 (O_3394,N_28862,N_29385);
or UO_3395 (O_3395,N_29990,N_29191);
xor UO_3396 (O_3396,N_29791,N_29542);
nand UO_3397 (O_3397,N_29416,N_29040);
nand UO_3398 (O_3398,N_29219,N_29139);
nor UO_3399 (O_3399,N_28870,N_29464);
or UO_3400 (O_3400,N_29874,N_29270);
nand UO_3401 (O_3401,N_29585,N_29867);
nand UO_3402 (O_3402,N_29296,N_29507);
nand UO_3403 (O_3403,N_29016,N_29043);
xor UO_3404 (O_3404,N_28975,N_28878);
nor UO_3405 (O_3405,N_29484,N_29493);
nor UO_3406 (O_3406,N_29129,N_28877);
nor UO_3407 (O_3407,N_29008,N_28918);
xnor UO_3408 (O_3408,N_29920,N_28821);
nor UO_3409 (O_3409,N_29873,N_28908);
or UO_3410 (O_3410,N_28857,N_29775);
or UO_3411 (O_3411,N_29349,N_29919);
and UO_3412 (O_3412,N_28874,N_29552);
and UO_3413 (O_3413,N_29106,N_29216);
and UO_3414 (O_3414,N_29044,N_29692);
nor UO_3415 (O_3415,N_29532,N_29228);
or UO_3416 (O_3416,N_29326,N_29353);
and UO_3417 (O_3417,N_28988,N_29022);
nand UO_3418 (O_3418,N_29644,N_29753);
nand UO_3419 (O_3419,N_29081,N_29602);
and UO_3420 (O_3420,N_29735,N_29626);
nor UO_3421 (O_3421,N_29295,N_29051);
and UO_3422 (O_3422,N_28948,N_29076);
nor UO_3423 (O_3423,N_29074,N_29158);
nand UO_3424 (O_3424,N_29790,N_29516);
xor UO_3425 (O_3425,N_29588,N_29436);
or UO_3426 (O_3426,N_28937,N_29860);
nand UO_3427 (O_3427,N_29249,N_28945);
nand UO_3428 (O_3428,N_29942,N_29201);
nand UO_3429 (O_3429,N_29133,N_29927);
and UO_3430 (O_3430,N_29017,N_29724);
nand UO_3431 (O_3431,N_29185,N_29274);
nand UO_3432 (O_3432,N_29502,N_29977);
nand UO_3433 (O_3433,N_29702,N_28888);
and UO_3434 (O_3434,N_28964,N_29566);
and UO_3435 (O_3435,N_28942,N_29772);
xor UO_3436 (O_3436,N_29517,N_29470);
nor UO_3437 (O_3437,N_29780,N_29024);
or UO_3438 (O_3438,N_29138,N_28919);
nand UO_3439 (O_3439,N_29687,N_29230);
and UO_3440 (O_3440,N_29331,N_29965);
nand UO_3441 (O_3441,N_28959,N_29839);
and UO_3442 (O_3442,N_28821,N_28901);
xor UO_3443 (O_3443,N_29101,N_29756);
xor UO_3444 (O_3444,N_29774,N_29050);
or UO_3445 (O_3445,N_29105,N_28945);
nand UO_3446 (O_3446,N_29026,N_29840);
nand UO_3447 (O_3447,N_29715,N_29300);
nand UO_3448 (O_3448,N_29269,N_28945);
and UO_3449 (O_3449,N_28880,N_29341);
and UO_3450 (O_3450,N_29457,N_29380);
or UO_3451 (O_3451,N_29568,N_29388);
xnor UO_3452 (O_3452,N_29975,N_29534);
or UO_3453 (O_3453,N_29206,N_29576);
xor UO_3454 (O_3454,N_29679,N_28907);
and UO_3455 (O_3455,N_28832,N_29223);
or UO_3456 (O_3456,N_29637,N_29810);
nor UO_3457 (O_3457,N_29767,N_29569);
xor UO_3458 (O_3458,N_29760,N_29078);
nor UO_3459 (O_3459,N_29785,N_29275);
nor UO_3460 (O_3460,N_29089,N_29630);
nand UO_3461 (O_3461,N_29196,N_28824);
and UO_3462 (O_3462,N_29841,N_29748);
or UO_3463 (O_3463,N_28880,N_29599);
xnor UO_3464 (O_3464,N_29374,N_29833);
nand UO_3465 (O_3465,N_29297,N_29262);
xor UO_3466 (O_3466,N_29590,N_29275);
and UO_3467 (O_3467,N_29879,N_29253);
and UO_3468 (O_3468,N_29745,N_29757);
nand UO_3469 (O_3469,N_29815,N_29609);
and UO_3470 (O_3470,N_29273,N_29827);
xnor UO_3471 (O_3471,N_29625,N_29972);
or UO_3472 (O_3472,N_28876,N_29619);
nor UO_3473 (O_3473,N_29817,N_29052);
xor UO_3474 (O_3474,N_29519,N_29138);
nor UO_3475 (O_3475,N_29739,N_29863);
nand UO_3476 (O_3476,N_29998,N_29523);
nand UO_3477 (O_3477,N_29775,N_29692);
nor UO_3478 (O_3478,N_29201,N_28840);
xnor UO_3479 (O_3479,N_29613,N_29186);
xnor UO_3480 (O_3480,N_29543,N_29774);
nand UO_3481 (O_3481,N_29915,N_29254);
nand UO_3482 (O_3482,N_28978,N_29783);
and UO_3483 (O_3483,N_29783,N_29420);
or UO_3484 (O_3484,N_29349,N_29951);
or UO_3485 (O_3485,N_29885,N_28949);
nand UO_3486 (O_3486,N_28946,N_28815);
nor UO_3487 (O_3487,N_29716,N_29396);
xor UO_3488 (O_3488,N_29337,N_29957);
nor UO_3489 (O_3489,N_28862,N_28997);
or UO_3490 (O_3490,N_28937,N_29862);
nand UO_3491 (O_3491,N_29591,N_29679);
or UO_3492 (O_3492,N_29978,N_29927);
or UO_3493 (O_3493,N_29280,N_29045);
nor UO_3494 (O_3494,N_28934,N_28827);
nand UO_3495 (O_3495,N_29862,N_29654);
xor UO_3496 (O_3496,N_29204,N_29487);
and UO_3497 (O_3497,N_29351,N_29857);
nor UO_3498 (O_3498,N_29892,N_29453);
xnor UO_3499 (O_3499,N_29421,N_29225);
endmodule