module basic_1000_10000_1500_4_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_461,In_130);
and U1 (N_1,In_47,In_348);
and U2 (N_2,In_413,In_531);
nor U3 (N_3,In_734,In_139);
nand U4 (N_4,In_396,In_924);
and U5 (N_5,In_470,In_925);
nand U6 (N_6,In_509,In_443);
or U7 (N_7,In_576,In_215);
xnor U8 (N_8,In_595,In_195);
nand U9 (N_9,In_326,In_119);
or U10 (N_10,In_568,In_567);
or U11 (N_11,In_952,In_503);
nor U12 (N_12,In_175,In_863);
xor U13 (N_13,In_279,In_214);
nor U14 (N_14,In_494,In_502);
nand U15 (N_15,In_76,In_23);
nor U16 (N_16,In_149,In_821);
and U17 (N_17,In_106,In_29);
and U18 (N_18,In_479,In_169);
nand U19 (N_19,In_517,In_935);
nand U20 (N_20,In_844,In_71);
nand U21 (N_21,In_220,In_719);
and U22 (N_22,In_336,In_242);
nand U23 (N_23,In_520,In_310);
or U24 (N_24,In_137,In_757);
and U25 (N_25,In_832,In_624);
or U26 (N_26,In_362,In_14);
or U27 (N_27,In_401,In_53);
nand U28 (N_28,In_392,In_825);
and U29 (N_29,In_616,In_631);
nor U30 (N_30,In_269,In_706);
or U31 (N_31,In_620,In_405);
nand U32 (N_32,In_113,In_627);
or U33 (N_33,In_493,In_906);
nand U34 (N_34,In_155,In_231);
or U35 (N_35,In_801,In_635);
xor U36 (N_36,In_30,In_355);
or U37 (N_37,In_538,In_417);
and U38 (N_38,In_94,In_575);
and U39 (N_39,In_323,In_835);
nor U40 (N_40,In_349,In_982);
and U41 (N_41,In_889,In_274);
nand U42 (N_42,In_448,In_344);
nor U43 (N_43,In_721,In_217);
or U44 (N_44,In_696,In_725);
or U45 (N_45,In_459,In_219);
and U46 (N_46,In_16,In_146);
nor U47 (N_47,In_630,In_668);
nor U48 (N_48,In_92,In_181);
nand U49 (N_49,In_587,In_415);
and U50 (N_50,In_34,In_565);
nor U51 (N_51,In_147,In_312);
nand U52 (N_52,In_903,In_720);
and U53 (N_53,In_643,In_255);
or U54 (N_54,In_601,In_177);
or U55 (N_55,In_171,In_954);
xor U56 (N_56,In_915,In_290);
and U57 (N_57,In_340,In_324);
or U58 (N_58,In_790,In_816);
nor U59 (N_59,In_506,In_179);
and U60 (N_60,In_875,In_841);
xor U61 (N_61,In_427,In_500);
or U62 (N_62,In_917,In_793);
nor U63 (N_63,In_986,In_868);
nor U64 (N_64,In_920,In_385);
and U65 (N_65,In_588,In_383);
and U66 (N_66,In_4,In_865);
and U67 (N_67,In_291,In_884);
nand U68 (N_68,In_619,In_846);
nor U69 (N_69,In_537,In_948);
or U70 (N_70,In_881,In_225);
and U71 (N_71,In_960,In_354);
nor U72 (N_72,In_745,In_968);
nand U73 (N_73,In_495,In_295);
and U74 (N_74,In_153,In_446);
nor U75 (N_75,In_22,In_545);
nand U76 (N_76,In_781,In_359);
and U77 (N_77,In_553,In_338);
or U78 (N_78,In_686,In_776);
and U79 (N_79,In_655,In_683);
and U80 (N_80,In_270,In_339);
nand U81 (N_81,In_398,In_423);
and U82 (N_82,In_899,In_918);
nor U83 (N_83,In_833,In_947);
and U84 (N_84,In_561,In_2);
nor U85 (N_85,In_484,In_133);
nor U86 (N_86,In_662,In_714);
nor U87 (N_87,In_964,In_300);
nand U88 (N_88,In_919,In_834);
or U89 (N_89,In_931,In_275);
or U90 (N_90,In_458,In_281);
or U91 (N_91,In_442,In_328);
nand U92 (N_92,In_411,In_285);
and U93 (N_93,In_582,In_513);
or U94 (N_94,In_792,In_928);
nand U95 (N_95,In_307,In_987);
nor U96 (N_96,In_700,In_253);
nand U97 (N_97,In_173,In_318);
nand U98 (N_98,In_89,In_969);
nor U99 (N_99,In_838,In_572);
xnor U100 (N_100,In_604,In_432);
and U101 (N_101,In_247,In_739);
or U102 (N_102,In_425,In_456);
nor U103 (N_103,In_967,In_439);
or U104 (N_104,In_334,In_901);
or U105 (N_105,In_638,In_666);
and U106 (N_106,In_994,In_806);
and U107 (N_107,In_970,In_262);
nand U108 (N_108,In_74,In_729);
nor U109 (N_109,In_202,In_100);
nor U110 (N_110,In_560,In_224);
nor U111 (N_111,In_164,In_775);
nor U112 (N_112,In_497,In_937);
and U113 (N_113,In_539,In_436);
xor U114 (N_114,In_356,In_43);
nand U115 (N_115,In_90,In_256);
or U116 (N_116,In_286,In_17);
nand U117 (N_117,In_434,In_910);
or U118 (N_118,In_187,In_867);
and U119 (N_119,In_52,In_56);
or U120 (N_120,In_777,In_883);
or U121 (N_121,In_73,In_407);
nand U122 (N_122,In_871,In_813);
nand U123 (N_123,In_730,In_496);
nor U124 (N_124,In_1,In_942);
and U125 (N_125,In_346,In_649);
or U126 (N_126,In_563,In_699);
or U127 (N_127,In_950,In_228);
nand U128 (N_128,In_264,In_268);
or U129 (N_129,In_266,In_756);
nand U130 (N_130,In_988,In_684);
nand U131 (N_131,In_91,In_112);
nand U132 (N_132,In_265,In_337);
xnor U133 (N_133,In_872,In_64);
nand U134 (N_134,In_449,In_261);
nor U135 (N_135,In_523,In_11);
nor U136 (N_136,In_465,In_70);
nor U137 (N_137,In_174,In_606);
and U138 (N_138,In_957,In_254);
or U139 (N_139,In_653,In_273);
nor U140 (N_140,In_753,In_235);
or U141 (N_141,In_898,In_276);
or U142 (N_142,In_140,In_232);
nor U143 (N_143,In_473,In_156);
or U144 (N_144,In_239,In_124);
nand U145 (N_145,In_380,In_311);
nand U146 (N_146,In_85,In_505);
or U147 (N_147,In_430,In_193);
nand U148 (N_148,In_573,In_977);
and U149 (N_149,In_900,In_783);
or U150 (N_150,In_626,In_812);
or U151 (N_151,In_934,In_599);
and U152 (N_152,In_853,In_851);
and U153 (N_153,In_404,In_460);
nor U154 (N_154,In_358,In_656);
or U155 (N_155,In_759,In_475);
nor U156 (N_156,In_543,In_804);
nand U157 (N_157,In_603,In_252);
nor U158 (N_158,In_305,In_444);
or U159 (N_159,In_250,In_972);
nor U160 (N_160,In_75,In_612);
nand U161 (N_161,In_379,In_660);
nand U162 (N_162,In_211,In_368);
or U163 (N_163,In_760,In_746);
and U164 (N_164,In_99,In_774);
or U165 (N_165,In_766,In_207);
nand U166 (N_166,In_319,In_611);
nand U167 (N_167,In_25,In_257);
or U168 (N_168,In_490,In_617);
xnor U169 (N_169,In_909,In_20);
or U170 (N_170,In_194,In_516);
or U171 (N_171,In_105,In_586);
nand U172 (N_172,In_514,In_571);
or U173 (N_173,In_912,In_787);
or U174 (N_174,In_382,In_747);
or U175 (N_175,In_882,In_6);
nand U176 (N_176,In_913,In_511);
nand U177 (N_177,In_679,In_839);
and U178 (N_178,In_546,In_88);
nand U179 (N_179,In_208,In_389);
nand U180 (N_180,In_40,In_908);
nand U181 (N_181,In_72,In_132);
and U182 (N_182,In_711,In_698);
nand U183 (N_183,In_372,In_751);
nor U184 (N_184,In_600,In_96);
nand U185 (N_185,In_188,In_245);
nand U186 (N_186,In_705,In_773);
nand U187 (N_187,In_707,In_938);
nor U188 (N_188,In_694,In_81);
nand U189 (N_189,In_42,In_672);
or U190 (N_190,In_248,In_157);
or U191 (N_191,In_975,In_243);
nand U192 (N_192,In_953,In_518);
or U193 (N_193,In_779,In_366);
or U194 (N_194,In_158,In_159);
nand U195 (N_195,In_750,In_763);
nand U196 (N_196,In_134,In_65);
nand U197 (N_197,In_229,In_690);
nor U198 (N_198,In_552,In_594);
nor U199 (N_199,In_384,In_284);
or U200 (N_200,In_670,In_847);
nand U201 (N_201,In_388,In_367);
nand U202 (N_202,In_877,In_689);
nor U203 (N_203,In_507,In_302);
and U204 (N_204,In_170,In_429);
or U205 (N_205,In_386,In_301);
and U206 (N_206,In_361,In_550);
or U207 (N_207,In_184,In_421);
and U208 (N_208,In_226,In_141);
nand U209 (N_209,In_549,In_309);
xnor U210 (N_210,In_870,In_980);
or U211 (N_211,In_559,In_457);
or U212 (N_212,In_765,In_412);
and U213 (N_213,In_722,In_534);
nand U214 (N_214,In_77,In_44);
nor U215 (N_215,In_165,In_657);
nor U216 (N_216,In_241,In_272);
and U217 (N_217,In_941,In_86);
or U218 (N_218,In_921,In_350);
or U219 (N_219,In_795,In_330);
or U220 (N_220,In_395,In_28);
nand U221 (N_221,In_422,In_916);
nor U222 (N_222,In_152,In_24);
nor U223 (N_223,In_732,In_907);
or U224 (N_224,In_403,In_237);
nand U225 (N_225,In_244,In_956);
or U226 (N_226,In_97,In_842);
nand U227 (N_227,In_393,In_370);
and U228 (N_228,In_451,In_201);
nand U229 (N_229,In_713,In_435);
nand U230 (N_230,In_84,In_373);
and U231 (N_231,In_431,In_428);
and U232 (N_232,In_930,In_377);
and U233 (N_233,In_15,In_823);
and U234 (N_234,In_827,In_166);
nor U235 (N_235,In_80,In_440);
nand U236 (N_236,In_331,In_961);
or U237 (N_237,In_267,In_597);
and U238 (N_238,In_332,In_569);
xnor U239 (N_239,In_778,In_196);
nand U240 (N_240,In_605,In_408);
or U241 (N_241,In_51,In_891);
and U242 (N_242,In_692,In_129);
or U243 (N_243,In_607,In_127);
nand U244 (N_244,In_817,In_876);
nand U245 (N_245,In_946,In_66);
nor U246 (N_246,In_914,In_79);
nor U247 (N_247,In_659,In_820);
or U248 (N_248,In_258,In_593);
nor U249 (N_249,In_136,In_249);
nor U250 (N_250,In_525,In_394);
and U251 (N_251,In_693,In_645);
nor U252 (N_252,In_399,In_259);
and U253 (N_253,In_848,In_789);
nor U254 (N_254,In_357,In_260);
nand U255 (N_255,In_993,In_117);
or U256 (N_256,In_618,In_862);
xnor U257 (N_257,In_168,In_973);
and U258 (N_258,In_271,In_676);
nor U259 (N_259,In_723,In_125);
and U260 (N_260,In_409,In_151);
nor U261 (N_261,In_251,In_880);
nor U262 (N_262,In_890,In_691);
and U263 (N_263,In_376,In_548);
or U264 (N_264,In_929,In_727);
nor U265 (N_265,In_658,In_850);
and U266 (N_266,In_740,In_221);
and U267 (N_267,In_62,In_210);
or U268 (N_268,In_297,In_426);
nor U269 (N_269,In_116,In_574);
or U270 (N_270,In_454,In_3);
nor U271 (N_271,In_788,In_533);
nand U272 (N_272,In_615,In_885);
nand U273 (N_273,In_752,In_845);
and U274 (N_274,In_621,In_866);
nor U275 (N_275,In_38,In_744);
and U276 (N_276,In_735,In_83);
and U277 (N_277,In_191,In_445);
nand U278 (N_278,In_512,In_628);
or U279 (N_279,In_748,In_375);
and U280 (N_280,In_887,In_489);
nor U281 (N_281,In_327,In_542);
nand U282 (N_282,In_785,In_222);
and U283 (N_283,In_837,In_410);
nand U284 (N_284,In_858,In_562);
and U285 (N_285,In_483,In_768);
and U286 (N_286,In_487,In_755);
nand U287 (N_287,In_37,In_308);
nor U288 (N_288,In_192,In_115);
and U289 (N_289,In_577,In_701);
nor U290 (N_290,In_855,In_936);
and U291 (N_291,In_227,In_161);
and U292 (N_292,In_927,In_182);
nand U293 (N_293,In_702,In_717);
or U294 (N_294,In_236,In_63);
and U295 (N_295,In_122,In_809);
or U296 (N_296,In_922,In_772);
nor U297 (N_297,In_68,In_18);
nor U298 (N_298,In_828,In_680);
nor U299 (N_299,In_992,In_642);
nand U300 (N_300,In_485,In_447);
nand U301 (N_301,In_737,In_144);
and U302 (N_302,In_478,In_59);
and U303 (N_303,In_976,In_61);
or U304 (N_304,In_498,In_200);
and U305 (N_305,In_945,In_78);
nand U306 (N_306,In_540,In_886);
nand U307 (N_307,In_704,In_861);
nand U308 (N_308,In_199,In_892);
nand U309 (N_309,In_761,In_49);
nand U310 (N_310,In_148,In_849);
and U311 (N_311,In_397,In_39);
nor U312 (N_312,In_360,In_613);
and U313 (N_313,In_904,In_424);
and U314 (N_314,In_869,In_767);
nor U315 (N_315,In_646,In_476);
or U316 (N_316,In_82,In_418);
or U317 (N_317,In_263,In_299);
xor U318 (N_318,In_598,In_374);
or U319 (N_319,In_27,In_864);
nand U320 (N_320,In_283,In_771);
nor U321 (N_321,In_897,In_536);
and U322 (N_322,In_715,In_831);
or U323 (N_323,In_710,In_530);
and U324 (N_324,In_278,In_304);
nand U325 (N_325,In_316,In_7);
nand U326 (N_326,In_9,In_280);
nor U327 (N_327,In_118,In_19);
nand U328 (N_328,In_547,In_488);
nor U329 (N_329,In_329,In_162);
or U330 (N_330,In_733,In_364);
nor U331 (N_331,In_321,In_60);
and U332 (N_332,In_230,In_145);
nand U333 (N_333,In_854,In_183);
or U334 (N_334,In_325,In_896);
and U335 (N_335,In_639,In_469);
and U336 (N_336,In_420,In_802);
and U337 (N_337,In_629,In_450);
or U338 (N_338,In_341,In_799);
or U339 (N_339,In_819,In_176);
or U340 (N_340,In_591,In_589);
or U341 (N_341,In_371,In_180);
and U342 (N_342,In_48,In_623);
nand U343 (N_343,In_622,In_36);
nand U344 (N_344,In_45,In_26);
nor U345 (N_345,In_979,In_138);
nand U346 (N_346,In_58,In_167);
nor U347 (N_347,In_189,In_570);
and U348 (N_348,In_87,In_579);
or U349 (N_349,In_741,In_492);
or U350 (N_350,In_32,In_682);
or U351 (N_351,In_378,In_762);
nand U352 (N_352,In_150,In_438);
nand U353 (N_353,In_142,In_528);
nor U354 (N_354,In_963,In_472);
nand U355 (N_355,In_69,In_474);
or U356 (N_356,In_654,In_209);
or U357 (N_357,In_716,In_240);
nand U358 (N_358,In_190,In_213);
or U359 (N_359,In_35,In_633);
or U360 (N_360,In_798,In_829);
nor U361 (N_361,In_135,In_958);
nand U362 (N_362,In_955,In_997);
xor U363 (N_363,In_160,In_856);
or U364 (N_364,In_402,In_471);
or U365 (N_365,In_31,In_218);
nand U366 (N_366,In_857,In_554);
nor U367 (N_367,In_671,In_452);
and U368 (N_368,In_102,In_453);
nand U369 (N_369,In_437,In_205);
or U370 (N_370,In_878,In_647);
nor U371 (N_371,In_555,In_313);
nand U372 (N_372,In_351,In_641);
or U373 (N_373,In_352,In_566);
or U374 (N_374,In_104,In_499);
nand U375 (N_375,In_126,In_998);
xor U376 (N_376,In_780,In_584);
or U377 (N_377,In_482,In_852);
nand U378 (N_378,In_894,In_664);
or U379 (N_379,In_681,In_669);
nor U380 (N_380,In_298,In_527);
nor U381 (N_381,In_650,In_433);
nand U382 (N_382,In_592,In_121);
nand U383 (N_383,In_640,In_808);
and U384 (N_384,In_932,In_971);
nand U385 (N_385,In_246,In_673);
nor U386 (N_386,In_55,In_455);
nand U387 (N_387,In_962,In_391);
nand U388 (N_388,In_983,In_108);
nor U389 (N_389,In_288,In_991);
nor U390 (N_390,In_50,In_365);
and U391 (N_391,In_466,In_416);
or U392 (N_392,In_462,In_46);
nand U393 (N_393,In_107,In_902);
and U394 (N_394,In_811,In_687);
nand U395 (N_395,In_708,In_728);
nor U396 (N_396,In_782,In_441);
nand U397 (N_397,In_840,In_933);
nor U398 (N_398,In_477,In_754);
nand U399 (N_399,In_178,In_709);
nor U400 (N_400,In_939,In_984);
nor U401 (N_401,In_419,In_342);
nand U402 (N_402,In_109,In_335);
nand U403 (N_403,In_390,In_926);
or U404 (N_404,In_414,In_712);
nor U405 (N_405,In_197,In_738);
nor U406 (N_406,In_749,In_667);
and U407 (N_407,In_726,In_282);
nor U408 (N_408,In_491,In_67);
nor U409 (N_409,In_363,In_293);
or U410 (N_410,In_836,In_648);
nor U411 (N_411,In_287,In_557);
nand U412 (N_412,In_843,In_791);
nor U413 (N_413,In_501,In_0);
nor U414 (N_414,In_532,In_508);
or U415 (N_415,In_602,In_524);
nor U416 (N_416,In_21,In_590);
or U417 (N_417,In_103,In_810);
or U418 (N_418,In_480,In_303);
and U419 (N_419,In_999,In_223);
and U420 (N_420,In_185,In_989);
nand U421 (N_421,In_685,In_204);
and U422 (N_422,In_541,In_625);
or U423 (N_423,In_556,In_238);
nand U424 (N_424,In_12,In_347);
nor U425 (N_425,In_292,In_203);
and U426 (N_426,In_381,In_990);
and U427 (N_427,In_911,In_564);
nand U428 (N_428,In_544,In_558);
and U429 (N_429,In_940,In_369);
nor U430 (N_430,In_10,In_526);
and U431 (N_431,In_551,In_467);
nor U432 (N_432,In_959,In_614);
or U433 (N_433,In_212,In_943);
nor U434 (N_434,In_172,In_296);
or U435 (N_435,In_110,In_873);
and U436 (N_436,In_859,In_944);
nand U437 (N_437,In_677,In_529);
or U438 (N_438,In_803,In_974);
nand U439 (N_439,In_981,In_652);
and U440 (N_440,In_128,In_784);
or U441 (N_441,In_826,In_805);
nor U442 (N_442,In_651,In_198);
nand U443 (N_443,In_54,In_665);
nand U444 (N_444,In_905,In_98);
and U445 (N_445,In_632,In_688);
nor U446 (N_446,In_521,In_233);
or U447 (N_447,In_95,In_695);
nand U448 (N_448,In_101,In_5);
or U449 (N_449,In_464,In_468);
nor U450 (N_450,In_277,In_731);
or U451 (N_451,In_515,In_736);
or U452 (N_452,In_874,In_41);
or U453 (N_453,In_504,In_314);
or U454 (N_454,In_661,In_797);
or U455 (N_455,In_345,In_578);
nand U456 (N_456,In_895,In_581);
or U457 (N_457,In_678,In_522);
and U458 (N_458,In_486,In_609);
nand U459 (N_459,In_758,In_343);
nor U460 (N_460,In_786,In_814);
or U461 (N_461,In_234,In_93);
nand U462 (N_462,In_718,In_674);
nor U463 (N_463,In_114,In_519);
or U464 (N_464,In_830,In_294);
nor U465 (N_465,In_923,In_996);
and U466 (N_466,In_57,In_965);
and U467 (N_467,In_800,In_610);
and U468 (N_468,In_123,In_703);
nor U469 (N_469,In_815,In_306);
nor U470 (N_470,In_966,In_13);
nand U471 (N_471,In_387,In_949);
and U472 (N_472,In_481,In_644);
nand U473 (N_473,In_636,In_216);
and U474 (N_474,In_697,In_580);
and U475 (N_475,In_317,In_186);
or U476 (N_476,In_995,In_807);
and U477 (N_477,In_608,In_888);
and U478 (N_478,In_206,In_353);
and U479 (N_479,In_315,In_879);
nand U480 (N_480,In_743,In_818);
and U481 (N_481,In_893,In_333);
nand U482 (N_482,In_33,In_724);
and U483 (N_483,In_583,In_860);
and U484 (N_484,In_794,In_663);
nand U485 (N_485,In_596,In_764);
nand U486 (N_486,In_796,In_742);
nor U487 (N_487,In_120,In_634);
nor U488 (N_488,In_322,In_985);
nor U489 (N_489,In_769,In_675);
nor U490 (N_490,In_637,In_289);
nor U491 (N_491,In_154,In_585);
nand U492 (N_492,In_400,In_978);
or U493 (N_493,In_951,In_111);
or U494 (N_494,In_463,In_143);
nor U495 (N_495,In_822,In_535);
or U496 (N_496,In_131,In_163);
or U497 (N_497,In_8,In_406);
and U498 (N_498,In_510,In_320);
and U499 (N_499,In_770,In_824);
nand U500 (N_500,In_488,In_928);
nand U501 (N_501,In_342,In_697);
or U502 (N_502,In_129,In_216);
or U503 (N_503,In_500,In_492);
or U504 (N_504,In_36,In_853);
nor U505 (N_505,In_137,In_539);
nor U506 (N_506,In_620,In_988);
nand U507 (N_507,In_653,In_639);
and U508 (N_508,In_660,In_977);
nor U509 (N_509,In_851,In_208);
nand U510 (N_510,In_439,In_670);
nor U511 (N_511,In_165,In_78);
nor U512 (N_512,In_827,In_964);
nor U513 (N_513,In_286,In_876);
and U514 (N_514,In_820,In_166);
or U515 (N_515,In_987,In_574);
nor U516 (N_516,In_581,In_973);
or U517 (N_517,In_183,In_631);
xor U518 (N_518,In_347,In_67);
or U519 (N_519,In_474,In_303);
nand U520 (N_520,In_139,In_310);
and U521 (N_521,In_869,In_892);
or U522 (N_522,In_341,In_490);
xor U523 (N_523,In_75,In_638);
nor U524 (N_524,In_796,In_921);
nand U525 (N_525,In_16,In_587);
nand U526 (N_526,In_670,In_65);
nor U527 (N_527,In_918,In_417);
nor U528 (N_528,In_178,In_259);
or U529 (N_529,In_770,In_336);
or U530 (N_530,In_436,In_456);
nand U531 (N_531,In_290,In_876);
nand U532 (N_532,In_253,In_855);
or U533 (N_533,In_227,In_756);
nand U534 (N_534,In_865,In_339);
nor U535 (N_535,In_694,In_127);
nor U536 (N_536,In_552,In_879);
xnor U537 (N_537,In_510,In_49);
nand U538 (N_538,In_894,In_778);
or U539 (N_539,In_889,In_336);
or U540 (N_540,In_719,In_37);
and U541 (N_541,In_212,In_299);
nor U542 (N_542,In_878,In_577);
and U543 (N_543,In_531,In_792);
or U544 (N_544,In_934,In_686);
nand U545 (N_545,In_328,In_45);
and U546 (N_546,In_745,In_782);
and U547 (N_547,In_457,In_742);
or U548 (N_548,In_190,In_41);
and U549 (N_549,In_615,In_382);
or U550 (N_550,In_911,In_358);
nand U551 (N_551,In_275,In_58);
or U552 (N_552,In_640,In_910);
and U553 (N_553,In_516,In_969);
and U554 (N_554,In_949,In_683);
and U555 (N_555,In_268,In_376);
or U556 (N_556,In_660,In_779);
nor U557 (N_557,In_315,In_309);
nand U558 (N_558,In_976,In_517);
or U559 (N_559,In_892,In_324);
and U560 (N_560,In_42,In_555);
or U561 (N_561,In_947,In_862);
and U562 (N_562,In_201,In_987);
and U563 (N_563,In_769,In_253);
xnor U564 (N_564,In_538,In_575);
or U565 (N_565,In_307,In_891);
and U566 (N_566,In_568,In_883);
nand U567 (N_567,In_487,In_500);
nor U568 (N_568,In_150,In_617);
or U569 (N_569,In_607,In_378);
and U570 (N_570,In_570,In_397);
nand U571 (N_571,In_925,In_444);
nand U572 (N_572,In_680,In_685);
nor U573 (N_573,In_297,In_520);
and U574 (N_574,In_79,In_672);
nand U575 (N_575,In_671,In_434);
or U576 (N_576,In_334,In_11);
or U577 (N_577,In_842,In_394);
and U578 (N_578,In_137,In_678);
and U579 (N_579,In_993,In_454);
nand U580 (N_580,In_673,In_542);
nor U581 (N_581,In_142,In_986);
nor U582 (N_582,In_230,In_630);
or U583 (N_583,In_738,In_408);
or U584 (N_584,In_851,In_166);
or U585 (N_585,In_672,In_848);
or U586 (N_586,In_566,In_911);
or U587 (N_587,In_788,In_91);
nor U588 (N_588,In_472,In_911);
nor U589 (N_589,In_251,In_281);
and U590 (N_590,In_26,In_413);
and U591 (N_591,In_490,In_577);
and U592 (N_592,In_153,In_480);
and U593 (N_593,In_842,In_366);
nand U594 (N_594,In_62,In_851);
xnor U595 (N_595,In_97,In_592);
nor U596 (N_596,In_968,In_343);
nor U597 (N_597,In_676,In_217);
or U598 (N_598,In_5,In_892);
and U599 (N_599,In_452,In_611);
and U600 (N_600,In_578,In_747);
and U601 (N_601,In_439,In_804);
or U602 (N_602,In_495,In_294);
nand U603 (N_603,In_785,In_879);
and U604 (N_604,In_997,In_638);
and U605 (N_605,In_828,In_755);
or U606 (N_606,In_530,In_936);
and U607 (N_607,In_236,In_798);
nor U608 (N_608,In_537,In_443);
and U609 (N_609,In_663,In_179);
nor U610 (N_610,In_745,In_25);
and U611 (N_611,In_506,In_589);
or U612 (N_612,In_402,In_501);
or U613 (N_613,In_113,In_528);
and U614 (N_614,In_600,In_402);
and U615 (N_615,In_95,In_412);
or U616 (N_616,In_896,In_903);
nor U617 (N_617,In_222,In_315);
and U618 (N_618,In_95,In_210);
nor U619 (N_619,In_129,In_56);
nor U620 (N_620,In_205,In_680);
and U621 (N_621,In_386,In_293);
and U622 (N_622,In_967,In_15);
or U623 (N_623,In_437,In_470);
and U624 (N_624,In_801,In_618);
and U625 (N_625,In_980,In_319);
or U626 (N_626,In_704,In_732);
and U627 (N_627,In_7,In_401);
or U628 (N_628,In_64,In_10);
nand U629 (N_629,In_933,In_884);
or U630 (N_630,In_964,In_170);
or U631 (N_631,In_597,In_940);
nand U632 (N_632,In_808,In_481);
nor U633 (N_633,In_776,In_870);
nor U634 (N_634,In_435,In_327);
nand U635 (N_635,In_203,In_600);
nor U636 (N_636,In_22,In_357);
or U637 (N_637,In_482,In_301);
nor U638 (N_638,In_414,In_390);
or U639 (N_639,In_320,In_153);
nand U640 (N_640,In_279,In_662);
nand U641 (N_641,In_407,In_109);
or U642 (N_642,In_759,In_303);
nor U643 (N_643,In_231,In_84);
xor U644 (N_644,In_916,In_349);
nand U645 (N_645,In_890,In_571);
and U646 (N_646,In_431,In_503);
and U647 (N_647,In_156,In_572);
or U648 (N_648,In_916,In_753);
nand U649 (N_649,In_808,In_329);
nor U650 (N_650,In_64,In_57);
nor U651 (N_651,In_421,In_101);
nand U652 (N_652,In_248,In_406);
and U653 (N_653,In_0,In_135);
nand U654 (N_654,In_177,In_896);
nand U655 (N_655,In_944,In_963);
and U656 (N_656,In_171,In_3);
or U657 (N_657,In_728,In_280);
nand U658 (N_658,In_409,In_169);
or U659 (N_659,In_122,In_213);
and U660 (N_660,In_323,In_348);
and U661 (N_661,In_115,In_842);
or U662 (N_662,In_866,In_994);
or U663 (N_663,In_787,In_264);
or U664 (N_664,In_678,In_378);
or U665 (N_665,In_311,In_435);
and U666 (N_666,In_558,In_506);
and U667 (N_667,In_343,In_225);
or U668 (N_668,In_487,In_581);
nor U669 (N_669,In_714,In_625);
and U670 (N_670,In_388,In_645);
nand U671 (N_671,In_50,In_74);
and U672 (N_672,In_937,In_407);
or U673 (N_673,In_974,In_863);
nor U674 (N_674,In_688,In_165);
and U675 (N_675,In_509,In_720);
nor U676 (N_676,In_124,In_791);
xor U677 (N_677,In_334,In_592);
nor U678 (N_678,In_13,In_368);
or U679 (N_679,In_567,In_465);
nor U680 (N_680,In_57,In_680);
nand U681 (N_681,In_768,In_210);
nand U682 (N_682,In_352,In_530);
nand U683 (N_683,In_213,In_818);
nor U684 (N_684,In_290,In_248);
nand U685 (N_685,In_150,In_927);
nor U686 (N_686,In_196,In_675);
nand U687 (N_687,In_74,In_253);
nand U688 (N_688,In_363,In_193);
or U689 (N_689,In_489,In_626);
or U690 (N_690,In_465,In_236);
nand U691 (N_691,In_451,In_370);
nor U692 (N_692,In_779,In_822);
nand U693 (N_693,In_333,In_214);
and U694 (N_694,In_840,In_581);
nand U695 (N_695,In_273,In_105);
and U696 (N_696,In_440,In_317);
nor U697 (N_697,In_609,In_716);
or U698 (N_698,In_663,In_956);
nor U699 (N_699,In_396,In_71);
nor U700 (N_700,In_355,In_510);
nand U701 (N_701,In_148,In_514);
and U702 (N_702,In_590,In_306);
nand U703 (N_703,In_198,In_173);
xnor U704 (N_704,In_441,In_740);
and U705 (N_705,In_646,In_462);
or U706 (N_706,In_74,In_689);
or U707 (N_707,In_484,In_168);
nand U708 (N_708,In_329,In_545);
and U709 (N_709,In_941,In_704);
or U710 (N_710,In_544,In_385);
nor U711 (N_711,In_741,In_811);
nand U712 (N_712,In_858,In_213);
or U713 (N_713,In_968,In_580);
or U714 (N_714,In_824,In_698);
nand U715 (N_715,In_257,In_603);
or U716 (N_716,In_937,In_801);
nand U717 (N_717,In_276,In_20);
nand U718 (N_718,In_367,In_996);
and U719 (N_719,In_430,In_387);
and U720 (N_720,In_67,In_709);
and U721 (N_721,In_428,In_732);
nand U722 (N_722,In_702,In_533);
nand U723 (N_723,In_400,In_93);
nand U724 (N_724,In_950,In_516);
nand U725 (N_725,In_839,In_75);
or U726 (N_726,In_957,In_786);
or U727 (N_727,In_288,In_306);
or U728 (N_728,In_491,In_462);
nor U729 (N_729,In_858,In_628);
nand U730 (N_730,In_376,In_740);
or U731 (N_731,In_286,In_423);
nand U732 (N_732,In_266,In_291);
nand U733 (N_733,In_198,In_905);
nor U734 (N_734,In_658,In_765);
and U735 (N_735,In_832,In_687);
nand U736 (N_736,In_289,In_791);
nand U737 (N_737,In_120,In_291);
nor U738 (N_738,In_188,In_164);
or U739 (N_739,In_753,In_925);
or U740 (N_740,In_886,In_448);
or U741 (N_741,In_427,In_401);
and U742 (N_742,In_250,In_882);
nand U743 (N_743,In_29,In_430);
and U744 (N_744,In_979,In_778);
or U745 (N_745,In_238,In_771);
nor U746 (N_746,In_696,In_239);
nor U747 (N_747,In_361,In_904);
or U748 (N_748,In_379,In_392);
nand U749 (N_749,In_551,In_319);
or U750 (N_750,In_677,In_769);
and U751 (N_751,In_363,In_665);
nor U752 (N_752,In_948,In_285);
or U753 (N_753,In_907,In_347);
nand U754 (N_754,In_753,In_596);
nor U755 (N_755,In_505,In_225);
nand U756 (N_756,In_724,In_545);
and U757 (N_757,In_607,In_848);
nor U758 (N_758,In_272,In_229);
or U759 (N_759,In_424,In_98);
nand U760 (N_760,In_610,In_52);
nand U761 (N_761,In_281,In_693);
or U762 (N_762,In_157,In_986);
and U763 (N_763,In_746,In_46);
xnor U764 (N_764,In_194,In_949);
or U765 (N_765,In_163,In_372);
nor U766 (N_766,In_686,In_287);
or U767 (N_767,In_589,In_537);
and U768 (N_768,In_878,In_640);
xnor U769 (N_769,In_346,In_693);
or U770 (N_770,In_755,In_883);
nor U771 (N_771,In_506,In_85);
and U772 (N_772,In_347,In_412);
nor U773 (N_773,In_331,In_650);
and U774 (N_774,In_939,In_130);
or U775 (N_775,In_380,In_782);
or U776 (N_776,In_145,In_113);
nand U777 (N_777,In_42,In_177);
or U778 (N_778,In_448,In_368);
or U779 (N_779,In_841,In_408);
nand U780 (N_780,In_902,In_25);
nand U781 (N_781,In_721,In_611);
or U782 (N_782,In_795,In_676);
nand U783 (N_783,In_274,In_360);
and U784 (N_784,In_306,In_312);
nand U785 (N_785,In_857,In_933);
or U786 (N_786,In_773,In_323);
xnor U787 (N_787,In_554,In_419);
and U788 (N_788,In_260,In_821);
nor U789 (N_789,In_926,In_391);
nor U790 (N_790,In_423,In_807);
nor U791 (N_791,In_240,In_362);
nand U792 (N_792,In_249,In_985);
nor U793 (N_793,In_682,In_823);
nor U794 (N_794,In_775,In_144);
nand U795 (N_795,In_547,In_897);
or U796 (N_796,In_150,In_970);
nor U797 (N_797,In_491,In_181);
and U798 (N_798,In_62,In_980);
nor U799 (N_799,In_483,In_122);
and U800 (N_800,In_722,In_899);
or U801 (N_801,In_944,In_867);
nand U802 (N_802,In_6,In_552);
or U803 (N_803,In_887,In_361);
nor U804 (N_804,In_807,In_33);
nor U805 (N_805,In_528,In_841);
nor U806 (N_806,In_586,In_493);
nor U807 (N_807,In_613,In_190);
nor U808 (N_808,In_279,In_803);
nand U809 (N_809,In_248,In_100);
or U810 (N_810,In_864,In_9);
nor U811 (N_811,In_619,In_524);
nor U812 (N_812,In_531,In_552);
nand U813 (N_813,In_330,In_962);
and U814 (N_814,In_583,In_743);
nand U815 (N_815,In_316,In_593);
and U816 (N_816,In_936,In_681);
nand U817 (N_817,In_912,In_250);
and U818 (N_818,In_972,In_596);
xnor U819 (N_819,In_603,In_290);
nor U820 (N_820,In_79,In_487);
and U821 (N_821,In_843,In_687);
nor U822 (N_822,In_24,In_986);
or U823 (N_823,In_325,In_476);
or U824 (N_824,In_6,In_832);
and U825 (N_825,In_857,In_213);
and U826 (N_826,In_895,In_204);
or U827 (N_827,In_994,In_460);
nand U828 (N_828,In_450,In_395);
or U829 (N_829,In_524,In_228);
or U830 (N_830,In_701,In_839);
and U831 (N_831,In_670,In_494);
nor U832 (N_832,In_178,In_634);
nand U833 (N_833,In_402,In_702);
or U834 (N_834,In_130,In_719);
and U835 (N_835,In_322,In_917);
nand U836 (N_836,In_775,In_476);
or U837 (N_837,In_302,In_328);
or U838 (N_838,In_824,In_540);
or U839 (N_839,In_390,In_55);
nand U840 (N_840,In_252,In_577);
or U841 (N_841,In_3,In_465);
or U842 (N_842,In_880,In_309);
nand U843 (N_843,In_844,In_985);
nand U844 (N_844,In_789,In_967);
and U845 (N_845,In_991,In_793);
nor U846 (N_846,In_172,In_369);
and U847 (N_847,In_916,In_999);
and U848 (N_848,In_335,In_788);
or U849 (N_849,In_117,In_818);
nor U850 (N_850,In_824,In_251);
nand U851 (N_851,In_835,In_500);
and U852 (N_852,In_881,In_981);
or U853 (N_853,In_991,In_563);
nand U854 (N_854,In_614,In_225);
and U855 (N_855,In_944,In_422);
or U856 (N_856,In_175,In_141);
nor U857 (N_857,In_739,In_74);
or U858 (N_858,In_716,In_942);
nor U859 (N_859,In_72,In_178);
nor U860 (N_860,In_353,In_479);
or U861 (N_861,In_562,In_321);
nor U862 (N_862,In_15,In_668);
and U863 (N_863,In_682,In_371);
nand U864 (N_864,In_578,In_545);
or U865 (N_865,In_375,In_257);
xor U866 (N_866,In_820,In_800);
xnor U867 (N_867,In_635,In_325);
nand U868 (N_868,In_964,In_444);
and U869 (N_869,In_21,In_505);
nand U870 (N_870,In_376,In_880);
or U871 (N_871,In_507,In_286);
or U872 (N_872,In_719,In_376);
nor U873 (N_873,In_251,In_438);
nand U874 (N_874,In_391,In_490);
nor U875 (N_875,In_899,In_373);
and U876 (N_876,In_192,In_403);
or U877 (N_877,In_251,In_817);
or U878 (N_878,In_36,In_337);
and U879 (N_879,In_248,In_331);
or U880 (N_880,In_289,In_953);
nand U881 (N_881,In_343,In_579);
nand U882 (N_882,In_970,In_899);
nand U883 (N_883,In_543,In_738);
nor U884 (N_884,In_90,In_710);
and U885 (N_885,In_451,In_417);
or U886 (N_886,In_885,In_801);
nor U887 (N_887,In_155,In_566);
nand U888 (N_888,In_229,In_168);
nand U889 (N_889,In_532,In_359);
nand U890 (N_890,In_458,In_4);
nand U891 (N_891,In_588,In_93);
nor U892 (N_892,In_311,In_960);
nand U893 (N_893,In_99,In_661);
and U894 (N_894,In_844,In_546);
and U895 (N_895,In_91,In_133);
nand U896 (N_896,In_901,In_943);
nor U897 (N_897,In_303,In_308);
or U898 (N_898,In_860,In_753);
nand U899 (N_899,In_229,In_194);
or U900 (N_900,In_656,In_167);
nor U901 (N_901,In_721,In_425);
nor U902 (N_902,In_85,In_193);
nor U903 (N_903,In_267,In_943);
nand U904 (N_904,In_638,In_482);
or U905 (N_905,In_596,In_783);
and U906 (N_906,In_666,In_928);
nor U907 (N_907,In_948,In_879);
and U908 (N_908,In_893,In_244);
and U909 (N_909,In_604,In_575);
nor U910 (N_910,In_657,In_513);
nor U911 (N_911,In_55,In_464);
and U912 (N_912,In_362,In_728);
nor U913 (N_913,In_119,In_415);
nand U914 (N_914,In_183,In_933);
and U915 (N_915,In_969,In_328);
nor U916 (N_916,In_328,In_635);
and U917 (N_917,In_91,In_20);
xnor U918 (N_918,In_5,In_834);
or U919 (N_919,In_641,In_285);
or U920 (N_920,In_909,In_819);
nand U921 (N_921,In_995,In_514);
nand U922 (N_922,In_964,In_69);
nor U923 (N_923,In_984,In_866);
and U924 (N_924,In_333,In_817);
nand U925 (N_925,In_714,In_342);
nand U926 (N_926,In_8,In_666);
and U927 (N_927,In_164,In_823);
and U928 (N_928,In_601,In_243);
or U929 (N_929,In_743,In_329);
and U930 (N_930,In_966,In_520);
nand U931 (N_931,In_693,In_612);
nand U932 (N_932,In_469,In_379);
or U933 (N_933,In_146,In_897);
and U934 (N_934,In_457,In_14);
nor U935 (N_935,In_580,In_748);
nor U936 (N_936,In_143,In_884);
nand U937 (N_937,In_123,In_926);
nand U938 (N_938,In_254,In_374);
nor U939 (N_939,In_65,In_900);
and U940 (N_940,In_363,In_904);
and U941 (N_941,In_769,In_268);
or U942 (N_942,In_160,In_133);
or U943 (N_943,In_333,In_211);
nor U944 (N_944,In_146,In_122);
xnor U945 (N_945,In_241,In_271);
nor U946 (N_946,In_488,In_238);
and U947 (N_947,In_605,In_808);
nor U948 (N_948,In_451,In_29);
nor U949 (N_949,In_537,In_2);
nor U950 (N_950,In_580,In_482);
nor U951 (N_951,In_788,In_83);
nor U952 (N_952,In_845,In_149);
nor U953 (N_953,In_681,In_900);
nand U954 (N_954,In_699,In_399);
and U955 (N_955,In_809,In_81);
nor U956 (N_956,In_755,In_102);
and U957 (N_957,In_378,In_148);
or U958 (N_958,In_872,In_215);
nor U959 (N_959,In_622,In_968);
and U960 (N_960,In_747,In_620);
nand U961 (N_961,In_167,In_464);
nand U962 (N_962,In_108,In_638);
nand U963 (N_963,In_750,In_547);
or U964 (N_964,In_625,In_610);
or U965 (N_965,In_322,In_261);
nor U966 (N_966,In_517,In_80);
and U967 (N_967,In_52,In_67);
nand U968 (N_968,In_730,In_632);
nand U969 (N_969,In_979,In_764);
nor U970 (N_970,In_7,In_71);
nor U971 (N_971,In_248,In_893);
or U972 (N_972,In_211,In_102);
and U973 (N_973,In_545,In_472);
nand U974 (N_974,In_213,In_198);
xor U975 (N_975,In_577,In_581);
and U976 (N_976,In_301,In_83);
and U977 (N_977,In_37,In_851);
and U978 (N_978,In_702,In_777);
or U979 (N_979,In_925,In_157);
nand U980 (N_980,In_920,In_279);
nor U981 (N_981,In_318,In_817);
or U982 (N_982,In_837,In_115);
nand U983 (N_983,In_257,In_69);
xnor U984 (N_984,In_47,In_890);
or U985 (N_985,In_114,In_598);
nand U986 (N_986,In_174,In_903);
xnor U987 (N_987,In_828,In_623);
or U988 (N_988,In_537,In_162);
and U989 (N_989,In_0,In_451);
nor U990 (N_990,In_338,In_572);
and U991 (N_991,In_690,In_232);
nand U992 (N_992,In_672,In_931);
nand U993 (N_993,In_424,In_583);
or U994 (N_994,In_726,In_716);
nand U995 (N_995,In_305,In_138);
nor U996 (N_996,In_724,In_188);
or U997 (N_997,In_810,In_609);
nor U998 (N_998,In_566,In_296);
nor U999 (N_999,In_173,In_413);
and U1000 (N_1000,In_678,In_592);
nand U1001 (N_1001,In_904,In_319);
or U1002 (N_1002,In_353,In_794);
or U1003 (N_1003,In_285,In_346);
nor U1004 (N_1004,In_1,In_925);
or U1005 (N_1005,In_800,In_749);
or U1006 (N_1006,In_514,In_937);
nor U1007 (N_1007,In_842,In_828);
or U1008 (N_1008,In_688,In_64);
and U1009 (N_1009,In_545,In_65);
and U1010 (N_1010,In_714,In_382);
and U1011 (N_1011,In_865,In_791);
or U1012 (N_1012,In_943,In_89);
nor U1013 (N_1013,In_25,In_147);
nor U1014 (N_1014,In_687,In_197);
and U1015 (N_1015,In_139,In_907);
nand U1016 (N_1016,In_7,In_551);
nand U1017 (N_1017,In_550,In_497);
nor U1018 (N_1018,In_939,In_329);
and U1019 (N_1019,In_628,In_925);
or U1020 (N_1020,In_672,In_471);
and U1021 (N_1021,In_114,In_3);
nor U1022 (N_1022,In_500,In_61);
or U1023 (N_1023,In_964,In_608);
or U1024 (N_1024,In_185,In_606);
or U1025 (N_1025,In_738,In_396);
nand U1026 (N_1026,In_965,In_819);
or U1027 (N_1027,In_58,In_796);
or U1028 (N_1028,In_783,In_700);
nand U1029 (N_1029,In_468,In_296);
nor U1030 (N_1030,In_222,In_292);
or U1031 (N_1031,In_671,In_148);
and U1032 (N_1032,In_837,In_768);
nor U1033 (N_1033,In_860,In_959);
nor U1034 (N_1034,In_167,In_867);
or U1035 (N_1035,In_604,In_858);
or U1036 (N_1036,In_541,In_94);
nand U1037 (N_1037,In_633,In_3);
nand U1038 (N_1038,In_630,In_920);
or U1039 (N_1039,In_555,In_489);
and U1040 (N_1040,In_406,In_652);
and U1041 (N_1041,In_67,In_220);
nor U1042 (N_1042,In_142,In_627);
or U1043 (N_1043,In_739,In_92);
xnor U1044 (N_1044,In_278,In_864);
or U1045 (N_1045,In_154,In_492);
and U1046 (N_1046,In_448,In_246);
or U1047 (N_1047,In_708,In_236);
and U1048 (N_1048,In_195,In_902);
or U1049 (N_1049,In_515,In_535);
nor U1050 (N_1050,In_400,In_146);
nor U1051 (N_1051,In_624,In_266);
and U1052 (N_1052,In_495,In_424);
and U1053 (N_1053,In_536,In_200);
and U1054 (N_1054,In_711,In_263);
nor U1055 (N_1055,In_484,In_446);
nor U1056 (N_1056,In_267,In_386);
and U1057 (N_1057,In_762,In_554);
or U1058 (N_1058,In_176,In_697);
nor U1059 (N_1059,In_423,In_731);
or U1060 (N_1060,In_451,In_532);
and U1061 (N_1061,In_748,In_621);
nor U1062 (N_1062,In_434,In_1);
nand U1063 (N_1063,In_607,In_523);
nor U1064 (N_1064,In_223,In_616);
nand U1065 (N_1065,In_751,In_625);
nand U1066 (N_1066,In_820,In_853);
nor U1067 (N_1067,In_75,In_485);
and U1068 (N_1068,In_649,In_91);
and U1069 (N_1069,In_303,In_577);
nand U1070 (N_1070,In_371,In_205);
and U1071 (N_1071,In_864,In_487);
and U1072 (N_1072,In_986,In_382);
or U1073 (N_1073,In_685,In_632);
nor U1074 (N_1074,In_75,In_309);
and U1075 (N_1075,In_858,In_688);
nor U1076 (N_1076,In_846,In_231);
xnor U1077 (N_1077,In_928,In_767);
and U1078 (N_1078,In_153,In_58);
and U1079 (N_1079,In_308,In_433);
and U1080 (N_1080,In_804,In_29);
nand U1081 (N_1081,In_293,In_179);
nand U1082 (N_1082,In_291,In_559);
and U1083 (N_1083,In_320,In_40);
nor U1084 (N_1084,In_605,In_456);
nor U1085 (N_1085,In_171,In_433);
nand U1086 (N_1086,In_537,In_200);
and U1087 (N_1087,In_274,In_728);
nand U1088 (N_1088,In_707,In_14);
nand U1089 (N_1089,In_938,In_734);
or U1090 (N_1090,In_937,In_505);
or U1091 (N_1091,In_191,In_690);
or U1092 (N_1092,In_360,In_199);
and U1093 (N_1093,In_512,In_191);
or U1094 (N_1094,In_342,In_135);
and U1095 (N_1095,In_439,In_503);
and U1096 (N_1096,In_939,In_77);
and U1097 (N_1097,In_718,In_533);
and U1098 (N_1098,In_147,In_805);
nor U1099 (N_1099,In_75,In_688);
nand U1100 (N_1100,In_96,In_398);
nor U1101 (N_1101,In_877,In_481);
and U1102 (N_1102,In_445,In_422);
nand U1103 (N_1103,In_198,In_706);
and U1104 (N_1104,In_390,In_777);
nand U1105 (N_1105,In_423,In_718);
xor U1106 (N_1106,In_613,In_152);
nor U1107 (N_1107,In_730,In_489);
nor U1108 (N_1108,In_379,In_47);
xor U1109 (N_1109,In_767,In_932);
nand U1110 (N_1110,In_981,In_376);
and U1111 (N_1111,In_248,In_894);
nand U1112 (N_1112,In_678,In_904);
nand U1113 (N_1113,In_927,In_782);
and U1114 (N_1114,In_396,In_389);
nor U1115 (N_1115,In_882,In_939);
and U1116 (N_1116,In_991,In_119);
nor U1117 (N_1117,In_262,In_357);
nand U1118 (N_1118,In_436,In_871);
nor U1119 (N_1119,In_536,In_155);
and U1120 (N_1120,In_13,In_181);
xnor U1121 (N_1121,In_411,In_896);
nor U1122 (N_1122,In_394,In_42);
or U1123 (N_1123,In_992,In_188);
or U1124 (N_1124,In_961,In_432);
xnor U1125 (N_1125,In_340,In_690);
and U1126 (N_1126,In_2,In_368);
nor U1127 (N_1127,In_628,In_137);
or U1128 (N_1128,In_936,In_887);
and U1129 (N_1129,In_249,In_633);
nand U1130 (N_1130,In_221,In_440);
or U1131 (N_1131,In_894,In_775);
and U1132 (N_1132,In_989,In_748);
and U1133 (N_1133,In_640,In_574);
nor U1134 (N_1134,In_358,In_36);
and U1135 (N_1135,In_744,In_837);
and U1136 (N_1136,In_521,In_164);
nand U1137 (N_1137,In_971,In_755);
nor U1138 (N_1138,In_551,In_405);
nor U1139 (N_1139,In_731,In_90);
or U1140 (N_1140,In_842,In_34);
or U1141 (N_1141,In_339,In_954);
nor U1142 (N_1142,In_316,In_866);
and U1143 (N_1143,In_463,In_607);
or U1144 (N_1144,In_545,In_961);
nor U1145 (N_1145,In_335,In_105);
nor U1146 (N_1146,In_797,In_451);
or U1147 (N_1147,In_259,In_466);
nand U1148 (N_1148,In_335,In_344);
xor U1149 (N_1149,In_136,In_971);
xor U1150 (N_1150,In_347,In_64);
nor U1151 (N_1151,In_316,In_726);
and U1152 (N_1152,In_731,In_727);
and U1153 (N_1153,In_770,In_197);
nor U1154 (N_1154,In_178,In_971);
nor U1155 (N_1155,In_313,In_773);
and U1156 (N_1156,In_105,In_641);
and U1157 (N_1157,In_988,In_283);
nand U1158 (N_1158,In_435,In_784);
or U1159 (N_1159,In_345,In_190);
nand U1160 (N_1160,In_297,In_838);
or U1161 (N_1161,In_34,In_899);
nand U1162 (N_1162,In_39,In_765);
xor U1163 (N_1163,In_527,In_649);
and U1164 (N_1164,In_744,In_451);
nor U1165 (N_1165,In_567,In_87);
and U1166 (N_1166,In_430,In_633);
and U1167 (N_1167,In_998,In_592);
nand U1168 (N_1168,In_642,In_94);
nor U1169 (N_1169,In_426,In_405);
or U1170 (N_1170,In_556,In_250);
or U1171 (N_1171,In_495,In_666);
nor U1172 (N_1172,In_508,In_600);
nor U1173 (N_1173,In_168,In_955);
nand U1174 (N_1174,In_633,In_235);
and U1175 (N_1175,In_462,In_400);
or U1176 (N_1176,In_258,In_868);
nor U1177 (N_1177,In_574,In_969);
nor U1178 (N_1178,In_464,In_192);
xnor U1179 (N_1179,In_714,In_92);
nand U1180 (N_1180,In_712,In_200);
and U1181 (N_1181,In_943,In_743);
nor U1182 (N_1182,In_368,In_934);
nand U1183 (N_1183,In_400,In_152);
or U1184 (N_1184,In_388,In_49);
or U1185 (N_1185,In_309,In_259);
and U1186 (N_1186,In_992,In_23);
nor U1187 (N_1187,In_284,In_531);
nand U1188 (N_1188,In_435,In_995);
or U1189 (N_1189,In_21,In_525);
nand U1190 (N_1190,In_996,In_170);
or U1191 (N_1191,In_114,In_320);
or U1192 (N_1192,In_105,In_697);
nand U1193 (N_1193,In_209,In_799);
and U1194 (N_1194,In_43,In_903);
nor U1195 (N_1195,In_169,In_884);
nand U1196 (N_1196,In_494,In_536);
nor U1197 (N_1197,In_355,In_21);
or U1198 (N_1198,In_115,In_890);
and U1199 (N_1199,In_697,In_608);
nand U1200 (N_1200,In_65,In_217);
or U1201 (N_1201,In_382,In_494);
nand U1202 (N_1202,In_773,In_271);
nor U1203 (N_1203,In_840,In_961);
nor U1204 (N_1204,In_522,In_939);
or U1205 (N_1205,In_644,In_997);
or U1206 (N_1206,In_48,In_592);
or U1207 (N_1207,In_770,In_516);
and U1208 (N_1208,In_853,In_838);
nand U1209 (N_1209,In_575,In_856);
or U1210 (N_1210,In_625,In_306);
nor U1211 (N_1211,In_638,In_418);
or U1212 (N_1212,In_147,In_72);
nand U1213 (N_1213,In_100,In_228);
and U1214 (N_1214,In_529,In_75);
nor U1215 (N_1215,In_643,In_37);
nand U1216 (N_1216,In_452,In_0);
nand U1217 (N_1217,In_630,In_672);
and U1218 (N_1218,In_65,In_972);
and U1219 (N_1219,In_885,In_722);
or U1220 (N_1220,In_559,In_593);
nand U1221 (N_1221,In_976,In_122);
nand U1222 (N_1222,In_900,In_15);
nor U1223 (N_1223,In_800,In_977);
and U1224 (N_1224,In_704,In_72);
nand U1225 (N_1225,In_37,In_918);
or U1226 (N_1226,In_922,In_627);
or U1227 (N_1227,In_447,In_260);
nand U1228 (N_1228,In_130,In_337);
nor U1229 (N_1229,In_299,In_714);
nor U1230 (N_1230,In_81,In_192);
or U1231 (N_1231,In_490,In_488);
nor U1232 (N_1232,In_423,In_631);
or U1233 (N_1233,In_898,In_23);
or U1234 (N_1234,In_391,In_703);
nand U1235 (N_1235,In_444,In_248);
xor U1236 (N_1236,In_937,In_899);
nor U1237 (N_1237,In_863,In_989);
or U1238 (N_1238,In_320,In_741);
nor U1239 (N_1239,In_431,In_48);
xnor U1240 (N_1240,In_457,In_649);
or U1241 (N_1241,In_318,In_665);
and U1242 (N_1242,In_960,In_873);
and U1243 (N_1243,In_682,In_784);
nand U1244 (N_1244,In_334,In_847);
or U1245 (N_1245,In_851,In_468);
nor U1246 (N_1246,In_992,In_386);
and U1247 (N_1247,In_740,In_999);
nand U1248 (N_1248,In_819,In_547);
or U1249 (N_1249,In_499,In_581);
nor U1250 (N_1250,In_827,In_606);
nor U1251 (N_1251,In_516,In_835);
nand U1252 (N_1252,In_592,In_948);
nor U1253 (N_1253,In_78,In_803);
and U1254 (N_1254,In_224,In_454);
nor U1255 (N_1255,In_961,In_914);
nand U1256 (N_1256,In_860,In_870);
and U1257 (N_1257,In_338,In_284);
nor U1258 (N_1258,In_760,In_105);
or U1259 (N_1259,In_949,In_23);
and U1260 (N_1260,In_835,In_295);
xnor U1261 (N_1261,In_345,In_783);
nand U1262 (N_1262,In_365,In_74);
xor U1263 (N_1263,In_974,In_405);
and U1264 (N_1264,In_112,In_310);
nor U1265 (N_1265,In_325,In_118);
nand U1266 (N_1266,In_950,In_795);
nand U1267 (N_1267,In_394,In_618);
xor U1268 (N_1268,In_922,In_715);
xnor U1269 (N_1269,In_809,In_592);
or U1270 (N_1270,In_254,In_595);
nor U1271 (N_1271,In_926,In_739);
nor U1272 (N_1272,In_399,In_616);
nor U1273 (N_1273,In_985,In_183);
and U1274 (N_1274,In_162,In_53);
and U1275 (N_1275,In_272,In_284);
and U1276 (N_1276,In_251,In_894);
and U1277 (N_1277,In_72,In_583);
nor U1278 (N_1278,In_899,In_547);
nand U1279 (N_1279,In_497,In_150);
nor U1280 (N_1280,In_844,In_406);
and U1281 (N_1281,In_282,In_805);
and U1282 (N_1282,In_644,In_855);
or U1283 (N_1283,In_401,In_653);
xnor U1284 (N_1284,In_226,In_616);
and U1285 (N_1285,In_703,In_113);
or U1286 (N_1286,In_134,In_110);
nor U1287 (N_1287,In_953,In_637);
nand U1288 (N_1288,In_821,In_64);
and U1289 (N_1289,In_160,In_816);
xnor U1290 (N_1290,In_631,In_278);
and U1291 (N_1291,In_599,In_414);
nor U1292 (N_1292,In_20,In_319);
nor U1293 (N_1293,In_704,In_893);
and U1294 (N_1294,In_761,In_457);
or U1295 (N_1295,In_9,In_370);
nand U1296 (N_1296,In_453,In_593);
or U1297 (N_1297,In_166,In_275);
nand U1298 (N_1298,In_946,In_534);
nand U1299 (N_1299,In_1,In_705);
nand U1300 (N_1300,In_509,In_361);
xor U1301 (N_1301,In_608,In_41);
xor U1302 (N_1302,In_831,In_155);
and U1303 (N_1303,In_39,In_984);
nand U1304 (N_1304,In_104,In_419);
and U1305 (N_1305,In_475,In_708);
and U1306 (N_1306,In_234,In_161);
nor U1307 (N_1307,In_352,In_529);
nor U1308 (N_1308,In_466,In_600);
or U1309 (N_1309,In_359,In_810);
and U1310 (N_1310,In_834,In_591);
nor U1311 (N_1311,In_869,In_28);
and U1312 (N_1312,In_199,In_415);
or U1313 (N_1313,In_305,In_483);
or U1314 (N_1314,In_51,In_818);
or U1315 (N_1315,In_233,In_435);
and U1316 (N_1316,In_659,In_366);
and U1317 (N_1317,In_326,In_174);
nand U1318 (N_1318,In_139,In_511);
or U1319 (N_1319,In_551,In_967);
nand U1320 (N_1320,In_625,In_40);
or U1321 (N_1321,In_581,In_187);
and U1322 (N_1322,In_247,In_635);
nor U1323 (N_1323,In_767,In_103);
xnor U1324 (N_1324,In_795,In_49);
or U1325 (N_1325,In_927,In_540);
nor U1326 (N_1326,In_10,In_285);
nor U1327 (N_1327,In_247,In_385);
nand U1328 (N_1328,In_361,In_638);
and U1329 (N_1329,In_77,In_52);
or U1330 (N_1330,In_578,In_686);
nor U1331 (N_1331,In_512,In_61);
nor U1332 (N_1332,In_96,In_310);
or U1333 (N_1333,In_362,In_723);
or U1334 (N_1334,In_213,In_86);
nand U1335 (N_1335,In_4,In_245);
nor U1336 (N_1336,In_967,In_298);
nand U1337 (N_1337,In_917,In_836);
and U1338 (N_1338,In_164,In_697);
and U1339 (N_1339,In_286,In_451);
nor U1340 (N_1340,In_233,In_141);
and U1341 (N_1341,In_256,In_3);
nand U1342 (N_1342,In_131,In_267);
nor U1343 (N_1343,In_468,In_272);
or U1344 (N_1344,In_408,In_109);
nand U1345 (N_1345,In_63,In_788);
nand U1346 (N_1346,In_341,In_600);
and U1347 (N_1347,In_203,In_249);
and U1348 (N_1348,In_230,In_144);
or U1349 (N_1349,In_312,In_356);
nor U1350 (N_1350,In_465,In_173);
nand U1351 (N_1351,In_350,In_355);
or U1352 (N_1352,In_542,In_491);
or U1353 (N_1353,In_261,In_727);
or U1354 (N_1354,In_630,In_742);
nor U1355 (N_1355,In_339,In_670);
nor U1356 (N_1356,In_404,In_790);
nor U1357 (N_1357,In_865,In_987);
nand U1358 (N_1358,In_543,In_386);
or U1359 (N_1359,In_775,In_193);
xnor U1360 (N_1360,In_515,In_802);
nand U1361 (N_1361,In_926,In_421);
nor U1362 (N_1362,In_766,In_646);
and U1363 (N_1363,In_375,In_659);
or U1364 (N_1364,In_794,In_58);
or U1365 (N_1365,In_426,In_321);
nand U1366 (N_1366,In_702,In_230);
nor U1367 (N_1367,In_957,In_944);
or U1368 (N_1368,In_233,In_774);
nor U1369 (N_1369,In_848,In_546);
nand U1370 (N_1370,In_17,In_881);
and U1371 (N_1371,In_967,In_225);
and U1372 (N_1372,In_546,In_319);
nor U1373 (N_1373,In_640,In_430);
or U1374 (N_1374,In_728,In_14);
and U1375 (N_1375,In_296,In_855);
or U1376 (N_1376,In_945,In_578);
or U1377 (N_1377,In_361,In_572);
xnor U1378 (N_1378,In_569,In_232);
and U1379 (N_1379,In_375,In_468);
or U1380 (N_1380,In_115,In_802);
xor U1381 (N_1381,In_810,In_574);
and U1382 (N_1382,In_665,In_978);
nand U1383 (N_1383,In_783,In_188);
nand U1384 (N_1384,In_736,In_316);
or U1385 (N_1385,In_894,In_818);
nor U1386 (N_1386,In_67,In_648);
nor U1387 (N_1387,In_684,In_289);
nand U1388 (N_1388,In_787,In_992);
or U1389 (N_1389,In_484,In_936);
and U1390 (N_1390,In_640,In_399);
nor U1391 (N_1391,In_185,In_137);
and U1392 (N_1392,In_312,In_201);
and U1393 (N_1393,In_137,In_401);
nor U1394 (N_1394,In_331,In_195);
nand U1395 (N_1395,In_647,In_937);
or U1396 (N_1396,In_707,In_828);
or U1397 (N_1397,In_791,In_256);
and U1398 (N_1398,In_761,In_671);
nor U1399 (N_1399,In_4,In_768);
and U1400 (N_1400,In_308,In_193);
nand U1401 (N_1401,In_978,In_222);
or U1402 (N_1402,In_875,In_953);
and U1403 (N_1403,In_378,In_412);
nor U1404 (N_1404,In_991,In_671);
nand U1405 (N_1405,In_317,In_647);
nand U1406 (N_1406,In_886,In_226);
and U1407 (N_1407,In_972,In_94);
nor U1408 (N_1408,In_643,In_147);
nor U1409 (N_1409,In_870,In_268);
nor U1410 (N_1410,In_643,In_471);
nor U1411 (N_1411,In_156,In_636);
or U1412 (N_1412,In_633,In_375);
or U1413 (N_1413,In_500,In_696);
nand U1414 (N_1414,In_901,In_24);
nand U1415 (N_1415,In_852,In_566);
nand U1416 (N_1416,In_793,In_253);
or U1417 (N_1417,In_118,In_837);
and U1418 (N_1418,In_854,In_813);
nor U1419 (N_1419,In_292,In_343);
and U1420 (N_1420,In_828,In_73);
and U1421 (N_1421,In_426,In_442);
or U1422 (N_1422,In_621,In_208);
or U1423 (N_1423,In_957,In_103);
or U1424 (N_1424,In_20,In_437);
nand U1425 (N_1425,In_445,In_262);
nor U1426 (N_1426,In_577,In_936);
or U1427 (N_1427,In_209,In_420);
and U1428 (N_1428,In_160,In_506);
nand U1429 (N_1429,In_655,In_352);
or U1430 (N_1430,In_374,In_111);
nand U1431 (N_1431,In_803,In_452);
nand U1432 (N_1432,In_779,In_515);
or U1433 (N_1433,In_732,In_713);
nor U1434 (N_1434,In_812,In_426);
nand U1435 (N_1435,In_852,In_681);
nand U1436 (N_1436,In_222,In_153);
and U1437 (N_1437,In_339,In_67);
and U1438 (N_1438,In_925,In_843);
or U1439 (N_1439,In_806,In_309);
or U1440 (N_1440,In_294,In_691);
nor U1441 (N_1441,In_487,In_214);
nand U1442 (N_1442,In_576,In_595);
nor U1443 (N_1443,In_539,In_801);
nor U1444 (N_1444,In_822,In_181);
or U1445 (N_1445,In_449,In_490);
or U1446 (N_1446,In_280,In_861);
or U1447 (N_1447,In_447,In_677);
nand U1448 (N_1448,In_6,In_140);
nand U1449 (N_1449,In_367,In_8);
and U1450 (N_1450,In_295,In_371);
or U1451 (N_1451,In_24,In_253);
or U1452 (N_1452,In_533,In_358);
or U1453 (N_1453,In_469,In_283);
nand U1454 (N_1454,In_282,In_960);
or U1455 (N_1455,In_299,In_909);
nand U1456 (N_1456,In_613,In_651);
or U1457 (N_1457,In_734,In_89);
and U1458 (N_1458,In_159,In_866);
nor U1459 (N_1459,In_122,In_40);
or U1460 (N_1460,In_996,In_990);
nor U1461 (N_1461,In_120,In_642);
and U1462 (N_1462,In_514,In_407);
nor U1463 (N_1463,In_791,In_730);
nand U1464 (N_1464,In_946,In_153);
and U1465 (N_1465,In_859,In_527);
nand U1466 (N_1466,In_88,In_866);
nand U1467 (N_1467,In_212,In_134);
nand U1468 (N_1468,In_150,In_624);
nand U1469 (N_1469,In_718,In_291);
nand U1470 (N_1470,In_184,In_905);
nor U1471 (N_1471,In_790,In_827);
and U1472 (N_1472,In_708,In_648);
nor U1473 (N_1473,In_863,In_621);
and U1474 (N_1474,In_330,In_631);
and U1475 (N_1475,In_330,In_152);
nor U1476 (N_1476,In_475,In_911);
or U1477 (N_1477,In_239,In_790);
or U1478 (N_1478,In_23,In_524);
or U1479 (N_1479,In_722,In_570);
nand U1480 (N_1480,In_734,In_307);
or U1481 (N_1481,In_200,In_291);
nor U1482 (N_1482,In_280,In_62);
and U1483 (N_1483,In_224,In_937);
nand U1484 (N_1484,In_848,In_329);
and U1485 (N_1485,In_410,In_915);
nor U1486 (N_1486,In_416,In_156);
nand U1487 (N_1487,In_669,In_142);
nor U1488 (N_1488,In_418,In_12);
or U1489 (N_1489,In_414,In_358);
and U1490 (N_1490,In_137,In_379);
nor U1491 (N_1491,In_246,In_489);
and U1492 (N_1492,In_448,In_229);
or U1493 (N_1493,In_633,In_528);
nor U1494 (N_1494,In_846,In_81);
and U1495 (N_1495,In_231,In_840);
and U1496 (N_1496,In_689,In_585);
nand U1497 (N_1497,In_181,In_569);
or U1498 (N_1498,In_982,In_636);
and U1499 (N_1499,In_521,In_431);
nand U1500 (N_1500,In_40,In_367);
and U1501 (N_1501,In_444,In_308);
or U1502 (N_1502,In_968,In_447);
nand U1503 (N_1503,In_100,In_33);
or U1504 (N_1504,In_624,In_108);
or U1505 (N_1505,In_341,In_394);
nand U1506 (N_1506,In_558,In_977);
and U1507 (N_1507,In_273,In_581);
nor U1508 (N_1508,In_208,In_424);
nor U1509 (N_1509,In_944,In_597);
nand U1510 (N_1510,In_535,In_238);
nor U1511 (N_1511,In_455,In_37);
nor U1512 (N_1512,In_701,In_400);
nor U1513 (N_1513,In_492,In_62);
nand U1514 (N_1514,In_348,In_595);
nand U1515 (N_1515,In_301,In_615);
or U1516 (N_1516,In_838,In_986);
nand U1517 (N_1517,In_533,In_608);
and U1518 (N_1518,In_580,In_265);
xor U1519 (N_1519,In_121,In_772);
or U1520 (N_1520,In_653,In_166);
or U1521 (N_1521,In_798,In_189);
or U1522 (N_1522,In_781,In_172);
and U1523 (N_1523,In_928,In_533);
nand U1524 (N_1524,In_366,In_278);
nor U1525 (N_1525,In_658,In_792);
and U1526 (N_1526,In_721,In_847);
and U1527 (N_1527,In_318,In_335);
or U1528 (N_1528,In_576,In_972);
or U1529 (N_1529,In_278,In_520);
nand U1530 (N_1530,In_610,In_978);
nand U1531 (N_1531,In_546,In_820);
nand U1532 (N_1532,In_996,In_499);
nand U1533 (N_1533,In_553,In_550);
and U1534 (N_1534,In_100,In_221);
nand U1535 (N_1535,In_455,In_108);
nor U1536 (N_1536,In_13,In_968);
nand U1537 (N_1537,In_927,In_449);
nand U1538 (N_1538,In_694,In_83);
xnor U1539 (N_1539,In_871,In_229);
and U1540 (N_1540,In_500,In_171);
nor U1541 (N_1541,In_571,In_93);
nand U1542 (N_1542,In_180,In_337);
nand U1543 (N_1543,In_48,In_439);
nand U1544 (N_1544,In_547,In_755);
and U1545 (N_1545,In_270,In_762);
nand U1546 (N_1546,In_886,In_126);
nor U1547 (N_1547,In_928,In_63);
nand U1548 (N_1548,In_185,In_747);
nand U1549 (N_1549,In_745,In_420);
and U1550 (N_1550,In_828,In_410);
or U1551 (N_1551,In_659,In_190);
nor U1552 (N_1552,In_960,In_322);
and U1553 (N_1553,In_476,In_723);
or U1554 (N_1554,In_65,In_345);
nand U1555 (N_1555,In_127,In_592);
xnor U1556 (N_1556,In_808,In_862);
and U1557 (N_1557,In_852,In_867);
xnor U1558 (N_1558,In_512,In_142);
nand U1559 (N_1559,In_567,In_712);
or U1560 (N_1560,In_949,In_7);
nand U1561 (N_1561,In_950,In_665);
and U1562 (N_1562,In_754,In_235);
nand U1563 (N_1563,In_725,In_499);
nand U1564 (N_1564,In_970,In_64);
xnor U1565 (N_1565,In_723,In_392);
and U1566 (N_1566,In_923,In_809);
and U1567 (N_1567,In_678,In_207);
nor U1568 (N_1568,In_21,In_864);
and U1569 (N_1569,In_667,In_254);
and U1570 (N_1570,In_219,In_326);
nor U1571 (N_1571,In_581,In_471);
and U1572 (N_1572,In_718,In_799);
nand U1573 (N_1573,In_202,In_55);
nor U1574 (N_1574,In_477,In_764);
or U1575 (N_1575,In_799,In_786);
nor U1576 (N_1576,In_348,In_865);
or U1577 (N_1577,In_356,In_675);
or U1578 (N_1578,In_733,In_741);
or U1579 (N_1579,In_800,In_768);
nand U1580 (N_1580,In_569,In_859);
nor U1581 (N_1581,In_943,In_339);
nor U1582 (N_1582,In_232,In_519);
nand U1583 (N_1583,In_806,In_636);
nor U1584 (N_1584,In_520,In_940);
and U1585 (N_1585,In_532,In_231);
or U1586 (N_1586,In_252,In_211);
or U1587 (N_1587,In_841,In_967);
and U1588 (N_1588,In_206,In_763);
nor U1589 (N_1589,In_244,In_657);
and U1590 (N_1590,In_533,In_786);
and U1591 (N_1591,In_321,In_941);
and U1592 (N_1592,In_501,In_780);
and U1593 (N_1593,In_564,In_594);
nor U1594 (N_1594,In_117,In_280);
nand U1595 (N_1595,In_502,In_945);
or U1596 (N_1596,In_534,In_211);
and U1597 (N_1597,In_392,In_144);
or U1598 (N_1598,In_448,In_406);
and U1599 (N_1599,In_689,In_442);
and U1600 (N_1600,In_504,In_33);
and U1601 (N_1601,In_330,In_687);
and U1602 (N_1602,In_230,In_952);
nand U1603 (N_1603,In_134,In_793);
nor U1604 (N_1604,In_47,In_149);
or U1605 (N_1605,In_214,In_868);
nand U1606 (N_1606,In_207,In_510);
xor U1607 (N_1607,In_230,In_441);
and U1608 (N_1608,In_119,In_758);
nor U1609 (N_1609,In_790,In_839);
nand U1610 (N_1610,In_592,In_614);
or U1611 (N_1611,In_415,In_184);
and U1612 (N_1612,In_989,In_696);
or U1613 (N_1613,In_942,In_746);
nor U1614 (N_1614,In_292,In_383);
nor U1615 (N_1615,In_333,In_629);
nor U1616 (N_1616,In_848,In_888);
nand U1617 (N_1617,In_627,In_508);
or U1618 (N_1618,In_992,In_116);
nand U1619 (N_1619,In_98,In_635);
or U1620 (N_1620,In_798,In_293);
or U1621 (N_1621,In_209,In_86);
nor U1622 (N_1622,In_874,In_765);
and U1623 (N_1623,In_301,In_432);
nand U1624 (N_1624,In_489,In_139);
or U1625 (N_1625,In_118,In_565);
nand U1626 (N_1626,In_398,In_668);
or U1627 (N_1627,In_29,In_785);
or U1628 (N_1628,In_756,In_374);
nor U1629 (N_1629,In_805,In_854);
nand U1630 (N_1630,In_952,In_585);
and U1631 (N_1631,In_641,In_749);
nand U1632 (N_1632,In_193,In_158);
or U1633 (N_1633,In_230,In_844);
and U1634 (N_1634,In_951,In_224);
or U1635 (N_1635,In_968,In_25);
and U1636 (N_1636,In_124,In_664);
or U1637 (N_1637,In_271,In_656);
nor U1638 (N_1638,In_371,In_909);
or U1639 (N_1639,In_50,In_635);
nand U1640 (N_1640,In_783,In_864);
nand U1641 (N_1641,In_220,In_648);
or U1642 (N_1642,In_558,In_891);
and U1643 (N_1643,In_865,In_498);
nand U1644 (N_1644,In_16,In_559);
nor U1645 (N_1645,In_708,In_254);
and U1646 (N_1646,In_53,In_145);
nor U1647 (N_1647,In_647,In_395);
and U1648 (N_1648,In_80,In_709);
nor U1649 (N_1649,In_666,In_515);
or U1650 (N_1650,In_54,In_649);
or U1651 (N_1651,In_908,In_697);
nor U1652 (N_1652,In_156,In_756);
and U1653 (N_1653,In_586,In_979);
or U1654 (N_1654,In_852,In_31);
nand U1655 (N_1655,In_308,In_293);
nor U1656 (N_1656,In_964,In_268);
nor U1657 (N_1657,In_695,In_363);
and U1658 (N_1658,In_368,In_891);
nand U1659 (N_1659,In_356,In_137);
nor U1660 (N_1660,In_135,In_594);
and U1661 (N_1661,In_339,In_726);
nor U1662 (N_1662,In_793,In_233);
nand U1663 (N_1663,In_800,In_911);
and U1664 (N_1664,In_500,In_504);
or U1665 (N_1665,In_487,In_970);
nand U1666 (N_1666,In_950,In_694);
nor U1667 (N_1667,In_104,In_229);
or U1668 (N_1668,In_407,In_451);
or U1669 (N_1669,In_302,In_749);
or U1670 (N_1670,In_333,In_421);
or U1671 (N_1671,In_670,In_295);
nor U1672 (N_1672,In_12,In_495);
and U1673 (N_1673,In_393,In_848);
and U1674 (N_1674,In_405,In_930);
or U1675 (N_1675,In_744,In_310);
and U1676 (N_1676,In_249,In_604);
and U1677 (N_1677,In_540,In_663);
xor U1678 (N_1678,In_894,In_711);
and U1679 (N_1679,In_491,In_717);
nor U1680 (N_1680,In_952,In_299);
or U1681 (N_1681,In_825,In_628);
and U1682 (N_1682,In_854,In_524);
nand U1683 (N_1683,In_482,In_751);
nand U1684 (N_1684,In_34,In_159);
nor U1685 (N_1685,In_298,In_352);
or U1686 (N_1686,In_701,In_594);
nand U1687 (N_1687,In_418,In_604);
nor U1688 (N_1688,In_297,In_841);
and U1689 (N_1689,In_85,In_161);
and U1690 (N_1690,In_306,In_716);
or U1691 (N_1691,In_74,In_761);
xor U1692 (N_1692,In_132,In_810);
or U1693 (N_1693,In_420,In_606);
or U1694 (N_1694,In_19,In_450);
nand U1695 (N_1695,In_816,In_101);
or U1696 (N_1696,In_675,In_521);
or U1697 (N_1697,In_866,In_174);
or U1698 (N_1698,In_924,In_300);
and U1699 (N_1699,In_48,In_441);
nand U1700 (N_1700,In_375,In_883);
nand U1701 (N_1701,In_572,In_950);
nor U1702 (N_1702,In_938,In_858);
or U1703 (N_1703,In_901,In_462);
nand U1704 (N_1704,In_179,In_518);
nor U1705 (N_1705,In_114,In_661);
xnor U1706 (N_1706,In_567,In_974);
and U1707 (N_1707,In_119,In_759);
nand U1708 (N_1708,In_790,In_821);
or U1709 (N_1709,In_180,In_465);
nand U1710 (N_1710,In_62,In_558);
nor U1711 (N_1711,In_524,In_969);
nor U1712 (N_1712,In_485,In_407);
nor U1713 (N_1713,In_361,In_380);
nand U1714 (N_1714,In_699,In_783);
and U1715 (N_1715,In_922,In_365);
and U1716 (N_1716,In_953,In_437);
nand U1717 (N_1717,In_497,In_785);
and U1718 (N_1718,In_992,In_934);
nor U1719 (N_1719,In_669,In_869);
and U1720 (N_1720,In_432,In_355);
nor U1721 (N_1721,In_348,In_539);
nor U1722 (N_1722,In_913,In_230);
and U1723 (N_1723,In_299,In_144);
xor U1724 (N_1724,In_807,In_187);
and U1725 (N_1725,In_953,In_89);
and U1726 (N_1726,In_378,In_29);
nand U1727 (N_1727,In_523,In_477);
nand U1728 (N_1728,In_623,In_720);
or U1729 (N_1729,In_985,In_14);
nand U1730 (N_1730,In_700,In_974);
and U1731 (N_1731,In_649,In_233);
and U1732 (N_1732,In_695,In_159);
and U1733 (N_1733,In_458,In_421);
or U1734 (N_1734,In_379,In_801);
or U1735 (N_1735,In_414,In_278);
or U1736 (N_1736,In_649,In_334);
nor U1737 (N_1737,In_614,In_927);
or U1738 (N_1738,In_423,In_40);
or U1739 (N_1739,In_861,In_57);
or U1740 (N_1740,In_46,In_801);
nor U1741 (N_1741,In_379,In_310);
and U1742 (N_1742,In_100,In_745);
nor U1743 (N_1743,In_659,In_640);
and U1744 (N_1744,In_504,In_710);
xnor U1745 (N_1745,In_633,In_194);
and U1746 (N_1746,In_735,In_529);
and U1747 (N_1747,In_176,In_448);
nand U1748 (N_1748,In_384,In_223);
nor U1749 (N_1749,In_231,In_83);
nor U1750 (N_1750,In_760,In_64);
and U1751 (N_1751,In_100,In_250);
or U1752 (N_1752,In_253,In_16);
or U1753 (N_1753,In_896,In_115);
and U1754 (N_1754,In_5,In_705);
nand U1755 (N_1755,In_710,In_880);
nor U1756 (N_1756,In_393,In_990);
or U1757 (N_1757,In_328,In_41);
and U1758 (N_1758,In_537,In_429);
nand U1759 (N_1759,In_474,In_392);
and U1760 (N_1760,In_203,In_744);
nand U1761 (N_1761,In_513,In_283);
and U1762 (N_1762,In_675,In_133);
nor U1763 (N_1763,In_892,In_435);
and U1764 (N_1764,In_74,In_831);
or U1765 (N_1765,In_884,In_450);
or U1766 (N_1766,In_569,In_989);
and U1767 (N_1767,In_137,In_416);
nand U1768 (N_1768,In_181,In_195);
nand U1769 (N_1769,In_491,In_722);
or U1770 (N_1770,In_876,In_807);
or U1771 (N_1771,In_518,In_31);
and U1772 (N_1772,In_947,In_969);
nand U1773 (N_1773,In_59,In_270);
nor U1774 (N_1774,In_649,In_566);
and U1775 (N_1775,In_620,In_27);
and U1776 (N_1776,In_715,In_333);
nor U1777 (N_1777,In_394,In_933);
nor U1778 (N_1778,In_203,In_45);
and U1779 (N_1779,In_990,In_16);
nand U1780 (N_1780,In_312,In_983);
nand U1781 (N_1781,In_614,In_546);
or U1782 (N_1782,In_523,In_129);
nor U1783 (N_1783,In_753,In_382);
and U1784 (N_1784,In_221,In_38);
nor U1785 (N_1785,In_535,In_836);
xor U1786 (N_1786,In_524,In_718);
and U1787 (N_1787,In_329,In_729);
nor U1788 (N_1788,In_375,In_851);
or U1789 (N_1789,In_467,In_303);
nor U1790 (N_1790,In_807,In_861);
nor U1791 (N_1791,In_278,In_355);
and U1792 (N_1792,In_344,In_173);
or U1793 (N_1793,In_847,In_565);
nor U1794 (N_1794,In_332,In_900);
nor U1795 (N_1795,In_383,In_84);
and U1796 (N_1796,In_746,In_301);
xnor U1797 (N_1797,In_495,In_932);
nor U1798 (N_1798,In_460,In_597);
nand U1799 (N_1799,In_492,In_564);
and U1800 (N_1800,In_516,In_651);
and U1801 (N_1801,In_635,In_923);
or U1802 (N_1802,In_390,In_986);
nor U1803 (N_1803,In_784,In_214);
nor U1804 (N_1804,In_76,In_992);
nand U1805 (N_1805,In_402,In_855);
nand U1806 (N_1806,In_770,In_200);
or U1807 (N_1807,In_510,In_864);
nor U1808 (N_1808,In_310,In_765);
nand U1809 (N_1809,In_479,In_708);
and U1810 (N_1810,In_577,In_381);
and U1811 (N_1811,In_413,In_473);
and U1812 (N_1812,In_144,In_16);
nand U1813 (N_1813,In_861,In_643);
or U1814 (N_1814,In_82,In_420);
nor U1815 (N_1815,In_845,In_541);
or U1816 (N_1816,In_112,In_597);
and U1817 (N_1817,In_897,In_203);
nand U1818 (N_1818,In_867,In_61);
and U1819 (N_1819,In_233,In_719);
nand U1820 (N_1820,In_304,In_364);
xnor U1821 (N_1821,In_607,In_728);
or U1822 (N_1822,In_165,In_432);
nor U1823 (N_1823,In_539,In_738);
nand U1824 (N_1824,In_816,In_730);
nand U1825 (N_1825,In_881,In_261);
nand U1826 (N_1826,In_627,In_772);
nand U1827 (N_1827,In_578,In_592);
or U1828 (N_1828,In_923,In_816);
nand U1829 (N_1829,In_694,In_112);
nor U1830 (N_1830,In_105,In_642);
nand U1831 (N_1831,In_910,In_631);
nand U1832 (N_1832,In_291,In_377);
nor U1833 (N_1833,In_453,In_435);
nand U1834 (N_1834,In_388,In_930);
or U1835 (N_1835,In_779,In_149);
nor U1836 (N_1836,In_82,In_372);
nor U1837 (N_1837,In_102,In_20);
nand U1838 (N_1838,In_999,In_571);
nand U1839 (N_1839,In_27,In_170);
xor U1840 (N_1840,In_486,In_945);
nor U1841 (N_1841,In_823,In_50);
and U1842 (N_1842,In_300,In_325);
or U1843 (N_1843,In_937,In_686);
or U1844 (N_1844,In_805,In_171);
nand U1845 (N_1845,In_668,In_489);
nand U1846 (N_1846,In_751,In_314);
nor U1847 (N_1847,In_87,In_562);
nor U1848 (N_1848,In_693,In_555);
nor U1849 (N_1849,In_410,In_298);
nor U1850 (N_1850,In_552,In_357);
nor U1851 (N_1851,In_133,In_670);
nor U1852 (N_1852,In_446,In_61);
and U1853 (N_1853,In_944,In_381);
nand U1854 (N_1854,In_692,In_322);
and U1855 (N_1855,In_15,In_222);
nand U1856 (N_1856,In_136,In_93);
nand U1857 (N_1857,In_924,In_993);
nor U1858 (N_1858,In_874,In_906);
nor U1859 (N_1859,In_868,In_611);
or U1860 (N_1860,In_728,In_499);
and U1861 (N_1861,In_445,In_692);
or U1862 (N_1862,In_9,In_325);
nand U1863 (N_1863,In_325,In_276);
and U1864 (N_1864,In_755,In_570);
or U1865 (N_1865,In_149,In_761);
and U1866 (N_1866,In_599,In_164);
and U1867 (N_1867,In_641,In_239);
or U1868 (N_1868,In_425,In_467);
nor U1869 (N_1869,In_645,In_4);
nand U1870 (N_1870,In_91,In_359);
nand U1871 (N_1871,In_839,In_58);
nand U1872 (N_1872,In_963,In_651);
nand U1873 (N_1873,In_63,In_764);
nor U1874 (N_1874,In_123,In_923);
and U1875 (N_1875,In_201,In_382);
nor U1876 (N_1876,In_549,In_427);
nor U1877 (N_1877,In_847,In_30);
and U1878 (N_1878,In_800,In_676);
and U1879 (N_1879,In_844,In_67);
and U1880 (N_1880,In_979,In_609);
nor U1881 (N_1881,In_454,In_487);
and U1882 (N_1882,In_113,In_52);
or U1883 (N_1883,In_889,In_377);
nor U1884 (N_1884,In_90,In_944);
nor U1885 (N_1885,In_64,In_751);
nor U1886 (N_1886,In_908,In_141);
nand U1887 (N_1887,In_142,In_138);
nand U1888 (N_1888,In_355,In_949);
nand U1889 (N_1889,In_935,In_717);
or U1890 (N_1890,In_909,In_555);
or U1891 (N_1891,In_595,In_11);
nor U1892 (N_1892,In_880,In_844);
or U1893 (N_1893,In_244,In_927);
and U1894 (N_1894,In_548,In_223);
xor U1895 (N_1895,In_180,In_325);
and U1896 (N_1896,In_979,In_853);
nand U1897 (N_1897,In_217,In_942);
nand U1898 (N_1898,In_734,In_149);
nand U1899 (N_1899,In_961,In_311);
nand U1900 (N_1900,In_167,In_674);
or U1901 (N_1901,In_450,In_468);
nand U1902 (N_1902,In_761,In_469);
and U1903 (N_1903,In_796,In_695);
and U1904 (N_1904,In_12,In_389);
or U1905 (N_1905,In_366,In_480);
and U1906 (N_1906,In_441,In_666);
nand U1907 (N_1907,In_772,In_359);
nand U1908 (N_1908,In_711,In_264);
nand U1909 (N_1909,In_225,In_932);
and U1910 (N_1910,In_295,In_173);
nor U1911 (N_1911,In_485,In_274);
and U1912 (N_1912,In_812,In_702);
or U1913 (N_1913,In_801,In_764);
or U1914 (N_1914,In_267,In_817);
nand U1915 (N_1915,In_702,In_679);
nand U1916 (N_1916,In_984,In_352);
nor U1917 (N_1917,In_832,In_390);
and U1918 (N_1918,In_382,In_514);
nand U1919 (N_1919,In_391,In_939);
and U1920 (N_1920,In_619,In_119);
nand U1921 (N_1921,In_483,In_225);
nor U1922 (N_1922,In_799,In_465);
and U1923 (N_1923,In_105,In_660);
nand U1924 (N_1924,In_871,In_277);
nand U1925 (N_1925,In_585,In_208);
nand U1926 (N_1926,In_57,In_221);
nor U1927 (N_1927,In_393,In_256);
nor U1928 (N_1928,In_974,In_78);
and U1929 (N_1929,In_903,In_241);
nand U1930 (N_1930,In_72,In_454);
and U1931 (N_1931,In_203,In_5);
nand U1932 (N_1932,In_107,In_295);
nor U1933 (N_1933,In_159,In_422);
xnor U1934 (N_1934,In_636,In_796);
nand U1935 (N_1935,In_146,In_796);
nor U1936 (N_1936,In_869,In_691);
or U1937 (N_1937,In_526,In_258);
nand U1938 (N_1938,In_303,In_765);
and U1939 (N_1939,In_144,In_124);
nor U1940 (N_1940,In_67,In_664);
nor U1941 (N_1941,In_813,In_853);
or U1942 (N_1942,In_317,In_826);
and U1943 (N_1943,In_353,In_267);
nor U1944 (N_1944,In_487,In_850);
or U1945 (N_1945,In_840,In_571);
and U1946 (N_1946,In_841,In_565);
nor U1947 (N_1947,In_531,In_696);
nor U1948 (N_1948,In_459,In_276);
nor U1949 (N_1949,In_871,In_449);
and U1950 (N_1950,In_187,In_484);
or U1951 (N_1951,In_777,In_109);
nor U1952 (N_1952,In_571,In_31);
nor U1953 (N_1953,In_853,In_837);
and U1954 (N_1954,In_962,In_571);
nand U1955 (N_1955,In_948,In_52);
or U1956 (N_1956,In_571,In_926);
nor U1957 (N_1957,In_177,In_567);
nor U1958 (N_1958,In_976,In_687);
nor U1959 (N_1959,In_934,In_125);
xor U1960 (N_1960,In_93,In_305);
nor U1961 (N_1961,In_829,In_19);
nor U1962 (N_1962,In_806,In_275);
or U1963 (N_1963,In_948,In_605);
nor U1964 (N_1964,In_618,In_502);
and U1965 (N_1965,In_49,In_895);
or U1966 (N_1966,In_166,In_918);
or U1967 (N_1967,In_756,In_92);
xnor U1968 (N_1968,In_317,In_524);
or U1969 (N_1969,In_509,In_30);
nor U1970 (N_1970,In_971,In_36);
or U1971 (N_1971,In_823,In_53);
and U1972 (N_1972,In_813,In_146);
nor U1973 (N_1973,In_28,In_647);
or U1974 (N_1974,In_508,In_807);
nand U1975 (N_1975,In_664,In_229);
nor U1976 (N_1976,In_782,In_981);
and U1977 (N_1977,In_423,In_220);
nor U1978 (N_1978,In_121,In_949);
nand U1979 (N_1979,In_980,In_65);
and U1980 (N_1980,In_429,In_512);
nand U1981 (N_1981,In_639,In_892);
and U1982 (N_1982,In_74,In_939);
nor U1983 (N_1983,In_11,In_247);
and U1984 (N_1984,In_635,In_702);
or U1985 (N_1985,In_495,In_597);
nand U1986 (N_1986,In_895,In_518);
nor U1987 (N_1987,In_348,In_588);
nand U1988 (N_1988,In_303,In_12);
nand U1989 (N_1989,In_801,In_323);
nand U1990 (N_1990,In_451,In_412);
nand U1991 (N_1991,In_318,In_978);
nor U1992 (N_1992,In_796,In_261);
nor U1993 (N_1993,In_358,In_231);
nor U1994 (N_1994,In_1,In_192);
or U1995 (N_1995,In_254,In_112);
xor U1996 (N_1996,In_71,In_981);
and U1997 (N_1997,In_45,In_56);
or U1998 (N_1998,In_797,In_589);
or U1999 (N_1999,In_930,In_502);
or U2000 (N_2000,In_9,In_17);
nor U2001 (N_2001,In_184,In_821);
and U2002 (N_2002,In_716,In_75);
nor U2003 (N_2003,In_127,In_606);
nor U2004 (N_2004,In_272,In_461);
and U2005 (N_2005,In_215,In_259);
or U2006 (N_2006,In_977,In_614);
or U2007 (N_2007,In_713,In_73);
or U2008 (N_2008,In_569,In_660);
xnor U2009 (N_2009,In_119,In_583);
nor U2010 (N_2010,In_404,In_29);
nor U2011 (N_2011,In_536,In_70);
nand U2012 (N_2012,In_573,In_203);
nand U2013 (N_2013,In_832,In_767);
nor U2014 (N_2014,In_849,In_756);
and U2015 (N_2015,In_491,In_932);
nor U2016 (N_2016,In_270,In_72);
or U2017 (N_2017,In_566,In_966);
nand U2018 (N_2018,In_713,In_538);
and U2019 (N_2019,In_873,In_105);
nand U2020 (N_2020,In_559,In_112);
and U2021 (N_2021,In_850,In_51);
nand U2022 (N_2022,In_200,In_408);
and U2023 (N_2023,In_602,In_329);
and U2024 (N_2024,In_777,In_876);
xnor U2025 (N_2025,In_152,In_147);
nor U2026 (N_2026,In_436,In_329);
nand U2027 (N_2027,In_563,In_142);
nor U2028 (N_2028,In_463,In_945);
and U2029 (N_2029,In_875,In_999);
or U2030 (N_2030,In_803,In_226);
or U2031 (N_2031,In_454,In_835);
and U2032 (N_2032,In_811,In_487);
and U2033 (N_2033,In_663,In_551);
or U2034 (N_2034,In_337,In_431);
and U2035 (N_2035,In_696,In_598);
and U2036 (N_2036,In_66,In_628);
and U2037 (N_2037,In_367,In_37);
nor U2038 (N_2038,In_549,In_749);
and U2039 (N_2039,In_523,In_176);
and U2040 (N_2040,In_944,In_49);
and U2041 (N_2041,In_983,In_1);
nand U2042 (N_2042,In_847,In_623);
and U2043 (N_2043,In_729,In_490);
nor U2044 (N_2044,In_132,In_807);
or U2045 (N_2045,In_839,In_65);
and U2046 (N_2046,In_574,In_178);
or U2047 (N_2047,In_800,In_167);
or U2048 (N_2048,In_988,In_271);
or U2049 (N_2049,In_758,In_105);
or U2050 (N_2050,In_191,In_93);
or U2051 (N_2051,In_776,In_559);
and U2052 (N_2052,In_16,In_591);
nand U2053 (N_2053,In_228,In_36);
nor U2054 (N_2054,In_495,In_601);
nor U2055 (N_2055,In_936,In_721);
or U2056 (N_2056,In_948,In_736);
nor U2057 (N_2057,In_868,In_954);
or U2058 (N_2058,In_949,In_479);
and U2059 (N_2059,In_824,In_693);
and U2060 (N_2060,In_488,In_393);
nand U2061 (N_2061,In_516,In_531);
or U2062 (N_2062,In_85,In_228);
and U2063 (N_2063,In_228,In_655);
nand U2064 (N_2064,In_791,In_280);
or U2065 (N_2065,In_748,In_292);
xor U2066 (N_2066,In_668,In_735);
and U2067 (N_2067,In_667,In_412);
nand U2068 (N_2068,In_925,In_259);
or U2069 (N_2069,In_738,In_112);
xnor U2070 (N_2070,In_601,In_635);
nor U2071 (N_2071,In_983,In_694);
xnor U2072 (N_2072,In_288,In_228);
nand U2073 (N_2073,In_909,In_271);
and U2074 (N_2074,In_413,In_497);
nand U2075 (N_2075,In_291,In_942);
nand U2076 (N_2076,In_836,In_560);
nor U2077 (N_2077,In_209,In_322);
nor U2078 (N_2078,In_238,In_41);
nor U2079 (N_2079,In_330,In_374);
or U2080 (N_2080,In_458,In_558);
and U2081 (N_2081,In_245,In_339);
nand U2082 (N_2082,In_810,In_853);
or U2083 (N_2083,In_485,In_691);
and U2084 (N_2084,In_746,In_529);
or U2085 (N_2085,In_683,In_118);
nor U2086 (N_2086,In_944,In_978);
or U2087 (N_2087,In_83,In_55);
and U2088 (N_2088,In_858,In_401);
nand U2089 (N_2089,In_897,In_340);
nor U2090 (N_2090,In_779,In_422);
and U2091 (N_2091,In_204,In_911);
and U2092 (N_2092,In_37,In_832);
nand U2093 (N_2093,In_330,In_887);
or U2094 (N_2094,In_3,In_158);
nor U2095 (N_2095,In_192,In_444);
nor U2096 (N_2096,In_449,In_866);
and U2097 (N_2097,In_571,In_4);
or U2098 (N_2098,In_109,In_871);
nand U2099 (N_2099,In_467,In_993);
xor U2100 (N_2100,In_102,In_62);
nor U2101 (N_2101,In_144,In_838);
or U2102 (N_2102,In_767,In_60);
nand U2103 (N_2103,In_845,In_788);
nor U2104 (N_2104,In_283,In_885);
xor U2105 (N_2105,In_347,In_105);
or U2106 (N_2106,In_546,In_164);
and U2107 (N_2107,In_609,In_13);
nand U2108 (N_2108,In_99,In_499);
nor U2109 (N_2109,In_122,In_285);
or U2110 (N_2110,In_471,In_787);
xor U2111 (N_2111,In_264,In_249);
or U2112 (N_2112,In_415,In_0);
and U2113 (N_2113,In_529,In_344);
and U2114 (N_2114,In_206,In_711);
nor U2115 (N_2115,In_659,In_628);
or U2116 (N_2116,In_318,In_489);
and U2117 (N_2117,In_451,In_736);
or U2118 (N_2118,In_460,In_159);
and U2119 (N_2119,In_122,In_812);
and U2120 (N_2120,In_781,In_978);
or U2121 (N_2121,In_409,In_268);
nand U2122 (N_2122,In_629,In_16);
nand U2123 (N_2123,In_451,In_678);
and U2124 (N_2124,In_267,In_554);
nand U2125 (N_2125,In_767,In_666);
or U2126 (N_2126,In_847,In_773);
and U2127 (N_2127,In_170,In_763);
nand U2128 (N_2128,In_212,In_991);
and U2129 (N_2129,In_197,In_533);
and U2130 (N_2130,In_539,In_492);
and U2131 (N_2131,In_882,In_677);
nand U2132 (N_2132,In_516,In_854);
or U2133 (N_2133,In_984,In_18);
xnor U2134 (N_2134,In_474,In_993);
and U2135 (N_2135,In_359,In_566);
and U2136 (N_2136,In_52,In_527);
or U2137 (N_2137,In_388,In_979);
nor U2138 (N_2138,In_920,In_13);
nor U2139 (N_2139,In_948,In_865);
and U2140 (N_2140,In_355,In_508);
nor U2141 (N_2141,In_33,In_164);
nor U2142 (N_2142,In_168,In_2);
nand U2143 (N_2143,In_726,In_865);
nor U2144 (N_2144,In_2,In_703);
nor U2145 (N_2145,In_894,In_796);
and U2146 (N_2146,In_241,In_792);
and U2147 (N_2147,In_600,In_184);
or U2148 (N_2148,In_767,In_873);
nor U2149 (N_2149,In_522,In_837);
nor U2150 (N_2150,In_488,In_333);
and U2151 (N_2151,In_872,In_923);
nand U2152 (N_2152,In_320,In_561);
and U2153 (N_2153,In_954,In_753);
nor U2154 (N_2154,In_171,In_990);
and U2155 (N_2155,In_979,In_913);
and U2156 (N_2156,In_809,In_485);
nand U2157 (N_2157,In_428,In_77);
and U2158 (N_2158,In_771,In_75);
nand U2159 (N_2159,In_418,In_477);
and U2160 (N_2160,In_635,In_398);
xor U2161 (N_2161,In_978,In_252);
or U2162 (N_2162,In_303,In_696);
or U2163 (N_2163,In_72,In_376);
nand U2164 (N_2164,In_851,In_496);
nor U2165 (N_2165,In_830,In_493);
and U2166 (N_2166,In_844,In_926);
nor U2167 (N_2167,In_71,In_31);
nand U2168 (N_2168,In_435,In_540);
nand U2169 (N_2169,In_278,In_543);
nor U2170 (N_2170,In_992,In_890);
or U2171 (N_2171,In_240,In_344);
and U2172 (N_2172,In_132,In_187);
and U2173 (N_2173,In_654,In_244);
nor U2174 (N_2174,In_170,In_598);
or U2175 (N_2175,In_850,In_555);
and U2176 (N_2176,In_38,In_358);
nor U2177 (N_2177,In_215,In_66);
nand U2178 (N_2178,In_739,In_828);
nor U2179 (N_2179,In_566,In_680);
or U2180 (N_2180,In_456,In_870);
nor U2181 (N_2181,In_819,In_308);
and U2182 (N_2182,In_76,In_418);
and U2183 (N_2183,In_527,In_29);
or U2184 (N_2184,In_100,In_470);
or U2185 (N_2185,In_46,In_455);
nor U2186 (N_2186,In_493,In_79);
nand U2187 (N_2187,In_493,In_527);
and U2188 (N_2188,In_44,In_968);
or U2189 (N_2189,In_102,In_484);
nand U2190 (N_2190,In_372,In_707);
nor U2191 (N_2191,In_808,In_547);
nand U2192 (N_2192,In_45,In_999);
xnor U2193 (N_2193,In_608,In_335);
and U2194 (N_2194,In_134,In_607);
nor U2195 (N_2195,In_108,In_21);
and U2196 (N_2196,In_145,In_725);
nor U2197 (N_2197,In_675,In_222);
nand U2198 (N_2198,In_318,In_233);
nor U2199 (N_2199,In_969,In_17);
nor U2200 (N_2200,In_294,In_323);
nand U2201 (N_2201,In_698,In_990);
nand U2202 (N_2202,In_720,In_721);
nor U2203 (N_2203,In_885,In_287);
or U2204 (N_2204,In_383,In_888);
and U2205 (N_2205,In_800,In_246);
and U2206 (N_2206,In_587,In_245);
and U2207 (N_2207,In_672,In_814);
nor U2208 (N_2208,In_687,In_416);
and U2209 (N_2209,In_46,In_658);
nor U2210 (N_2210,In_491,In_276);
and U2211 (N_2211,In_594,In_754);
and U2212 (N_2212,In_108,In_204);
nor U2213 (N_2213,In_569,In_383);
nand U2214 (N_2214,In_426,In_792);
or U2215 (N_2215,In_592,In_676);
nand U2216 (N_2216,In_424,In_627);
nor U2217 (N_2217,In_570,In_647);
and U2218 (N_2218,In_384,In_622);
nor U2219 (N_2219,In_404,In_227);
xnor U2220 (N_2220,In_22,In_594);
nand U2221 (N_2221,In_794,In_39);
and U2222 (N_2222,In_162,In_868);
nand U2223 (N_2223,In_348,In_59);
nor U2224 (N_2224,In_399,In_4);
nand U2225 (N_2225,In_777,In_350);
nand U2226 (N_2226,In_891,In_935);
nand U2227 (N_2227,In_973,In_333);
nand U2228 (N_2228,In_279,In_644);
and U2229 (N_2229,In_594,In_632);
or U2230 (N_2230,In_933,In_731);
nor U2231 (N_2231,In_846,In_868);
nand U2232 (N_2232,In_189,In_695);
or U2233 (N_2233,In_387,In_0);
nor U2234 (N_2234,In_282,In_447);
nand U2235 (N_2235,In_802,In_282);
or U2236 (N_2236,In_359,In_394);
and U2237 (N_2237,In_6,In_120);
nor U2238 (N_2238,In_590,In_765);
nand U2239 (N_2239,In_586,In_578);
and U2240 (N_2240,In_551,In_589);
nand U2241 (N_2241,In_487,In_588);
nand U2242 (N_2242,In_642,In_821);
xor U2243 (N_2243,In_695,In_524);
nor U2244 (N_2244,In_770,In_221);
nand U2245 (N_2245,In_123,In_144);
nand U2246 (N_2246,In_882,In_706);
nand U2247 (N_2247,In_66,In_792);
nand U2248 (N_2248,In_639,In_168);
or U2249 (N_2249,In_804,In_904);
nor U2250 (N_2250,In_937,In_888);
nor U2251 (N_2251,In_176,In_558);
nor U2252 (N_2252,In_18,In_837);
and U2253 (N_2253,In_728,In_996);
nand U2254 (N_2254,In_874,In_21);
nand U2255 (N_2255,In_73,In_225);
or U2256 (N_2256,In_181,In_413);
or U2257 (N_2257,In_446,In_714);
or U2258 (N_2258,In_421,In_461);
nor U2259 (N_2259,In_636,In_353);
and U2260 (N_2260,In_219,In_202);
nor U2261 (N_2261,In_315,In_5);
nor U2262 (N_2262,In_46,In_684);
nand U2263 (N_2263,In_467,In_293);
or U2264 (N_2264,In_865,In_953);
nand U2265 (N_2265,In_825,In_250);
nor U2266 (N_2266,In_818,In_459);
and U2267 (N_2267,In_540,In_218);
nor U2268 (N_2268,In_171,In_579);
and U2269 (N_2269,In_708,In_193);
xor U2270 (N_2270,In_264,In_707);
nand U2271 (N_2271,In_523,In_773);
nand U2272 (N_2272,In_83,In_593);
and U2273 (N_2273,In_397,In_742);
or U2274 (N_2274,In_568,In_474);
nand U2275 (N_2275,In_628,In_456);
nand U2276 (N_2276,In_817,In_200);
and U2277 (N_2277,In_789,In_238);
or U2278 (N_2278,In_305,In_319);
and U2279 (N_2279,In_675,In_740);
nor U2280 (N_2280,In_698,In_977);
nor U2281 (N_2281,In_101,In_56);
and U2282 (N_2282,In_715,In_234);
or U2283 (N_2283,In_780,In_509);
nand U2284 (N_2284,In_501,In_493);
nor U2285 (N_2285,In_533,In_693);
or U2286 (N_2286,In_547,In_156);
nand U2287 (N_2287,In_97,In_77);
and U2288 (N_2288,In_722,In_421);
or U2289 (N_2289,In_164,In_359);
nor U2290 (N_2290,In_351,In_167);
xor U2291 (N_2291,In_557,In_342);
nand U2292 (N_2292,In_30,In_716);
nand U2293 (N_2293,In_703,In_553);
nor U2294 (N_2294,In_784,In_719);
or U2295 (N_2295,In_244,In_792);
or U2296 (N_2296,In_305,In_677);
nand U2297 (N_2297,In_175,In_228);
nor U2298 (N_2298,In_520,In_312);
or U2299 (N_2299,In_317,In_660);
and U2300 (N_2300,In_398,In_426);
nor U2301 (N_2301,In_392,In_506);
nor U2302 (N_2302,In_486,In_569);
nor U2303 (N_2303,In_991,In_81);
and U2304 (N_2304,In_955,In_128);
nor U2305 (N_2305,In_440,In_312);
and U2306 (N_2306,In_305,In_705);
nor U2307 (N_2307,In_599,In_511);
nand U2308 (N_2308,In_850,In_382);
nor U2309 (N_2309,In_810,In_199);
nand U2310 (N_2310,In_314,In_668);
or U2311 (N_2311,In_596,In_761);
or U2312 (N_2312,In_843,In_88);
or U2313 (N_2313,In_807,In_337);
nor U2314 (N_2314,In_316,In_759);
or U2315 (N_2315,In_52,In_977);
nand U2316 (N_2316,In_391,In_91);
or U2317 (N_2317,In_533,In_560);
nor U2318 (N_2318,In_550,In_845);
nor U2319 (N_2319,In_514,In_144);
and U2320 (N_2320,In_256,In_823);
nand U2321 (N_2321,In_832,In_203);
or U2322 (N_2322,In_374,In_914);
or U2323 (N_2323,In_344,In_679);
and U2324 (N_2324,In_324,In_57);
or U2325 (N_2325,In_274,In_486);
nor U2326 (N_2326,In_643,In_935);
nor U2327 (N_2327,In_6,In_341);
nor U2328 (N_2328,In_681,In_944);
or U2329 (N_2329,In_323,In_51);
and U2330 (N_2330,In_379,In_368);
or U2331 (N_2331,In_733,In_128);
nor U2332 (N_2332,In_637,In_833);
nor U2333 (N_2333,In_477,In_605);
nand U2334 (N_2334,In_153,In_333);
nor U2335 (N_2335,In_545,In_248);
or U2336 (N_2336,In_739,In_349);
nor U2337 (N_2337,In_261,In_780);
nor U2338 (N_2338,In_290,In_278);
and U2339 (N_2339,In_292,In_642);
nor U2340 (N_2340,In_247,In_5);
or U2341 (N_2341,In_153,In_974);
and U2342 (N_2342,In_660,In_999);
nand U2343 (N_2343,In_382,In_684);
or U2344 (N_2344,In_198,In_11);
nor U2345 (N_2345,In_804,In_365);
nand U2346 (N_2346,In_687,In_699);
nand U2347 (N_2347,In_109,In_258);
nor U2348 (N_2348,In_499,In_927);
nand U2349 (N_2349,In_689,In_407);
and U2350 (N_2350,In_101,In_718);
or U2351 (N_2351,In_905,In_731);
nor U2352 (N_2352,In_842,In_891);
nor U2353 (N_2353,In_148,In_769);
nor U2354 (N_2354,In_131,In_899);
and U2355 (N_2355,In_473,In_277);
or U2356 (N_2356,In_131,In_833);
or U2357 (N_2357,In_406,In_907);
and U2358 (N_2358,In_960,In_102);
nand U2359 (N_2359,In_928,In_173);
or U2360 (N_2360,In_805,In_418);
nand U2361 (N_2361,In_822,In_810);
nor U2362 (N_2362,In_268,In_831);
and U2363 (N_2363,In_897,In_976);
and U2364 (N_2364,In_675,In_766);
nand U2365 (N_2365,In_61,In_909);
nor U2366 (N_2366,In_713,In_895);
and U2367 (N_2367,In_956,In_117);
nand U2368 (N_2368,In_363,In_1);
nor U2369 (N_2369,In_384,In_428);
or U2370 (N_2370,In_751,In_736);
nor U2371 (N_2371,In_501,In_150);
and U2372 (N_2372,In_568,In_524);
nor U2373 (N_2373,In_294,In_384);
and U2374 (N_2374,In_803,In_708);
and U2375 (N_2375,In_532,In_872);
xor U2376 (N_2376,In_399,In_623);
nor U2377 (N_2377,In_669,In_96);
nor U2378 (N_2378,In_822,In_373);
nand U2379 (N_2379,In_938,In_10);
nand U2380 (N_2380,In_188,In_209);
or U2381 (N_2381,In_866,In_343);
nor U2382 (N_2382,In_678,In_47);
and U2383 (N_2383,In_91,In_794);
nand U2384 (N_2384,In_719,In_538);
or U2385 (N_2385,In_894,In_835);
or U2386 (N_2386,In_818,In_766);
and U2387 (N_2387,In_421,In_878);
nand U2388 (N_2388,In_180,In_764);
or U2389 (N_2389,In_466,In_954);
or U2390 (N_2390,In_906,In_203);
and U2391 (N_2391,In_365,In_704);
xor U2392 (N_2392,In_321,In_139);
nand U2393 (N_2393,In_781,In_194);
nor U2394 (N_2394,In_453,In_650);
or U2395 (N_2395,In_265,In_395);
nor U2396 (N_2396,In_103,In_930);
xnor U2397 (N_2397,In_256,In_770);
or U2398 (N_2398,In_604,In_564);
xnor U2399 (N_2399,In_847,In_837);
or U2400 (N_2400,In_859,In_739);
nor U2401 (N_2401,In_38,In_969);
nor U2402 (N_2402,In_396,In_553);
nor U2403 (N_2403,In_678,In_953);
nand U2404 (N_2404,In_310,In_492);
or U2405 (N_2405,In_148,In_108);
nand U2406 (N_2406,In_409,In_476);
or U2407 (N_2407,In_981,In_310);
nand U2408 (N_2408,In_96,In_615);
or U2409 (N_2409,In_637,In_538);
and U2410 (N_2410,In_647,In_994);
or U2411 (N_2411,In_368,In_248);
nor U2412 (N_2412,In_925,In_209);
nand U2413 (N_2413,In_355,In_846);
and U2414 (N_2414,In_684,In_496);
nand U2415 (N_2415,In_809,In_620);
nor U2416 (N_2416,In_138,In_383);
or U2417 (N_2417,In_485,In_144);
nand U2418 (N_2418,In_43,In_527);
and U2419 (N_2419,In_162,In_324);
nor U2420 (N_2420,In_461,In_156);
or U2421 (N_2421,In_386,In_122);
nand U2422 (N_2422,In_637,In_303);
nor U2423 (N_2423,In_16,In_302);
or U2424 (N_2424,In_79,In_52);
nor U2425 (N_2425,In_176,In_859);
nor U2426 (N_2426,In_993,In_910);
nor U2427 (N_2427,In_496,In_64);
or U2428 (N_2428,In_940,In_896);
and U2429 (N_2429,In_889,In_802);
or U2430 (N_2430,In_844,In_10);
nand U2431 (N_2431,In_835,In_618);
nor U2432 (N_2432,In_919,In_344);
nand U2433 (N_2433,In_124,In_892);
nand U2434 (N_2434,In_962,In_4);
or U2435 (N_2435,In_620,In_293);
nor U2436 (N_2436,In_614,In_41);
nor U2437 (N_2437,In_866,In_229);
or U2438 (N_2438,In_362,In_227);
and U2439 (N_2439,In_134,In_653);
or U2440 (N_2440,In_120,In_630);
xnor U2441 (N_2441,In_764,In_309);
or U2442 (N_2442,In_723,In_621);
or U2443 (N_2443,In_136,In_143);
nor U2444 (N_2444,In_757,In_630);
or U2445 (N_2445,In_605,In_968);
and U2446 (N_2446,In_695,In_507);
nand U2447 (N_2447,In_436,In_620);
or U2448 (N_2448,In_580,In_928);
nand U2449 (N_2449,In_720,In_475);
or U2450 (N_2450,In_694,In_992);
nor U2451 (N_2451,In_925,In_487);
nand U2452 (N_2452,In_583,In_408);
or U2453 (N_2453,In_595,In_826);
nor U2454 (N_2454,In_313,In_84);
and U2455 (N_2455,In_958,In_921);
or U2456 (N_2456,In_625,In_635);
nor U2457 (N_2457,In_90,In_803);
nand U2458 (N_2458,In_194,In_978);
nor U2459 (N_2459,In_571,In_753);
and U2460 (N_2460,In_493,In_995);
or U2461 (N_2461,In_69,In_681);
nand U2462 (N_2462,In_848,In_770);
nor U2463 (N_2463,In_78,In_991);
nand U2464 (N_2464,In_464,In_525);
nand U2465 (N_2465,In_648,In_339);
or U2466 (N_2466,In_163,In_360);
nand U2467 (N_2467,In_274,In_41);
and U2468 (N_2468,In_708,In_551);
nand U2469 (N_2469,In_239,In_998);
nand U2470 (N_2470,In_691,In_657);
or U2471 (N_2471,In_938,In_310);
or U2472 (N_2472,In_299,In_41);
nor U2473 (N_2473,In_286,In_565);
nand U2474 (N_2474,In_500,In_268);
and U2475 (N_2475,In_492,In_773);
nand U2476 (N_2476,In_999,In_302);
nor U2477 (N_2477,In_130,In_532);
and U2478 (N_2478,In_902,In_828);
and U2479 (N_2479,In_279,In_523);
and U2480 (N_2480,In_71,In_255);
and U2481 (N_2481,In_432,In_228);
nor U2482 (N_2482,In_926,In_827);
or U2483 (N_2483,In_710,In_429);
nand U2484 (N_2484,In_603,In_666);
or U2485 (N_2485,In_94,In_720);
and U2486 (N_2486,In_602,In_922);
xor U2487 (N_2487,In_212,In_31);
nand U2488 (N_2488,In_769,In_501);
nor U2489 (N_2489,In_424,In_910);
xnor U2490 (N_2490,In_203,In_6);
or U2491 (N_2491,In_428,In_313);
nand U2492 (N_2492,In_465,In_398);
nand U2493 (N_2493,In_874,In_242);
or U2494 (N_2494,In_720,In_152);
and U2495 (N_2495,In_840,In_518);
nor U2496 (N_2496,In_796,In_83);
or U2497 (N_2497,In_759,In_197);
or U2498 (N_2498,In_34,In_182);
nand U2499 (N_2499,In_649,In_310);
or U2500 (N_2500,N_1191,N_2293);
nand U2501 (N_2501,N_211,N_1149);
nand U2502 (N_2502,N_836,N_870);
xnor U2503 (N_2503,N_1095,N_527);
nor U2504 (N_2504,N_1481,N_926);
and U2505 (N_2505,N_472,N_1530);
xnor U2506 (N_2506,N_1336,N_2290);
or U2507 (N_2507,N_646,N_1741);
and U2508 (N_2508,N_980,N_993);
nor U2509 (N_2509,N_754,N_1726);
or U2510 (N_2510,N_25,N_501);
or U2511 (N_2511,N_1935,N_1843);
or U2512 (N_2512,N_453,N_1126);
nor U2513 (N_2513,N_1491,N_1584);
or U2514 (N_2514,N_948,N_908);
or U2515 (N_2515,N_1267,N_1066);
nand U2516 (N_2516,N_264,N_945);
or U2517 (N_2517,N_1916,N_462);
or U2518 (N_2518,N_1179,N_1732);
nand U2519 (N_2519,N_481,N_2103);
or U2520 (N_2520,N_77,N_246);
nor U2521 (N_2521,N_519,N_1711);
nor U2522 (N_2522,N_2335,N_1475);
or U2523 (N_2523,N_1,N_2368);
or U2524 (N_2524,N_379,N_1437);
nand U2525 (N_2525,N_225,N_876);
and U2526 (N_2526,N_1197,N_856);
nor U2527 (N_2527,N_721,N_1998);
nor U2528 (N_2528,N_1470,N_1506);
or U2529 (N_2529,N_2246,N_1482);
nor U2530 (N_2530,N_2468,N_1782);
nor U2531 (N_2531,N_2304,N_404);
nand U2532 (N_2532,N_414,N_855);
nor U2533 (N_2533,N_605,N_405);
nand U2534 (N_2534,N_1487,N_2187);
nand U2535 (N_2535,N_2313,N_1942);
nor U2536 (N_2536,N_1721,N_969);
and U2537 (N_2537,N_1501,N_1708);
or U2538 (N_2538,N_804,N_1462);
nand U2539 (N_2539,N_1838,N_2161);
nand U2540 (N_2540,N_111,N_800);
or U2541 (N_2541,N_2004,N_1093);
nor U2542 (N_2542,N_1166,N_739);
and U2543 (N_2543,N_71,N_1381);
and U2544 (N_2544,N_1019,N_2277);
nor U2545 (N_2545,N_851,N_2491);
or U2546 (N_2546,N_1103,N_2346);
nor U2547 (N_2547,N_2417,N_2244);
or U2548 (N_2548,N_2184,N_1900);
nand U2549 (N_2549,N_2216,N_2116);
nand U2550 (N_2550,N_1348,N_2312);
nor U2551 (N_2551,N_2279,N_1361);
or U2552 (N_2552,N_606,N_640);
nor U2553 (N_2553,N_1633,N_2493);
nor U2554 (N_2554,N_1368,N_2150);
nand U2555 (N_2555,N_2385,N_2220);
or U2556 (N_2556,N_1966,N_1547);
nor U2557 (N_2557,N_1814,N_2331);
nor U2558 (N_2558,N_229,N_554);
nand U2559 (N_2559,N_192,N_1080);
nand U2560 (N_2560,N_869,N_2364);
nand U2561 (N_2561,N_571,N_78);
or U2562 (N_2562,N_1586,N_1785);
and U2563 (N_2563,N_1333,N_2265);
nor U2564 (N_2564,N_23,N_708);
nand U2565 (N_2565,N_1376,N_1196);
nand U2566 (N_2566,N_1923,N_2367);
nand U2567 (N_2567,N_2301,N_2081);
or U2568 (N_2568,N_716,N_538);
or U2569 (N_2569,N_2432,N_1279);
or U2570 (N_2570,N_639,N_844);
and U2571 (N_2571,N_442,N_1284);
and U2572 (N_2572,N_144,N_1129);
or U2573 (N_2573,N_1011,N_1753);
or U2574 (N_2574,N_123,N_1562);
or U2575 (N_2575,N_2118,N_638);
and U2576 (N_2576,N_1985,N_261);
nor U2577 (N_2577,N_43,N_2452);
and U2578 (N_2578,N_916,N_879);
or U2579 (N_2579,N_841,N_320);
nor U2580 (N_2580,N_1884,N_999);
nand U2581 (N_2581,N_1121,N_432);
or U2582 (N_2582,N_2496,N_2238);
and U2583 (N_2583,N_1370,N_408);
nor U2584 (N_2584,N_1097,N_216);
and U2585 (N_2585,N_126,N_893);
nand U2586 (N_2586,N_971,N_1394);
and U2587 (N_2587,N_2155,N_1213);
nor U2588 (N_2588,N_2386,N_203);
nand U2589 (N_2589,N_746,N_1388);
and U2590 (N_2590,N_936,N_2242);
and U2591 (N_2591,N_2267,N_1519);
nand U2592 (N_2592,N_236,N_1846);
or U2593 (N_2593,N_2424,N_2451);
nand U2594 (N_2594,N_2002,N_2429);
or U2595 (N_2595,N_1316,N_1430);
nand U2596 (N_2596,N_915,N_878);
nor U2597 (N_2597,N_441,N_1687);
or U2598 (N_2598,N_1277,N_130);
nor U2599 (N_2599,N_1099,N_748);
or U2600 (N_2600,N_904,N_52);
and U2601 (N_2601,N_1690,N_382);
nand U2602 (N_2602,N_2160,N_476);
nand U2603 (N_2603,N_179,N_169);
nor U2604 (N_2604,N_507,N_1142);
nand U2605 (N_2605,N_2143,N_1391);
nor U2606 (N_2606,N_1762,N_1406);
nor U2607 (N_2607,N_1178,N_989);
and U2608 (N_2608,N_955,N_2024);
nand U2609 (N_2609,N_2445,N_1335);
nand U2610 (N_2610,N_975,N_875);
or U2611 (N_2611,N_486,N_2034);
or U2612 (N_2612,N_1013,N_831);
or U2613 (N_2613,N_1797,N_2145);
xor U2614 (N_2614,N_1398,N_2461);
nor U2615 (N_2615,N_2077,N_1401);
nand U2616 (N_2616,N_331,N_949);
nor U2617 (N_2617,N_124,N_1531);
nand U2618 (N_2618,N_1358,N_257);
and U2619 (N_2619,N_2221,N_987);
and U2620 (N_2620,N_2087,N_1715);
nand U2621 (N_2621,N_1385,N_1044);
nand U2622 (N_2622,N_1311,N_401);
nor U2623 (N_2623,N_188,N_1622);
or U2624 (N_2624,N_1466,N_475);
or U2625 (N_2625,N_2270,N_1453);
and U2626 (N_2626,N_352,N_317);
and U2627 (N_2627,N_1521,N_2498);
xnor U2628 (N_2628,N_725,N_1631);
nor U2629 (N_2629,N_131,N_1342);
or U2630 (N_2630,N_337,N_2106);
nor U2631 (N_2631,N_2140,N_1035);
nand U2632 (N_2632,N_2311,N_2377);
and U2633 (N_2633,N_674,N_296);
or U2634 (N_2634,N_1635,N_397);
nor U2635 (N_2635,N_351,N_350);
and U2636 (N_2636,N_2091,N_894);
or U2637 (N_2637,N_2305,N_2436);
or U2638 (N_2638,N_1655,N_637);
nand U2639 (N_2639,N_1452,N_2254);
or U2640 (N_2640,N_1789,N_504);
xor U2641 (N_2641,N_468,N_1334);
and U2642 (N_2642,N_1374,N_2192);
nor U2643 (N_2643,N_992,N_1702);
nor U2644 (N_2644,N_1249,N_1664);
nor U2645 (N_2645,N_1139,N_371);
nor U2646 (N_2646,N_570,N_2049);
and U2647 (N_2647,N_839,N_1040);
nand U2648 (N_2648,N_711,N_1984);
or U2649 (N_2649,N_1717,N_347);
nand U2650 (N_2650,N_2234,N_1761);
nor U2651 (N_2651,N_60,N_1112);
nand U2652 (N_2652,N_2455,N_2181);
nor U2653 (N_2653,N_114,N_645);
nor U2654 (N_2654,N_1583,N_1891);
or U2655 (N_2655,N_2210,N_1295);
and U2656 (N_2656,N_1600,N_906);
nand U2657 (N_2657,N_817,N_167);
nand U2658 (N_2658,N_631,N_1557);
nor U2659 (N_2659,N_2015,N_1955);
nor U2660 (N_2660,N_49,N_622);
and U2661 (N_2661,N_2344,N_1629);
and U2662 (N_2662,N_1345,N_176);
nand U2663 (N_2663,N_1852,N_724);
nor U2664 (N_2664,N_1668,N_595);
nor U2665 (N_2665,N_872,N_1204);
nor U2666 (N_2666,N_1565,N_2366);
and U2667 (N_2667,N_1329,N_1774);
nor U2668 (N_2668,N_420,N_540);
or U2669 (N_2669,N_2297,N_2402);
and U2670 (N_2670,N_1420,N_1014);
nand U2671 (N_2671,N_151,N_2029);
or U2672 (N_2672,N_1844,N_1173);
nor U2673 (N_2673,N_277,N_559);
or U2674 (N_2674,N_707,N_26);
nor U2675 (N_2675,N_2476,N_1484);
nor U2676 (N_2676,N_944,N_1949);
and U2677 (N_2677,N_1569,N_79);
or U2678 (N_2678,N_1479,N_342);
nand U2679 (N_2679,N_1210,N_1324);
nand U2680 (N_2680,N_510,N_564);
or U2681 (N_2681,N_1777,N_1449);
nor U2682 (N_2682,N_2176,N_1587);
nand U2683 (N_2683,N_1034,N_127);
or U2684 (N_2684,N_2412,N_1575);
and U2685 (N_2685,N_1938,N_2391);
and U2686 (N_2686,N_200,N_436);
nand U2687 (N_2687,N_2153,N_888);
or U2688 (N_2688,N_2361,N_1218);
nand U2689 (N_2689,N_853,N_1418);
and U2690 (N_2690,N_51,N_2052);
nand U2691 (N_2691,N_2051,N_2308);
or U2692 (N_2692,N_2164,N_780);
or U2693 (N_2693,N_1544,N_2115);
nor U2694 (N_2694,N_1554,N_979);
and U2695 (N_2695,N_2405,N_1555);
or U2696 (N_2696,N_961,N_332);
and U2697 (N_2697,N_1070,N_2253);
nor U2698 (N_2698,N_513,N_1498);
nand U2699 (N_2699,N_1386,N_1275);
nand U2700 (N_2700,N_1076,N_1661);
or U2701 (N_2701,N_1198,N_2310);
or U2702 (N_2702,N_1104,N_1281);
nand U2703 (N_2703,N_905,N_59);
nor U2704 (N_2704,N_2442,N_349);
or U2705 (N_2705,N_2411,N_649);
and U2706 (N_2706,N_621,N_2454);
and U2707 (N_2707,N_1893,N_819);
nand U2708 (N_2708,N_2355,N_618);
nor U2709 (N_2709,N_1956,N_2247);
nand U2710 (N_2710,N_1445,N_2146);
nand U2711 (N_2711,N_2166,N_221);
or U2712 (N_2712,N_943,N_32);
or U2713 (N_2713,N_690,N_1051);
and U2714 (N_2714,N_435,N_165);
nor U2715 (N_2715,N_1793,N_1004);
nand U2716 (N_2716,N_1958,N_1351);
and U2717 (N_2717,N_2497,N_1349);
and U2718 (N_2718,N_2157,N_2440);
nand U2719 (N_2719,N_2348,N_2014);
xnor U2720 (N_2720,N_1323,N_2151);
and U2721 (N_2721,N_2190,N_1647);
and U2722 (N_2722,N_1674,N_2264);
nor U2723 (N_2723,N_458,N_1839);
nand U2724 (N_2724,N_895,N_2203);
nand U2725 (N_2725,N_2175,N_1500);
nand U2726 (N_2726,N_1207,N_561);
or U2727 (N_2727,N_97,N_22);
nand U2728 (N_2728,N_2207,N_1536);
nand U2729 (N_2729,N_898,N_1003);
and U2730 (N_2730,N_1122,N_642);
or U2731 (N_2731,N_365,N_280);
or U2732 (N_2732,N_2185,N_1795);
or U2733 (N_2733,N_709,N_1199);
nor U2734 (N_2734,N_1634,N_1450);
or U2735 (N_2735,N_1170,N_1654);
nand U2736 (N_2736,N_2033,N_1410);
nor U2737 (N_2737,N_2063,N_41);
and U2738 (N_2738,N_344,N_2101);
or U2739 (N_2739,N_1048,N_2482);
and U2740 (N_2740,N_951,N_1181);
and U2741 (N_2741,N_2378,N_1176);
xor U2742 (N_2742,N_2397,N_1653);
nor U2743 (N_2743,N_187,N_1948);
nor U2744 (N_2744,N_1613,N_191);
nand U2745 (N_2745,N_492,N_399);
and U2746 (N_2746,N_148,N_89);
nand U2747 (N_2747,N_1068,N_737);
xnor U2748 (N_2748,N_530,N_1508);
nor U2749 (N_2749,N_1623,N_548);
and U2750 (N_2750,N_1941,N_2459);
nand U2751 (N_2751,N_129,N_553);
or U2752 (N_2752,N_1303,N_620);
nand U2753 (N_2753,N_784,N_1988);
nand U2754 (N_2754,N_1085,N_2307);
and U2755 (N_2755,N_2382,N_1957);
nand U2756 (N_2756,N_2082,N_962);
nand U2757 (N_2757,N_1617,N_2007);
nand U2758 (N_2758,N_226,N_2055);
nand U2759 (N_2759,N_2258,N_1389);
or U2760 (N_2760,N_306,N_512);
nand U2761 (N_2761,N_1180,N_198);
nand U2762 (N_2762,N_985,N_1274);
nor U2763 (N_2763,N_103,N_1880);
and U2764 (N_2764,N_2068,N_372);
nand U2765 (N_2765,N_137,N_1823);
and U2766 (N_2766,N_2433,N_574);
and U2767 (N_2767,N_2375,N_1953);
or U2768 (N_2768,N_275,N_1723);
or U2769 (N_2769,N_139,N_2136);
nand U2770 (N_2770,N_24,N_1174);
nor U2771 (N_2771,N_966,N_1913);
nand U2772 (N_2772,N_1766,N_1148);
or U2773 (N_2773,N_40,N_1026);
nor U2774 (N_2774,N_155,N_1287);
or U2775 (N_2775,N_2449,N_1863);
and U2776 (N_2776,N_838,N_2197);
or U2777 (N_2777,N_847,N_2434);
or U2778 (N_2778,N_482,N_1892);
nor U2779 (N_2779,N_1610,N_568);
nor U2780 (N_2780,N_1413,N_28);
nor U2781 (N_2781,N_164,N_431);
nand U2782 (N_2782,N_1440,N_301);
nand U2783 (N_2783,N_1270,N_2100);
xor U2784 (N_2784,N_2095,N_1379);
xor U2785 (N_2785,N_582,N_417);
or U2786 (N_2786,N_1424,N_499);
nor U2787 (N_2787,N_1509,N_1087);
and U2788 (N_2788,N_2439,N_974);
and U2789 (N_2789,N_1781,N_1384);
or U2790 (N_2790,N_670,N_1786);
nor U2791 (N_2791,N_2096,N_1593);
and U2792 (N_2792,N_1169,N_2248);
nand U2793 (N_2793,N_1714,N_508);
and U2794 (N_2794,N_429,N_822);
nand U2795 (N_2795,N_956,N_1006);
and U2796 (N_2796,N_616,N_312);
nand U2797 (N_2797,N_1110,N_1772);
or U2798 (N_2798,N_2406,N_1644);
or U2799 (N_2799,N_1096,N_1881);
or U2800 (N_2800,N_1867,N_1527);
nand U2801 (N_2801,N_30,N_632);
and U2802 (N_2802,N_1225,N_2255);
and U2803 (N_2803,N_2225,N_1124);
xnor U2804 (N_2804,N_1262,N_141);
and U2805 (N_2805,N_195,N_558);
nand U2806 (N_2806,N_892,N_995);
or U2807 (N_2807,N_929,N_850);
nor U2808 (N_2808,N_2065,N_2032);
and U2809 (N_2809,N_2174,N_1858);
nand U2810 (N_2810,N_1339,N_656);
and U2811 (N_2811,N_2127,N_336);
nor U2812 (N_2812,N_650,N_415);
and U2813 (N_2813,N_2462,N_653);
or U2814 (N_2814,N_1513,N_1670);
and U2815 (N_2815,N_938,N_13);
and U2816 (N_2816,N_1659,N_2485);
nand U2817 (N_2817,N_896,N_837);
or U2818 (N_2818,N_981,N_1614);
and U2819 (N_2819,N_1626,N_807);
or U2820 (N_2820,N_1257,N_821);
nand U2821 (N_2821,N_1423,N_1594);
nand U2822 (N_2822,N_1483,N_1220);
nor U2823 (N_2823,N_396,N_2430);
nand U2824 (N_2824,N_2189,N_666);
nand U2825 (N_2825,N_427,N_890);
and U2826 (N_2826,N_1175,N_2040);
and U2827 (N_2827,N_1268,N_292);
nand U2828 (N_2828,N_1697,N_1234);
nor U2829 (N_2829,N_1754,N_88);
or U2830 (N_2830,N_752,N_627);
or U2831 (N_2831,N_166,N_1028);
or U2832 (N_2832,N_80,N_223);
nor U2833 (N_2833,N_2026,N_1252);
nand U2834 (N_2834,N_2338,N_1673);
or U2835 (N_2835,N_914,N_500);
nand U2836 (N_2836,N_318,N_1549);
and U2837 (N_2837,N_1514,N_1739);
nor U2838 (N_2838,N_823,N_232);
nor U2839 (N_2839,N_2021,N_2414);
nand U2840 (N_2840,N_735,N_923);
nand U2841 (N_2841,N_687,N_580);
or U2842 (N_2842,N_1172,N_2171);
nor U2843 (N_2843,N_1157,N_1609);
nand U2844 (N_2844,N_727,N_72);
or U2845 (N_2845,N_487,N_2419);
or U2846 (N_2846,N_366,N_451);
nand U2847 (N_2847,N_1933,N_8);
and U2848 (N_2848,N_2232,N_1105);
or U2849 (N_2849,N_815,N_498);
nand U2850 (N_2850,N_1522,N_830);
and U2851 (N_2851,N_2269,N_1618);
nor U2852 (N_2852,N_2019,N_920);
nor U2853 (N_2853,N_2109,N_1184);
and U2854 (N_2854,N_1108,N_1399);
and U2855 (N_2855,N_2113,N_147);
nand U2856 (N_2856,N_294,N_394);
or U2857 (N_2857,N_1253,N_1827);
xor U2858 (N_2858,N_1457,N_329);
nor U2859 (N_2859,N_609,N_270);
nor U2860 (N_2860,N_887,N_145);
or U2861 (N_2861,N_658,N_134);
nand U2862 (N_2862,N_353,N_18);
and U2863 (N_2863,N_1133,N_1412);
nor U2864 (N_2864,N_2369,N_1993);
and U2865 (N_2865,N_219,N_788);
or U2866 (N_2866,N_884,N_1826);
or U2867 (N_2867,N_313,N_2401);
and U2868 (N_2868,N_1309,N_589);
or U2869 (N_2869,N_133,N_753);
xnor U2870 (N_2870,N_2239,N_2050);
nand U2871 (N_2871,N_1371,N_1350);
and U2872 (N_2872,N_1053,N_2130);
nor U2873 (N_2873,N_16,N_506);
or U2874 (N_2874,N_1845,N_1959);
or U2875 (N_2875,N_994,N_541);
nor U2876 (N_2876,N_1232,N_1638);
nor U2877 (N_2877,N_174,N_864);
nand U2878 (N_2878,N_803,N_1704);
nand U2879 (N_2879,N_1650,N_719);
and U2880 (N_2880,N_1043,N_2104);
nor U2881 (N_2881,N_551,N_2283);
nand U2882 (N_2882,N_1305,N_566);
nand U2883 (N_2883,N_2172,N_1778);
and U2884 (N_2884,N_1662,N_437);
nand U2885 (N_2885,N_1224,N_1947);
and U2886 (N_2886,N_2320,N_1929);
and U2887 (N_2887,N_2167,N_1152);
or U2888 (N_2888,N_555,N_1190);
or U2889 (N_2889,N_1493,N_1119);
nor U2890 (N_2890,N_170,N_732);
and U2891 (N_2891,N_1203,N_39);
nor U2892 (N_2892,N_1925,N_2235);
nor U2893 (N_2893,N_2045,N_45);
nor U2894 (N_2894,N_1005,N_1735);
and U2895 (N_2895,N_1510,N_1700);
or U2896 (N_2896,N_1109,N_231);
xnor U2897 (N_2897,N_1943,N_1293);
nand U2898 (N_2898,N_2183,N_65);
nand U2899 (N_2899,N_720,N_1327);
and U2900 (N_2900,N_871,N_1646);
nand U2901 (N_2901,N_931,N_9);
nand U2902 (N_2902,N_2403,N_284);
nor U2903 (N_2903,N_1658,N_1405);
nand U2904 (N_2904,N_2022,N_2404);
and U2905 (N_2905,N_1136,N_263);
nand U2906 (N_2906,N_479,N_1969);
nand U2907 (N_2907,N_1002,N_1469);
nand U2908 (N_2908,N_2273,N_1579);
or U2909 (N_2909,N_612,N_952);
xor U2910 (N_2910,N_2198,N_1691);
and U2911 (N_2911,N_505,N_1448);
and U2912 (N_2912,N_2230,N_918);
and U2913 (N_2913,N_186,N_965);
or U2914 (N_2914,N_300,N_789);
nor U2915 (N_2915,N_2374,N_1288);
nor U2916 (N_2916,N_1128,N_1961);
nor U2917 (N_2917,N_1822,N_1314);
or U2918 (N_2918,N_2111,N_1815);
and U2919 (N_2919,N_2178,N_1595);
or U2920 (N_2920,N_552,N_36);
or U2921 (N_2921,N_64,N_113);
nor U2922 (N_2922,N_2046,N_101);
and U2923 (N_2923,N_1436,N_825);
and U2924 (N_2924,N_325,N_1564);
nor U2925 (N_2925,N_214,N_1041);
or U2926 (N_2926,N_522,N_1317);
nand U2927 (N_2927,N_689,N_1903);
nor U2928 (N_2928,N_1459,N_2473);
or U2929 (N_2929,N_2078,N_2205);
and U2930 (N_2930,N_1032,N_1601);
nand U2931 (N_2931,N_1116,N_1425);
nand U2932 (N_2932,N_1576,N_1752);
nand U2933 (N_2933,N_48,N_1542);
or U2934 (N_2934,N_2010,N_1141);
nand U2935 (N_2935,N_2149,N_1417);
nand U2936 (N_2936,N_2036,N_1018);
or U2937 (N_2937,N_1981,N_1832);
and U2938 (N_2938,N_597,N_793);
or U2939 (N_2939,N_86,N_867);
nor U2940 (N_2940,N_1625,N_440);
or U2941 (N_2941,N_12,N_227);
or U2942 (N_2942,N_1012,N_303);
nand U2943 (N_2943,N_322,N_272);
nand U2944 (N_2944,N_1382,N_1532);
nand U2945 (N_2945,N_369,N_673);
and U2946 (N_2946,N_805,N_824);
or U2947 (N_2947,N_1719,N_484);
nand U2948 (N_2948,N_1446,N_594);
xor U2949 (N_2949,N_2098,N_1695);
xor U2950 (N_2950,N_2437,N_210);
nor U2951 (N_2951,N_2300,N_340);
nand U2952 (N_2952,N_1915,N_854);
or U2953 (N_2953,N_565,N_2325);
and U2954 (N_2954,N_346,N_1950);
nand U2955 (N_2955,N_692,N_465);
nor U2956 (N_2956,N_2243,N_1496);
nor U2957 (N_2957,N_2259,N_321);
or U2958 (N_2958,N_2001,N_2306);
or U2959 (N_2959,N_902,N_1680);
nor U2960 (N_2960,N_1049,N_1090);
and U2961 (N_2961,N_668,N_1086);
and U2962 (N_2962,N_880,N_2107);
or U2963 (N_2963,N_1098,N_1320);
and U2964 (N_2964,N_1123,N_1447);
nand U2965 (N_2965,N_536,N_87);
nand U2966 (N_2966,N_521,N_1499);
nand U2967 (N_2967,N_228,N_4);
nor U2968 (N_2968,N_1686,N_1058);
nand U2969 (N_2969,N_407,N_2363);
nand U2970 (N_2970,N_1015,N_626);
nand U2971 (N_2971,N_1486,N_46);
and U2972 (N_2972,N_808,N_2241);
or U2973 (N_2973,N_783,N_91);
or U2974 (N_2974,N_2324,N_1485);
nand U2975 (N_2975,N_1296,N_157);
and U2976 (N_2976,N_2373,N_269);
or U2977 (N_2977,N_293,N_1763);
and U2978 (N_2978,N_1050,N_2315);
or U2979 (N_2979,N_1936,N_2356);
nor U2980 (N_2980,N_1990,N_792);
and U2981 (N_2981,N_135,N_276);
nand U2982 (N_2982,N_260,N_2477);
and U2983 (N_2983,N_1675,N_683);
and U2984 (N_2984,N_411,N_652);
nand U2985 (N_2985,N_775,N_1082);
and U2986 (N_2986,N_2370,N_463);
and U2987 (N_2987,N_1241,N_617);
nor U2988 (N_2988,N_2121,N_1147);
nor U2989 (N_2989,N_1372,N_1895);
and U2990 (N_2990,N_2226,N_5);
nand U2991 (N_2991,N_1980,N_921);
or U2992 (N_2992,N_390,N_2392);
or U2993 (N_2993,N_1724,N_1404);
nand U2994 (N_2994,N_573,N_1454);
nand U2995 (N_2995,N_218,N_577);
and U2996 (N_2996,N_1716,N_1037);
and U2997 (N_2997,N_206,N_2105);
nor U2998 (N_2998,N_866,N_490);
and U2999 (N_2999,N_54,N_425);
or U3000 (N_3000,N_1831,N_745);
and U3001 (N_3001,N_1983,N_2008);
and U3002 (N_3002,N_2389,N_1533);
nand U3003 (N_3003,N_654,N_1703);
nor U3004 (N_3004,N_874,N_302);
nor U3005 (N_3005,N_1052,N_897);
nor U3006 (N_3006,N_1811,N_782);
nand U3007 (N_3007,N_2499,N_1813);
and U3008 (N_3008,N_781,N_2148);
nand U3009 (N_3009,N_509,N_1725);
or U3010 (N_3010,N_278,N_664);
or U3011 (N_3011,N_799,N_1922);
nand U3012 (N_3012,N_1432,N_1373);
or U3013 (N_3013,N_1874,N_2137);
nand U3014 (N_3014,N_2289,N_354);
or U3015 (N_3015,N_2018,N_1408);
or U3016 (N_3016,N_833,N_1009);
or U3017 (N_3017,N_1889,N_1063);
nand U3018 (N_3018,N_1236,N_403);
nand U3019 (N_3019,N_1878,N_1291);
or U3020 (N_3020,N_592,N_751);
or U3021 (N_3021,N_970,N_2464);
nand U3022 (N_3022,N_1573,N_1836);
or U3023 (N_3023,N_2492,N_0);
and U3024 (N_3024,N_1528,N_1393);
or U3025 (N_3025,N_445,N_1285);
and U3026 (N_3026,N_168,N_723);
nor U3027 (N_3027,N_1411,N_1830);
nor U3028 (N_3028,N_1474,N_1226);
nor U3029 (N_3029,N_583,N_2354);
nand U3030 (N_3030,N_604,N_758);
nand U3031 (N_3031,N_265,N_1255);
and U3032 (N_3032,N_1952,N_1857);
or U3033 (N_3033,N_1855,N_1606);
nor U3034 (N_3034,N_873,N_2394);
and U3035 (N_3035,N_2071,N_1696);
and U3036 (N_3036,N_1768,N_556);
nor U3037 (N_3037,N_1489,N_1362);
nand U3038 (N_3038,N_1894,N_2457);
nand U3039 (N_3039,N_1850,N_816);
or U3040 (N_3040,N_245,N_1566);
and U3041 (N_3041,N_1115,N_282);
and U3042 (N_3042,N_1201,N_1960);
nor U3043 (N_3043,N_591,N_1540);
and U3044 (N_3044,N_2222,N_271);
or U3045 (N_3045,N_2169,N_1997);
nand U3046 (N_3046,N_2060,N_2112);
or U3047 (N_3047,N_903,N_1870);
nor U3048 (N_3048,N_2206,N_1365);
or U3049 (N_3049,N_518,N_2211);
nand U3050 (N_3050,N_1887,N_477);
or U3051 (N_3051,N_1918,N_706);
nand U3052 (N_3052,N_900,N_1643);
and U3053 (N_3053,N_1776,N_2275);
nand U3054 (N_3054,N_2067,N_1666);
nor U3055 (N_3055,N_2302,N_1572);
and U3056 (N_3056,N_2467,N_734);
or U3057 (N_3057,N_705,N_927);
or U3058 (N_3058,N_2215,N_419);
and U3059 (N_3059,N_2003,N_2028);
or U3060 (N_3060,N_1699,N_2163);
nand U3061 (N_3061,N_2005,N_1962);
or U3062 (N_3062,N_972,N_1208);
and U3063 (N_3063,N_1869,N_1709);
nand U3064 (N_3064,N_728,N_1861);
or U3065 (N_3065,N_1828,N_940);
and U3066 (N_3066,N_2341,N_2035);
nor U3067 (N_3067,N_1042,N_934);
or U3068 (N_3068,N_2410,N_2418);
or U3069 (N_3069,N_2069,N_2177);
or U3070 (N_3070,N_1206,N_798);
nor U3071 (N_3071,N_557,N_563);
and U3072 (N_3072,N_1344,N_1548);
nor U3073 (N_3073,N_67,N_307);
nor U3074 (N_3074,N_1182,N_1899);
and U3075 (N_3075,N_1987,N_2345);
and U3076 (N_3076,N_1227,N_1140);
nand U3077 (N_3077,N_1229,N_285);
nor U3078 (N_3078,N_1520,N_2245);
nor U3079 (N_3079,N_496,N_1387);
nand U3080 (N_3080,N_1627,N_598);
nand U3081 (N_3081,N_889,N_1074);
or U3082 (N_3082,N_2428,N_2075);
and U3083 (N_3083,N_2483,N_1392);
nand U3084 (N_3084,N_2044,N_603);
and U3085 (N_3085,N_763,N_964);
or U3086 (N_3086,N_1931,N_69);
and U3087 (N_3087,N_1965,N_1266);
nand U3088 (N_3088,N_109,N_533);
and U3089 (N_3089,N_1017,N_1456);
and U3090 (N_3090,N_702,N_1286);
and U3091 (N_3091,N_1677,N_572);
nand U3092 (N_3092,N_1167,N_1737);
and U3093 (N_3093,N_1230,N_1775);
and U3094 (N_3094,N_1100,N_588);
nor U3095 (N_3095,N_254,N_1054);
and U3096 (N_3096,N_1265,N_644);
nor U3097 (N_3097,N_651,N_355);
or U3098 (N_3098,N_585,N_607);
nor U3099 (N_3099,N_1146,N_37);
or U3100 (N_3100,N_450,N_1473);
and U3101 (N_3101,N_102,N_1636);
and U3102 (N_3102,N_785,N_1438);
or U3103 (N_3103,N_1089,N_930);
or U3104 (N_3104,N_99,N_835);
or U3105 (N_3105,N_1264,N_2233);
or U3106 (N_3106,N_1750,N_599);
nor U3107 (N_3107,N_1835,N_1442);
nand U3108 (N_3108,N_398,N_545);
and U3109 (N_3109,N_478,N_2123);
and U3110 (N_3110,N_801,N_459);
nand U3111 (N_3111,N_2413,N_2453);
nor U3112 (N_3112,N_1490,N_1964);
or U3113 (N_3113,N_811,N_2085);
or U3114 (N_3114,N_1022,N_988);
and U3115 (N_3115,N_1395,N_1021);
and U3116 (N_3116,N_986,N_375);
and U3117 (N_3117,N_1865,N_1061);
and U3118 (N_3118,N_1541,N_576);
and U3119 (N_3119,N_1992,N_2062);
and U3120 (N_3120,N_524,N_881);
or U3121 (N_3121,N_70,N_1607);
or U3122 (N_3122,N_1143,N_1810);
and U3123 (N_3123,N_843,N_611);
and U3124 (N_3124,N_146,N_330);
or U3125 (N_3125,N_2227,N_2124);
or U3126 (N_3126,N_1944,N_502);
or U3127 (N_3127,N_1630,N_1346);
or U3128 (N_3128,N_1193,N_740);
nor U3129 (N_3129,N_1151,N_1701);
nor U3130 (N_3130,N_1332,N_2090);
and U3131 (N_3131,N_996,N_1117);
nor U3132 (N_3132,N_773,N_2132);
and U3133 (N_3133,N_55,N_249);
nor U3134 (N_3134,N_204,N_1312);
and U3135 (N_3135,N_2296,N_2427);
or U3136 (N_3136,N_1315,N_2083);
and U3137 (N_3137,N_1665,N_2463);
or U3138 (N_3138,N_466,N_1582);
nor U3139 (N_3139,N_1046,N_2281);
and U3140 (N_3140,N_2446,N_712);
nor U3141 (N_3141,N_984,N_777);
nand U3142 (N_3142,N_1559,N_2490);
or U3143 (N_3143,N_2379,N_2387);
and U3144 (N_3144,N_2357,N_1792);
and U3145 (N_3145,N_1188,N_1212);
nand U3146 (N_3146,N_2388,N_1879);
and U3147 (N_3147,N_2135,N_255);
or U3148 (N_3148,N_1840,N_861);
nor U3149 (N_3149,N_143,N_62);
nor U3150 (N_3150,N_659,N_1897);
nand U3151 (N_3151,N_623,N_295);
nor U3152 (N_3152,N_1738,N_932);
or U3153 (N_3153,N_6,N_2390);
xnor U3154 (N_3154,N_1860,N_175);
nor U3155 (N_3155,N_1127,N_1621);
xnor U3156 (N_3156,N_309,N_1694);
or U3157 (N_3157,N_266,N_2224);
nor U3158 (N_3158,N_2299,N_2475);
and U3159 (N_3159,N_2489,N_1886);
and U3160 (N_3160,N_1808,N_1278);
or U3161 (N_3161,N_660,N_217);
nand U3162 (N_3162,N_1301,N_1186);
nand U3163 (N_3163,N_1672,N_430);
or U3164 (N_3164,N_1896,N_1106);
and U3165 (N_3165,N_1337,N_1803);
and U3166 (N_3166,N_2017,N_2126);
nand U3167 (N_3167,N_154,N_208);
and U3168 (N_3168,N_315,N_2231);
nor U3169 (N_3169,N_1556,N_662);
or U3170 (N_3170,N_1156,N_2195);
nor U3171 (N_3171,N_2426,N_2381);
and U3172 (N_3172,N_1906,N_1568);
and U3173 (N_3173,N_1194,N_1771);
nand U3174 (N_3174,N_2336,N_2086);
and U3175 (N_3175,N_584,N_928);
nor U3176 (N_3176,N_2383,N_770);
or U3177 (N_3177,N_1325,N_1036);
or U3178 (N_3178,N_1338,N_1546);
or U3179 (N_3179,N_1722,N_587);
nor U3180 (N_3180,N_1968,N_2059);
or U3181 (N_3181,N_2494,N_1000);
or U3182 (N_3182,N_2237,N_682);
and U3183 (N_3183,N_376,N_1260);
nor U3184 (N_3184,N_1409,N_1589);
or U3185 (N_3185,N_1901,N_1047);
and U3186 (N_3186,N_1231,N_1125);
and U3187 (N_3187,N_1801,N_201);
and U3188 (N_3188,N_238,N_1632);
nor U3189 (N_3189,N_388,N_1693);
or U3190 (N_3190,N_361,N_511);
nand U3191 (N_3191,N_2142,N_911);
nor U3192 (N_3192,N_1414,N_1824);
or U3193 (N_3193,N_967,N_1578);
nand U3194 (N_3194,N_485,N_2333);
or U3195 (N_3195,N_1937,N_1250);
nor U3196 (N_3196,N_2252,N_532);
nand U3197 (N_3197,N_2080,N_447);
or U3198 (N_3198,N_1535,N_1476);
or U3199 (N_3199,N_909,N_1107);
or U3200 (N_3200,N_1258,N_2097);
nor U3201 (N_3201,N_1328,N_234);
nand U3202 (N_3202,N_1366,N_2425);
or U3203 (N_3203,N_1882,N_326);
and U3204 (N_3204,N_2000,N_2420);
or U3205 (N_3205,N_1507,N_1580);
nand U3206 (N_3206,N_1403,N_1161);
nand U3207 (N_3207,N_550,N_546);
nand U3208 (N_3208,N_1341,N_11);
and U3209 (N_3209,N_1728,N_2251);
nor U3210 (N_3210,N_444,N_657);
nand U3211 (N_3211,N_31,N_1145);
nand U3212 (N_3212,N_387,N_209);
and U3213 (N_3213,N_1624,N_1353);
nand U3214 (N_3214,N_1800,N_212);
xor U3215 (N_3215,N_2326,N_776);
nor U3216 (N_3216,N_865,N_2196);
nand U3217 (N_3217,N_413,N_1088);
and U3218 (N_3218,N_2360,N_2292);
nand U3219 (N_3219,N_153,N_963);
nand U3220 (N_3220,N_790,N_806);
or U3221 (N_3221,N_2456,N_672);
and U3222 (N_3222,N_691,N_562);
nand U3223 (N_3223,N_1598,N_207);
nand U3224 (N_3224,N_942,N_1272);
nor U3225 (N_3225,N_1560,N_389);
and U3226 (N_3226,N_858,N_1492);
nor U3227 (N_3227,N_291,N_2173);
nand U3228 (N_3228,N_818,N_2322);
nor U3229 (N_3229,N_1729,N_973);
and U3230 (N_3230,N_1787,N_1439);
and U3231 (N_3231,N_237,N_177);
nor U3232 (N_3232,N_1604,N_1134);
nor U3233 (N_3233,N_1856,N_2236);
nand U3234 (N_3234,N_1946,N_182);
or U3235 (N_3235,N_122,N_2191);
nand U3236 (N_3236,N_181,N_2288);
or U3237 (N_3237,N_222,N_1467);
and U3238 (N_3238,N_1751,N_1713);
nand U3239 (N_3239,N_968,N_602);
nand U3240 (N_3240,N_239,N_2212);
and U3241 (N_3241,N_575,N_287);
nand U3242 (N_3242,N_1978,N_601);
and U3243 (N_3243,N_1619,N_1657);
nor U3244 (N_3244,N_324,N_2158);
nand U3245 (N_3245,N_56,N_663);
or U3246 (N_3246,N_852,N_1577);
xnor U3247 (N_3247,N_1921,N_1628);
nand U3248 (N_3248,N_925,N_515);
or U3249 (N_3249,N_1712,N_1177);
or U3250 (N_3250,N_197,N_1912);
or U3251 (N_3251,N_240,N_1300);
nor U3252 (N_3252,N_750,N_220);
and U3253 (N_3253,N_717,N_1760);
xnor U3254 (N_3254,N_2278,N_1319);
or U3255 (N_3255,N_681,N_2208);
nor U3256 (N_3256,N_1038,N_1571);
and U3257 (N_3257,N_1558,N_648);
and U3258 (N_3258,N_701,N_901);
or U3259 (N_3259,N_1282,N_2327);
or U3260 (N_3260,N_1790,N_1154);
nor U3261 (N_3261,N_2488,N_743);
or U3262 (N_3262,N_1421,N_1433);
nand U3263 (N_3263,N_802,N_250);
nand U3264 (N_3264,N_730,N_1645);
and U3265 (N_3265,N_2084,N_224);
and U3266 (N_3266,N_733,N_1130);
or U3267 (N_3267,N_1471,N_460);
nand U3268 (N_3268,N_2240,N_402);
nand U3269 (N_3269,N_686,N_2061);
or U3270 (N_3270,N_1242,N_2162);
nand U3271 (N_3271,N_1783,N_832);
or U3272 (N_3272,N_1131,N_862);
xor U3273 (N_3273,N_1648,N_2250);
and U3274 (N_3274,N_159,N_1849);
nor U3275 (N_3275,N_1364,N_813);
nand U3276 (N_3276,N_2487,N_3);
nor U3277 (N_3277,N_163,N_1596);
and U3278 (N_3278,N_1045,N_578);
or U3279 (N_3279,N_17,N_1667);
or U3280 (N_3280,N_1426,N_304);
xor U3281 (N_3281,N_107,N_1534);
and U3282 (N_3282,N_1503,N_1299);
nand U3283 (N_3283,N_1165,N_1698);
and U3284 (N_3284,N_1383,N_1187);
nand U3285 (N_3285,N_1357,N_1254);
nor U3286 (N_3286,N_883,N_34);
and U3287 (N_3287,N_1238,N_171);
and U3288 (N_3288,N_2053,N_308);
and U3289 (N_3289,N_196,N_1989);
nor U3290 (N_3290,N_2263,N_2125);
nand U3291 (N_3291,N_715,N_1010);
nand U3292 (N_3292,N_1681,N_1217);
and U3293 (N_3293,N_456,N_1359);
nor U3294 (N_3294,N_1773,N_2444);
nand U3295 (N_3295,N_1330,N_58);
or U3296 (N_3296,N_1720,N_1158);
nand U3297 (N_3297,N_1495,N_2303);
nand U3298 (N_3298,N_1977,N_1240);
nor U3299 (N_3299,N_2094,N_494);
and U3300 (N_3300,N_1380,N_299);
nand U3301 (N_3301,N_755,N_83);
nand U3302 (N_3302,N_138,N_2108);
or U3303 (N_3303,N_2321,N_1072);
nor U3304 (N_3304,N_319,N_434);
or U3305 (N_3305,N_1574,N_443);
or U3306 (N_3306,N_2340,N_2159);
or U3307 (N_3307,N_2041,N_1064);
or U3308 (N_3308,N_1331,N_671);
and U3309 (N_3309,N_2470,N_235);
nand U3310 (N_3310,N_1039,N_1821);
nor U3311 (N_3311,N_796,N_1927);
nand U3312 (N_3312,N_1612,N_1727);
or U3313 (N_3313,N_455,N_762);
or U3314 (N_3314,N_2266,N_2330);
nor U3315 (N_3315,N_1367,N_549);
and U3316 (N_3316,N_1740,N_1755);
nor U3317 (N_3317,N_1745,N_1932);
and U3318 (N_3318,N_1620,N_410);
and U3319 (N_3319,N_1637,N_1669);
nand U3320 (N_3320,N_1642,N_428);
and U3321 (N_3321,N_392,N_108);
and U3322 (N_3322,N_112,N_439);
or U3323 (N_3323,N_991,N_1245);
and U3324 (N_3324,N_1736,N_917);
nand U3325 (N_3325,N_713,N_744);
nor U3326 (N_3326,N_2030,N_1991);
nor U3327 (N_3327,N_613,N_1407);
nand U3328 (N_3328,N_1511,N_860);
xnor U3329 (N_3329,N_998,N_1347);
nor U3330 (N_3330,N_886,N_1660);
and U3331 (N_3331,N_2012,N_1866);
and U3332 (N_3332,N_421,N_1926);
or U3333 (N_3333,N_2229,N_2179);
nor U3334 (N_3334,N_121,N_2287);
and U3335 (N_3335,N_205,N_119);
nand U3336 (N_3336,N_543,N_173);
xnor U3337 (N_3337,N_1917,N_2393);
and U3338 (N_3338,N_826,N_1458);
nor U3339 (N_3339,N_378,N_1705);
nor U3340 (N_3340,N_787,N_2438);
or U3341 (N_3341,N_2037,N_2043);
nor U3342 (N_3342,N_1605,N_63);
or U3343 (N_3343,N_2272,N_281);
and U3344 (N_3344,N_82,N_1444);
nor U3345 (N_3345,N_1999,N_452);
nand U3346 (N_3346,N_1590,N_1427);
nor U3347 (N_3347,N_2249,N_96);
nand U3348 (N_3348,N_1302,N_1524);
nor U3349 (N_3349,N_1016,N_1798);
and U3350 (N_3350,N_2219,N_2039);
nor U3351 (N_3351,N_1819,N_73);
and U3352 (N_3352,N_1092,N_2152);
or U3353 (N_3353,N_809,N_2134);
and U3354 (N_3354,N_395,N_2416);
or U3355 (N_3355,N_1872,N_105);
nor U3356 (N_3356,N_1817,N_747);
or U3357 (N_3357,N_1537,N_2102);
nor U3358 (N_3358,N_467,N_1237);
nor U3359 (N_3359,N_1435,N_1055);
nand U3360 (N_3360,N_1794,N_547);
nor U3361 (N_3361,N_2217,N_2271);
xnor U3362 (N_3362,N_820,N_503);
nor U3363 (N_3363,N_1497,N_643);
and U3364 (N_3364,N_1280,N_1062);
or U3365 (N_3365,N_1974,N_92);
nand U3366 (N_3366,N_1463,N_1431);
nand U3367 (N_3367,N_400,N_1940);
nand U3368 (N_3368,N_1402,N_2339);
nand U3369 (N_3369,N_368,N_514);
nor U3370 (N_3370,N_367,N_1355);
or U3371 (N_3371,N_1976,N_471);
nand U3372 (N_3372,N_1543,N_1748);
nand U3373 (N_3373,N_1159,N_1354);
nor U3374 (N_3374,N_2372,N_1885);
nor U3375 (N_3375,N_696,N_1764);
nor U3376 (N_3376,N_2193,N_2286);
and U3377 (N_3377,N_935,N_1215);
and U3378 (N_3378,N_677,N_426);
or U3379 (N_3379,N_377,N_859);
and U3380 (N_3380,N_464,N_156);
nor U3381 (N_3381,N_1829,N_116);
nand U3382 (N_3382,N_2458,N_190);
nor U3383 (N_3383,N_233,N_2280);
and U3384 (N_3384,N_526,N_1567);
or U3385 (N_3385,N_1788,N_1890);
nor U3386 (N_3386,N_2114,N_766);
and U3387 (N_3387,N_1078,N_1185);
nor U3388 (N_3388,N_669,N_150);
and U3389 (N_3389,N_1599,N_741);
and U3390 (N_3390,N_2365,N_95);
nand U3391 (N_3391,N_774,N_2353);
nor U3392 (N_3392,N_1029,N_947);
nand U3393 (N_3393,N_1907,N_978);
nor U3394 (N_3394,N_53,N_1970);
nor U3395 (N_3395,N_323,N_383);
nor U3396 (N_3396,N_2423,N_1995);
and U3397 (N_3397,N_2396,N_528);
nand U3398 (N_3398,N_1102,N_2110);
xor U3399 (N_3399,N_2099,N_422);
nand U3400 (N_3400,N_615,N_409);
and U3401 (N_3401,N_1477,N_1294);
or U3402 (N_3402,N_910,N_757);
or U3403 (N_3403,N_1689,N_812);
nand U3404 (N_3404,N_2268,N_1276);
or U3405 (N_3405,N_2479,N_172);
nor U3406 (N_3406,N_534,N_1375);
nor U3407 (N_3407,N_2156,N_1603);
nand U3408 (N_3408,N_132,N_1075);
or U3409 (N_3409,N_1876,N_1008);
nor U3410 (N_3410,N_1244,N_128);
and U3411 (N_3411,N_1963,N_311);
nand U3412 (N_3412,N_1707,N_2466);
and U3413 (N_3413,N_1919,N_1552);
nor U3414 (N_3414,N_1292,N_117);
and U3415 (N_3415,N_629,N_765);
nand U3416 (N_3416,N_2469,N_959);
nand U3417 (N_3417,N_1135,N_1488);
nand U3418 (N_3418,N_1585,N_178);
nand U3419 (N_3419,N_1263,N_193);
or U3420 (N_3420,N_756,N_1928);
nor U3421 (N_3421,N_958,N_2228);
nand U3422 (N_3422,N_1834,N_2474);
or U3423 (N_3423,N_579,N_1113);
nor U3424 (N_3424,N_1975,N_289);
nor U3425 (N_3425,N_1663,N_1924);
nand U3426 (N_3426,N_2415,N_1526);
nor U3427 (N_3427,N_953,N_1416);
or U3428 (N_3428,N_1195,N_125);
nor U3429 (N_3429,N_243,N_1163);
xor U3430 (N_3430,N_779,N_2337);
or U3431 (N_3431,N_2057,N_2371);
nor U3432 (N_3432,N_2362,N_21);
xor U3433 (N_3433,N_1219,N_829);
nor U3434 (N_3434,N_230,N_675);
and U3435 (N_3435,N_1945,N_842);
nor U3436 (N_3436,N_2460,N_726);
or U3437 (N_3437,N_449,N_525);
nand U3438 (N_3438,N_1796,N_423);
nor U3439 (N_3439,N_1352,N_1001);
nand U3440 (N_3440,N_1057,N_385);
or U3441 (N_3441,N_685,N_194);
and U3442 (N_3442,N_2076,N_241);
or U3443 (N_3443,N_2073,N_339);
or U3444 (N_3444,N_2400,N_1862);
or U3445 (N_3445,N_1377,N_1025);
nand U3446 (N_3446,N_1251,N_1326);
and U3447 (N_3447,N_2256,N_678);
nor U3448 (N_3448,N_539,N_635);
nor U3449 (N_3449,N_2352,N_1898);
nand U3450 (N_3450,N_1920,N_1007);
nand U3451 (N_3451,N_983,N_2329);
nand U3452 (N_3452,N_1640,N_2223);
and U3453 (N_3453,N_247,N_535);
or U3454 (N_3454,N_1073,N_710);
or U3455 (N_3455,N_1307,N_74);
or U3456 (N_3456,N_1067,N_1805);
and U3457 (N_3457,N_1847,N_882);
nor U3458 (N_3458,N_749,N_359);
nand U3459 (N_3459,N_1806,N_778);
and U3460 (N_3460,N_316,N_863);
nand U3461 (N_3461,N_273,N_2380);
nand U3462 (N_3462,N_1758,N_2117);
or U3463 (N_3463,N_76,N_2282);
nand U3464 (N_3464,N_1480,N_2328);
nand U3465 (N_3465,N_1939,N_364);
and U3466 (N_3466,N_891,N_268);
nor U3467 (N_3467,N_1415,N_795);
nand U3468 (N_3468,N_66,N_1419);
and U3469 (N_3469,N_1441,N_2465);
and U3470 (N_3470,N_2154,N_2284);
nand U3471 (N_3471,N_960,N_1202);
nand U3472 (N_3472,N_19,N_693);
and U3473 (N_3473,N_2170,N_1749);
nor U3474 (N_3474,N_1360,N_655);
and U3475 (N_3475,N_2421,N_845);
nand U3476 (N_3476,N_1779,N_457);
or U3477 (N_3477,N_199,N_1155);
nor U3478 (N_3478,N_1400,N_256);
and U3479 (N_3479,N_2486,N_937);
or U3480 (N_3480,N_94,N_1211);
nand U3481 (N_3481,N_1322,N_1243);
nor U3482 (N_3482,N_267,N_544);
nand U3483 (N_3483,N_767,N_2180);
or U3484 (N_3484,N_2129,N_258);
nand U3485 (N_3485,N_1027,N_81);
nor U3486 (N_3486,N_338,N_694);
nor U3487 (N_3487,N_1460,N_1468);
and U3488 (N_3488,N_2260,N_2079);
nor U3489 (N_3489,N_497,N_461);
xnor U3490 (N_3490,N_2186,N_2011);
and U3491 (N_3491,N_149,N_2194);
and U3492 (N_3492,N_2471,N_1273);
nor U3493 (N_3493,N_373,N_2218);
and U3494 (N_3494,N_1545,N_1734);
xnor U3495 (N_3495,N_567,N_1505);
nor U3496 (N_3496,N_480,N_1651);
or U3497 (N_3497,N_1318,N_160);
nor U3498 (N_3498,N_61,N_684);
or U3499 (N_3499,N_161,N_424);
or U3500 (N_3500,N_2314,N_520);
nor U3501 (N_3501,N_416,N_2274);
and U3502 (N_3502,N_1461,N_1083);
and U3503 (N_3503,N_1369,N_2316);
and U3504 (N_3504,N_2350,N_1615);
or U3505 (N_3505,N_697,N_1221);
and U3506 (N_3506,N_244,N_1081);
nor U3507 (N_3507,N_769,N_68);
and U3508 (N_3508,N_184,N_2495);
or U3509 (N_3509,N_2332,N_1304);
nor U3510 (N_3510,N_1422,N_215);
nor U3511 (N_3511,N_1616,N_1770);
nand U3512 (N_3512,N_1023,N_2480);
and U3513 (N_3513,N_2351,N_380);
nor U3514 (N_3514,N_310,N_877);
nand U3515 (N_3515,N_474,N_1222);
nor U3516 (N_3516,N_1464,N_2319);
and U3517 (N_3517,N_42,N_1859);
nor U3518 (N_3518,N_1837,N_2);
nor U3519 (N_3519,N_115,N_625);
nor U3520 (N_3520,N_1563,N_680);
nand U3521 (N_3521,N_699,N_1588);
or U3522 (N_3522,N_140,N_665);
or U3523 (N_3523,N_771,N_2200);
nor U3524 (N_3524,N_760,N_977);
nor U3525 (N_3525,N_27,N_1079);
nand U3526 (N_3526,N_764,N_2025);
nand U3527 (N_3527,N_1930,N_957);
and U3528 (N_3528,N_47,N_1118);
nor U3529 (N_3529,N_1812,N_1854);
nor U3530 (N_3530,N_1570,N_1216);
nor U3531 (N_3531,N_531,N_849);
or U3532 (N_3532,N_406,N_954);
or U3533 (N_3533,N_183,N_15);
or U3534 (N_3534,N_1247,N_57);
or U3535 (N_3535,N_1030,N_493);
or U3536 (N_3536,N_2435,N_1767);
xor U3537 (N_3537,N_1683,N_814);
and U3538 (N_3538,N_262,N_297);
or U3539 (N_3539,N_2144,N_44);
or U3540 (N_3540,N_990,N_834);
or U3541 (N_3541,N_1747,N_1971);
nor U3542 (N_3542,N_1162,N_1256);
nor U3543 (N_3543,N_2334,N_158);
nor U3544 (N_3544,N_2214,N_688);
xor U3545 (N_3545,N_700,N_152);
and U3546 (N_3546,N_667,N_90);
nand U3547 (N_3547,N_1523,N_469);
or U3548 (N_3548,N_1784,N_35);
or U3549 (N_3549,N_2199,N_1451);
or U3550 (N_3550,N_1306,N_1671);
xor U3551 (N_3551,N_950,N_253);
nand U3552 (N_3552,N_704,N_1429);
nand U3553 (N_3553,N_641,N_1111);
and U3554 (N_3554,N_2399,N_248);
nor U3555 (N_3555,N_1059,N_1780);
and U3556 (N_3556,N_85,N_695);
nand U3557 (N_3557,N_1682,N_110);
xor U3558 (N_3558,N_722,N_2138);
nand U3559 (N_3559,N_1235,N_630);
and U3560 (N_3560,N_314,N_1094);
nor U3561 (N_3561,N_33,N_848);
or U3562 (N_3562,N_251,N_1652);
or U3563 (N_3563,N_679,N_1223);
or U3564 (N_3564,N_772,N_1730);
and U3565 (N_3565,N_2070,N_2042);
nor U3566 (N_3566,N_391,N_1551);
nor U3567 (N_3567,N_924,N_470);
xnor U3568 (N_3568,N_1340,N_2088);
nor U3569 (N_3569,N_1472,N_1804);
and U3570 (N_3570,N_1871,N_100);
xor U3571 (N_3571,N_647,N_1200);
nand U3572 (N_3572,N_1688,N_729);
nand U3573 (N_3573,N_768,N_1308);
or U3574 (N_3574,N_1060,N_10);
or U3575 (N_3575,N_596,N_1825);
or U3576 (N_3576,N_327,N_529);
nand U3577 (N_3577,N_1908,N_333);
or U3578 (N_3578,N_2295,N_1071);
and U3579 (N_3579,N_142,N_2168);
and U3580 (N_3580,N_2072,N_614);
and U3581 (N_3581,N_857,N_1743);
and U3582 (N_3582,N_433,N_1914);
nand U3583 (N_3583,N_328,N_1649);
nand U3584 (N_3584,N_1816,N_1077);
and U3585 (N_3585,N_2408,N_1259);
nand U3586 (N_3586,N_698,N_106);
nor U3587 (N_3587,N_1592,N_2202);
and U3588 (N_3588,N_274,N_933);
nand U3589 (N_3589,N_370,N_634);
or U3590 (N_3590,N_1525,N_2347);
xnor U3591 (N_3591,N_1742,N_1904);
nor U3592 (N_3592,N_1909,N_1676);
or U3593 (N_3593,N_454,N_1132);
or U3594 (N_3594,N_2147,N_1967);
nand U3595 (N_3595,N_288,N_305);
nor U3596 (N_3596,N_1757,N_120);
nor U3597 (N_3597,N_2213,N_1343);
nand U3598 (N_3598,N_1137,N_919);
nor U3599 (N_3599,N_2359,N_1678);
nand U3600 (N_3600,N_356,N_412);
nor U3601 (N_3601,N_1171,N_2298);
or U3602 (N_3602,N_242,N_2323);
nor U3603 (N_3603,N_386,N_982);
nor U3604 (N_3604,N_2201,N_1972);
nand U3605 (N_3605,N_1321,N_384);
nand U3606 (N_3606,N_676,N_1710);
or U3607 (N_3607,N_2047,N_1160);
nor U3608 (N_3608,N_345,N_593);
nand U3609 (N_3609,N_885,N_1759);
nand U3610 (N_3610,N_718,N_868);
nand U3611 (N_3611,N_1138,N_1214);
xor U3612 (N_3612,N_1982,N_1791);
nand U3613 (N_3613,N_517,N_489);
nand U3614 (N_3614,N_1853,N_1396);
and U3615 (N_3615,N_1397,N_446);
nor U3616 (N_3616,N_1611,N_38);
nand U3617 (N_3617,N_7,N_633);
xor U3618 (N_3618,N_393,N_448);
or U3619 (N_3619,N_495,N_343);
nor U3620 (N_3620,N_1084,N_2472);
or U3621 (N_3621,N_810,N_290);
nor U3622 (N_3622,N_2484,N_2407);
and U3623 (N_3623,N_2038,N_1428);
or U3624 (N_3624,N_899,N_537);
nor U3625 (N_3625,N_2120,N_1283);
or U3626 (N_3626,N_1841,N_2122);
or U3627 (N_3627,N_1973,N_1756);
nor U3628 (N_3628,N_2409,N_1246);
and U3629 (N_3629,N_93,N_279);
or U3630 (N_3630,N_98,N_2056);
nor U3631 (N_3631,N_1228,N_797);
nand U3632 (N_3632,N_162,N_2141);
and U3633 (N_3633,N_298,N_1809);
and U3634 (N_3634,N_1851,N_590);
or U3635 (N_3635,N_374,N_2431);
nor U3636 (N_3636,N_438,N_1561);
or U3637 (N_3637,N_488,N_1455);
and U3638 (N_3638,N_189,N_608);
and U3639 (N_3639,N_2066,N_1144);
and U3640 (N_3640,N_381,N_1934);
xnor U3641 (N_3641,N_2450,N_2031);
and U3642 (N_3642,N_2131,N_1833);
and U3643 (N_3643,N_1363,N_1209);
nand U3644 (N_3644,N_2133,N_1807);
and U3645 (N_3645,N_1602,N_939);
or U3646 (N_3646,N_1539,N_2318);
or U3647 (N_3647,N_1517,N_2398);
nand U3648 (N_3648,N_1020,N_1733);
nand U3649 (N_3649,N_661,N_1883);
nor U3650 (N_3650,N_283,N_976);
xnor U3651 (N_3651,N_542,N_2048);
nor U3652 (N_3652,N_1205,N_912);
nor U3653 (N_3653,N_1192,N_1641);
or U3654 (N_3654,N_1313,N_2188);
nor U3655 (N_3655,N_362,N_104);
or U3656 (N_3656,N_1164,N_1289);
nand U3657 (N_3657,N_1597,N_1518);
nand U3658 (N_3658,N_2481,N_358);
and U3659 (N_3659,N_2093,N_2376);
nor U3660 (N_3660,N_2262,N_2257);
nor U3661 (N_3661,N_1297,N_2285);
or U3662 (N_3662,N_1718,N_1538);
and U3663 (N_3663,N_2119,N_491);
and U3664 (N_3664,N_2165,N_761);
nand U3665 (N_3665,N_1692,N_1261);
and U3666 (N_3666,N_1168,N_1056);
nand U3667 (N_3667,N_483,N_1378);
nor U3668 (N_3668,N_736,N_1091);
nor U3669 (N_3669,N_1290,N_180);
or U3670 (N_3670,N_1494,N_75);
xor U3671 (N_3671,N_913,N_2276);
nor U3672 (N_3672,N_1502,N_2020);
and U3673 (N_3673,N_1954,N_1516);
or U3674 (N_3674,N_136,N_759);
or U3675 (N_3675,N_2261,N_1239);
nand U3676 (N_3676,N_2128,N_1434);
nand U3677 (N_3677,N_1996,N_1765);
xor U3678 (N_3678,N_1706,N_473);
or U3679 (N_3679,N_2342,N_1820);
or U3680 (N_3680,N_2441,N_2139);
nor U3681 (N_3681,N_2009,N_1684);
nor U3682 (N_3682,N_1478,N_348);
and U3683 (N_3683,N_1746,N_600);
and U3684 (N_3684,N_1744,N_286);
nand U3685 (N_3685,N_610,N_2291);
nand U3686 (N_3686,N_1818,N_2478);
nor U3687 (N_3687,N_1731,N_2089);
and U3688 (N_3688,N_1512,N_1465);
nor U3689 (N_3689,N_624,N_252);
and U3690 (N_3690,N_1994,N_2074);
and U3691 (N_3691,N_357,N_1656);
and U3692 (N_3692,N_1189,N_2064);
nand U3693 (N_3693,N_20,N_2013);
or U3694 (N_3694,N_941,N_1842);
and U3695 (N_3695,N_334,N_341);
and U3696 (N_3696,N_2358,N_1911);
nand U3697 (N_3697,N_1553,N_997);
nor U3698 (N_3698,N_1685,N_846);
or U3699 (N_3699,N_2395,N_828);
nor U3700 (N_3700,N_560,N_703);
nand U3701 (N_3701,N_1848,N_1390);
xnor U3702 (N_3702,N_360,N_586);
and U3703 (N_3703,N_581,N_1769);
and U3704 (N_3704,N_1591,N_731);
nor U3705 (N_3705,N_2209,N_2317);
nor U3706 (N_3706,N_1986,N_1183);
or U3707 (N_3707,N_1065,N_2054);
nor U3708 (N_3708,N_2016,N_1799);
nand U3709 (N_3709,N_619,N_213);
or U3710 (N_3710,N_335,N_50);
nor U3711 (N_3711,N_202,N_516);
nand U3712 (N_3712,N_786,N_569);
nor U3713 (N_3713,N_1504,N_1679);
nand U3714 (N_3714,N_2204,N_1529);
nand U3715 (N_3715,N_2343,N_259);
nor U3716 (N_3716,N_794,N_2309);
nor U3717 (N_3717,N_29,N_636);
nor U3718 (N_3718,N_1271,N_1101);
nand U3719 (N_3719,N_1356,N_2182);
nor U3720 (N_3720,N_1515,N_1910);
nor U3721 (N_3721,N_1248,N_1608);
nor U3722 (N_3722,N_922,N_1550);
nand U3723 (N_3723,N_791,N_118);
or U3724 (N_3724,N_1868,N_2058);
nor U3725 (N_3725,N_2384,N_1233);
or U3726 (N_3726,N_1024,N_1443);
nor U3727 (N_3727,N_840,N_1120);
nand U3728 (N_3728,N_2349,N_1114);
nor U3729 (N_3729,N_523,N_1864);
or U3730 (N_3730,N_738,N_1873);
nand U3731 (N_3731,N_2443,N_827);
and U3732 (N_3732,N_1905,N_1875);
or U3733 (N_3733,N_628,N_946);
nor U3734 (N_3734,N_363,N_2092);
or U3735 (N_3735,N_1153,N_2448);
nor U3736 (N_3736,N_2027,N_1979);
and U3737 (N_3737,N_1310,N_2422);
or U3738 (N_3738,N_84,N_2294);
nand U3739 (N_3739,N_1802,N_1581);
nand U3740 (N_3740,N_1069,N_1033);
and U3741 (N_3741,N_1902,N_1877);
nand U3742 (N_3742,N_907,N_1031);
or U3743 (N_3743,N_2023,N_14);
nand U3744 (N_3744,N_185,N_2447);
or U3745 (N_3745,N_418,N_742);
xnor U3746 (N_3746,N_1639,N_2006);
and U3747 (N_3747,N_1298,N_1150);
or U3748 (N_3748,N_714,N_1269);
and U3749 (N_3749,N_1951,N_1888);
and U3750 (N_3750,N_349,N_2245);
or U3751 (N_3751,N_2307,N_2433);
nand U3752 (N_3752,N_1834,N_762);
nor U3753 (N_3753,N_1132,N_738);
and U3754 (N_3754,N_242,N_2106);
nor U3755 (N_3755,N_651,N_271);
nor U3756 (N_3756,N_1684,N_2200);
nor U3757 (N_3757,N_1133,N_1654);
and U3758 (N_3758,N_275,N_416);
nor U3759 (N_3759,N_1492,N_230);
and U3760 (N_3760,N_985,N_1378);
nor U3761 (N_3761,N_975,N_1854);
nand U3762 (N_3762,N_106,N_36);
nor U3763 (N_3763,N_358,N_1268);
nand U3764 (N_3764,N_540,N_1697);
and U3765 (N_3765,N_326,N_2271);
or U3766 (N_3766,N_746,N_12);
nor U3767 (N_3767,N_1171,N_2032);
and U3768 (N_3768,N_2308,N_660);
or U3769 (N_3769,N_1806,N_2363);
or U3770 (N_3770,N_1582,N_1953);
nand U3771 (N_3771,N_894,N_665);
nand U3772 (N_3772,N_972,N_72);
nand U3773 (N_3773,N_28,N_339);
xor U3774 (N_3774,N_1896,N_730);
and U3775 (N_3775,N_214,N_903);
or U3776 (N_3776,N_2336,N_1408);
nand U3777 (N_3777,N_743,N_85);
or U3778 (N_3778,N_1931,N_698);
and U3779 (N_3779,N_1344,N_236);
nand U3780 (N_3780,N_2318,N_2406);
xnor U3781 (N_3781,N_291,N_2268);
or U3782 (N_3782,N_1607,N_1137);
nor U3783 (N_3783,N_2055,N_1205);
or U3784 (N_3784,N_658,N_450);
and U3785 (N_3785,N_177,N_2136);
and U3786 (N_3786,N_1184,N_2075);
and U3787 (N_3787,N_458,N_641);
or U3788 (N_3788,N_2003,N_311);
nand U3789 (N_3789,N_1882,N_859);
nand U3790 (N_3790,N_1195,N_1181);
nand U3791 (N_3791,N_1538,N_351);
nand U3792 (N_3792,N_276,N_595);
nand U3793 (N_3793,N_1731,N_374);
nor U3794 (N_3794,N_1766,N_1647);
and U3795 (N_3795,N_12,N_519);
xnor U3796 (N_3796,N_2184,N_961);
nand U3797 (N_3797,N_485,N_1410);
nand U3798 (N_3798,N_1696,N_923);
nand U3799 (N_3799,N_1888,N_2273);
nor U3800 (N_3800,N_1934,N_2467);
nor U3801 (N_3801,N_329,N_2058);
nor U3802 (N_3802,N_1274,N_1977);
nor U3803 (N_3803,N_2333,N_2136);
and U3804 (N_3804,N_272,N_277);
or U3805 (N_3805,N_938,N_1306);
or U3806 (N_3806,N_1309,N_1097);
nand U3807 (N_3807,N_1838,N_83);
or U3808 (N_3808,N_356,N_123);
and U3809 (N_3809,N_8,N_1719);
and U3810 (N_3810,N_1718,N_176);
nand U3811 (N_3811,N_1922,N_1547);
nand U3812 (N_3812,N_2278,N_1303);
and U3813 (N_3813,N_957,N_1607);
and U3814 (N_3814,N_2300,N_1475);
and U3815 (N_3815,N_928,N_2035);
nand U3816 (N_3816,N_113,N_762);
and U3817 (N_3817,N_1039,N_345);
nor U3818 (N_3818,N_1680,N_1196);
or U3819 (N_3819,N_1908,N_2006);
or U3820 (N_3820,N_1087,N_2329);
nand U3821 (N_3821,N_447,N_2044);
nand U3822 (N_3822,N_1169,N_1152);
and U3823 (N_3823,N_1472,N_1857);
nand U3824 (N_3824,N_242,N_347);
nand U3825 (N_3825,N_584,N_2385);
nor U3826 (N_3826,N_1361,N_752);
nand U3827 (N_3827,N_1955,N_2395);
and U3828 (N_3828,N_479,N_52);
and U3829 (N_3829,N_424,N_1218);
nor U3830 (N_3830,N_2364,N_1595);
and U3831 (N_3831,N_1672,N_1222);
or U3832 (N_3832,N_93,N_238);
and U3833 (N_3833,N_10,N_730);
or U3834 (N_3834,N_2046,N_517);
nand U3835 (N_3835,N_1729,N_2450);
nor U3836 (N_3836,N_1007,N_112);
nand U3837 (N_3837,N_1784,N_765);
and U3838 (N_3838,N_2225,N_1369);
or U3839 (N_3839,N_754,N_671);
and U3840 (N_3840,N_1026,N_504);
nand U3841 (N_3841,N_313,N_950);
or U3842 (N_3842,N_1795,N_373);
and U3843 (N_3843,N_247,N_2072);
and U3844 (N_3844,N_1428,N_2477);
nor U3845 (N_3845,N_2173,N_1474);
or U3846 (N_3846,N_85,N_757);
nand U3847 (N_3847,N_635,N_534);
nand U3848 (N_3848,N_1720,N_569);
nor U3849 (N_3849,N_2048,N_1563);
and U3850 (N_3850,N_1,N_9);
or U3851 (N_3851,N_2425,N_980);
nor U3852 (N_3852,N_1945,N_2006);
nor U3853 (N_3853,N_2402,N_216);
and U3854 (N_3854,N_1667,N_201);
nand U3855 (N_3855,N_1631,N_1064);
nor U3856 (N_3856,N_616,N_101);
and U3857 (N_3857,N_354,N_1550);
xnor U3858 (N_3858,N_712,N_2196);
xnor U3859 (N_3859,N_2235,N_1449);
nor U3860 (N_3860,N_542,N_598);
xor U3861 (N_3861,N_1239,N_2497);
and U3862 (N_3862,N_2100,N_148);
and U3863 (N_3863,N_2244,N_2192);
or U3864 (N_3864,N_1165,N_2175);
nor U3865 (N_3865,N_1882,N_1840);
and U3866 (N_3866,N_642,N_1281);
or U3867 (N_3867,N_438,N_1607);
or U3868 (N_3868,N_2455,N_1792);
and U3869 (N_3869,N_1879,N_1367);
and U3870 (N_3870,N_2437,N_2392);
nand U3871 (N_3871,N_892,N_1291);
nand U3872 (N_3872,N_388,N_2142);
nor U3873 (N_3873,N_631,N_668);
nor U3874 (N_3874,N_1815,N_956);
or U3875 (N_3875,N_2054,N_412);
or U3876 (N_3876,N_1665,N_691);
and U3877 (N_3877,N_843,N_2122);
nand U3878 (N_3878,N_1596,N_2239);
nor U3879 (N_3879,N_592,N_842);
or U3880 (N_3880,N_2211,N_1859);
nor U3881 (N_3881,N_1978,N_1582);
nand U3882 (N_3882,N_1910,N_1116);
or U3883 (N_3883,N_288,N_1643);
and U3884 (N_3884,N_1188,N_2148);
or U3885 (N_3885,N_1803,N_80);
or U3886 (N_3886,N_1383,N_212);
or U3887 (N_3887,N_1978,N_1350);
nand U3888 (N_3888,N_1721,N_336);
or U3889 (N_3889,N_1342,N_2494);
nor U3890 (N_3890,N_1399,N_375);
and U3891 (N_3891,N_1445,N_1992);
and U3892 (N_3892,N_152,N_2140);
xor U3893 (N_3893,N_1110,N_793);
or U3894 (N_3894,N_2076,N_1979);
or U3895 (N_3895,N_2107,N_2165);
nor U3896 (N_3896,N_1136,N_1112);
or U3897 (N_3897,N_589,N_1040);
and U3898 (N_3898,N_1884,N_305);
nor U3899 (N_3899,N_1935,N_150);
xnor U3900 (N_3900,N_2103,N_348);
nand U3901 (N_3901,N_471,N_1015);
nor U3902 (N_3902,N_2390,N_1030);
nand U3903 (N_3903,N_1487,N_2453);
and U3904 (N_3904,N_1379,N_1871);
nor U3905 (N_3905,N_1664,N_1153);
nand U3906 (N_3906,N_644,N_2470);
and U3907 (N_3907,N_1389,N_1962);
or U3908 (N_3908,N_856,N_1593);
and U3909 (N_3909,N_1526,N_192);
or U3910 (N_3910,N_955,N_1126);
nor U3911 (N_3911,N_462,N_582);
xor U3912 (N_3912,N_1482,N_1572);
nor U3913 (N_3913,N_1891,N_2024);
xnor U3914 (N_3914,N_2271,N_2343);
nand U3915 (N_3915,N_1588,N_1313);
nand U3916 (N_3916,N_1415,N_910);
nand U3917 (N_3917,N_686,N_1636);
nand U3918 (N_3918,N_348,N_1375);
or U3919 (N_3919,N_1151,N_640);
and U3920 (N_3920,N_2426,N_830);
nand U3921 (N_3921,N_2483,N_221);
or U3922 (N_3922,N_2274,N_599);
nor U3923 (N_3923,N_1131,N_2167);
nor U3924 (N_3924,N_792,N_247);
nand U3925 (N_3925,N_867,N_455);
nand U3926 (N_3926,N_2031,N_1880);
and U3927 (N_3927,N_638,N_2164);
nor U3928 (N_3928,N_1554,N_171);
or U3929 (N_3929,N_2091,N_204);
nor U3930 (N_3930,N_1809,N_1185);
or U3931 (N_3931,N_1552,N_1258);
and U3932 (N_3932,N_2309,N_2003);
nand U3933 (N_3933,N_830,N_1890);
xor U3934 (N_3934,N_2152,N_1857);
nor U3935 (N_3935,N_1124,N_129);
nor U3936 (N_3936,N_1926,N_1154);
and U3937 (N_3937,N_1185,N_508);
and U3938 (N_3938,N_1437,N_1868);
and U3939 (N_3939,N_453,N_2443);
and U3940 (N_3940,N_1763,N_1495);
and U3941 (N_3941,N_584,N_1340);
nor U3942 (N_3942,N_1565,N_259);
nor U3943 (N_3943,N_1041,N_230);
nor U3944 (N_3944,N_170,N_1633);
and U3945 (N_3945,N_1236,N_2365);
and U3946 (N_3946,N_2100,N_1508);
nor U3947 (N_3947,N_2351,N_683);
or U3948 (N_3948,N_494,N_2473);
nor U3949 (N_3949,N_1651,N_1260);
or U3950 (N_3950,N_1762,N_356);
nor U3951 (N_3951,N_1056,N_600);
nand U3952 (N_3952,N_2000,N_1331);
nor U3953 (N_3953,N_1272,N_254);
and U3954 (N_3954,N_2493,N_2443);
nand U3955 (N_3955,N_158,N_855);
and U3956 (N_3956,N_229,N_1127);
nand U3957 (N_3957,N_824,N_1681);
or U3958 (N_3958,N_1260,N_1316);
or U3959 (N_3959,N_437,N_1725);
nand U3960 (N_3960,N_1779,N_1003);
nor U3961 (N_3961,N_942,N_1403);
nor U3962 (N_3962,N_1465,N_875);
or U3963 (N_3963,N_589,N_1052);
or U3964 (N_3964,N_527,N_417);
nor U3965 (N_3965,N_1429,N_177);
nand U3966 (N_3966,N_195,N_2309);
or U3967 (N_3967,N_1221,N_1784);
nand U3968 (N_3968,N_1852,N_1407);
and U3969 (N_3969,N_1311,N_1875);
nor U3970 (N_3970,N_1655,N_2419);
and U3971 (N_3971,N_2044,N_906);
and U3972 (N_3972,N_2325,N_1241);
nor U3973 (N_3973,N_1408,N_1978);
or U3974 (N_3974,N_363,N_701);
or U3975 (N_3975,N_2344,N_1404);
nand U3976 (N_3976,N_357,N_1725);
or U3977 (N_3977,N_2048,N_2385);
or U3978 (N_3978,N_753,N_723);
and U3979 (N_3979,N_30,N_1757);
and U3980 (N_3980,N_1050,N_1323);
nand U3981 (N_3981,N_1695,N_728);
nand U3982 (N_3982,N_1642,N_1806);
and U3983 (N_3983,N_2009,N_533);
nor U3984 (N_3984,N_1838,N_1701);
or U3985 (N_3985,N_1446,N_1318);
or U3986 (N_3986,N_395,N_134);
or U3987 (N_3987,N_2214,N_957);
or U3988 (N_3988,N_1259,N_2048);
nand U3989 (N_3989,N_2204,N_1545);
nand U3990 (N_3990,N_1089,N_916);
and U3991 (N_3991,N_1604,N_460);
nand U3992 (N_3992,N_1738,N_2163);
or U3993 (N_3993,N_732,N_2206);
or U3994 (N_3994,N_148,N_846);
nor U3995 (N_3995,N_507,N_682);
nand U3996 (N_3996,N_975,N_2342);
nand U3997 (N_3997,N_1110,N_2045);
and U3998 (N_3998,N_214,N_912);
or U3999 (N_3999,N_1420,N_930);
nand U4000 (N_4000,N_1533,N_1323);
and U4001 (N_4001,N_1395,N_2355);
or U4002 (N_4002,N_1499,N_1772);
xnor U4003 (N_4003,N_2115,N_790);
or U4004 (N_4004,N_443,N_1060);
xor U4005 (N_4005,N_522,N_1958);
nor U4006 (N_4006,N_623,N_1522);
xnor U4007 (N_4007,N_2347,N_1528);
or U4008 (N_4008,N_811,N_57);
and U4009 (N_4009,N_1183,N_537);
nand U4010 (N_4010,N_1643,N_2025);
and U4011 (N_4011,N_746,N_1076);
and U4012 (N_4012,N_925,N_1118);
nand U4013 (N_4013,N_679,N_342);
nor U4014 (N_4014,N_1072,N_1475);
and U4015 (N_4015,N_1974,N_616);
nor U4016 (N_4016,N_1014,N_1591);
and U4017 (N_4017,N_987,N_1780);
and U4018 (N_4018,N_2306,N_246);
nor U4019 (N_4019,N_2078,N_2082);
and U4020 (N_4020,N_1923,N_2195);
nor U4021 (N_4021,N_637,N_651);
nor U4022 (N_4022,N_1560,N_2240);
nor U4023 (N_4023,N_313,N_2485);
or U4024 (N_4024,N_612,N_1294);
and U4025 (N_4025,N_2346,N_163);
nor U4026 (N_4026,N_2481,N_1027);
or U4027 (N_4027,N_821,N_208);
nor U4028 (N_4028,N_2259,N_1094);
nand U4029 (N_4029,N_1272,N_1245);
and U4030 (N_4030,N_1147,N_733);
nand U4031 (N_4031,N_665,N_1583);
or U4032 (N_4032,N_1037,N_557);
or U4033 (N_4033,N_2041,N_1806);
nor U4034 (N_4034,N_1320,N_495);
xnor U4035 (N_4035,N_947,N_2486);
nor U4036 (N_4036,N_1174,N_621);
nand U4037 (N_4037,N_246,N_2275);
and U4038 (N_4038,N_227,N_1361);
and U4039 (N_4039,N_2411,N_2404);
nor U4040 (N_4040,N_1474,N_1995);
or U4041 (N_4041,N_2350,N_498);
and U4042 (N_4042,N_495,N_577);
nor U4043 (N_4043,N_1359,N_947);
or U4044 (N_4044,N_2155,N_95);
nand U4045 (N_4045,N_749,N_1974);
xnor U4046 (N_4046,N_978,N_2382);
and U4047 (N_4047,N_1459,N_2328);
nor U4048 (N_4048,N_200,N_1507);
or U4049 (N_4049,N_2089,N_144);
xor U4050 (N_4050,N_1639,N_2431);
nand U4051 (N_4051,N_2121,N_1221);
and U4052 (N_4052,N_934,N_197);
and U4053 (N_4053,N_916,N_90);
and U4054 (N_4054,N_1579,N_485);
nand U4055 (N_4055,N_2190,N_133);
and U4056 (N_4056,N_1782,N_2334);
nor U4057 (N_4057,N_2488,N_1140);
nand U4058 (N_4058,N_2078,N_87);
nand U4059 (N_4059,N_2460,N_105);
or U4060 (N_4060,N_221,N_1454);
nor U4061 (N_4061,N_443,N_1926);
nand U4062 (N_4062,N_519,N_2224);
nor U4063 (N_4063,N_680,N_13);
and U4064 (N_4064,N_1018,N_1151);
nor U4065 (N_4065,N_363,N_669);
nor U4066 (N_4066,N_650,N_1970);
nor U4067 (N_4067,N_1318,N_1689);
and U4068 (N_4068,N_980,N_1355);
nor U4069 (N_4069,N_1844,N_1580);
xnor U4070 (N_4070,N_2272,N_2395);
or U4071 (N_4071,N_1387,N_920);
nor U4072 (N_4072,N_2035,N_621);
or U4073 (N_4073,N_961,N_115);
nand U4074 (N_4074,N_562,N_1168);
nor U4075 (N_4075,N_1218,N_868);
or U4076 (N_4076,N_1838,N_1979);
and U4077 (N_4077,N_223,N_1262);
nor U4078 (N_4078,N_2436,N_685);
nand U4079 (N_4079,N_983,N_2001);
nor U4080 (N_4080,N_2096,N_1216);
nand U4081 (N_4081,N_2452,N_2325);
and U4082 (N_4082,N_896,N_115);
or U4083 (N_4083,N_1038,N_1774);
xnor U4084 (N_4084,N_934,N_10);
and U4085 (N_4085,N_1179,N_1858);
nand U4086 (N_4086,N_2113,N_2267);
nand U4087 (N_4087,N_2414,N_2129);
or U4088 (N_4088,N_399,N_2358);
nand U4089 (N_4089,N_507,N_1810);
nor U4090 (N_4090,N_1294,N_1791);
nor U4091 (N_4091,N_2461,N_1597);
nor U4092 (N_4092,N_1756,N_243);
or U4093 (N_4093,N_2164,N_106);
and U4094 (N_4094,N_290,N_2159);
or U4095 (N_4095,N_1045,N_2260);
or U4096 (N_4096,N_861,N_559);
nor U4097 (N_4097,N_1352,N_1584);
and U4098 (N_4098,N_1919,N_155);
and U4099 (N_4099,N_1785,N_1285);
and U4100 (N_4100,N_1393,N_274);
or U4101 (N_4101,N_1142,N_1721);
nand U4102 (N_4102,N_786,N_2063);
and U4103 (N_4103,N_1184,N_725);
nor U4104 (N_4104,N_684,N_1297);
or U4105 (N_4105,N_746,N_1048);
or U4106 (N_4106,N_1582,N_1377);
nand U4107 (N_4107,N_1015,N_2286);
and U4108 (N_4108,N_958,N_1811);
xnor U4109 (N_4109,N_1475,N_353);
and U4110 (N_4110,N_1386,N_1753);
nor U4111 (N_4111,N_2246,N_656);
nor U4112 (N_4112,N_184,N_867);
or U4113 (N_4113,N_2147,N_895);
or U4114 (N_4114,N_213,N_573);
nand U4115 (N_4115,N_2272,N_1969);
or U4116 (N_4116,N_458,N_32);
nor U4117 (N_4117,N_584,N_1681);
or U4118 (N_4118,N_179,N_1859);
or U4119 (N_4119,N_1260,N_166);
or U4120 (N_4120,N_1016,N_108);
xor U4121 (N_4121,N_1466,N_1882);
and U4122 (N_4122,N_2018,N_1681);
nor U4123 (N_4123,N_2123,N_1516);
nand U4124 (N_4124,N_697,N_1746);
nand U4125 (N_4125,N_2379,N_1066);
or U4126 (N_4126,N_774,N_1900);
and U4127 (N_4127,N_2311,N_764);
nor U4128 (N_4128,N_326,N_485);
or U4129 (N_4129,N_1852,N_1124);
nor U4130 (N_4130,N_1071,N_53);
nand U4131 (N_4131,N_694,N_1021);
nand U4132 (N_4132,N_107,N_1639);
nor U4133 (N_4133,N_983,N_33);
nor U4134 (N_4134,N_1653,N_2198);
nand U4135 (N_4135,N_1153,N_5);
and U4136 (N_4136,N_2365,N_937);
and U4137 (N_4137,N_2206,N_570);
and U4138 (N_4138,N_1150,N_218);
and U4139 (N_4139,N_1182,N_1100);
xnor U4140 (N_4140,N_2230,N_224);
nand U4141 (N_4141,N_452,N_801);
nand U4142 (N_4142,N_1686,N_855);
and U4143 (N_4143,N_1819,N_856);
nor U4144 (N_4144,N_1583,N_1008);
nand U4145 (N_4145,N_731,N_2300);
nor U4146 (N_4146,N_2168,N_2407);
or U4147 (N_4147,N_108,N_360);
nand U4148 (N_4148,N_871,N_1510);
and U4149 (N_4149,N_89,N_212);
nand U4150 (N_4150,N_375,N_1022);
nor U4151 (N_4151,N_886,N_1921);
nand U4152 (N_4152,N_167,N_1918);
or U4153 (N_4153,N_698,N_144);
or U4154 (N_4154,N_1706,N_399);
nand U4155 (N_4155,N_219,N_1090);
nand U4156 (N_4156,N_2368,N_442);
nand U4157 (N_4157,N_2486,N_616);
nor U4158 (N_4158,N_292,N_539);
and U4159 (N_4159,N_668,N_558);
nor U4160 (N_4160,N_168,N_1053);
and U4161 (N_4161,N_581,N_359);
and U4162 (N_4162,N_509,N_212);
nor U4163 (N_4163,N_2473,N_1385);
or U4164 (N_4164,N_1054,N_1209);
or U4165 (N_4165,N_2395,N_2071);
nand U4166 (N_4166,N_548,N_1911);
nor U4167 (N_4167,N_248,N_433);
nand U4168 (N_4168,N_1585,N_2413);
nor U4169 (N_4169,N_1322,N_1608);
or U4170 (N_4170,N_1370,N_1612);
or U4171 (N_4171,N_1917,N_2295);
or U4172 (N_4172,N_1525,N_462);
nand U4173 (N_4173,N_1117,N_975);
or U4174 (N_4174,N_275,N_1870);
and U4175 (N_4175,N_2365,N_1284);
and U4176 (N_4176,N_512,N_593);
nand U4177 (N_4177,N_58,N_2063);
and U4178 (N_4178,N_1560,N_1920);
and U4179 (N_4179,N_735,N_333);
nor U4180 (N_4180,N_185,N_1950);
nor U4181 (N_4181,N_1659,N_530);
or U4182 (N_4182,N_2200,N_2497);
and U4183 (N_4183,N_1882,N_2065);
nand U4184 (N_4184,N_864,N_2478);
or U4185 (N_4185,N_1760,N_1311);
or U4186 (N_4186,N_903,N_2123);
or U4187 (N_4187,N_2344,N_437);
nor U4188 (N_4188,N_2230,N_1434);
and U4189 (N_4189,N_21,N_2330);
and U4190 (N_4190,N_2274,N_1500);
nand U4191 (N_4191,N_760,N_1847);
or U4192 (N_4192,N_611,N_125);
or U4193 (N_4193,N_1782,N_1683);
nor U4194 (N_4194,N_1232,N_7);
nor U4195 (N_4195,N_1338,N_2239);
or U4196 (N_4196,N_1,N_1428);
or U4197 (N_4197,N_848,N_1698);
or U4198 (N_4198,N_2366,N_1275);
xor U4199 (N_4199,N_1250,N_2246);
nor U4200 (N_4200,N_2436,N_1084);
nor U4201 (N_4201,N_170,N_1982);
nor U4202 (N_4202,N_822,N_1406);
nor U4203 (N_4203,N_1616,N_2250);
and U4204 (N_4204,N_486,N_925);
xnor U4205 (N_4205,N_1330,N_2150);
or U4206 (N_4206,N_1642,N_951);
nand U4207 (N_4207,N_2192,N_2080);
and U4208 (N_4208,N_275,N_947);
nand U4209 (N_4209,N_118,N_1564);
nor U4210 (N_4210,N_1760,N_1386);
and U4211 (N_4211,N_87,N_1106);
and U4212 (N_4212,N_2057,N_483);
and U4213 (N_4213,N_765,N_516);
and U4214 (N_4214,N_444,N_1113);
and U4215 (N_4215,N_2155,N_751);
or U4216 (N_4216,N_728,N_1236);
nor U4217 (N_4217,N_2171,N_2395);
and U4218 (N_4218,N_802,N_149);
nor U4219 (N_4219,N_2055,N_541);
or U4220 (N_4220,N_440,N_2352);
or U4221 (N_4221,N_1411,N_1550);
xnor U4222 (N_4222,N_1188,N_1157);
nor U4223 (N_4223,N_1903,N_2263);
and U4224 (N_4224,N_1034,N_1182);
or U4225 (N_4225,N_2249,N_919);
nor U4226 (N_4226,N_1228,N_472);
nand U4227 (N_4227,N_1034,N_2446);
and U4228 (N_4228,N_1012,N_77);
nor U4229 (N_4229,N_527,N_1231);
or U4230 (N_4230,N_2125,N_1075);
or U4231 (N_4231,N_2338,N_398);
nor U4232 (N_4232,N_26,N_1750);
and U4233 (N_4233,N_421,N_61);
nand U4234 (N_4234,N_1502,N_760);
nand U4235 (N_4235,N_769,N_791);
nand U4236 (N_4236,N_864,N_1267);
nand U4237 (N_4237,N_182,N_153);
nand U4238 (N_4238,N_1538,N_1886);
nand U4239 (N_4239,N_88,N_2040);
nor U4240 (N_4240,N_1157,N_576);
nor U4241 (N_4241,N_1745,N_2421);
and U4242 (N_4242,N_1227,N_2176);
or U4243 (N_4243,N_894,N_1010);
nand U4244 (N_4244,N_2187,N_124);
nand U4245 (N_4245,N_2423,N_2161);
and U4246 (N_4246,N_1828,N_427);
nand U4247 (N_4247,N_2360,N_1716);
or U4248 (N_4248,N_5,N_1400);
and U4249 (N_4249,N_2474,N_34);
nand U4250 (N_4250,N_1383,N_1246);
or U4251 (N_4251,N_843,N_1531);
xnor U4252 (N_4252,N_859,N_384);
nand U4253 (N_4253,N_517,N_2318);
and U4254 (N_4254,N_1618,N_2156);
or U4255 (N_4255,N_501,N_2388);
nor U4256 (N_4256,N_2339,N_92);
nor U4257 (N_4257,N_1125,N_125);
or U4258 (N_4258,N_1282,N_1498);
nor U4259 (N_4259,N_1821,N_226);
nand U4260 (N_4260,N_2345,N_672);
nand U4261 (N_4261,N_1318,N_2467);
nand U4262 (N_4262,N_123,N_2310);
nor U4263 (N_4263,N_1940,N_2189);
nor U4264 (N_4264,N_2408,N_869);
xnor U4265 (N_4265,N_2056,N_1873);
nor U4266 (N_4266,N_566,N_2097);
or U4267 (N_4267,N_2259,N_2349);
or U4268 (N_4268,N_303,N_1589);
or U4269 (N_4269,N_177,N_1551);
or U4270 (N_4270,N_559,N_1335);
or U4271 (N_4271,N_2099,N_1031);
or U4272 (N_4272,N_1101,N_702);
and U4273 (N_4273,N_985,N_96);
or U4274 (N_4274,N_1544,N_2224);
and U4275 (N_4275,N_216,N_2285);
or U4276 (N_4276,N_2318,N_911);
and U4277 (N_4277,N_1060,N_2143);
and U4278 (N_4278,N_912,N_2231);
nor U4279 (N_4279,N_2463,N_1425);
nand U4280 (N_4280,N_1894,N_2266);
or U4281 (N_4281,N_729,N_2109);
and U4282 (N_4282,N_995,N_2064);
nor U4283 (N_4283,N_1445,N_634);
nand U4284 (N_4284,N_1124,N_2308);
and U4285 (N_4285,N_2038,N_214);
or U4286 (N_4286,N_1171,N_347);
nor U4287 (N_4287,N_761,N_380);
nor U4288 (N_4288,N_928,N_923);
and U4289 (N_4289,N_925,N_1174);
nand U4290 (N_4290,N_1614,N_2207);
xor U4291 (N_4291,N_492,N_827);
nor U4292 (N_4292,N_1654,N_68);
nor U4293 (N_4293,N_1633,N_1679);
nor U4294 (N_4294,N_483,N_1250);
or U4295 (N_4295,N_1222,N_695);
and U4296 (N_4296,N_848,N_1959);
nand U4297 (N_4297,N_1998,N_372);
nand U4298 (N_4298,N_862,N_484);
nor U4299 (N_4299,N_1414,N_660);
or U4300 (N_4300,N_1165,N_1917);
nand U4301 (N_4301,N_2204,N_16);
nand U4302 (N_4302,N_2410,N_1942);
and U4303 (N_4303,N_622,N_1640);
or U4304 (N_4304,N_1515,N_2031);
nor U4305 (N_4305,N_1460,N_967);
or U4306 (N_4306,N_1760,N_2206);
nor U4307 (N_4307,N_2454,N_1584);
nand U4308 (N_4308,N_1045,N_506);
or U4309 (N_4309,N_671,N_201);
nor U4310 (N_4310,N_1397,N_653);
nor U4311 (N_4311,N_1237,N_2335);
or U4312 (N_4312,N_327,N_1891);
or U4313 (N_4313,N_1616,N_1578);
nor U4314 (N_4314,N_164,N_1003);
or U4315 (N_4315,N_1992,N_2033);
nor U4316 (N_4316,N_1034,N_1736);
or U4317 (N_4317,N_990,N_2031);
or U4318 (N_4318,N_75,N_23);
or U4319 (N_4319,N_1224,N_1640);
nor U4320 (N_4320,N_174,N_452);
or U4321 (N_4321,N_943,N_2170);
or U4322 (N_4322,N_2069,N_371);
or U4323 (N_4323,N_1071,N_1567);
nor U4324 (N_4324,N_2266,N_1492);
nand U4325 (N_4325,N_867,N_2460);
nor U4326 (N_4326,N_2065,N_592);
nand U4327 (N_4327,N_221,N_765);
or U4328 (N_4328,N_703,N_1466);
and U4329 (N_4329,N_290,N_745);
nor U4330 (N_4330,N_2092,N_432);
nor U4331 (N_4331,N_2074,N_801);
and U4332 (N_4332,N_2149,N_1150);
or U4333 (N_4333,N_2221,N_1249);
nand U4334 (N_4334,N_245,N_836);
nor U4335 (N_4335,N_626,N_427);
nand U4336 (N_4336,N_2175,N_341);
and U4337 (N_4337,N_744,N_1716);
nor U4338 (N_4338,N_2259,N_884);
nand U4339 (N_4339,N_1763,N_1675);
nor U4340 (N_4340,N_175,N_1185);
nor U4341 (N_4341,N_438,N_570);
and U4342 (N_4342,N_1959,N_2277);
and U4343 (N_4343,N_2313,N_1323);
or U4344 (N_4344,N_2308,N_903);
nand U4345 (N_4345,N_2093,N_751);
and U4346 (N_4346,N_1217,N_1123);
nor U4347 (N_4347,N_2193,N_399);
or U4348 (N_4348,N_1540,N_165);
and U4349 (N_4349,N_22,N_383);
or U4350 (N_4350,N_1243,N_325);
nor U4351 (N_4351,N_1538,N_1668);
or U4352 (N_4352,N_1420,N_251);
xnor U4353 (N_4353,N_2141,N_1948);
and U4354 (N_4354,N_1055,N_1744);
nor U4355 (N_4355,N_2106,N_1807);
xor U4356 (N_4356,N_2194,N_1881);
and U4357 (N_4357,N_2475,N_2260);
nand U4358 (N_4358,N_1994,N_2111);
or U4359 (N_4359,N_1165,N_922);
or U4360 (N_4360,N_1158,N_1793);
and U4361 (N_4361,N_1586,N_1467);
or U4362 (N_4362,N_2231,N_230);
or U4363 (N_4363,N_908,N_758);
and U4364 (N_4364,N_264,N_1792);
xor U4365 (N_4365,N_855,N_423);
nand U4366 (N_4366,N_740,N_1053);
nand U4367 (N_4367,N_1696,N_836);
and U4368 (N_4368,N_9,N_963);
or U4369 (N_4369,N_1567,N_475);
nand U4370 (N_4370,N_323,N_125);
nand U4371 (N_4371,N_372,N_795);
and U4372 (N_4372,N_2029,N_1820);
nand U4373 (N_4373,N_1900,N_539);
nor U4374 (N_4374,N_2225,N_1483);
or U4375 (N_4375,N_1533,N_1373);
nor U4376 (N_4376,N_1832,N_7);
and U4377 (N_4377,N_2154,N_1688);
nor U4378 (N_4378,N_1363,N_1392);
and U4379 (N_4379,N_70,N_2382);
nand U4380 (N_4380,N_2257,N_1941);
and U4381 (N_4381,N_1620,N_1051);
nor U4382 (N_4382,N_962,N_1231);
nand U4383 (N_4383,N_2354,N_2057);
nand U4384 (N_4384,N_805,N_1769);
xnor U4385 (N_4385,N_1995,N_2000);
or U4386 (N_4386,N_1157,N_1864);
nand U4387 (N_4387,N_929,N_1490);
nor U4388 (N_4388,N_123,N_646);
nor U4389 (N_4389,N_187,N_158);
nand U4390 (N_4390,N_192,N_161);
and U4391 (N_4391,N_1538,N_1910);
nand U4392 (N_4392,N_2265,N_2435);
or U4393 (N_4393,N_1471,N_1407);
and U4394 (N_4394,N_1806,N_2096);
nor U4395 (N_4395,N_38,N_1978);
and U4396 (N_4396,N_300,N_2358);
or U4397 (N_4397,N_448,N_1986);
nand U4398 (N_4398,N_163,N_525);
nor U4399 (N_4399,N_1134,N_1368);
and U4400 (N_4400,N_2199,N_1384);
or U4401 (N_4401,N_2387,N_2355);
nor U4402 (N_4402,N_1903,N_430);
or U4403 (N_4403,N_1421,N_1947);
nor U4404 (N_4404,N_804,N_1417);
and U4405 (N_4405,N_1414,N_340);
or U4406 (N_4406,N_380,N_729);
xnor U4407 (N_4407,N_1179,N_599);
xor U4408 (N_4408,N_263,N_2136);
xor U4409 (N_4409,N_1941,N_1660);
and U4410 (N_4410,N_2206,N_648);
or U4411 (N_4411,N_336,N_1726);
nand U4412 (N_4412,N_1819,N_118);
and U4413 (N_4413,N_1568,N_913);
or U4414 (N_4414,N_1788,N_1262);
nor U4415 (N_4415,N_1318,N_1935);
nor U4416 (N_4416,N_1194,N_2048);
nor U4417 (N_4417,N_2275,N_1331);
nand U4418 (N_4418,N_2061,N_331);
or U4419 (N_4419,N_1968,N_1641);
xnor U4420 (N_4420,N_1858,N_857);
and U4421 (N_4421,N_1095,N_69);
nor U4422 (N_4422,N_862,N_1845);
nor U4423 (N_4423,N_1043,N_2174);
nand U4424 (N_4424,N_912,N_1260);
or U4425 (N_4425,N_1419,N_228);
nor U4426 (N_4426,N_740,N_435);
or U4427 (N_4427,N_631,N_540);
and U4428 (N_4428,N_2436,N_556);
or U4429 (N_4429,N_1646,N_1809);
nand U4430 (N_4430,N_2175,N_2260);
and U4431 (N_4431,N_973,N_228);
and U4432 (N_4432,N_277,N_758);
nand U4433 (N_4433,N_248,N_546);
nand U4434 (N_4434,N_1675,N_832);
nand U4435 (N_4435,N_1576,N_488);
and U4436 (N_4436,N_1073,N_598);
or U4437 (N_4437,N_2057,N_0);
nor U4438 (N_4438,N_882,N_1938);
nor U4439 (N_4439,N_2327,N_774);
nor U4440 (N_4440,N_289,N_466);
nand U4441 (N_4441,N_1251,N_2346);
or U4442 (N_4442,N_1890,N_1905);
nand U4443 (N_4443,N_1057,N_1361);
nor U4444 (N_4444,N_2443,N_986);
nor U4445 (N_4445,N_1722,N_715);
and U4446 (N_4446,N_1663,N_904);
nand U4447 (N_4447,N_648,N_238);
nand U4448 (N_4448,N_1351,N_1827);
nor U4449 (N_4449,N_685,N_398);
nor U4450 (N_4450,N_987,N_952);
nor U4451 (N_4451,N_2098,N_2224);
or U4452 (N_4452,N_2370,N_916);
and U4453 (N_4453,N_2450,N_336);
nor U4454 (N_4454,N_114,N_336);
nor U4455 (N_4455,N_2477,N_2337);
nor U4456 (N_4456,N_2488,N_1772);
and U4457 (N_4457,N_1363,N_1636);
nand U4458 (N_4458,N_1015,N_806);
or U4459 (N_4459,N_2295,N_759);
nand U4460 (N_4460,N_1464,N_2387);
nand U4461 (N_4461,N_1299,N_317);
nand U4462 (N_4462,N_521,N_2261);
or U4463 (N_4463,N_16,N_1895);
or U4464 (N_4464,N_1855,N_985);
nor U4465 (N_4465,N_175,N_2245);
and U4466 (N_4466,N_1772,N_1490);
nand U4467 (N_4467,N_1532,N_1513);
nand U4468 (N_4468,N_1816,N_2115);
nand U4469 (N_4469,N_2262,N_1975);
nor U4470 (N_4470,N_1958,N_1821);
and U4471 (N_4471,N_272,N_1902);
nor U4472 (N_4472,N_294,N_439);
or U4473 (N_4473,N_1538,N_325);
nand U4474 (N_4474,N_2274,N_2218);
and U4475 (N_4475,N_875,N_549);
nor U4476 (N_4476,N_81,N_1439);
and U4477 (N_4477,N_361,N_1101);
or U4478 (N_4478,N_1538,N_113);
or U4479 (N_4479,N_410,N_2160);
nand U4480 (N_4480,N_718,N_1414);
nor U4481 (N_4481,N_928,N_2198);
and U4482 (N_4482,N_1956,N_1182);
or U4483 (N_4483,N_442,N_225);
nand U4484 (N_4484,N_1328,N_1509);
nor U4485 (N_4485,N_2214,N_1545);
nor U4486 (N_4486,N_113,N_1205);
or U4487 (N_4487,N_2080,N_937);
nor U4488 (N_4488,N_1290,N_754);
and U4489 (N_4489,N_1983,N_86);
and U4490 (N_4490,N_1274,N_36);
nand U4491 (N_4491,N_594,N_1916);
or U4492 (N_4492,N_2259,N_1168);
or U4493 (N_4493,N_71,N_915);
or U4494 (N_4494,N_2472,N_2079);
or U4495 (N_4495,N_1649,N_1531);
nor U4496 (N_4496,N_1094,N_437);
nand U4497 (N_4497,N_157,N_1531);
or U4498 (N_4498,N_555,N_870);
and U4499 (N_4499,N_2394,N_624);
and U4500 (N_4500,N_279,N_1316);
nor U4501 (N_4501,N_1881,N_351);
or U4502 (N_4502,N_2046,N_1330);
nor U4503 (N_4503,N_966,N_677);
nor U4504 (N_4504,N_404,N_2164);
and U4505 (N_4505,N_286,N_507);
or U4506 (N_4506,N_1409,N_2432);
nand U4507 (N_4507,N_2468,N_741);
and U4508 (N_4508,N_514,N_1659);
or U4509 (N_4509,N_1068,N_2111);
nor U4510 (N_4510,N_1015,N_761);
nor U4511 (N_4511,N_598,N_1710);
nand U4512 (N_4512,N_1807,N_61);
nor U4513 (N_4513,N_903,N_1592);
nor U4514 (N_4514,N_828,N_648);
and U4515 (N_4515,N_1445,N_1413);
nand U4516 (N_4516,N_1962,N_1175);
or U4517 (N_4517,N_2121,N_1677);
xor U4518 (N_4518,N_2106,N_789);
or U4519 (N_4519,N_1354,N_307);
and U4520 (N_4520,N_1689,N_1904);
nand U4521 (N_4521,N_277,N_278);
and U4522 (N_4522,N_1822,N_1812);
and U4523 (N_4523,N_1005,N_979);
or U4524 (N_4524,N_66,N_18);
nand U4525 (N_4525,N_1130,N_848);
or U4526 (N_4526,N_9,N_1492);
or U4527 (N_4527,N_1524,N_2273);
and U4528 (N_4528,N_2047,N_1330);
and U4529 (N_4529,N_1502,N_1697);
xor U4530 (N_4530,N_1358,N_2490);
or U4531 (N_4531,N_544,N_1538);
and U4532 (N_4532,N_475,N_1008);
nand U4533 (N_4533,N_385,N_655);
xor U4534 (N_4534,N_2197,N_823);
and U4535 (N_4535,N_1364,N_258);
or U4536 (N_4536,N_863,N_1311);
and U4537 (N_4537,N_1278,N_250);
nor U4538 (N_4538,N_637,N_2060);
nor U4539 (N_4539,N_2177,N_2410);
or U4540 (N_4540,N_422,N_577);
nand U4541 (N_4541,N_1522,N_416);
nor U4542 (N_4542,N_1838,N_213);
or U4543 (N_4543,N_1618,N_1053);
or U4544 (N_4544,N_2098,N_1078);
nor U4545 (N_4545,N_1910,N_256);
nand U4546 (N_4546,N_902,N_355);
nor U4547 (N_4547,N_751,N_1759);
nor U4548 (N_4548,N_1572,N_912);
and U4549 (N_4549,N_769,N_155);
nor U4550 (N_4550,N_823,N_1427);
and U4551 (N_4551,N_804,N_2026);
nor U4552 (N_4552,N_1725,N_1435);
or U4553 (N_4553,N_1121,N_1194);
or U4554 (N_4554,N_661,N_425);
and U4555 (N_4555,N_2470,N_2277);
nand U4556 (N_4556,N_789,N_1341);
and U4557 (N_4557,N_64,N_1328);
and U4558 (N_4558,N_2230,N_2263);
nor U4559 (N_4559,N_195,N_2393);
nor U4560 (N_4560,N_266,N_1585);
or U4561 (N_4561,N_1219,N_1734);
and U4562 (N_4562,N_1564,N_1450);
nand U4563 (N_4563,N_2489,N_1047);
nand U4564 (N_4564,N_1660,N_735);
nand U4565 (N_4565,N_468,N_2092);
nor U4566 (N_4566,N_818,N_2329);
and U4567 (N_4567,N_367,N_356);
and U4568 (N_4568,N_921,N_719);
or U4569 (N_4569,N_1264,N_1374);
nor U4570 (N_4570,N_1894,N_406);
nand U4571 (N_4571,N_773,N_1438);
and U4572 (N_4572,N_2199,N_1302);
nor U4573 (N_4573,N_983,N_1642);
xor U4574 (N_4574,N_1226,N_1577);
and U4575 (N_4575,N_1861,N_1327);
nand U4576 (N_4576,N_1203,N_1704);
nor U4577 (N_4577,N_1499,N_1047);
nand U4578 (N_4578,N_1005,N_1813);
and U4579 (N_4579,N_1942,N_1020);
nand U4580 (N_4580,N_1404,N_3);
nor U4581 (N_4581,N_1716,N_2385);
nand U4582 (N_4582,N_1750,N_1218);
nor U4583 (N_4583,N_2361,N_433);
and U4584 (N_4584,N_1672,N_2324);
nor U4585 (N_4585,N_1010,N_2266);
or U4586 (N_4586,N_707,N_2039);
and U4587 (N_4587,N_2022,N_2383);
nor U4588 (N_4588,N_1556,N_583);
nand U4589 (N_4589,N_173,N_982);
nor U4590 (N_4590,N_382,N_47);
nor U4591 (N_4591,N_600,N_1929);
nor U4592 (N_4592,N_1311,N_2238);
and U4593 (N_4593,N_1718,N_663);
nor U4594 (N_4594,N_216,N_2339);
and U4595 (N_4595,N_480,N_2218);
nor U4596 (N_4596,N_2251,N_724);
nor U4597 (N_4597,N_325,N_2026);
nand U4598 (N_4598,N_701,N_1770);
and U4599 (N_4599,N_148,N_1753);
nand U4600 (N_4600,N_145,N_676);
or U4601 (N_4601,N_55,N_1060);
nor U4602 (N_4602,N_1813,N_1404);
xnor U4603 (N_4603,N_1761,N_2405);
nand U4604 (N_4604,N_123,N_77);
nand U4605 (N_4605,N_2491,N_274);
and U4606 (N_4606,N_2214,N_886);
nand U4607 (N_4607,N_1329,N_2204);
nor U4608 (N_4608,N_543,N_2015);
nor U4609 (N_4609,N_1944,N_2315);
nand U4610 (N_4610,N_2407,N_1912);
nand U4611 (N_4611,N_577,N_759);
nor U4612 (N_4612,N_251,N_2363);
or U4613 (N_4613,N_556,N_1111);
nor U4614 (N_4614,N_1615,N_536);
or U4615 (N_4615,N_2322,N_981);
and U4616 (N_4616,N_1688,N_1857);
or U4617 (N_4617,N_1761,N_2381);
or U4618 (N_4618,N_1581,N_2045);
and U4619 (N_4619,N_842,N_128);
and U4620 (N_4620,N_1520,N_2017);
nor U4621 (N_4621,N_11,N_1196);
and U4622 (N_4622,N_105,N_101);
or U4623 (N_4623,N_941,N_715);
nor U4624 (N_4624,N_2335,N_1703);
and U4625 (N_4625,N_157,N_656);
nor U4626 (N_4626,N_1836,N_2275);
nor U4627 (N_4627,N_1119,N_225);
nor U4628 (N_4628,N_27,N_742);
nand U4629 (N_4629,N_1096,N_1209);
and U4630 (N_4630,N_1223,N_2484);
nor U4631 (N_4631,N_243,N_1893);
nand U4632 (N_4632,N_1964,N_2473);
nand U4633 (N_4633,N_1432,N_87);
and U4634 (N_4634,N_211,N_2401);
and U4635 (N_4635,N_922,N_988);
nand U4636 (N_4636,N_2113,N_1310);
or U4637 (N_4637,N_372,N_251);
and U4638 (N_4638,N_2253,N_89);
xor U4639 (N_4639,N_2475,N_1623);
nand U4640 (N_4640,N_2362,N_1935);
nand U4641 (N_4641,N_2190,N_771);
and U4642 (N_4642,N_1089,N_165);
nor U4643 (N_4643,N_1969,N_2317);
nand U4644 (N_4644,N_162,N_243);
and U4645 (N_4645,N_1035,N_2332);
nand U4646 (N_4646,N_161,N_254);
or U4647 (N_4647,N_272,N_1875);
and U4648 (N_4648,N_564,N_209);
nor U4649 (N_4649,N_1602,N_1585);
nand U4650 (N_4650,N_971,N_2365);
or U4651 (N_4651,N_951,N_1265);
nor U4652 (N_4652,N_2153,N_2248);
and U4653 (N_4653,N_1667,N_2185);
nor U4654 (N_4654,N_1714,N_2316);
and U4655 (N_4655,N_679,N_1246);
xnor U4656 (N_4656,N_1212,N_1771);
and U4657 (N_4657,N_228,N_1857);
and U4658 (N_4658,N_1587,N_1040);
and U4659 (N_4659,N_143,N_1310);
nand U4660 (N_4660,N_1042,N_341);
nor U4661 (N_4661,N_1764,N_216);
or U4662 (N_4662,N_165,N_2157);
nor U4663 (N_4663,N_1576,N_1175);
or U4664 (N_4664,N_1357,N_1403);
or U4665 (N_4665,N_1372,N_1726);
and U4666 (N_4666,N_2326,N_619);
or U4667 (N_4667,N_587,N_931);
and U4668 (N_4668,N_1603,N_724);
xor U4669 (N_4669,N_1069,N_1556);
and U4670 (N_4670,N_2144,N_1141);
and U4671 (N_4671,N_1851,N_379);
and U4672 (N_4672,N_899,N_1513);
or U4673 (N_4673,N_2027,N_2055);
or U4674 (N_4674,N_2290,N_0);
xnor U4675 (N_4675,N_508,N_1445);
and U4676 (N_4676,N_2127,N_1248);
and U4677 (N_4677,N_848,N_650);
nor U4678 (N_4678,N_363,N_940);
nor U4679 (N_4679,N_792,N_31);
nand U4680 (N_4680,N_367,N_1327);
or U4681 (N_4681,N_1113,N_643);
nand U4682 (N_4682,N_714,N_924);
and U4683 (N_4683,N_164,N_1923);
or U4684 (N_4684,N_1343,N_1005);
nand U4685 (N_4685,N_1441,N_61);
and U4686 (N_4686,N_2087,N_1742);
or U4687 (N_4687,N_91,N_724);
nand U4688 (N_4688,N_2058,N_2306);
nor U4689 (N_4689,N_26,N_792);
nor U4690 (N_4690,N_1586,N_1354);
and U4691 (N_4691,N_1122,N_2341);
or U4692 (N_4692,N_833,N_227);
nor U4693 (N_4693,N_1925,N_540);
nor U4694 (N_4694,N_216,N_2472);
nand U4695 (N_4695,N_1074,N_2232);
nand U4696 (N_4696,N_1055,N_2070);
nand U4697 (N_4697,N_2412,N_2379);
and U4698 (N_4698,N_439,N_722);
and U4699 (N_4699,N_898,N_526);
nor U4700 (N_4700,N_26,N_488);
nor U4701 (N_4701,N_347,N_1947);
nand U4702 (N_4702,N_423,N_687);
or U4703 (N_4703,N_1019,N_899);
or U4704 (N_4704,N_464,N_535);
or U4705 (N_4705,N_889,N_2004);
xnor U4706 (N_4706,N_700,N_1653);
or U4707 (N_4707,N_724,N_1460);
or U4708 (N_4708,N_1553,N_1753);
and U4709 (N_4709,N_196,N_255);
and U4710 (N_4710,N_1400,N_1575);
or U4711 (N_4711,N_2335,N_755);
nand U4712 (N_4712,N_1688,N_1862);
and U4713 (N_4713,N_1734,N_2338);
nor U4714 (N_4714,N_20,N_1758);
and U4715 (N_4715,N_1473,N_1973);
nand U4716 (N_4716,N_1649,N_2053);
or U4717 (N_4717,N_1868,N_1422);
or U4718 (N_4718,N_1641,N_2317);
nor U4719 (N_4719,N_1426,N_1434);
or U4720 (N_4720,N_2166,N_1926);
xor U4721 (N_4721,N_988,N_632);
or U4722 (N_4722,N_2456,N_1296);
nand U4723 (N_4723,N_1114,N_599);
nand U4724 (N_4724,N_266,N_1155);
and U4725 (N_4725,N_142,N_1203);
or U4726 (N_4726,N_1915,N_1638);
and U4727 (N_4727,N_954,N_426);
nand U4728 (N_4728,N_293,N_31);
and U4729 (N_4729,N_491,N_1561);
nand U4730 (N_4730,N_1601,N_1785);
nand U4731 (N_4731,N_256,N_2376);
nand U4732 (N_4732,N_2249,N_2468);
and U4733 (N_4733,N_2127,N_2195);
or U4734 (N_4734,N_1206,N_2064);
nand U4735 (N_4735,N_231,N_755);
or U4736 (N_4736,N_805,N_1729);
and U4737 (N_4737,N_1151,N_2161);
nor U4738 (N_4738,N_602,N_1313);
and U4739 (N_4739,N_419,N_2368);
nor U4740 (N_4740,N_847,N_296);
nor U4741 (N_4741,N_1752,N_2207);
and U4742 (N_4742,N_979,N_691);
and U4743 (N_4743,N_2486,N_319);
nor U4744 (N_4744,N_1570,N_307);
or U4745 (N_4745,N_613,N_1090);
or U4746 (N_4746,N_1920,N_1355);
or U4747 (N_4747,N_2135,N_826);
nand U4748 (N_4748,N_1747,N_1727);
nand U4749 (N_4749,N_1502,N_1543);
and U4750 (N_4750,N_1011,N_696);
and U4751 (N_4751,N_1021,N_2109);
and U4752 (N_4752,N_380,N_35);
nor U4753 (N_4753,N_1435,N_1263);
or U4754 (N_4754,N_56,N_622);
nand U4755 (N_4755,N_1961,N_1176);
nor U4756 (N_4756,N_1939,N_2464);
or U4757 (N_4757,N_1022,N_2062);
and U4758 (N_4758,N_1600,N_1793);
and U4759 (N_4759,N_2249,N_855);
nand U4760 (N_4760,N_2326,N_2041);
or U4761 (N_4761,N_2311,N_991);
nor U4762 (N_4762,N_1615,N_644);
and U4763 (N_4763,N_147,N_2106);
or U4764 (N_4764,N_2090,N_1140);
and U4765 (N_4765,N_542,N_1725);
or U4766 (N_4766,N_1313,N_370);
and U4767 (N_4767,N_2028,N_1674);
or U4768 (N_4768,N_1266,N_1796);
or U4769 (N_4769,N_2117,N_2203);
nor U4770 (N_4770,N_459,N_363);
nand U4771 (N_4771,N_18,N_1087);
or U4772 (N_4772,N_1286,N_286);
nand U4773 (N_4773,N_1866,N_823);
nor U4774 (N_4774,N_2406,N_1225);
or U4775 (N_4775,N_442,N_2293);
or U4776 (N_4776,N_22,N_2470);
nor U4777 (N_4777,N_2363,N_889);
and U4778 (N_4778,N_282,N_1314);
nand U4779 (N_4779,N_1242,N_651);
nor U4780 (N_4780,N_55,N_864);
nor U4781 (N_4781,N_2030,N_2429);
nor U4782 (N_4782,N_1596,N_2280);
nand U4783 (N_4783,N_1531,N_436);
nor U4784 (N_4784,N_642,N_1677);
nor U4785 (N_4785,N_210,N_395);
and U4786 (N_4786,N_1893,N_254);
nor U4787 (N_4787,N_1479,N_2083);
nand U4788 (N_4788,N_66,N_1281);
nor U4789 (N_4789,N_1528,N_464);
or U4790 (N_4790,N_1996,N_1428);
or U4791 (N_4791,N_1768,N_2257);
nor U4792 (N_4792,N_460,N_777);
and U4793 (N_4793,N_1675,N_1570);
or U4794 (N_4794,N_831,N_114);
nor U4795 (N_4795,N_680,N_941);
or U4796 (N_4796,N_2382,N_2229);
or U4797 (N_4797,N_604,N_1222);
and U4798 (N_4798,N_1724,N_2116);
or U4799 (N_4799,N_1385,N_955);
nand U4800 (N_4800,N_660,N_592);
or U4801 (N_4801,N_1327,N_194);
nand U4802 (N_4802,N_261,N_1103);
and U4803 (N_4803,N_1156,N_1215);
nand U4804 (N_4804,N_462,N_250);
nor U4805 (N_4805,N_1872,N_569);
and U4806 (N_4806,N_1810,N_465);
nand U4807 (N_4807,N_1459,N_1863);
nor U4808 (N_4808,N_589,N_1076);
nor U4809 (N_4809,N_1799,N_2034);
and U4810 (N_4810,N_449,N_1350);
nand U4811 (N_4811,N_2468,N_618);
and U4812 (N_4812,N_2225,N_191);
and U4813 (N_4813,N_830,N_942);
or U4814 (N_4814,N_1311,N_2216);
and U4815 (N_4815,N_792,N_1052);
nand U4816 (N_4816,N_1418,N_1015);
and U4817 (N_4817,N_1539,N_480);
nor U4818 (N_4818,N_2179,N_1289);
nor U4819 (N_4819,N_335,N_2333);
nand U4820 (N_4820,N_1743,N_235);
or U4821 (N_4821,N_714,N_2399);
and U4822 (N_4822,N_2212,N_181);
or U4823 (N_4823,N_904,N_179);
or U4824 (N_4824,N_356,N_81);
or U4825 (N_4825,N_850,N_335);
nor U4826 (N_4826,N_2150,N_2260);
nor U4827 (N_4827,N_1651,N_2324);
xor U4828 (N_4828,N_1396,N_1050);
or U4829 (N_4829,N_1611,N_656);
and U4830 (N_4830,N_379,N_1980);
nand U4831 (N_4831,N_1196,N_291);
or U4832 (N_4832,N_2066,N_41);
nor U4833 (N_4833,N_2199,N_790);
xnor U4834 (N_4834,N_269,N_6);
and U4835 (N_4835,N_861,N_2407);
nand U4836 (N_4836,N_1509,N_695);
and U4837 (N_4837,N_60,N_407);
nor U4838 (N_4838,N_695,N_867);
and U4839 (N_4839,N_2279,N_15);
nand U4840 (N_4840,N_1493,N_629);
nor U4841 (N_4841,N_1684,N_604);
or U4842 (N_4842,N_818,N_957);
xnor U4843 (N_4843,N_2382,N_2255);
or U4844 (N_4844,N_631,N_1708);
nand U4845 (N_4845,N_1850,N_200);
or U4846 (N_4846,N_903,N_1708);
and U4847 (N_4847,N_1805,N_358);
and U4848 (N_4848,N_900,N_425);
nor U4849 (N_4849,N_168,N_1416);
nand U4850 (N_4850,N_2017,N_1611);
or U4851 (N_4851,N_270,N_545);
nand U4852 (N_4852,N_1349,N_948);
and U4853 (N_4853,N_466,N_71);
or U4854 (N_4854,N_2342,N_729);
or U4855 (N_4855,N_366,N_2313);
nor U4856 (N_4856,N_987,N_744);
or U4857 (N_4857,N_2077,N_368);
nor U4858 (N_4858,N_1879,N_1011);
xnor U4859 (N_4859,N_1538,N_1318);
and U4860 (N_4860,N_1498,N_1782);
or U4861 (N_4861,N_115,N_641);
and U4862 (N_4862,N_1928,N_1625);
and U4863 (N_4863,N_1280,N_1635);
and U4864 (N_4864,N_1719,N_1745);
nand U4865 (N_4865,N_1647,N_1150);
nor U4866 (N_4866,N_343,N_1556);
nand U4867 (N_4867,N_1070,N_2202);
and U4868 (N_4868,N_850,N_1643);
nor U4869 (N_4869,N_1617,N_1267);
and U4870 (N_4870,N_709,N_729);
or U4871 (N_4871,N_1386,N_1743);
and U4872 (N_4872,N_687,N_1143);
or U4873 (N_4873,N_1323,N_643);
or U4874 (N_4874,N_1063,N_2492);
and U4875 (N_4875,N_468,N_2032);
or U4876 (N_4876,N_822,N_668);
nor U4877 (N_4877,N_798,N_379);
and U4878 (N_4878,N_432,N_1378);
and U4879 (N_4879,N_2286,N_1542);
or U4880 (N_4880,N_1634,N_325);
nand U4881 (N_4881,N_1998,N_215);
nor U4882 (N_4882,N_968,N_28);
and U4883 (N_4883,N_1755,N_283);
and U4884 (N_4884,N_1268,N_2060);
and U4885 (N_4885,N_1883,N_2407);
and U4886 (N_4886,N_1449,N_369);
nand U4887 (N_4887,N_2156,N_2420);
nor U4888 (N_4888,N_1161,N_1827);
and U4889 (N_4889,N_1571,N_869);
nor U4890 (N_4890,N_1100,N_693);
nor U4891 (N_4891,N_2445,N_2296);
nand U4892 (N_4892,N_1716,N_2158);
and U4893 (N_4893,N_970,N_373);
or U4894 (N_4894,N_2251,N_650);
nor U4895 (N_4895,N_467,N_121);
or U4896 (N_4896,N_136,N_111);
nand U4897 (N_4897,N_1524,N_656);
nor U4898 (N_4898,N_1426,N_35);
and U4899 (N_4899,N_1258,N_371);
and U4900 (N_4900,N_574,N_1192);
nand U4901 (N_4901,N_688,N_1709);
nand U4902 (N_4902,N_1639,N_195);
nand U4903 (N_4903,N_2285,N_2376);
and U4904 (N_4904,N_1617,N_1402);
or U4905 (N_4905,N_222,N_1077);
nand U4906 (N_4906,N_2411,N_2382);
and U4907 (N_4907,N_1081,N_1490);
or U4908 (N_4908,N_1637,N_396);
nor U4909 (N_4909,N_2345,N_2220);
or U4910 (N_4910,N_1070,N_357);
or U4911 (N_4911,N_1669,N_237);
or U4912 (N_4912,N_1482,N_209);
xor U4913 (N_4913,N_1716,N_79);
or U4914 (N_4914,N_2054,N_602);
nor U4915 (N_4915,N_782,N_732);
nor U4916 (N_4916,N_311,N_937);
and U4917 (N_4917,N_425,N_1020);
nor U4918 (N_4918,N_1878,N_1825);
nor U4919 (N_4919,N_1622,N_2027);
or U4920 (N_4920,N_1338,N_1598);
or U4921 (N_4921,N_1523,N_350);
and U4922 (N_4922,N_528,N_352);
or U4923 (N_4923,N_974,N_1280);
nand U4924 (N_4924,N_1180,N_2183);
xnor U4925 (N_4925,N_27,N_485);
nand U4926 (N_4926,N_1141,N_1623);
or U4927 (N_4927,N_124,N_2366);
nor U4928 (N_4928,N_414,N_1153);
nor U4929 (N_4929,N_998,N_1310);
nor U4930 (N_4930,N_1274,N_407);
nand U4931 (N_4931,N_1280,N_1214);
and U4932 (N_4932,N_776,N_2007);
or U4933 (N_4933,N_777,N_1855);
nor U4934 (N_4934,N_213,N_376);
nor U4935 (N_4935,N_1977,N_1141);
or U4936 (N_4936,N_1793,N_587);
and U4937 (N_4937,N_490,N_1299);
and U4938 (N_4938,N_610,N_186);
or U4939 (N_4939,N_1229,N_529);
or U4940 (N_4940,N_792,N_2435);
or U4941 (N_4941,N_1904,N_750);
and U4942 (N_4942,N_1223,N_566);
nand U4943 (N_4943,N_1941,N_30);
nor U4944 (N_4944,N_1065,N_845);
and U4945 (N_4945,N_73,N_2355);
or U4946 (N_4946,N_1690,N_1605);
or U4947 (N_4947,N_1634,N_973);
nand U4948 (N_4948,N_1333,N_676);
nor U4949 (N_4949,N_669,N_1258);
or U4950 (N_4950,N_2422,N_1651);
or U4951 (N_4951,N_1508,N_2054);
nand U4952 (N_4952,N_185,N_753);
nand U4953 (N_4953,N_17,N_1625);
and U4954 (N_4954,N_1168,N_1706);
or U4955 (N_4955,N_2207,N_579);
nand U4956 (N_4956,N_835,N_1970);
nand U4957 (N_4957,N_609,N_817);
nand U4958 (N_4958,N_1745,N_2229);
or U4959 (N_4959,N_1903,N_1119);
nor U4960 (N_4960,N_990,N_507);
nand U4961 (N_4961,N_690,N_1419);
nor U4962 (N_4962,N_434,N_1977);
or U4963 (N_4963,N_745,N_2481);
nor U4964 (N_4964,N_1784,N_1954);
or U4965 (N_4965,N_2194,N_577);
and U4966 (N_4966,N_1632,N_318);
and U4967 (N_4967,N_485,N_966);
and U4968 (N_4968,N_1261,N_739);
nand U4969 (N_4969,N_2017,N_1723);
and U4970 (N_4970,N_2486,N_1024);
or U4971 (N_4971,N_1231,N_1926);
nor U4972 (N_4972,N_422,N_1324);
nor U4973 (N_4973,N_990,N_1603);
nor U4974 (N_4974,N_1304,N_2314);
nand U4975 (N_4975,N_1962,N_1722);
and U4976 (N_4976,N_1518,N_130);
nor U4977 (N_4977,N_116,N_950);
and U4978 (N_4978,N_391,N_1187);
and U4979 (N_4979,N_1924,N_1405);
and U4980 (N_4980,N_611,N_0);
nand U4981 (N_4981,N_935,N_659);
or U4982 (N_4982,N_2478,N_355);
nand U4983 (N_4983,N_1217,N_445);
nand U4984 (N_4984,N_2267,N_1001);
xor U4985 (N_4985,N_118,N_1917);
or U4986 (N_4986,N_1885,N_2090);
or U4987 (N_4987,N_2430,N_361);
nor U4988 (N_4988,N_2188,N_559);
or U4989 (N_4989,N_2299,N_745);
nand U4990 (N_4990,N_1914,N_1875);
nor U4991 (N_4991,N_1462,N_924);
xnor U4992 (N_4992,N_683,N_2177);
nand U4993 (N_4993,N_1783,N_1042);
or U4994 (N_4994,N_2164,N_2283);
nand U4995 (N_4995,N_711,N_2031);
and U4996 (N_4996,N_728,N_1716);
or U4997 (N_4997,N_552,N_335);
nand U4998 (N_4998,N_2399,N_1540);
or U4999 (N_4999,N_598,N_1899);
and U5000 (N_5000,N_2926,N_4175);
and U5001 (N_5001,N_2554,N_4383);
and U5002 (N_5002,N_3325,N_4786);
and U5003 (N_5003,N_3867,N_3689);
and U5004 (N_5004,N_2628,N_3944);
or U5005 (N_5005,N_3139,N_4106);
xor U5006 (N_5006,N_4111,N_4589);
or U5007 (N_5007,N_3847,N_4975);
nor U5008 (N_5008,N_3853,N_2869);
and U5009 (N_5009,N_3544,N_3252);
nand U5010 (N_5010,N_3825,N_4161);
and U5011 (N_5011,N_3212,N_3426);
and U5012 (N_5012,N_4810,N_2975);
nand U5013 (N_5013,N_4882,N_4136);
or U5014 (N_5014,N_2698,N_3726);
nor U5015 (N_5015,N_3534,N_4060);
and U5016 (N_5016,N_4177,N_4283);
nand U5017 (N_5017,N_4115,N_2893);
nand U5018 (N_5018,N_4925,N_4675);
nor U5019 (N_5019,N_4313,N_4344);
nor U5020 (N_5020,N_4578,N_3064);
or U5021 (N_5021,N_4842,N_2643);
nor U5022 (N_5022,N_3894,N_2883);
nand U5023 (N_5023,N_4173,N_4054);
xor U5024 (N_5024,N_3671,N_3472);
or U5025 (N_5025,N_3257,N_2703);
nor U5026 (N_5026,N_3103,N_4889);
and U5027 (N_5027,N_4271,N_2702);
or U5028 (N_5028,N_3844,N_3326);
nand U5029 (N_5029,N_3583,N_4191);
nor U5030 (N_5030,N_4576,N_4659);
or U5031 (N_5031,N_2745,N_3943);
and U5032 (N_5032,N_3304,N_3864);
or U5033 (N_5033,N_3842,N_3204);
nand U5034 (N_5034,N_4680,N_2566);
and U5035 (N_5035,N_2856,N_3085);
nand U5036 (N_5036,N_3196,N_3210);
nand U5037 (N_5037,N_4089,N_3801);
and U5038 (N_5038,N_4284,N_4160);
nor U5039 (N_5039,N_3585,N_4204);
nor U5040 (N_5040,N_4379,N_3947);
or U5041 (N_5041,N_4276,N_4065);
and U5042 (N_5042,N_4821,N_3056);
nand U5043 (N_5043,N_2622,N_3955);
and U5044 (N_5044,N_3623,N_3399);
or U5045 (N_5045,N_3039,N_3415);
or U5046 (N_5046,N_4309,N_3497);
nand U5047 (N_5047,N_3413,N_2931);
nand U5048 (N_5048,N_2900,N_3496);
nand U5049 (N_5049,N_2736,N_4965);
nand U5050 (N_5050,N_2571,N_4755);
or U5051 (N_5051,N_4979,N_3068);
nor U5052 (N_5052,N_4792,N_3876);
nor U5053 (N_5053,N_4015,N_4042);
and U5054 (N_5054,N_3873,N_2828);
and U5055 (N_5055,N_4628,N_3023);
or U5056 (N_5056,N_2639,N_3004);
nand U5057 (N_5057,N_3438,N_3254);
nor U5058 (N_5058,N_4819,N_2667);
and U5059 (N_5059,N_4728,N_3779);
and U5060 (N_5060,N_2610,N_3348);
and U5061 (N_5061,N_3655,N_2956);
and U5062 (N_5062,N_4367,N_3140);
or U5063 (N_5063,N_2606,N_3372);
and U5064 (N_5064,N_3375,N_4021);
and U5065 (N_5065,N_3235,N_4359);
and U5066 (N_5066,N_2965,N_3150);
or U5067 (N_5067,N_4652,N_3259);
nand U5068 (N_5068,N_4326,N_4634);
or U5069 (N_5069,N_4741,N_3597);
and U5070 (N_5070,N_3333,N_2678);
nor U5071 (N_5071,N_3940,N_3117);
nand U5072 (N_5072,N_4027,N_2929);
nand U5073 (N_5073,N_3667,N_3613);
nor U5074 (N_5074,N_3697,N_4132);
nand U5075 (N_5075,N_3060,N_2930);
or U5076 (N_5076,N_3404,N_4010);
nand U5077 (N_5077,N_2857,N_3767);
and U5078 (N_5078,N_3449,N_4017);
nand U5079 (N_5079,N_4000,N_2559);
or U5080 (N_5080,N_2860,N_4079);
nand U5081 (N_5081,N_3255,N_3549);
nor U5082 (N_5082,N_4813,N_3687);
nand U5083 (N_5083,N_2699,N_3848);
or U5084 (N_5084,N_4411,N_2783);
xnor U5085 (N_5085,N_4114,N_4006);
nor U5086 (N_5086,N_4637,N_3281);
or U5087 (N_5087,N_4936,N_4227);
nand U5088 (N_5088,N_3498,N_4828);
nand U5089 (N_5089,N_4710,N_3527);
nand U5090 (N_5090,N_3939,N_2612);
nor U5091 (N_5091,N_2630,N_3546);
nor U5092 (N_5092,N_2729,N_3112);
or U5093 (N_5093,N_4881,N_3231);
or U5094 (N_5094,N_3843,N_3714);
and U5095 (N_5095,N_4030,N_2831);
or U5096 (N_5096,N_4339,N_4094);
and U5097 (N_5097,N_3475,N_4343);
nor U5098 (N_5098,N_3081,N_3615);
or U5099 (N_5099,N_4037,N_4614);
and U5100 (N_5100,N_4702,N_4389);
or U5101 (N_5101,N_4892,N_2876);
or U5102 (N_5102,N_3209,N_3719);
or U5103 (N_5103,N_3678,N_3566);
nor U5104 (N_5104,N_3849,N_3436);
nand U5105 (N_5105,N_4559,N_3759);
nor U5106 (N_5106,N_4855,N_3595);
nor U5107 (N_5107,N_3308,N_4839);
nor U5108 (N_5108,N_4214,N_4219);
nand U5109 (N_5109,N_3272,N_4534);
and U5110 (N_5110,N_3635,N_4729);
nor U5111 (N_5111,N_2598,N_3012);
nand U5112 (N_5112,N_3884,N_4513);
xnor U5113 (N_5113,N_4818,N_4325);
nand U5114 (N_5114,N_2662,N_3906);
nor U5115 (N_5115,N_4218,N_3991);
and U5116 (N_5116,N_2582,N_3818);
or U5117 (N_5117,N_2543,N_4942);
nand U5118 (N_5118,N_3479,N_3754);
and U5119 (N_5119,N_2905,N_2776);
and U5120 (N_5120,N_4645,N_4356);
nand U5121 (N_5121,N_2907,N_4186);
or U5122 (N_5122,N_3590,N_3523);
nand U5123 (N_5123,N_4905,N_3556);
nor U5124 (N_5124,N_3531,N_3402);
and U5125 (N_5125,N_2539,N_4888);
or U5126 (N_5126,N_3401,N_2726);
nor U5127 (N_5127,N_4758,N_2684);
or U5128 (N_5128,N_3875,N_4131);
and U5129 (N_5129,N_2906,N_3161);
or U5130 (N_5130,N_3238,N_4759);
and U5131 (N_5131,N_3006,N_2895);
nand U5132 (N_5132,N_3761,N_4119);
and U5133 (N_5133,N_3727,N_4725);
nand U5134 (N_5134,N_4714,N_3494);
nand U5135 (N_5135,N_3237,N_2800);
or U5136 (N_5136,N_4558,N_4328);
nand U5137 (N_5137,N_3540,N_2819);
and U5138 (N_5138,N_4629,N_4508);
and U5139 (N_5139,N_2742,N_4791);
or U5140 (N_5140,N_3770,N_2955);
nor U5141 (N_5141,N_2894,N_3747);
nand U5142 (N_5142,N_2780,N_3014);
and U5143 (N_5143,N_4803,N_4019);
nand U5144 (N_5144,N_3772,N_4996);
or U5145 (N_5145,N_3278,N_2769);
nor U5146 (N_5146,N_3820,N_4859);
and U5147 (N_5147,N_2743,N_4785);
and U5148 (N_5148,N_4701,N_4222);
nand U5149 (N_5149,N_4352,N_3493);
and U5150 (N_5150,N_3397,N_3710);
nand U5151 (N_5151,N_3920,N_4387);
and U5152 (N_5152,N_4216,N_2749);
nand U5153 (N_5153,N_2875,N_3086);
or U5154 (N_5154,N_3158,N_3422);
or U5155 (N_5155,N_4435,N_3244);
and U5156 (N_5156,N_3491,N_4621);
or U5157 (N_5157,N_4503,N_3190);
nand U5158 (N_5158,N_3838,N_3097);
nand U5159 (N_5159,N_4399,N_3587);
nand U5160 (N_5160,N_3879,N_4431);
nand U5161 (N_5161,N_4290,N_2530);
nor U5162 (N_5162,N_4931,N_4945);
or U5163 (N_5163,N_2790,N_3706);
nand U5164 (N_5164,N_4442,N_4455);
nand U5165 (N_5165,N_3358,N_4823);
nor U5166 (N_5166,N_2578,N_3594);
nor U5167 (N_5167,N_4212,N_3798);
and U5168 (N_5168,N_3685,N_3092);
nor U5169 (N_5169,N_2514,N_4670);
and U5170 (N_5170,N_4413,N_2794);
nand U5171 (N_5171,N_4564,N_3223);
nand U5172 (N_5172,N_3049,N_3808);
and U5173 (N_5173,N_4754,N_3619);
nor U5174 (N_5174,N_2944,N_3677);
and U5175 (N_5175,N_4141,N_4051);
nand U5176 (N_5176,N_2880,N_2627);
or U5177 (N_5177,N_2551,N_4949);
nor U5178 (N_5178,N_2533,N_4857);
or U5179 (N_5179,N_3020,N_4647);
nand U5180 (N_5180,N_4968,N_4631);
and U5181 (N_5181,N_4380,N_3810);
and U5182 (N_5182,N_3777,N_4928);
nor U5183 (N_5183,N_4189,N_4269);
nand U5184 (N_5184,N_4337,N_3153);
nand U5185 (N_5185,N_2933,N_4427);
or U5186 (N_5186,N_2588,N_4172);
nand U5187 (N_5187,N_4843,N_3684);
nor U5188 (N_5188,N_3447,N_4144);
and U5189 (N_5189,N_3392,N_4583);
nand U5190 (N_5190,N_2918,N_4124);
nor U5191 (N_5191,N_4028,N_3164);
or U5192 (N_5192,N_4976,N_3769);
or U5193 (N_5193,N_4993,N_3837);
xnor U5194 (N_5194,N_4310,N_3784);
or U5195 (N_5195,N_3532,N_4194);
and U5196 (N_5196,N_3990,N_3606);
and U5197 (N_5197,N_4463,N_4750);
and U5198 (N_5198,N_3709,N_3007);
nand U5199 (N_5199,N_2672,N_4672);
nand U5200 (N_5200,N_3206,N_2989);
nor U5201 (N_5201,N_4980,N_3188);
and U5202 (N_5202,N_2656,N_4777);
or U5203 (N_5203,N_4544,N_3700);
nand U5204 (N_5204,N_3050,N_3680);
nand U5205 (N_5205,N_4001,N_4814);
or U5206 (N_5206,N_2505,N_3079);
nand U5207 (N_5207,N_4994,N_4642);
or U5208 (N_5208,N_4306,N_4291);
or U5209 (N_5209,N_2567,N_3067);
nand U5210 (N_5210,N_2820,N_4409);
or U5211 (N_5211,N_3292,N_4962);
and U5212 (N_5212,N_3119,N_3854);
xnor U5213 (N_5213,N_3126,N_2990);
or U5214 (N_5214,N_3197,N_3291);
and U5215 (N_5215,N_3351,N_4904);
and U5216 (N_5216,N_4068,N_3541);
nand U5217 (N_5217,N_3013,N_3800);
nor U5218 (N_5218,N_2544,N_4987);
and U5219 (N_5219,N_3242,N_3130);
nor U5220 (N_5220,N_3312,N_4510);
nor U5221 (N_5221,N_4224,N_2710);
or U5222 (N_5222,N_2773,N_3274);
and U5223 (N_5223,N_4880,N_4587);
or U5224 (N_5224,N_4836,N_2673);
nand U5225 (N_5225,N_2771,N_4013);
and U5226 (N_5226,N_4333,N_4081);
or U5227 (N_5227,N_3214,N_3460);
and U5228 (N_5228,N_2658,N_3057);
or U5229 (N_5229,N_2679,N_4043);
nor U5230 (N_5230,N_3315,N_4527);
or U5231 (N_5231,N_3976,N_4462);
and U5232 (N_5232,N_3189,N_3768);
nor U5233 (N_5233,N_3495,N_2705);
or U5234 (N_5234,N_2635,N_3831);
and U5235 (N_5235,N_4676,N_2838);
nor U5236 (N_5236,N_4057,N_4530);
or U5237 (N_5237,N_2837,N_3025);
or U5238 (N_5238,N_3649,N_3914);
nor U5239 (N_5239,N_3478,N_4196);
nor U5240 (N_5240,N_4292,N_3696);
and U5241 (N_5241,N_3617,N_2813);
nor U5242 (N_5242,N_4529,N_3405);
and U5243 (N_5243,N_4386,N_2558);
nand U5244 (N_5244,N_3787,N_4581);
and U5245 (N_5245,N_4890,N_4778);
and U5246 (N_5246,N_3988,N_3444);
and U5247 (N_5247,N_3878,N_4384);
xor U5248 (N_5248,N_2936,N_4234);
or U5249 (N_5249,N_4388,N_3732);
nand U5250 (N_5250,N_3824,N_4466);
nor U5251 (N_5251,N_3860,N_4902);
nor U5252 (N_5252,N_3986,N_3390);
and U5253 (N_5253,N_4561,N_4850);
nor U5254 (N_5254,N_3387,N_4151);
or U5255 (N_5255,N_2862,N_3143);
or U5256 (N_5256,N_2650,N_4648);
nand U5257 (N_5257,N_3846,N_2728);
and U5258 (N_5258,N_2885,N_2802);
nand U5259 (N_5259,N_2932,N_2889);
nand U5260 (N_5260,N_2892,N_4095);
nor U5261 (N_5261,N_4126,N_3483);
and U5262 (N_5262,N_4447,N_2850);
nand U5263 (N_5263,N_3135,N_4484);
nor U5264 (N_5264,N_2943,N_4891);
nor U5265 (N_5265,N_2696,N_3224);
nor U5266 (N_5266,N_2919,N_3396);
nor U5267 (N_5267,N_3412,N_3902);
nand U5268 (N_5268,N_4341,N_4390);
nand U5269 (N_5269,N_4594,N_3945);
or U5270 (N_5270,N_3567,N_4727);
nor U5271 (N_5271,N_3071,N_4516);
nand U5272 (N_5272,N_3218,N_3341);
nand U5273 (N_5273,N_3746,N_2520);
and U5274 (N_5274,N_2793,N_4649);
and U5275 (N_5275,N_2810,N_4147);
xor U5276 (N_5276,N_4963,N_2879);
nor U5277 (N_5277,N_3423,N_3155);
nand U5278 (N_5278,N_3877,N_2952);
nand U5279 (N_5279,N_4319,N_4560);
and U5280 (N_5280,N_4860,N_3248);
or U5281 (N_5281,N_3822,N_4619);
or U5282 (N_5282,N_2806,N_4489);
or U5283 (N_5283,N_4229,N_2519);
or U5284 (N_5284,N_2980,N_3264);
or U5285 (N_5285,N_2941,N_3699);
nor U5286 (N_5286,N_3486,N_4206);
and U5287 (N_5287,N_3339,N_4789);
nand U5288 (N_5288,N_4375,N_4154);
nand U5289 (N_5289,N_4443,N_3120);
or U5290 (N_5290,N_4166,N_4526);
and U5291 (N_5291,N_2546,N_3167);
and U5292 (N_5292,N_2945,N_3336);
nor U5293 (N_5293,N_3323,N_4072);
or U5294 (N_5294,N_4723,N_4123);
xnor U5295 (N_5295,N_3031,N_4113);
nor U5296 (N_5296,N_4597,N_3037);
and U5297 (N_5297,N_2508,N_4591);
nor U5298 (N_5298,N_2823,N_3658);
and U5299 (N_5299,N_3106,N_4116);
and U5300 (N_5300,N_2787,N_3428);
or U5301 (N_5301,N_3251,N_3954);
nand U5302 (N_5302,N_4139,N_2704);
and U5303 (N_5303,N_2604,N_3434);
nand U5304 (N_5304,N_4008,N_2642);
and U5305 (N_5305,N_3736,N_4677);
nor U5306 (N_5306,N_4432,N_3192);
nand U5307 (N_5307,N_4615,N_4300);
or U5308 (N_5308,N_2881,N_2506);
or U5309 (N_5309,N_3017,N_2739);
nor U5310 (N_5310,N_4428,N_3221);
and U5311 (N_5311,N_2765,N_3895);
nand U5312 (N_5312,N_3324,N_3601);
and U5313 (N_5313,N_3885,N_3528);
or U5314 (N_5314,N_4549,N_4253);
and U5315 (N_5315,N_4417,N_2763);
and U5316 (N_5316,N_3195,N_4694);
nor U5317 (N_5317,N_3187,N_2865);
or U5318 (N_5318,N_2963,N_4209);
xnor U5319 (N_5319,N_3724,N_3273);
nor U5320 (N_5320,N_4509,N_2999);
and U5321 (N_5321,N_4125,N_4520);
nor U5322 (N_5322,N_2573,N_2518);
or U5323 (N_5323,N_4033,N_4371);
or U5324 (N_5324,N_3880,N_4596);
xnor U5325 (N_5325,N_4248,N_4408);
nor U5326 (N_5326,N_4854,N_3015);
or U5327 (N_5327,N_4764,N_4215);
or U5328 (N_5328,N_2966,N_3668);
nand U5329 (N_5329,N_3510,N_3216);
and U5330 (N_5330,N_3384,N_3100);
nor U5331 (N_5331,N_3931,N_3113);
or U5332 (N_5332,N_3370,N_3917);
or U5333 (N_5333,N_4316,N_3116);
nand U5334 (N_5334,N_3427,N_3430);
nor U5335 (N_5335,N_4268,N_3804);
nand U5336 (N_5336,N_4971,N_4988);
nand U5337 (N_5337,N_3124,N_3950);
nor U5338 (N_5338,N_3215,N_3773);
xor U5339 (N_5339,N_4236,N_2803);
nor U5340 (N_5340,N_4689,N_3461);
or U5341 (N_5341,N_3547,N_3579);
and U5342 (N_5342,N_3425,N_3589);
nand U5343 (N_5343,N_3271,N_2830);
or U5344 (N_5344,N_4293,N_4546);
nand U5345 (N_5345,N_4127,N_4301);
nand U5346 (N_5346,N_4226,N_3093);
and U5347 (N_5347,N_3865,N_4012);
nand U5348 (N_5348,N_3347,N_4536);
or U5349 (N_5349,N_2910,N_2951);
and U5350 (N_5350,N_3887,N_4270);
or U5351 (N_5351,N_4239,N_3698);
nor U5352 (N_5352,N_2560,N_4448);
and U5353 (N_5353,N_3035,N_2576);
nand U5354 (N_5354,N_4769,N_3090);
nand U5355 (N_5355,N_4586,N_4872);
or U5356 (N_5356,N_3753,N_3815);
nand U5357 (N_5357,N_3536,N_4972);
and U5358 (N_5358,N_2607,N_4217);
nor U5359 (N_5359,N_3077,N_3382);
or U5360 (N_5360,N_4364,N_2624);
nand U5361 (N_5361,N_3319,N_4070);
xor U5362 (N_5362,N_4743,N_3075);
nor U5363 (N_5363,N_2674,N_4871);
and U5364 (N_5364,N_4721,N_3355);
and U5365 (N_5365,N_3171,N_4726);
or U5366 (N_5366,N_3136,N_3764);
nand U5367 (N_5367,N_4278,N_4656);
xor U5368 (N_5368,N_3276,N_2561);
nor U5369 (N_5369,N_4492,N_3095);
nand U5370 (N_5370,N_3733,N_4009);
nand U5371 (N_5371,N_3518,N_2600);
and U5372 (N_5372,N_3938,N_2616);
or U5373 (N_5373,N_3421,N_2614);
and U5374 (N_5374,N_4610,N_2748);
xor U5375 (N_5375,N_4922,N_3925);
nor U5376 (N_5376,N_3279,N_4137);
or U5377 (N_5377,N_4285,N_2653);
nand U5378 (N_5378,N_4308,N_2912);
and U5379 (N_5379,N_3984,N_4109);
and U5380 (N_5380,N_3640,N_4868);
nand U5381 (N_5381,N_4961,N_4099);
and U5382 (N_5382,N_2882,N_4152);
nand U5383 (N_5383,N_4445,N_4496);
nor U5384 (N_5384,N_3408,N_3855);
or U5385 (N_5385,N_4201,N_3132);
and U5386 (N_5386,N_4307,N_4471);
and U5387 (N_5387,N_3612,N_4487);
or U5388 (N_5388,N_2870,N_3448);
nor U5389 (N_5389,N_4391,N_2503);
and U5390 (N_5390,N_4956,N_3376);
nand U5391 (N_5391,N_4523,N_4895);
xnor U5392 (N_5392,N_3839,N_4883);
or U5393 (N_5393,N_4967,N_3561);
nor U5394 (N_5394,N_3501,N_4372);
and U5395 (N_5395,N_4446,N_3780);
nand U5396 (N_5396,N_3829,N_3476);
or U5397 (N_5397,N_4440,N_3563);
nand U5398 (N_5398,N_4749,N_4335);
nor U5399 (N_5399,N_4479,N_3835);
and U5400 (N_5400,N_3998,N_3702);
or U5401 (N_5401,N_3234,N_4575);
or U5402 (N_5402,N_4362,N_3827);
nand U5403 (N_5403,N_4260,N_4877);
or U5404 (N_5404,N_4497,N_3748);
nor U5405 (N_5405,N_4437,N_4745);
nand U5406 (N_5406,N_2608,N_2564);
nor U5407 (N_5407,N_2834,N_3091);
and U5408 (N_5408,N_4995,N_3073);
nand U5409 (N_5409,N_3972,N_4704);
or U5410 (N_5410,N_2785,N_4198);
nor U5411 (N_5411,N_2997,N_2996);
nand U5412 (N_5412,N_4368,N_4184);
xor U5413 (N_5413,N_2751,N_4910);
or U5414 (N_5414,N_3352,N_4453);
nand U5415 (N_5415,N_3146,N_3651);
nand U5416 (N_5416,N_3181,N_4524);
and U5417 (N_5417,N_4679,N_4932);
nor U5418 (N_5418,N_2647,N_2593);
and U5419 (N_5419,N_3809,N_4712);
or U5420 (N_5420,N_4064,N_3836);
nand U5421 (N_5421,N_3788,N_4318);
nor U5422 (N_5422,N_4552,N_2701);
nor U5423 (N_5423,N_3555,N_2632);
nand U5424 (N_5424,N_2676,N_3716);
nand U5425 (N_5425,N_3052,N_2871);
and U5426 (N_5426,N_3394,N_2690);
or U5427 (N_5427,N_4174,N_4235);
or U5428 (N_5428,N_2994,N_2967);
and U5429 (N_5429,N_3058,N_4545);
or U5430 (N_5430,N_3647,N_4709);
xnor U5431 (N_5431,N_2959,N_4632);
nand U5432 (N_5432,N_4288,N_4066);
nand U5433 (N_5433,N_4024,N_4879);
nor U5434 (N_5434,N_3128,N_4858);
xor U5435 (N_5435,N_3785,N_4566);
nand U5436 (N_5436,N_2580,N_2511);
nor U5437 (N_5437,N_2948,N_3080);
or U5438 (N_5438,N_3817,N_4303);
and U5439 (N_5439,N_4381,N_4840);
nand U5440 (N_5440,N_4122,N_4921);
or U5441 (N_5441,N_3907,N_3138);
and U5442 (N_5442,N_3662,N_3573);
nor U5443 (N_5443,N_4103,N_2526);
or U5444 (N_5444,N_4180,N_4277);
nor U5445 (N_5445,N_3713,N_4767);
nor U5446 (N_5446,N_2623,N_3318);
nand U5447 (N_5447,N_4415,N_4007);
and U5448 (N_5448,N_3965,N_3265);
nor U5449 (N_5449,N_2740,N_3163);
or U5450 (N_5450,N_3165,N_3638);
and U5451 (N_5451,N_3560,N_2599);
or U5452 (N_5452,N_3929,N_4346);
nor U5453 (N_5453,N_4167,N_4711);
nor U5454 (N_5454,N_4869,N_3608);
nor U5455 (N_5455,N_4220,N_3949);
and U5456 (N_5456,N_3888,N_2528);
and U5457 (N_5457,N_3270,N_4535);
and U5458 (N_5458,N_4469,N_3040);
and U5459 (N_5459,N_2849,N_4203);
nor U5460 (N_5460,N_4938,N_4294);
or U5461 (N_5461,N_3369,N_3470);
and U5462 (N_5462,N_2553,N_2922);
xnor U5463 (N_5463,N_3115,N_2960);
or U5464 (N_5464,N_3942,N_4686);
or U5465 (N_5465,N_3791,N_3314);
or U5466 (N_5466,N_4329,N_3280);
and U5467 (N_5467,N_3366,N_2847);
and U5468 (N_5468,N_4193,N_3870);
nand U5469 (N_5469,N_4422,N_2808);
and U5470 (N_5470,N_3708,N_3858);
or U5471 (N_5471,N_2515,N_3852);
nor U5472 (N_5472,N_3028,N_3591);
nor U5473 (N_5473,N_4402,N_4826);
nor U5474 (N_5474,N_4385,N_2668);
and U5475 (N_5475,N_3360,N_3042);
and U5476 (N_5476,N_2646,N_3695);
or U5477 (N_5477,N_4838,N_3203);
and U5478 (N_5478,N_4360,N_2845);
or U5479 (N_5479,N_3686,N_3863);
and U5480 (N_5480,N_3123,N_3592);
or U5481 (N_5481,N_4423,N_4110);
or U5482 (N_5482,N_3900,N_3286);
nand U5483 (N_5483,N_3760,N_2523);
nand U5484 (N_5484,N_2886,N_4678);
nand U5485 (N_5485,N_4772,N_3750);
and U5486 (N_5486,N_4851,N_4093);
or U5487 (N_5487,N_3922,N_4475);
and U5488 (N_5488,N_4358,N_3099);
and U5489 (N_5489,N_3811,N_2782);
nand U5490 (N_5490,N_4092,N_3602);
nor U5491 (N_5491,N_3230,N_4719);
or U5492 (N_5492,N_3356,N_3469);
or U5493 (N_5493,N_3083,N_4311);
nand U5494 (N_5494,N_3180,N_4580);
nand U5495 (N_5495,N_3946,N_3346);
or U5496 (N_5496,N_4816,N_2902);
nor U5497 (N_5497,N_4481,N_4722);
or U5498 (N_5498,N_4638,N_3681);
and U5499 (N_5499,N_3416,N_3634);
or U5500 (N_5500,N_3841,N_2545);
or U5501 (N_5501,N_3633,N_4603);
nor U5502 (N_5502,N_2770,N_3969);
and U5503 (N_5503,N_3373,N_4003);
and U5504 (N_5504,N_4584,N_4718);
nor U5505 (N_5505,N_2709,N_4188);
xnor U5506 (N_5506,N_4538,N_2618);
or U5507 (N_5507,N_3033,N_4739);
and U5508 (N_5508,N_3474,N_3503);
xnor U5509 (N_5509,N_4504,N_3144);
nor U5510 (N_5510,N_3407,N_3309);
and U5511 (N_5511,N_3311,N_3047);
nand U5512 (N_5512,N_3285,N_3982);
or U5513 (N_5513,N_2711,N_4230);
nand U5514 (N_5514,N_4289,N_4327);
and U5515 (N_5515,N_4480,N_2500);
nand U5516 (N_5516,N_3284,N_4623);
or U5517 (N_5517,N_3539,N_4083);
and U5518 (N_5518,N_4062,N_4863);
and U5519 (N_5519,N_4740,N_4460);
xnor U5520 (N_5520,N_3320,N_3928);
and U5521 (N_5521,N_4644,N_2877);
nand U5522 (N_5522,N_4178,N_2715);
or U5523 (N_5523,N_4022,N_4138);
nor U5524 (N_5524,N_4334,N_2985);
and U5525 (N_5525,N_2961,N_3997);
nor U5526 (N_5526,N_2677,N_3987);
or U5527 (N_5527,N_2693,N_2651);
and U5528 (N_5528,N_4195,N_2654);
nor U5529 (N_5529,N_4815,N_4747);
or U5530 (N_5530,N_4071,N_3513);
or U5531 (N_5531,N_4627,N_4695);
nor U5532 (N_5532,N_2818,N_3022);
or U5533 (N_5533,N_2764,N_4543);
nor U5534 (N_5534,N_2501,N_3786);
or U5535 (N_5535,N_4133,N_3909);
or U5536 (N_5536,N_2937,N_3456);
and U5537 (N_5537,N_3066,N_2868);
and U5538 (N_5538,N_3983,N_3652);
nor U5539 (N_5539,N_4420,N_4715);
nor U5540 (N_5540,N_3419,N_2781);
nand U5541 (N_5541,N_3443,N_3548);
or U5542 (N_5542,N_3564,N_4811);
nor U5543 (N_5543,N_4698,N_4511);
and U5544 (N_5544,N_2611,N_4425);
and U5545 (N_5545,N_2666,N_3962);
nand U5546 (N_5546,N_2664,N_4493);
nor U5547 (N_5547,N_3641,N_4599);
nor U5548 (N_5548,N_2947,N_3996);
or U5549 (N_5549,N_3675,N_3883);
nor U5550 (N_5550,N_4087,N_3310);
nand U5551 (N_5551,N_4342,N_3065);
or U5552 (N_5552,N_4550,N_2669);
nor U5553 (N_5553,N_4713,N_4588);
and U5554 (N_5554,N_4595,N_4799);
and U5555 (N_5555,N_3582,N_3168);
or U5556 (N_5556,N_3463,N_3505);
or U5557 (N_5557,N_3749,N_3871);
nand U5558 (N_5558,N_3912,N_3213);
or U5559 (N_5559,N_3256,N_3802);
nand U5560 (N_5560,N_4029,N_2852);
and U5561 (N_5561,N_4050,N_4756);
nor U5562 (N_5562,N_2940,N_4395);
nor U5563 (N_5563,N_4901,N_2649);
nand U5564 (N_5564,N_4917,N_2707);
or U5565 (N_5565,N_3952,N_3201);
nand U5566 (N_5566,N_4746,N_4039);
or U5567 (N_5567,N_2942,N_4795);
nand U5568 (N_5568,N_3796,N_3266);
nand U5569 (N_5569,N_4716,N_3923);
or U5570 (N_5570,N_3530,N_4512);
nor U5571 (N_5571,N_4914,N_4404);
xor U5572 (N_5572,N_3936,N_4494);
nand U5573 (N_5573,N_4477,N_4783);
and U5574 (N_5574,N_4419,N_2510);
nand U5575 (N_5575,N_4732,N_3845);
and U5576 (N_5576,N_4822,N_4034);
nor U5577 (N_5577,N_3519,N_3473);
nor U5578 (N_5578,N_3395,N_2786);
nand U5579 (N_5579,N_3104,N_4086);
and U5580 (N_5580,N_3711,N_3391);
nand U5581 (N_5581,N_3026,N_4102);
nor U5582 (N_5582,N_3935,N_4554);
nand U5583 (N_5583,N_4059,N_3797);
nor U5584 (N_5584,N_3956,N_2671);
xor U5585 (N_5585,N_3765,N_2824);
nor U5586 (N_5586,N_3169,N_3621);
and U5587 (N_5587,N_2805,N_4365);
or U5588 (N_5588,N_4556,N_3993);
xnor U5589 (N_5589,N_3293,N_2538);
and U5590 (N_5590,N_2601,N_3908);
and U5591 (N_5591,N_2502,N_3964);
nand U5592 (N_5592,N_3559,N_3137);
nor U5593 (N_5593,N_3913,N_4969);
nor U5594 (N_5594,N_3045,N_3737);
or U5595 (N_5595,N_3620,N_2688);
nand U5596 (N_5596,N_4286,N_4129);
and U5597 (N_5597,N_3850,N_4374);
and U5598 (N_5598,N_2574,N_3490);
or U5599 (N_5599,N_2755,N_3666);
nor U5600 (N_5600,N_3961,N_4369);
nor U5601 (N_5601,N_3317,N_4183);
or U5602 (N_5602,N_3512,N_3330);
or U5603 (N_5603,N_4005,N_3905);
nand U5604 (N_5604,N_3364,N_4495);
or U5605 (N_5605,N_2998,N_3899);
nand U5606 (N_5606,N_4958,N_3061);
and U5607 (N_5607,N_2884,N_2691);
or U5608 (N_5608,N_4941,N_4458);
and U5609 (N_5609,N_3432,N_4320);
nor U5610 (N_5610,N_3268,N_4893);
or U5611 (N_5611,N_4221,N_3618);
or U5612 (N_5612,N_4846,N_4911);
or U5613 (N_5613,N_2858,N_4955);
nand U5614 (N_5614,N_3565,N_3290);
and U5615 (N_5615,N_4848,N_4997);
nand U5616 (N_5616,N_2953,N_2851);
nand U5617 (N_5617,N_2934,N_3869);
nand U5618 (N_5618,N_4082,N_3721);
nand U5619 (N_5619,N_3492,N_4620);
nand U5620 (N_5620,N_3792,N_3411);
nand U5621 (N_5621,N_3645,N_3414);
nand U5622 (N_5622,N_4242,N_2717);
or U5623 (N_5623,N_2957,N_3584);
and U5624 (N_5624,N_3823,N_4964);
nor U5625 (N_5625,N_4787,N_2887);
and U5626 (N_5626,N_4498,N_3970);
and U5627 (N_5627,N_3776,N_3166);
and U5628 (N_5628,N_2602,N_3889);
nor U5629 (N_5629,N_3400,N_2836);
and U5630 (N_5630,N_2814,N_4240);
nor U5631 (N_5631,N_4681,N_3628);
nand U5632 (N_5632,N_2759,N_3298);
nor U5633 (N_5633,N_4537,N_4806);
and U5634 (N_5634,N_4055,N_3593);
nand U5635 (N_5635,N_4067,N_2822);
nand U5636 (N_5636,N_3451,N_2788);
nand U5637 (N_5637,N_3806,N_4401);
nand U5638 (N_5638,N_3217,N_3705);
nand U5639 (N_5639,N_3134,N_3378);
nand U5640 (N_5640,N_4250,N_4225);
nand U5641 (N_5641,N_3533,N_2631);
or U5642 (N_5642,N_4622,N_3643);
and U5643 (N_5643,N_4668,N_3198);
and U5644 (N_5644,N_3979,N_2692);
xnor U5645 (N_5645,N_2716,N_4377);
nand U5646 (N_5646,N_3739,N_4258);
or U5647 (N_5647,N_3874,N_4244);
and U5648 (N_5648,N_3890,N_4633);
or U5649 (N_5649,N_4096,N_3799);
nor U5650 (N_5650,N_3703,N_4332);
or U5651 (N_5651,N_2577,N_3377);
nor U5652 (N_5652,N_4461,N_4939);
nand U5653 (N_5653,N_4354,N_4870);
or U5654 (N_5654,N_4906,N_3131);
and U5655 (N_5655,N_2752,N_2565);
nor U5656 (N_5656,N_4797,N_3814);
nand U5657 (N_5657,N_2853,N_3866);
nor U5658 (N_5658,N_4439,N_4370);
or U5659 (N_5659,N_3043,N_4145);
and U5660 (N_5660,N_2970,N_3420);
nand U5661 (N_5661,N_4100,N_4582);
nor U5662 (N_5662,N_3568,N_4153);
or U5663 (N_5663,N_4565,N_2562);
and U5664 (N_5664,N_3245,N_4837);
nand U5665 (N_5665,N_4827,N_4674);
or U5666 (N_5666,N_4363,N_3322);
nand U5667 (N_5667,N_3160,N_2841);
nor U5668 (N_5668,N_4041,N_4366);
nor U5669 (N_5669,N_3239,N_3000);
nand U5670 (N_5670,N_3431,N_3669);
and U5671 (N_5671,N_3967,N_2556);
nand U5672 (N_5672,N_3228,N_4085);
nor U5673 (N_5673,N_2584,N_2744);
nand U5674 (N_5674,N_2552,N_4148);
nor U5675 (N_5675,N_3926,N_2792);
or U5676 (N_5676,N_2914,N_4687);
or U5677 (N_5677,N_4165,N_4563);
or U5678 (N_5678,N_3030,N_3639);
and U5679 (N_5679,N_3915,N_4651);
nand U5680 (N_5680,N_2640,N_4540);
or U5681 (N_5681,N_4667,N_3794);
or U5682 (N_5682,N_3287,N_3771);
nor U5683 (N_5683,N_4456,N_2978);
nand U5684 (N_5684,N_3762,N_3622);
nand U5685 (N_5685,N_4982,N_4765);
nand U5686 (N_5686,N_3344,N_3283);
nand U5687 (N_5687,N_3636,N_3715);
or U5688 (N_5688,N_4832,N_4078);
nand U5689 (N_5689,N_4555,N_2904);
nand U5690 (N_5690,N_3805,N_3793);
and U5691 (N_5691,N_2591,N_4407);
nand U5692 (N_5692,N_3019,N_4616);
or U5693 (N_5693,N_3220,N_4809);
nand U5694 (N_5694,N_2784,N_3054);
and U5695 (N_5695,N_3380,N_2550);
nor U5696 (N_5696,N_4989,N_2540);
nor U5697 (N_5697,N_3087,N_3409);
nand U5698 (N_5698,N_4817,N_2652);
nor U5699 (N_5699,N_4532,N_2921);
or U5700 (N_5700,N_3735,N_4025);
nor U5701 (N_5701,N_3442,N_3515);
nor U5702 (N_5702,N_3299,N_4593);
and U5703 (N_5703,N_2757,N_4052);
nand U5704 (N_5704,N_4521,N_4673);
or U5705 (N_5705,N_4170,N_4211);
nor U5706 (N_5706,N_3653,N_2768);
or U5707 (N_5707,N_3893,N_2899);
nor U5708 (N_5708,N_2722,N_4002);
or U5709 (N_5709,N_3226,N_3362);
or U5710 (N_5710,N_3371,N_4467);
nand U5711 (N_5711,N_4053,N_4853);
or U5712 (N_5712,N_4541,N_4393);
nand U5713 (N_5713,N_4742,N_4405);
and U5714 (N_5714,N_4522,N_4579);
or U5715 (N_5715,N_2909,N_4473);
and U5716 (N_5716,N_3755,N_4084);
nor U5717 (N_5717,N_4699,N_4011);
nor U5718 (N_5718,N_4903,N_3300);
or U5719 (N_5719,N_2542,N_4261);
nand U5720 (N_5720,N_3386,N_4465);
nand U5721 (N_5721,N_4098,N_4187);
or U5722 (N_5722,N_3648,N_2586);
or U5723 (N_5723,N_4149,N_2670);
nand U5724 (N_5724,N_4773,N_4424);
nand U5725 (N_5725,N_4483,N_3142);
nand U5726 (N_5726,N_2758,N_4760);
or U5727 (N_5727,N_4200,N_4533);
nand U5728 (N_5728,N_4434,N_2714);
nand U5729 (N_5729,N_4373,N_3159);
or U5730 (N_5730,N_3157,N_3807);
and U5731 (N_5731,N_4977,N_4805);
or U5732 (N_5732,N_4252,N_4899);
nand U5733 (N_5733,N_2891,N_3538);
and U5734 (N_5734,N_3588,N_4952);
nand U5735 (N_5735,N_3021,N_3741);
and U5736 (N_5736,N_4801,N_4074);
nand U5737 (N_5737,N_3118,N_4990);
xnor U5738 (N_5738,N_4948,N_2825);
nor U5739 (N_5739,N_3101,N_3712);
or U5740 (N_5740,N_4592,N_3891);
or U5741 (N_5741,N_2585,N_4018);
nand U5742 (N_5742,N_3379,N_2986);
or U5743 (N_5743,N_3663,N_4751);
xnor U5744 (N_5744,N_2982,N_3828);
and U5745 (N_5745,N_4800,N_3029);
xor U5746 (N_5746,N_4047,N_3529);
or U5747 (N_5747,N_4763,N_3577);
and U5748 (N_5748,N_2621,N_2863);
nor U5749 (N_5749,N_3172,N_2829);
nor U5750 (N_5750,N_2839,N_4831);
or U5751 (N_5751,N_2681,N_4076);
nor U5752 (N_5752,N_4159,N_4357);
nand U5753 (N_5753,N_4429,N_3783);
or U5754 (N_5754,N_2516,N_4752);
nand U5755 (N_5755,N_4761,N_3176);
or U5756 (N_5756,N_4876,N_2572);
and U5757 (N_5757,N_2817,N_2594);
and U5758 (N_5758,N_3610,N_3338);
nor U5759 (N_5759,N_4661,N_3657);
nand U5760 (N_5760,N_3516,N_2916);
nor U5761 (N_5761,N_3034,N_2655);
nor U5762 (N_5762,N_4397,N_4951);
nor U5763 (N_5763,N_2747,N_2644);
xnor U5764 (N_5764,N_3282,N_4981);
nand U5765 (N_5765,N_4197,N_4950);
and U5766 (N_5766,N_4738,N_4426);
nand U5767 (N_5767,N_3367,N_3693);
and U5768 (N_5768,N_3477,N_3114);
or U5769 (N_5769,N_3125,N_4213);
nor U5770 (N_5770,N_4608,N_4724);
nor U5771 (N_5771,N_4478,N_3892);
and U5772 (N_5772,N_4682,N_3916);
or U5773 (N_5773,N_3148,N_2797);
or U5774 (N_5774,N_3403,N_2746);
nand U5775 (N_5775,N_3349,N_2971);
or U5776 (N_5776,N_3183,N_2779);
or U5777 (N_5777,N_2821,N_4782);
nand U5778 (N_5778,N_4336,N_2816);
and U5779 (N_5779,N_3999,N_4692);
nand U5780 (N_5780,N_3520,N_4451);
and U5781 (N_5781,N_4158,N_3459);
and U5782 (N_5782,N_3331,N_4243);
and U5783 (N_5783,N_4457,N_3757);
nor U5784 (N_5784,N_2827,N_3297);
nor U5785 (N_5785,N_3694,N_4654);
nor U5786 (N_5786,N_3948,N_4302);
and U5787 (N_5787,N_4345,N_2753);
nor U5788 (N_5788,N_3236,N_4697);
and U5789 (N_5789,N_2958,N_4049);
nor U5790 (N_5790,N_4032,N_3233);
nor U5791 (N_5791,N_4474,N_4983);
nand U5792 (N_5792,N_4528,N_3327);
nor U5793 (N_5793,N_2527,N_3162);
or U5794 (N_5794,N_2974,N_4574);
nand U5795 (N_5795,N_3243,N_2723);
nor U5796 (N_5796,N_3661,N_4835);
nand U5797 (N_5797,N_3464,N_3343);
nor U5798 (N_5798,N_3637,N_3574);
nand U5799 (N_5799,N_4097,N_3055);
or U5800 (N_5800,N_3193,N_3173);
nand U5801 (N_5801,N_4257,N_4490);
and U5802 (N_5802,N_3289,N_3729);
or U5803 (N_5803,N_3522,N_4666);
or U5804 (N_5804,N_2762,N_2568);
and U5805 (N_5805,N_2920,N_3614);
nor U5806 (N_5806,N_3790,N_4824);
xnor U5807 (N_5807,N_3725,N_3959);
or U5808 (N_5808,N_4693,N_4794);
and U5809 (N_5809,N_4607,N_3084);
and U5810 (N_5810,N_3457,N_4600);
nand U5811 (N_5811,N_3455,N_2925);
and U5812 (N_5812,N_3604,N_2605);
or U5813 (N_5813,N_4245,N_3525);
xor U5814 (N_5814,N_2991,N_4943);
and U5815 (N_5815,N_4612,N_2617);
nand U5816 (N_5816,N_2626,N_4350);
nor U5817 (N_5817,N_3435,N_4768);
and U5818 (N_5818,N_3345,N_3506);
or U5819 (N_5819,N_3521,N_4829);
and U5820 (N_5820,N_3313,N_3051);
nor U5821 (N_5821,N_4886,N_3078);
nand U5822 (N_5822,N_4421,N_3429);
or U5823 (N_5823,N_4091,N_4798);
or U5824 (N_5824,N_2968,N_4878);
or U5825 (N_5825,N_3774,N_4412);
nor U5826 (N_5826,N_2992,N_3968);
or U5827 (N_5827,N_4731,N_4205);
nor U5828 (N_5828,N_4472,N_4757);
nor U5829 (N_5829,N_4924,N_3417);
and U5830 (N_5830,N_3507,N_2583);
or U5831 (N_5831,N_3978,N_2659);
nand U5832 (N_5832,N_3334,N_4601);
and U5833 (N_5833,N_4897,N_3896);
nor U5834 (N_5834,N_3263,N_3354);
nor U5835 (N_5835,N_2719,N_2778);
and U5836 (N_5836,N_2799,N_3337);
xnor U5837 (N_5837,N_4105,N_2927);
nand U5838 (N_5838,N_4992,N_4459);
nand U5839 (N_5839,N_2609,N_3720);
nand U5840 (N_5840,N_2804,N_3288);
nand U5841 (N_5841,N_3751,N_3151);
nor U5842 (N_5842,N_4351,N_4862);
or U5843 (N_5843,N_4775,N_3763);
or U5844 (N_5844,N_4266,N_4918);
and U5845 (N_5845,N_3819,N_3886);
or U5846 (N_5846,N_4488,N_4331);
or U5847 (N_5847,N_4444,N_4812);
or U5848 (N_5848,N_2682,N_4040);
xnor U5849 (N_5849,N_4322,N_3552);
nand U5850 (N_5850,N_4430,N_3048);
and U5851 (N_5851,N_4887,N_4916);
and U5852 (N_5852,N_4120,N_4705);
nand U5853 (N_5853,N_2735,N_4830);
and U5854 (N_5854,N_4577,N_3296);
or U5855 (N_5855,N_3191,N_4403);
nor U5856 (N_5856,N_4023,N_4080);
nor U5857 (N_5857,N_4920,N_3170);
nand U5858 (N_5858,N_4121,N_4232);
or U5859 (N_5859,N_2911,N_3570);
or U5860 (N_5860,N_3781,N_3670);
or U5861 (N_5861,N_3062,N_4088);
or U5862 (N_5862,N_4491,N_4650);
and U5863 (N_5863,N_4653,N_4118);
nand U5864 (N_5864,N_4181,N_4016);
nor U5865 (N_5865,N_4700,N_3966);
nor U5866 (N_5866,N_2570,N_3005);
or U5867 (N_5867,N_3467,N_3960);
nor U5868 (N_5868,N_2812,N_3149);
nand U5869 (N_5869,N_3660,N_3207);
nor U5870 (N_5870,N_2939,N_2809);
or U5871 (N_5871,N_3795,N_2737);
nand U5872 (N_5872,N_4077,N_3572);
or U5873 (N_5873,N_3665,N_4048);
nor U5874 (N_5874,N_3389,N_2525);
nor U5875 (N_5875,N_3003,N_4609);
nor U5876 (N_5876,N_4793,N_3277);
nand U5877 (N_5877,N_2620,N_4784);
and U5878 (N_5878,N_4531,N_3742);
or U5879 (N_5879,N_3691,N_3937);
xnor U5880 (N_5880,N_3446,N_4323);
and U5881 (N_5881,N_4338,N_2615);
or U5882 (N_5882,N_3267,N_4199);
or U5883 (N_5883,N_4636,N_4753);
nor U5884 (N_5884,N_2867,N_2859);
and U5885 (N_5885,N_3227,N_3098);
nand U5886 (N_5886,N_3307,N_3335);
nand U5887 (N_5887,N_4960,N_3607);
nand U5888 (N_5888,N_4696,N_3738);
nand U5889 (N_5889,N_4135,N_4263);
and U5890 (N_5890,N_2694,N_3656);
nor U5891 (N_5891,N_4542,N_3241);
and U5892 (N_5892,N_2772,N_2720);
nor U5893 (N_5893,N_3951,N_3826);
and U5894 (N_5894,N_3901,N_2854);
or U5895 (N_5895,N_3232,N_4376);
xnor U5896 (N_5896,N_4735,N_3105);
nor U5897 (N_5897,N_4450,N_3328);
xnor U5898 (N_5898,N_4073,N_4590);
nor U5899 (N_5899,N_4433,N_4884);
and U5900 (N_5900,N_3069,N_2724);
or U5901 (N_5901,N_4296,N_2555);
nand U5902 (N_5902,N_4247,N_2807);
and U5903 (N_5903,N_3517,N_4282);
nand U5904 (N_5904,N_2897,N_2924);
or U5905 (N_5905,N_4984,N_3924);
and U5906 (N_5906,N_4568,N_3575);
nor U5907 (N_5907,N_3911,N_4279);
and U5908 (N_5908,N_3365,N_4382);
and U5909 (N_5909,N_4298,N_4690);
or U5910 (N_5910,N_3406,N_2861);
nand U5911 (N_5911,N_3973,N_4361);
nand U5912 (N_5912,N_4970,N_3758);
nor U5913 (N_5913,N_4557,N_3046);
nand U5914 (N_5914,N_3557,N_3717);
nor U5915 (N_5915,N_3089,N_2532);
xor U5916 (N_5916,N_2791,N_3654);
xor U5917 (N_5917,N_3745,N_4254);
nor U5918 (N_5918,N_2675,N_4507);
nand U5919 (N_5919,N_2522,N_2795);
or U5920 (N_5920,N_4171,N_3631);
and U5921 (N_5921,N_4436,N_3219);
xnor U5922 (N_5922,N_2521,N_3963);
and U5923 (N_5923,N_2928,N_3778);
nor U5924 (N_5924,N_4834,N_3109);
nor U5925 (N_5925,N_3932,N_3357);
nand U5926 (N_5926,N_3205,N_4182);
nor U5927 (N_5927,N_3526,N_4305);
nor U5928 (N_5928,N_4685,N_4207);
and U5929 (N_5929,N_2509,N_2513);
or U5930 (N_5930,N_3175,N_3471);
nand U5931 (N_5931,N_4915,N_3301);
nor U5932 (N_5932,N_4978,N_3179);
or U5933 (N_5933,N_3186,N_3624);
nand U5934 (N_5934,N_2733,N_2625);
nand U5935 (N_5935,N_3578,N_4185);
or U5936 (N_5936,N_4671,N_4449);
xor U5937 (N_5937,N_3868,N_3342);
nand U5938 (N_5938,N_4355,N_3044);
and U5939 (N_5939,N_4625,N_4957);
or U5940 (N_5940,N_2756,N_2547);
or U5941 (N_5941,N_4169,N_4392);
or U5942 (N_5942,N_3605,N_3260);
nand U5943 (N_5943,N_4312,N_3974);
nor U5944 (N_5944,N_3229,N_4155);
and U5945 (N_5945,N_4163,N_3141);
nand U5946 (N_5946,N_3683,N_4844);
and U5947 (N_5947,N_2846,N_3789);
and U5948 (N_5948,N_3630,N_4069);
nand U5949 (N_5949,N_4396,N_4340);
or U5950 (N_5950,N_3812,N_4874);
nor U5951 (N_5951,N_3452,N_4944);
or U5952 (N_5952,N_4688,N_3921);
or U5953 (N_5953,N_3861,N_4157);
nand U5954 (N_5954,N_3194,N_4506);
or U5955 (N_5955,N_2713,N_3018);
or U5956 (N_5956,N_4233,N_3642);
nand U5957 (N_5957,N_2833,N_3743);
and U5958 (N_5958,N_2563,N_3011);
nand U5959 (N_5959,N_4611,N_4605);
nand U5960 (N_5960,N_2766,N_2706);
nor U5961 (N_5961,N_4748,N_4825);
and U5962 (N_5962,N_3250,N_4861);
or U5963 (N_5963,N_4999,N_4210);
nand U5964 (N_5964,N_4849,N_4031);
xor U5965 (N_5965,N_4852,N_3596);
or U5966 (N_5966,N_4929,N_3481);
and U5967 (N_5967,N_3985,N_3659);
nand U5968 (N_5968,N_3989,N_2541);
xnor U5969 (N_5969,N_3545,N_3551);
nand U5970 (N_5970,N_3851,N_3919);
and U5971 (N_5971,N_4347,N_4841);
nor U5972 (N_5972,N_3718,N_4933);
or U5973 (N_5973,N_3302,N_4486);
or U5974 (N_5974,N_3766,N_4406);
and U5975 (N_5975,N_4518,N_2581);
xor U5976 (N_5976,N_3903,N_3450);
nor U5977 (N_5977,N_4164,N_3393);
or U5978 (N_5978,N_2592,N_3731);
or U5979 (N_5979,N_2775,N_2796);
nor U5980 (N_5980,N_2977,N_3038);
nand U5981 (N_5981,N_3918,N_2908);
nor U5982 (N_5982,N_2984,N_3485);
nand U5983 (N_5983,N_3580,N_3053);
and U5984 (N_5984,N_4864,N_2730);
nor U5985 (N_5985,N_4255,N_4604);
nor U5986 (N_5986,N_3688,N_3558);
or U5987 (N_5987,N_2629,N_3111);
or U5988 (N_5988,N_2569,N_4223);
and U5989 (N_5989,N_2935,N_4249);
and U5990 (N_5990,N_3509,N_4662);
nor U5991 (N_5991,N_4639,N_3581);
and U5992 (N_5992,N_4912,N_4517);
or U5993 (N_5993,N_3740,N_4202);
or U5994 (N_5994,N_3728,N_3070);
and U5995 (N_5995,N_4867,N_4262);
or U5996 (N_5996,N_4669,N_4176);
nand U5997 (N_5997,N_3857,N_2537);
or U5998 (N_5998,N_3388,N_4986);
or U5999 (N_5999,N_4602,N_3995);
or U6000 (N_6000,N_3832,N_3208);
nand U6001 (N_6001,N_4953,N_4500);
or U6002 (N_6002,N_4416,N_3553);
or U6003 (N_6003,N_3240,N_2954);
or U6004 (N_6004,N_4804,N_4394);
nor U6005 (N_6005,N_2603,N_4567);
nor U6006 (N_6006,N_4954,N_2725);
and U6007 (N_6007,N_4572,N_2534);
or U6008 (N_6008,N_4856,N_4935);
nand U6009 (N_6009,N_3074,N_3480);
nor U6010 (N_6010,N_2634,N_3554);
and U6011 (N_6011,N_3361,N_2536);
nand U6012 (N_6012,N_4934,N_3489);
or U6013 (N_6013,N_4907,N_3830);
nand U6014 (N_6014,N_4476,N_2798);
nor U6015 (N_6015,N_3350,N_3211);
and U6016 (N_6016,N_4790,N_3782);
and U6017 (N_6017,N_4045,N_3910);
nor U6018 (N_6018,N_4272,N_4730);
nand U6019 (N_6019,N_2890,N_4259);
and U6020 (N_6020,N_3482,N_2901);
nor U6021 (N_6021,N_2754,N_2949);
nand U6022 (N_6022,N_3514,N_3321);
nor U6023 (N_6023,N_4112,N_2915);
nand U6024 (N_6024,N_3133,N_3121);
nand U6025 (N_6025,N_4438,N_3009);
and U6026 (N_6026,N_2721,N_4734);
nand U6027 (N_6027,N_4900,N_3690);
and U6028 (N_6028,N_2964,N_3598);
nand U6029 (N_6029,N_4485,N_4691);
and U6030 (N_6030,N_4452,N_3303);
nor U6031 (N_6031,N_4613,N_2596);
and U6032 (N_6032,N_3316,N_4927);
and U6033 (N_6033,N_3562,N_4134);
or U6034 (N_6034,N_4464,N_4117);
nand U6035 (N_6035,N_3002,N_3672);
or U6036 (N_6036,N_4548,N_4314);
and U6037 (N_6037,N_4499,N_4468);
or U6038 (N_6038,N_2680,N_4418);
and U6039 (N_6039,N_4626,N_4299);
and U6040 (N_6040,N_4985,N_4707);
and U6041 (N_6041,N_2835,N_3882);
or U6042 (N_6042,N_4937,N_4378);
nor U6043 (N_6043,N_3008,N_2531);
and U6044 (N_6044,N_2946,N_3294);
and U6045 (N_6045,N_4781,N_2727);
xor U6046 (N_6046,N_3332,N_4706);
nor U6047 (N_6047,N_3182,N_3424);
nand U6048 (N_6048,N_4808,N_2987);
or U6049 (N_6049,N_3980,N_3082);
nand U6050 (N_6050,N_3941,N_2549);
nand U6051 (N_6051,N_3488,N_4655);
and U6052 (N_6052,N_2983,N_3453);
nand U6053 (N_6053,N_3975,N_3156);
nand U6054 (N_6054,N_4241,N_3992);
nand U6055 (N_6055,N_2950,N_4974);
nor U6056 (N_6056,N_3041,N_2981);
nand U6057 (N_6057,N_2842,N_3247);
and U6058 (N_6058,N_3862,N_3859);
and U6059 (N_6059,N_4762,N_3543);
or U6060 (N_6060,N_2708,N_2979);
nor U6061 (N_6061,N_2637,N_3383);
and U6062 (N_6062,N_4273,N_2826);
nand U6063 (N_6063,N_4281,N_2815);
nand U6064 (N_6064,N_3001,N_3462);
nor U6065 (N_6065,N_3502,N_3275);
nor U6066 (N_6066,N_3484,N_3550);
nor U6067 (N_6067,N_3499,N_3542);
nor U6068 (N_6068,N_2761,N_4525);
nand U6069 (N_6069,N_2801,N_2988);
or U6070 (N_6070,N_2683,N_4179);
nor U6071 (N_6071,N_3305,N_2633);
and U6072 (N_6072,N_2686,N_3625);
or U6073 (N_6073,N_2657,N_3107);
nor U6074 (N_6074,N_2777,N_2888);
and U6075 (N_6075,N_4502,N_4796);
or U6076 (N_6076,N_4774,N_4414);
nor U6077 (N_6077,N_4720,N_4238);
nor U6078 (N_6078,N_2687,N_4297);
nor U6079 (N_6079,N_3258,N_3174);
and U6080 (N_6080,N_3756,N_4501);
nand U6081 (N_6081,N_3856,N_3904);
xnor U6082 (N_6082,N_2595,N_3122);
or U6083 (N_6083,N_3752,N_4646);
nand U6084 (N_6084,N_4926,N_4295);
and U6085 (N_6085,N_2613,N_4410);
nor U6086 (N_6086,N_4606,N_3441);
nand U6087 (N_6087,N_2866,N_4802);
or U6088 (N_6088,N_2832,N_4562);
nor U6089 (N_6089,N_4470,N_3930);
nand U6090 (N_6090,N_3127,N_4237);
nor U6091 (N_6091,N_3500,N_3569);
nand U6092 (N_6092,N_3524,N_3898);
nor U6093 (N_6093,N_3246,N_2993);
nor U6094 (N_6094,N_4973,N_2645);
or U6095 (N_6095,N_3222,N_2638);
nor U6096 (N_6096,N_3368,N_2619);
or U6097 (N_6097,N_4569,N_4657);
nand U6098 (N_6098,N_4665,N_2969);
nor U6099 (N_6099,N_3353,N_3410);
nand U6100 (N_6100,N_3734,N_4026);
nor U6101 (N_6101,N_4908,N_4020);
or U6102 (N_6102,N_2663,N_4885);
or U6103 (N_6103,N_4947,N_3644);
or U6104 (N_6104,N_3834,N_4287);
nand U6105 (N_6105,N_3466,N_4733);
nand U6106 (N_6106,N_3676,N_4776);
and U6107 (N_6107,N_4991,N_4143);
nor U6108 (N_6108,N_3059,N_4146);
and U6109 (N_6109,N_2840,N_2557);
nand U6110 (N_6110,N_3440,N_2661);
nor U6111 (N_6111,N_4684,N_4635);
nor U6112 (N_6112,N_4063,N_4128);
nor U6113 (N_6113,N_4779,N_4573);
nand U6114 (N_6114,N_4737,N_3632);
and U6115 (N_6115,N_4875,N_4348);
nor U6116 (N_6116,N_4398,N_3129);
nor U6117 (N_6117,N_4736,N_4708);
xor U6118 (N_6118,N_3701,N_2718);
nor U6119 (N_6119,N_3108,N_3872);
or U6120 (N_6120,N_3994,N_4044);
nor U6121 (N_6121,N_4108,N_4571);
or U6122 (N_6122,N_2689,N_3094);
and U6123 (N_6123,N_3381,N_3674);
nand U6124 (N_6124,N_4441,N_3199);
nor U6125 (N_6125,N_4315,N_4058);
or U6126 (N_6126,N_4321,N_2903);
nand U6127 (N_6127,N_3730,N_3707);
nor U6128 (N_6128,N_4101,N_2848);
nor U6129 (N_6129,N_2732,N_4585);
and U6130 (N_6130,N_4660,N_4514);
nand U6131 (N_6131,N_4035,N_3269);
nand U6132 (N_6132,N_3437,N_2995);
and U6133 (N_6133,N_3682,N_3664);
nor U6134 (N_6134,N_4866,N_4847);
nand U6135 (N_6135,N_2973,N_3184);
and U6136 (N_6136,N_4598,N_2734);
nor U6137 (N_6137,N_4643,N_4515);
or U6138 (N_6138,N_3586,N_2898);
or U6139 (N_6139,N_2587,N_3145);
or U6140 (N_6140,N_3821,N_4873);
and U6141 (N_6141,N_4780,N_3418);
and U6142 (N_6142,N_4833,N_3249);
nand U6143 (N_6143,N_2872,N_3535);
nand U6144 (N_6144,N_4959,N_3202);
nor U6145 (N_6145,N_4156,N_4275);
nor U6146 (N_6146,N_3504,N_2896);
nor U6147 (N_6147,N_3576,N_2590);
and U6148 (N_6148,N_3627,N_3537);
and U6149 (N_6149,N_4349,N_3359);
nor U6150 (N_6150,N_3295,N_2789);
or U6151 (N_6151,N_3508,N_4788);
and U6152 (N_6152,N_4353,N_3152);
nor U6153 (N_6153,N_4150,N_3971);
or U6154 (N_6154,N_4142,N_3454);
and U6155 (N_6155,N_4256,N_4038);
and U6156 (N_6156,N_2636,N_4162);
and U6157 (N_6157,N_4913,N_4246);
and U6158 (N_6158,N_2504,N_3692);
nand U6159 (N_6159,N_4807,N_3147);
nand U6160 (N_6160,N_4703,N_2695);
or U6161 (N_6161,N_2864,N_2697);
or U6162 (N_6162,N_2843,N_3840);
nand U6163 (N_6163,N_3032,N_4770);
and U6164 (N_6164,N_3833,N_3487);
or U6165 (N_6165,N_3363,N_3933);
nor U6166 (N_6166,N_4454,N_2548);
and U6167 (N_6167,N_4036,N_3154);
or U6168 (N_6168,N_4683,N_4551);
or U6169 (N_6169,N_2575,N_3468);
and U6170 (N_6170,N_4046,N_3096);
nor U6171 (N_6171,N_2760,N_4168);
or U6172 (N_6172,N_2512,N_4190);
nand U6173 (N_6173,N_4766,N_4744);
nand U6174 (N_6174,N_4898,N_4966);
or U6175 (N_6175,N_4641,N_4624);
nor U6176 (N_6176,N_4482,N_3603);
nand U6177 (N_6177,N_4140,N_3977);
nor U6178 (N_6178,N_2917,N_4664);
nand U6179 (N_6179,N_4004,N_4400);
or U6180 (N_6180,N_4547,N_4630);
or U6181 (N_6181,N_4663,N_3010);
nor U6182 (N_6182,N_4539,N_3881);
and U6183 (N_6183,N_2972,N_3813);
nand U6184 (N_6184,N_3374,N_3704);
or U6185 (N_6185,N_3629,N_4264);
nand U6186 (N_6186,N_2738,N_4570);
nor U6187 (N_6187,N_4274,N_3178);
and U6188 (N_6188,N_3803,N_3027);
nor U6189 (N_6189,N_4617,N_4658);
nand U6190 (N_6190,N_4061,N_3609);
and U6191 (N_6191,N_3600,N_4505);
nand U6192 (N_6192,N_4228,N_3511);
nand U6193 (N_6193,N_4130,N_2648);
nor U6194 (N_6194,N_2976,N_3088);
nor U6195 (N_6195,N_4923,N_4267);
nand U6196 (N_6196,N_2811,N_3072);
or U6197 (N_6197,N_4090,N_3063);
and U6198 (N_6198,N_3398,N_2685);
or U6199 (N_6199,N_2913,N_2579);
or U6200 (N_6200,N_3110,N_3934);
and U6201 (N_6201,N_3439,N_3673);
or U6202 (N_6202,N_3816,N_4717);
nor U6203 (N_6203,N_3036,N_2741);
nor U6204 (N_6204,N_2700,N_3253);
and U6205 (N_6205,N_4771,N_3744);
or U6206 (N_6206,N_2750,N_3650);
and U6207 (N_6207,N_2529,N_4640);
nor U6208 (N_6208,N_4265,N_2844);
nor U6209 (N_6209,N_4845,N_4304);
nand U6210 (N_6210,N_4192,N_3177);
and U6211 (N_6211,N_2712,N_2641);
and U6212 (N_6212,N_3306,N_3957);
nor U6213 (N_6213,N_4998,N_3981);
nor U6214 (N_6214,N_3262,N_2660);
or U6215 (N_6215,N_2507,N_3646);
and U6216 (N_6216,N_2524,N_2878);
and U6217 (N_6217,N_4909,N_4251);
nor U6218 (N_6218,N_4231,N_4107);
nand U6219 (N_6219,N_3185,N_3722);
xor U6220 (N_6220,N_4519,N_2874);
nand U6221 (N_6221,N_3076,N_4618);
or U6222 (N_6222,N_4208,N_4280);
and U6223 (N_6223,N_3225,N_3775);
nand U6224 (N_6224,N_3433,N_2938);
nor U6225 (N_6225,N_3261,N_4865);
and U6226 (N_6226,N_2517,N_4894);
nor U6227 (N_6227,N_2873,N_2731);
nor U6228 (N_6228,N_3571,N_4820);
or U6229 (N_6229,N_4330,N_4930);
or U6230 (N_6230,N_3723,N_3927);
nor U6231 (N_6231,N_3445,N_3329);
nor U6232 (N_6232,N_3458,N_4075);
and U6233 (N_6233,N_4553,N_3385);
nor U6234 (N_6234,N_2589,N_4104);
nand U6235 (N_6235,N_2774,N_4317);
and U6236 (N_6236,N_3953,N_2767);
nand U6237 (N_6237,N_3616,N_4919);
and U6238 (N_6238,N_3102,N_3340);
and U6239 (N_6239,N_3599,N_4940);
nand U6240 (N_6240,N_3958,N_2923);
nor U6241 (N_6241,N_4324,N_3626);
nand U6242 (N_6242,N_2597,N_4946);
nor U6243 (N_6243,N_3016,N_4056);
or U6244 (N_6244,N_2855,N_3897);
or U6245 (N_6245,N_4014,N_3200);
and U6246 (N_6246,N_4896,N_3611);
nand U6247 (N_6247,N_3679,N_2535);
and U6248 (N_6248,N_2665,N_3024);
or U6249 (N_6249,N_3465,N_2962);
nor U6250 (N_6250,N_3851,N_3603);
nor U6251 (N_6251,N_4921,N_4057);
nor U6252 (N_6252,N_4810,N_4641);
and U6253 (N_6253,N_4610,N_4605);
or U6254 (N_6254,N_3639,N_4223);
or U6255 (N_6255,N_2824,N_4612);
nand U6256 (N_6256,N_4916,N_4379);
nand U6257 (N_6257,N_3452,N_4760);
nor U6258 (N_6258,N_3858,N_3338);
nor U6259 (N_6259,N_4021,N_4833);
or U6260 (N_6260,N_4474,N_4636);
or U6261 (N_6261,N_3614,N_3575);
or U6262 (N_6262,N_4165,N_3058);
nor U6263 (N_6263,N_3692,N_4605);
or U6264 (N_6264,N_4396,N_3791);
and U6265 (N_6265,N_2847,N_4361);
or U6266 (N_6266,N_3639,N_4252);
nor U6267 (N_6267,N_4480,N_3790);
nand U6268 (N_6268,N_3762,N_4430);
nor U6269 (N_6269,N_3804,N_4882);
or U6270 (N_6270,N_3545,N_2667);
or U6271 (N_6271,N_3752,N_4238);
and U6272 (N_6272,N_2898,N_3915);
nand U6273 (N_6273,N_4893,N_3457);
and U6274 (N_6274,N_4848,N_4008);
nor U6275 (N_6275,N_4833,N_4559);
and U6276 (N_6276,N_3107,N_2719);
nand U6277 (N_6277,N_3601,N_2921);
or U6278 (N_6278,N_2692,N_2796);
and U6279 (N_6279,N_3290,N_3884);
nand U6280 (N_6280,N_4930,N_2595);
nor U6281 (N_6281,N_3983,N_3559);
and U6282 (N_6282,N_4642,N_4691);
and U6283 (N_6283,N_4268,N_3091);
or U6284 (N_6284,N_4670,N_4357);
nand U6285 (N_6285,N_4626,N_2642);
nand U6286 (N_6286,N_4452,N_3312);
and U6287 (N_6287,N_2731,N_4167);
nand U6288 (N_6288,N_4349,N_3109);
nor U6289 (N_6289,N_3685,N_3036);
and U6290 (N_6290,N_3149,N_3789);
nand U6291 (N_6291,N_3280,N_3519);
or U6292 (N_6292,N_4827,N_3372);
or U6293 (N_6293,N_2905,N_3116);
nand U6294 (N_6294,N_2873,N_4268);
nor U6295 (N_6295,N_3127,N_4009);
or U6296 (N_6296,N_3207,N_3034);
nand U6297 (N_6297,N_4668,N_4601);
xor U6298 (N_6298,N_3239,N_3272);
nor U6299 (N_6299,N_4762,N_4400);
nand U6300 (N_6300,N_4050,N_2984);
nor U6301 (N_6301,N_4520,N_2758);
nor U6302 (N_6302,N_4633,N_2554);
nand U6303 (N_6303,N_3007,N_3098);
xnor U6304 (N_6304,N_4493,N_2646);
and U6305 (N_6305,N_3406,N_3674);
xnor U6306 (N_6306,N_3298,N_3026);
and U6307 (N_6307,N_3532,N_3445);
nand U6308 (N_6308,N_4779,N_4578);
and U6309 (N_6309,N_2541,N_4248);
nor U6310 (N_6310,N_2857,N_2862);
and U6311 (N_6311,N_3154,N_4413);
nor U6312 (N_6312,N_3022,N_4243);
xnor U6313 (N_6313,N_2677,N_4274);
and U6314 (N_6314,N_3583,N_4543);
and U6315 (N_6315,N_4272,N_3467);
and U6316 (N_6316,N_3183,N_4152);
nor U6317 (N_6317,N_2903,N_3179);
nor U6318 (N_6318,N_4689,N_4140);
xor U6319 (N_6319,N_4617,N_3709);
nand U6320 (N_6320,N_4644,N_2890);
nand U6321 (N_6321,N_2702,N_3188);
or U6322 (N_6322,N_4386,N_3343);
nand U6323 (N_6323,N_3426,N_2535);
and U6324 (N_6324,N_3706,N_4233);
nor U6325 (N_6325,N_4827,N_2818);
nand U6326 (N_6326,N_3590,N_4250);
nand U6327 (N_6327,N_3396,N_4443);
and U6328 (N_6328,N_4118,N_2676);
xnor U6329 (N_6329,N_4663,N_4121);
nor U6330 (N_6330,N_2862,N_3176);
and U6331 (N_6331,N_3764,N_3373);
nor U6332 (N_6332,N_3066,N_4185);
xor U6333 (N_6333,N_3345,N_2786);
and U6334 (N_6334,N_2969,N_4276);
nand U6335 (N_6335,N_3610,N_3755);
and U6336 (N_6336,N_2948,N_3427);
and U6337 (N_6337,N_3804,N_4074);
and U6338 (N_6338,N_3468,N_4330);
nand U6339 (N_6339,N_3800,N_4181);
nand U6340 (N_6340,N_4544,N_4711);
nand U6341 (N_6341,N_2586,N_3332);
or U6342 (N_6342,N_3037,N_3692);
nor U6343 (N_6343,N_4837,N_4979);
nor U6344 (N_6344,N_3824,N_4524);
and U6345 (N_6345,N_3142,N_3341);
nand U6346 (N_6346,N_2659,N_4643);
and U6347 (N_6347,N_4696,N_2824);
or U6348 (N_6348,N_4132,N_4175);
nor U6349 (N_6349,N_2798,N_4492);
and U6350 (N_6350,N_2625,N_4778);
nor U6351 (N_6351,N_3909,N_3644);
or U6352 (N_6352,N_4468,N_4540);
nor U6353 (N_6353,N_3178,N_3832);
or U6354 (N_6354,N_4298,N_3046);
nor U6355 (N_6355,N_4776,N_3662);
nand U6356 (N_6356,N_3093,N_2643);
or U6357 (N_6357,N_4217,N_3100);
and U6358 (N_6358,N_4085,N_3001);
or U6359 (N_6359,N_3906,N_3639);
nand U6360 (N_6360,N_3439,N_4142);
nand U6361 (N_6361,N_4357,N_3599);
nor U6362 (N_6362,N_4086,N_4040);
nand U6363 (N_6363,N_4131,N_3469);
and U6364 (N_6364,N_2970,N_3104);
nor U6365 (N_6365,N_3987,N_4220);
and U6366 (N_6366,N_4616,N_3332);
or U6367 (N_6367,N_4494,N_4708);
nor U6368 (N_6368,N_3902,N_4433);
or U6369 (N_6369,N_4978,N_3380);
nand U6370 (N_6370,N_3956,N_3057);
nor U6371 (N_6371,N_4496,N_4939);
or U6372 (N_6372,N_4971,N_2714);
nor U6373 (N_6373,N_3896,N_3072);
and U6374 (N_6374,N_4398,N_4496);
and U6375 (N_6375,N_4612,N_2840);
and U6376 (N_6376,N_3471,N_3347);
or U6377 (N_6377,N_3028,N_4823);
nor U6378 (N_6378,N_2546,N_4385);
and U6379 (N_6379,N_4882,N_4827);
and U6380 (N_6380,N_4695,N_4853);
nand U6381 (N_6381,N_4091,N_4440);
nand U6382 (N_6382,N_3253,N_4761);
nor U6383 (N_6383,N_4945,N_3260);
and U6384 (N_6384,N_2577,N_4243);
or U6385 (N_6385,N_3816,N_3019);
and U6386 (N_6386,N_2554,N_4802);
or U6387 (N_6387,N_4624,N_4120);
and U6388 (N_6388,N_2725,N_4880);
or U6389 (N_6389,N_4058,N_3568);
nor U6390 (N_6390,N_3122,N_3829);
and U6391 (N_6391,N_4389,N_4803);
nand U6392 (N_6392,N_3461,N_2775);
and U6393 (N_6393,N_3821,N_4059);
nor U6394 (N_6394,N_4790,N_4772);
nor U6395 (N_6395,N_3125,N_4366);
nor U6396 (N_6396,N_4466,N_3583);
nor U6397 (N_6397,N_3096,N_4216);
nand U6398 (N_6398,N_4143,N_3763);
xnor U6399 (N_6399,N_3710,N_4369);
xnor U6400 (N_6400,N_2740,N_4420);
and U6401 (N_6401,N_3222,N_2707);
and U6402 (N_6402,N_4128,N_3828);
and U6403 (N_6403,N_2593,N_2847);
or U6404 (N_6404,N_4111,N_3901);
nand U6405 (N_6405,N_4644,N_4943);
xnor U6406 (N_6406,N_2681,N_2779);
nor U6407 (N_6407,N_4451,N_4679);
or U6408 (N_6408,N_2601,N_2879);
or U6409 (N_6409,N_4849,N_4597);
nor U6410 (N_6410,N_3981,N_4165);
nor U6411 (N_6411,N_3848,N_4860);
nor U6412 (N_6412,N_3169,N_4445);
nor U6413 (N_6413,N_4645,N_3399);
nand U6414 (N_6414,N_4074,N_4665);
and U6415 (N_6415,N_2876,N_2860);
nor U6416 (N_6416,N_3171,N_3389);
nand U6417 (N_6417,N_3780,N_4459);
nand U6418 (N_6418,N_2824,N_3576);
nor U6419 (N_6419,N_3561,N_4832);
nand U6420 (N_6420,N_4260,N_3519);
or U6421 (N_6421,N_2596,N_2548);
or U6422 (N_6422,N_3397,N_3047);
nor U6423 (N_6423,N_3439,N_4466);
nor U6424 (N_6424,N_4966,N_3525);
or U6425 (N_6425,N_3208,N_2511);
and U6426 (N_6426,N_2696,N_4999);
nor U6427 (N_6427,N_4069,N_3835);
nand U6428 (N_6428,N_2984,N_2771);
nand U6429 (N_6429,N_3472,N_4032);
nand U6430 (N_6430,N_2743,N_4515);
nor U6431 (N_6431,N_2632,N_4928);
nand U6432 (N_6432,N_2805,N_4308);
or U6433 (N_6433,N_3698,N_2803);
xnor U6434 (N_6434,N_2895,N_3578);
and U6435 (N_6435,N_2526,N_3555);
or U6436 (N_6436,N_4689,N_4026);
or U6437 (N_6437,N_3313,N_2623);
nor U6438 (N_6438,N_3750,N_4833);
nor U6439 (N_6439,N_4954,N_3987);
nor U6440 (N_6440,N_4199,N_2673);
xor U6441 (N_6441,N_4732,N_3689);
or U6442 (N_6442,N_4155,N_3889);
or U6443 (N_6443,N_4169,N_4829);
nand U6444 (N_6444,N_4175,N_3153);
or U6445 (N_6445,N_3914,N_2716);
or U6446 (N_6446,N_3806,N_4680);
xor U6447 (N_6447,N_4418,N_4050);
or U6448 (N_6448,N_4098,N_4112);
nand U6449 (N_6449,N_4825,N_4249);
and U6450 (N_6450,N_2754,N_3392);
or U6451 (N_6451,N_4880,N_2702);
nor U6452 (N_6452,N_3346,N_3823);
and U6453 (N_6453,N_3967,N_4045);
and U6454 (N_6454,N_2540,N_3932);
nor U6455 (N_6455,N_2961,N_2806);
and U6456 (N_6456,N_3334,N_4851);
and U6457 (N_6457,N_3070,N_4475);
nand U6458 (N_6458,N_4233,N_4197);
nor U6459 (N_6459,N_2758,N_3762);
nand U6460 (N_6460,N_3040,N_3006);
nand U6461 (N_6461,N_3988,N_3768);
and U6462 (N_6462,N_3229,N_4045);
nand U6463 (N_6463,N_2659,N_4686);
or U6464 (N_6464,N_4103,N_3164);
nand U6465 (N_6465,N_3263,N_4814);
nor U6466 (N_6466,N_3358,N_2809);
nand U6467 (N_6467,N_4641,N_4167);
nand U6468 (N_6468,N_3029,N_4787);
nor U6469 (N_6469,N_3176,N_4922);
or U6470 (N_6470,N_2542,N_3693);
nor U6471 (N_6471,N_4877,N_3155);
nor U6472 (N_6472,N_2738,N_3398);
nand U6473 (N_6473,N_4255,N_4801);
nand U6474 (N_6474,N_4667,N_4024);
nor U6475 (N_6475,N_2671,N_2616);
nand U6476 (N_6476,N_3621,N_4625);
nor U6477 (N_6477,N_4244,N_2982);
nand U6478 (N_6478,N_3811,N_3324);
nor U6479 (N_6479,N_3469,N_2962);
nor U6480 (N_6480,N_2967,N_3816);
nor U6481 (N_6481,N_4931,N_2785);
xnor U6482 (N_6482,N_3547,N_4814);
or U6483 (N_6483,N_4719,N_3792);
or U6484 (N_6484,N_3599,N_4748);
and U6485 (N_6485,N_3623,N_2643);
nand U6486 (N_6486,N_4104,N_3382);
nor U6487 (N_6487,N_4595,N_2755);
and U6488 (N_6488,N_4848,N_2808);
nor U6489 (N_6489,N_4629,N_3477);
or U6490 (N_6490,N_2838,N_2588);
nand U6491 (N_6491,N_3214,N_4706);
nand U6492 (N_6492,N_3491,N_4546);
or U6493 (N_6493,N_2627,N_3141);
or U6494 (N_6494,N_2830,N_2955);
or U6495 (N_6495,N_3460,N_3988);
and U6496 (N_6496,N_2776,N_3090);
or U6497 (N_6497,N_3206,N_4129);
nor U6498 (N_6498,N_2862,N_4042);
nand U6499 (N_6499,N_2907,N_3298);
and U6500 (N_6500,N_3813,N_3077);
and U6501 (N_6501,N_3032,N_3778);
nor U6502 (N_6502,N_4711,N_2980);
nand U6503 (N_6503,N_3489,N_2824);
nor U6504 (N_6504,N_4702,N_2605);
and U6505 (N_6505,N_4538,N_4827);
nand U6506 (N_6506,N_4993,N_3574);
and U6507 (N_6507,N_4967,N_4528);
nand U6508 (N_6508,N_3814,N_3153);
and U6509 (N_6509,N_4674,N_3654);
or U6510 (N_6510,N_3532,N_3788);
nand U6511 (N_6511,N_3560,N_4951);
nor U6512 (N_6512,N_4063,N_4135);
nor U6513 (N_6513,N_4143,N_2741);
or U6514 (N_6514,N_3868,N_3196);
and U6515 (N_6515,N_3869,N_3123);
xnor U6516 (N_6516,N_4006,N_3970);
and U6517 (N_6517,N_3812,N_2968);
nor U6518 (N_6518,N_4295,N_3121);
or U6519 (N_6519,N_4107,N_4867);
and U6520 (N_6520,N_4577,N_4235);
nor U6521 (N_6521,N_2865,N_3714);
nand U6522 (N_6522,N_4178,N_3373);
and U6523 (N_6523,N_4312,N_4754);
and U6524 (N_6524,N_4339,N_2854);
nand U6525 (N_6525,N_2530,N_4925);
or U6526 (N_6526,N_3586,N_3644);
and U6527 (N_6527,N_4763,N_3489);
nand U6528 (N_6528,N_2747,N_3748);
or U6529 (N_6529,N_2640,N_4552);
or U6530 (N_6530,N_2711,N_2666);
or U6531 (N_6531,N_2858,N_3379);
nand U6532 (N_6532,N_2576,N_3811);
and U6533 (N_6533,N_4391,N_2774);
and U6534 (N_6534,N_3918,N_4563);
nor U6535 (N_6535,N_2952,N_3057);
and U6536 (N_6536,N_3322,N_4801);
nand U6537 (N_6537,N_4598,N_2986);
nor U6538 (N_6538,N_4345,N_4305);
and U6539 (N_6539,N_2775,N_3607);
or U6540 (N_6540,N_4832,N_3715);
or U6541 (N_6541,N_3702,N_3284);
nor U6542 (N_6542,N_3681,N_2550);
or U6543 (N_6543,N_4585,N_3901);
and U6544 (N_6544,N_2954,N_3613);
nand U6545 (N_6545,N_4566,N_4069);
and U6546 (N_6546,N_4359,N_3183);
nor U6547 (N_6547,N_3634,N_4597);
nand U6548 (N_6548,N_3351,N_3472);
or U6549 (N_6549,N_3392,N_3447);
or U6550 (N_6550,N_2650,N_2870);
or U6551 (N_6551,N_4355,N_3489);
nor U6552 (N_6552,N_4049,N_4597);
and U6553 (N_6553,N_2948,N_3836);
and U6554 (N_6554,N_2617,N_3105);
nor U6555 (N_6555,N_3310,N_3429);
nand U6556 (N_6556,N_4301,N_4817);
nand U6557 (N_6557,N_3215,N_3908);
nand U6558 (N_6558,N_2879,N_4626);
nor U6559 (N_6559,N_4661,N_3176);
nor U6560 (N_6560,N_4722,N_3166);
nand U6561 (N_6561,N_3836,N_4401);
and U6562 (N_6562,N_4090,N_4531);
nand U6563 (N_6563,N_2516,N_4784);
and U6564 (N_6564,N_2846,N_2663);
and U6565 (N_6565,N_4546,N_2565);
and U6566 (N_6566,N_3106,N_3034);
nand U6567 (N_6567,N_3467,N_3754);
xor U6568 (N_6568,N_4098,N_3372);
nand U6569 (N_6569,N_2712,N_4891);
nand U6570 (N_6570,N_2601,N_4768);
nand U6571 (N_6571,N_2629,N_4686);
nand U6572 (N_6572,N_2519,N_3607);
and U6573 (N_6573,N_4001,N_2752);
nor U6574 (N_6574,N_4064,N_4538);
and U6575 (N_6575,N_2717,N_3724);
or U6576 (N_6576,N_3150,N_2866);
and U6577 (N_6577,N_4245,N_4888);
and U6578 (N_6578,N_3863,N_3827);
nor U6579 (N_6579,N_3705,N_4038);
nand U6580 (N_6580,N_3114,N_3998);
nand U6581 (N_6581,N_3565,N_4454);
or U6582 (N_6582,N_3164,N_4303);
xnor U6583 (N_6583,N_4064,N_3100);
or U6584 (N_6584,N_2687,N_4311);
nand U6585 (N_6585,N_2658,N_4442);
xor U6586 (N_6586,N_2979,N_3193);
nor U6587 (N_6587,N_4744,N_4385);
xor U6588 (N_6588,N_4484,N_3420);
nand U6589 (N_6589,N_3955,N_3772);
nand U6590 (N_6590,N_4725,N_2753);
nor U6591 (N_6591,N_2967,N_3168);
and U6592 (N_6592,N_2527,N_2994);
and U6593 (N_6593,N_2870,N_3771);
nand U6594 (N_6594,N_3304,N_3036);
and U6595 (N_6595,N_4017,N_4615);
or U6596 (N_6596,N_4787,N_3354);
nand U6597 (N_6597,N_3688,N_4266);
and U6598 (N_6598,N_4650,N_3066);
and U6599 (N_6599,N_3796,N_3054);
xnor U6600 (N_6600,N_2887,N_4086);
nor U6601 (N_6601,N_3574,N_3556);
nand U6602 (N_6602,N_3794,N_3678);
nand U6603 (N_6603,N_3059,N_4133);
and U6604 (N_6604,N_2529,N_2614);
nand U6605 (N_6605,N_3305,N_3672);
and U6606 (N_6606,N_3636,N_3104);
or U6607 (N_6607,N_2523,N_4909);
or U6608 (N_6608,N_3979,N_3599);
and U6609 (N_6609,N_3110,N_4939);
nor U6610 (N_6610,N_4610,N_3338);
and U6611 (N_6611,N_2573,N_2542);
or U6612 (N_6612,N_2753,N_4410);
nand U6613 (N_6613,N_3296,N_3818);
nand U6614 (N_6614,N_4050,N_3341);
nor U6615 (N_6615,N_3201,N_3176);
nor U6616 (N_6616,N_2672,N_4812);
nor U6617 (N_6617,N_4837,N_4787);
and U6618 (N_6618,N_3132,N_4546);
nor U6619 (N_6619,N_3974,N_4323);
or U6620 (N_6620,N_3688,N_3614);
and U6621 (N_6621,N_4157,N_3424);
nand U6622 (N_6622,N_3177,N_3191);
nor U6623 (N_6623,N_4693,N_4544);
nor U6624 (N_6624,N_2754,N_4395);
nand U6625 (N_6625,N_2839,N_3087);
and U6626 (N_6626,N_3718,N_4165);
or U6627 (N_6627,N_4171,N_3931);
or U6628 (N_6628,N_4131,N_4411);
nor U6629 (N_6629,N_2869,N_3421);
nor U6630 (N_6630,N_3408,N_4413);
or U6631 (N_6631,N_4016,N_4359);
or U6632 (N_6632,N_3902,N_4978);
nor U6633 (N_6633,N_3300,N_4980);
nand U6634 (N_6634,N_3192,N_4349);
and U6635 (N_6635,N_3192,N_4905);
and U6636 (N_6636,N_3229,N_2945);
nor U6637 (N_6637,N_4470,N_2982);
nand U6638 (N_6638,N_2579,N_3086);
or U6639 (N_6639,N_2914,N_4290);
or U6640 (N_6640,N_3972,N_4483);
and U6641 (N_6641,N_3234,N_3775);
and U6642 (N_6642,N_4096,N_3626);
nor U6643 (N_6643,N_2637,N_2793);
nand U6644 (N_6644,N_3241,N_4795);
or U6645 (N_6645,N_2741,N_2684);
nand U6646 (N_6646,N_4357,N_4833);
xnor U6647 (N_6647,N_4394,N_3382);
or U6648 (N_6648,N_4187,N_2680);
or U6649 (N_6649,N_2968,N_3462);
and U6650 (N_6650,N_3073,N_4670);
nand U6651 (N_6651,N_3663,N_3770);
nand U6652 (N_6652,N_4529,N_3181);
nor U6653 (N_6653,N_4067,N_4171);
and U6654 (N_6654,N_3638,N_4654);
nand U6655 (N_6655,N_4626,N_4180);
and U6656 (N_6656,N_4314,N_4305);
or U6657 (N_6657,N_3350,N_2596);
or U6658 (N_6658,N_3959,N_2506);
xnor U6659 (N_6659,N_3611,N_3867);
nand U6660 (N_6660,N_4048,N_2832);
or U6661 (N_6661,N_4052,N_4317);
nor U6662 (N_6662,N_4610,N_2905);
nor U6663 (N_6663,N_3282,N_4607);
and U6664 (N_6664,N_3776,N_3779);
or U6665 (N_6665,N_4035,N_3874);
nand U6666 (N_6666,N_3066,N_2767);
nor U6667 (N_6667,N_3205,N_4956);
and U6668 (N_6668,N_3777,N_4870);
or U6669 (N_6669,N_3200,N_3412);
and U6670 (N_6670,N_3822,N_4508);
nand U6671 (N_6671,N_3126,N_3103);
and U6672 (N_6672,N_4954,N_4840);
and U6673 (N_6673,N_3571,N_4241);
or U6674 (N_6674,N_3854,N_2732);
or U6675 (N_6675,N_4565,N_3206);
nor U6676 (N_6676,N_3390,N_2805);
and U6677 (N_6677,N_2750,N_4132);
and U6678 (N_6678,N_3730,N_2794);
nor U6679 (N_6679,N_4275,N_3626);
and U6680 (N_6680,N_4301,N_2822);
and U6681 (N_6681,N_4813,N_4006);
nand U6682 (N_6682,N_4402,N_3548);
nand U6683 (N_6683,N_4585,N_3162);
xor U6684 (N_6684,N_3195,N_2814);
nor U6685 (N_6685,N_2731,N_2887);
nand U6686 (N_6686,N_3094,N_2661);
or U6687 (N_6687,N_3979,N_4976);
and U6688 (N_6688,N_3776,N_3789);
or U6689 (N_6689,N_4999,N_3999);
xnor U6690 (N_6690,N_3848,N_4498);
or U6691 (N_6691,N_4519,N_4100);
or U6692 (N_6692,N_2513,N_4161);
and U6693 (N_6693,N_4701,N_3522);
and U6694 (N_6694,N_2845,N_2516);
or U6695 (N_6695,N_4951,N_4051);
and U6696 (N_6696,N_3348,N_3846);
or U6697 (N_6697,N_4737,N_4905);
or U6698 (N_6698,N_4155,N_4109);
xnor U6699 (N_6699,N_4647,N_4880);
or U6700 (N_6700,N_3862,N_2610);
and U6701 (N_6701,N_4052,N_4662);
nand U6702 (N_6702,N_4811,N_3465);
and U6703 (N_6703,N_3978,N_2749);
nor U6704 (N_6704,N_2633,N_2914);
and U6705 (N_6705,N_4075,N_3861);
nand U6706 (N_6706,N_3856,N_4689);
nor U6707 (N_6707,N_3432,N_3157);
and U6708 (N_6708,N_4049,N_3836);
and U6709 (N_6709,N_3261,N_2707);
xor U6710 (N_6710,N_2662,N_3007);
and U6711 (N_6711,N_3759,N_3303);
or U6712 (N_6712,N_3019,N_2858);
nor U6713 (N_6713,N_3705,N_4549);
and U6714 (N_6714,N_4457,N_3288);
and U6715 (N_6715,N_4376,N_4104);
nand U6716 (N_6716,N_3093,N_4026);
nand U6717 (N_6717,N_2769,N_3266);
or U6718 (N_6718,N_4276,N_3017);
or U6719 (N_6719,N_3186,N_4194);
nand U6720 (N_6720,N_4819,N_4513);
xor U6721 (N_6721,N_4407,N_4394);
nand U6722 (N_6722,N_4271,N_3594);
nor U6723 (N_6723,N_4941,N_4965);
and U6724 (N_6724,N_3613,N_3557);
nand U6725 (N_6725,N_4970,N_3067);
nor U6726 (N_6726,N_2807,N_2667);
nor U6727 (N_6727,N_3790,N_2776);
or U6728 (N_6728,N_3003,N_4687);
nor U6729 (N_6729,N_4713,N_4502);
or U6730 (N_6730,N_3602,N_4135);
and U6731 (N_6731,N_4619,N_3071);
nand U6732 (N_6732,N_3891,N_3105);
nand U6733 (N_6733,N_3880,N_3681);
nand U6734 (N_6734,N_2636,N_3114);
nand U6735 (N_6735,N_4053,N_2686);
and U6736 (N_6736,N_4893,N_3884);
and U6737 (N_6737,N_3033,N_4632);
or U6738 (N_6738,N_3659,N_3268);
nand U6739 (N_6739,N_4841,N_3868);
nand U6740 (N_6740,N_3649,N_3397);
nor U6741 (N_6741,N_2875,N_3911);
nor U6742 (N_6742,N_2583,N_4796);
or U6743 (N_6743,N_2504,N_4172);
nand U6744 (N_6744,N_4387,N_3986);
nand U6745 (N_6745,N_2908,N_2841);
nor U6746 (N_6746,N_3995,N_2893);
nand U6747 (N_6747,N_3403,N_3267);
or U6748 (N_6748,N_3790,N_3327);
nand U6749 (N_6749,N_4446,N_3858);
nor U6750 (N_6750,N_4678,N_3884);
and U6751 (N_6751,N_4116,N_4848);
nor U6752 (N_6752,N_3011,N_4568);
nand U6753 (N_6753,N_2549,N_4537);
or U6754 (N_6754,N_3453,N_3834);
nor U6755 (N_6755,N_4669,N_2590);
and U6756 (N_6756,N_3510,N_2708);
and U6757 (N_6757,N_2740,N_2732);
nand U6758 (N_6758,N_2889,N_3821);
nor U6759 (N_6759,N_3294,N_4585);
or U6760 (N_6760,N_3674,N_4685);
nand U6761 (N_6761,N_2593,N_3341);
nor U6762 (N_6762,N_4018,N_4225);
or U6763 (N_6763,N_4513,N_4694);
nor U6764 (N_6764,N_3595,N_2656);
or U6765 (N_6765,N_4057,N_4404);
nor U6766 (N_6766,N_2755,N_3910);
nand U6767 (N_6767,N_2946,N_2583);
nor U6768 (N_6768,N_3279,N_3653);
nor U6769 (N_6769,N_3389,N_3631);
and U6770 (N_6770,N_3722,N_3943);
nand U6771 (N_6771,N_4532,N_4276);
nor U6772 (N_6772,N_3809,N_4654);
nand U6773 (N_6773,N_2530,N_2771);
nand U6774 (N_6774,N_3051,N_2905);
nor U6775 (N_6775,N_4084,N_3145);
nand U6776 (N_6776,N_4619,N_4424);
nor U6777 (N_6777,N_4198,N_3307);
or U6778 (N_6778,N_3407,N_4578);
and U6779 (N_6779,N_2964,N_4830);
nand U6780 (N_6780,N_3282,N_4460);
nand U6781 (N_6781,N_4839,N_3305);
nand U6782 (N_6782,N_2995,N_2861);
and U6783 (N_6783,N_3626,N_4637);
nand U6784 (N_6784,N_3550,N_4994);
or U6785 (N_6785,N_2501,N_4464);
nand U6786 (N_6786,N_3324,N_4919);
nand U6787 (N_6787,N_3185,N_2966);
or U6788 (N_6788,N_4378,N_4915);
nand U6789 (N_6789,N_4244,N_3632);
and U6790 (N_6790,N_4732,N_3366);
and U6791 (N_6791,N_2583,N_4715);
and U6792 (N_6792,N_3648,N_4210);
nor U6793 (N_6793,N_3442,N_3549);
or U6794 (N_6794,N_3920,N_4612);
nand U6795 (N_6795,N_4374,N_4476);
or U6796 (N_6796,N_2924,N_3771);
nor U6797 (N_6797,N_2986,N_4349);
or U6798 (N_6798,N_3364,N_2909);
nand U6799 (N_6799,N_2830,N_4832);
nand U6800 (N_6800,N_2588,N_2847);
or U6801 (N_6801,N_3651,N_4712);
or U6802 (N_6802,N_3636,N_4311);
or U6803 (N_6803,N_2946,N_3567);
nand U6804 (N_6804,N_3232,N_3298);
or U6805 (N_6805,N_3065,N_3948);
nor U6806 (N_6806,N_4885,N_4055);
xor U6807 (N_6807,N_3130,N_3427);
and U6808 (N_6808,N_4769,N_4366);
or U6809 (N_6809,N_3204,N_2971);
or U6810 (N_6810,N_4743,N_3758);
nand U6811 (N_6811,N_2665,N_4303);
xor U6812 (N_6812,N_3674,N_4747);
nor U6813 (N_6813,N_3746,N_4482);
and U6814 (N_6814,N_3370,N_4432);
or U6815 (N_6815,N_3307,N_2916);
nand U6816 (N_6816,N_3578,N_3547);
or U6817 (N_6817,N_4417,N_3000);
nor U6818 (N_6818,N_4969,N_2582);
and U6819 (N_6819,N_3485,N_2663);
or U6820 (N_6820,N_4998,N_3216);
nor U6821 (N_6821,N_3412,N_3407);
nor U6822 (N_6822,N_2879,N_4277);
and U6823 (N_6823,N_2765,N_2648);
nand U6824 (N_6824,N_4229,N_4771);
nand U6825 (N_6825,N_2891,N_4743);
nor U6826 (N_6826,N_4398,N_4201);
or U6827 (N_6827,N_3924,N_4618);
or U6828 (N_6828,N_3131,N_4036);
nand U6829 (N_6829,N_4340,N_3857);
nand U6830 (N_6830,N_3479,N_2553);
nand U6831 (N_6831,N_3365,N_4815);
and U6832 (N_6832,N_2792,N_3405);
or U6833 (N_6833,N_4616,N_3360);
and U6834 (N_6834,N_2631,N_3414);
nor U6835 (N_6835,N_3020,N_3500);
and U6836 (N_6836,N_2701,N_3106);
nor U6837 (N_6837,N_3075,N_4573);
or U6838 (N_6838,N_3445,N_3781);
or U6839 (N_6839,N_4441,N_2944);
nor U6840 (N_6840,N_4579,N_4426);
nand U6841 (N_6841,N_4229,N_4375);
or U6842 (N_6842,N_3871,N_3662);
and U6843 (N_6843,N_3315,N_4204);
xor U6844 (N_6844,N_2911,N_4604);
or U6845 (N_6845,N_3969,N_3841);
or U6846 (N_6846,N_3349,N_2673);
and U6847 (N_6847,N_3345,N_4532);
nor U6848 (N_6848,N_4728,N_2721);
or U6849 (N_6849,N_4988,N_2985);
and U6850 (N_6850,N_2729,N_4462);
nor U6851 (N_6851,N_4743,N_4267);
nor U6852 (N_6852,N_3916,N_3285);
nand U6853 (N_6853,N_4354,N_3337);
or U6854 (N_6854,N_4816,N_3234);
or U6855 (N_6855,N_2643,N_3051);
nor U6856 (N_6856,N_4663,N_3667);
nand U6857 (N_6857,N_4104,N_2890);
xor U6858 (N_6858,N_3311,N_2953);
nand U6859 (N_6859,N_3797,N_4605);
or U6860 (N_6860,N_3356,N_2855);
nor U6861 (N_6861,N_3353,N_4466);
nand U6862 (N_6862,N_2587,N_3882);
or U6863 (N_6863,N_3788,N_4485);
and U6864 (N_6864,N_2933,N_4614);
nor U6865 (N_6865,N_4854,N_3701);
nor U6866 (N_6866,N_3884,N_4578);
nand U6867 (N_6867,N_4456,N_3109);
xor U6868 (N_6868,N_2846,N_4005);
nand U6869 (N_6869,N_3409,N_3344);
or U6870 (N_6870,N_3483,N_3745);
nor U6871 (N_6871,N_4972,N_3643);
xnor U6872 (N_6872,N_4330,N_3417);
or U6873 (N_6873,N_3833,N_2638);
nand U6874 (N_6874,N_4801,N_2894);
and U6875 (N_6875,N_2890,N_3787);
xor U6876 (N_6876,N_3572,N_4101);
nor U6877 (N_6877,N_2567,N_4601);
nor U6878 (N_6878,N_2555,N_2581);
or U6879 (N_6879,N_3743,N_2939);
nor U6880 (N_6880,N_4353,N_3646);
and U6881 (N_6881,N_4339,N_4506);
or U6882 (N_6882,N_4057,N_4323);
nand U6883 (N_6883,N_3153,N_4290);
or U6884 (N_6884,N_4888,N_3621);
or U6885 (N_6885,N_4328,N_4735);
or U6886 (N_6886,N_4994,N_4636);
or U6887 (N_6887,N_3916,N_4298);
or U6888 (N_6888,N_2685,N_4058);
nand U6889 (N_6889,N_3608,N_3373);
nor U6890 (N_6890,N_2833,N_3926);
or U6891 (N_6891,N_4754,N_4710);
or U6892 (N_6892,N_4769,N_3368);
nand U6893 (N_6893,N_4302,N_3248);
or U6894 (N_6894,N_4658,N_4809);
or U6895 (N_6895,N_2595,N_3904);
xor U6896 (N_6896,N_3387,N_3573);
or U6897 (N_6897,N_3870,N_3349);
and U6898 (N_6898,N_2562,N_4794);
and U6899 (N_6899,N_2533,N_3215);
or U6900 (N_6900,N_4885,N_3400);
or U6901 (N_6901,N_2540,N_2585);
nor U6902 (N_6902,N_3992,N_3617);
or U6903 (N_6903,N_2702,N_4748);
and U6904 (N_6904,N_4652,N_3827);
nor U6905 (N_6905,N_4591,N_2933);
xnor U6906 (N_6906,N_2714,N_3787);
nand U6907 (N_6907,N_4941,N_4587);
or U6908 (N_6908,N_3220,N_4467);
xnor U6909 (N_6909,N_3164,N_4272);
or U6910 (N_6910,N_3309,N_3907);
nor U6911 (N_6911,N_3520,N_4794);
or U6912 (N_6912,N_4268,N_3162);
and U6913 (N_6913,N_3476,N_3295);
or U6914 (N_6914,N_4396,N_4270);
or U6915 (N_6915,N_3018,N_4264);
nor U6916 (N_6916,N_4726,N_4186);
nor U6917 (N_6917,N_4666,N_2648);
nand U6918 (N_6918,N_2518,N_4396);
nor U6919 (N_6919,N_2879,N_2731);
or U6920 (N_6920,N_2877,N_4519);
or U6921 (N_6921,N_4023,N_4878);
or U6922 (N_6922,N_2764,N_4350);
xnor U6923 (N_6923,N_2626,N_3433);
and U6924 (N_6924,N_3034,N_3984);
nand U6925 (N_6925,N_4727,N_3828);
nand U6926 (N_6926,N_3678,N_3359);
and U6927 (N_6927,N_2874,N_3432);
and U6928 (N_6928,N_4337,N_4478);
or U6929 (N_6929,N_2879,N_3247);
or U6930 (N_6930,N_3934,N_2596);
nor U6931 (N_6931,N_2895,N_4730);
nor U6932 (N_6932,N_2626,N_4859);
and U6933 (N_6933,N_4860,N_4474);
and U6934 (N_6934,N_4467,N_3442);
or U6935 (N_6935,N_4235,N_4782);
nand U6936 (N_6936,N_3398,N_2749);
nand U6937 (N_6937,N_3663,N_3131);
nand U6938 (N_6938,N_3529,N_2546);
and U6939 (N_6939,N_3592,N_4365);
and U6940 (N_6940,N_2796,N_2660);
and U6941 (N_6941,N_3555,N_4812);
nor U6942 (N_6942,N_3782,N_4856);
or U6943 (N_6943,N_2675,N_3760);
and U6944 (N_6944,N_3090,N_2650);
and U6945 (N_6945,N_3774,N_4687);
or U6946 (N_6946,N_4611,N_3523);
and U6947 (N_6947,N_2920,N_4915);
nand U6948 (N_6948,N_3578,N_3248);
nand U6949 (N_6949,N_3826,N_4269);
and U6950 (N_6950,N_3117,N_4124);
or U6951 (N_6951,N_4014,N_2946);
or U6952 (N_6952,N_3905,N_2676);
or U6953 (N_6953,N_3248,N_2709);
nor U6954 (N_6954,N_4101,N_3901);
and U6955 (N_6955,N_2816,N_3926);
or U6956 (N_6956,N_2913,N_2543);
or U6957 (N_6957,N_4912,N_4264);
or U6958 (N_6958,N_2621,N_2742);
and U6959 (N_6959,N_3171,N_4195);
and U6960 (N_6960,N_2777,N_4668);
and U6961 (N_6961,N_3488,N_2716);
nor U6962 (N_6962,N_3270,N_3988);
nor U6963 (N_6963,N_4141,N_4263);
nand U6964 (N_6964,N_2698,N_3982);
or U6965 (N_6965,N_3599,N_3168);
and U6966 (N_6966,N_4995,N_3906);
nor U6967 (N_6967,N_3934,N_2769);
nand U6968 (N_6968,N_3939,N_2604);
nor U6969 (N_6969,N_3454,N_3846);
and U6970 (N_6970,N_3681,N_4307);
and U6971 (N_6971,N_4252,N_3501);
and U6972 (N_6972,N_4030,N_2779);
or U6973 (N_6973,N_3666,N_4488);
and U6974 (N_6974,N_3004,N_4227);
and U6975 (N_6975,N_3374,N_4146);
nand U6976 (N_6976,N_3047,N_3938);
and U6977 (N_6977,N_3615,N_4934);
and U6978 (N_6978,N_4362,N_3127);
nand U6979 (N_6979,N_3184,N_3913);
and U6980 (N_6980,N_3501,N_4832);
or U6981 (N_6981,N_2927,N_3780);
nor U6982 (N_6982,N_3211,N_2942);
nor U6983 (N_6983,N_3214,N_3989);
or U6984 (N_6984,N_4670,N_4441);
or U6985 (N_6985,N_4806,N_4670);
xnor U6986 (N_6986,N_2678,N_2850);
and U6987 (N_6987,N_4521,N_2574);
or U6988 (N_6988,N_4404,N_3885);
or U6989 (N_6989,N_3071,N_4179);
and U6990 (N_6990,N_2686,N_4468);
or U6991 (N_6991,N_4889,N_3812);
nor U6992 (N_6992,N_3772,N_3324);
and U6993 (N_6993,N_4376,N_4203);
nand U6994 (N_6994,N_2579,N_3909);
or U6995 (N_6995,N_4795,N_2765);
nor U6996 (N_6996,N_4311,N_4733);
or U6997 (N_6997,N_3809,N_4932);
and U6998 (N_6998,N_2937,N_3198);
and U6999 (N_6999,N_2522,N_4901);
nor U7000 (N_7000,N_2986,N_4554);
nand U7001 (N_7001,N_2927,N_4098);
or U7002 (N_7002,N_4178,N_4244);
and U7003 (N_7003,N_4949,N_2828);
nand U7004 (N_7004,N_4942,N_3560);
or U7005 (N_7005,N_2512,N_2535);
or U7006 (N_7006,N_3248,N_3142);
or U7007 (N_7007,N_3902,N_4919);
nand U7008 (N_7008,N_4660,N_4701);
nand U7009 (N_7009,N_2949,N_4884);
xnor U7010 (N_7010,N_4598,N_3215);
or U7011 (N_7011,N_4891,N_2919);
or U7012 (N_7012,N_4797,N_3198);
nand U7013 (N_7013,N_2968,N_2750);
nand U7014 (N_7014,N_3950,N_4455);
nor U7015 (N_7015,N_3029,N_3222);
or U7016 (N_7016,N_4742,N_4502);
or U7017 (N_7017,N_2509,N_3585);
nand U7018 (N_7018,N_2580,N_3854);
nand U7019 (N_7019,N_4080,N_3884);
and U7020 (N_7020,N_4220,N_2927);
nand U7021 (N_7021,N_4532,N_3510);
or U7022 (N_7022,N_3164,N_3142);
nor U7023 (N_7023,N_3518,N_3574);
and U7024 (N_7024,N_3575,N_4729);
and U7025 (N_7025,N_2975,N_4453);
or U7026 (N_7026,N_2829,N_3282);
or U7027 (N_7027,N_3506,N_2899);
nor U7028 (N_7028,N_4582,N_4648);
or U7029 (N_7029,N_2840,N_4734);
nor U7030 (N_7030,N_4418,N_4163);
nor U7031 (N_7031,N_3526,N_2856);
nor U7032 (N_7032,N_3044,N_4219);
and U7033 (N_7033,N_3446,N_2714);
nand U7034 (N_7034,N_2717,N_4092);
and U7035 (N_7035,N_3027,N_3387);
and U7036 (N_7036,N_4543,N_3039);
nand U7037 (N_7037,N_4347,N_4894);
or U7038 (N_7038,N_4806,N_4957);
nor U7039 (N_7039,N_4445,N_4215);
xnor U7040 (N_7040,N_3120,N_3575);
nor U7041 (N_7041,N_3194,N_4713);
nand U7042 (N_7042,N_3854,N_2944);
nand U7043 (N_7043,N_4153,N_2868);
or U7044 (N_7044,N_2551,N_4668);
nand U7045 (N_7045,N_3600,N_2632);
nand U7046 (N_7046,N_2845,N_2510);
nand U7047 (N_7047,N_4602,N_4089);
and U7048 (N_7048,N_4718,N_4750);
and U7049 (N_7049,N_2598,N_4806);
or U7050 (N_7050,N_4559,N_3698);
and U7051 (N_7051,N_4899,N_2641);
nand U7052 (N_7052,N_4828,N_4045);
or U7053 (N_7053,N_3075,N_2736);
and U7054 (N_7054,N_4650,N_4421);
nand U7055 (N_7055,N_3941,N_3761);
nand U7056 (N_7056,N_4054,N_3350);
and U7057 (N_7057,N_3941,N_2840);
nand U7058 (N_7058,N_3511,N_3999);
nor U7059 (N_7059,N_3549,N_3385);
nor U7060 (N_7060,N_3045,N_3048);
or U7061 (N_7061,N_3474,N_4595);
nor U7062 (N_7062,N_2565,N_2898);
nand U7063 (N_7063,N_3431,N_2531);
nand U7064 (N_7064,N_2520,N_4120);
or U7065 (N_7065,N_2738,N_4556);
nor U7066 (N_7066,N_4089,N_3458);
or U7067 (N_7067,N_4290,N_3818);
nor U7068 (N_7068,N_4128,N_4883);
nand U7069 (N_7069,N_4268,N_4602);
or U7070 (N_7070,N_2671,N_3309);
and U7071 (N_7071,N_4729,N_3493);
nand U7072 (N_7072,N_3400,N_3960);
and U7073 (N_7073,N_4918,N_2577);
nor U7074 (N_7074,N_2816,N_4961);
or U7075 (N_7075,N_2554,N_3422);
and U7076 (N_7076,N_3650,N_2853);
or U7077 (N_7077,N_2613,N_2572);
nor U7078 (N_7078,N_4852,N_3118);
and U7079 (N_7079,N_3758,N_2594);
and U7080 (N_7080,N_4855,N_3234);
or U7081 (N_7081,N_2870,N_4418);
nand U7082 (N_7082,N_3254,N_3878);
nand U7083 (N_7083,N_2648,N_4460);
xor U7084 (N_7084,N_3854,N_2584);
nand U7085 (N_7085,N_4759,N_3170);
and U7086 (N_7086,N_2917,N_3122);
and U7087 (N_7087,N_2961,N_2804);
nor U7088 (N_7088,N_4662,N_3252);
nor U7089 (N_7089,N_3907,N_3634);
or U7090 (N_7090,N_3659,N_2565);
nand U7091 (N_7091,N_3990,N_3609);
and U7092 (N_7092,N_3229,N_3649);
and U7093 (N_7093,N_4566,N_3230);
and U7094 (N_7094,N_3258,N_4806);
nand U7095 (N_7095,N_4468,N_4331);
and U7096 (N_7096,N_3609,N_4343);
or U7097 (N_7097,N_3609,N_4241);
and U7098 (N_7098,N_3219,N_3774);
nand U7099 (N_7099,N_4401,N_3520);
and U7100 (N_7100,N_3215,N_3528);
nand U7101 (N_7101,N_2874,N_4599);
or U7102 (N_7102,N_2712,N_2663);
or U7103 (N_7103,N_2779,N_2770);
or U7104 (N_7104,N_3457,N_4784);
nor U7105 (N_7105,N_3721,N_3744);
nand U7106 (N_7106,N_2996,N_3638);
nand U7107 (N_7107,N_4226,N_3594);
nand U7108 (N_7108,N_4798,N_3269);
or U7109 (N_7109,N_3247,N_4341);
and U7110 (N_7110,N_4887,N_2656);
or U7111 (N_7111,N_3155,N_2998);
nand U7112 (N_7112,N_4167,N_4263);
nor U7113 (N_7113,N_2923,N_3199);
or U7114 (N_7114,N_4717,N_3784);
and U7115 (N_7115,N_3412,N_4173);
and U7116 (N_7116,N_3730,N_4645);
nand U7117 (N_7117,N_3447,N_3040);
nand U7118 (N_7118,N_4315,N_4871);
nand U7119 (N_7119,N_3845,N_2771);
or U7120 (N_7120,N_4837,N_4018);
and U7121 (N_7121,N_2713,N_4928);
nand U7122 (N_7122,N_2951,N_4853);
or U7123 (N_7123,N_2552,N_2921);
nand U7124 (N_7124,N_3998,N_4650);
nor U7125 (N_7125,N_3742,N_4276);
and U7126 (N_7126,N_4506,N_3751);
or U7127 (N_7127,N_4484,N_4381);
xor U7128 (N_7128,N_3932,N_2817);
nor U7129 (N_7129,N_4938,N_3471);
or U7130 (N_7130,N_2648,N_4808);
and U7131 (N_7131,N_4055,N_2980);
nor U7132 (N_7132,N_4642,N_3086);
xnor U7133 (N_7133,N_4722,N_4894);
and U7134 (N_7134,N_2915,N_2503);
nand U7135 (N_7135,N_4076,N_4025);
nand U7136 (N_7136,N_3047,N_4315);
nor U7137 (N_7137,N_3628,N_2790);
and U7138 (N_7138,N_4660,N_3292);
nand U7139 (N_7139,N_4273,N_3637);
nand U7140 (N_7140,N_3542,N_4031);
and U7141 (N_7141,N_3005,N_3965);
and U7142 (N_7142,N_3179,N_2703);
or U7143 (N_7143,N_4555,N_3729);
and U7144 (N_7144,N_3686,N_4496);
or U7145 (N_7145,N_4315,N_3740);
nand U7146 (N_7146,N_2840,N_3537);
nor U7147 (N_7147,N_2912,N_4112);
or U7148 (N_7148,N_3772,N_4501);
nand U7149 (N_7149,N_3456,N_4999);
nand U7150 (N_7150,N_3235,N_4294);
and U7151 (N_7151,N_2997,N_4782);
nand U7152 (N_7152,N_3491,N_2872);
and U7153 (N_7153,N_3641,N_2938);
nand U7154 (N_7154,N_3751,N_3889);
xnor U7155 (N_7155,N_4838,N_2888);
nand U7156 (N_7156,N_4593,N_4153);
or U7157 (N_7157,N_3510,N_2718);
nor U7158 (N_7158,N_3201,N_3867);
nor U7159 (N_7159,N_2519,N_3077);
or U7160 (N_7160,N_4191,N_2504);
nand U7161 (N_7161,N_2820,N_4331);
nor U7162 (N_7162,N_4791,N_2956);
nand U7163 (N_7163,N_3373,N_2670);
or U7164 (N_7164,N_2747,N_3970);
xnor U7165 (N_7165,N_4195,N_4983);
nand U7166 (N_7166,N_2852,N_4206);
nand U7167 (N_7167,N_3024,N_4245);
nor U7168 (N_7168,N_3454,N_3574);
nor U7169 (N_7169,N_4437,N_3074);
nand U7170 (N_7170,N_3071,N_2830);
and U7171 (N_7171,N_2559,N_2534);
nand U7172 (N_7172,N_3424,N_2600);
and U7173 (N_7173,N_4085,N_2750);
nand U7174 (N_7174,N_2961,N_2785);
and U7175 (N_7175,N_3807,N_3035);
and U7176 (N_7176,N_3121,N_3351);
or U7177 (N_7177,N_2887,N_4841);
nor U7178 (N_7178,N_4884,N_3034);
or U7179 (N_7179,N_4831,N_4326);
and U7180 (N_7180,N_2666,N_3913);
or U7181 (N_7181,N_3526,N_3621);
and U7182 (N_7182,N_3623,N_3775);
and U7183 (N_7183,N_3431,N_4778);
nor U7184 (N_7184,N_4729,N_2788);
nand U7185 (N_7185,N_4407,N_2904);
and U7186 (N_7186,N_2618,N_4589);
or U7187 (N_7187,N_4767,N_2739);
or U7188 (N_7188,N_3118,N_4822);
nand U7189 (N_7189,N_4525,N_2975);
or U7190 (N_7190,N_4927,N_4477);
and U7191 (N_7191,N_2741,N_4206);
or U7192 (N_7192,N_2788,N_3387);
or U7193 (N_7193,N_3836,N_3410);
nor U7194 (N_7194,N_2634,N_4019);
and U7195 (N_7195,N_4093,N_2804);
and U7196 (N_7196,N_3577,N_4541);
and U7197 (N_7197,N_2579,N_3809);
and U7198 (N_7198,N_2967,N_3606);
and U7199 (N_7199,N_2793,N_4362);
nand U7200 (N_7200,N_4705,N_3673);
and U7201 (N_7201,N_3826,N_4699);
nand U7202 (N_7202,N_4903,N_3986);
nor U7203 (N_7203,N_4898,N_2656);
nand U7204 (N_7204,N_2915,N_4021);
and U7205 (N_7205,N_2876,N_4832);
or U7206 (N_7206,N_4296,N_3929);
and U7207 (N_7207,N_2526,N_3475);
and U7208 (N_7208,N_4551,N_3896);
and U7209 (N_7209,N_4754,N_4554);
xor U7210 (N_7210,N_3315,N_4976);
and U7211 (N_7211,N_4936,N_3082);
or U7212 (N_7212,N_3576,N_2719);
and U7213 (N_7213,N_4617,N_3310);
or U7214 (N_7214,N_4648,N_4686);
and U7215 (N_7215,N_2910,N_4461);
nor U7216 (N_7216,N_3461,N_4470);
nor U7217 (N_7217,N_2960,N_3444);
nor U7218 (N_7218,N_4113,N_4998);
nand U7219 (N_7219,N_4737,N_4515);
or U7220 (N_7220,N_3271,N_3868);
nand U7221 (N_7221,N_4955,N_2975);
nor U7222 (N_7222,N_4865,N_4573);
nand U7223 (N_7223,N_3222,N_4648);
and U7224 (N_7224,N_4306,N_4093);
or U7225 (N_7225,N_2798,N_3329);
nor U7226 (N_7226,N_4944,N_3933);
nand U7227 (N_7227,N_3784,N_4658);
nor U7228 (N_7228,N_4089,N_3635);
nor U7229 (N_7229,N_4336,N_4998);
nand U7230 (N_7230,N_3265,N_4471);
nand U7231 (N_7231,N_3756,N_2787);
and U7232 (N_7232,N_2967,N_4386);
nand U7233 (N_7233,N_3664,N_4648);
nor U7234 (N_7234,N_2504,N_3214);
nor U7235 (N_7235,N_2868,N_2960);
nor U7236 (N_7236,N_3452,N_2975);
or U7237 (N_7237,N_3348,N_3525);
nand U7238 (N_7238,N_4162,N_4844);
nand U7239 (N_7239,N_3353,N_3595);
nor U7240 (N_7240,N_4292,N_3891);
nand U7241 (N_7241,N_2733,N_3251);
nand U7242 (N_7242,N_3049,N_4147);
or U7243 (N_7243,N_3632,N_4926);
nor U7244 (N_7244,N_2988,N_4785);
and U7245 (N_7245,N_3489,N_3761);
nand U7246 (N_7246,N_4673,N_2809);
and U7247 (N_7247,N_2670,N_2604);
nor U7248 (N_7248,N_2957,N_2988);
nand U7249 (N_7249,N_3854,N_4905);
or U7250 (N_7250,N_3152,N_4101);
and U7251 (N_7251,N_2861,N_4483);
or U7252 (N_7252,N_3079,N_3667);
nand U7253 (N_7253,N_3429,N_3932);
and U7254 (N_7254,N_2734,N_3491);
nor U7255 (N_7255,N_4260,N_4953);
nand U7256 (N_7256,N_3721,N_3560);
or U7257 (N_7257,N_3374,N_3300);
nand U7258 (N_7258,N_4308,N_3477);
nor U7259 (N_7259,N_2654,N_4853);
or U7260 (N_7260,N_4720,N_4943);
nand U7261 (N_7261,N_4880,N_3775);
nor U7262 (N_7262,N_2965,N_3612);
xnor U7263 (N_7263,N_3571,N_4858);
nor U7264 (N_7264,N_3504,N_2535);
nand U7265 (N_7265,N_3016,N_3002);
or U7266 (N_7266,N_2563,N_3777);
nand U7267 (N_7267,N_2685,N_3394);
and U7268 (N_7268,N_3339,N_4402);
or U7269 (N_7269,N_2905,N_3272);
and U7270 (N_7270,N_2879,N_3592);
and U7271 (N_7271,N_3216,N_3369);
nand U7272 (N_7272,N_3217,N_4809);
nor U7273 (N_7273,N_3773,N_3139);
nor U7274 (N_7274,N_3452,N_3613);
xor U7275 (N_7275,N_4259,N_4489);
or U7276 (N_7276,N_3011,N_3901);
nand U7277 (N_7277,N_4480,N_2952);
nor U7278 (N_7278,N_4834,N_4686);
or U7279 (N_7279,N_4852,N_3683);
or U7280 (N_7280,N_3367,N_3652);
nor U7281 (N_7281,N_3813,N_3108);
or U7282 (N_7282,N_3155,N_4540);
nor U7283 (N_7283,N_4858,N_4013);
nand U7284 (N_7284,N_3586,N_3067);
and U7285 (N_7285,N_2903,N_3842);
nand U7286 (N_7286,N_3683,N_3669);
nand U7287 (N_7287,N_3845,N_4248);
nor U7288 (N_7288,N_2702,N_3562);
xor U7289 (N_7289,N_2709,N_2541);
or U7290 (N_7290,N_3475,N_3012);
nor U7291 (N_7291,N_2843,N_3008);
nand U7292 (N_7292,N_4159,N_4651);
or U7293 (N_7293,N_3928,N_3366);
nand U7294 (N_7294,N_4715,N_3172);
xnor U7295 (N_7295,N_3836,N_3433);
nor U7296 (N_7296,N_3025,N_2887);
and U7297 (N_7297,N_3512,N_3282);
or U7298 (N_7298,N_4615,N_4342);
or U7299 (N_7299,N_4842,N_3647);
and U7300 (N_7300,N_4069,N_3228);
and U7301 (N_7301,N_4689,N_4822);
and U7302 (N_7302,N_3266,N_4838);
nand U7303 (N_7303,N_3782,N_2552);
nor U7304 (N_7304,N_4741,N_4675);
xnor U7305 (N_7305,N_2812,N_4991);
nor U7306 (N_7306,N_4532,N_4983);
and U7307 (N_7307,N_3595,N_2991);
nand U7308 (N_7308,N_2687,N_2715);
nor U7309 (N_7309,N_4881,N_2561);
and U7310 (N_7310,N_4443,N_4315);
nand U7311 (N_7311,N_2544,N_2715);
xor U7312 (N_7312,N_4391,N_4489);
and U7313 (N_7313,N_3662,N_3570);
nor U7314 (N_7314,N_4745,N_4040);
or U7315 (N_7315,N_3817,N_3031);
nand U7316 (N_7316,N_4921,N_4914);
nand U7317 (N_7317,N_4167,N_4893);
nand U7318 (N_7318,N_3727,N_4249);
or U7319 (N_7319,N_4042,N_4801);
nor U7320 (N_7320,N_3186,N_3453);
and U7321 (N_7321,N_4267,N_3160);
and U7322 (N_7322,N_2683,N_4335);
nor U7323 (N_7323,N_2590,N_4534);
nand U7324 (N_7324,N_4556,N_3897);
or U7325 (N_7325,N_2941,N_4489);
nand U7326 (N_7326,N_4513,N_4952);
nand U7327 (N_7327,N_2883,N_4386);
and U7328 (N_7328,N_2644,N_3403);
nand U7329 (N_7329,N_4834,N_4934);
nor U7330 (N_7330,N_4709,N_2609);
or U7331 (N_7331,N_3359,N_4132);
nor U7332 (N_7332,N_4547,N_4037);
nand U7333 (N_7333,N_4856,N_3846);
and U7334 (N_7334,N_2627,N_3558);
nand U7335 (N_7335,N_3279,N_2822);
nand U7336 (N_7336,N_4072,N_4515);
nor U7337 (N_7337,N_3399,N_4318);
nor U7338 (N_7338,N_2914,N_4784);
nor U7339 (N_7339,N_3922,N_4198);
or U7340 (N_7340,N_4078,N_4164);
nand U7341 (N_7341,N_2501,N_4870);
or U7342 (N_7342,N_3402,N_4747);
nand U7343 (N_7343,N_3285,N_4835);
nor U7344 (N_7344,N_4576,N_2938);
or U7345 (N_7345,N_4034,N_4325);
nor U7346 (N_7346,N_2547,N_3850);
and U7347 (N_7347,N_4670,N_4534);
nor U7348 (N_7348,N_4374,N_4858);
nand U7349 (N_7349,N_3442,N_2607);
and U7350 (N_7350,N_2588,N_4120);
and U7351 (N_7351,N_3045,N_4580);
or U7352 (N_7352,N_4300,N_4748);
nand U7353 (N_7353,N_4377,N_2817);
nand U7354 (N_7354,N_3566,N_2752);
and U7355 (N_7355,N_2908,N_2566);
nor U7356 (N_7356,N_4249,N_4601);
nand U7357 (N_7357,N_4054,N_3611);
nor U7358 (N_7358,N_3302,N_2653);
and U7359 (N_7359,N_3423,N_2692);
or U7360 (N_7360,N_4771,N_3459);
nor U7361 (N_7361,N_4435,N_2677);
nor U7362 (N_7362,N_3580,N_3611);
or U7363 (N_7363,N_3247,N_4988);
nor U7364 (N_7364,N_2756,N_2507);
and U7365 (N_7365,N_2624,N_2836);
nor U7366 (N_7366,N_2799,N_3764);
or U7367 (N_7367,N_3397,N_3738);
nand U7368 (N_7368,N_2847,N_2880);
and U7369 (N_7369,N_3191,N_3823);
and U7370 (N_7370,N_4156,N_3559);
nor U7371 (N_7371,N_3851,N_3931);
nor U7372 (N_7372,N_2827,N_4216);
and U7373 (N_7373,N_3446,N_4212);
and U7374 (N_7374,N_3608,N_4100);
and U7375 (N_7375,N_4556,N_3027);
and U7376 (N_7376,N_4081,N_3558);
and U7377 (N_7377,N_3427,N_3346);
or U7378 (N_7378,N_3365,N_4905);
nor U7379 (N_7379,N_4776,N_4628);
or U7380 (N_7380,N_4458,N_4270);
and U7381 (N_7381,N_4106,N_4074);
nand U7382 (N_7382,N_3376,N_4355);
nand U7383 (N_7383,N_2618,N_2581);
nand U7384 (N_7384,N_4659,N_4186);
nor U7385 (N_7385,N_2666,N_3954);
or U7386 (N_7386,N_4594,N_3406);
nand U7387 (N_7387,N_3259,N_3159);
and U7388 (N_7388,N_4877,N_4796);
nand U7389 (N_7389,N_3243,N_3002);
nor U7390 (N_7390,N_3881,N_2665);
nor U7391 (N_7391,N_2653,N_2998);
or U7392 (N_7392,N_3065,N_3112);
nand U7393 (N_7393,N_3595,N_3112);
and U7394 (N_7394,N_4648,N_2848);
and U7395 (N_7395,N_3496,N_3462);
nand U7396 (N_7396,N_4624,N_2817);
or U7397 (N_7397,N_3204,N_3297);
and U7398 (N_7398,N_4369,N_3321);
nand U7399 (N_7399,N_4682,N_3429);
or U7400 (N_7400,N_4656,N_4953);
nor U7401 (N_7401,N_4715,N_4601);
and U7402 (N_7402,N_3908,N_3363);
nor U7403 (N_7403,N_4404,N_4281);
xor U7404 (N_7404,N_3631,N_3677);
or U7405 (N_7405,N_2946,N_4507);
and U7406 (N_7406,N_3165,N_3962);
or U7407 (N_7407,N_2757,N_2882);
and U7408 (N_7408,N_4428,N_3275);
or U7409 (N_7409,N_4079,N_4768);
nand U7410 (N_7410,N_4716,N_2868);
nor U7411 (N_7411,N_3488,N_4065);
nand U7412 (N_7412,N_3108,N_3238);
and U7413 (N_7413,N_2647,N_3247);
nand U7414 (N_7414,N_4604,N_4832);
and U7415 (N_7415,N_3955,N_3265);
or U7416 (N_7416,N_3267,N_4999);
and U7417 (N_7417,N_4454,N_4705);
xnor U7418 (N_7418,N_2623,N_4749);
and U7419 (N_7419,N_3181,N_3994);
nor U7420 (N_7420,N_4317,N_4034);
nor U7421 (N_7421,N_4660,N_4170);
nor U7422 (N_7422,N_2898,N_4484);
nor U7423 (N_7423,N_2890,N_4250);
nand U7424 (N_7424,N_3957,N_3610);
or U7425 (N_7425,N_4488,N_3490);
nor U7426 (N_7426,N_4447,N_3344);
nand U7427 (N_7427,N_3656,N_4583);
nand U7428 (N_7428,N_2933,N_3717);
nand U7429 (N_7429,N_2924,N_4076);
or U7430 (N_7430,N_3024,N_3309);
nor U7431 (N_7431,N_4534,N_2810);
nand U7432 (N_7432,N_3979,N_4034);
and U7433 (N_7433,N_4945,N_4622);
and U7434 (N_7434,N_4854,N_4108);
or U7435 (N_7435,N_4294,N_2643);
nor U7436 (N_7436,N_3675,N_2823);
nand U7437 (N_7437,N_3330,N_3414);
and U7438 (N_7438,N_2707,N_2846);
nand U7439 (N_7439,N_3388,N_3054);
and U7440 (N_7440,N_3485,N_3043);
and U7441 (N_7441,N_4260,N_2627);
or U7442 (N_7442,N_4687,N_3967);
xor U7443 (N_7443,N_3746,N_2612);
or U7444 (N_7444,N_3570,N_3858);
nor U7445 (N_7445,N_3550,N_4883);
and U7446 (N_7446,N_3835,N_3595);
and U7447 (N_7447,N_3811,N_3229);
or U7448 (N_7448,N_3421,N_4226);
nand U7449 (N_7449,N_4323,N_4687);
or U7450 (N_7450,N_4964,N_3398);
nor U7451 (N_7451,N_3329,N_3310);
nand U7452 (N_7452,N_3522,N_4654);
nand U7453 (N_7453,N_3808,N_2611);
nand U7454 (N_7454,N_4645,N_4423);
nand U7455 (N_7455,N_3649,N_4016);
and U7456 (N_7456,N_3665,N_4108);
and U7457 (N_7457,N_4351,N_4922);
nor U7458 (N_7458,N_3354,N_2729);
nor U7459 (N_7459,N_2768,N_4148);
or U7460 (N_7460,N_4234,N_2598);
nand U7461 (N_7461,N_3038,N_4068);
and U7462 (N_7462,N_2890,N_4295);
and U7463 (N_7463,N_3043,N_3164);
nor U7464 (N_7464,N_4531,N_4858);
nand U7465 (N_7465,N_3059,N_4639);
nand U7466 (N_7466,N_3031,N_4615);
or U7467 (N_7467,N_4092,N_3264);
or U7468 (N_7468,N_4757,N_3519);
or U7469 (N_7469,N_3291,N_3593);
and U7470 (N_7470,N_2937,N_3951);
and U7471 (N_7471,N_2900,N_2747);
or U7472 (N_7472,N_4115,N_3115);
nor U7473 (N_7473,N_3250,N_2762);
nor U7474 (N_7474,N_3634,N_3475);
nor U7475 (N_7475,N_4468,N_3733);
nand U7476 (N_7476,N_3736,N_3848);
nor U7477 (N_7477,N_4063,N_4716);
nor U7478 (N_7478,N_4037,N_2622);
nor U7479 (N_7479,N_3855,N_3171);
nor U7480 (N_7480,N_3366,N_3234);
nand U7481 (N_7481,N_2976,N_3653);
nor U7482 (N_7482,N_4029,N_4615);
nand U7483 (N_7483,N_3863,N_3186);
nand U7484 (N_7484,N_4328,N_4659);
nor U7485 (N_7485,N_2821,N_2698);
or U7486 (N_7486,N_4050,N_3943);
nand U7487 (N_7487,N_2611,N_4863);
and U7488 (N_7488,N_3554,N_2549);
nor U7489 (N_7489,N_4691,N_2990);
and U7490 (N_7490,N_2645,N_4153);
and U7491 (N_7491,N_3163,N_3629);
nor U7492 (N_7492,N_3543,N_3878);
nor U7493 (N_7493,N_3619,N_3411);
and U7494 (N_7494,N_3713,N_3424);
nand U7495 (N_7495,N_3639,N_2894);
nor U7496 (N_7496,N_3623,N_2948);
nor U7497 (N_7497,N_2916,N_4639);
and U7498 (N_7498,N_3258,N_3840);
and U7499 (N_7499,N_3512,N_3261);
nor U7500 (N_7500,N_5751,N_6267);
or U7501 (N_7501,N_5122,N_6899);
nor U7502 (N_7502,N_6600,N_5794);
nor U7503 (N_7503,N_5601,N_6652);
nand U7504 (N_7504,N_6726,N_5205);
nor U7505 (N_7505,N_6729,N_6614);
nor U7506 (N_7506,N_6035,N_6367);
nor U7507 (N_7507,N_6002,N_6365);
and U7508 (N_7508,N_7052,N_5088);
nor U7509 (N_7509,N_6366,N_7144);
or U7510 (N_7510,N_6655,N_6838);
nand U7511 (N_7511,N_5425,N_6373);
or U7512 (N_7512,N_5333,N_6973);
and U7513 (N_7513,N_5991,N_5606);
nand U7514 (N_7514,N_7388,N_5298);
or U7515 (N_7515,N_5743,N_7016);
nand U7516 (N_7516,N_7148,N_5220);
and U7517 (N_7517,N_5550,N_6124);
nor U7518 (N_7518,N_7230,N_5233);
nand U7519 (N_7519,N_7385,N_6402);
nor U7520 (N_7520,N_6239,N_7464);
and U7521 (N_7521,N_5157,N_5741);
xnor U7522 (N_7522,N_5130,N_5961);
and U7523 (N_7523,N_6480,N_6881);
xnor U7524 (N_7524,N_6371,N_7374);
and U7525 (N_7525,N_7287,N_6242);
nand U7526 (N_7526,N_6471,N_5868);
and U7527 (N_7527,N_5717,N_7219);
nor U7528 (N_7528,N_5624,N_7102);
or U7529 (N_7529,N_5109,N_5043);
xor U7530 (N_7530,N_5324,N_5971);
nand U7531 (N_7531,N_5163,N_5642);
or U7532 (N_7532,N_5394,N_7140);
nand U7533 (N_7533,N_5870,N_6657);
nor U7534 (N_7534,N_5716,N_6406);
and U7535 (N_7535,N_5808,N_7400);
nand U7536 (N_7536,N_5223,N_7019);
xor U7537 (N_7537,N_6725,N_7261);
nor U7538 (N_7538,N_7014,N_7325);
nand U7539 (N_7539,N_5629,N_6268);
nor U7540 (N_7540,N_5346,N_5029);
nor U7541 (N_7541,N_6063,N_6156);
or U7542 (N_7542,N_5709,N_5864);
nor U7543 (N_7543,N_5761,N_6615);
and U7544 (N_7544,N_5231,N_5575);
and U7545 (N_7545,N_6562,N_6601);
or U7546 (N_7546,N_7168,N_5781);
nor U7547 (N_7547,N_5668,N_6554);
nand U7548 (N_7548,N_5962,N_5616);
or U7549 (N_7549,N_7130,N_6887);
and U7550 (N_7550,N_6428,N_6689);
nor U7551 (N_7551,N_5318,N_7202);
nand U7552 (N_7552,N_6344,N_5738);
or U7553 (N_7553,N_6651,N_6106);
nand U7554 (N_7554,N_5327,N_7236);
or U7555 (N_7555,N_6741,N_5412);
or U7556 (N_7556,N_6000,N_5311);
nor U7557 (N_7557,N_7250,N_6575);
nor U7558 (N_7558,N_7440,N_6003);
nand U7559 (N_7559,N_5909,N_5025);
nor U7560 (N_7560,N_6164,N_6686);
xor U7561 (N_7561,N_5368,N_5496);
xor U7562 (N_7562,N_5865,N_6389);
and U7563 (N_7563,N_5524,N_6151);
and U7564 (N_7564,N_6841,N_7496);
or U7565 (N_7565,N_5871,N_5982);
nor U7566 (N_7566,N_7387,N_6659);
nand U7567 (N_7567,N_5734,N_6360);
nand U7568 (N_7568,N_7193,N_5742);
or U7569 (N_7569,N_6456,N_5730);
nor U7570 (N_7570,N_6880,N_7286);
nand U7571 (N_7571,N_7311,N_5426);
and U7572 (N_7572,N_5521,N_6091);
nor U7573 (N_7573,N_7295,N_6611);
nand U7574 (N_7574,N_5973,N_5893);
xor U7575 (N_7575,N_6446,N_7483);
nand U7576 (N_7576,N_6265,N_5495);
and U7577 (N_7577,N_5546,N_7481);
nor U7578 (N_7578,N_6858,N_5446);
or U7579 (N_7579,N_6811,N_5490);
and U7580 (N_7580,N_5920,N_5753);
nand U7581 (N_7581,N_6102,N_6101);
nand U7582 (N_7582,N_6270,N_6177);
or U7583 (N_7583,N_6429,N_7376);
nand U7584 (N_7584,N_6421,N_7223);
or U7585 (N_7585,N_6308,N_7488);
nor U7586 (N_7586,N_7184,N_6044);
nand U7587 (N_7587,N_6178,N_7065);
nand U7588 (N_7588,N_6807,N_5792);
nor U7589 (N_7589,N_7313,N_6910);
nand U7590 (N_7590,N_5360,N_5643);
nor U7591 (N_7591,N_5699,N_7208);
nand U7592 (N_7592,N_5929,N_5778);
nand U7593 (N_7593,N_5478,N_7017);
nand U7594 (N_7594,N_5848,N_5613);
or U7595 (N_7595,N_6870,N_6381);
nor U7596 (N_7596,N_6412,N_6771);
or U7597 (N_7597,N_5283,N_5416);
and U7598 (N_7598,N_5802,N_6119);
nand U7599 (N_7599,N_5976,N_6587);
nand U7600 (N_7600,N_6081,N_5403);
xnor U7601 (N_7601,N_5434,N_6936);
nand U7602 (N_7602,N_5296,N_5193);
or U7603 (N_7603,N_5209,N_6136);
nor U7604 (N_7604,N_5051,N_5228);
nor U7605 (N_7605,N_6604,N_6410);
and U7606 (N_7606,N_6258,N_6801);
nor U7607 (N_7607,N_5352,N_6742);
xnor U7608 (N_7608,N_5070,N_5143);
and U7609 (N_7609,N_5072,N_5455);
and U7610 (N_7610,N_6219,N_6945);
and U7611 (N_7611,N_5115,N_5978);
and U7612 (N_7612,N_6922,N_5097);
or U7613 (N_7613,N_5469,N_6160);
nand U7614 (N_7614,N_5790,N_6276);
or U7615 (N_7615,N_5789,N_6162);
nand U7616 (N_7616,N_6279,N_6590);
or U7617 (N_7617,N_5650,N_5195);
and U7618 (N_7618,N_6730,N_5869);
nor U7619 (N_7619,N_7369,N_7039);
and U7620 (N_7620,N_5112,N_5138);
and U7621 (N_7621,N_6054,N_7162);
nand U7622 (N_7622,N_5128,N_6888);
nand U7623 (N_7623,N_5999,N_5652);
nand U7624 (N_7624,N_6161,N_6200);
nand U7625 (N_7625,N_7224,N_5161);
and U7626 (N_7626,N_5291,N_7431);
nand U7627 (N_7627,N_5366,N_6581);
nor U7628 (N_7628,N_6169,N_7106);
or U7629 (N_7629,N_5471,N_5382);
nand U7630 (N_7630,N_6301,N_5438);
and U7631 (N_7631,N_5987,N_6877);
nand U7632 (N_7632,N_5702,N_5242);
nor U7633 (N_7633,N_6719,N_6041);
nand U7634 (N_7634,N_7458,N_5451);
nor U7635 (N_7635,N_7046,N_6603);
nor U7636 (N_7636,N_5456,N_6721);
nor U7637 (N_7637,N_5441,N_7490);
or U7638 (N_7638,N_6008,N_6746);
nor U7639 (N_7639,N_7105,N_5019);
nand U7640 (N_7640,N_5306,N_7329);
nand U7641 (N_7641,N_6397,N_6089);
nor U7642 (N_7642,N_6364,N_5757);
or U7643 (N_7643,N_5281,N_6468);
nand U7644 (N_7644,N_7346,N_5911);
nand U7645 (N_7645,N_5289,N_6439);
and U7646 (N_7646,N_5907,N_6920);
and U7647 (N_7647,N_6690,N_5486);
nand U7648 (N_7648,N_5473,N_7421);
and U7649 (N_7649,N_7428,N_5940);
or U7650 (N_7650,N_6188,N_5439);
or U7651 (N_7651,N_6370,N_6049);
or U7652 (N_7652,N_6812,N_6891);
nor U7653 (N_7653,N_5856,N_6931);
or U7654 (N_7654,N_7343,N_6525);
or U7655 (N_7655,N_5960,N_7389);
xor U7656 (N_7656,N_7079,N_6324);
and U7657 (N_7657,N_7264,N_7284);
nor U7658 (N_7658,N_6249,N_6739);
or U7659 (N_7659,N_7354,N_6470);
xor U7660 (N_7660,N_5079,N_5218);
or U7661 (N_7661,N_5661,N_7394);
or U7662 (N_7662,N_6847,N_7439);
and U7663 (N_7663,N_7066,N_6745);
and U7664 (N_7664,N_7268,N_5357);
nor U7665 (N_7665,N_6213,N_6783);
nand U7666 (N_7666,N_6948,N_6459);
nor U7667 (N_7667,N_6758,N_6722);
nor U7668 (N_7668,N_7392,N_6304);
and U7669 (N_7669,N_5304,N_5227);
nor U7670 (N_7670,N_7175,N_6782);
nand U7671 (N_7671,N_6767,N_7301);
and U7672 (N_7672,N_5264,N_5934);
and U7673 (N_7673,N_5532,N_6806);
and U7674 (N_7674,N_5599,N_5012);
nand U7675 (N_7675,N_6735,N_6481);
and U7676 (N_7676,N_6499,N_5016);
nor U7677 (N_7677,N_5736,N_6254);
nor U7678 (N_7678,N_5234,N_5615);
and U7679 (N_7679,N_7060,N_5747);
nor U7680 (N_7680,N_6385,N_7338);
nor U7681 (N_7681,N_5877,N_5854);
and U7682 (N_7682,N_6039,N_5052);
nor U7683 (N_7683,N_5622,N_5817);
or U7684 (N_7684,N_6329,N_7018);
nor U7685 (N_7685,N_5312,N_7249);
or U7686 (N_7686,N_7429,N_5194);
nand U7687 (N_7687,N_6204,N_5090);
nand U7688 (N_7688,N_5140,N_6335);
and U7689 (N_7689,N_5832,N_5659);
nand U7690 (N_7690,N_7247,N_6997);
nor U7691 (N_7691,N_6768,N_6191);
nand U7692 (N_7692,N_6792,N_6504);
and U7693 (N_7693,N_7020,N_6430);
and U7694 (N_7694,N_5252,N_6498);
and U7695 (N_7695,N_7067,N_5913);
nor U7696 (N_7696,N_6065,N_6356);
nor U7697 (N_7697,N_6750,N_5073);
xnor U7698 (N_7698,N_6100,N_6307);
nor U7699 (N_7699,N_5968,N_6450);
or U7700 (N_7700,N_6999,N_5873);
and U7701 (N_7701,N_5400,N_7081);
or U7702 (N_7702,N_6048,N_5034);
nor U7703 (N_7703,N_5837,N_6814);
nand U7704 (N_7704,N_6112,N_5829);
nor U7705 (N_7705,N_5506,N_5388);
or U7706 (N_7706,N_6129,N_5901);
nor U7707 (N_7707,N_5764,N_6586);
nor U7708 (N_7708,N_6170,N_7234);
or U7709 (N_7709,N_5300,N_5098);
or U7710 (N_7710,N_7161,N_5621);
nor U7711 (N_7711,N_6157,N_6970);
and U7712 (N_7712,N_5767,N_5396);
or U7713 (N_7713,N_6789,N_5755);
nand U7714 (N_7714,N_6720,N_7266);
nand U7715 (N_7715,N_7372,N_5876);
nand U7716 (N_7716,N_7181,N_6336);
and U7717 (N_7717,N_5216,N_6103);
and U7718 (N_7718,N_5154,N_5891);
and U7719 (N_7719,N_6195,N_6140);
and U7720 (N_7720,N_5586,N_6666);
nor U7721 (N_7721,N_6946,N_7013);
nand U7722 (N_7722,N_7159,N_7221);
or U7723 (N_7723,N_5830,N_7258);
nor U7724 (N_7724,N_7408,N_6363);
and U7725 (N_7725,N_5551,N_5512);
nand U7726 (N_7726,N_6232,N_7073);
or U7727 (N_7727,N_5749,N_6663);
and U7728 (N_7728,N_5598,N_5579);
or U7729 (N_7729,N_6808,N_5503);
nor U7730 (N_7730,N_6055,N_5349);
or U7731 (N_7731,N_6082,N_6411);
nand U7732 (N_7732,N_6104,N_5574);
nor U7733 (N_7733,N_7356,N_5042);
or U7734 (N_7734,N_6211,N_7406);
and U7735 (N_7735,N_6701,N_5279);
nor U7736 (N_7736,N_5248,N_5656);
nor U7737 (N_7737,N_5383,N_6975);
or U7738 (N_7738,N_5492,N_6911);
and U7739 (N_7739,N_6951,N_6928);
and U7740 (N_7740,N_5822,N_5316);
nor U7741 (N_7741,N_5818,N_5545);
nand U7742 (N_7742,N_7164,N_6935);
nand U7743 (N_7743,N_6248,N_7152);
and U7744 (N_7744,N_7112,N_5099);
nand U7745 (N_7745,N_6833,N_6068);
and U7746 (N_7746,N_6486,N_5011);
or U7747 (N_7747,N_6202,N_5370);
and U7748 (N_7748,N_7195,N_7349);
and U7749 (N_7749,N_7333,N_5219);
and U7750 (N_7750,N_6705,N_6298);
nand U7751 (N_7751,N_5255,N_5898);
nand U7752 (N_7752,N_6774,N_7163);
and U7753 (N_7753,N_6455,N_5897);
and U7754 (N_7754,N_6541,N_7450);
nand U7755 (N_7755,N_5080,N_5113);
or U7756 (N_7756,N_6190,N_5750);
nor U7757 (N_7757,N_5703,N_6776);
nand U7758 (N_7758,N_6558,N_6185);
and U7759 (N_7759,N_6037,N_6872);
nand U7760 (N_7760,N_5697,N_5930);
nand U7761 (N_7761,N_7024,N_5430);
nor U7762 (N_7762,N_6293,N_7445);
or U7763 (N_7763,N_6264,N_6024);
nand U7764 (N_7764,N_7289,N_5733);
nand U7765 (N_7765,N_6777,N_6165);
nor U7766 (N_7766,N_5625,N_5827);
nand U7767 (N_7767,N_7364,N_5341);
nand U7768 (N_7768,N_6890,N_5254);
nand U7769 (N_7769,N_6377,N_7273);
or U7770 (N_7770,N_6475,N_5863);
nor U7771 (N_7771,N_7327,N_5995);
xor U7772 (N_7772,N_5124,N_5121);
and U7773 (N_7773,N_6284,N_6571);
and U7774 (N_7774,N_7393,N_6913);
or U7775 (N_7775,N_5297,N_6488);
nand U7776 (N_7776,N_6206,N_6597);
or U7777 (N_7777,N_5914,N_6023);
nor U7778 (N_7778,N_6795,N_5558);
and U7779 (N_7779,N_6095,N_7143);
and U7780 (N_7780,N_7326,N_5938);
and U7781 (N_7781,N_7368,N_5385);
nor U7782 (N_7782,N_7154,N_5942);
nand U7783 (N_7783,N_5384,N_5453);
and U7784 (N_7784,N_6013,N_5038);
and U7785 (N_7785,N_7272,N_5986);
nor U7786 (N_7786,N_5939,N_5239);
nor U7787 (N_7787,N_6493,N_6749);
nand U7788 (N_7788,N_6009,N_6821);
or U7789 (N_7789,N_5293,N_6660);
nor U7790 (N_7790,N_6226,N_5395);
or U7791 (N_7791,N_6633,N_5520);
nor U7792 (N_7792,N_7489,N_7413);
nor U7793 (N_7793,N_6531,N_7452);
nor U7794 (N_7794,N_6438,N_7379);
nand U7795 (N_7795,N_5107,N_7056);
or U7796 (N_7796,N_7128,N_6046);
and U7797 (N_7797,N_7075,N_6699);
and U7798 (N_7798,N_6275,N_5036);
or U7799 (N_7799,N_5513,N_6507);
nor U7800 (N_7800,N_6463,N_5049);
and U7801 (N_7801,N_5246,N_5762);
or U7802 (N_7802,N_6334,N_7253);
or U7803 (N_7803,N_6673,N_7142);
and U7804 (N_7804,N_5947,N_5782);
nand U7805 (N_7805,N_7321,N_6122);
nor U7806 (N_7806,N_5129,N_5258);
nand U7807 (N_7807,N_6339,N_7274);
nand U7808 (N_7808,N_7093,N_7475);
and U7809 (N_7809,N_6569,N_6793);
nand U7810 (N_7810,N_5603,N_6019);
and U7811 (N_7811,N_5531,N_6593);
nor U7812 (N_7812,N_5373,N_5746);
nor U7813 (N_7813,N_6754,N_6845);
xor U7814 (N_7814,N_6863,N_5890);
or U7815 (N_7815,N_7005,N_5718);
nor U7816 (N_7816,N_6126,N_6451);
nor U7817 (N_7817,N_7353,N_6574);
nand U7818 (N_7818,N_5347,N_6692);
or U7819 (N_7819,N_5980,N_5263);
nor U7820 (N_7820,N_6245,N_6413);
nand U7821 (N_7821,N_5917,N_6552);
nor U7822 (N_7822,N_5433,N_6416);
or U7823 (N_7823,N_5542,N_7331);
and U7824 (N_7824,N_7006,N_7251);
and U7825 (N_7825,N_5886,N_7312);
and U7826 (N_7826,N_5713,N_5567);
nand U7827 (N_7827,N_5057,N_6403);
and U7828 (N_7828,N_5437,N_6479);
nor U7829 (N_7829,N_5238,N_6010);
nand U7830 (N_7830,N_6251,N_7141);
nor U7831 (N_7831,N_5452,N_6810);
nor U7832 (N_7832,N_5657,N_5340);
nand U7833 (N_7833,N_7160,N_6519);
nor U7834 (N_7834,N_5196,N_6128);
nand U7835 (N_7835,N_5308,N_7373);
nor U7836 (N_7836,N_5149,N_5847);
nor U7837 (N_7837,N_5466,N_5752);
or U7838 (N_7838,N_5724,N_6332);
and U7839 (N_7839,N_6193,N_6386);
nor U7840 (N_7840,N_6235,N_6223);
nand U7841 (N_7841,N_6523,N_6760);
nand U7842 (N_7842,N_7486,N_6109);
nor U7843 (N_7843,N_7177,N_5570);
nor U7844 (N_7844,N_7293,N_5949);
nand U7845 (N_7845,N_7189,N_6932);
and U7846 (N_7846,N_7091,N_7196);
nor U7847 (N_7847,N_6214,N_5075);
xor U7848 (N_7848,N_5435,N_7398);
and U7849 (N_7849,N_5895,N_5103);
nor U7850 (N_7850,N_5226,N_6353);
xor U7851 (N_7851,N_7239,N_7188);
or U7852 (N_7852,N_7199,N_7165);
nand U7853 (N_7853,N_6839,N_5564);
nand U7854 (N_7854,N_5292,N_5838);
and U7855 (N_7855,N_5553,N_7461);
and U7856 (N_7856,N_6555,N_6289);
nor U7857 (N_7857,N_5502,N_5843);
nand U7858 (N_7858,N_5636,N_6067);
nand U7859 (N_7859,N_5266,N_5731);
xor U7860 (N_7860,N_7232,N_5766);
and U7861 (N_7861,N_5803,N_5569);
and U7862 (N_7862,N_6658,N_7001);
nand U7863 (N_7863,N_5320,N_6461);
nor U7864 (N_7864,N_5759,N_6797);
nand U7865 (N_7865,N_5580,N_5776);
nand U7866 (N_7866,N_7324,N_5737);
and U7867 (N_7867,N_5780,N_6506);
and U7868 (N_7868,N_6892,N_5664);
and U7869 (N_7869,N_6836,N_6457);
nor U7870 (N_7870,N_7011,N_5253);
and U7871 (N_7871,N_5728,N_6595);
nand U7872 (N_7872,N_7340,N_5573);
nor U7873 (N_7873,N_5533,N_7146);
or U7874 (N_7874,N_6950,N_7077);
and U7875 (N_7875,N_5970,N_5607);
nand U7876 (N_7876,N_6622,N_7315);
nand U7877 (N_7877,N_5609,N_7416);
nor U7878 (N_7878,N_5082,N_6034);
nor U7879 (N_7879,N_5379,N_6415);
or U7880 (N_7880,N_7497,N_6153);
nand U7881 (N_7881,N_7305,N_5957);
nor U7882 (N_7882,N_6283,N_7336);
or U7883 (N_7883,N_6991,N_5666);
nor U7884 (N_7884,N_7100,N_6553);
or U7885 (N_7885,N_6354,N_6196);
nand U7886 (N_7886,N_7228,N_6866);
nand U7887 (N_7887,N_6709,N_5708);
or U7888 (N_7888,N_5969,N_5463);
nor U7889 (N_7889,N_5572,N_5244);
nor U7890 (N_7890,N_5595,N_6704);
or U7891 (N_7891,N_7367,N_5758);
and U7892 (N_7892,N_7213,N_6111);
nand U7893 (N_7893,N_5114,N_6585);
nor U7894 (N_7894,N_6616,N_6957);
and U7895 (N_7895,N_6362,N_5627);
nand U7896 (N_7896,N_6864,N_6478);
nor U7897 (N_7897,N_7211,N_6988);
nor U7898 (N_7898,N_5994,N_5325);
nand U7899 (N_7899,N_5348,N_6320);
and U7900 (N_7900,N_5924,N_5065);
xor U7901 (N_7901,N_6820,N_6800);
xor U7902 (N_7902,N_5105,N_7110);
nor U7903 (N_7903,N_5861,N_7276);
or U7904 (N_7904,N_7363,N_7412);
nor U7905 (N_7905,N_5389,N_7466);
nor U7906 (N_7906,N_7116,N_5319);
xor U7907 (N_7907,N_6691,N_5033);
or U7908 (N_7908,N_5372,N_6683);
or U7909 (N_7909,N_6277,N_7279);
and U7910 (N_7910,N_6984,N_5714);
nor U7911 (N_7911,N_6234,N_6306);
or U7912 (N_7912,N_6943,N_6056);
nor U7913 (N_7913,N_5884,N_7257);
and U7914 (N_7914,N_5640,N_5021);
or U7915 (N_7915,N_7457,N_6250);
nand U7916 (N_7916,N_5100,N_6236);
nand U7917 (N_7917,N_6390,N_6786);
or U7918 (N_7918,N_6465,N_6661);
nand U7919 (N_7919,N_6059,N_6824);
or U7920 (N_7920,N_6038,N_6647);
nor U7921 (N_7921,N_6404,N_6565);
nor U7922 (N_7922,N_5605,N_6773);
nor U7923 (N_7923,N_5271,N_5582);
nor U7924 (N_7924,N_6542,N_6001);
nor U7925 (N_7925,N_7082,N_7447);
and U7926 (N_7926,N_6294,N_7064);
and U7927 (N_7927,N_6247,N_5068);
or U7928 (N_7928,N_5529,N_5588);
and U7929 (N_7929,N_7167,N_6693);
and U7930 (N_7930,N_5375,N_6532);
and U7931 (N_7931,N_5007,N_7045);
and U7932 (N_7932,N_6732,N_6288);
and U7933 (N_7933,N_6543,N_5885);
nor U7934 (N_7934,N_5044,N_6515);
nand U7935 (N_7935,N_6072,N_6099);
or U7936 (N_7936,N_6007,N_6222);
nand U7937 (N_7937,N_6476,N_5450);
nor U7938 (N_7938,N_6987,N_7114);
nor U7939 (N_7939,N_5398,N_7149);
nor U7940 (N_7940,N_5413,N_6016);
and U7941 (N_7941,N_7265,N_7021);
and U7942 (N_7942,N_6036,N_6272);
nor U7943 (N_7943,N_6454,N_5141);
and U7944 (N_7944,N_6583,N_6189);
nor U7945 (N_7945,N_5883,N_6028);
nor U7946 (N_7946,N_6173,N_6285);
or U7947 (N_7947,N_7480,N_6959);
and U7948 (N_7948,N_6359,N_6733);
xnor U7949 (N_7949,N_6664,N_7068);
and U7950 (N_7950,N_6350,N_6075);
nand U7951 (N_7951,N_5959,N_5210);
and U7952 (N_7952,N_6460,N_6340);
or U7953 (N_7953,N_5882,N_6005);
nand U7954 (N_7954,N_7347,N_5156);
or U7955 (N_7955,N_5247,N_5002);
nor U7956 (N_7956,N_5517,N_5853);
nand U7957 (N_7957,N_5775,N_5423);
and U7958 (N_7958,N_6623,N_7104);
or U7959 (N_7959,N_5680,N_6395);
xnor U7960 (N_7960,N_5826,N_6835);
nor U7961 (N_7961,N_6425,N_6570);
nand U7962 (N_7962,N_6452,N_6310);
and U7963 (N_7963,N_6526,N_6904);
nand U7964 (N_7964,N_5592,N_7405);
xnor U7965 (N_7965,N_5685,N_5303);
nand U7966 (N_7966,N_5040,N_5457);
or U7967 (N_7967,N_6097,N_6867);
nand U7968 (N_7968,N_5559,N_6755);
nand U7969 (N_7969,N_5147,N_5996);
nand U7970 (N_7970,N_5711,N_5377);
and U7971 (N_7971,N_6155,N_7139);
nor U7972 (N_7972,N_6968,N_7237);
and U7973 (N_7973,N_6492,N_7095);
nand U7974 (N_7974,N_5662,N_6414);
and U7975 (N_7975,N_5276,N_5027);
and U7976 (N_7976,N_5221,N_6854);
and U7977 (N_7977,N_7215,N_6556);
nand U7978 (N_7978,N_6047,N_5783);
and U7979 (N_7979,N_5626,N_5793);
or U7980 (N_7980,N_5535,N_5317);
nor U7981 (N_7981,N_7150,N_6436);
or U7982 (N_7982,N_7092,N_7197);
nor U7983 (N_7983,N_6637,N_6426);
nand U7984 (N_7984,N_6912,N_6131);
nor U7985 (N_7985,N_7337,N_6640);
and U7986 (N_7986,N_7484,N_7062);
or U7987 (N_7987,N_7216,N_7442);
nor U7988 (N_7988,N_6629,N_6751);
nor U7989 (N_7989,N_5171,N_6440);
nand U7990 (N_7990,N_5874,N_6924);
or U7991 (N_7991,N_6848,N_7302);
or U7992 (N_7992,N_7157,N_5367);
nor U7993 (N_7993,N_5427,N_5811);
nor U7994 (N_7994,N_6823,N_7298);
xnor U7995 (N_7995,N_6628,N_5777);
nor U7996 (N_7996,N_7332,N_6955);
and U7997 (N_7997,N_6256,N_6322);
nand U7998 (N_7998,N_6859,N_7424);
and U7999 (N_7999,N_6895,N_5229);
and U8000 (N_8000,N_6757,N_7493);
nor U8001 (N_8001,N_6923,N_7007);
or U8002 (N_8002,N_7494,N_6078);
or U8003 (N_8003,N_5094,N_6560);
and U8004 (N_8004,N_6458,N_6512);
nor U8005 (N_8005,N_5707,N_6550);
nor U8006 (N_8006,N_6042,N_6018);
xnor U8007 (N_8007,N_6772,N_6163);
nand U8008 (N_8008,N_5307,N_6233);
or U8009 (N_8009,N_5354,N_5436);
nand U8010 (N_8010,N_5151,N_7474);
and U8011 (N_8011,N_6917,N_5788);
or U8012 (N_8012,N_5726,N_6143);
and U8013 (N_8013,N_5272,N_5204);
nand U8014 (N_8014,N_6840,N_6916);
nor U8015 (N_8015,N_5197,N_7131);
xnor U8016 (N_8016,N_5326,N_7359);
and U8017 (N_8017,N_6342,N_6607);
and U8018 (N_8018,N_7097,N_6869);
nor U8019 (N_8019,N_6731,N_6201);
and U8020 (N_8020,N_7201,N_6317);
nor U8021 (N_8021,N_6295,N_6516);
nor U8022 (N_8022,N_7036,N_7402);
and U8023 (N_8023,N_6224,N_6330);
nor U8024 (N_8024,N_6901,N_6740);
and U8025 (N_8025,N_5988,N_5363);
and U8026 (N_8026,N_6736,N_7218);
or U8027 (N_8027,N_6765,N_5063);
nor U8028 (N_8028,N_5632,N_6842);
and U8029 (N_8029,N_5800,N_5145);
nor U8030 (N_8030,N_6702,N_6971);
nand U8031 (N_8031,N_6229,N_6761);
and U8032 (N_8032,N_5862,N_5872);
xnor U8033 (N_8033,N_6407,N_7304);
and U8034 (N_8034,N_5344,N_5700);
nor U8035 (N_8035,N_7185,N_7255);
xnor U8036 (N_8036,N_6361,N_5686);
or U8037 (N_8037,N_7147,N_5504);
or U8038 (N_8038,N_5321,N_5785);
or U8039 (N_8039,N_6645,N_6194);
and U8040 (N_8040,N_6929,N_5878);
nand U8041 (N_8041,N_5462,N_6021);
nor U8042 (N_8042,N_6278,N_6958);
nand U8043 (N_8043,N_6280,N_6966);
and U8044 (N_8044,N_6688,N_6915);
nor U8045 (N_8045,N_6168,N_6107);
nor U8046 (N_8046,N_7375,N_5402);
nor U8047 (N_8047,N_7410,N_7101);
nand U8048 (N_8048,N_5235,N_5390);
nor U8049 (N_8049,N_6582,N_5162);
nor U8050 (N_8050,N_5760,N_5181);
or U8051 (N_8051,N_5179,N_7296);
xor U8052 (N_8052,N_5295,N_6706);
nor U8053 (N_8053,N_6608,N_5445);
nand U8054 (N_8054,N_6853,N_6409);
nand U8055 (N_8055,N_5217,N_5715);
xnor U8056 (N_8056,N_6496,N_7470);
nor U8057 (N_8057,N_6529,N_5912);
nor U8058 (N_8058,N_6674,N_7459);
nand U8059 (N_8059,N_6026,N_6885);
nor U8060 (N_8060,N_6393,N_6313);
and U8061 (N_8061,N_7226,N_7449);
nand U8062 (N_8062,N_7425,N_7487);
or U8063 (N_8063,N_7222,N_6259);
and U8064 (N_8064,N_6779,N_6941);
and U8065 (N_8065,N_5620,N_6266);
nand U8066 (N_8066,N_5284,N_5965);
nor U8067 (N_8067,N_6894,N_6120);
and U8068 (N_8068,N_5910,N_6850);
nor U8069 (N_8069,N_5528,N_6564);
nand U8070 (N_8070,N_5144,N_6724);
or U8071 (N_8071,N_6626,N_5260);
or U8072 (N_8072,N_6684,N_5189);
and U8073 (N_8073,N_6568,N_5501);
nor U8074 (N_8074,N_5131,N_6713);
nor U8075 (N_8075,N_7207,N_6352);
nor U8076 (N_8076,N_7023,N_6592);
and U8077 (N_8077,N_5386,N_5740);
nand U8078 (N_8078,N_5449,N_5146);
or U8079 (N_8079,N_6817,N_7187);
and U8080 (N_8080,N_5812,N_5474);
nor U8081 (N_8081,N_6981,N_5359);
xnor U8082 (N_8082,N_6011,N_7035);
or U8083 (N_8083,N_5017,N_6752);
nor U8084 (N_8084,N_5055,N_5555);
and U8085 (N_8085,N_7397,N_6613);
nor U8086 (N_8086,N_6624,N_5168);
nand U8087 (N_8087,N_7117,N_7469);
or U8088 (N_8088,N_6347,N_7032);
nand U8089 (N_8089,N_7127,N_7087);
or U8090 (N_8090,N_5534,N_6207);
or U8091 (N_8091,N_5069,N_7126);
and U8092 (N_8092,N_5526,N_7441);
and U8093 (N_8093,N_5023,N_6369);
nand U8094 (N_8094,N_6012,N_6127);
nand U8095 (N_8095,N_5026,N_6986);
nor U8096 (N_8096,N_6282,N_6832);
or U8097 (N_8097,N_5493,N_6376);
or U8098 (N_8098,N_5815,N_5798);
nand U8099 (N_8099,N_5561,N_6738);
or U8100 (N_8100,N_5108,N_5840);
nor U8101 (N_8101,N_5310,N_7260);
or U8102 (N_8102,N_5381,N_7055);
nor U8103 (N_8103,N_5475,N_5923);
or U8104 (N_8104,N_5118,N_6252);
and U8105 (N_8105,N_6716,N_6572);
nand U8106 (N_8106,N_5819,N_7033);
xnor U8107 (N_8107,N_5461,N_6671);
and U8108 (N_8108,N_5468,N_5314);
and U8109 (N_8109,N_6826,N_6383);
xnor U8110 (N_8110,N_7134,N_7477);
and U8111 (N_8111,N_7138,N_7047);
or U8112 (N_8112,N_6031,N_5786);
nand U8113 (N_8113,N_6780,N_5820);
nor U8114 (N_8114,N_6632,N_6635);
and U8115 (N_8115,N_6802,N_7120);
nand U8116 (N_8116,N_6520,N_6314);
nand U8117 (N_8117,N_5066,N_7050);
nor U8118 (N_8118,N_5249,N_5251);
and U8119 (N_8119,N_5277,N_5411);
nand U8120 (N_8120,N_6967,N_6960);
nor U8121 (N_8121,N_6228,N_6545);
or U8122 (N_8122,N_7094,N_6822);
nand U8123 (N_8123,N_7245,N_5508);
or U8124 (N_8124,N_5207,N_5587);
nand U8125 (N_8125,N_6505,N_6672);
or U8126 (N_8126,N_5270,N_6299);
or U8127 (N_8127,N_7417,N_5085);
nor U8128 (N_8128,N_6927,N_6680);
nand U8129 (N_8129,N_5334,N_6539);
nor U8130 (N_8130,N_6064,N_5153);
nor U8131 (N_8131,N_7334,N_5224);
or U8132 (N_8132,N_7022,N_5795);
or U8133 (N_8133,N_7323,N_5180);
nor U8134 (N_8134,N_6710,N_6382);
and U8135 (N_8135,N_6908,N_5404);
and U8136 (N_8136,N_6942,N_6114);
nand U8137 (N_8137,N_5290,N_6548);
nand U8138 (N_8138,N_5015,N_7172);
nor U8139 (N_8139,N_6096,N_5071);
nand U8140 (N_8140,N_5116,N_5268);
nor U8141 (N_8141,N_5673,N_7209);
nand U8142 (N_8142,N_5639,N_5024);
nor U8143 (N_8143,N_5984,N_5692);
nand U8144 (N_8144,N_6796,N_7361);
nor U8145 (N_8145,N_5712,N_6387);
and U8146 (N_8146,N_5084,N_5351);
nand U8147 (N_8147,N_6154,N_6237);
nor U8148 (N_8148,N_7446,N_7109);
nor U8149 (N_8149,N_5833,N_7000);
nor U8150 (N_8150,N_5169,N_5754);
nand U8151 (N_8151,N_6778,N_6949);
and U8152 (N_8152,N_7174,N_6105);
nand U8153 (N_8153,N_5378,N_7238);
and U8154 (N_8154,N_5589,N_5301);
nor U8155 (N_8155,N_5269,N_5259);
nand U8156 (N_8156,N_6074,N_6580);
or U8157 (N_8157,N_7297,N_5671);
nor U8158 (N_8158,N_5152,N_6311);
and U8159 (N_8159,N_6567,N_6513);
nand U8160 (N_8160,N_6076,N_6142);
and U8161 (N_8161,N_5522,N_5556);
nor U8162 (N_8162,N_6775,N_6985);
or U8163 (N_8163,N_6546,N_5612);
nand U8164 (N_8164,N_6472,N_6500);
nor U8165 (N_8165,N_6069,N_5241);
nand U8166 (N_8166,N_6110,N_7319);
or U8167 (N_8167,N_6357,N_7409);
or U8168 (N_8168,N_5428,N_5600);
nand U8169 (N_8169,N_5250,N_6271);
and U8170 (N_8170,N_6547,N_6281);
nor U8171 (N_8171,N_5164,N_5213);
nor U8172 (N_8172,N_6179,N_5998);
nor U8173 (N_8173,N_5975,N_5892);
or U8174 (N_8174,N_6084,N_5515);
nor U8175 (N_8175,N_5850,N_5581);
or U8176 (N_8176,N_5081,N_6584);
and U8177 (N_8177,N_5653,N_6871);
or U8178 (N_8178,N_5391,N_6345);
nor U8179 (N_8179,N_7433,N_5660);
nand U8180 (N_8180,N_7010,N_7434);
nor U8181 (N_8181,N_5593,N_7436);
nand U8182 (N_8182,N_6152,N_6399);
nor U8183 (N_8183,N_7342,N_6695);
and U8184 (N_8184,N_6612,N_6868);
or U8185 (N_8185,N_6183,N_6788);
or U8186 (N_8186,N_6599,N_5841);
and U8187 (N_8187,N_6963,N_7084);
and U8188 (N_8188,N_5637,N_7124);
and U8189 (N_8189,N_5165,N_5405);
nor U8190 (N_8190,N_5645,N_5200);
or U8191 (N_8191,N_6490,N_6435);
nand U8192 (N_8192,N_5614,N_5117);
and U8193 (N_8193,N_6711,N_5866);
nor U8194 (N_8194,N_5842,N_6394);
or U8195 (N_8195,N_5240,N_5274);
and U8196 (N_8196,N_6670,N_5393);
or U8197 (N_8197,N_6205,N_7269);
nand U8198 (N_8198,N_7212,N_5721);
or U8199 (N_8199,N_6631,N_6723);
nand U8200 (N_8200,N_6873,N_5813);
xnor U8201 (N_8201,N_5483,N_6925);
nand U8202 (N_8202,N_5454,N_7448);
or U8203 (N_8203,N_6718,N_6857);
nor U8204 (N_8204,N_5432,N_7242);
or U8205 (N_8205,N_7037,N_7419);
nor U8206 (N_8206,N_6947,N_7028);
nor U8207 (N_8207,N_6681,N_7170);
nor U8208 (N_8208,N_5825,N_5062);
or U8209 (N_8209,N_6368,N_6938);
nand U8210 (N_8210,N_6325,N_5136);
or U8211 (N_8211,N_6509,N_7133);
nor U8212 (N_8212,N_7380,N_7029);
or U8213 (N_8213,N_5212,N_6135);
nor U8214 (N_8214,N_5584,N_7383);
nand U8215 (N_8215,N_5192,N_6053);
or U8216 (N_8216,N_6343,N_6083);
nand U8217 (N_8217,N_7183,N_6818);
or U8218 (N_8218,N_6437,N_5089);
nand U8219 (N_8219,N_7430,N_6132);
nor U8220 (N_8220,N_6326,N_5232);
or U8221 (N_8221,N_6905,N_6855);
or U8222 (N_8222,N_7294,N_5365);
nor U8223 (N_8223,N_5676,N_5688);
and U8224 (N_8224,N_6535,N_6090);
nor U8225 (N_8225,N_5763,N_7437);
and U8226 (N_8226,N_6400,N_5696);
nor U8227 (N_8227,N_6464,N_7220);
and U8228 (N_8228,N_6315,N_6115);
or U8229 (N_8229,N_5560,N_6926);
or U8230 (N_8230,N_6875,N_5339);
and U8231 (N_8231,N_6918,N_6829);
nor U8232 (N_8232,N_7089,N_6502);
or U8233 (N_8233,N_5353,N_7435);
nor U8234 (N_8234,N_5211,N_5979);
nand U8235 (N_8235,N_6551,N_6990);
nor U8236 (N_8236,N_6508,N_7460);
nor U8237 (N_8237,N_6032,N_7341);
nor U8238 (N_8238,N_6816,N_5119);
nand U8239 (N_8239,N_5675,N_5476);
nor U8240 (N_8240,N_6333,N_5682);
and U8241 (N_8241,N_7108,N_5003);
and U8242 (N_8242,N_5665,N_5086);
nor U8243 (N_8243,N_5004,N_7227);
nor U8244 (N_8244,N_5739,N_6388);
and U8245 (N_8245,N_7348,N_6896);
nor U8246 (N_8246,N_6378,N_7169);
nand U8247 (N_8247,N_5689,N_5336);
nand U8248 (N_8248,N_5399,N_5137);
or U8249 (N_8249,N_5485,N_7217);
and U8250 (N_8250,N_5967,N_5465);
nor U8251 (N_8251,N_6052,N_6982);
or U8252 (N_8252,N_5173,N_5337);
or U8253 (N_8253,N_5936,N_6125);
nand U8254 (N_8254,N_5925,N_6448);
and U8255 (N_8255,N_7070,N_6538);
or U8256 (N_8256,N_5681,N_6939);
nand U8257 (N_8257,N_6148,N_6676);
or U8258 (N_8258,N_5932,N_7283);
nor U8259 (N_8259,N_7012,N_5663);
and U8260 (N_8260,N_7080,N_5649);
and U8261 (N_8261,N_6238,N_6442);
or U8262 (N_8262,N_7378,N_7478);
nand U8263 (N_8263,N_6804,N_6737);
nand U8264 (N_8264,N_6244,N_6215);
or U8265 (N_8265,N_6969,N_6521);
nor U8266 (N_8266,N_7040,N_6384);
nor U8267 (N_8267,N_6418,N_5345);
nor U8268 (N_8268,N_5447,N_6909);
nand U8269 (N_8269,N_6762,N_6837);
nor U8270 (N_8270,N_5409,N_5470);
and U8271 (N_8271,N_5376,N_6117);
and U8272 (N_8272,N_6318,N_5635);
or U8273 (N_8273,N_5201,N_6844);
xor U8274 (N_8274,N_5568,N_6027);
and U8275 (N_8275,N_6594,N_6212);
or U8276 (N_8276,N_7491,N_6605);
nand U8277 (N_8277,N_6121,N_5926);
nand U8278 (N_8278,N_6708,N_5768);
nand U8279 (N_8279,N_5974,N_7229);
and U8280 (N_8280,N_6933,N_5810);
and U8281 (N_8281,N_6591,N_5880);
nand U8282 (N_8282,N_5058,N_5821);
or U8283 (N_8283,N_6994,N_6287);
nand U8284 (N_8284,N_7074,N_7194);
nor U8285 (N_8285,N_5944,N_6596);
nor U8286 (N_8286,N_5406,N_5167);
and U8287 (N_8287,N_5875,N_5361);
or U8288 (N_8288,N_6218,N_5860);
and U8289 (N_8289,N_6998,N_5797);
nand U8290 (N_8290,N_5387,N_7241);
nor U8291 (N_8291,N_5032,N_5155);
and U8292 (N_8292,N_7119,N_5594);
nand U8293 (N_8293,N_6874,N_7404);
nand U8294 (N_8294,N_5623,N_7288);
or U8295 (N_8295,N_5028,N_6243);
nand U8296 (N_8296,N_5530,N_7085);
nand U8297 (N_8297,N_7355,N_5104);
nand U8298 (N_8298,N_5010,N_5591);
or U8299 (N_8299,N_5647,N_6328);
nand U8300 (N_8300,N_7377,N_5059);
and U8301 (N_8301,N_7034,N_5288);
nand U8302 (N_8302,N_6022,N_5687);
and U8303 (N_8303,N_6220,N_5509);
nand U8304 (N_8304,N_5918,N_6240);
and U8305 (N_8305,N_6602,N_6092);
nor U8306 (N_8306,N_7498,N_6473);
or U8307 (N_8307,N_5610,N_7407);
and U8308 (N_8308,N_7335,N_5540);
and U8309 (N_8309,N_6113,N_5510);
and U8310 (N_8310,N_6893,N_6401);
or U8311 (N_8311,N_7482,N_7002);
or U8312 (N_8312,N_5602,N_6006);
or U8313 (N_8313,N_7086,N_6687);
nand U8314 (N_8314,N_5172,N_6497);
nand U8315 (N_8315,N_5937,N_7351);
nand U8316 (N_8316,N_6494,N_5464);
nand U8317 (N_8317,N_7262,N_7137);
or U8318 (N_8318,N_5966,N_5669);
or U8319 (N_8319,N_7420,N_5106);
nor U8320 (N_8320,N_7352,N_6589);
nand U8321 (N_8321,N_6787,N_6753);
nand U8322 (N_8322,N_6717,N_5578);
xor U8323 (N_8323,N_5380,N_6372);
or U8324 (N_8324,N_5732,N_5037);
nand U8325 (N_8325,N_6790,N_5543);
nand U8326 (N_8326,N_5287,N_5765);
nand U8327 (N_8327,N_6954,N_5744);
nand U8328 (N_8328,N_7370,N_5651);
xor U8329 (N_8329,N_7121,N_7476);
nor U8330 (N_8330,N_5020,N_7307);
nor U8331 (N_8331,N_7155,N_6902);
nand U8332 (N_8332,N_5646,N_6530);
nand U8333 (N_8333,N_5364,N_5479);
xor U8334 (N_8334,N_7465,N_6649);
nand U8335 (N_8335,N_5771,N_6208);
or U8336 (N_8336,N_6791,N_7200);
nand U8337 (N_8337,N_6712,N_5444);
nand U8338 (N_8338,N_6351,N_7135);
or U8339 (N_8339,N_7365,N_6549);
and U8340 (N_8340,N_6305,N_5539);
nand U8341 (N_8341,N_5514,N_7358);
nand U8342 (N_8342,N_6123,N_6441);
and U8343 (N_8343,N_5824,N_6086);
xnor U8344 (N_8344,N_5611,N_7422);
and U8345 (N_8345,N_5851,N_5677);
nand U8346 (N_8346,N_5963,N_5905);
or U8347 (N_8347,N_5844,N_7015);
xnor U8348 (N_8348,N_5041,N_5022);
or U8349 (N_8349,N_6819,N_7072);
nand U8350 (N_8350,N_6033,N_6434);
nand U8351 (N_8351,N_6544,N_5013);
nor U8352 (N_8352,N_7129,N_6654);
nor U8353 (N_8353,N_5678,N_5487);
and U8354 (N_8354,N_7205,N_6993);
or U8355 (N_8355,N_5505,N_7041);
or U8356 (N_8356,N_6176,N_6665);
and U8357 (N_8357,N_6487,N_7309);
nand U8358 (N_8358,N_6398,N_5127);
or U8359 (N_8359,N_5989,N_5185);
xor U8360 (N_8360,N_6953,N_7246);
and U8361 (N_8361,N_5335,N_6559);
and U8362 (N_8362,N_5849,N_7078);
nand U8363 (N_8363,N_5719,N_6338);
nand U8364 (N_8364,N_5009,N_7214);
nor U8365 (N_8365,N_6781,N_6830);
nand U8366 (N_8366,N_5857,N_5356);
nor U8367 (N_8367,N_5215,N_6974);
and U8368 (N_8368,N_5667,N_7357);
and U8369 (N_8369,N_5773,N_7198);
nor U8370 (N_8370,N_7099,N_7038);
nor U8371 (N_8371,N_7003,N_6700);
or U8372 (N_8372,N_5630,N_5309);
and U8373 (N_8373,N_5735,N_6563);
and U8374 (N_8374,N_5981,N_7061);
nand U8375 (N_8375,N_5518,N_6514);
nor U8376 (N_8376,N_5641,N_7096);
nand U8377 (N_8377,N_5160,N_7009);
and U8378 (N_8378,N_5093,N_5807);
and U8379 (N_8379,N_5001,N_6983);
and U8380 (N_8380,N_7362,N_5322);
nor U8381 (N_8381,N_5683,N_6759);
or U8382 (N_8382,N_5074,N_6257);
nor U8383 (N_8383,N_6852,N_6621);
and U8384 (N_8384,N_6697,N_7360);
and U8385 (N_8385,N_7322,N_6166);
xor U8386 (N_8386,N_7300,N_6419);
nor U8387 (N_8387,N_6020,N_5985);
or U8388 (N_8388,N_6805,N_7113);
nand U8389 (N_8389,N_5519,N_7455);
or U8390 (N_8390,N_5198,N_5177);
nor U8391 (N_8391,N_7292,N_5566);
nor U8392 (N_8392,N_5928,N_6141);
and U8393 (N_8393,N_5723,N_7054);
or U8394 (N_8394,N_5867,N_5946);
nor U8395 (N_8395,N_5060,N_6108);
or U8396 (N_8396,N_5618,N_7290);
or U8397 (N_8397,N_5896,N_7317);
xor U8398 (N_8398,N_5927,N_7076);
and U8399 (N_8399,N_5125,N_6694);
or U8400 (N_8400,N_6656,N_7225);
and U8401 (N_8401,N_5919,N_6348);
or U8402 (N_8402,N_5904,N_5008);
and U8403 (N_8403,N_5695,N_6186);
and U8404 (N_8404,N_6846,N_7418);
and U8405 (N_8405,N_6914,N_7027);
nand U8406 (N_8406,N_6828,N_6653);
nor U8407 (N_8407,N_6462,N_6561);
nor U8408 (N_8408,N_6618,N_6501);
or U8409 (N_8409,N_5648,N_5787);
or U8410 (N_8410,N_5256,N_6184);
nor U8411 (N_8411,N_6444,N_5362);
or U8412 (N_8412,N_6045,N_6355);
or U8413 (N_8413,N_5342,N_5701);
nor U8414 (N_8414,N_7244,N_7330);
and U8415 (N_8415,N_5906,N_6619);
nor U8416 (N_8416,N_6668,N_5111);
nand U8417 (N_8417,N_6077,N_6715);
or U8418 (N_8418,N_5338,N_5374);
nand U8419 (N_8419,N_7384,N_7438);
nand U8420 (N_8420,N_6528,N_6187);
xor U8421 (N_8421,N_5477,N_5415);
or U8422 (N_8422,N_6375,N_6292);
nand U8423 (N_8423,N_6972,N_5500);
or U8424 (N_8424,N_7391,N_7125);
nand U8425 (N_8425,N_5178,N_5414);
nor U8426 (N_8426,N_7098,N_6769);
or U8427 (N_8427,N_7048,N_5684);
or U8428 (N_8428,N_5305,N_5633);
and U8429 (N_8429,N_6474,N_5706);
or U8430 (N_8430,N_5691,N_5031);
nand U8431 (N_8431,N_6087,N_6849);
and U8432 (N_8432,N_5018,N_7318);
or U8433 (N_8433,N_6405,N_6261);
and U8434 (N_8434,N_5527,N_6876);
or U8435 (N_8435,N_5067,N_5132);
and U8436 (N_8436,N_6172,N_7176);
or U8437 (N_8437,N_5908,N_5956);
nand U8438 (N_8438,N_7473,N_7179);
and U8439 (N_8439,N_7118,N_7453);
nor U8440 (N_8440,N_5267,N_6192);
nor U8441 (N_8441,N_5954,N_6094);
nor U8442 (N_8442,N_6040,N_6743);
or U8443 (N_8443,N_6210,N_5805);
nor U8444 (N_8444,N_6898,N_5355);
and U8445 (N_8445,N_5491,N_6511);
nand U8446 (N_8446,N_5407,N_6630);
xor U8447 (N_8447,N_6199,N_6015);
and U8448 (N_8448,N_5299,N_5330);
or U8449 (N_8449,N_5922,N_5030);
nor U8450 (N_8450,N_6296,N_7451);
nand U8451 (N_8451,N_5679,N_7366);
nor U8452 (N_8452,N_6907,N_5046);
nor U8453 (N_8453,N_6262,N_6273);
and U8454 (N_8454,N_5148,N_6995);
or U8455 (N_8455,N_5889,N_6447);
or U8456 (N_8456,N_7495,N_7485);
xor U8457 (N_8457,N_5748,N_6643);
nand U8458 (N_8458,N_5421,N_7115);
nand U8459 (N_8459,N_7203,N_6940);
or U8460 (N_8460,N_6198,N_7443);
and U8461 (N_8461,N_5729,N_5076);
or U8462 (N_8462,N_5442,N_5460);
nand U8463 (N_8463,N_6662,N_7151);
xor U8464 (N_8464,N_6756,N_5576);
nand U8465 (N_8465,N_6088,N_5583);
nand U8466 (N_8466,N_5536,N_6467);
nor U8467 (N_8467,N_7263,N_5562);
or U8468 (N_8468,N_5237,N_6346);
and U8469 (N_8469,N_5604,N_5343);
nand U8470 (N_8470,N_6639,N_7345);
nand U8471 (N_8471,N_7004,N_6794);
nor U8472 (N_8472,N_6297,N_7310);
and U8473 (N_8473,N_5182,N_6482);
and U8474 (N_8474,N_7173,N_5654);
nand U8475 (N_8475,N_6573,N_7206);
nand U8476 (N_8476,N_5804,N_6133);
nor U8477 (N_8477,N_6707,N_7395);
nor U8478 (N_8478,N_7059,N_6396);
and U8479 (N_8479,N_7462,N_6677);
and U8480 (N_8480,N_6518,N_7371);
nor U8481 (N_8481,N_6060,N_6331);
or U8482 (N_8482,N_5756,N_7231);
nor U8483 (N_8483,N_7158,N_6432);
and U8484 (N_8484,N_6831,N_6253);
or U8485 (N_8485,N_6420,N_6085);
or U8486 (N_8486,N_5993,N_5332);
nor U8487 (N_8487,N_5997,N_5784);
nand U8488 (N_8488,N_6650,N_6748);
and U8489 (N_8489,N_5772,N_5166);
nor U8490 (N_8490,N_6358,N_6004);
and U8491 (N_8491,N_6646,N_5690);
and U8492 (N_8492,N_5879,N_7057);
nor U8493 (N_8493,N_6862,N_6221);
or U8494 (N_8494,N_5774,N_5230);
nor U8495 (N_8495,N_7252,N_5547);
nor U8496 (N_8496,N_5191,N_7306);
nand U8497 (N_8497,N_5931,N_5064);
and U8498 (N_8498,N_6495,N_5903);
nor U8499 (N_8499,N_5537,N_6537);
and U8500 (N_8500,N_6527,N_5548);
nand U8501 (N_8501,N_6174,N_5101);
and U8502 (N_8502,N_5634,N_5710);
and U8503 (N_8503,N_5631,N_5183);
or U8504 (N_8504,N_5796,N_6116);
and U8505 (N_8505,N_6379,N_6679);
nor U8506 (N_8506,N_6834,N_6134);
nand U8507 (N_8507,N_6809,N_5953);
nand U8508 (N_8508,N_6682,N_7204);
nor U8509 (N_8509,N_5408,N_5608);
and U8510 (N_8510,N_7171,N_7280);
nand U8511 (N_8511,N_5720,N_6517);
nor U8512 (N_8512,N_5315,N_5053);
or U8513 (N_8513,N_6043,N_5516);
and U8514 (N_8514,N_6231,N_6209);
or U8515 (N_8515,N_5206,N_5459);
and U8516 (N_8516,N_7153,N_6827);
nand U8517 (N_8517,N_6255,N_6641);
and U8518 (N_8518,N_5941,N_7471);
nand U8519 (N_8519,N_7044,N_6445);
or U8520 (N_8520,N_5257,N_7090);
or U8521 (N_8521,N_5418,N_5499);
and U8522 (N_8522,N_5199,N_5693);
and U8523 (N_8523,N_5494,N_7314);
nor U8524 (N_8524,N_7479,N_5597);
or U8525 (N_8525,N_5816,N_7210);
and U8526 (N_8526,N_5126,N_5175);
or U8527 (N_8527,N_6764,N_5831);
nand U8528 (N_8528,N_6050,N_5852);
and U8529 (N_8529,N_5050,N_5498);
nand U8530 (N_8530,N_6181,N_5488);
or U8531 (N_8531,N_5590,N_5282);
nand U8532 (N_8532,N_6098,N_6080);
or U8533 (N_8533,N_5401,N_7281);
nand U8534 (N_8534,N_5577,N_6617);
nand U8535 (N_8535,N_6522,N_6610);
or U8536 (N_8536,N_6203,N_6302);
nor U8537 (N_8537,N_5948,N_5331);
nor U8538 (N_8538,N_6906,N_6260);
or U8539 (N_8539,N_5056,N_5839);
and U8540 (N_8540,N_6427,N_5809);
and U8541 (N_8541,N_5135,N_5563);
and U8542 (N_8542,N_7132,N_5846);
and U8543 (N_8543,N_5039,N_7396);
or U8544 (N_8544,N_7233,N_5188);
and U8545 (N_8545,N_6171,N_5915);
and U8546 (N_8546,N_6491,N_5431);
or U8547 (N_8547,N_5855,N_6728);
nand U8548 (N_8548,N_6977,N_6534);
and U8549 (N_8549,N_7103,N_6431);
and U8550 (N_8550,N_7053,N_5828);
nand U8551 (N_8551,N_6485,N_5054);
nor U8552 (N_8552,N_5899,N_6992);
nor U8553 (N_8553,N_7156,N_7049);
nand U8554 (N_8554,N_6747,N_5170);
nor U8555 (N_8555,N_6274,N_7278);
nor U8556 (N_8556,N_5972,N_5933);
and U8557 (N_8557,N_5000,N_6763);
or U8558 (N_8558,N_7058,N_7107);
nand U8559 (N_8559,N_5095,N_6139);
nand U8560 (N_8560,N_5845,N_5420);
nor U8561 (N_8561,N_5698,N_5087);
or U8562 (N_8562,N_7426,N_5565);
nand U8563 (N_8563,N_5617,N_6062);
and U8564 (N_8564,N_7415,N_7468);
xor U8565 (N_8565,N_5133,N_6634);
and U8566 (N_8566,N_6856,N_5472);
and U8567 (N_8567,N_6620,N_6453);
or U8568 (N_8568,N_6225,N_6934);
nor U8569 (N_8569,N_5704,N_6300);
nor U8570 (N_8570,N_6058,N_5313);
and U8571 (N_8571,N_7042,N_7432);
nor U8572 (N_8572,N_6557,N_6785);
nand U8573 (N_8573,N_6449,N_5186);
nand U8574 (N_8574,N_5261,N_5779);
nand U8575 (N_8575,N_5429,N_7308);
nor U8576 (N_8576,N_6976,N_6609);
and U8577 (N_8577,N_5078,N_5048);
and U8578 (N_8578,N_6734,N_6309);
nor U8579 (N_8579,N_6879,N_7444);
and U8580 (N_8580,N_6230,N_5329);
and U8581 (N_8581,N_5571,N_5139);
and U8582 (N_8582,N_5945,N_7069);
and U8583 (N_8583,N_6477,N_5894);
nor U8584 (N_8584,N_5552,N_6269);
and U8585 (N_8585,N_5190,N_6627);
or U8586 (N_8586,N_5203,N_7271);
xnor U8587 (N_8587,N_6291,N_7328);
nor U8588 (N_8588,N_6374,N_6698);
nor U8589 (N_8589,N_6489,N_6312);
nand U8590 (N_8590,N_6057,N_5958);
and U8591 (N_8591,N_6073,N_5507);
or U8592 (N_8592,N_7492,N_7282);
and U8593 (N_8593,N_6703,N_6965);
or U8594 (N_8594,N_6962,N_6349);
nor U8595 (N_8595,N_7192,N_6216);
nor U8596 (N_8596,N_6766,N_5801);
or U8597 (N_8597,N_6341,N_5448);
or U8598 (N_8598,N_6423,N_6989);
or U8599 (N_8599,N_6469,N_5014);
xor U8600 (N_8600,N_5858,N_5538);
nand U8601 (N_8601,N_6483,N_5881);
nand U8602 (N_8602,N_5725,N_6130);
nor U8603 (N_8603,N_6051,N_6466);
nand U8604 (N_8604,N_7026,N_6648);
or U8605 (N_8605,N_6919,N_5655);
or U8606 (N_8606,N_5285,N_6577);
nand U8607 (N_8607,N_6669,N_6158);
nand U8608 (N_8608,N_5123,N_5275);
or U8609 (N_8609,N_6303,N_5628);
nor U8610 (N_8610,N_6061,N_6897);
or U8611 (N_8611,N_5983,N_5814);
nand U8612 (N_8612,N_6167,N_6878);
or U8613 (N_8613,N_6029,N_6071);
and U8614 (N_8614,N_5791,N_6145);
xor U8615 (N_8615,N_5424,N_5280);
or U8616 (N_8616,N_6327,N_6017);
or U8617 (N_8617,N_5410,N_5417);
nand U8618 (N_8618,N_6138,N_5120);
nand U8619 (N_8619,N_6484,N_5371);
nor U8620 (N_8620,N_6770,N_6964);
and U8621 (N_8621,N_5397,N_6137);
and U8622 (N_8622,N_6900,N_5888);
and U8623 (N_8623,N_5102,N_5419);
nor U8624 (N_8624,N_6606,N_7390);
nor U8625 (N_8625,N_6392,N_7382);
nor U8626 (N_8626,N_6079,N_7456);
nand U8627 (N_8627,N_6433,N_5458);
nand U8628 (N_8628,N_6798,N_6996);
or U8629 (N_8629,N_5262,N_5943);
and U8630 (N_8630,N_7499,N_7463);
and U8631 (N_8631,N_5921,N_6685);
nor U8632 (N_8632,N_5091,N_6588);
nor U8633 (N_8633,N_6321,N_7111);
nor U8634 (N_8634,N_5835,N_6510);
and U8635 (N_8635,N_6417,N_5836);
and U8636 (N_8636,N_7454,N_7472);
xor U8637 (N_8637,N_6337,N_6696);
nand U8638 (N_8638,N_5273,N_7299);
nor U8639 (N_8639,N_6290,N_5549);
nor U8640 (N_8640,N_5061,N_7043);
nor U8641 (N_8641,N_5369,N_7277);
xor U8642 (N_8642,N_7180,N_6930);
or U8643 (N_8643,N_5245,N_6727);
nor U8644 (N_8644,N_6149,N_5952);
or U8645 (N_8645,N_5541,N_5674);
nand U8646 (N_8646,N_6443,N_6813);
nand U8647 (N_8647,N_7303,N_6524);
nor U8648 (N_8648,N_5243,N_7291);
nor U8649 (N_8649,N_7381,N_5096);
nor U8650 (N_8650,N_6815,N_6678);
nand U8651 (N_8651,N_6625,N_6579);
or U8652 (N_8652,N_5977,N_7423);
or U8653 (N_8653,N_7316,N_7166);
and U8654 (N_8654,N_6803,N_5727);
and U8655 (N_8655,N_5202,N_6175);
and U8656 (N_8656,N_6882,N_5134);
nor U8657 (N_8657,N_5214,N_5480);
or U8658 (N_8658,N_5544,N_6150);
nor U8659 (N_8659,N_6851,N_7123);
or U8660 (N_8660,N_6424,N_6159);
and U8661 (N_8661,N_6865,N_6598);
nor U8662 (N_8662,N_5328,N_6956);
nand U8663 (N_8663,N_5077,N_7083);
or U8664 (N_8664,N_5859,N_5722);
or U8665 (N_8665,N_6286,N_6578);
and U8666 (N_8666,N_7191,N_5142);
and U8667 (N_8667,N_6197,N_5392);
nor U8668 (N_8668,N_5286,N_6536);
and U8669 (N_8669,N_6883,N_6636);
or U8670 (N_8670,N_5294,N_7008);
nand U8671 (N_8671,N_5497,N_7051);
or U8672 (N_8672,N_7235,N_6825);
nand U8673 (N_8673,N_6884,N_6861);
nor U8674 (N_8674,N_6784,N_5902);
or U8675 (N_8675,N_5422,N_5208);
or U8676 (N_8676,N_7270,N_5006);
xnor U8677 (N_8677,N_5158,N_5176);
and U8678 (N_8678,N_7275,N_7243);
nor U8679 (N_8679,N_7182,N_7240);
or U8680 (N_8680,N_5159,N_6391);
nand U8681 (N_8681,N_5951,N_5236);
and U8682 (N_8682,N_5557,N_6182);
nor U8683 (N_8683,N_7145,N_5658);
nor U8684 (N_8684,N_5992,N_6025);
nand U8685 (N_8685,N_6144,N_6980);
nor U8686 (N_8686,N_6503,N_6380);
and U8687 (N_8687,N_7467,N_5964);
nand U8688 (N_8688,N_6566,N_6030);
nor U8689 (N_8689,N_5955,N_6961);
or U8690 (N_8690,N_5083,N_5834);
nand U8691 (N_8691,N_5187,N_7254);
and U8692 (N_8692,N_5935,N_7030);
and U8693 (N_8693,N_5745,N_6146);
or U8694 (N_8694,N_5350,N_5047);
or U8695 (N_8695,N_7320,N_6638);
nand U8696 (N_8696,N_6316,N_6217);
xnor U8697 (N_8697,N_5705,N_5554);
and U8698 (N_8698,N_5694,N_6323);
and U8699 (N_8699,N_5184,N_6118);
xor U8700 (N_8700,N_5644,N_6540);
nor U8701 (N_8701,N_6644,N_6014);
nand U8702 (N_8702,N_7178,N_6860);
and U8703 (N_8703,N_5806,N_6744);
and U8704 (N_8704,N_6979,N_5990);
nor U8705 (N_8705,N_5900,N_6667);
nand U8706 (N_8706,N_6843,N_6147);
nor U8707 (N_8707,N_5045,N_6799);
nor U8708 (N_8708,N_6903,N_6066);
or U8709 (N_8709,N_7344,N_7339);
or U8710 (N_8710,N_5265,N_7411);
nand U8711 (N_8711,N_6952,N_7256);
and U8712 (N_8712,N_7248,N_6978);
and U8713 (N_8713,N_5278,N_7403);
or U8714 (N_8714,N_5222,N_6263);
nor U8715 (N_8715,N_5440,N_6886);
xor U8716 (N_8716,N_7031,N_7414);
nor U8717 (N_8717,N_5489,N_5484);
nor U8718 (N_8718,N_7186,N_5150);
and U8719 (N_8719,N_5110,N_6241);
xnor U8720 (N_8720,N_6533,N_6422);
or U8721 (N_8721,N_7259,N_6937);
and U8722 (N_8722,N_5887,N_5035);
nand U8723 (N_8723,N_6319,N_6227);
and U8724 (N_8724,N_7190,N_5916);
nand U8725 (N_8725,N_5525,N_5174);
nand U8726 (N_8726,N_6675,N_6408);
nor U8727 (N_8727,N_6889,N_5302);
nand U8728 (N_8728,N_7386,N_5482);
nor U8729 (N_8729,N_7088,N_6714);
xnor U8730 (N_8730,N_5585,N_5225);
and U8731 (N_8731,N_6246,N_5596);
xor U8732 (N_8732,N_6576,N_5619);
nand U8733 (N_8733,N_6070,N_7136);
and U8734 (N_8734,N_5769,N_5323);
nor U8735 (N_8735,N_5092,N_5358);
or U8736 (N_8736,N_7063,N_7399);
and U8737 (N_8737,N_7350,N_7285);
nor U8738 (N_8738,N_5770,N_5511);
nor U8739 (N_8739,N_7267,N_5523);
and U8740 (N_8740,N_5638,N_6921);
and U8741 (N_8741,N_6944,N_6642);
nor U8742 (N_8742,N_5005,N_5670);
nor U8743 (N_8743,N_6093,N_5443);
and U8744 (N_8744,N_6180,N_5467);
and U8745 (N_8745,N_7122,N_5823);
nor U8746 (N_8746,N_7071,N_5672);
and U8747 (N_8747,N_7401,N_5950);
nor U8748 (N_8748,N_7025,N_5481);
nor U8749 (N_8749,N_5799,N_7427);
and U8750 (N_8750,N_6644,N_6025);
or U8751 (N_8751,N_5949,N_6336);
and U8752 (N_8752,N_6609,N_5335);
nand U8753 (N_8753,N_6329,N_7273);
or U8754 (N_8754,N_5662,N_6720);
xor U8755 (N_8755,N_7047,N_6262);
nand U8756 (N_8756,N_5233,N_7184);
nand U8757 (N_8757,N_6024,N_7015);
and U8758 (N_8758,N_7132,N_6813);
or U8759 (N_8759,N_6611,N_6932);
and U8760 (N_8760,N_7439,N_5409);
nor U8761 (N_8761,N_5687,N_7454);
nor U8762 (N_8762,N_5954,N_7402);
or U8763 (N_8763,N_7438,N_5747);
and U8764 (N_8764,N_6683,N_6807);
or U8765 (N_8765,N_6639,N_7297);
nor U8766 (N_8766,N_6413,N_6117);
nor U8767 (N_8767,N_7018,N_7480);
nor U8768 (N_8768,N_5991,N_5021);
nand U8769 (N_8769,N_6241,N_5362);
or U8770 (N_8770,N_5370,N_6943);
xor U8771 (N_8771,N_5517,N_5450);
or U8772 (N_8772,N_6343,N_6373);
and U8773 (N_8773,N_5778,N_5649);
and U8774 (N_8774,N_5007,N_6184);
nand U8775 (N_8775,N_7298,N_6841);
nor U8776 (N_8776,N_7326,N_6304);
nand U8777 (N_8777,N_5016,N_5762);
and U8778 (N_8778,N_5920,N_6094);
or U8779 (N_8779,N_6039,N_6742);
and U8780 (N_8780,N_6188,N_7153);
or U8781 (N_8781,N_5778,N_5877);
and U8782 (N_8782,N_6961,N_7064);
or U8783 (N_8783,N_5709,N_6937);
and U8784 (N_8784,N_5166,N_5082);
or U8785 (N_8785,N_7028,N_7351);
and U8786 (N_8786,N_5847,N_6993);
nor U8787 (N_8787,N_5845,N_6160);
nor U8788 (N_8788,N_7037,N_6903);
or U8789 (N_8789,N_7190,N_6703);
and U8790 (N_8790,N_5080,N_5767);
and U8791 (N_8791,N_5735,N_7172);
or U8792 (N_8792,N_6307,N_7232);
and U8793 (N_8793,N_5271,N_7212);
nand U8794 (N_8794,N_7198,N_5125);
nor U8795 (N_8795,N_7160,N_6205);
and U8796 (N_8796,N_5330,N_5917);
and U8797 (N_8797,N_6754,N_7306);
and U8798 (N_8798,N_6827,N_5109);
nor U8799 (N_8799,N_5167,N_7024);
nor U8800 (N_8800,N_5177,N_7408);
nand U8801 (N_8801,N_6789,N_5531);
or U8802 (N_8802,N_5254,N_5121);
and U8803 (N_8803,N_5271,N_5640);
nor U8804 (N_8804,N_6949,N_5878);
nor U8805 (N_8805,N_5724,N_6540);
nor U8806 (N_8806,N_6570,N_5302);
nand U8807 (N_8807,N_6696,N_5608);
nand U8808 (N_8808,N_7026,N_6154);
nor U8809 (N_8809,N_5849,N_5906);
nand U8810 (N_8810,N_5066,N_5038);
or U8811 (N_8811,N_6762,N_6251);
nand U8812 (N_8812,N_5951,N_5078);
nand U8813 (N_8813,N_6851,N_5320);
or U8814 (N_8814,N_5334,N_5550);
or U8815 (N_8815,N_5574,N_5348);
and U8816 (N_8816,N_5996,N_7296);
nand U8817 (N_8817,N_7450,N_7273);
nand U8818 (N_8818,N_5249,N_6246);
or U8819 (N_8819,N_6574,N_5862);
or U8820 (N_8820,N_6210,N_6151);
and U8821 (N_8821,N_7385,N_5839);
nand U8822 (N_8822,N_7310,N_6689);
or U8823 (N_8823,N_5324,N_7473);
and U8824 (N_8824,N_6492,N_5000);
nand U8825 (N_8825,N_5781,N_5155);
nor U8826 (N_8826,N_5659,N_5007);
nor U8827 (N_8827,N_6719,N_5709);
nor U8828 (N_8828,N_5091,N_5262);
nand U8829 (N_8829,N_7277,N_6616);
or U8830 (N_8830,N_6977,N_6442);
nand U8831 (N_8831,N_6248,N_6392);
nand U8832 (N_8832,N_7382,N_6995);
nand U8833 (N_8833,N_7409,N_7393);
or U8834 (N_8834,N_5442,N_5606);
nand U8835 (N_8835,N_5216,N_6682);
and U8836 (N_8836,N_6931,N_7253);
nor U8837 (N_8837,N_5827,N_7001);
nor U8838 (N_8838,N_5108,N_5373);
and U8839 (N_8839,N_6829,N_6774);
or U8840 (N_8840,N_5785,N_7105);
nor U8841 (N_8841,N_6030,N_7063);
nor U8842 (N_8842,N_5085,N_5187);
or U8843 (N_8843,N_5766,N_5498);
nor U8844 (N_8844,N_6979,N_6864);
and U8845 (N_8845,N_5013,N_5340);
xnor U8846 (N_8846,N_5583,N_7168);
or U8847 (N_8847,N_5757,N_6105);
and U8848 (N_8848,N_6281,N_5945);
or U8849 (N_8849,N_7218,N_5615);
and U8850 (N_8850,N_6673,N_7413);
and U8851 (N_8851,N_5708,N_6716);
or U8852 (N_8852,N_6188,N_6536);
nor U8853 (N_8853,N_6247,N_6109);
and U8854 (N_8854,N_6637,N_5786);
nor U8855 (N_8855,N_5091,N_6154);
and U8856 (N_8856,N_6071,N_5514);
or U8857 (N_8857,N_7108,N_6224);
nor U8858 (N_8858,N_5327,N_5796);
and U8859 (N_8859,N_5480,N_5871);
and U8860 (N_8860,N_5399,N_6495);
and U8861 (N_8861,N_5885,N_5770);
and U8862 (N_8862,N_7485,N_6771);
nor U8863 (N_8863,N_5147,N_7348);
and U8864 (N_8864,N_5413,N_5061);
nand U8865 (N_8865,N_7376,N_5965);
nand U8866 (N_8866,N_7250,N_6055);
nand U8867 (N_8867,N_6546,N_6226);
nand U8868 (N_8868,N_6037,N_5214);
or U8869 (N_8869,N_6334,N_5736);
or U8870 (N_8870,N_5473,N_7160);
and U8871 (N_8871,N_6437,N_6226);
or U8872 (N_8872,N_5327,N_5927);
nor U8873 (N_8873,N_6206,N_7301);
or U8874 (N_8874,N_7233,N_5691);
or U8875 (N_8875,N_7207,N_6567);
and U8876 (N_8876,N_5748,N_5771);
nand U8877 (N_8877,N_6327,N_7004);
nand U8878 (N_8878,N_5038,N_5995);
or U8879 (N_8879,N_5017,N_5034);
or U8880 (N_8880,N_5726,N_5831);
nand U8881 (N_8881,N_6128,N_6318);
or U8882 (N_8882,N_7493,N_5234);
and U8883 (N_8883,N_5728,N_6385);
nand U8884 (N_8884,N_5390,N_6613);
nor U8885 (N_8885,N_7224,N_6116);
nand U8886 (N_8886,N_7258,N_5177);
nor U8887 (N_8887,N_6169,N_5709);
or U8888 (N_8888,N_5046,N_6735);
nor U8889 (N_8889,N_6662,N_6735);
nor U8890 (N_8890,N_6670,N_6523);
or U8891 (N_8891,N_6493,N_6299);
nand U8892 (N_8892,N_5695,N_6346);
nor U8893 (N_8893,N_5910,N_5236);
nand U8894 (N_8894,N_6127,N_6643);
nor U8895 (N_8895,N_5486,N_5793);
nor U8896 (N_8896,N_5259,N_7279);
or U8897 (N_8897,N_6027,N_6716);
and U8898 (N_8898,N_6261,N_5214);
or U8899 (N_8899,N_6547,N_5365);
or U8900 (N_8900,N_5919,N_5501);
and U8901 (N_8901,N_6215,N_5207);
and U8902 (N_8902,N_7416,N_5709);
and U8903 (N_8903,N_7192,N_6861);
or U8904 (N_8904,N_5440,N_6983);
and U8905 (N_8905,N_5566,N_6792);
nand U8906 (N_8906,N_5540,N_6597);
or U8907 (N_8907,N_5650,N_7028);
xnor U8908 (N_8908,N_6873,N_5044);
nand U8909 (N_8909,N_6586,N_7363);
or U8910 (N_8910,N_5515,N_7112);
or U8911 (N_8911,N_6713,N_7109);
and U8912 (N_8912,N_5165,N_6035);
nand U8913 (N_8913,N_5020,N_6553);
or U8914 (N_8914,N_6438,N_6215);
and U8915 (N_8915,N_5897,N_7358);
nor U8916 (N_8916,N_5988,N_6048);
or U8917 (N_8917,N_5198,N_5550);
or U8918 (N_8918,N_7422,N_5532);
nor U8919 (N_8919,N_6289,N_6097);
and U8920 (N_8920,N_5832,N_6263);
nor U8921 (N_8921,N_5206,N_5103);
nor U8922 (N_8922,N_5302,N_6151);
nand U8923 (N_8923,N_6379,N_5220);
nand U8924 (N_8924,N_6443,N_6932);
and U8925 (N_8925,N_5889,N_7179);
or U8926 (N_8926,N_5399,N_6431);
and U8927 (N_8927,N_6426,N_6241);
and U8928 (N_8928,N_5799,N_6289);
xnor U8929 (N_8929,N_6988,N_5433);
nand U8930 (N_8930,N_5038,N_5538);
nor U8931 (N_8931,N_7090,N_5364);
nand U8932 (N_8932,N_7488,N_7338);
and U8933 (N_8933,N_6160,N_5678);
or U8934 (N_8934,N_5882,N_6346);
nand U8935 (N_8935,N_6454,N_5181);
or U8936 (N_8936,N_5249,N_5755);
or U8937 (N_8937,N_7424,N_5624);
or U8938 (N_8938,N_6358,N_5847);
nor U8939 (N_8939,N_7243,N_6296);
nor U8940 (N_8940,N_6090,N_5549);
and U8941 (N_8941,N_7048,N_5557);
nor U8942 (N_8942,N_5539,N_6342);
nand U8943 (N_8943,N_6531,N_6870);
nor U8944 (N_8944,N_5494,N_6712);
and U8945 (N_8945,N_5644,N_5590);
and U8946 (N_8946,N_7299,N_5344);
nor U8947 (N_8947,N_6630,N_6121);
xnor U8948 (N_8948,N_5390,N_5004);
and U8949 (N_8949,N_6409,N_5047);
xnor U8950 (N_8950,N_6823,N_5939);
nand U8951 (N_8951,N_6444,N_7145);
nor U8952 (N_8952,N_6698,N_6162);
nand U8953 (N_8953,N_5783,N_5026);
nand U8954 (N_8954,N_6043,N_5363);
nor U8955 (N_8955,N_6835,N_6158);
or U8956 (N_8956,N_7281,N_6561);
nand U8957 (N_8957,N_5870,N_5751);
nand U8958 (N_8958,N_5316,N_6720);
xnor U8959 (N_8959,N_6228,N_6270);
nor U8960 (N_8960,N_5081,N_5134);
and U8961 (N_8961,N_7207,N_6942);
or U8962 (N_8962,N_6137,N_5656);
nor U8963 (N_8963,N_6840,N_6413);
and U8964 (N_8964,N_7077,N_6936);
nor U8965 (N_8965,N_6322,N_6730);
nand U8966 (N_8966,N_7200,N_5729);
nor U8967 (N_8967,N_5338,N_5639);
or U8968 (N_8968,N_5767,N_6673);
and U8969 (N_8969,N_6379,N_6820);
and U8970 (N_8970,N_5120,N_5360);
nand U8971 (N_8971,N_5141,N_6696);
and U8972 (N_8972,N_5023,N_7186);
or U8973 (N_8973,N_5786,N_6782);
nand U8974 (N_8974,N_5000,N_5081);
or U8975 (N_8975,N_5518,N_6103);
and U8976 (N_8976,N_6055,N_7464);
or U8977 (N_8977,N_5175,N_5689);
nand U8978 (N_8978,N_5936,N_7139);
or U8979 (N_8979,N_6274,N_6061);
and U8980 (N_8980,N_5722,N_6974);
and U8981 (N_8981,N_7459,N_6875);
nand U8982 (N_8982,N_6563,N_6807);
or U8983 (N_8983,N_7325,N_6827);
and U8984 (N_8984,N_6875,N_6522);
nor U8985 (N_8985,N_7275,N_5853);
and U8986 (N_8986,N_6824,N_7176);
nand U8987 (N_8987,N_7366,N_6397);
or U8988 (N_8988,N_6540,N_5700);
xor U8989 (N_8989,N_7363,N_5155);
nor U8990 (N_8990,N_5718,N_6594);
nand U8991 (N_8991,N_7105,N_7318);
nand U8992 (N_8992,N_5564,N_7447);
nor U8993 (N_8993,N_6956,N_5453);
nand U8994 (N_8994,N_5092,N_6656);
and U8995 (N_8995,N_5041,N_5931);
and U8996 (N_8996,N_5378,N_6066);
nor U8997 (N_8997,N_6445,N_6782);
nand U8998 (N_8998,N_7280,N_7251);
nand U8999 (N_8999,N_5554,N_7223);
or U9000 (N_9000,N_5509,N_7488);
nor U9001 (N_9001,N_7074,N_5654);
nand U9002 (N_9002,N_6667,N_6589);
or U9003 (N_9003,N_6300,N_7187);
nor U9004 (N_9004,N_5613,N_5034);
nor U9005 (N_9005,N_5804,N_5416);
xor U9006 (N_9006,N_6383,N_6979);
nor U9007 (N_9007,N_7360,N_5063);
and U9008 (N_9008,N_5520,N_7095);
nor U9009 (N_9009,N_6331,N_5631);
nor U9010 (N_9010,N_7180,N_5947);
nand U9011 (N_9011,N_5193,N_5645);
nand U9012 (N_9012,N_7342,N_7134);
or U9013 (N_9013,N_6358,N_7018);
nand U9014 (N_9014,N_5496,N_6781);
nor U9015 (N_9015,N_6473,N_5722);
nor U9016 (N_9016,N_6898,N_7438);
nor U9017 (N_9017,N_5988,N_7453);
nor U9018 (N_9018,N_5188,N_5713);
nand U9019 (N_9019,N_5754,N_6067);
nor U9020 (N_9020,N_6567,N_5872);
and U9021 (N_9021,N_5674,N_7089);
or U9022 (N_9022,N_7352,N_7274);
or U9023 (N_9023,N_5077,N_6157);
or U9024 (N_9024,N_5302,N_6768);
or U9025 (N_9025,N_5853,N_5886);
nor U9026 (N_9026,N_6205,N_5685);
nor U9027 (N_9027,N_6720,N_7029);
and U9028 (N_9028,N_5294,N_6871);
nand U9029 (N_9029,N_6415,N_5997);
or U9030 (N_9030,N_6900,N_6023);
and U9031 (N_9031,N_6140,N_6666);
nand U9032 (N_9032,N_5229,N_5417);
xnor U9033 (N_9033,N_6835,N_7240);
nor U9034 (N_9034,N_6126,N_6961);
nor U9035 (N_9035,N_5841,N_5129);
and U9036 (N_9036,N_7311,N_5390);
or U9037 (N_9037,N_5537,N_7168);
nand U9038 (N_9038,N_6576,N_7066);
or U9039 (N_9039,N_7256,N_5497);
nand U9040 (N_9040,N_7474,N_5578);
nand U9041 (N_9041,N_7388,N_6331);
and U9042 (N_9042,N_6021,N_7276);
nand U9043 (N_9043,N_6985,N_6420);
or U9044 (N_9044,N_7048,N_5565);
nand U9045 (N_9045,N_6235,N_7134);
nor U9046 (N_9046,N_6760,N_6059);
or U9047 (N_9047,N_5465,N_7229);
nand U9048 (N_9048,N_7292,N_7428);
and U9049 (N_9049,N_7149,N_5850);
nor U9050 (N_9050,N_6771,N_6564);
nor U9051 (N_9051,N_5060,N_6744);
or U9052 (N_9052,N_7377,N_5312);
or U9053 (N_9053,N_7206,N_7009);
nand U9054 (N_9054,N_6932,N_7282);
nand U9055 (N_9055,N_5287,N_5442);
and U9056 (N_9056,N_6132,N_5166);
nor U9057 (N_9057,N_6132,N_5601);
and U9058 (N_9058,N_6926,N_5342);
and U9059 (N_9059,N_6869,N_6403);
or U9060 (N_9060,N_6956,N_5014);
nand U9061 (N_9061,N_6408,N_6634);
and U9062 (N_9062,N_6981,N_5008);
and U9063 (N_9063,N_6344,N_5225);
nand U9064 (N_9064,N_5532,N_7205);
or U9065 (N_9065,N_5338,N_5805);
or U9066 (N_9066,N_6700,N_6296);
or U9067 (N_9067,N_5102,N_6037);
or U9068 (N_9068,N_7149,N_6103);
nor U9069 (N_9069,N_6990,N_5754);
nand U9070 (N_9070,N_6267,N_6002);
nand U9071 (N_9071,N_5759,N_6293);
nand U9072 (N_9072,N_6886,N_5008);
or U9073 (N_9073,N_6107,N_6824);
and U9074 (N_9074,N_6401,N_5947);
nand U9075 (N_9075,N_7247,N_5662);
and U9076 (N_9076,N_5552,N_6344);
and U9077 (N_9077,N_6083,N_7411);
and U9078 (N_9078,N_5379,N_5116);
or U9079 (N_9079,N_5225,N_5579);
nand U9080 (N_9080,N_6172,N_5484);
and U9081 (N_9081,N_5517,N_6439);
and U9082 (N_9082,N_5465,N_6397);
nand U9083 (N_9083,N_7061,N_5051);
nor U9084 (N_9084,N_7220,N_5366);
nand U9085 (N_9085,N_5090,N_5491);
and U9086 (N_9086,N_5143,N_7016);
nand U9087 (N_9087,N_5453,N_7462);
nand U9088 (N_9088,N_5349,N_7021);
nand U9089 (N_9089,N_7294,N_6739);
or U9090 (N_9090,N_5373,N_5110);
nor U9091 (N_9091,N_6288,N_6503);
and U9092 (N_9092,N_6177,N_5123);
and U9093 (N_9093,N_6373,N_6781);
and U9094 (N_9094,N_5878,N_6274);
and U9095 (N_9095,N_5675,N_6986);
nor U9096 (N_9096,N_7356,N_7236);
nor U9097 (N_9097,N_6597,N_5060);
nand U9098 (N_9098,N_7436,N_5521);
nand U9099 (N_9099,N_5300,N_5046);
xnor U9100 (N_9100,N_7453,N_7428);
nand U9101 (N_9101,N_6341,N_6633);
nand U9102 (N_9102,N_5912,N_7408);
nand U9103 (N_9103,N_5452,N_6130);
and U9104 (N_9104,N_6984,N_5564);
nand U9105 (N_9105,N_5967,N_5749);
and U9106 (N_9106,N_6754,N_5951);
nand U9107 (N_9107,N_7159,N_7108);
nor U9108 (N_9108,N_5116,N_5160);
and U9109 (N_9109,N_6685,N_5923);
and U9110 (N_9110,N_5154,N_5445);
or U9111 (N_9111,N_7153,N_7071);
or U9112 (N_9112,N_5160,N_6164);
nand U9113 (N_9113,N_6462,N_7006);
or U9114 (N_9114,N_6208,N_6306);
or U9115 (N_9115,N_5941,N_7150);
nand U9116 (N_9116,N_7475,N_5719);
and U9117 (N_9117,N_7126,N_6504);
or U9118 (N_9118,N_5825,N_6757);
nor U9119 (N_9119,N_5872,N_6681);
or U9120 (N_9120,N_5166,N_6535);
nor U9121 (N_9121,N_6233,N_7322);
nor U9122 (N_9122,N_5387,N_5698);
nor U9123 (N_9123,N_6632,N_6925);
nand U9124 (N_9124,N_5952,N_5805);
nor U9125 (N_9125,N_7181,N_5770);
or U9126 (N_9126,N_6959,N_6733);
and U9127 (N_9127,N_6363,N_7406);
nor U9128 (N_9128,N_7208,N_6258);
nand U9129 (N_9129,N_5744,N_7476);
or U9130 (N_9130,N_7004,N_5004);
nand U9131 (N_9131,N_6362,N_7124);
or U9132 (N_9132,N_7078,N_7160);
and U9133 (N_9133,N_5466,N_5609);
nand U9134 (N_9134,N_6806,N_7209);
or U9135 (N_9135,N_7024,N_5645);
nor U9136 (N_9136,N_6827,N_6651);
nor U9137 (N_9137,N_5760,N_7285);
xor U9138 (N_9138,N_5211,N_6443);
nor U9139 (N_9139,N_5316,N_5391);
or U9140 (N_9140,N_5068,N_6185);
and U9141 (N_9141,N_7142,N_6624);
nand U9142 (N_9142,N_6181,N_5266);
nand U9143 (N_9143,N_6907,N_6996);
or U9144 (N_9144,N_6355,N_6673);
nor U9145 (N_9145,N_5093,N_5981);
nor U9146 (N_9146,N_6413,N_7163);
nand U9147 (N_9147,N_6318,N_7069);
and U9148 (N_9148,N_5028,N_7030);
and U9149 (N_9149,N_5264,N_5658);
nor U9150 (N_9150,N_6669,N_7128);
or U9151 (N_9151,N_7445,N_5582);
and U9152 (N_9152,N_7101,N_5571);
nor U9153 (N_9153,N_6663,N_6054);
nand U9154 (N_9154,N_5723,N_6881);
or U9155 (N_9155,N_5736,N_6800);
or U9156 (N_9156,N_7165,N_5306);
nand U9157 (N_9157,N_5244,N_6932);
xnor U9158 (N_9158,N_7357,N_5527);
nor U9159 (N_9159,N_5467,N_6623);
and U9160 (N_9160,N_5716,N_6431);
or U9161 (N_9161,N_6205,N_7245);
or U9162 (N_9162,N_6762,N_7384);
or U9163 (N_9163,N_5346,N_5043);
and U9164 (N_9164,N_7472,N_7423);
nand U9165 (N_9165,N_6964,N_5159);
or U9166 (N_9166,N_7114,N_7117);
nand U9167 (N_9167,N_5244,N_5210);
nand U9168 (N_9168,N_6933,N_6879);
and U9169 (N_9169,N_6018,N_5946);
and U9170 (N_9170,N_5680,N_7055);
xnor U9171 (N_9171,N_5924,N_6521);
and U9172 (N_9172,N_5610,N_6452);
nor U9173 (N_9173,N_5411,N_5089);
or U9174 (N_9174,N_7321,N_5770);
or U9175 (N_9175,N_7163,N_6073);
or U9176 (N_9176,N_5864,N_5773);
nand U9177 (N_9177,N_6261,N_7160);
or U9178 (N_9178,N_6296,N_5920);
or U9179 (N_9179,N_5063,N_7372);
or U9180 (N_9180,N_7236,N_7253);
nand U9181 (N_9181,N_5229,N_5287);
nor U9182 (N_9182,N_6946,N_5070);
nand U9183 (N_9183,N_5668,N_6351);
or U9184 (N_9184,N_6340,N_5605);
nand U9185 (N_9185,N_5040,N_5050);
or U9186 (N_9186,N_6538,N_6130);
nor U9187 (N_9187,N_5286,N_6249);
and U9188 (N_9188,N_6315,N_5757);
or U9189 (N_9189,N_5022,N_6694);
or U9190 (N_9190,N_6540,N_7242);
and U9191 (N_9191,N_6158,N_5988);
and U9192 (N_9192,N_6320,N_7360);
nand U9193 (N_9193,N_6088,N_6180);
nor U9194 (N_9194,N_6023,N_6463);
nand U9195 (N_9195,N_5736,N_6431);
nor U9196 (N_9196,N_5985,N_5967);
nor U9197 (N_9197,N_7168,N_6893);
nor U9198 (N_9198,N_6237,N_5071);
nor U9199 (N_9199,N_5811,N_6523);
or U9200 (N_9200,N_5097,N_6968);
nand U9201 (N_9201,N_6989,N_7301);
xor U9202 (N_9202,N_6580,N_6203);
or U9203 (N_9203,N_7057,N_6480);
nor U9204 (N_9204,N_7235,N_5498);
and U9205 (N_9205,N_5895,N_6708);
nor U9206 (N_9206,N_6764,N_5271);
nor U9207 (N_9207,N_7480,N_5897);
nand U9208 (N_9208,N_7491,N_6820);
nand U9209 (N_9209,N_6647,N_5352);
or U9210 (N_9210,N_6231,N_5616);
or U9211 (N_9211,N_7493,N_5392);
nand U9212 (N_9212,N_5433,N_5949);
or U9213 (N_9213,N_6770,N_6629);
or U9214 (N_9214,N_7075,N_6602);
or U9215 (N_9215,N_6080,N_6927);
and U9216 (N_9216,N_6313,N_7307);
nand U9217 (N_9217,N_7167,N_5656);
and U9218 (N_9218,N_6955,N_5956);
and U9219 (N_9219,N_6959,N_6186);
nor U9220 (N_9220,N_6268,N_5756);
and U9221 (N_9221,N_6480,N_5449);
nand U9222 (N_9222,N_7209,N_5776);
or U9223 (N_9223,N_5355,N_5503);
xnor U9224 (N_9224,N_6532,N_5424);
and U9225 (N_9225,N_5980,N_7030);
and U9226 (N_9226,N_5154,N_7248);
nor U9227 (N_9227,N_5429,N_7400);
nand U9228 (N_9228,N_5272,N_5982);
nand U9229 (N_9229,N_6673,N_5788);
nor U9230 (N_9230,N_5345,N_6261);
nand U9231 (N_9231,N_5823,N_7045);
or U9232 (N_9232,N_7104,N_6466);
nor U9233 (N_9233,N_5770,N_6043);
and U9234 (N_9234,N_7226,N_6841);
and U9235 (N_9235,N_6758,N_7466);
and U9236 (N_9236,N_6060,N_6515);
and U9237 (N_9237,N_6210,N_5649);
nand U9238 (N_9238,N_7365,N_5919);
nand U9239 (N_9239,N_5386,N_6167);
nor U9240 (N_9240,N_7435,N_7375);
nor U9241 (N_9241,N_5621,N_6348);
nand U9242 (N_9242,N_5759,N_5529);
nand U9243 (N_9243,N_5216,N_6313);
and U9244 (N_9244,N_5507,N_6873);
nand U9245 (N_9245,N_5299,N_7232);
and U9246 (N_9246,N_5225,N_6271);
nor U9247 (N_9247,N_7274,N_6962);
or U9248 (N_9248,N_7304,N_6070);
or U9249 (N_9249,N_5449,N_6386);
nor U9250 (N_9250,N_6145,N_5683);
or U9251 (N_9251,N_6958,N_5946);
nand U9252 (N_9252,N_6071,N_6743);
nand U9253 (N_9253,N_5509,N_6328);
and U9254 (N_9254,N_7372,N_6520);
and U9255 (N_9255,N_7101,N_5284);
or U9256 (N_9256,N_7097,N_7300);
nor U9257 (N_9257,N_5559,N_6466);
or U9258 (N_9258,N_6764,N_6164);
and U9259 (N_9259,N_6470,N_5329);
nand U9260 (N_9260,N_6738,N_6863);
nand U9261 (N_9261,N_7067,N_5897);
nor U9262 (N_9262,N_6408,N_5821);
or U9263 (N_9263,N_6658,N_5008);
or U9264 (N_9264,N_6333,N_6210);
nand U9265 (N_9265,N_5710,N_6616);
or U9266 (N_9266,N_5073,N_5198);
and U9267 (N_9267,N_5594,N_6311);
and U9268 (N_9268,N_5395,N_6396);
or U9269 (N_9269,N_6725,N_7197);
or U9270 (N_9270,N_6217,N_6419);
and U9271 (N_9271,N_7377,N_6470);
nor U9272 (N_9272,N_6120,N_7233);
or U9273 (N_9273,N_7347,N_5340);
nand U9274 (N_9274,N_5070,N_5095);
nor U9275 (N_9275,N_6314,N_7315);
and U9276 (N_9276,N_6289,N_5358);
nand U9277 (N_9277,N_5038,N_7058);
or U9278 (N_9278,N_5583,N_5579);
nand U9279 (N_9279,N_7409,N_6495);
xor U9280 (N_9280,N_6691,N_7263);
nand U9281 (N_9281,N_5203,N_5174);
nand U9282 (N_9282,N_7025,N_6159);
nand U9283 (N_9283,N_5682,N_5539);
nand U9284 (N_9284,N_6618,N_5225);
and U9285 (N_9285,N_6917,N_5264);
nand U9286 (N_9286,N_6062,N_6773);
nor U9287 (N_9287,N_5790,N_5380);
and U9288 (N_9288,N_5639,N_6391);
nor U9289 (N_9289,N_5325,N_5866);
or U9290 (N_9290,N_5375,N_5056);
and U9291 (N_9291,N_5130,N_6333);
nand U9292 (N_9292,N_7071,N_7257);
or U9293 (N_9293,N_6813,N_6052);
nand U9294 (N_9294,N_6525,N_5129);
nand U9295 (N_9295,N_7207,N_6423);
nand U9296 (N_9296,N_6938,N_7477);
or U9297 (N_9297,N_5728,N_6677);
nand U9298 (N_9298,N_5305,N_7186);
nand U9299 (N_9299,N_5433,N_5293);
or U9300 (N_9300,N_5685,N_7206);
and U9301 (N_9301,N_5417,N_6682);
nand U9302 (N_9302,N_7391,N_5001);
xor U9303 (N_9303,N_5834,N_6518);
or U9304 (N_9304,N_5926,N_6204);
xnor U9305 (N_9305,N_7056,N_6999);
and U9306 (N_9306,N_6425,N_6917);
nor U9307 (N_9307,N_5107,N_6747);
and U9308 (N_9308,N_5852,N_7491);
nand U9309 (N_9309,N_6917,N_6937);
or U9310 (N_9310,N_6653,N_6286);
nand U9311 (N_9311,N_5493,N_6362);
nor U9312 (N_9312,N_6044,N_5013);
nor U9313 (N_9313,N_6543,N_6792);
nor U9314 (N_9314,N_6943,N_7312);
and U9315 (N_9315,N_6710,N_6754);
nand U9316 (N_9316,N_6882,N_6940);
nor U9317 (N_9317,N_6964,N_7092);
and U9318 (N_9318,N_5455,N_6710);
nor U9319 (N_9319,N_6122,N_6095);
nor U9320 (N_9320,N_6582,N_7081);
nand U9321 (N_9321,N_5330,N_5855);
nand U9322 (N_9322,N_7368,N_5517);
xnor U9323 (N_9323,N_5707,N_6716);
and U9324 (N_9324,N_6941,N_5409);
nor U9325 (N_9325,N_7154,N_7313);
and U9326 (N_9326,N_7375,N_5627);
nand U9327 (N_9327,N_5573,N_5345);
nand U9328 (N_9328,N_5784,N_7282);
and U9329 (N_9329,N_6843,N_6625);
and U9330 (N_9330,N_5511,N_5575);
nand U9331 (N_9331,N_6185,N_6723);
nor U9332 (N_9332,N_5205,N_6043);
and U9333 (N_9333,N_5575,N_5919);
nor U9334 (N_9334,N_5533,N_5632);
and U9335 (N_9335,N_6266,N_5688);
nand U9336 (N_9336,N_6794,N_7076);
nor U9337 (N_9337,N_5589,N_6851);
xor U9338 (N_9338,N_5869,N_5376);
nand U9339 (N_9339,N_6986,N_7298);
and U9340 (N_9340,N_6545,N_6539);
nand U9341 (N_9341,N_6833,N_6997);
and U9342 (N_9342,N_7429,N_6986);
nor U9343 (N_9343,N_6081,N_5496);
nand U9344 (N_9344,N_6944,N_7041);
or U9345 (N_9345,N_6681,N_6038);
and U9346 (N_9346,N_6166,N_6745);
nand U9347 (N_9347,N_7497,N_6245);
nor U9348 (N_9348,N_7140,N_7124);
or U9349 (N_9349,N_6151,N_6709);
and U9350 (N_9350,N_6277,N_5720);
nand U9351 (N_9351,N_5606,N_5744);
nor U9352 (N_9352,N_5788,N_6383);
nand U9353 (N_9353,N_6090,N_6290);
and U9354 (N_9354,N_5192,N_5734);
or U9355 (N_9355,N_5464,N_7076);
nor U9356 (N_9356,N_6603,N_5020);
nor U9357 (N_9357,N_7110,N_7193);
or U9358 (N_9358,N_7227,N_5256);
and U9359 (N_9359,N_6419,N_6448);
or U9360 (N_9360,N_7316,N_5673);
and U9361 (N_9361,N_7340,N_7421);
and U9362 (N_9362,N_5465,N_7286);
or U9363 (N_9363,N_5520,N_6912);
nor U9364 (N_9364,N_6428,N_6382);
and U9365 (N_9365,N_5902,N_5160);
and U9366 (N_9366,N_7088,N_6534);
or U9367 (N_9367,N_5572,N_6337);
or U9368 (N_9368,N_6363,N_6215);
or U9369 (N_9369,N_7140,N_5826);
or U9370 (N_9370,N_5640,N_7168);
nand U9371 (N_9371,N_6151,N_5986);
nand U9372 (N_9372,N_5242,N_7455);
nor U9373 (N_9373,N_5133,N_5300);
or U9374 (N_9374,N_5060,N_5604);
and U9375 (N_9375,N_6104,N_5945);
nor U9376 (N_9376,N_5800,N_5099);
and U9377 (N_9377,N_6107,N_5331);
nand U9378 (N_9378,N_7407,N_5394);
nor U9379 (N_9379,N_5741,N_7449);
or U9380 (N_9380,N_6694,N_6593);
or U9381 (N_9381,N_5495,N_6466);
nor U9382 (N_9382,N_6119,N_6185);
and U9383 (N_9383,N_5810,N_5805);
nand U9384 (N_9384,N_6336,N_6539);
or U9385 (N_9385,N_6353,N_5185);
nor U9386 (N_9386,N_5404,N_5115);
nand U9387 (N_9387,N_6647,N_6054);
nand U9388 (N_9388,N_6658,N_5740);
nand U9389 (N_9389,N_6124,N_6094);
nand U9390 (N_9390,N_6317,N_6851);
or U9391 (N_9391,N_5550,N_5630);
and U9392 (N_9392,N_7240,N_6103);
or U9393 (N_9393,N_7386,N_6465);
nand U9394 (N_9394,N_6103,N_5646);
nor U9395 (N_9395,N_6581,N_6133);
nor U9396 (N_9396,N_7022,N_6523);
and U9397 (N_9397,N_7215,N_5416);
or U9398 (N_9398,N_5856,N_7451);
nor U9399 (N_9399,N_5469,N_5098);
and U9400 (N_9400,N_6054,N_7091);
and U9401 (N_9401,N_5434,N_6848);
or U9402 (N_9402,N_5114,N_7062);
and U9403 (N_9403,N_6397,N_6727);
nor U9404 (N_9404,N_7358,N_6244);
nand U9405 (N_9405,N_5235,N_6275);
nand U9406 (N_9406,N_6420,N_6469);
or U9407 (N_9407,N_6329,N_6565);
nand U9408 (N_9408,N_6569,N_5467);
nor U9409 (N_9409,N_6306,N_6805);
and U9410 (N_9410,N_5632,N_5599);
nor U9411 (N_9411,N_5517,N_6353);
or U9412 (N_9412,N_6351,N_7332);
and U9413 (N_9413,N_5320,N_6427);
nand U9414 (N_9414,N_6443,N_6216);
nand U9415 (N_9415,N_6340,N_6762);
nand U9416 (N_9416,N_5244,N_7245);
nor U9417 (N_9417,N_5813,N_6440);
nor U9418 (N_9418,N_5606,N_7448);
or U9419 (N_9419,N_5798,N_7160);
or U9420 (N_9420,N_5505,N_5063);
nand U9421 (N_9421,N_6347,N_6272);
nand U9422 (N_9422,N_6557,N_7474);
nand U9423 (N_9423,N_5782,N_5002);
nor U9424 (N_9424,N_5086,N_7270);
nand U9425 (N_9425,N_7142,N_5618);
or U9426 (N_9426,N_5640,N_7097);
and U9427 (N_9427,N_7026,N_5328);
and U9428 (N_9428,N_5090,N_7175);
and U9429 (N_9429,N_7301,N_6469);
nor U9430 (N_9430,N_7488,N_5174);
or U9431 (N_9431,N_6743,N_5511);
nor U9432 (N_9432,N_6918,N_6201);
nor U9433 (N_9433,N_7101,N_5938);
nor U9434 (N_9434,N_6779,N_6520);
or U9435 (N_9435,N_6724,N_6363);
nand U9436 (N_9436,N_7264,N_6780);
and U9437 (N_9437,N_5423,N_5910);
nor U9438 (N_9438,N_6516,N_5613);
or U9439 (N_9439,N_7328,N_7318);
nand U9440 (N_9440,N_6971,N_6476);
and U9441 (N_9441,N_5278,N_7071);
or U9442 (N_9442,N_6537,N_5023);
or U9443 (N_9443,N_7267,N_7083);
and U9444 (N_9444,N_6757,N_6460);
or U9445 (N_9445,N_6235,N_6306);
and U9446 (N_9446,N_5995,N_7330);
nand U9447 (N_9447,N_5795,N_7170);
or U9448 (N_9448,N_5354,N_6750);
or U9449 (N_9449,N_6262,N_6527);
xor U9450 (N_9450,N_5467,N_5383);
and U9451 (N_9451,N_6194,N_7421);
nor U9452 (N_9452,N_5744,N_5947);
and U9453 (N_9453,N_7211,N_7461);
nand U9454 (N_9454,N_6393,N_7457);
or U9455 (N_9455,N_5543,N_5704);
and U9456 (N_9456,N_6797,N_6427);
and U9457 (N_9457,N_6460,N_7424);
and U9458 (N_9458,N_5099,N_5827);
or U9459 (N_9459,N_5821,N_7300);
nand U9460 (N_9460,N_5072,N_7055);
and U9461 (N_9461,N_6678,N_5461);
xor U9462 (N_9462,N_5080,N_7388);
xor U9463 (N_9463,N_7247,N_7230);
or U9464 (N_9464,N_5223,N_5775);
nor U9465 (N_9465,N_5933,N_7069);
nor U9466 (N_9466,N_5599,N_6831);
nand U9467 (N_9467,N_5805,N_6814);
nand U9468 (N_9468,N_6740,N_7418);
or U9469 (N_9469,N_6469,N_5887);
nand U9470 (N_9470,N_6638,N_5117);
nand U9471 (N_9471,N_6612,N_6516);
or U9472 (N_9472,N_5056,N_5172);
nor U9473 (N_9473,N_6057,N_5316);
and U9474 (N_9474,N_7316,N_5220);
or U9475 (N_9475,N_5558,N_7369);
or U9476 (N_9476,N_5909,N_5647);
and U9477 (N_9477,N_6710,N_7246);
nor U9478 (N_9478,N_5898,N_5559);
and U9479 (N_9479,N_6503,N_6624);
nor U9480 (N_9480,N_5445,N_6741);
nor U9481 (N_9481,N_6757,N_5046);
nand U9482 (N_9482,N_6419,N_5056);
and U9483 (N_9483,N_5462,N_7321);
nand U9484 (N_9484,N_5102,N_5878);
or U9485 (N_9485,N_5975,N_5105);
or U9486 (N_9486,N_7478,N_6073);
nand U9487 (N_9487,N_5358,N_6808);
and U9488 (N_9488,N_6279,N_5036);
nand U9489 (N_9489,N_5987,N_5067);
nor U9490 (N_9490,N_5691,N_5122);
nand U9491 (N_9491,N_5046,N_5290);
nand U9492 (N_9492,N_7489,N_5729);
xor U9493 (N_9493,N_6661,N_5740);
nor U9494 (N_9494,N_7487,N_6148);
nand U9495 (N_9495,N_5309,N_5108);
nand U9496 (N_9496,N_6557,N_5141);
and U9497 (N_9497,N_7163,N_7213);
or U9498 (N_9498,N_5991,N_6172);
nor U9499 (N_9499,N_6331,N_7269);
and U9500 (N_9500,N_7108,N_6547);
or U9501 (N_9501,N_5671,N_5804);
or U9502 (N_9502,N_6774,N_5888);
or U9503 (N_9503,N_6273,N_5050);
and U9504 (N_9504,N_6309,N_5543);
and U9505 (N_9505,N_7098,N_6207);
nand U9506 (N_9506,N_6351,N_7108);
nor U9507 (N_9507,N_6300,N_6428);
nand U9508 (N_9508,N_5382,N_5094);
xor U9509 (N_9509,N_5543,N_5007);
or U9510 (N_9510,N_6664,N_5392);
and U9511 (N_9511,N_5004,N_5426);
or U9512 (N_9512,N_6186,N_6902);
and U9513 (N_9513,N_5291,N_7459);
nand U9514 (N_9514,N_6108,N_6641);
nand U9515 (N_9515,N_5474,N_5238);
nor U9516 (N_9516,N_5658,N_6893);
and U9517 (N_9517,N_5392,N_5329);
nand U9518 (N_9518,N_5701,N_5821);
and U9519 (N_9519,N_6950,N_6566);
nand U9520 (N_9520,N_5227,N_6960);
nor U9521 (N_9521,N_6655,N_7474);
or U9522 (N_9522,N_5870,N_7061);
or U9523 (N_9523,N_5589,N_5884);
nand U9524 (N_9524,N_6975,N_5289);
nor U9525 (N_9525,N_6988,N_6557);
and U9526 (N_9526,N_6217,N_6479);
or U9527 (N_9527,N_7329,N_5931);
and U9528 (N_9528,N_7342,N_6926);
and U9529 (N_9529,N_7256,N_7153);
and U9530 (N_9530,N_7498,N_5121);
or U9531 (N_9531,N_6132,N_6706);
nand U9532 (N_9532,N_5166,N_7345);
xor U9533 (N_9533,N_6823,N_6068);
nand U9534 (N_9534,N_5545,N_5003);
nor U9535 (N_9535,N_7007,N_5397);
nor U9536 (N_9536,N_5061,N_7231);
or U9537 (N_9537,N_7244,N_7019);
or U9538 (N_9538,N_6792,N_5912);
nor U9539 (N_9539,N_7235,N_5177);
nor U9540 (N_9540,N_5869,N_6279);
nand U9541 (N_9541,N_6761,N_5762);
nor U9542 (N_9542,N_7437,N_7235);
nand U9543 (N_9543,N_6562,N_7260);
or U9544 (N_9544,N_5805,N_5512);
or U9545 (N_9545,N_5967,N_6486);
and U9546 (N_9546,N_5511,N_5126);
or U9547 (N_9547,N_6097,N_6152);
nand U9548 (N_9548,N_5521,N_7420);
or U9549 (N_9549,N_5246,N_6025);
or U9550 (N_9550,N_6444,N_7038);
nor U9551 (N_9551,N_7239,N_5811);
or U9552 (N_9552,N_5323,N_5634);
nand U9553 (N_9553,N_5344,N_6404);
nand U9554 (N_9554,N_6114,N_7238);
and U9555 (N_9555,N_5158,N_7454);
or U9556 (N_9556,N_5203,N_5510);
or U9557 (N_9557,N_5841,N_6253);
or U9558 (N_9558,N_5353,N_5022);
and U9559 (N_9559,N_7065,N_5367);
nand U9560 (N_9560,N_5608,N_6223);
or U9561 (N_9561,N_5562,N_6680);
nand U9562 (N_9562,N_6978,N_6182);
nor U9563 (N_9563,N_7376,N_6527);
and U9564 (N_9564,N_5042,N_6337);
nor U9565 (N_9565,N_5898,N_5892);
nor U9566 (N_9566,N_6221,N_5748);
nand U9567 (N_9567,N_6196,N_5659);
or U9568 (N_9568,N_5184,N_6395);
nor U9569 (N_9569,N_6080,N_6307);
or U9570 (N_9570,N_6574,N_6493);
nand U9571 (N_9571,N_6924,N_5582);
nor U9572 (N_9572,N_6035,N_6434);
or U9573 (N_9573,N_5253,N_6623);
and U9574 (N_9574,N_5280,N_6530);
or U9575 (N_9575,N_7474,N_6187);
or U9576 (N_9576,N_5858,N_5881);
xnor U9577 (N_9577,N_7081,N_6331);
and U9578 (N_9578,N_6580,N_5813);
or U9579 (N_9579,N_5990,N_5044);
nor U9580 (N_9580,N_6733,N_6267);
nand U9581 (N_9581,N_5730,N_5179);
nor U9582 (N_9582,N_6864,N_7456);
nand U9583 (N_9583,N_6288,N_5039);
and U9584 (N_9584,N_6674,N_6540);
nor U9585 (N_9585,N_5300,N_7187);
or U9586 (N_9586,N_5583,N_6515);
nand U9587 (N_9587,N_5109,N_5196);
and U9588 (N_9588,N_5796,N_5227);
nand U9589 (N_9589,N_5434,N_7035);
or U9590 (N_9590,N_6725,N_5538);
nand U9591 (N_9591,N_6967,N_5354);
nand U9592 (N_9592,N_7223,N_7017);
xnor U9593 (N_9593,N_7300,N_7122);
and U9594 (N_9594,N_6065,N_6254);
nor U9595 (N_9595,N_5337,N_6337);
nand U9596 (N_9596,N_6908,N_5662);
xnor U9597 (N_9597,N_6286,N_7495);
and U9598 (N_9598,N_5010,N_6046);
and U9599 (N_9599,N_5968,N_7484);
or U9600 (N_9600,N_7237,N_5362);
nor U9601 (N_9601,N_6732,N_6431);
or U9602 (N_9602,N_6987,N_5607);
or U9603 (N_9603,N_6427,N_5024);
nand U9604 (N_9604,N_5309,N_6033);
nand U9605 (N_9605,N_6831,N_6054);
nand U9606 (N_9606,N_5370,N_5222);
or U9607 (N_9607,N_5961,N_6972);
and U9608 (N_9608,N_5796,N_6956);
nand U9609 (N_9609,N_5160,N_6262);
and U9610 (N_9610,N_5803,N_5609);
nor U9611 (N_9611,N_6097,N_7086);
and U9612 (N_9612,N_6384,N_7062);
nand U9613 (N_9613,N_5637,N_7361);
nor U9614 (N_9614,N_6803,N_5226);
and U9615 (N_9615,N_6386,N_6414);
nand U9616 (N_9616,N_7365,N_5418);
and U9617 (N_9617,N_5517,N_7230);
and U9618 (N_9618,N_6528,N_6803);
nand U9619 (N_9619,N_5295,N_6324);
nand U9620 (N_9620,N_5318,N_7390);
nor U9621 (N_9621,N_5836,N_7400);
nand U9622 (N_9622,N_7084,N_6854);
and U9623 (N_9623,N_6685,N_5268);
or U9624 (N_9624,N_7359,N_7425);
nor U9625 (N_9625,N_6119,N_7206);
nand U9626 (N_9626,N_7187,N_5727);
nor U9627 (N_9627,N_7264,N_6706);
and U9628 (N_9628,N_5344,N_6354);
and U9629 (N_9629,N_6972,N_5119);
and U9630 (N_9630,N_5484,N_5093);
nand U9631 (N_9631,N_6920,N_5190);
nand U9632 (N_9632,N_6359,N_6291);
nand U9633 (N_9633,N_6242,N_6222);
and U9634 (N_9634,N_5405,N_5143);
and U9635 (N_9635,N_5486,N_7202);
or U9636 (N_9636,N_5272,N_7321);
or U9637 (N_9637,N_6191,N_7035);
nand U9638 (N_9638,N_5896,N_6327);
nand U9639 (N_9639,N_5889,N_5298);
nor U9640 (N_9640,N_5200,N_5572);
or U9641 (N_9641,N_6611,N_6722);
nand U9642 (N_9642,N_6136,N_6664);
nor U9643 (N_9643,N_5764,N_5711);
and U9644 (N_9644,N_7462,N_6587);
nand U9645 (N_9645,N_6376,N_6307);
nand U9646 (N_9646,N_5383,N_6741);
or U9647 (N_9647,N_6876,N_6319);
nand U9648 (N_9648,N_5036,N_5966);
nand U9649 (N_9649,N_5497,N_5470);
and U9650 (N_9650,N_5081,N_7237);
nor U9651 (N_9651,N_5669,N_5889);
or U9652 (N_9652,N_6275,N_6038);
and U9653 (N_9653,N_6412,N_6073);
and U9654 (N_9654,N_5308,N_7036);
nand U9655 (N_9655,N_7357,N_7028);
or U9656 (N_9656,N_5182,N_6639);
or U9657 (N_9657,N_5255,N_6418);
nor U9658 (N_9658,N_6123,N_7016);
nand U9659 (N_9659,N_5839,N_5454);
and U9660 (N_9660,N_6402,N_6794);
nor U9661 (N_9661,N_5184,N_5676);
or U9662 (N_9662,N_6410,N_7359);
or U9663 (N_9663,N_6944,N_5303);
nand U9664 (N_9664,N_6342,N_5853);
nand U9665 (N_9665,N_5304,N_5553);
or U9666 (N_9666,N_7225,N_6528);
nand U9667 (N_9667,N_5019,N_7266);
or U9668 (N_9668,N_5958,N_5050);
xnor U9669 (N_9669,N_7043,N_5382);
nand U9670 (N_9670,N_6260,N_6567);
or U9671 (N_9671,N_7387,N_6365);
and U9672 (N_9672,N_6117,N_5157);
nor U9673 (N_9673,N_5839,N_5180);
nand U9674 (N_9674,N_5996,N_6230);
nand U9675 (N_9675,N_5220,N_6679);
or U9676 (N_9676,N_5024,N_7102);
and U9677 (N_9677,N_6373,N_5904);
nand U9678 (N_9678,N_6516,N_5570);
and U9679 (N_9679,N_6403,N_5784);
or U9680 (N_9680,N_6095,N_6406);
nand U9681 (N_9681,N_5305,N_6247);
and U9682 (N_9682,N_7246,N_6288);
or U9683 (N_9683,N_6692,N_5198);
xor U9684 (N_9684,N_6454,N_6429);
nand U9685 (N_9685,N_5395,N_6375);
and U9686 (N_9686,N_6494,N_5257);
or U9687 (N_9687,N_6315,N_6264);
nor U9688 (N_9688,N_5856,N_5114);
and U9689 (N_9689,N_6819,N_5544);
nand U9690 (N_9690,N_5761,N_7394);
xnor U9691 (N_9691,N_5765,N_6827);
and U9692 (N_9692,N_5912,N_6017);
or U9693 (N_9693,N_5099,N_5239);
nand U9694 (N_9694,N_7349,N_7272);
nand U9695 (N_9695,N_6194,N_6536);
nand U9696 (N_9696,N_7185,N_5727);
and U9697 (N_9697,N_6167,N_6039);
nand U9698 (N_9698,N_6537,N_5561);
nor U9699 (N_9699,N_7421,N_6225);
nor U9700 (N_9700,N_5882,N_5164);
nand U9701 (N_9701,N_6484,N_7457);
nand U9702 (N_9702,N_7080,N_7454);
nor U9703 (N_9703,N_5658,N_7479);
nand U9704 (N_9704,N_7269,N_6654);
nand U9705 (N_9705,N_5930,N_5895);
or U9706 (N_9706,N_6210,N_5068);
nor U9707 (N_9707,N_5174,N_5101);
xor U9708 (N_9708,N_7166,N_5385);
or U9709 (N_9709,N_7408,N_6479);
nor U9710 (N_9710,N_6910,N_5665);
or U9711 (N_9711,N_6275,N_7140);
nor U9712 (N_9712,N_7486,N_7345);
nor U9713 (N_9713,N_6143,N_5333);
and U9714 (N_9714,N_7235,N_7109);
or U9715 (N_9715,N_7189,N_5787);
and U9716 (N_9716,N_5162,N_6148);
and U9717 (N_9717,N_6491,N_6831);
nand U9718 (N_9718,N_5178,N_5772);
and U9719 (N_9719,N_5478,N_5443);
xnor U9720 (N_9720,N_5418,N_6085);
nor U9721 (N_9721,N_5303,N_5477);
or U9722 (N_9722,N_7270,N_6363);
nor U9723 (N_9723,N_6881,N_6887);
nand U9724 (N_9724,N_5599,N_6807);
and U9725 (N_9725,N_6147,N_6447);
and U9726 (N_9726,N_7282,N_7009);
nor U9727 (N_9727,N_6986,N_6600);
nand U9728 (N_9728,N_5853,N_5045);
and U9729 (N_9729,N_5618,N_6128);
nor U9730 (N_9730,N_5186,N_6742);
or U9731 (N_9731,N_6790,N_6233);
and U9732 (N_9732,N_6366,N_6799);
xnor U9733 (N_9733,N_5917,N_6131);
nand U9734 (N_9734,N_6462,N_5624);
or U9735 (N_9735,N_6010,N_6668);
nor U9736 (N_9736,N_6641,N_7052);
nand U9737 (N_9737,N_6918,N_6907);
xor U9738 (N_9738,N_5950,N_6378);
and U9739 (N_9739,N_6610,N_5635);
nor U9740 (N_9740,N_7199,N_5390);
nand U9741 (N_9741,N_6104,N_5147);
nand U9742 (N_9742,N_5958,N_6027);
xnor U9743 (N_9743,N_5730,N_6591);
or U9744 (N_9744,N_6545,N_6115);
xnor U9745 (N_9745,N_7297,N_5679);
nor U9746 (N_9746,N_6469,N_7045);
nand U9747 (N_9747,N_5989,N_7498);
and U9748 (N_9748,N_6046,N_5768);
and U9749 (N_9749,N_5490,N_7285);
and U9750 (N_9750,N_6738,N_6866);
nor U9751 (N_9751,N_5922,N_7484);
nor U9752 (N_9752,N_6366,N_6591);
nor U9753 (N_9753,N_5897,N_5059);
and U9754 (N_9754,N_5125,N_6933);
nand U9755 (N_9755,N_5596,N_5331);
nor U9756 (N_9756,N_6392,N_6764);
xnor U9757 (N_9757,N_6532,N_5087);
or U9758 (N_9758,N_7400,N_6966);
nor U9759 (N_9759,N_5455,N_5850);
nand U9760 (N_9760,N_7199,N_7104);
nand U9761 (N_9761,N_5961,N_6160);
or U9762 (N_9762,N_6628,N_7197);
and U9763 (N_9763,N_5874,N_6192);
nor U9764 (N_9764,N_7378,N_7251);
nand U9765 (N_9765,N_5661,N_6089);
and U9766 (N_9766,N_5216,N_7152);
and U9767 (N_9767,N_5940,N_6954);
nand U9768 (N_9768,N_5401,N_5735);
nor U9769 (N_9769,N_6393,N_6936);
nor U9770 (N_9770,N_5034,N_6721);
or U9771 (N_9771,N_7371,N_6407);
and U9772 (N_9772,N_6681,N_6562);
and U9773 (N_9773,N_6002,N_7144);
or U9774 (N_9774,N_6845,N_5046);
nand U9775 (N_9775,N_5087,N_5372);
or U9776 (N_9776,N_6587,N_6958);
nand U9777 (N_9777,N_6132,N_7414);
or U9778 (N_9778,N_5909,N_7364);
or U9779 (N_9779,N_6482,N_6695);
and U9780 (N_9780,N_5249,N_5059);
nor U9781 (N_9781,N_6832,N_5022);
nand U9782 (N_9782,N_5003,N_5184);
nand U9783 (N_9783,N_5061,N_7449);
or U9784 (N_9784,N_7326,N_7417);
or U9785 (N_9785,N_6952,N_5772);
nand U9786 (N_9786,N_6725,N_6291);
or U9787 (N_9787,N_7176,N_5985);
and U9788 (N_9788,N_6714,N_5120);
or U9789 (N_9789,N_5510,N_6897);
or U9790 (N_9790,N_5454,N_5678);
or U9791 (N_9791,N_5823,N_5362);
nand U9792 (N_9792,N_7230,N_6947);
nand U9793 (N_9793,N_5528,N_7451);
nor U9794 (N_9794,N_6744,N_5529);
xor U9795 (N_9795,N_6447,N_6029);
and U9796 (N_9796,N_5456,N_7491);
and U9797 (N_9797,N_5204,N_6992);
and U9798 (N_9798,N_6099,N_5886);
and U9799 (N_9799,N_5241,N_6263);
nor U9800 (N_9800,N_5278,N_7321);
nor U9801 (N_9801,N_6587,N_5396);
nand U9802 (N_9802,N_5541,N_5706);
nand U9803 (N_9803,N_6415,N_6942);
or U9804 (N_9804,N_6921,N_5913);
nand U9805 (N_9805,N_7267,N_7257);
xnor U9806 (N_9806,N_5685,N_6462);
xnor U9807 (N_9807,N_6683,N_6977);
or U9808 (N_9808,N_5319,N_7451);
or U9809 (N_9809,N_5554,N_6381);
or U9810 (N_9810,N_6925,N_6939);
and U9811 (N_9811,N_7346,N_5026);
nand U9812 (N_9812,N_6381,N_7143);
nand U9813 (N_9813,N_5534,N_7242);
and U9814 (N_9814,N_6587,N_6994);
nor U9815 (N_9815,N_6860,N_6315);
nand U9816 (N_9816,N_6471,N_6822);
nor U9817 (N_9817,N_5047,N_5454);
nor U9818 (N_9818,N_5143,N_5615);
or U9819 (N_9819,N_5635,N_7086);
nand U9820 (N_9820,N_5603,N_5192);
nand U9821 (N_9821,N_5007,N_6327);
and U9822 (N_9822,N_7106,N_7201);
or U9823 (N_9823,N_5582,N_5726);
nor U9824 (N_9824,N_5463,N_7462);
and U9825 (N_9825,N_5016,N_6096);
and U9826 (N_9826,N_6704,N_6602);
or U9827 (N_9827,N_6895,N_7477);
nor U9828 (N_9828,N_6770,N_5251);
nand U9829 (N_9829,N_5344,N_6125);
and U9830 (N_9830,N_5169,N_6313);
nand U9831 (N_9831,N_6575,N_7334);
nor U9832 (N_9832,N_7159,N_6156);
or U9833 (N_9833,N_7257,N_6951);
nor U9834 (N_9834,N_6416,N_5231);
nand U9835 (N_9835,N_6479,N_5839);
nor U9836 (N_9836,N_6819,N_6592);
nor U9837 (N_9837,N_5106,N_5488);
and U9838 (N_9838,N_6507,N_6171);
nor U9839 (N_9839,N_6893,N_6053);
and U9840 (N_9840,N_5763,N_6753);
or U9841 (N_9841,N_6281,N_5298);
or U9842 (N_9842,N_7454,N_5563);
and U9843 (N_9843,N_6597,N_5621);
and U9844 (N_9844,N_6409,N_7272);
nand U9845 (N_9845,N_6089,N_6724);
nand U9846 (N_9846,N_6380,N_5910);
nor U9847 (N_9847,N_6072,N_6859);
and U9848 (N_9848,N_6230,N_5573);
or U9849 (N_9849,N_6378,N_7084);
nand U9850 (N_9850,N_6843,N_6840);
or U9851 (N_9851,N_6190,N_7109);
nand U9852 (N_9852,N_5342,N_6086);
or U9853 (N_9853,N_7114,N_5041);
or U9854 (N_9854,N_6525,N_5268);
or U9855 (N_9855,N_6559,N_5066);
or U9856 (N_9856,N_7459,N_6082);
nor U9857 (N_9857,N_5547,N_6457);
xor U9858 (N_9858,N_6372,N_7187);
or U9859 (N_9859,N_5072,N_5706);
and U9860 (N_9860,N_6233,N_5573);
and U9861 (N_9861,N_7053,N_6894);
and U9862 (N_9862,N_5704,N_5461);
nand U9863 (N_9863,N_6797,N_6121);
or U9864 (N_9864,N_5812,N_5452);
and U9865 (N_9865,N_5857,N_6735);
or U9866 (N_9866,N_6653,N_7464);
nand U9867 (N_9867,N_5834,N_6299);
nand U9868 (N_9868,N_7127,N_5016);
nor U9869 (N_9869,N_5108,N_5853);
xnor U9870 (N_9870,N_5733,N_5788);
or U9871 (N_9871,N_6916,N_5154);
and U9872 (N_9872,N_6051,N_6533);
or U9873 (N_9873,N_6158,N_5501);
nand U9874 (N_9874,N_5639,N_6191);
nor U9875 (N_9875,N_5722,N_5689);
nand U9876 (N_9876,N_7012,N_6800);
and U9877 (N_9877,N_6646,N_7303);
nor U9878 (N_9878,N_6745,N_6821);
or U9879 (N_9879,N_7047,N_5689);
and U9880 (N_9880,N_5052,N_6387);
nor U9881 (N_9881,N_5110,N_5023);
and U9882 (N_9882,N_7340,N_5935);
and U9883 (N_9883,N_6037,N_5371);
or U9884 (N_9884,N_5200,N_7143);
nand U9885 (N_9885,N_5622,N_7369);
or U9886 (N_9886,N_6183,N_5732);
and U9887 (N_9887,N_5943,N_7343);
nor U9888 (N_9888,N_6221,N_7047);
nor U9889 (N_9889,N_7446,N_5068);
and U9890 (N_9890,N_5190,N_5707);
nand U9891 (N_9891,N_5272,N_5791);
or U9892 (N_9892,N_5132,N_6464);
xnor U9893 (N_9893,N_6195,N_6016);
nand U9894 (N_9894,N_6133,N_5547);
or U9895 (N_9895,N_7277,N_5642);
or U9896 (N_9896,N_5213,N_6965);
nor U9897 (N_9897,N_6324,N_5890);
nand U9898 (N_9898,N_6380,N_7493);
or U9899 (N_9899,N_5722,N_5565);
nor U9900 (N_9900,N_6784,N_6577);
nand U9901 (N_9901,N_5899,N_6845);
nand U9902 (N_9902,N_6635,N_6420);
nand U9903 (N_9903,N_7205,N_7291);
or U9904 (N_9904,N_5364,N_5796);
nand U9905 (N_9905,N_7461,N_7199);
or U9906 (N_9906,N_6757,N_7306);
or U9907 (N_9907,N_6406,N_6423);
nand U9908 (N_9908,N_5216,N_5283);
or U9909 (N_9909,N_5661,N_6291);
or U9910 (N_9910,N_7183,N_6136);
and U9911 (N_9911,N_7296,N_6355);
and U9912 (N_9912,N_5563,N_5769);
nor U9913 (N_9913,N_6863,N_7161);
nand U9914 (N_9914,N_5873,N_6333);
nand U9915 (N_9915,N_5588,N_6280);
or U9916 (N_9916,N_7058,N_7010);
or U9917 (N_9917,N_5845,N_6632);
nor U9918 (N_9918,N_6194,N_7261);
and U9919 (N_9919,N_7176,N_6280);
and U9920 (N_9920,N_6738,N_5287);
nand U9921 (N_9921,N_6223,N_5034);
nor U9922 (N_9922,N_7128,N_5816);
nor U9923 (N_9923,N_5378,N_5115);
and U9924 (N_9924,N_7447,N_6509);
and U9925 (N_9925,N_5889,N_6822);
and U9926 (N_9926,N_5189,N_6478);
nor U9927 (N_9927,N_6513,N_7031);
nor U9928 (N_9928,N_7201,N_7499);
xnor U9929 (N_9929,N_5113,N_6749);
and U9930 (N_9930,N_6080,N_6824);
or U9931 (N_9931,N_6264,N_6053);
nor U9932 (N_9932,N_7120,N_5696);
nand U9933 (N_9933,N_5734,N_6087);
or U9934 (N_9934,N_6546,N_5019);
and U9935 (N_9935,N_6719,N_7379);
and U9936 (N_9936,N_5929,N_6215);
nor U9937 (N_9937,N_5811,N_6675);
or U9938 (N_9938,N_6384,N_5853);
and U9939 (N_9939,N_6280,N_7128);
or U9940 (N_9940,N_5664,N_6666);
or U9941 (N_9941,N_6282,N_6911);
nand U9942 (N_9942,N_7036,N_5625);
nand U9943 (N_9943,N_7407,N_5724);
or U9944 (N_9944,N_6618,N_6306);
or U9945 (N_9945,N_5604,N_5626);
and U9946 (N_9946,N_6207,N_5296);
nor U9947 (N_9947,N_5392,N_6773);
xnor U9948 (N_9948,N_6863,N_5496);
and U9949 (N_9949,N_5738,N_5076);
and U9950 (N_9950,N_5149,N_6236);
nor U9951 (N_9951,N_7437,N_5124);
and U9952 (N_9952,N_5989,N_5707);
and U9953 (N_9953,N_5306,N_6449);
nor U9954 (N_9954,N_6582,N_5603);
nand U9955 (N_9955,N_5090,N_6715);
nand U9956 (N_9956,N_6027,N_6244);
nand U9957 (N_9957,N_5037,N_5670);
nand U9958 (N_9958,N_5125,N_5071);
xnor U9959 (N_9959,N_6651,N_6543);
and U9960 (N_9960,N_5584,N_5730);
and U9961 (N_9961,N_5765,N_5256);
and U9962 (N_9962,N_5853,N_6655);
nand U9963 (N_9963,N_5464,N_6705);
and U9964 (N_9964,N_6804,N_5105);
nand U9965 (N_9965,N_5531,N_6910);
nand U9966 (N_9966,N_5272,N_6094);
nor U9967 (N_9967,N_6513,N_5014);
and U9968 (N_9968,N_6498,N_6527);
nor U9969 (N_9969,N_5550,N_6293);
nand U9970 (N_9970,N_7028,N_5514);
nor U9971 (N_9971,N_5891,N_6841);
xor U9972 (N_9972,N_7320,N_5896);
or U9973 (N_9973,N_6782,N_7082);
nand U9974 (N_9974,N_7088,N_5279);
nor U9975 (N_9975,N_5767,N_7104);
nand U9976 (N_9976,N_5473,N_6399);
nor U9977 (N_9977,N_6945,N_5994);
nand U9978 (N_9978,N_5667,N_6223);
or U9979 (N_9979,N_6636,N_5266);
and U9980 (N_9980,N_5223,N_5573);
nor U9981 (N_9981,N_6254,N_6232);
xnor U9982 (N_9982,N_7193,N_5142);
or U9983 (N_9983,N_6637,N_6983);
xnor U9984 (N_9984,N_6420,N_6973);
nand U9985 (N_9985,N_6127,N_6542);
or U9986 (N_9986,N_6369,N_7032);
nand U9987 (N_9987,N_7172,N_6447);
or U9988 (N_9988,N_6440,N_6323);
or U9989 (N_9989,N_5954,N_6149);
nor U9990 (N_9990,N_7301,N_5757);
nand U9991 (N_9991,N_6265,N_5030);
nor U9992 (N_9992,N_7484,N_5937);
or U9993 (N_9993,N_5142,N_7363);
nor U9994 (N_9994,N_6741,N_7443);
or U9995 (N_9995,N_5020,N_5097);
nor U9996 (N_9996,N_6432,N_5693);
nor U9997 (N_9997,N_5585,N_5005);
and U9998 (N_9998,N_7123,N_5469);
nor U9999 (N_9999,N_7163,N_5215);
or UO_0 (O_0,N_7917,N_9492);
or UO_1 (O_1,N_9286,N_7520);
and UO_2 (O_2,N_8121,N_8655);
and UO_3 (O_3,N_9763,N_9281);
and UO_4 (O_4,N_9124,N_7674);
nor UO_5 (O_5,N_8256,N_7809);
or UO_6 (O_6,N_9835,N_9275);
nor UO_7 (O_7,N_9323,N_7949);
or UO_8 (O_8,N_8985,N_9503);
nand UO_9 (O_9,N_9787,N_9938);
or UO_10 (O_10,N_8957,N_8844);
nand UO_11 (O_11,N_8005,N_9188);
xor UO_12 (O_12,N_8541,N_8824);
nand UO_13 (O_13,N_7661,N_8275);
and UO_14 (O_14,N_8817,N_8069);
nand UO_15 (O_15,N_9197,N_7933);
nor UO_16 (O_16,N_8424,N_9999);
and UO_17 (O_17,N_9804,N_7766);
nand UO_18 (O_18,N_8015,N_9156);
nor UO_19 (O_19,N_8033,N_8970);
or UO_20 (O_20,N_7592,N_9261);
nand UO_21 (O_21,N_9382,N_8514);
and UO_22 (O_22,N_8523,N_7926);
or UO_23 (O_23,N_9596,N_8040);
or UO_24 (O_24,N_9218,N_9844);
nor UO_25 (O_25,N_8476,N_9003);
and UO_26 (O_26,N_9166,N_8140);
and UO_27 (O_27,N_8757,N_8306);
and UO_28 (O_28,N_9950,N_9768);
and UO_29 (O_29,N_8609,N_9330);
or UO_30 (O_30,N_7544,N_9241);
or UO_31 (O_31,N_9376,N_9072);
and UO_32 (O_32,N_7738,N_9774);
or UO_33 (O_33,N_7744,N_9269);
nor UO_34 (O_34,N_9054,N_9164);
nand UO_35 (O_35,N_8084,N_8616);
nand UO_36 (O_36,N_8872,N_8848);
or UO_37 (O_37,N_7792,N_7854);
or UO_38 (O_38,N_9012,N_8077);
xnor UO_39 (O_39,N_8968,N_9355);
nor UO_40 (O_40,N_9413,N_8746);
and UO_41 (O_41,N_7846,N_8645);
and UO_42 (O_42,N_7988,N_8176);
nor UO_43 (O_43,N_7627,N_8338);
nand UO_44 (O_44,N_8224,N_9408);
or UO_45 (O_45,N_9818,N_8611);
nor UO_46 (O_46,N_8950,N_7785);
and UO_47 (O_47,N_9460,N_7756);
or UO_48 (O_48,N_8528,N_8255);
or UO_49 (O_49,N_7973,N_9442);
and UO_50 (O_50,N_9163,N_9521);
or UO_51 (O_51,N_8703,N_9739);
nor UO_52 (O_52,N_9671,N_9904);
nand UO_53 (O_53,N_7908,N_9992);
nor UO_54 (O_54,N_8557,N_8928);
and UO_55 (O_55,N_8829,N_9077);
and UO_56 (O_56,N_9029,N_7543);
nor UO_57 (O_57,N_9038,N_8912);
or UO_58 (O_58,N_9506,N_9094);
or UO_59 (O_59,N_9707,N_9445);
and UO_60 (O_60,N_9761,N_8346);
and UO_61 (O_61,N_9320,N_8761);
or UO_62 (O_62,N_8971,N_9510);
and UO_63 (O_63,N_9337,N_7565);
and UO_64 (O_64,N_7847,N_9374);
and UO_65 (O_65,N_9562,N_8204);
nor UO_66 (O_66,N_8249,N_8152);
and UO_67 (O_67,N_9549,N_8963);
or UO_68 (O_68,N_8258,N_7745);
nor UO_69 (O_69,N_8764,N_7542);
nor UO_70 (O_70,N_9430,N_8840);
or UO_71 (O_71,N_9595,N_7778);
and UO_72 (O_72,N_8406,N_8931);
nand UO_73 (O_73,N_8842,N_7811);
nor UO_74 (O_74,N_7964,N_9890);
or UO_75 (O_75,N_8362,N_9883);
and UO_76 (O_76,N_9783,N_7887);
and UO_77 (O_77,N_8075,N_8486);
or UO_78 (O_78,N_9173,N_9368);
or UO_79 (O_79,N_8187,N_8414);
and UO_80 (O_80,N_8952,N_8702);
and UO_81 (O_81,N_8421,N_8850);
xor UO_82 (O_82,N_7659,N_8477);
nor UO_83 (O_83,N_8560,N_9842);
or UO_84 (O_84,N_8567,N_9016);
or UO_85 (O_85,N_9296,N_8737);
xor UO_86 (O_86,N_9934,N_9378);
nor UO_87 (O_87,N_8522,N_9803);
nor UO_88 (O_88,N_7883,N_8007);
nor UO_89 (O_89,N_9878,N_8061);
nand UO_90 (O_90,N_8464,N_8626);
and UO_91 (O_91,N_7660,N_8876);
nand UO_92 (O_92,N_8624,N_9869);
nor UO_93 (O_93,N_7708,N_8649);
nand UO_94 (O_94,N_9654,N_8054);
nand UO_95 (O_95,N_9105,N_9597);
nor UO_96 (O_96,N_8489,N_9843);
and UO_97 (O_97,N_9381,N_9748);
or UO_98 (O_98,N_9479,N_8169);
nand UO_99 (O_99,N_9634,N_7812);
nor UO_100 (O_100,N_7976,N_9556);
nor UO_101 (O_101,N_9558,N_8496);
nor UO_102 (O_102,N_9082,N_9910);
nor UO_103 (O_103,N_7572,N_9840);
nand UO_104 (O_104,N_7995,N_8181);
and UO_105 (O_105,N_9980,N_8045);
nand UO_106 (O_106,N_8094,N_9954);
nor UO_107 (O_107,N_8303,N_9245);
or UO_108 (O_108,N_8559,N_9712);
nor UO_109 (O_109,N_8922,N_8293);
and UO_110 (O_110,N_8881,N_9951);
and UO_111 (O_111,N_8854,N_8975);
or UO_112 (O_112,N_7678,N_9021);
and UO_113 (O_113,N_8715,N_7965);
or UO_114 (O_114,N_9185,N_7638);
nor UO_115 (O_115,N_9387,N_8288);
nor UO_116 (O_116,N_8240,N_8895);
or UO_117 (O_117,N_8283,N_8235);
nor UO_118 (O_118,N_8276,N_8847);
and UO_119 (O_119,N_9342,N_9443);
nand UO_120 (O_120,N_9974,N_8602);
nand UO_121 (O_121,N_7611,N_8022);
nor UO_122 (O_122,N_8372,N_9489);
or UO_123 (O_123,N_9401,N_8843);
or UO_124 (O_124,N_9664,N_9554);
or UO_125 (O_125,N_9970,N_9274);
xor UO_126 (O_126,N_8774,N_9502);
or UO_127 (O_127,N_9723,N_8704);
xor UO_128 (O_128,N_9577,N_8127);
or UO_129 (O_129,N_8991,N_7959);
nand UO_130 (O_130,N_8631,N_9217);
and UO_131 (O_131,N_9514,N_9935);
or UO_132 (O_132,N_9621,N_8646);
nand UO_133 (O_133,N_8753,N_7914);
nor UO_134 (O_134,N_7508,N_8793);
or UO_135 (O_135,N_7907,N_8336);
nand UO_136 (O_136,N_7866,N_8961);
and UO_137 (O_137,N_9372,N_8735);
nand UO_138 (O_138,N_7863,N_7799);
nor UO_139 (O_139,N_9110,N_9733);
nand UO_140 (O_140,N_8225,N_9973);
and UO_141 (O_141,N_8013,N_8179);
and UO_142 (O_142,N_7862,N_7993);
and UO_143 (O_143,N_8683,N_7786);
xnor UO_144 (O_144,N_8729,N_9256);
nand UO_145 (O_145,N_9717,N_9540);
and UO_146 (O_146,N_9919,N_8815);
nor UO_147 (O_147,N_8691,N_9699);
or UO_148 (O_148,N_8593,N_8837);
nor UO_149 (O_149,N_7900,N_9501);
nor UO_150 (O_150,N_8906,N_9161);
nor UO_151 (O_151,N_9244,N_8266);
or UO_152 (O_152,N_9734,N_9548);
nand UO_153 (O_153,N_9066,N_8792);
nand UO_154 (O_154,N_8590,N_9364);
xor UO_155 (O_155,N_8380,N_9670);
and UO_156 (O_156,N_8877,N_9478);
nor UO_157 (O_157,N_9452,N_9302);
nor UO_158 (O_158,N_9627,N_9174);
or UO_159 (O_159,N_9068,N_9799);
nor UO_160 (O_160,N_8413,N_8647);
and UO_161 (O_161,N_8600,N_7823);
and UO_162 (O_162,N_9569,N_8025);
and UO_163 (O_163,N_7950,N_8196);
or UO_164 (O_164,N_7712,N_8816);
xor UO_165 (O_165,N_8940,N_8603);
nand UO_166 (O_166,N_8891,N_8699);
and UO_167 (O_167,N_7967,N_8500);
nor UO_168 (O_168,N_7984,N_9658);
or UO_169 (O_169,N_7918,N_8893);
nand UO_170 (O_170,N_8767,N_7579);
and UO_171 (O_171,N_9095,N_8946);
or UO_172 (O_172,N_9139,N_9019);
nor UO_173 (O_173,N_7833,N_8763);
nand UO_174 (O_174,N_8955,N_8493);
or UO_175 (O_175,N_7956,N_8031);
nand UO_176 (O_176,N_9130,N_8599);
nand UO_177 (O_177,N_8951,N_9921);
nor UO_178 (O_178,N_9945,N_8897);
nor UO_179 (O_179,N_7511,N_8163);
or UO_180 (O_180,N_8430,N_9705);
or UO_181 (O_181,N_9099,N_8066);
or UO_182 (O_182,N_8065,N_8941);
nor UO_183 (O_183,N_9856,N_9065);
and UO_184 (O_184,N_7616,N_8860);
nor UO_185 (O_185,N_8526,N_8542);
and UO_186 (O_186,N_9039,N_8727);
or UO_187 (O_187,N_8589,N_8419);
or UO_188 (O_188,N_9192,N_7527);
nor UO_189 (O_189,N_8131,N_8597);
and UO_190 (O_190,N_8156,N_8976);
nor UO_191 (O_191,N_8294,N_8823);
nand UO_192 (O_192,N_8502,N_8900);
or UO_193 (O_193,N_9398,N_8123);
and UO_194 (O_194,N_9092,N_9399);
and UO_195 (O_195,N_9905,N_9583);
and UO_196 (O_196,N_8021,N_9624);
nand UO_197 (O_197,N_9885,N_7763);
nor UO_198 (O_198,N_8518,N_7741);
or UO_199 (O_199,N_8902,N_8911);
nor UO_200 (O_200,N_9559,N_8819);
nand UO_201 (O_201,N_9874,N_7706);
or UO_202 (O_202,N_9643,N_9700);
and UO_203 (O_203,N_9948,N_8651);
nand UO_204 (O_204,N_8714,N_7780);
or UO_205 (O_205,N_9766,N_9880);
and UO_206 (O_206,N_9071,N_9147);
and UO_207 (O_207,N_7961,N_8549);
and UO_208 (O_208,N_7551,N_7979);
nor UO_209 (O_209,N_8278,N_9291);
nor UO_210 (O_210,N_8863,N_8676);
or UO_211 (O_211,N_8873,N_7768);
and UO_212 (O_212,N_9609,N_8207);
nor UO_213 (O_213,N_7997,N_9606);
or UO_214 (O_214,N_8724,N_9416);
nand UO_215 (O_215,N_9715,N_8265);
nand UO_216 (O_216,N_8707,N_8828);
nand UO_217 (O_217,N_9441,N_8908);
nand UO_218 (O_218,N_8554,N_7895);
and UO_219 (O_219,N_9882,N_9417);
nor UO_220 (O_220,N_8544,N_7526);
nand UO_221 (O_221,N_9133,N_9747);
nand UO_222 (O_222,N_8312,N_8708);
nor UO_223 (O_223,N_8109,N_9340);
or UO_224 (O_224,N_8478,N_9287);
or UO_225 (O_225,N_7723,N_9555);
or UO_226 (O_226,N_8359,N_9805);
and UO_227 (O_227,N_8324,N_7770);
and UO_228 (O_228,N_9622,N_7636);
and UO_229 (O_229,N_9070,N_9119);
nor UO_230 (O_230,N_7943,N_8286);
or UO_231 (O_231,N_7981,N_7603);
and UO_232 (O_232,N_9819,N_8450);
or UO_233 (O_233,N_7919,N_7937);
and UO_234 (O_234,N_8495,N_9711);
nand UO_235 (O_235,N_8068,N_8411);
nand UO_236 (O_236,N_7673,N_8247);
nand UO_237 (O_237,N_9650,N_8635);
and UO_238 (O_238,N_8861,N_8457);
or UO_239 (O_239,N_9385,N_8375);
xnor UO_240 (O_240,N_8453,N_9465);
or UO_241 (O_241,N_7597,N_9531);
nor UO_242 (O_242,N_9030,N_8423);
and UO_243 (O_243,N_8841,N_9893);
or UO_244 (O_244,N_9745,N_8042);
or UO_245 (O_245,N_7690,N_8012);
or UO_246 (O_246,N_8331,N_8371);
and UO_247 (O_247,N_9022,N_7662);
nand UO_248 (O_248,N_8182,N_7632);
nor UO_249 (O_249,N_9204,N_9299);
nor UO_250 (O_250,N_7676,N_9267);
nand UO_251 (O_251,N_9630,N_9638);
or UO_252 (O_252,N_7618,N_9311);
nor UO_253 (O_253,N_9131,N_7670);
nand UO_254 (O_254,N_9963,N_9779);
and UO_255 (O_255,N_7873,N_9966);
nor UO_256 (O_256,N_8487,N_9719);
or UO_257 (O_257,N_8171,N_7549);
and UO_258 (O_258,N_9911,N_9474);
or UO_259 (O_259,N_9500,N_7582);
or UO_260 (O_260,N_8571,N_9590);
or UO_261 (O_261,N_7535,N_8525);
nand UO_262 (O_262,N_9272,N_9143);
nor UO_263 (O_263,N_9572,N_8009);
and UO_264 (O_264,N_9931,N_9611);
or UO_265 (O_265,N_8512,N_9150);
or UO_266 (O_266,N_8710,N_9743);
or UO_267 (O_267,N_9265,N_7695);
nand UO_268 (O_268,N_9876,N_9626);
nor UO_269 (O_269,N_8806,N_7782);
nor UO_270 (O_270,N_8245,N_9455);
nor UO_271 (O_271,N_9231,N_8122);
nand UO_272 (O_272,N_9181,N_7672);
nor UO_273 (O_273,N_9551,N_9873);
and UO_274 (O_274,N_7947,N_9369);
or UO_275 (O_275,N_8982,N_9657);
or UO_276 (O_276,N_8079,N_9917);
nand UO_277 (O_277,N_9675,N_8128);
or UO_278 (O_278,N_9132,N_8041);
nand UO_279 (O_279,N_9426,N_9560);
nand UO_280 (O_280,N_7539,N_8565);
nand UO_281 (O_281,N_9239,N_9854);
nor UO_282 (O_282,N_7901,N_9446);
nor UO_283 (O_283,N_9209,N_8277);
nor UO_284 (O_284,N_8638,N_8096);
nor UO_285 (O_285,N_9160,N_7510);
and UO_286 (O_286,N_8801,N_7894);
or UO_287 (O_287,N_8345,N_8488);
nand UO_288 (O_288,N_8504,N_8713);
nand UO_289 (O_289,N_9008,N_9867);
nand UO_290 (O_290,N_9729,N_8799);
and UO_291 (O_291,N_7939,N_8956);
nor UO_292 (O_292,N_9464,N_8973);
nor UO_293 (O_293,N_8378,N_8264);
and UO_294 (O_294,N_8779,N_8505);
nand UO_295 (O_295,N_8775,N_9914);
and UO_296 (O_296,N_8995,N_7932);
or UO_297 (O_297,N_9920,N_8773);
or UO_298 (O_298,N_7634,N_9737);
or UO_299 (O_299,N_7668,N_8325);
and UO_300 (O_300,N_8916,N_7850);
and UO_301 (O_301,N_9149,N_9794);
nor UO_302 (O_302,N_9993,N_9069);
and UO_303 (O_303,N_9480,N_7599);
or UO_304 (O_304,N_7775,N_9254);
and UO_305 (O_305,N_9491,N_9995);
nand UO_306 (O_306,N_9316,N_8846);
nand UO_307 (O_307,N_9352,N_9112);
xor UO_308 (O_308,N_9073,N_8370);
nor UO_309 (O_309,N_9676,N_9109);
and UO_310 (O_310,N_7604,N_7516);
and UO_311 (O_311,N_9341,N_9258);
or UO_312 (O_312,N_8728,N_7675);
nor UO_313 (O_313,N_7881,N_7601);
nor UO_314 (O_314,N_8297,N_9248);
and UO_315 (O_315,N_8272,N_7892);
nor UO_316 (O_316,N_9986,N_7643);
or UO_317 (O_317,N_9391,N_8326);
or UO_318 (O_318,N_9079,N_7821);
and UO_319 (O_319,N_7613,N_9425);
or UO_320 (O_320,N_8481,N_9567);
and UO_321 (O_321,N_8016,N_9709);
nand UO_322 (O_322,N_8527,N_9894);
nor UO_323 (O_323,N_9250,N_9326);
nor UO_324 (O_324,N_8408,N_9651);
nand UO_325 (O_325,N_9866,N_8654);
or UO_326 (O_326,N_7889,N_7925);
and UO_327 (O_327,N_9653,N_8510);
or UO_328 (O_328,N_8190,N_9824);
nand UO_329 (O_329,N_8177,N_9755);
and UO_330 (O_330,N_8513,N_8390);
or UO_331 (O_331,N_8731,N_7897);
or UO_332 (O_332,N_8339,N_9394);
or UO_333 (O_333,N_7752,N_9405);
or UO_334 (O_334,N_8055,N_8234);
nor UO_335 (O_335,N_8778,N_8323);
or UO_336 (O_336,N_7834,N_7577);
nand UO_337 (O_337,N_7586,N_8664);
and UO_338 (O_338,N_9001,N_8583);
nand UO_339 (O_339,N_9075,N_7912);
nor UO_340 (O_340,N_8756,N_7842);
or UO_341 (O_341,N_7711,N_9578);
nor UO_342 (O_342,N_8352,N_7583);
and UO_343 (O_343,N_9206,N_8959);
and UO_344 (O_344,N_8804,N_7621);
or UO_345 (O_345,N_7623,N_9359);
and UO_346 (O_346,N_8458,N_9081);
or UO_347 (O_347,N_8680,N_8434);
xor UO_348 (O_348,N_8930,N_8194);
and UO_349 (O_349,N_7924,N_9182);
or UO_350 (O_350,N_9319,N_9698);
or UO_351 (O_351,N_8029,N_9850);
and UO_352 (O_352,N_8316,N_8648);
nand UO_353 (O_353,N_7808,N_7774);
nor UO_354 (O_354,N_8428,N_8330);
nor UO_355 (O_355,N_8839,N_9176);
nor UO_356 (O_356,N_7653,N_9710);
nor UO_357 (O_357,N_8448,N_8994);
or UO_358 (O_358,N_8690,N_8723);
and UO_359 (O_359,N_9023,N_8174);
or UO_360 (O_360,N_7578,N_9177);
nor UO_361 (O_361,N_7920,N_7825);
or UO_362 (O_362,N_8112,N_9695);
and UO_363 (O_363,N_9448,N_9047);
xor UO_364 (O_364,N_9198,N_8962);
and UO_365 (O_365,N_7739,N_9046);
nor UO_366 (O_366,N_9607,N_8834);
and UO_367 (O_367,N_9541,N_9601);
or UO_368 (O_368,N_7714,N_9224);
nand UO_369 (O_369,N_8948,N_8533);
nand UO_370 (O_370,N_9584,N_9329);
nand UO_371 (O_371,N_8856,N_7888);
or UO_372 (O_372,N_9550,N_8536);
or UO_373 (O_373,N_7595,N_7628);
and UO_374 (O_374,N_8657,N_8093);
nor UO_375 (O_375,N_9453,N_9871);
nor UO_376 (O_376,N_7861,N_9570);
nand UO_377 (O_377,N_8894,N_8335);
and UO_378 (O_378,N_7787,N_8321);
and UO_379 (O_379,N_9884,N_8028);
nand UO_380 (O_380,N_8550,N_8832);
nor UO_381 (O_381,N_8261,N_9477);
and UO_382 (O_382,N_9058,N_9773);
and UO_383 (O_383,N_8712,N_9051);
nor UO_384 (O_384,N_9196,N_9539);
or UO_385 (O_385,N_9930,N_8284);
or UO_386 (O_386,N_7879,N_9263);
and UO_387 (O_387,N_7591,N_8064);
nand UO_388 (O_388,N_8984,N_9529);
and UO_389 (O_389,N_8791,N_7721);
nor UO_390 (O_390,N_9259,N_8665);
nor UO_391 (O_391,N_9222,N_8102);
nor UO_392 (O_392,N_9586,N_9350);
nor UO_393 (O_393,N_9832,N_9214);
nor UO_394 (O_394,N_8289,N_7767);
nor UO_395 (O_395,N_9137,N_9598);
nand UO_396 (O_396,N_7802,N_8446);
and UO_397 (O_397,N_9947,N_9436);
and UO_398 (O_398,N_9831,N_9406);
or UO_399 (O_399,N_8780,N_8569);
nand UO_400 (O_400,N_9348,N_8092);
nor UO_401 (O_401,N_7941,N_9235);
nand UO_402 (O_402,N_7598,N_8909);
or UO_403 (O_403,N_9328,N_8798);
and UO_404 (O_404,N_9288,N_8422);
and UO_405 (O_405,N_7975,N_9178);
or UO_406 (O_406,N_9701,N_8106);
and UO_407 (O_407,N_7664,N_7588);
nand UO_408 (O_408,N_7585,N_9210);
or UO_409 (O_409,N_9015,N_8784);
or UO_410 (O_410,N_9795,N_9785);
nor UO_411 (O_411,N_8178,N_9536);
nand UO_412 (O_412,N_9716,N_8257);
and UO_413 (O_413,N_7777,N_9419);
nand UO_414 (O_414,N_8287,N_9498);
and UO_415 (O_415,N_8067,N_8564);
nor UO_416 (O_416,N_7729,N_7563);
or UO_417 (O_417,N_8251,N_9037);
or UO_418 (O_418,N_8578,N_9321);
nor UO_419 (O_419,N_7971,N_8271);
or UO_420 (O_420,N_9546,N_8866);
nor UO_421 (O_421,N_8148,N_7703);
and UO_422 (O_422,N_8442,N_8643);
or UO_423 (O_423,N_8814,N_8134);
nor UO_424 (O_424,N_9410,N_8974);
nand UO_425 (O_425,N_7783,N_8919);
nand UO_426 (O_426,N_9014,N_9042);
or UO_427 (O_427,N_9414,N_8686);
and UO_428 (O_428,N_7798,N_9511);
or UO_429 (O_429,N_9765,N_9706);
or UO_430 (O_430,N_9184,N_7719);
or UO_431 (O_431,N_7574,N_9730);
and UO_432 (O_432,N_9524,N_8351);
nand UO_433 (O_433,N_9264,N_9450);
and UO_434 (O_434,N_8006,N_9989);
nand UO_435 (O_435,N_8246,N_7764);
or UO_436 (O_436,N_9409,N_9565);
or UO_437 (O_437,N_9845,N_8089);
nand UO_438 (O_438,N_9772,N_8818);
nor UO_439 (O_439,N_8270,N_9988);
or UO_440 (O_440,N_9020,N_8787);
and UO_441 (O_441,N_9395,N_9249);
or UO_442 (O_442,N_8935,N_8465);
nand UO_443 (O_443,N_8738,N_7612);
and UO_444 (O_444,N_9220,N_9673);
or UO_445 (O_445,N_8101,N_8307);
nand UO_446 (O_446,N_8805,N_9821);
nand UO_447 (O_447,N_7515,N_9924);
nor UO_448 (O_448,N_9468,N_9096);
or UO_449 (O_449,N_9226,N_8302);
nand UO_450 (O_450,N_8074,N_9396);
nor UO_451 (O_451,N_8548,N_7718);
xor UO_452 (O_452,N_9542,N_8228);
nand UO_453 (O_453,N_8168,N_9308);
nor UO_454 (O_454,N_8802,N_8992);
and UO_455 (O_455,N_9152,N_9044);
and UO_456 (O_456,N_8011,N_9505);
nor UO_457 (O_457,N_8620,N_9614);
nor UO_458 (O_458,N_8770,N_9537);
nor UO_459 (O_459,N_8198,N_9052);
or UO_460 (O_460,N_8851,N_8725);
and UO_461 (O_461,N_7843,N_9338);
and UO_462 (O_462,N_8745,N_9767);
nand UO_463 (O_463,N_8087,N_8340);
nand UO_464 (O_464,N_9041,N_9530);
or UO_465 (O_465,N_9113,N_9581);
nand UO_466 (O_466,N_9106,N_8923);
or UO_467 (O_467,N_7795,N_7500);
nand UO_468 (O_468,N_9668,N_8594);
and UO_469 (O_469,N_9903,N_8242);
nand UO_470 (O_470,N_9366,N_8639);
nor UO_471 (O_471,N_8003,N_9162);
or UO_472 (O_472,N_7594,N_8592);
nor UO_473 (O_473,N_7755,N_9897);
or UO_474 (O_474,N_9900,N_8534);
and UO_475 (O_475,N_9786,N_8389);
nor UO_476 (O_476,N_7877,N_8322);
and UO_477 (O_477,N_7518,N_8173);
nor UO_478 (O_478,N_8768,N_9255);
and UO_479 (O_479,N_7702,N_8572);
or UO_480 (O_480,N_7528,N_7838);
or UO_481 (O_481,N_7960,N_8200);
or UO_482 (O_482,N_9433,N_9290);
nand UO_483 (O_483,N_8263,N_8996);
or UO_484 (O_484,N_9758,N_9508);
nor UO_485 (O_485,N_7832,N_7637);
nor UO_486 (O_486,N_9512,N_7987);
or UO_487 (O_487,N_7750,N_8693);
nor UO_488 (O_488,N_9440,N_9193);
nand UO_489 (O_489,N_7870,N_8561);
and UO_490 (O_490,N_8803,N_8095);
nand UO_491 (O_491,N_8468,N_9543);
or UO_492 (O_492,N_7751,N_8315);
or UO_493 (O_493,N_9488,N_9813);
nand UO_494 (O_494,N_9762,N_9062);
nor UO_495 (O_495,N_7633,N_8501);
or UO_496 (O_496,N_7909,N_7966);
nand UO_497 (O_497,N_9862,N_7816);
nand UO_498 (O_498,N_7587,N_7771);
and UO_499 (O_499,N_9295,N_9683);
nand UO_500 (O_500,N_9397,N_8865);
nand UO_501 (O_501,N_8333,N_7710);
or UO_502 (O_502,N_7720,N_9778);
and UO_503 (O_503,N_9659,N_9728);
nand UO_504 (O_504,N_7608,N_8681);
or UO_505 (O_505,N_9306,N_8138);
nand UO_506 (O_506,N_9889,N_9981);
nor UO_507 (O_507,N_7757,N_8073);
nand UO_508 (O_508,N_9025,N_7635);
nand UO_509 (O_509,N_9088,N_8469);
or UO_510 (O_510,N_7725,N_9183);
nor UO_511 (O_511,N_8099,N_9371);
nor UO_512 (O_512,N_9688,N_7733);
and UO_513 (O_513,N_8749,N_9278);
nor UO_514 (O_514,N_8701,N_8595);
or UO_515 (O_515,N_8998,N_8880);
nor UO_516 (O_516,N_8416,N_8107);
nor UO_517 (O_517,N_8517,N_8835);
or UO_518 (O_518,N_9545,N_9045);
nor UO_519 (O_519,N_9823,N_7835);
or UO_520 (O_520,N_7682,N_8314);
and UO_521 (O_521,N_7698,N_9532);
and UO_522 (O_522,N_9916,N_7805);
nand UO_523 (O_523,N_9312,N_9741);
or UO_524 (O_524,N_8479,N_8588);
and UO_525 (O_525,N_8260,N_9852);
or UO_526 (O_526,N_8212,N_8553);
and UO_527 (O_527,N_9941,N_9444);
and UO_528 (O_528,N_7998,N_7970);
nand UO_529 (O_529,N_9357,N_8766);
and UO_530 (O_530,N_8132,N_9400);
nor UO_531 (O_531,N_9246,N_8933);
or UO_532 (O_532,N_9179,N_9034);
nor UO_533 (O_533,N_9744,N_7974);
or UO_534 (O_534,N_8607,N_8360);
and UO_535 (O_535,N_9157,N_8080);
nand UO_536 (O_536,N_8395,N_8387);
nand UO_537 (O_537,N_9365,N_9853);
nand UO_538 (O_538,N_8601,N_9434);
nand UO_539 (O_539,N_9937,N_8215);
nand UO_540 (O_540,N_7781,N_9236);
and UO_541 (O_541,N_9200,N_8043);
nand UO_542 (O_542,N_9327,N_8402);
and UO_543 (O_543,N_9703,N_9064);
nand UO_544 (O_544,N_9775,N_9470);
or UO_545 (O_545,N_8216,N_9825);
or UO_546 (O_546,N_9589,N_7958);
and UO_547 (O_547,N_9153,N_8202);
or UO_548 (O_548,N_8184,N_8547);
nand UO_549 (O_549,N_8205,N_9571);
nor UO_550 (O_550,N_8896,N_8890);
and UO_551 (O_551,N_8452,N_9807);
or UO_552 (O_552,N_7867,N_9449);
or UO_553 (O_553,N_9764,N_8660);
and UO_554 (O_554,N_9507,N_9361);
and UO_555 (O_555,N_9788,N_9170);
nor UO_556 (O_556,N_9965,N_9107);
or UO_557 (O_557,N_7696,N_8162);
nand UO_558 (O_558,N_9238,N_7837);
and UO_559 (O_559,N_8199,N_8598);
nand UO_560 (O_560,N_7650,N_7512);
and UO_561 (O_561,N_9946,N_9393);
or UO_562 (O_562,N_9770,N_9144);
and UO_563 (O_563,N_9146,N_8466);
or UO_564 (O_564,N_9771,N_8243);
nor UO_565 (O_565,N_8296,N_9944);
and UO_566 (O_566,N_9742,N_8776);
or UO_567 (O_567,N_7651,N_8618);
or UO_568 (O_568,N_9485,N_9661);
nor UO_569 (O_569,N_8081,N_7576);
nor UO_570 (O_570,N_9279,N_7533);
or UO_571 (O_571,N_9509,N_9942);
nor UO_572 (O_572,N_7685,N_8480);
or UO_573 (O_573,N_9985,N_9936);
and UO_574 (O_574,N_8892,N_7957);
and UO_575 (O_575,N_8915,N_8250);
nor UO_576 (O_576,N_9836,N_7831);
and UO_577 (O_577,N_9702,N_9816);
nor UO_578 (O_578,N_9674,N_8644);
or UO_579 (O_579,N_9459,N_7828);
nor UO_580 (O_580,N_8197,N_9922);
or UO_581 (O_581,N_7826,N_7614);
and UO_582 (O_582,N_9526,N_9677);
nand UO_583 (O_583,N_9411,N_8105);
nor UO_584 (O_584,N_7550,N_7640);
and UO_585 (O_585,N_8530,N_7540);
nand UO_586 (O_586,N_9967,N_9221);
nand UO_587 (O_587,N_9240,N_8467);
and UO_588 (O_588,N_8661,N_7911);
nor UO_589 (O_589,N_8490,N_8608);
or UO_590 (O_590,N_8188,N_9685);
and UO_591 (O_591,N_8788,N_7546);
nor UO_592 (O_592,N_7902,N_9848);
nand UO_593 (O_593,N_8070,N_7532);
nor UO_594 (O_594,N_9428,N_8936);
and UO_595 (O_595,N_9696,N_8899);
nor UO_596 (O_596,N_7564,N_8393);
or UO_597 (O_597,N_9839,N_9252);
nand UO_598 (O_598,N_9203,N_7642);
and UO_599 (O_599,N_9093,N_8456);
nor UO_600 (O_600,N_8300,N_7807);
and UO_601 (O_601,N_9718,N_7715);
or UO_602 (O_602,N_7830,N_9587);
and UO_603 (O_603,N_9633,N_8157);
and UO_604 (O_604,N_9566,N_8304);
nor UO_605 (O_605,N_8621,N_7891);
or UO_606 (O_606,N_8129,N_9298);
nor UO_607 (O_607,N_9605,N_7874);
nor UO_608 (O_608,N_8666,N_9297);
or UO_609 (O_609,N_8396,N_9289);
nor UO_610 (O_610,N_8214,N_9050);
nor UO_611 (O_611,N_8605,N_7991);
nor UO_612 (O_612,N_7938,N_9881);
nor UO_613 (O_613,N_8509,N_7502);
nand UO_614 (O_614,N_8443,N_8953);
nand UO_615 (O_615,N_8049,N_8274);
nor UO_616 (O_616,N_9083,N_8407);
nor UO_617 (O_617,N_9984,N_7688);
or UO_618 (O_618,N_8153,N_7827);
or UO_619 (O_619,N_8625,N_9864);
nor UO_620 (O_620,N_9956,N_7904);
and UO_621 (O_621,N_8241,N_8986);
or UO_622 (O_622,N_8158,N_8219);
or UO_623 (O_623,N_9090,N_7882);
nor UO_624 (O_624,N_9603,N_7927);
nand UO_625 (O_625,N_8627,N_7584);
and UO_626 (O_626,N_7989,N_7878);
and UO_627 (O_627,N_9610,N_8350);
and UO_628 (O_628,N_8273,N_7880);
nand UO_629 (O_629,N_8870,N_8679);
or UO_630 (O_630,N_8400,N_7936);
and UO_631 (O_631,N_7626,N_8034);
or UO_632 (O_632,N_8853,N_9827);
or UO_633 (O_633,N_7607,N_8142);
or UO_634 (O_634,N_9140,N_8309);
nor UO_635 (O_635,N_9828,N_7906);
nor UO_636 (O_636,N_9086,N_9447);
or UO_637 (O_637,N_7657,N_8568);
and UO_638 (O_638,N_9456,N_8248);
nand UO_639 (O_639,N_7665,N_9538);
and UO_640 (O_640,N_8821,N_8721);
nor UO_641 (O_641,N_9009,N_8417);
or UO_642 (O_642,N_8000,N_9102);
nand UO_643 (O_643,N_9122,N_9806);
nor UO_644 (O_644,N_8811,N_9789);
or UO_645 (O_645,N_7605,N_9915);
and UO_646 (O_646,N_8736,N_8642);
nor UO_647 (O_647,N_8349,N_7704);
nor UO_648 (O_648,N_7731,N_8613);
nor UO_649 (O_649,N_7513,N_8368);
nand UO_650 (O_650,N_9943,N_7713);
or UO_651 (O_651,N_9036,N_8332);
nor UO_652 (O_652,N_7829,N_9004);
and UO_653 (O_653,N_8001,N_8010);
xnor UO_654 (O_654,N_9604,N_9476);
or UO_655 (O_655,N_7884,N_7545);
and UO_656 (O_656,N_9314,N_9721);
nand UO_657 (O_657,N_9078,N_9666);
and UO_658 (O_658,N_8392,N_8855);
nand UO_659 (O_659,N_9678,N_9349);
nand UO_660 (O_660,N_8540,N_8825);
and UO_661 (O_661,N_8612,N_7994);
xor UO_662 (O_662,N_9817,N_8385);
and UO_663 (O_663,N_7724,N_9751);
or UO_664 (O_664,N_8146,N_8301);
nand UO_665 (O_665,N_9720,N_8059);
and UO_666 (O_666,N_8772,N_7820);
nand UO_667 (O_667,N_9544,N_8218);
or UO_668 (O_668,N_8135,N_8675);
nand UO_669 (O_669,N_9781,N_7876);
nor UO_670 (O_670,N_9168,N_8999);
nand UO_671 (O_671,N_9339,N_9632);
and UO_672 (O_672,N_8857,N_7554);
nor UO_673 (O_673,N_8383,N_7727);
or UO_674 (O_674,N_8754,N_8038);
or UO_675 (O_675,N_8026,N_9964);
nor UO_676 (O_676,N_9482,N_9262);
xor UO_677 (O_677,N_8524,N_8869);
xnor UO_678 (O_678,N_8849,N_9462);
and UO_679 (O_679,N_7930,N_9644);
and UO_680 (O_680,N_9169,N_7841);
nor UO_681 (O_681,N_9228,N_7915);
or UO_682 (O_682,N_8328,N_9483);
nor UO_683 (O_683,N_7951,N_9351);
and UO_684 (O_684,N_9219,N_8381);
nand UO_685 (O_685,N_8410,N_8913);
nand UO_686 (O_686,N_9648,N_8960);
and UO_687 (O_687,N_8499,N_8845);
nor UO_688 (O_688,N_8209,N_7972);
or UO_689 (O_689,N_9860,N_9123);
or UO_690 (O_690,N_7794,N_8221);
and UO_691 (O_691,N_9642,N_8658);
nor UO_692 (O_692,N_8483,N_9939);
or UO_693 (O_693,N_8440,N_8193);
nand UO_694 (O_694,N_8104,N_8934);
or UO_695 (O_695,N_8388,N_8630);
and UO_696 (O_696,N_8606,N_8475);
or UO_697 (O_697,N_9976,N_9877);
nor UO_698 (O_698,N_7615,N_9983);
and UO_699 (O_699,N_8144,N_8455);
nand UO_700 (O_700,N_9379,N_8983);
nand UO_701 (O_701,N_9516,N_8687);
and UO_702 (O_702,N_8425,N_7600);
nand UO_703 (O_703,N_9517,N_8361);
or UO_704 (O_704,N_9660,N_8903);
or UO_705 (O_705,N_9018,N_8800);
and UO_706 (O_706,N_7982,N_8027);
nor UO_707 (O_707,N_8685,N_9418);
xnor UO_708 (O_708,N_8344,N_9892);
or UO_709 (O_709,N_9332,N_7522);
and UO_710 (O_710,N_8119,N_9929);
nand UO_711 (O_711,N_8826,N_8917);
and UO_712 (O_712,N_9708,N_7580);
nand UO_713 (O_713,N_9849,N_7800);
nor UO_714 (O_714,N_8538,N_8223);
xnor UO_715 (O_715,N_7644,N_9802);
nor UO_716 (O_716,N_8619,N_9997);
or UO_717 (O_717,N_9334,N_7602);
or UO_718 (O_718,N_7680,N_7619);
and UO_719 (O_719,N_9487,N_9031);
and UO_720 (O_720,N_9191,N_8532);
nor UO_721 (O_721,N_9757,N_8684);
and UO_722 (O_722,N_9114,N_9855);
and UO_723 (O_723,N_8398,N_8290);
and UO_724 (O_724,N_7791,N_7728);
xor UO_725 (O_725,N_9344,N_9953);
and UO_726 (O_726,N_7609,N_9694);
or UO_727 (O_727,N_7856,N_8432);
nand UO_728 (O_728,N_9791,N_9955);
nand UO_729 (O_729,N_8978,N_9284);
nand UO_730 (O_730,N_9002,N_8310);
xnor UO_731 (O_731,N_8110,N_8515);
or UO_732 (O_732,N_8910,N_9463);
nand UO_733 (O_733,N_9769,N_9208);
and UO_734 (O_734,N_9972,N_8615);
and UO_735 (O_735,N_8318,N_7885);
or UO_736 (O_736,N_8114,N_8192);
or UO_737 (O_737,N_9300,N_8208);
nor UO_738 (O_738,N_9135,N_7709);
and UO_739 (O_739,N_9722,N_8947);
nor UO_740 (O_740,N_8017,N_7742);
nand UO_741 (O_741,N_9367,N_8697);
nor UO_742 (O_742,N_9613,N_9115);
nor UO_743 (O_743,N_7722,N_7596);
or UO_744 (O_744,N_8926,N_9151);
or UO_745 (O_745,N_8743,N_9576);
and UO_746 (O_746,N_8020,N_9793);
nor UO_747 (O_747,N_7523,N_8374);
nor UO_748 (O_748,N_9525,N_8126);
nand UO_749 (O_749,N_9753,N_7990);
nand UO_750 (O_750,N_7617,N_8581);
nand UO_751 (O_751,N_8718,N_8357);
nand UO_752 (O_752,N_7684,N_9594);
nor UO_753 (O_753,N_9563,N_9407);
nor UO_754 (O_754,N_9809,N_9879);
and UO_755 (O_755,N_9043,N_9402);
and UO_756 (O_756,N_9097,N_9968);
nor UO_757 (O_757,N_9579,N_9704);
and UO_758 (O_758,N_7529,N_7624);
and UO_759 (O_759,N_8875,N_8373);
nor UO_760 (O_760,N_8008,N_8717);
and UO_761 (O_761,N_9667,N_7652);
or UO_762 (O_762,N_9714,N_9053);
or UO_763 (O_763,N_7553,N_9421);
xor UO_764 (O_764,N_9148,N_9377);
xor UO_765 (O_765,N_9912,N_9582);
xor UO_766 (O_766,N_7740,N_8752);
nand UO_767 (O_767,N_8943,N_7560);
nor UO_768 (O_768,N_8694,N_8765);
nand UO_769 (O_769,N_8604,N_9592);
nor UO_770 (O_770,N_8972,N_8348);
or UO_771 (O_771,N_9901,N_9949);
nand UO_772 (O_772,N_9969,N_9175);
or UO_773 (O_773,N_8969,N_9631);
and UO_774 (O_774,N_8211,N_8989);
nand UO_775 (O_775,N_8091,N_8267);
or UO_776 (O_776,N_7691,N_9665);
and UO_777 (O_777,N_7556,N_8124);
nor UO_778 (O_778,N_9625,N_7589);
or UO_779 (O_779,N_8556,N_7818);
nand UO_780 (O_780,N_9136,N_8019);
or UO_781 (O_781,N_9098,N_9028);
and UO_782 (O_782,N_7504,N_8742);
nor UO_783 (O_783,N_8566,N_7852);
nand UO_784 (O_784,N_9154,N_7506);
or UO_785 (O_785,N_8584,N_8734);
and UO_786 (O_786,N_8751,N_8641);
nor UO_787 (O_787,N_9356,N_9280);
or UO_788 (O_788,N_8451,N_8471);
and UO_789 (O_789,N_9846,N_9007);
and UO_790 (O_790,N_9962,N_9756);
nor UO_791 (O_791,N_9782,N_8636);
nand UO_792 (O_792,N_9437,N_8640);
nand UO_793 (O_793,N_9335,N_8698);
and UO_794 (O_794,N_8945,N_7946);
and UO_795 (O_795,N_9907,N_9116);
nand UO_796 (O_796,N_7701,N_9363);
or UO_797 (O_797,N_9089,N_8669);
and UO_798 (O_798,N_9987,N_8369);
nand UO_799 (O_799,N_9750,N_8436);
nand UO_800 (O_800,N_8186,N_9027);
nand UO_801 (O_801,N_8036,N_8964);
nor UO_802 (O_802,N_9724,N_8150);
nor UO_803 (O_803,N_7824,N_7726);
nand UO_804 (O_804,N_7694,N_8797);
nand UO_805 (O_805,N_8575,N_8253);
or UO_806 (O_806,N_8706,N_8795);
and UO_807 (O_807,N_9815,N_9347);
and UO_808 (O_808,N_9424,N_9687);
or UO_809 (O_809,N_9294,N_8720);
nor UO_810 (O_810,N_9211,N_9732);
or UO_811 (O_811,N_8577,N_9458);
nor UO_812 (O_812,N_7983,N_9243);
or UO_813 (O_813,N_8213,N_7999);
or UO_814 (O_814,N_7590,N_8460);
nor UO_815 (O_815,N_9207,N_9847);
or UO_816 (O_816,N_8794,N_9268);
nand UO_817 (O_817,N_7839,N_8653);
nor UO_818 (O_818,N_8470,N_8166);
and UO_819 (O_819,N_9373,N_7683);
nor UO_820 (O_820,N_8125,N_9467);
xor UO_821 (O_821,N_8147,N_8161);
or UO_822 (O_822,N_9909,N_8552);
or UO_823 (O_823,N_9790,N_8543);
or UO_824 (O_824,N_9834,N_9875);
nor UO_825 (O_825,N_9796,N_7575);
or UO_826 (O_826,N_9471,N_7630);
nor UO_827 (O_827,N_7648,N_9725);
or UO_828 (O_828,N_8927,N_8570);
or UO_829 (O_829,N_9223,N_9229);
nor UO_830 (O_830,N_9684,N_9412);
nand UO_831 (O_831,N_7606,N_9812);
and UO_832 (O_832,N_9513,N_7747);
nor UO_833 (O_833,N_7759,N_9232);
and UO_834 (O_834,N_8907,N_7865);
nand UO_835 (O_835,N_8591,N_7753);
and UO_836 (O_836,N_8790,N_9872);
nor UO_837 (O_837,N_9689,N_9345);
or UO_838 (O_838,N_8937,N_8886);
nor UO_839 (O_839,N_8229,N_8227);
and UO_840 (O_840,N_8462,N_7992);
and UO_841 (O_841,N_8252,N_7845);
or UO_842 (O_842,N_7622,N_9429);
xor UO_843 (O_843,N_9777,N_8337);
and UO_844 (O_844,N_9740,N_9655);
nor UO_845 (O_845,N_8507,N_9800);
or UO_846 (O_846,N_7779,N_7806);
and UO_847 (O_847,N_7663,N_8014);
nand UO_848 (O_848,N_7679,N_9599);
xor UO_849 (O_849,N_8342,N_8889);
nor UO_850 (O_850,N_8164,N_9189);
nor UO_851 (O_851,N_7559,N_8461);
nand UO_852 (O_852,N_9383,N_9959);
or UO_853 (O_853,N_8420,N_7803);
and UO_854 (O_854,N_9528,N_8537);
nand UO_855 (O_855,N_9861,N_7872);
or UO_856 (O_856,N_8586,N_7692);
nor UO_857 (O_857,N_7996,N_7913);
and UO_858 (O_858,N_9612,N_8454);
nand UO_859 (O_859,N_7509,N_8862);
and UO_860 (O_860,N_7804,N_8587);
nor UO_861 (O_861,N_9575,N_8852);
nand UO_862 (O_862,N_7658,N_7687);
nor UO_863 (O_863,N_9829,N_7858);
nand UO_864 (O_864,N_8827,N_8405);
xor UO_865 (O_865,N_7537,N_8579);
and UO_866 (O_866,N_7505,N_8921);
and UO_867 (O_867,N_8520,N_8004);
nor UO_868 (O_868,N_9049,N_9518);
nand UO_869 (O_869,N_7944,N_8474);
or UO_870 (O_870,N_9325,N_9360);
nand UO_871 (O_871,N_8183,N_7521);
or UO_872 (O_872,N_8279,N_8427);
nand UO_873 (O_873,N_9990,N_8313);
or UO_874 (O_874,N_8437,N_8663);
nor UO_875 (O_875,N_9353,N_7916);
or UO_876 (O_876,N_8088,N_7784);
nor UO_877 (O_877,N_9126,N_7686);
nand UO_878 (O_878,N_7524,N_8060);
nand UO_879 (O_879,N_8696,N_7836);
or UO_880 (O_880,N_9637,N_7928);
nor UO_881 (O_881,N_7758,N_9979);
or UO_882 (O_882,N_9087,N_8233);
and UO_883 (O_883,N_8130,N_8932);
and UO_884 (O_884,N_7954,N_7853);
nor UO_885 (O_885,N_9978,N_9271);
nand UO_886 (O_886,N_9055,N_9669);
or UO_887 (O_887,N_7761,N_9602);
and UO_888 (O_888,N_8629,N_7571);
nor UO_889 (O_889,N_7593,N_8531);
and UO_890 (O_890,N_8391,N_9736);
nor UO_891 (O_891,N_9574,N_8682);
and UO_892 (O_892,N_8771,N_9461);
or UO_893 (O_893,N_7952,N_7769);
and UO_894 (O_894,N_9121,N_8191);
or UO_895 (O_895,N_8018,N_8628);
nand UO_896 (O_896,N_9888,N_8796);
nor UO_897 (O_897,N_9040,N_9273);
or UO_898 (O_898,N_9032,N_9557);
nor UO_899 (O_899,N_8232,N_7552);
nor UO_900 (O_900,N_9282,N_8175);
or UO_901 (O_901,N_9403,N_8988);
and UO_902 (O_902,N_8170,N_8546);
nand UO_903 (O_903,N_9649,N_8473);
or UO_904 (O_904,N_9165,N_8165);
nand UO_905 (O_905,N_7980,N_8888);
nand UO_906 (O_906,N_9749,N_8329);
or UO_907 (O_907,N_9310,N_8090);
or UO_908 (O_908,N_9693,N_8057);
nand UO_909 (O_909,N_8494,N_9117);
nor UO_910 (O_910,N_9420,N_8172);
nor UO_911 (O_911,N_9552,N_9908);
and UO_912 (O_912,N_8482,N_9000);
nor UO_913 (O_913,N_8023,N_8596);
or UO_914 (O_914,N_8634,N_8149);
nor UO_915 (O_915,N_7765,N_8115);
nand UO_916 (O_916,N_9746,N_9681);
and UO_917 (O_917,N_8238,N_7736);
or UO_918 (O_918,N_8516,N_8563);
nor UO_919 (O_919,N_9158,N_8050);
nor UO_920 (O_920,N_9380,N_9629);
nand UO_921 (O_921,N_9899,N_9647);
or UO_922 (O_922,N_8677,N_8511);
and UO_923 (O_923,N_9195,N_9858);
nand UO_924 (O_924,N_8812,N_9808);
nand UO_925 (O_925,N_7531,N_9155);
nand UO_926 (O_926,N_9568,N_8435);
nand UO_927 (O_927,N_8674,N_9084);
nor UO_928 (O_928,N_8722,N_9331);
and UO_929 (O_929,N_8269,N_8048);
and UO_930 (O_930,N_8347,N_8695);
and UO_931 (O_931,N_7558,N_9841);
nor UO_932 (O_932,N_8262,N_8305);
nor UO_933 (O_933,N_9386,N_7538);
nand UO_934 (O_934,N_7962,N_8063);
or UO_935 (O_935,N_9277,N_7760);
nor UO_936 (O_936,N_7922,N_9784);
nand UO_937 (O_937,N_9215,N_9754);
nor UO_938 (O_938,N_9466,N_7569);
or UO_939 (O_939,N_9145,N_9336);
or UO_940 (O_940,N_9731,N_8944);
or UO_941 (O_941,N_9977,N_8813);
and UO_942 (O_942,N_8981,N_8334);
or UO_943 (O_943,N_9333,N_7813);
or UO_944 (O_944,N_9960,N_9190);
or UO_945 (O_945,N_9033,N_9251);
nor UO_946 (O_946,N_9830,N_8415);
nand UO_947 (O_947,N_8117,N_9063);
nor UO_948 (O_948,N_8280,N_9591);
or UO_949 (O_949,N_9451,N_8418);
nand UO_950 (O_950,N_8399,N_8762);
nand UO_951 (O_951,N_9475,N_7797);
or UO_952 (O_952,N_8426,N_8047);
nor UO_953 (O_953,N_9370,N_7905);
or UO_954 (O_954,N_9358,N_7507);
nor UO_955 (O_955,N_9438,N_7776);
nand UO_956 (O_956,N_8052,N_7953);
nand UO_957 (O_957,N_9317,N_9010);
and UO_958 (O_958,N_9134,N_9227);
and UO_959 (O_959,N_9618,N_9975);
nand UO_960 (O_960,N_9898,N_8445);
or UO_961 (O_961,N_8268,N_8113);
nor UO_962 (O_962,N_7746,N_8141);
or UO_963 (O_963,N_8298,N_7689);
or UO_964 (O_964,N_7705,N_9495);
nor UO_965 (O_965,N_9404,N_7655);
and UO_966 (O_966,N_9108,N_8394);
nand UO_967 (O_967,N_8519,N_9129);
or UO_968 (O_968,N_7849,N_8379);
or UO_969 (O_969,N_7848,N_8447);
nor UO_970 (O_970,N_9616,N_9682);
nor UO_971 (O_971,N_7893,N_7717);
nand UO_972 (O_972,N_8491,N_9225);
and UO_973 (O_973,N_9048,N_7541);
nand UO_974 (O_974,N_8071,N_9833);
and UO_975 (O_975,N_9324,N_8747);
or UO_976 (O_976,N_7666,N_8343);
nand UO_977 (O_977,N_9958,N_9535);
nand UO_978 (O_978,N_8758,N_9857);
nor UO_979 (O_979,N_9564,N_7986);
nor UO_980 (O_980,N_8990,N_9600);
or UO_981 (O_981,N_8610,N_7547);
nor UO_982 (O_982,N_8444,N_9527);
nand UO_983 (O_983,N_9423,N_9167);
nand UO_984 (O_984,N_9304,N_8887);
nor UO_985 (O_985,N_9301,N_9141);
nor UO_986 (O_986,N_9887,N_9838);
nor UO_987 (O_987,N_9473,N_8498);
nor UO_988 (O_988,N_8580,N_8189);
and UO_989 (O_989,N_7737,N_7693);
nor UO_990 (O_990,N_9390,N_7977);
and UO_991 (O_991,N_8401,N_8929);
or UO_992 (O_992,N_7871,N_8439);
or UO_993 (O_993,N_9111,N_7963);
nor UO_994 (O_994,N_9519,N_7514);
nor UO_995 (O_995,N_8429,N_7625);
nor UO_996 (O_996,N_9776,N_8898);
nor UO_997 (O_997,N_8692,N_8431);
nand UO_998 (O_998,N_8748,N_8295);
or UO_999 (O_999,N_7530,N_8097);
nand UO_1000 (O_1000,N_9076,N_7735);
nand UO_1001 (O_1001,N_8459,N_9013);
and UO_1002 (O_1002,N_9636,N_8376);
and UO_1003 (O_1003,N_9180,N_9305);
and UO_1004 (O_1004,N_9293,N_8716);
xor UO_1005 (O_1005,N_7940,N_8024);
nand UO_1006 (O_1006,N_9759,N_8650);
nand UO_1007 (O_1007,N_8281,N_8555);
or UO_1008 (O_1008,N_9142,N_9057);
or UO_1009 (O_1009,N_9247,N_9313);
and UO_1010 (O_1010,N_9932,N_9957);
and UO_1011 (O_1011,N_7567,N_8382);
and UO_1012 (O_1012,N_8226,N_9292);
and UO_1013 (O_1013,N_8143,N_8492);
or UO_1014 (O_1014,N_8086,N_8836);
and UO_1015 (O_1015,N_9260,N_9925);
or UO_1016 (O_1016,N_8667,N_7503);
or UO_1017 (O_1017,N_8901,N_9375);
nor UO_1018 (O_1018,N_8485,N_7631);
nor UO_1019 (O_1019,N_9212,N_8292);
nor UO_1020 (O_1020,N_8210,N_8133);
nor UO_1021 (O_1021,N_9792,N_7581);
or UO_1022 (O_1022,N_9902,N_9496);
nor UO_1023 (O_1023,N_8155,N_9309);
nand UO_1024 (O_1024,N_9952,N_8868);
nand UO_1025 (O_1025,N_8769,N_9645);
or UO_1026 (O_1026,N_8918,N_7548);
and UO_1027 (O_1027,N_7570,N_7730);
nand UO_1028 (O_1028,N_9918,N_7896);
or UO_1029 (O_1029,N_9253,N_7978);
nor UO_1030 (O_1030,N_9005,N_9486);
nor UO_1031 (O_1031,N_8404,N_9201);
nor UO_1032 (O_1032,N_7743,N_7762);
xnor UO_1033 (O_1033,N_9998,N_7573);
nor UO_1034 (O_1034,N_7700,N_8358);
or UO_1035 (O_1035,N_8741,N_7793);
and UO_1036 (O_1036,N_8949,N_7645);
and UO_1037 (O_1037,N_7814,N_9283);
or UO_1038 (O_1038,N_7801,N_7557);
nand UO_1039 (O_1039,N_8659,N_9056);
nand UO_1040 (O_1040,N_9814,N_9691);
nor UO_1041 (O_1041,N_9457,N_9923);
and UO_1042 (O_1042,N_8355,N_8920);
nand UO_1043 (O_1043,N_9672,N_9727);
or UO_1044 (O_1044,N_7534,N_7669);
xor UO_1045 (O_1045,N_9186,N_9801);
or UO_1046 (O_1046,N_9573,N_8672);
xor UO_1047 (O_1047,N_7641,N_8883);
nand UO_1048 (O_1048,N_8299,N_8497);
or UO_1049 (O_1049,N_9125,N_7501);
or UO_1050 (O_1050,N_8924,N_8822);
nand UO_1051 (O_1051,N_8558,N_7819);
and UO_1052 (O_1052,N_7864,N_9230);
nand UO_1053 (O_1053,N_9504,N_9100);
nor UO_1054 (O_1054,N_9006,N_7519);
nor UO_1055 (O_1055,N_9991,N_9679);
or UO_1056 (O_1056,N_8789,N_8585);
nor UO_1057 (O_1057,N_7561,N_9863);
nor UO_1058 (O_1058,N_9202,N_9522);
and UO_1059 (O_1059,N_8777,N_8366);
nand UO_1060 (O_1060,N_9494,N_8403);
and UO_1061 (O_1061,N_7620,N_9628);
and UO_1062 (O_1062,N_9896,N_8154);
nor UO_1063 (O_1063,N_9270,N_8882);
or UO_1064 (O_1064,N_8904,N_9895);
nand UO_1065 (O_1065,N_8237,N_8623);
or UO_1066 (O_1066,N_9118,N_8433);
or UO_1067 (O_1067,N_8539,N_9663);
and UO_1068 (O_1068,N_9454,N_9389);
nor UO_1069 (O_1069,N_8449,N_9686);
nor UO_1070 (O_1070,N_9138,N_8062);
nand UO_1071 (O_1071,N_8954,N_8167);
and UO_1072 (O_1072,N_8838,N_9523);
and UO_1073 (O_1073,N_8574,N_9837);
and UO_1074 (O_1074,N_7646,N_8759);
xor UO_1075 (O_1075,N_8700,N_8750);
nor UO_1076 (O_1076,N_9580,N_9484);
nand UO_1077 (O_1077,N_7629,N_8965);
nor UO_1078 (O_1078,N_9171,N_9128);
and UO_1079 (O_1079,N_9307,N_8807);
nand UO_1080 (O_1080,N_9797,N_9891);
and UO_1081 (O_1081,N_9617,N_7517);
and UO_1082 (O_1082,N_8632,N_8858);
and UO_1083 (O_1083,N_8809,N_8688);
nand UO_1084 (O_1084,N_8206,N_8409);
nand UO_1085 (O_1085,N_8116,N_8874);
and UO_1086 (O_1086,N_8726,N_9472);
nand UO_1087 (O_1087,N_8076,N_8878);
nor UO_1088 (O_1088,N_8885,N_8291);
or UO_1089 (O_1089,N_9104,N_7772);
or UO_1090 (O_1090,N_8082,N_8002);
and UO_1091 (O_1091,N_9641,N_7647);
or UO_1092 (O_1092,N_8652,N_8662);
nor UO_1093 (O_1093,N_9652,N_8353);
or UO_1094 (O_1094,N_7748,N_7942);
or UO_1095 (O_1095,N_8056,N_8217);
nand UO_1096 (O_1096,N_9561,N_8032);
nand UO_1097 (O_1097,N_8535,N_9276);
and UO_1098 (O_1098,N_9469,N_9933);
nor UO_1099 (O_1099,N_9427,N_7860);
nand UO_1100 (O_1100,N_9415,N_7859);
nand UO_1101 (O_1101,N_8035,N_8195);
or UO_1102 (O_1102,N_9822,N_8864);
nor UO_1103 (O_1103,N_9620,N_7840);
or UO_1104 (O_1104,N_9194,N_9384);
nor UO_1105 (O_1105,N_8386,N_8656);
nand UO_1106 (O_1106,N_9322,N_7934);
and UO_1107 (O_1107,N_7869,N_9303);
nor UO_1108 (O_1108,N_9553,N_9913);
nor UO_1109 (O_1109,N_8103,N_7851);
nor UO_1110 (O_1110,N_8078,N_9865);
nand UO_1111 (O_1111,N_7929,N_8254);
and UO_1112 (O_1112,N_8397,N_9927);
and UO_1113 (O_1113,N_7875,N_7610);
or UO_1114 (O_1114,N_8058,N_9060);
or UO_1115 (O_1115,N_8958,N_9615);
and UO_1116 (O_1116,N_8966,N_8222);
nand UO_1117 (O_1117,N_8236,N_7815);
or UO_1118 (O_1118,N_9481,N_9926);
nand UO_1119 (O_1119,N_8051,N_9690);
or UO_1120 (O_1120,N_8508,N_9392);
and UO_1121 (O_1121,N_8503,N_7789);
xnor UO_1122 (O_1122,N_7525,N_9646);
or UO_1123 (O_1123,N_8709,N_7749);
or UO_1124 (O_1124,N_7699,N_9593);
or UO_1125 (O_1125,N_8705,N_7857);
or UO_1126 (O_1126,N_8377,N_7868);
nor UO_1127 (O_1127,N_8046,N_8879);
nor UO_1128 (O_1128,N_8438,N_7923);
nor UO_1129 (O_1129,N_7890,N_7844);
nand UO_1130 (O_1130,N_8185,N_8884);
nand UO_1131 (O_1131,N_7948,N_8942);
nand UO_1132 (O_1132,N_9635,N_9886);
nand UO_1133 (O_1133,N_9266,N_9091);
or UO_1134 (O_1134,N_8098,N_7562);
and UO_1135 (O_1135,N_7985,N_8151);
or UO_1136 (O_1136,N_9026,N_8820);
nand UO_1137 (O_1137,N_8484,N_9692);
and UO_1138 (O_1138,N_9074,N_7790);
nand UO_1139 (O_1139,N_9780,N_9085);
nand UO_1140 (O_1140,N_9237,N_7716);
xnor UO_1141 (O_1141,N_9101,N_7649);
and UO_1142 (O_1142,N_9172,N_9608);
nand UO_1143 (O_1143,N_8072,N_8711);
and UO_1144 (O_1144,N_8786,N_8867);
nor UO_1145 (O_1145,N_9059,N_7671);
and UO_1146 (O_1146,N_8545,N_9547);
and UO_1147 (O_1147,N_8085,N_8039);
nor UO_1148 (O_1148,N_9798,N_9493);
or UO_1149 (O_1149,N_9639,N_8744);
and UO_1150 (O_1150,N_8914,N_9928);
or UO_1151 (O_1151,N_9080,N_8120);
and UO_1152 (O_1152,N_7555,N_8311);
nor UO_1153 (O_1153,N_7945,N_8668);
and UO_1154 (O_1154,N_8967,N_8993);
nor UO_1155 (O_1155,N_7677,N_8979);
nor UO_1156 (O_1156,N_9738,N_9011);
or UO_1157 (O_1157,N_8833,N_8363);
nand UO_1158 (O_1158,N_9242,N_7566);
nand UO_1159 (O_1159,N_9017,N_9315);
or UO_1160 (O_1160,N_9680,N_8506);
and UO_1161 (O_1161,N_9127,N_8320);
nor UO_1162 (O_1162,N_8782,N_9490);
or UO_1163 (O_1163,N_9061,N_8384);
and UO_1164 (O_1164,N_8030,N_9199);
or UO_1165 (O_1165,N_8905,N_8633);
or UO_1166 (O_1166,N_7910,N_9354);
nor UO_1167 (O_1167,N_9859,N_8137);
or UO_1168 (O_1168,N_8044,N_9760);
and UO_1169 (O_1169,N_8576,N_8760);
or UO_1170 (O_1170,N_8938,N_9996);
nor UO_1171 (O_1171,N_9640,N_8139);
and UO_1172 (O_1172,N_9810,N_8108);
xor UO_1173 (O_1173,N_9713,N_8145);
nand UO_1174 (O_1174,N_9362,N_7968);
or UO_1175 (O_1175,N_8781,N_8859);
nand UO_1176 (O_1176,N_7817,N_7931);
nand UO_1177 (O_1177,N_7899,N_8939);
nor UO_1178 (O_1178,N_9035,N_9697);
nand UO_1179 (O_1179,N_9994,N_8111);
or UO_1180 (O_1180,N_7788,N_8785);
nand UO_1181 (O_1181,N_7822,N_9233);
nor UO_1182 (O_1182,N_8341,N_8319);
and UO_1183 (O_1183,N_8614,N_9431);
or UO_1184 (O_1184,N_7855,N_8203);
nand UO_1185 (O_1185,N_8529,N_8980);
nand UO_1186 (O_1186,N_8100,N_8259);
or UO_1187 (O_1187,N_8472,N_8730);
or UO_1188 (O_1188,N_9205,N_9318);
nand UO_1189 (O_1189,N_9343,N_8678);
nor UO_1190 (O_1190,N_9515,N_8637);
nor UO_1191 (O_1191,N_8118,N_9120);
and UO_1192 (O_1192,N_8622,N_8830);
or UO_1193 (O_1193,N_9432,N_8808);
or UO_1194 (O_1194,N_9961,N_8180);
and UO_1195 (O_1195,N_9067,N_7681);
and UO_1196 (O_1196,N_8201,N_8783);
and UO_1197 (O_1197,N_8582,N_9103);
or UO_1198 (O_1198,N_9820,N_8925);
nand UO_1199 (O_1199,N_8673,N_9533);
xor UO_1200 (O_1200,N_7732,N_8733);
nor UO_1201 (O_1201,N_9585,N_8367);
xor UO_1202 (O_1202,N_9826,N_7810);
and UO_1203 (O_1203,N_7734,N_9435);
or UO_1204 (O_1204,N_9870,N_8755);
nor UO_1205 (O_1205,N_9971,N_9499);
or UO_1206 (O_1206,N_7536,N_9868);
or UO_1207 (O_1207,N_7955,N_7898);
xor UO_1208 (O_1208,N_8521,N_8230);
and UO_1209 (O_1209,N_8354,N_9662);
or UO_1210 (O_1210,N_7568,N_8412);
or UO_1211 (O_1211,N_9940,N_9213);
nand UO_1212 (O_1212,N_9752,N_8810);
and UO_1213 (O_1213,N_7969,N_8441);
or UO_1214 (O_1214,N_9257,N_7639);
or UO_1215 (O_1215,N_7707,N_8617);
nand UO_1216 (O_1216,N_9619,N_8244);
nand UO_1217 (O_1217,N_8573,N_8671);
nand UO_1218 (O_1218,N_8053,N_7796);
and UO_1219 (O_1219,N_9656,N_9216);
or UO_1220 (O_1220,N_8871,N_8037);
nor UO_1221 (O_1221,N_8231,N_8239);
nor UO_1222 (O_1222,N_8739,N_8732);
nor UO_1223 (O_1223,N_8083,N_8160);
nand UO_1224 (O_1224,N_9234,N_8356);
nand UO_1225 (O_1225,N_9735,N_8364);
and UO_1226 (O_1226,N_8285,N_9346);
or UO_1227 (O_1227,N_7654,N_9422);
and UO_1228 (O_1228,N_8159,N_9285);
nand UO_1229 (O_1229,N_7903,N_8689);
nand UO_1230 (O_1230,N_8327,N_7656);
nor UO_1231 (O_1231,N_8719,N_8463);
and UO_1232 (O_1232,N_8670,N_9388);
nand UO_1233 (O_1233,N_8282,N_9623);
or UO_1234 (O_1234,N_7921,N_7773);
nand UO_1235 (O_1235,N_7935,N_8831);
and UO_1236 (O_1236,N_9024,N_8562);
and UO_1237 (O_1237,N_9906,N_8365);
and UO_1238 (O_1238,N_7697,N_9439);
nor UO_1239 (O_1239,N_9159,N_7754);
or UO_1240 (O_1240,N_8987,N_7667);
nor UO_1241 (O_1241,N_9726,N_8977);
and UO_1242 (O_1242,N_9534,N_9811);
or UO_1243 (O_1243,N_8308,N_8136);
nand UO_1244 (O_1244,N_9497,N_9588);
or UO_1245 (O_1245,N_8551,N_8740);
or UO_1246 (O_1246,N_8997,N_9187);
nor UO_1247 (O_1247,N_8220,N_9982);
or UO_1248 (O_1248,N_9851,N_8317);
nand UO_1249 (O_1249,N_9520,N_7886);
or UO_1250 (O_1250,N_8389,N_9131);
and UO_1251 (O_1251,N_8985,N_9679);
nor UO_1252 (O_1252,N_9709,N_8782);
nor UO_1253 (O_1253,N_8686,N_9694);
nor UO_1254 (O_1254,N_8447,N_7615);
xnor UO_1255 (O_1255,N_9818,N_8008);
and UO_1256 (O_1256,N_9128,N_9318);
or UO_1257 (O_1257,N_7747,N_9029);
and UO_1258 (O_1258,N_9317,N_9715);
or UO_1259 (O_1259,N_9858,N_9839);
nand UO_1260 (O_1260,N_7517,N_9728);
nor UO_1261 (O_1261,N_7819,N_9672);
or UO_1262 (O_1262,N_9327,N_8300);
nor UO_1263 (O_1263,N_9184,N_9463);
and UO_1264 (O_1264,N_9052,N_9009);
nor UO_1265 (O_1265,N_8219,N_8813);
nand UO_1266 (O_1266,N_8341,N_8707);
nor UO_1267 (O_1267,N_8495,N_9411);
and UO_1268 (O_1268,N_9047,N_8705);
or UO_1269 (O_1269,N_9602,N_9264);
and UO_1270 (O_1270,N_8656,N_8042);
nor UO_1271 (O_1271,N_8935,N_7677);
or UO_1272 (O_1272,N_7812,N_7855);
nor UO_1273 (O_1273,N_8787,N_8167);
or UO_1274 (O_1274,N_9307,N_9677);
nor UO_1275 (O_1275,N_8004,N_8372);
nor UO_1276 (O_1276,N_8041,N_9262);
nor UO_1277 (O_1277,N_9345,N_8637);
nand UO_1278 (O_1278,N_8451,N_9780);
nand UO_1279 (O_1279,N_9480,N_7689);
nand UO_1280 (O_1280,N_7789,N_9958);
nand UO_1281 (O_1281,N_7791,N_9324);
xnor UO_1282 (O_1282,N_8437,N_8256);
or UO_1283 (O_1283,N_9820,N_9248);
nand UO_1284 (O_1284,N_9015,N_9742);
or UO_1285 (O_1285,N_9919,N_8739);
nand UO_1286 (O_1286,N_8133,N_8505);
or UO_1287 (O_1287,N_8180,N_9713);
xor UO_1288 (O_1288,N_8583,N_9441);
nor UO_1289 (O_1289,N_8186,N_9458);
nand UO_1290 (O_1290,N_9799,N_8705);
nand UO_1291 (O_1291,N_8344,N_9309);
or UO_1292 (O_1292,N_8904,N_8361);
and UO_1293 (O_1293,N_7529,N_8519);
nor UO_1294 (O_1294,N_8129,N_9577);
nor UO_1295 (O_1295,N_7716,N_8475);
nor UO_1296 (O_1296,N_7848,N_8078);
nand UO_1297 (O_1297,N_7847,N_9894);
or UO_1298 (O_1298,N_8162,N_7558);
nand UO_1299 (O_1299,N_9348,N_8732);
nand UO_1300 (O_1300,N_7559,N_9072);
or UO_1301 (O_1301,N_9777,N_8716);
nor UO_1302 (O_1302,N_8079,N_7864);
or UO_1303 (O_1303,N_7514,N_8198);
or UO_1304 (O_1304,N_7930,N_9538);
nand UO_1305 (O_1305,N_7953,N_7885);
or UO_1306 (O_1306,N_9660,N_9947);
and UO_1307 (O_1307,N_7503,N_9180);
nor UO_1308 (O_1308,N_8530,N_7962);
or UO_1309 (O_1309,N_8107,N_8834);
or UO_1310 (O_1310,N_7672,N_9375);
or UO_1311 (O_1311,N_9326,N_7935);
and UO_1312 (O_1312,N_7515,N_9724);
or UO_1313 (O_1313,N_9769,N_8526);
nand UO_1314 (O_1314,N_9506,N_8845);
xor UO_1315 (O_1315,N_8779,N_9872);
nor UO_1316 (O_1316,N_8995,N_7823);
and UO_1317 (O_1317,N_8614,N_9017);
xor UO_1318 (O_1318,N_9030,N_9976);
nor UO_1319 (O_1319,N_9865,N_8880);
or UO_1320 (O_1320,N_8662,N_9900);
and UO_1321 (O_1321,N_7983,N_9211);
nand UO_1322 (O_1322,N_7956,N_8659);
nor UO_1323 (O_1323,N_9101,N_7771);
nand UO_1324 (O_1324,N_7653,N_8610);
nor UO_1325 (O_1325,N_9750,N_7675);
nand UO_1326 (O_1326,N_9176,N_8668);
or UO_1327 (O_1327,N_8961,N_7543);
and UO_1328 (O_1328,N_9790,N_9422);
or UO_1329 (O_1329,N_9977,N_9816);
nand UO_1330 (O_1330,N_9401,N_8018);
nor UO_1331 (O_1331,N_9178,N_9153);
and UO_1332 (O_1332,N_9054,N_8745);
and UO_1333 (O_1333,N_7988,N_8868);
and UO_1334 (O_1334,N_9229,N_9185);
and UO_1335 (O_1335,N_7680,N_9732);
and UO_1336 (O_1336,N_8631,N_7988);
nand UO_1337 (O_1337,N_8375,N_7806);
nor UO_1338 (O_1338,N_9962,N_9277);
or UO_1339 (O_1339,N_8055,N_8143);
and UO_1340 (O_1340,N_9430,N_9282);
and UO_1341 (O_1341,N_8748,N_8032);
and UO_1342 (O_1342,N_7853,N_8622);
or UO_1343 (O_1343,N_8867,N_8245);
and UO_1344 (O_1344,N_8464,N_9050);
nand UO_1345 (O_1345,N_9149,N_9260);
or UO_1346 (O_1346,N_8843,N_7776);
or UO_1347 (O_1347,N_7501,N_7969);
nand UO_1348 (O_1348,N_8243,N_9212);
nand UO_1349 (O_1349,N_8769,N_7597);
and UO_1350 (O_1350,N_9331,N_8665);
nand UO_1351 (O_1351,N_8238,N_7843);
nand UO_1352 (O_1352,N_8699,N_8634);
nand UO_1353 (O_1353,N_8469,N_9740);
nor UO_1354 (O_1354,N_8803,N_9373);
xnor UO_1355 (O_1355,N_9481,N_8442);
or UO_1356 (O_1356,N_9042,N_8001);
nand UO_1357 (O_1357,N_8979,N_8477);
nor UO_1358 (O_1358,N_8515,N_9397);
nand UO_1359 (O_1359,N_8403,N_9178);
nand UO_1360 (O_1360,N_8819,N_8797);
or UO_1361 (O_1361,N_8457,N_7807);
nand UO_1362 (O_1362,N_8139,N_9265);
or UO_1363 (O_1363,N_8813,N_9077);
or UO_1364 (O_1364,N_9008,N_8591);
nand UO_1365 (O_1365,N_8729,N_8889);
nand UO_1366 (O_1366,N_7662,N_8957);
nor UO_1367 (O_1367,N_9717,N_7669);
or UO_1368 (O_1368,N_9379,N_9417);
and UO_1369 (O_1369,N_8631,N_8568);
nand UO_1370 (O_1370,N_8439,N_9209);
nor UO_1371 (O_1371,N_8460,N_7975);
nor UO_1372 (O_1372,N_9420,N_7992);
and UO_1373 (O_1373,N_8228,N_9089);
nand UO_1374 (O_1374,N_8656,N_7564);
or UO_1375 (O_1375,N_9870,N_9877);
xnor UO_1376 (O_1376,N_9481,N_8747);
nand UO_1377 (O_1377,N_8189,N_9980);
or UO_1378 (O_1378,N_8776,N_7656);
nor UO_1379 (O_1379,N_9490,N_9091);
nand UO_1380 (O_1380,N_9267,N_7716);
or UO_1381 (O_1381,N_9598,N_9498);
and UO_1382 (O_1382,N_8688,N_9239);
nand UO_1383 (O_1383,N_9269,N_9400);
nor UO_1384 (O_1384,N_8266,N_9143);
and UO_1385 (O_1385,N_9000,N_9154);
nand UO_1386 (O_1386,N_8300,N_7962);
nor UO_1387 (O_1387,N_8744,N_7533);
nand UO_1388 (O_1388,N_8607,N_7945);
or UO_1389 (O_1389,N_8893,N_9619);
nand UO_1390 (O_1390,N_7564,N_8819);
and UO_1391 (O_1391,N_9638,N_8109);
nand UO_1392 (O_1392,N_8980,N_7982);
and UO_1393 (O_1393,N_9540,N_8141);
nand UO_1394 (O_1394,N_9156,N_7797);
or UO_1395 (O_1395,N_8265,N_9173);
or UO_1396 (O_1396,N_8732,N_8089);
nand UO_1397 (O_1397,N_9957,N_9601);
nor UO_1398 (O_1398,N_9581,N_9280);
nand UO_1399 (O_1399,N_9153,N_8919);
nand UO_1400 (O_1400,N_9304,N_9929);
or UO_1401 (O_1401,N_7701,N_8824);
nor UO_1402 (O_1402,N_9856,N_7680);
nand UO_1403 (O_1403,N_8234,N_9720);
xor UO_1404 (O_1404,N_9967,N_9474);
nor UO_1405 (O_1405,N_8809,N_9409);
nor UO_1406 (O_1406,N_8970,N_9693);
nand UO_1407 (O_1407,N_7983,N_8153);
and UO_1408 (O_1408,N_9561,N_8646);
and UO_1409 (O_1409,N_9698,N_7997);
nor UO_1410 (O_1410,N_9971,N_9675);
or UO_1411 (O_1411,N_9091,N_8065);
and UO_1412 (O_1412,N_8259,N_8851);
and UO_1413 (O_1413,N_9977,N_7915);
nand UO_1414 (O_1414,N_8726,N_8894);
nand UO_1415 (O_1415,N_8436,N_8082);
nor UO_1416 (O_1416,N_8825,N_9748);
nand UO_1417 (O_1417,N_8144,N_7504);
or UO_1418 (O_1418,N_7892,N_8206);
and UO_1419 (O_1419,N_9788,N_7572);
and UO_1420 (O_1420,N_8163,N_9097);
nand UO_1421 (O_1421,N_8641,N_8619);
nor UO_1422 (O_1422,N_9958,N_8452);
xnor UO_1423 (O_1423,N_9648,N_8443);
nand UO_1424 (O_1424,N_9454,N_8562);
nand UO_1425 (O_1425,N_8783,N_8649);
and UO_1426 (O_1426,N_8104,N_8747);
and UO_1427 (O_1427,N_9189,N_8946);
and UO_1428 (O_1428,N_7651,N_8599);
or UO_1429 (O_1429,N_9107,N_8094);
nand UO_1430 (O_1430,N_9603,N_8885);
and UO_1431 (O_1431,N_7758,N_8194);
xnor UO_1432 (O_1432,N_9206,N_8950);
nand UO_1433 (O_1433,N_9639,N_9308);
nand UO_1434 (O_1434,N_8645,N_9184);
xor UO_1435 (O_1435,N_9313,N_9388);
or UO_1436 (O_1436,N_8042,N_8480);
or UO_1437 (O_1437,N_7713,N_7510);
or UO_1438 (O_1438,N_7987,N_9360);
or UO_1439 (O_1439,N_9391,N_9535);
or UO_1440 (O_1440,N_9595,N_7942);
nand UO_1441 (O_1441,N_9847,N_9531);
or UO_1442 (O_1442,N_9584,N_7791);
or UO_1443 (O_1443,N_9968,N_7640);
xnor UO_1444 (O_1444,N_9691,N_7951);
nand UO_1445 (O_1445,N_8891,N_8150);
nor UO_1446 (O_1446,N_7752,N_9218);
or UO_1447 (O_1447,N_8357,N_9240);
nand UO_1448 (O_1448,N_7574,N_8951);
and UO_1449 (O_1449,N_8897,N_7808);
nand UO_1450 (O_1450,N_9172,N_7519);
nor UO_1451 (O_1451,N_8529,N_9488);
nand UO_1452 (O_1452,N_8402,N_9704);
nor UO_1453 (O_1453,N_7599,N_9648);
nand UO_1454 (O_1454,N_9488,N_9845);
nor UO_1455 (O_1455,N_8762,N_9925);
nor UO_1456 (O_1456,N_8071,N_9239);
nor UO_1457 (O_1457,N_9953,N_9208);
and UO_1458 (O_1458,N_7742,N_8152);
or UO_1459 (O_1459,N_9618,N_9913);
nand UO_1460 (O_1460,N_9054,N_8068);
nand UO_1461 (O_1461,N_9385,N_8336);
or UO_1462 (O_1462,N_9549,N_8332);
or UO_1463 (O_1463,N_9337,N_8255);
or UO_1464 (O_1464,N_9750,N_7758);
nor UO_1465 (O_1465,N_8965,N_8176);
or UO_1466 (O_1466,N_7508,N_7682);
xnor UO_1467 (O_1467,N_7896,N_9793);
or UO_1468 (O_1468,N_8143,N_8012);
and UO_1469 (O_1469,N_8653,N_8705);
and UO_1470 (O_1470,N_9718,N_7810);
nand UO_1471 (O_1471,N_9750,N_9770);
and UO_1472 (O_1472,N_9316,N_8619);
or UO_1473 (O_1473,N_9919,N_8012);
nand UO_1474 (O_1474,N_7900,N_8677);
and UO_1475 (O_1475,N_7639,N_9436);
or UO_1476 (O_1476,N_9981,N_9680);
and UO_1477 (O_1477,N_9381,N_7772);
nand UO_1478 (O_1478,N_8054,N_7858);
nand UO_1479 (O_1479,N_9877,N_9015);
nand UO_1480 (O_1480,N_9230,N_9590);
nor UO_1481 (O_1481,N_8498,N_9063);
or UO_1482 (O_1482,N_8001,N_8596);
or UO_1483 (O_1483,N_9011,N_8659);
or UO_1484 (O_1484,N_9946,N_8448);
xor UO_1485 (O_1485,N_8464,N_9924);
or UO_1486 (O_1486,N_9052,N_8632);
nor UO_1487 (O_1487,N_8049,N_9699);
nand UO_1488 (O_1488,N_8179,N_8634);
and UO_1489 (O_1489,N_7854,N_9947);
nand UO_1490 (O_1490,N_7801,N_8450);
or UO_1491 (O_1491,N_9879,N_9457);
or UO_1492 (O_1492,N_7616,N_8869);
nor UO_1493 (O_1493,N_8146,N_9939);
nand UO_1494 (O_1494,N_8848,N_8394);
nand UO_1495 (O_1495,N_8655,N_8683);
nor UO_1496 (O_1496,N_9131,N_9729);
nor UO_1497 (O_1497,N_8957,N_7584);
and UO_1498 (O_1498,N_9856,N_9029);
or UO_1499 (O_1499,N_9951,N_8922);
endmodule