module basic_750_5000_1000_25_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_103,In_145);
or U1 (N_1,In_226,In_546);
and U2 (N_2,In_218,In_306);
nor U3 (N_3,In_224,In_187);
and U4 (N_4,In_619,In_432);
or U5 (N_5,In_469,In_393);
nor U6 (N_6,In_150,In_685);
nor U7 (N_7,In_732,In_292);
and U8 (N_8,In_714,In_472);
and U9 (N_9,In_112,In_45);
and U10 (N_10,In_166,In_128);
and U11 (N_11,In_744,In_19);
nor U12 (N_12,In_660,In_505);
or U13 (N_13,In_533,In_184);
and U14 (N_14,In_658,In_480);
nand U15 (N_15,In_31,In_503);
nand U16 (N_16,In_559,In_681);
nand U17 (N_17,In_671,In_334);
and U18 (N_18,In_264,In_81);
nor U19 (N_19,In_713,In_326);
and U20 (N_20,In_720,In_21);
nor U21 (N_21,In_143,In_599);
nand U22 (N_22,In_353,In_510);
nand U23 (N_23,In_213,In_701);
nand U24 (N_24,In_664,In_277);
or U25 (N_25,In_57,In_651);
nor U26 (N_26,In_182,In_349);
nor U27 (N_27,In_662,In_422);
or U28 (N_28,In_611,In_745);
or U29 (N_29,In_108,In_598);
and U30 (N_30,In_567,In_729);
nor U31 (N_31,In_552,In_425);
and U32 (N_32,In_133,In_52);
or U33 (N_33,In_32,In_227);
nor U34 (N_34,In_618,In_613);
nor U35 (N_35,In_276,In_125);
nand U36 (N_36,In_444,In_426);
nor U37 (N_37,In_244,In_414);
nor U38 (N_38,In_54,In_581);
and U39 (N_39,In_449,In_233);
nand U40 (N_40,In_424,In_616);
xor U41 (N_41,In_695,In_48);
nor U42 (N_42,In_396,In_286);
nor U43 (N_43,In_465,In_604);
xnor U44 (N_44,In_17,In_439);
nand U45 (N_45,In_595,In_607);
or U46 (N_46,In_263,In_560);
or U47 (N_47,In_105,In_614);
nor U48 (N_48,In_654,In_222);
or U49 (N_49,In_268,In_545);
nor U50 (N_50,In_247,In_578);
nor U51 (N_51,In_78,In_121);
and U52 (N_52,In_137,In_433);
or U53 (N_53,In_294,In_482);
nand U54 (N_54,In_562,In_229);
nand U55 (N_55,In_295,In_409);
nor U56 (N_56,In_576,In_223);
nor U57 (N_57,In_82,In_259);
or U58 (N_58,In_169,In_316);
nand U59 (N_59,In_149,In_44);
and U60 (N_60,In_35,In_257);
or U61 (N_61,In_258,In_285);
and U62 (N_62,In_568,In_636);
nor U63 (N_63,In_293,In_666);
nand U64 (N_64,In_158,In_649);
nor U65 (N_65,In_534,In_357);
and U66 (N_66,In_402,In_436);
nand U67 (N_67,In_712,In_728);
nor U68 (N_68,In_127,In_321);
nor U69 (N_69,In_267,In_428);
nand U70 (N_70,In_354,In_404);
nand U71 (N_71,In_741,In_300);
nor U72 (N_72,In_352,In_629);
and U73 (N_73,In_468,In_160);
or U74 (N_74,In_39,In_539);
nor U75 (N_75,In_372,In_362);
or U76 (N_76,In_410,In_291);
or U77 (N_77,In_721,In_710);
nand U78 (N_78,In_596,In_446);
nor U79 (N_79,In_7,In_719);
and U80 (N_80,In_43,In_153);
and U81 (N_81,In_514,In_461);
nor U82 (N_82,In_711,In_689);
nand U83 (N_83,In_392,In_221);
and U84 (N_84,In_208,In_602);
or U85 (N_85,In_246,In_217);
or U86 (N_86,In_412,In_358);
and U87 (N_87,In_477,In_361);
nor U88 (N_88,In_283,In_89);
and U89 (N_89,In_189,In_168);
nor U90 (N_90,In_261,In_99);
nand U91 (N_91,In_457,In_674);
nor U92 (N_92,In_167,In_634);
nor U93 (N_93,In_415,In_517);
or U94 (N_94,In_346,In_206);
nor U95 (N_95,In_491,In_434);
nor U96 (N_96,In_110,In_542);
nand U97 (N_97,In_537,In_524);
and U98 (N_98,In_638,In_394);
nand U99 (N_99,In_126,In_216);
or U100 (N_100,In_297,In_525);
nand U101 (N_101,In_245,In_195);
or U102 (N_102,In_679,In_549);
nor U103 (N_103,In_60,In_580);
and U104 (N_104,In_579,In_210);
and U105 (N_105,In_648,In_113);
and U106 (N_106,In_156,In_502);
and U107 (N_107,In_256,In_675);
nor U108 (N_108,In_319,In_51);
and U109 (N_109,In_730,In_389);
and U110 (N_110,In_200,In_573);
and U111 (N_111,In_470,In_390);
xor U112 (N_112,In_553,In_307);
or U113 (N_113,In_355,In_138);
xor U114 (N_114,In_492,In_59);
or U115 (N_115,In_451,In_692);
nand U116 (N_116,In_521,In_661);
and U117 (N_117,In_65,In_388);
and U118 (N_118,In_459,In_11);
nor U119 (N_119,In_398,In_56);
or U120 (N_120,In_298,In_360);
and U121 (N_121,In_305,In_339);
and U122 (N_122,In_350,In_212);
nand U123 (N_123,In_38,In_624);
nand U124 (N_124,In_280,In_281);
or U125 (N_125,In_485,In_202);
and U126 (N_126,In_543,In_209);
nand U127 (N_127,In_387,In_640);
nor U128 (N_128,In_269,In_438);
and U129 (N_129,In_84,In_370);
or U130 (N_130,In_673,In_430);
or U131 (N_131,In_600,In_199);
nor U132 (N_132,In_623,In_347);
nor U133 (N_133,In_255,In_107);
nand U134 (N_134,In_464,In_344);
nand U135 (N_135,In_737,In_445);
or U136 (N_136,In_739,In_376);
nor U137 (N_137,In_136,In_76);
nor U138 (N_138,In_122,In_163);
nor U139 (N_139,In_135,In_500);
xor U140 (N_140,In_87,In_42);
and U141 (N_141,In_735,In_515);
nand U142 (N_142,In_667,In_453);
nand U143 (N_143,In_499,In_93);
and U144 (N_144,In_572,In_483);
and U145 (N_145,In_722,In_252);
nand U146 (N_146,In_192,In_141);
nand U147 (N_147,In_67,In_157);
or U148 (N_148,In_345,In_707);
nor U149 (N_149,In_311,In_119);
nor U150 (N_150,In_617,In_63);
nand U151 (N_151,In_250,In_642);
and U152 (N_152,In_518,In_315);
or U153 (N_153,In_118,In_320);
xor U154 (N_154,In_102,In_519);
nor U155 (N_155,In_249,In_2);
nor U156 (N_156,In_74,In_395);
or U157 (N_157,In_486,In_558);
or U158 (N_158,In_234,In_625);
nand U159 (N_159,In_341,In_228);
nor U160 (N_160,In_129,In_375);
and U161 (N_161,In_708,In_36);
or U162 (N_162,In_550,In_379);
nor U163 (N_163,In_363,In_70);
or U164 (N_164,In_351,In_716);
and U165 (N_165,In_6,In_225);
and U166 (N_166,In_696,In_656);
or U167 (N_167,In_570,In_565);
nor U168 (N_168,In_382,In_513);
or U169 (N_169,In_365,In_621);
nor U170 (N_170,In_639,In_569);
xnor U171 (N_171,In_597,In_338);
nand U172 (N_172,In_380,In_566);
nand U173 (N_173,In_130,In_30);
or U174 (N_174,In_232,In_207);
nand U175 (N_175,In_690,In_747);
or U176 (N_176,In_612,In_678);
nand U177 (N_177,In_564,In_5);
nand U178 (N_178,In_152,In_235);
or U179 (N_179,In_725,In_463);
nor U180 (N_180,In_717,In_508);
nand U181 (N_181,In_726,In_520);
or U182 (N_182,In_563,In_556);
or U183 (N_183,In_495,In_85);
and U184 (N_184,In_700,In_179);
and U185 (N_185,In_659,In_652);
or U186 (N_186,In_541,In_83);
and U187 (N_187,In_740,In_348);
and U188 (N_188,In_238,In_385);
or U189 (N_189,In_622,In_582);
and U190 (N_190,In_115,In_176);
nor U191 (N_191,In_254,In_475);
nand U192 (N_192,In_241,In_544);
nand U193 (N_193,In_403,In_18);
and U194 (N_194,In_615,In_274);
or U195 (N_195,In_586,In_309);
nor U196 (N_196,In_368,In_191);
and U197 (N_197,In_687,In_400);
or U198 (N_198,In_68,In_680);
nand U199 (N_199,In_683,In_460);
and U200 (N_200,In_655,In_104);
and U201 (N_201,In_72,In_62);
nand U202 (N_202,N_175,N_136);
nor U203 (N_203,In_527,In_588);
and U204 (N_204,In_427,In_496);
nand U205 (N_205,In_676,N_85);
nand U206 (N_206,In_327,In_165);
or U207 (N_207,In_738,In_69);
or U208 (N_208,N_178,N_122);
nor U209 (N_209,N_194,In_587);
nor U210 (N_210,N_33,N_142);
nor U211 (N_211,N_12,In_561);
and U212 (N_212,In_456,In_584);
or U213 (N_213,N_101,N_54);
or U214 (N_214,N_83,N_140);
nand U215 (N_215,N_191,In_507);
nor U216 (N_216,N_38,In_440);
or U217 (N_217,In_646,N_105);
or U218 (N_218,N_57,In_516);
nor U219 (N_219,In_506,In_190);
and U220 (N_220,In_605,In_201);
and U221 (N_221,In_455,N_171);
and U222 (N_222,N_126,In_431);
nor U223 (N_223,N_146,N_168);
or U224 (N_224,In_33,N_30);
or U225 (N_225,N_53,In_694);
or U226 (N_226,In_509,In_733);
and U227 (N_227,N_4,In_384);
or U228 (N_228,In_585,In_734);
and U229 (N_229,In_554,In_53);
xor U230 (N_230,In_452,In_248);
or U231 (N_231,In_178,In_330);
or U232 (N_232,In_635,In_139);
nand U233 (N_233,In_94,In_220);
or U234 (N_234,In_253,N_177);
and U235 (N_235,In_260,N_3);
nor U236 (N_236,In_219,In_186);
or U237 (N_237,In_650,N_42);
nor U238 (N_238,N_111,In_237);
and U239 (N_239,In_723,In_251);
nand U240 (N_240,In_663,In_325);
nor U241 (N_241,In_55,In_275);
or U242 (N_242,N_77,N_63);
nor U243 (N_243,In_736,N_130);
nand U244 (N_244,N_184,In_114);
or U245 (N_245,N_160,N_75);
nor U246 (N_246,In_159,N_0);
or U247 (N_247,In_287,In_462);
xor U248 (N_248,N_19,N_134);
nor U249 (N_249,In_407,N_133);
nor U250 (N_250,In_626,N_98);
and U251 (N_251,In_147,In_95);
xnor U252 (N_252,In_632,In_657);
nor U253 (N_253,N_114,N_108);
and U254 (N_254,N_107,N_155);
nand U255 (N_255,N_137,In_279);
and U256 (N_256,In_271,In_265);
nand U257 (N_257,In_479,N_127);
nor U258 (N_258,In_9,N_169);
and U259 (N_259,N_21,N_58);
and U260 (N_260,In_91,In_437);
or U261 (N_261,In_270,In_413);
and U262 (N_262,N_147,In_4);
or U263 (N_263,In_374,In_80);
nand U264 (N_264,In_644,N_123);
and U265 (N_265,In_630,In_12);
nor U266 (N_266,In_405,In_164);
nor U267 (N_267,N_56,In_501);
xnor U268 (N_268,In_243,In_124);
or U269 (N_269,In_148,N_182);
and U270 (N_270,In_123,In_131);
nor U271 (N_271,N_39,In_132);
nor U272 (N_272,In_448,In_669);
nand U273 (N_273,N_199,N_106);
and U274 (N_274,In_106,N_100);
or U275 (N_275,In_466,N_31);
and U276 (N_276,In_670,In_71);
or U277 (N_277,In_535,In_289);
or U278 (N_278,In_369,N_115);
and U279 (N_279,In_748,In_197);
nor U280 (N_280,In_242,In_704);
nor U281 (N_281,In_418,N_185);
nor U282 (N_282,In_397,In_530);
or U283 (N_283,In_627,N_102);
xnor U284 (N_284,N_196,N_35);
and U285 (N_285,In_15,In_117);
nand U286 (N_286,In_173,In_411);
nand U287 (N_287,In_272,N_188);
and U288 (N_288,N_24,N_71);
nor U289 (N_289,In_526,In_40);
nand U290 (N_290,In_668,N_153);
xor U291 (N_291,In_682,In_547);
nand U292 (N_292,In_378,N_117);
nor U293 (N_293,N_192,N_131);
nor U294 (N_294,N_65,In_196);
or U295 (N_295,In_743,In_193);
and U296 (N_296,N_64,In_447);
and U297 (N_297,N_88,In_749);
and U298 (N_298,N_23,In_24);
or U299 (N_299,In_706,In_278);
and U300 (N_300,N_72,N_70);
xnor U301 (N_301,In_46,In_308);
and U302 (N_302,In_342,In_386);
nor U303 (N_303,N_2,In_98);
and U304 (N_304,In_417,In_367);
xor U305 (N_305,In_134,N_197);
and U306 (N_306,N_44,In_49);
nand U307 (N_307,In_601,In_161);
nand U308 (N_308,In_79,In_47);
or U309 (N_309,In_691,In_312);
nor U310 (N_310,N_103,N_59);
nand U311 (N_311,N_189,In_288);
and U312 (N_312,In_188,N_14);
or U313 (N_313,In_536,N_135);
nand U314 (N_314,N_68,N_91);
or U315 (N_315,N_150,N_25);
nand U316 (N_316,In_474,In_356);
or U317 (N_317,In_609,In_577);
nand U318 (N_318,In_154,In_631);
nand U319 (N_319,In_364,In_574);
nand U320 (N_320,In_203,In_684);
nor U321 (N_321,In_467,In_481);
or U322 (N_322,In_120,In_140);
nand U323 (N_323,N_84,N_148);
or U324 (N_324,In_16,N_13);
nor U325 (N_325,In_296,In_693);
xor U326 (N_326,N_129,In_155);
and U327 (N_327,In_419,In_8);
nand U328 (N_328,N_93,In_540);
nand U329 (N_329,N_37,In_647);
and U330 (N_330,N_139,N_66);
or U331 (N_331,N_1,In_100);
and U332 (N_332,N_97,N_40);
nor U333 (N_333,N_48,N_164);
nand U334 (N_334,In_555,In_686);
and U335 (N_335,In_603,N_112);
nor U336 (N_336,N_26,In_331);
nand U337 (N_337,In_215,N_20);
nand U338 (N_338,N_159,In_0);
and U339 (N_339,In_589,In_142);
or U340 (N_340,In_214,In_284);
nand U341 (N_341,N_87,N_80);
and U342 (N_342,In_177,In_420);
nand U343 (N_343,In_512,In_231);
nand U344 (N_344,In_408,In_677);
and U345 (N_345,In_593,N_165);
nor U346 (N_346,In_435,N_173);
nand U347 (N_347,In_653,N_128);
and U348 (N_348,N_96,In_181);
nor U349 (N_349,N_69,N_181);
nand U350 (N_350,In_377,In_494);
and U351 (N_351,In_606,N_34);
nor U352 (N_352,In_273,N_156);
or U353 (N_353,N_89,In_34);
nand U354 (N_354,N_174,In_672);
or U355 (N_355,N_187,In_366);
nor U356 (N_356,In_337,In_633);
and U357 (N_357,N_198,N_158);
nand U358 (N_358,N_86,N_82);
nand U359 (N_359,N_11,In_383);
and U360 (N_360,N_49,In_10);
or U361 (N_361,In_531,In_194);
nor U362 (N_362,In_724,In_302);
or U363 (N_363,N_52,In_73);
and U364 (N_364,In_511,In_406);
nand U365 (N_365,N_79,In_443);
nand U366 (N_366,N_76,In_328);
and U367 (N_367,In_37,N_145);
and U368 (N_368,In_172,In_637);
nor U369 (N_369,In_335,In_198);
or U370 (N_370,In_340,In_594);
or U371 (N_371,N_16,In_571);
and U372 (N_372,N_152,N_17);
nor U373 (N_373,In_96,N_47);
and U374 (N_374,N_113,In_529);
nand U375 (N_375,In_14,In_471);
nand U376 (N_376,In_727,In_476);
or U377 (N_377,N_180,In_591);
nor U378 (N_378,In_109,In_92);
and U379 (N_379,In_27,In_423);
nand U380 (N_380,In_488,In_487);
or U381 (N_381,N_172,In_583);
and U382 (N_382,N_43,In_26);
or U383 (N_383,In_313,In_688);
or U384 (N_384,In_421,In_473);
nor U385 (N_385,N_67,In_75);
nand U386 (N_386,In_303,In_643);
and U387 (N_387,In_318,N_104);
nand U388 (N_388,In_641,In_211);
and U389 (N_389,In_490,In_29);
or U390 (N_390,In_329,In_262);
and U391 (N_391,N_166,In_538);
and U392 (N_392,In_180,N_183);
nor U393 (N_393,In_718,N_121);
and U394 (N_394,In_116,N_7);
nor U395 (N_395,In_175,In_266);
nand U396 (N_396,In_371,In_41);
nor U397 (N_397,In_441,In_498);
or U398 (N_398,In_322,In_25);
and U399 (N_399,N_179,In_230);
nor U400 (N_400,N_207,N_345);
nand U401 (N_401,In_282,N_301);
or U402 (N_402,N_203,N_225);
and U403 (N_403,N_318,N_341);
nand U404 (N_404,In_528,N_226);
nor U405 (N_405,N_354,In_665);
nand U406 (N_406,N_399,In_310);
nand U407 (N_407,In_58,In_183);
and U408 (N_408,In_381,N_176);
or U409 (N_409,N_190,N_235);
or U410 (N_410,In_240,N_230);
nor U411 (N_411,N_363,N_239);
nand U412 (N_412,N_227,N_283);
and U413 (N_413,In_620,N_167);
nor U414 (N_414,N_27,N_36);
or U415 (N_415,In_551,N_204);
or U416 (N_416,N_277,N_266);
nand U417 (N_417,In_504,N_248);
nor U418 (N_418,N_60,N_393);
nor U419 (N_419,N_236,N_250);
and U420 (N_420,N_157,N_374);
or U421 (N_421,In_458,N_328);
or U422 (N_422,N_347,In_359);
nor U423 (N_423,N_276,N_311);
or U424 (N_424,N_312,N_41);
and U425 (N_425,N_119,In_144);
nand U426 (N_426,N_331,N_259);
nor U427 (N_427,N_6,In_239);
nand U428 (N_428,In_592,N_219);
and U429 (N_429,N_109,N_310);
nor U430 (N_430,In_101,In_715);
nand U431 (N_431,N_395,N_270);
nand U432 (N_432,In_323,N_186);
nor U433 (N_433,N_81,N_272);
or U434 (N_434,In_66,N_246);
nor U435 (N_435,N_210,In_742);
and U436 (N_436,N_384,N_293);
or U437 (N_437,N_381,In_697);
nor U438 (N_438,N_382,In_705);
nor U439 (N_439,N_304,N_303);
or U440 (N_440,N_327,N_261);
and U441 (N_441,N_305,In_416);
and U442 (N_442,N_333,N_234);
or U443 (N_443,N_110,In_236);
nor U444 (N_444,In_343,In_628);
and U445 (N_445,N_322,N_90);
nand U446 (N_446,In_698,N_78);
nor U447 (N_447,N_221,N_255);
nor U448 (N_448,N_350,N_5);
xor U449 (N_449,N_264,N_379);
and U450 (N_450,N_398,In_548);
nor U451 (N_451,N_61,In_497);
nand U452 (N_452,N_209,In_522);
and U453 (N_453,N_278,N_380);
nor U454 (N_454,N_55,In_64);
nor U455 (N_455,N_376,N_397);
nand U456 (N_456,In_429,N_202);
nand U457 (N_457,N_271,N_231);
or U458 (N_458,N_289,In_77);
nand U459 (N_459,N_99,N_214);
nor U460 (N_460,In_699,In_317);
or U461 (N_461,N_262,N_62);
or U462 (N_462,N_299,N_257);
nand U463 (N_463,In_746,In_336);
and U464 (N_464,N_161,N_208);
nand U465 (N_465,N_233,N_280);
nand U466 (N_466,N_260,N_390);
or U467 (N_467,N_263,In_332);
and U468 (N_468,In_391,N_200);
or U469 (N_469,N_8,In_523);
and U470 (N_470,N_392,N_144);
and U471 (N_471,N_193,N_370);
or U472 (N_472,N_294,In_23);
and U473 (N_473,N_338,N_377);
or U474 (N_474,N_286,In_731);
or U475 (N_475,N_279,N_92);
nand U476 (N_476,N_275,In_608);
nand U477 (N_477,N_389,N_319);
nand U478 (N_478,In_442,N_335);
or U479 (N_479,In_703,N_375);
nand U480 (N_480,N_228,In_28);
and U481 (N_481,In_557,N_244);
and U482 (N_482,N_372,N_138);
xnor U483 (N_483,N_368,In_532);
or U484 (N_484,N_297,N_201);
and U485 (N_485,N_269,N_360);
and U486 (N_486,N_344,N_124);
nand U487 (N_487,N_18,N_290);
or U488 (N_488,N_251,N_132);
or U489 (N_489,N_274,In_299);
nor U490 (N_490,N_332,N_46);
or U491 (N_491,In_13,N_316);
or U492 (N_492,In_170,N_258);
and U493 (N_493,N_383,N_369);
xor U494 (N_494,N_391,In_61);
nor U495 (N_495,In_97,N_281);
nand U496 (N_496,In_1,In_90);
or U497 (N_497,In_709,N_321);
or U498 (N_498,N_334,N_296);
nor U499 (N_499,N_151,N_29);
xnor U500 (N_500,N_143,N_215);
nand U501 (N_501,N_359,In_645);
or U502 (N_502,N_141,In_304);
nand U503 (N_503,N_352,N_298);
and U504 (N_504,N_120,In_333);
nand U505 (N_505,N_95,N_238);
and U506 (N_506,N_254,N_306);
nor U507 (N_507,In_373,N_162);
or U508 (N_508,N_73,In_301);
nand U509 (N_509,N_163,N_116);
nor U510 (N_510,N_232,N_315);
nor U511 (N_511,N_287,N_346);
nor U512 (N_512,In_50,N_320);
and U513 (N_513,N_224,N_367);
nand U514 (N_514,N_330,N_15);
nand U515 (N_515,N_340,N_273);
and U516 (N_516,N_339,In_146);
or U517 (N_517,N_343,In_185);
nor U518 (N_518,N_282,N_229);
nand U519 (N_519,N_324,N_216);
nand U520 (N_520,N_342,N_364);
or U521 (N_521,N_74,N_241);
nor U522 (N_522,In_204,N_206);
nand U523 (N_523,N_317,In_290);
or U524 (N_524,N_348,N_240);
xor U525 (N_525,N_291,N_326);
nand U526 (N_526,N_385,N_223);
or U527 (N_527,In_151,N_212);
nor U528 (N_528,N_356,N_373);
and U529 (N_529,In_399,N_237);
nand U530 (N_530,N_351,N_355);
nand U531 (N_531,N_195,N_357);
nor U532 (N_532,In_610,N_211);
or U533 (N_533,N_51,N_336);
and U534 (N_534,In_401,In_3);
and U535 (N_535,N_362,N_245);
and U536 (N_536,N_267,N_149);
nand U537 (N_537,N_323,N_118);
nand U538 (N_538,N_394,N_378);
or U539 (N_539,In_174,N_265);
nand U540 (N_540,N_247,N_32);
or U541 (N_541,N_313,N_314);
or U542 (N_542,N_349,N_154);
nand U543 (N_543,N_371,N_329);
nor U544 (N_544,N_288,N_387);
xnor U545 (N_545,N_217,N_220);
and U546 (N_546,N_308,N_309);
or U547 (N_547,N_365,N_213);
nor U548 (N_548,N_256,In_20);
nor U549 (N_549,In_205,In_702);
nand U550 (N_550,In_450,N_388);
and U551 (N_551,N_292,N_302);
nor U552 (N_552,N_243,N_10);
and U553 (N_553,N_396,N_307);
nand U554 (N_554,N_366,N_252);
or U555 (N_555,N_28,N_218);
or U556 (N_556,N_285,N_358);
and U557 (N_557,N_170,In_590);
nand U558 (N_558,N_386,N_300);
or U559 (N_559,N_9,N_205);
and U560 (N_560,In_454,In_489);
nand U561 (N_561,In_493,In_111);
and U562 (N_562,N_22,N_268);
nor U563 (N_563,In_478,N_50);
or U564 (N_564,In_575,In_22);
nand U565 (N_565,N_284,N_242);
or U566 (N_566,In_86,In_314);
and U567 (N_567,N_249,N_325);
nand U568 (N_568,In_324,N_45);
nor U569 (N_569,In_162,N_295);
nor U570 (N_570,In_171,N_337);
and U571 (N_571,N_125,N_361);
nand U572 (N_572,N_222,In_484);
or U573 (N_573,N_94,N_353);
and U574 (N_574,In_88,N_253);
and U575 (N_575,N_349,N_90);
or U576 (N_576,In_698,N_41);
or U577 (N_577,In_645,N_236);
or U578 (N_578,N_8,In_493);
and U579 (N_579,N_125,N_372);
and U580 (N_580,In_454,N_220);
nand U581 (N_581,N_366,N_356);
and U582 (N_582,N_241,N_216);
nand U583 (N_583,N_279,N_395);
and U584 (N_584,N_255,N_398);
and U585 (N_585,N_193,In_88);
and U586 (N_586,N_398,In_22);
nand U587 (N_587,In_702,N_389);
nor U588 (N_588,In_170,In_705);
nor U589 (N_589,N_293,In_323);
nand U590 (N_590,In_523,N_249);
or U591 (N_591,N_15,N_338);
and U592 (N_592,N_299,N_154);
nand U593 (N_593,N_29,N_355);
nand U594 (N_594,N_167,N_190);
nor U595 (N_595,In_282,In_204);
and U596 (N_596,N_343,N_269);
nor U597 (N_597,N_288,N_335);
and U598 (N_598,In_88,N_46);
nor U599 (N_599,N_73,N_353);
nor U600 (N_600,N_588,N_501);
nor U601 (N_601,N_509,N_493);
or U602 (N_602,N_498,N_490);
nor U603 (N_603,N_596,N_423);
nor U604 (N_604,N_465,N_591);
or U605 (N_605,N_497,N_451);
nor U606 (N_606,N_507,N_479);
and U607 (N_607,N_569,N_529);
nand U608 (N_608,N_422,N_562);
nor U609 (N_609,N_444,N_469);
nor U610 (N_610,N_522,N_579);
or U611 (N_611,N_426,N_477);
and U612 (N_612,N_432,N_467);
xnor U613 (N_613,N_427,N_471);
and U614 (N_614,N_440,N_535);
nand U615 (N_615,N_434,N_573);
or U616 (N_616,N_474,N_534);
nand U617 (N_617,N_595,N_411);
nor U618 (N_618,N_516,N_408);
nand U619 (N_619,N_540,N_499);
or U620 (N_620,N_594,N_476);
and U621 (N_621,N_442,N_530);
and U622 (N_622,N_566,N_458);
or U623 (N_623,N_578,N_593);
nand U624 (N_624,N_407,N_401);
or U625 (N_625,N_548,N_470);
xnor U626 (N_626,N_413,N_488);
nor U627 (N_627,N_406,N_536);
nor U628 (N_628,N_544,N_425);
nor U629 (N_629,N_492,N_505);
or U630 (N_630,N_515,N_452);
nor U631 (N_631,N_478,N_409);
nand U632 (N_632,N_545,N_552);
and U633 (N_633,N_527,N_599);
nor U634 (N_634,N_561,N_405);
nand U635 (N_635,N_424,N_570);
or U636 (N_636,N_568,N_462);
nand U637 (N_637,N_495,N_463);
and U638 (N_638,N_441,N_439);
and U639 (N_639,N_494,N_503);
nand U640 (N_640,N_461,N_550);
nand U641 (N_641,N_576,N_583);
nand U642 (N_642,N_475,N_559);
nand U643 (N_643,N_485,N_443);
nor U644 (N_644,N_519,N_459);
and U645 (N_645,N_582,N_521);
or U646 (N_646,N_532,N_506);
and U647 (N_647,N_524,N_445);
nand U648 (N_648,N_400,N_549);
and U649 (N_649,N_523,N_543);
nand U650 (N_650,N_429,N_489);
or U651 (N_651,N_416,N_419);
nor U652 (N_652,N_403,N_418);
or U653 (N_653,N_435,N_455);
xor U654 (N_654,N_417,N_464);
xnor U655 (N_655,N_421,N_546);
and U656 (N_656,N_520,N_404);
and U657 (N_657,N_564,N_531);
and U658 (N_658,N_500,N_547);
and U659 (N_659,N_514,N_551);
or U660 (N_660,N_450,N_481);
nor U661 (N_661,N_597,N_473);
nor U662 (N_662,N_517,N_437);
nand U663 (N_663,N_586,N_446);
nor U664 (N_664,N_453,N_504);
and U665 (N_665,N_575,N_589);
and U666 (N_666,N_584,N_487);
and U667 (N_667,N_468,N_496);
and U668 (N_668,N_430,N_482);
and U669 (N_669,N_480,N_460);
or U670 (N_670,N_572,N_402);
nor U671 (N_671,N_454,N_431);
nor U672 (N_672,N_581,N_541);
nor U673 (N_673,N_525,N_555);
nor U674 (N_674,N_537,N_448);
or U675 (N_675,N_486,N_466);
nor U676 (N_676,N_420,N_598);
nor U677 (N_677,N_436,N_585);
nand U678 (N_678,N_574,N_433);
or U679 (N_679,N_587,N_526);
nor U680 (N_680,N_538,N_449);
and U681 (N_681,N_554,N_571);
nand U682 (N_682,N_412,N_590);
or U683 (N_683,N_428,N_491);
or U684 (N_684,N_513,N_512);
nor U685 (N_685,N_533,N_565);
or U686 (N_686,N_502,N_438);
and U687 (N_687,N_563,N_456);
nor U688 (N_688,N_560,N_483);
xor U689 (N_689,N_558,N_410);
and U690 (N_690,N_592,N_472);
nor U691 (N_691,N_556,N_415);
or U692 (N_692,N_542,N_539);
nand U693 (N_693,N_511,N_557);
nor U694 (N_694,N_577,N_553);
or U695 (N_695,N_457,N_414);
and U696 (N_696,N_567,N_484);
nand U697 (N_697,N_508,N_510);
and U698 (N_698,N_528,N_580);
nand U699 (N_699,N_447,N_518);
nand U700 (N_700,N_591,N_407);
nand U701 (N_701,N_521,N_569);
nor U702 (N_702,N_529,N_572);
and U703 (N_703,N_457,N_485);
nor U704 (N_704,N_473,N_483);
and U705 (N_705,N_553,N_430);
nor U706 (N_706,N_407,N_442);
nand U707 (N_707,N_505,N_485);
nor U708 (N_708,N_544,N_565);
and U709 (N_709,N_449,N_570);
nor U710 (N_710,N_459,N_503);
nand U711 (N_711,N_583,N_496);
nor U712 (N_712,N_505,N_405);
or U713 (N_713,N_599,N_558);
nand U714 (N_714,N_438,N_597);
and U715 (N_715,N_496,N_451);
nand U716 (N_716,N_549,N_555);
or U717 (N_717,N_456,N_544);
nand U718 (N_718,N_447,N_430);
nand U719 (N_719,N_527,N_432);
nand U720 (N_720,N_541,N_523);
and U721 (N_721,N_481,N_434);
nor U722 (N_722,N_534,N_405);
nand U723 (N_723,N_542,N_496);
nor U724 (N_724,N_528,N_408);
or U725 (N_725,N_454,N_417);
nand U726 (N_726,N_575,N_454);
nor U727 (N_727,N_478,N_562);
and U728 (N_728,N_595,N_445);
and U729 (N_729,N_507,N_412);
and U730 (N_730,N_466,N_520);
and U731 (N_731,N_552,N_405);
nor U732 (N_732,N_568,N_425);
or U733 (N_733,N_562,N_453);
nor U734 (N_734,N_578,N_464);
or U735 (N_735,N_581,N_438);
or U736 (N_736,N_551,N_473);
and U737 (N_737,N_578,N_502);
nand U738 (N_738,N_425,N_575);
nand U739 (N_739,N_525,N_488);
or U740 (N_740,N_421,N_594);
nand U741 (N_741,N_419,N_534);
and U742 (N_742,N_428,N_526);
or U743 (N_743,N_564,N_471);
or U744 (N_744,N_525,N_504);
nor U745 (N_745,N_496,N_483);
or U746 (N_746,N_570,N_419);
nand U747 (N_747,N_522,N_446);
nand U748 (N_748,N_573,N_506);
and U749 (N_749,N_508,N_482);
and U750 (N_750,N_557,N_402);
and U751 (N_751,N_544,N_525);
nor U752 (N_752,N_440,N_478);
or U753 (N_753,N_480,N_582);
and U754 (N_754,N_488,N_453);
nor U755 (N_755,N_466,N_491);
nor U756 (N_756,N_504,N_549);
nand U757 (N_757,N_565,N_597);
nand U758 (N_758,N_521,N_465);
nor U759 (N_759,N_440,N_525);
nand U760 (N_760,N_529,N_435);
or U761 (N_761,N_536,N_402);
and U762 (N_762,N_544,N_476);
or U763 (N_763,N_574,N_550);
and U764 (N_764,N_456,N_524);
or U765 (N_765,N_438,N_454);
xnor U766 (N_766,N_565,N_567);
and U767 (N_767,N_599,N_417);
or U768 (N_768,N_574,N_487);
nor U769 (N_769,N_412,N_480);
nand U770 (N_770,N_515,N_425);
or U771 (N_771,N_534,N_456);
nand U772 (N_772,N_579,N_597);
and U773 (N_773,N_515,N_531);
nand U774 (N_774,N_566,N_520);
and U775 (N_775,N_598,N_591);
nor U776 (N_776,N_589,N_400);
and U777 (N_777,N_578,N_480);
nand U778 (N_778,N_491,N_579);
nand U779 (N_779,N_520,N_436);
and U780 (N_780,N_534,N_526);
and U781 (N_781,N_531,N_566);
nor U782 (N_782,N_571,N_511);
nand U783 (N_783,N_528,N_575);
or U784 (N_784,N_511,N_580);
and U785 (N_785,N_522,N_560);
or U786 (N_786,N_434,N_459);
and U787 (N_787,N_407,N_549);
and U788 (N_788,N_574,N_563);
nand U789 (N_789,N_450,N_433);
nor U790 (N_790,N_550,N_591);
or U791 (N_791,N_547,N_414);
nand U792 (N_792,N_563,N_445);
or U793 (N_793,N_462,N_573);
nand U794 (N_794,N_523,N_419);
and U795 (N_795,N_576,N_573);
and U796 (N_796,N_424,N_544);
or U797 (N_797,N_446,N_569);
nor U798 (N_798,N_413,N_558);
nor U799 (N_799,N_447,N_588);
or U800 (N_800,N_633,N_732);
or U801 (N_801,N_673,N_710);
nand U802 (N_802,N_608,N_646);
and U803 (N_803,N_730,N_672);
nor U804 (N_804,N_799,N_707);
and U805 (N_805,N_602,N_686);
xnor U806 (N_806,N_768,N_720);
and U807 (N_807,N_795,N_688);
or U808 (N_808,N_696,N_671);
or U809 (N_809,N_796,N_702);
or U810 (N_810,N_737,N_723);
nor U811 (N_811,N_731,N_791);
nor U812 (N_812,N_647,N_625);
nor U813 (N_813,N_772,N_721);
xnor U814 (N_814,N_724,N_618);
or U815 (N_815,N_619,N_758);
nand U816 (N_816,N_783,N_652);
and U817 (N_817,N_660,N_760);
nand U818 (N_818,N_697,N_678);
nor U819 (N_819,N_653,N_711);
nor U820 (N_820,N_709,N_641);
nand U821 (N_821,N_659,N_656);
nor U822 (N_822,N_675,N_609);
nor U823 (N_823,N_769,N_704);
xor U824 (N_824,N_708,N_712);
and U825 (N_825,N_770,N_612);
nand U826 (N_826,N_606,N_763);
or U827 (N_827,N_775,N_767);
nand U828 (N_828,N_748,N_692);
and U829 (N_829,N_685,N_781);
nand U830 (N_830,N_699,N_747);
or U831 (N_831,N_741,N_668);
nor U832 (N_832,N_638,N_725);
and U833 (N_833,N_777,N_634);
nand U834 (N_834,N_687,N_679);
or U835 (N_835,N_742,N_666);
and U836 (N_836,N_753,N_705);
nor U837 (N_837,N_663,N_621);
or U838 (N_838,N_765,N_746);
or U839 (N_839,N_648,N_657);
xnor U840 (N_840,N_669,N_654);
nand U841 (N_841,N_736,N_698);
nand U842 (N_842,N_701,N_645);
and U843 (N_843,N_693,N_750);
nand U844 (N_844,N_726,N_738);
or U845 (N_845,N_745,N_706);
nor U846 (N_846,N_751,N_637);
nand U847 (N_847,N_670,N_655);
nand U848 (N_848,N_644,N_676);
or U849 (N_849,N_716,N_600);
nor U850 (N_850,N_622,N_694);
or U851 (N_851,N_623,N_662);
nor U852 (N_852,N_626,N_752);
or U853 (N_853,N_635,N_787);
or U854 (N_854,N_617,N_743);
and U855 (N_855,N_661,N_727);
nand U856 (N_856,N_757,N_689);
nor U857 (N_857,N_629,N_793);
nand U858 (N_858,N_762,N_682);
nand U859 (N_859,N_649,N_691);
or U860 (N_860,N_680,N_789);
or U861 (N_861,N_667,N_739);
nand U862 (N_862,N_761,N_613);
nor U863 (N_863,N_780,N_778);
and U864 (N_864,N_784,N_700);
nand U865 (N_865,N_722,N_630);
nand U866 (N_866,N_603,N_771);
or U867 (N_867,N_642,N_601);
nor U868 (N_868,N_733,N_684);
or U869 (N_869,N_651,N_658);
nor U870 (N_870,N_779,N_624);
or U871 (N_871,N_665,N_755);
nor U872 (N_872,N_744,N_643);
and U873 (N_873,N_610,N_766);
or U874 (N_874,N_759,N_794);
and U875 (N_875,N_632,N_614);
and U876 (N_876,N_631,N_756);
and U877 (N_877,N_717,N_628);
nor U878 (N_878,N_674,N_797);
nor U879 (N_879,N_703,N_719);
nor U880 (N_880,N_754,N_650);
or U881 (N_881,N_790,N_611);
or U882 (N_882,N_695,N_677);
and U883 (N_883,N_607,N_620);
nor U884 (N_884,N_683,N_627);
or U885 (N_885,N_639,N_798);
nand U886 (N_886,N_664,N_636);
nand U887 (N_887,N_718,N_713);
or U888 (N_888,N_640,N_735);
or U889 (N_889,N_605,N_728);
and U890 (N_890,N_792,N_788);
nand U891 (N_891,N_785,N_715);
nor U892 (N_892,N_764,N_786);
or U893 (N_893,N_734,N_681);
or U894 (N_894,N_729,N_615);
nor U895 (N_895,N_774,N_690);
and U896 (N_896,N_616,N_776);
xnor U897 (N_897,N_714,N_604);
nand U898 (N_898,N_773,N_782);
or U899 (N_899,N_740,N_749);
and U900 (N_900,N_734,N_770);
nor U901 (N_901,N_659,N_641);
nand U902 (N_902,N_656,N_679);
nor U903 (N_903,N_628,N_758);
and U904 (N_904,N_726,N_743);
and U905 (N_905,N_749,N_738);
nor U906 (N_906,N_651,N_784);
and U907 (N_907,N_780,N_664);
or U908 (N_908,N_772,N_739);
xnor U909 (N_909,N_713,N_735);
or U910 (N_910,N_743,N_644);
nor U911 (N_911,N_746,N_693);
and U912 (N_912,N_721,N_706);
nor U913 (N_913,N_729,N_719);
and U914 (N_914,N_786,N_625);
and U915 (N_915,N_751,N_709);
xnor U916 (N_916,N_684,N_708);
nand U917 (N_917,N_664,N_701);
nor U918 (N_918,N_695,N_714);
nand U919 (N_919,N_723,N_626);
nor U920 (N_920,N_730,N_627);
nor U921 (N_921,N_738,N_677);
xor U922 (N_922,N_762,N_692);
and U923 (N_923,N_775,N_654);
nor U924 (N_924,N_661,N_674);
or U925 (N_925,N_690,N_729);
or U926 (N_926,N_655,N_621);
nor U927 (N_927,N_615,N_613);
nor U928 (N_928,N_692,N_649);
nand U929 (N_929,N_729,N_663);
nor U930 (N_930,N_771,N_758);
nor U931 (N_931,N_606,N_717);
and U932 (N_932,N_793,N_657);
and U933 (N_933,N_663,N_603);
nand U934 (N_934,N_625,N_712);
nand U935 (N_935,N_614,N_654);
or U936 (N_936,N_631,N_685);
nand U937 (N_937,N_758,N_751);
or U938 (N_938,N_609,N_611);
or U939 (N_939,N_651,N_719);
nor U940 (N_940,N_724,N_613);
and U941 (N_941,N_773,N_768);
and U942 (N_942,N_784,N_786);
and U943 (N_943,N_735,N_714);
or U944 (N_944,N_717,N_635);
nor U945 (N_945,N_653,N_712);
and U946 (N_946,N_722,N_700);
nor U947 (N_947,N_718,N_795);
and U948 (N_948,N_747,N_694);
or U949 (N_949,N_683,N_795);
nor U950 (N_950,N_722,N_698);
nand U951 (N_951,N_725,N_646);
or U952 (N_952,N_610,N_746);
nor U953 (N_953,N_608,N_602);
nand U954 (N_954,N_727,N_799);
nand U955 (N_955,N_625,N_798);
or U956 (N_956,N_638,N_752);
nand U957 (N_957,N_633,N_662);
and U958 (N_958,N_765,N_684);
and U959 (N_959,N_689,N_785);
and U960 (N_960,N_690,N_742);
nor U961 (N_961,N_786,N_779);
xor U962 (N_962,N_768,N_797);
and U963 (N_963,N_752,N_727);
nor U964 (N_964,N_619,N_647);
nor U965 (N_965,N_716,N_720);
or U966 (N_966,N_683,N_727);
nor U967 (N_967,N_627,N_682);
nand U968 (N_968,N_680,N_734);
nor U969 (N_969,N_725,N_639);
nor U970 (N_970,N_634,N_607);
and U971 (N_971,N_704,N_781);
nand U972 (N_972,N_782,N_673);
nor U973 (N_973,N_726,N_774);
or U974 (N_974,N_691,N_752);
and U975 (N_975,N_755,N_774);
nand U976 (N_976,N_754,N_643);
nand U977 (N_977,N_709,N_661);
nand U978 (N_978,N_609,N_638);
nand U979 (N_979,N_708,N_738);
or U980 (N_980,N_620,N_638);
nand U981 (N_981,N_787,N_679);
and U982 (N_982,N_693,N_615);
nand U983 (N_983,N_792,N_780);
and U984 (N_984,N_605,N_730);
or U985 (N_985,N_790,N_758);
or U986 (N_986,N_607,N_771);
nand U987 (N_987,N_725,N_657);
or U988 (N_988,N_677,N_739);
and U989 (N_989,N_712,N_680);
and U990 (N_990,N_638,N_716);
nor U991 (N_991,N_700,N_746);
or U992 (N_992,N_620,N_744);
and U993 (N_993,N_728,N_759);
nand U994 (N_994,N_622,N_780);
nor U995 (N_995,N_743,N_603);
and U996 (N_996,N_679,N_711);
nand U997 (N_997,N_703,N_714);
or U998 (N_998,N_694,N_781);
nor U999 (N_999,N_620,N_735);
nor U1000 (N_1000,N_929,N_924);
and U1001 (N_1001,N_812,N_806);
or U1002 (N_1002,N_965,N_999);
or U1003 (N_1003,N_882,N_844);
nor U1004 (N_1004,N_908,N_982);
nor U1005 (N_1005,N_960,N_961);
and U1006 (N_1006,N_885,N_940);
and U1007 (N_1007,N_825,N_968);
or U1008 (N_1008,N_958,N_926);
and U1009 (N_1009,N_843,N_955);
or U1010 (N_1010,N_850,N_811);
or U1011 (N_1011,N_840,N_801);
nand U1012 (N_1012,N_925,N_935);
nor U1013 (N_1013,N_993,N_969);
and U1014 (N_1014,N_934,N_866);
nor U1015 (N_1015,N_847,N_890);
nand U1016 (N_1016,N_983,N_984);
or U1017 (N_1017,N_829,N_883);
and U1018 (N_1018,N_970,N_837);
nor U1019 (N_1019,N_985,N_978);
and U1020 (N_1020,N_810,N_942);
and U1021 (N_1021,N_817,N_859);
or U1022 (N_1022,N_876,N_899);
and U1023 (N_1023,N_887,N_805);
and U1024 (N_1024,N_877,N_977);
nor U1025 (N_1025,N_851,N_992);
and U1026 (N_1026,N_881,N_901);
nand U1027 (N_1027,N_870,N_932);
nor U1028 (N_1028,N_952,N_864);
or U1029 (N_1029,N_892,N_996);
and U1030 (N_1030,N_895,N_863);
and U1031 (N_1031,N_845,N_927);
and U1032 (N_1032,N_897,N_972);
nor U1033 (N_1033,N_914,N_893);
or U1034 (N_1034,N_944,N_909);
and U1035 (N_1035,N_994,N_918);
or U1036 (N_1036,N_900,N_808);
or U1037 (N_1037,N_821,N_902);
nor U1038 (N_1038,N_997,N_907);
or U1039 (N_1039,N_826,N_986);
nor U1040 (N_1040,N_867,N_981);
and U1041 (N_1041,N_822,N_941);
and U1042 (N_1042,N_875,N_830);
or U1043 (N_1043,N_922,N_930);
and U1044 (N_1044,N_988,N_857);
nand U1045 (N_1045,N_824,N_962);
nor U1046 (N_1046,N_838,N_879);
nand U1047 (N_1047,N_820,N_998);
and U1048 (N_1048,N_860,N_943);
and U1049 (N_1049,N_891,N_818);
and U1050 (N_1050,N_936,N_919);
or U1051 (N_1051,N_833,N_906);
nand U1052 (N_1052,N_905,N_991);
or U1053 (N_1053,N_848,N_896);
and U1054 (N_1054,N_819,N_937);
or U1055 (N_1055,N_979,N_949);
or U1056 (N_1056,N_995,N_854);
nand U1057 (N_1057,N_846,N_871);
nand U1058 (N_1058,N_974,N_976);
or U1059 (N_1059,N_853,N_872);
nand U1060 (N_1060,N_975,N_950);
nor U1061 (N_1061,N_832,N_912);
or U1062 (N_1062,N_917,N_931);
or U1063 (N_1063,N_967,N_886);
nand U1064 (N_1064,N_939,N_803);
or U1065 (N_1065,N_898,N_928);
and U1066 (N_1066,N_836,N_878);
or U1067 (N_1067,N_957,N_933);
nor U1068 (N_1068,N_959,N_880);
nand U1069 (N_1069,N_816,N_938);
and U1070 (N_1070,N_874,N_989);
or U1071 (N_1071,N_948,N_954);
nor U1072 (N_1072,N_827,N_865);
nor U1073 (N_1073,N_815,N_971);
and U1074 (N_1074,N_964,N_990);
nor U1075 (N_1075,N_868,N_953);
or U1076 (N_1076,N_894,N_921);
and U1077 (N_1077,N_861,N_945);
nand U1078 (N_1078,N_980,N_913);
and U1079 (N_1079,N_963,N_862);
or U1080 (N_1080,N_911,N_973);
and U1081 (N_1081,N_802,N_809);
and U1082 (N_1082,N_813,N_903);
nand U1083 (N_1083,N_966,N_855);
nand U1084 (N_1084,N_849,N_915);
nor U1085 (N_1085,N_923,N_807);
nand U1086 (N_1086,N_920,N_884);
nand U1087 (N_1087,N_873,N_951);
nor U1088 (N_1088,N_904,N_916);
xnor U1089 (N_1089,N_888,N_834);
nand U1090 (N_1090,N_835,N_889);
nand U1091 (N_1091,N_947,N_910);
nand U1092 (N_1092,N_956,N_852);
or U1093 (N_1093,N_814,N_987);
or U1094 (N_1094,N_800,N_842);
and U1095 (N_1095,N_841,N_839);
nor U1096 (N_1096,N_856,N_828);
or U1097 (N_1097,N_804,N_831);
and U1098 (N_1098,N_869,N_823);
nand U1099 (N_1099,N_858,N_946);
and U1100 (N_1100,N_978,N_917);
or U1101 (N_1101,N_840,N_904);
nor U1102 (N_1102,N_975,N_903);
or U1103 (N_1103,N_869,N_831);
nand U1104 (N_1104,N_947,N_908);
and U1105 (N_1105,N_944,N_922);
or U1106 (N_1106,N_825,N_996);
nor U1107 (N_1107,N_842,N_968);
xnor U1108 (N_1108,N_927,N_855);
nor U1109 (N_1109,N_908,N_939);
nand U1110 (N_1110,N_869,N_965);
or U1111 (N_1111,N_819,N_862);
nor U1112 (N_1112,N_895,N_892);
and U1113 (N_1113,N_855,N_996);
or U1114 (N_1114,N_833,N_873);
and U1115 (N_1115,N_983,N_895);
and U1116 (N_1116,N_940,N_872);
and U1117 (N_1117,N_812,N_889);
nor U1118 (N_1118,N_892,N_825);
nor U1119 (N_1119,N_893,N_998);
nand U1120 (N_1120,N_825,N_817);
nand U1121 (N_1121,N_990,N_940);
and U1122 (N_1122,N_978,N_885);
or U1123 (N_1123,N_800,N_802);
nand U1124 (N_1124,N_894,N_823);
and U1125 (N_1125,N_842,N_970);
and U1126 (N_1126,N_833,N_920);
or U1127 (N_1127,N_942,N_886);
nand U1128 (N_1128,N_936,N_810);
nor U1129 (N_1129,N_977,N_838);
or U1130 (N_1130,N_804,N_946);
nor U1131 (N_1131,N_968,N_998);
and U1132 (N_1132,N_845,N_963);
and U1133 (N_1133,N_993,N_814);
and U1134 (N_1134,N_900,N_842);
and U1135 (N_1135,N_948,N_894);
nor U1136 (N_1136,N_898,N_833);
nand U1137 (N_1137,N_954,N_883);
and U1138 (N_1138,N_956,N_920);
xnor U1139 (N_1139,N_956,N_891);
nand U1140 (N_1140,N_802,N_814);
and U1141 (N_1141,N_843,N_904);
and U1142 (N_1142,N_955,N_888);
and U1143 (N_1143,N_815,N_828);
nand U1144 (N_1144,N_951,N_827);
or U1145 (N_1145,N_850,N_831);
nor U1146 (N_1146,N_901,N_934);
xnor U1147 (N_1147,N_910,N_943);
and U1148 (N_1148,N_930,N_883);
and U1149 (N_1149,N_968,N_896);
or U1150 (N_1150,N_877,N_899);
nand U1151 (N_1151,N_822,N_931);
and U1152 (N_1152,N_830,N_911);
or U1153 (N_1153,N_957,N_863);
nand U1154 (N_1154,N_918,N_957);
and U1155 (N_1155,N_956,N_841);
or U1156 (N_1156,N_851,N_839);
nand U1157 (N_1157,N_853,N_891);
nor U1158 (N_1158,N_986,N_936);
nor U1159 (N_1159,N_924,N_933);
nor U1160 (N_1160,N_829,N_855);
or U1161 (N_1161,N_996,N_817);
nand U1162 (N_1162,N_913,N_802);
xor U1163 (N_1163,N_934,N_889);
nor U1164 (N_1164,N_812,N_929);
and U1165 (N_1165,N_853,N_918);
nand U1166 (N_1166,N_980,N_942);
or U1167 (N_1167,N_922,N_836);
xnor U1168 (N_1168,N_919,N_899);
nor U1169 (N_1169,N_849,N_803);
or U1170 (N_1170,N_866,N_833);
and U1171 (N_1171,N_956,N_948);
or U1172 (N_1172,N_890,N_920);
or U1173 (N_1173,N_856,N_928);
nand U1174 (N_1174,N_965,N_907);
nand U1175 (N_1175,N_863,N_848);
and U1176 (N_1176,N_903,N_976);
nand U1177 (N_1177,N_840,N_994);
and U1178 (N_1178,N_874,N_862);
or U1179 (N_1179,N_990,N_884);
xor U1180 (N_1180,N_936,N_918);
nand U1181 (N_1181,N_927,N_900);
or U1182 (N_1182,N_972,N_993);
and U1183 (N_1183,N_813,N_816);
or U1184 (N_1184,N_886,N_803);
nand U1185 (N_1185,N_985,N_935);
or U1186 (N_1186,N_865,N_922);
nand U1187 (N_1187,N_815,N_903);
nor U1188 (N_1188,N_982,N_901);
nand U1189 (N_1189,N_887,N_852);
nor U1190 (N_1190,N_992,N_908);
or U1191 (N_1191,N_861,N_959);
and U1192 (N_1192,N_993,N_880);
nand U1193 (N_1193,N_991,N_884);
or U1194 (N_1194,N_960,N_801);
nor U1195 (N_1195,N_977,N_870);
nand U1196 (N_1196,N_837,N_990);
nor U1197 (N_1197,N_827,N_985);
nor U1198 (N_1198,N_886,N_969);
nand U1199 (N_1199,N_897,N_828);
or U1200 (N_1200,N_1018,N_1128);
or U1201 (N_1201,N_1179,N_1173);
nand U1202 (N_1202,N_1096,N_1176);
nor U1203 (N_1203,N_1042,N_1119);
or U1204 (N_1204,N_1150,N_1022);
and U1205 (N_1205,N_1078,N_1058);
or U1206 (N_1206,N_1144,N_1052);
and U1207 (N_1207,N_1178,N_1134);
and U1208 (N_1208,N_1185,N_1064);
and U1209 (N_1209,N_1183,N_1095);
nand U1210 (N_1210,N_1169,N_1057);
nor U1211 (N_1211,N_1123,N_1067);
nand U1212 (N_1212,N_1082,N_1101);
and U1213 (N_1213,N_1046,N_1015);
nor U1214 (N_1214,N_1195,N_1040);
or U1215 (N_1215,N_1103,N_1047);
nor U1216 (N_1216,N_1072,N_1126);
nor U1217 (N_1217,N_1062,N_1154);
nor U1218 (N_1218,N_1143,N_1087);
nand U1219 (N_1219,N_1177,N_1013);
nor U1220 (N_1220,N_1085,N_1030);
nor U1221 (N_1221,N_1148,N_1175);
or U1222 (N_1222,N_1117,N_1125);
nor U1223 (N_1223,N_1019,N_1184);
and U1224 (N_1224,N_1031,N_1146);
or U1225 (N_1225,N_1011,N_1180);
or U1226 (N_1226,N_1049,N_1166);
or U1227 (N_1227,N_1159,N_1155);
nand U1228 (N_1228,N_1120,N_1055);
or U1229 (N_1229,N_1116,N_1107);
xnor U1230 (N_1230,N_1152,N_1097);
nand U1231 (N_1231,N_1182,N_1026);
nor U1232 (N_1232,N_1197,N_1017);
and U1233 (N_1233,N_1113,N_1020);
nand U1234 (N_1234,N_1187,N_1109);
nand U1235 (N_1235,N_1006,N_1198);
or U1236 (N_1236,N_1024,N_1059);
nand U1237 (N_1237,N_1135,N_1073);
nor U1238 (N_1238,N_1081,N_1147);
or U1239 (N_1239,N_1171,N_1088);
nand U1240 (N_1240,N_1194,N_1091);
nand U1241 (N_1241,N_1039,N_1048);
nor U1242 (N_1242,N_1189,N_1153);
or U1243 (N_1243,N_1043,N_1145);
nor U1244 (N_1244,N_1115,N_1190);
and U1245 (N_1245,N_1193,N_1138);
nand U1246 (N_1246,N_1075,N_1099);
nand U1247 (N_1247,N_1133,N_1137);
nor U1248 (N_1248,N_1164,N_1041);
xnor U1249 (N_1249,N_1192,N_1086);
nor U1250 (N_1250,N_1105,N_1053);
nor U1251 (N_1251,N_1002,N_1035);
or U1252 (N_1252,N_1127,N_1181);
nand U1253 (N_1253,N_1070,N_1033);
nor U1254 (N_1254,N_1162,N_1136);
nand U1255 (N_1255,N_1079,N_1151);
nand U1256 (N_1256,N_1131,N_1121);
and U1257 (N_1257,N_1023,N_1014);
nor U1258 (N_1258,N_1004,N_1060);
and U1259 (N_1259,N_1029,N_1007);
or U1260 (N_1260,N_1158,N_1037);
nor U1261 (N_1261,N_1063,N_1172);
and U1262 (N_1262,N_1074,N_1092);
nand U1263 (N_1263,N_1149,N_1094);
nand U1264 (N_1264,N_1114,N_1130);
or U1265 (N_1265,N_1199,N_1157);
and U1266 (N_1266,N_1050,N_1038);
nor U1267 (N_1267,N_1168,N_1044);
nand U1268 (N_1268,N_1084,N_1051);
nor U1269 (N_1269,N_1140,N_1065);
xor U1270 (N_1270,N_1196,N_1156);
or U1271 (N_1271,N_1142,N_1036);
nand U1272 (N_1272,N_1112,N_1139);
nand U1273 (N_1273,N_1032,N_1170);
and U1274 (N_1274,N_1005,N_1071);
nor U1275 (N_1275,N_1000,N_1034);
nand U1276 (N_1276,N_1100,N_1025);
nand U1277 (N_1277,N_1045,N_1129);
nor U1278 (N_1278,N_1161,N_1106);
nand U1279 (N_1279,N_1083,N_1098);
nand U1280 (N_1280,N_1080,N_1001);
and U1281 (N_1281,N_1016,N_1012);
nand U1282 (N_1282,N_1160,N_1104);
nor U1283 (N_1283,N_1141,N_1008);
or U1284 (N_1284,N_1054,N_1163);
and U1285 (N_1285,N_1188,N_1093);
nor U1286 (N_1286,N_1102,N_1027);
and U1287 (N_1287,N_1174,N_1028);
nand U1288 (N_1288,N_1110,N_1077);
or U1289 (N_1289,N_1010,N_1118);
or U1290 (N_1290,N_1056,N_1089);
and U1291 (N_1291,N_1124,N_1122);
nor U1292 (N_1292,N_1068,N_1167);
nand U1293 (N_1293,N_1108,N_1066);
and U1294 (N_1294,N_1090,N_1132);
or U1295 (N_1295,N_1003,N_1069);
and U1296 (N_1296,N_1076,N_1111);
and U1297 (N_1297,N_1009,N_1061);
nor U1298 (N_1298,N_1191,N_1186);
nand U1299 (N_1299,N_1021,N_1165);
and U1300 (N_1300,N_1098,N_1040);
nor U1301 (N_1301,N_1158,N_1019);
or U1302 (N_1302,N_1113,N_1150);
or U1303 (N_1303,N_1080,N_1092);
and U1304 (N_1304,N_1018,N_1150);
or U1305 (N_1305,N_1043,N_1121);
or U1306 (N_1306,N_1184,N_1068);
nand U1307 (N_1307,N_1100,N_1033);
and U1308 (N_1308,N_1043,N_1152);
nand U1309 (N_1309,N_1010,N_1162);
and U1310 (N_1310,N_1016,N_1071);
or U1311 (N_1311,N_1142,N_1034);
and U1312 (N_1312,N_1117,N_1112);
and U1313 (N_1313,N_1112,N_1099);
nor U1314 (N_1314,N_1024,N_1044);
or U1315 (N_1315,N_1149,N_1037);
nor U1316 (N_1316,N_1051,N_1080);
nor U1317 (N_1317,N_1022,N_1067);
or U1318 (N_1318,N_1041,N_1167);
and U1319 (N_1319,N_1006,N_1148);
and U1320 (N_1320,N_1100,N_1013);
or U1321 (N_1321,N_1134,N_1095);
nand U1322 (N_1322,N_1088,N_1057);
nor U1323 (N_1323,N_1031,N_1053);
nor U1324 (N_1324,N_1008,N_1029);
or U1325 (N_1325,N_1122,N_1114);
and U1326 (N_1326,N_1141,N_1187);
or U1327 (N_1327,N_1033,N_1165);
or U1328 (N_1328,N_1018,N_1035);
nor U1329 (N_1329,N_1159,N_1198);
or U1330 (N_1330,N_1145,N_1009);
nand U1331 (N_1331,N_1067,N_1050);
nor U1332 (N_1332,N_1023,N_1051);
nor U1333 (N_1333,N_1057,N_1123);
or U1334 (N_1334,N_1153,N_1193);
and U1335 (N_1335,N_1055,N_1130);
or U1336 (N_1336,N_1007,N_1069);
and U1337 (N_1337,N_1159,N_1130);
nand U1338 (N_1338,N_1112,N_1069);
nand U1339 (N_1339,N_1032,N_1113);
or U1340 (N_1340,N_1119,N_1076);
or U1341 (N_1341,N_1038,N_1088);
nor U1342 (N_1342,N_1032,N_1152);
nor U1343 (N_1343,N_1066,N_1179);
and U1344 (N_1344,N_1102,N_1089);
nor U1345 (N_1345,N_1009,N_1094);
nand U1346 (N_1346,N_1180,N_1103);
nand U1347 (N_1347,N_1024,N_1006);
nor U1348 (N_1348,N_1008,N_1167);
nor U1349 (N_1349,N_1076,N_1153);
and U1350 (N_1350,N_1093,N_1019);
nor U1351 (N_1351,N_1161,N_1179);
xor U1352 (N_1352,N_1164,N_1174);
or U1353 (N_1353,N_1010,N_1121);
or U1354 (N_1354,N_1193,N_1165);
or U1355 (N_1355,N_1108,N_1009);
nand U1356 (N_1356,N_1052,N_1167);
nand U1357 (N_1357,N_1019,N_1047);
and U1358 (N_1358,N_1086,N_1099);
or U1359 (N_1359,N_1053,N_1070);
nand U1360 (N_1360,N_1193,N_1027);
or U1361 (N_1361,N_1172,N_1029);
nand U1362 (N_1362,N_1197,N_1192);
nand U1363 (N_1363,N_1115,N_1031);
or U1364 (N_1364,N_1024,N_1035);
nor U1365 (N_1365,N_1156,N_1068);
or U1366 (N_1366,N_1042,N_1125);
or U1367 (N_1367,N_1140,N_1091);
and U1368 (N_1368,N_1154,N_1027);
or U1369 (N_1369,N_1116,N_1069);
nor U1370 (N_1370,N_1105,N_1159);
nand U1371 (N_1371,N_1086,N_1164);
nor U1372 (N_1372,N_1126,N_1178);
nor U1373 (N_1373,N_1186,N_1171);
or U1374 (N_1374,N_1051,N_1065);
nand U1375 (N_1375,N_1029,N_1017);
nor U1376 (N_1376,N_1089,N_1002);
and U1377 (N_1377,N_1149,N_1099);
nand U1378 (N_1378,N_1127,N_1068);
and U1379 (N_1379,N_1145,N_1053);
and U1380 (N_1380,N_1143,N_1198);
nand U1381 (N_1381,N_1031,N_1097);
or U1382 (N_1382,N_1162,N_1042);
and U1383 (N_1383,N_1138,N_1159);
nor U1384 (N_1384,N_1089,N_1059);
nand U1385 (N_1385,N_1163,N_1188);
nand U1386 (N_1386,N_1146,N_1076);
and U1387 (N_1387,N_1018,N_1130);
nand U1388 (N_1388,N_1028,N_1002);
or U1389 (N_1389,N_1186,N_1170);
and U1390 (N_1390,N_1167,N_1165);
or U1391 (N_1391,N_1061,N_1057);
nand U1392 (N_1392,N_1166,N_1169);
and U1393 (N_1393,N_1046,N_1109);
or U1394 (N_1394,N_1005,N_1032);
xor U1395 (N_1395,N_1150,N_1116);
or U1396 (N_1396,N_1123,N_1065);
or U1397 (N_1397,N_1055,N_1099);
nor U1398 (N_1398,N_1010,N_1094);
and U1399 (N_1399,N_1065,N_1145);
or U1400 (N_1400,N_1280,N_1241);
nor U1401 (N_1401,N_1245,N_1300);
nor U1402 (N_1402,N_1308,N_1362);
or U1403 (N_1403,N_1265,N_1311);
nor U1404 (N_1404,N_1333,N_1388);
and U1405 (N_1405,N_1361,N_1310);
nand U1406 (N_1406,N_1324,N_1318);
or U1407 (N_1407,N_1255,N_1273);
and U1408 (N_1408,N_1363,N_1332);
nand U1409 (N_1409,N_1347,N_1306);
nand U1410 (N_1410,N_1222,N_1254);
and U1411 (N_1411,N_1210,N_1367);
nor U1412 (N_1412,N_1248,N_1389);
and U1413 (N_1413,N_1329,N_1223);
nand U1414 (N_1414,N_1215,N_1337);
nor U1415 (N_1415,N_1326,N_1357);
or U1416 (N_1416,N_1396,N_1325);
nor U1417 (N_1417,N_1383,N_1239);
nand U1418 (N_1418,N_1247,N_1294);
nor U1419 (N_1419,N_1227,N_1378);
nor U1420 (N_1420,N_1240,N_1201);
and U1421 (N_1421,N_1246,N_1202);
or U1422 (N_1422,N_1236,N_1206);
or U1423 (N_1423,N_1351,N_1376);
or U1424 (N_1424,N_1216,N_1371);
or U1425 (N_1425,N_1285,N_1224);
nor U1426 (N_1426,N_1207,N_1200);
or U1427 (N_1427,N_1374,N_1252);
or U1428 (N_1428,N_1268,N_1386);
or U1429 (N_1429,N_1225,N_1307);
and U1430 (N_1430,N_1365,N_1243);
nor U1431 (N_1431,N_1276,N_1369);
nand U1432 (N_1432,N_1256,N_1314);
xor U1433 (N_1433,N_1233,N_1260);
and U1434 (N_1434,N_1286,N_1262);
or U1435 (N_1435,N_1313,N_1238);
and U1436 (N_1436,N_1397,N_1353);
nand U1437 (N_1437,N_1299,N_1282);
or U1438 (N_1438,N_1283,N_1373);
nand U1439 (N_1439,N_1387,N_1336);
nor U1440 (N_1440,N_1359,N_1334);
or U1441 (N_1441,N_1263,N_1249);
or U1442 (N_1442,N_1323,N_1296);
and U1443 (N_1443,N_1375,N_1257);
nor U1444 (N_1444,N_1281,N_1355);
nand U1445 (N_1445,N_1278,N_1392);
nand U1446 (N_1446,N_1218,N_1364);
or U1447 (N_1447,N_1350,N_1309);
and U1448 (N_1448,N_1237,N_1370);
nand U1449 (N_1449,N_1377,N_1354);
nor U1450 (N_1450,N_1228,N_1331);
nand U1451 (N_1451,N_1348,N_1208);
and U1452 (N_1452,N_1372,N_1235);
nand U1453 (N_1453,N_1293,N_1349);
and U1454 (N_1454,N_1391,N_1275);
or U1455 (N_1455,N_1244,N_1343);
nand U1456 (N_1456,N_1342,N_1279);
or U1457 (N_1457,N_1288,N_1303);
and U1458 (N_1458,N_1315,N_1234);
and U1459 (N_1459,N_1322,N_1385);
or U1460 (N_1460,N_1317,N_1312);
nor U1461 (N_1461,N_1221,N_1382);
nor U1462 (N_1462,N_1289,N_1290);
and U1463 (N_1463,N_1328,N_1345);
nor U1464 (N_1464,N_1330,N_1394);
or U1465 (N_1465,N_1226,N_1301);
and U1466 (N_1466,N_1274,N_1320);
xnor U1467 (N_1467,N_1302,N_1253);
nand U1468 (N_1468,N_1209,N_1251);
nor U1469 (N_1469,N_1380,N_1217);
nor U1470 (N_1470,N_1298,N_1214);
nor U1471 (N_1471,N_1211,N_1316);
or U1472 (N_1472,N_1384,N_1229);
xnor U1473 (N_1473,N_1203,N_1340);
or U1474 (N_1474,N_1259,N_1395);
and U1475 (N_1475,N_1284,N_1267);
nand U1476 (N_1476,N_1277,N_1272);
nor U1477 (N_1477,N_1356,N_1242);
nand U1478 (N_1478,N_1270,N_1360);
nor U1479 (N_1479,N_1379,N_1231);
nor U1480 (N_1480,N_1220,N_1258);
nand U1481 (N_1481,N_1338,N_1335);
or U1482 (N_1482,N_1297,N_1204);
nand U1483 (N_1483,N_1390,N_1381);
nor U1484 (N_1484,N_1368,N_1399);
nor U1485 (N_1485,N_1232,N_1292);
nand U1486 (N_1486,N_1269,N_1264);
and U1487 (N_1487,N_1271,N_1319);
nand U1488 (N_1488,N_1304,N_1205);
and U1489 (N_1489,N_1398,N_1341);
or U1490 (N_1490,N_1266,N_1291);
and U1491 (N_1491,N_1358,N_1230);
xnor U1492 (N_1492,N_1321,N_1261);
and U1493 (N_1493,N_1305,N_1250);
or U1494 (N_1494,N_1393,N_1339);
nand U1495 (N_1495,N_1295,N_1352);
nand U1496 (N_1496,N_1287,N_1219);
nor U1497 (N_1497,N_1213,N_1327);
nor U1498 (N_1498,N_1346,N_1212);
nand U1499 (N_1499,N_1344,N_1366);
nand U1500 (N_1500,N_1288,N_1336);
or U1501 (N_1501,N_1224,N_1391);
nand U1502 (N_1502,N_1350,N_1334);
or U1503 (N_1503,N_1328,N_1367);
nor U1504 (N_1504,N_1374,N_1213);
nand U1505 (N_1505,N_1312,N_1204);
or U1506 (N_1506,N_1366,N_1367);
nand U1507 (N_1507,N_1227,N_1217);
nand U1508 (N_1508,N_1223,N_1297);
or U1509 (N_1509,N_1334,N_1266);
or U1510 (N_1510,N_1359,N_1246);
nor U1511 (N_1511,N_1335,N_1278);
nand U1512 (N_1512,N_1361,N_1257);
or U1513 (N_1513,N_1326,N_1244);
nor U1514 (N_1514,N_1274,N_1256);
xnor U1515 (N_1515,N_1388,N_1217);
and U1516 (N_1516,N_1365,N_1258);
nand U1517 (N_1517,N_1275,N_1280);
or U1518 (N_1518,N_1277,N_1205);
and U1519 (N_1519,N_1362,N_1364);
nor U1520 (N_1520,N_1287,N_1324);
nor U1521 (N_1521,N_1369,N_1305);
nand U1522 (N_1522,N_1216,N_1339);
xor U1523 (N_1523,N_1360,N_1299);
or U1524 (N_1524,N_1224,N_1343);
nand U1525 (N_1525,N_1220,N_1348);
or U1526 (N_1526,N_1317,N_1267);
and U1527 (N_1527,N_1216,N_1281);
or U1528 (N_1528,N_1378,N_1364);
and U1529 (N_1529,N_1353,N_1243);
or U1530 (N_1530,N_1216,N_1384);
or U1531 (N_1531,N_1206,N_1391);
nor U1532 (N_1532,N_1349,N_1286);
nor U1533 (N_1533,N_1349,N_1276);
nand U1534 (N_1534,N_1271,N_1213);
nand U1535 (N_1535,N_1369,N_1215);
xnor U1536 (N_1536,N_1342,N_1240);
nand U1537 (N_1537,N_1259,N_1279);
nand U1538 (N_1538,N_1265,N_1213);
nor U1539 (N_1539,N_1320,N_1270);
nor U1540 (N_1540,N_1296,N_1398);
nand U1541 (N_1541,N_1228,N_1257);
or U1542 (N_1542,N_1226,N_1372);
nor U1543 (N_1543,N_1234,N_1349);
or U1544 (N_1544,N_1342,N_1247);
nor U1545 (N_1545,N_1367,N_1264);
nand U1546 (N_1546,N_1383,N_1357);
or U1547 (N_1547,N_1339,N_1394);
or U1548 (N_1548,N_1364,N_1379);
and U1549 (N_1549,N_1249,N_1352);
or U1550 (N_1550,N_1229,N_1396);
or U1551 (N_1551,N_1340,N_1292);
and U1552 (N_1552,N_1294,N_1357);
or U1553 (N_1553,N_1286,N_1203);
nor U1554 (N_1554,N_1257,N_1300);
nor U1555 (N_1555,N_1207,N_1362);
nor U1556 (N_1556,N_1399,N_1354);
nand U1557 (N_1557,N_1293,N_1340);
and U1558 (N_1558,N_1231,N_1206);
nor U1559 (N_1559,N_1296,N_1389);
nand U1560 (N_1560,N_1377,N_1348);
nor U1561 (N_1561,N_1383,N_1339);
and U1562 (N_1562,N_1250,N_1341);
nand U1563 (N_1563,N_1321,N_1331);
and U1564 (N_1564,N_1279,N_1234);
or U1565 (N_1565,N_1341,N_1383);
nor U1566 (N_1566,N_1392,N_1350);
xnor U1567 (N_1567,N_1379,N_1393);
nand U1568 (N_1568,N_1325,N_1226);
nand U1569 (N_1569,N_1240,N_1225);
nor U1570 (N_1570,N_1223,N_1361);
nand U1571 (N_1571,N_1292,N_1217);
or U1572 (N_1572,N_1323,N_1242);
and U1573 (N_1573,N_1286,N_1273);
and U1574 (N_1574,N_1226,N_1205);
nand U1575 (N_1575,N_1356,N_1390);
or U1576 (N_1576,N_1250,N_1232);
and U1577 (N_1577,N_1318,N_1204);
nor U1578 (N_1578,N_1311,N_1224);
nand U1579 (N_1579,N_1353,N_1263);
nand U1580 (N_1580,N_1322,N_1219);
or U1581 (N_1581,N_1384,N_1353);
and U1582 (N_1582,N_1298,N_1307);
and U1583 (N_1583,N_1261,N_1285);
and U1584 (N_1584,N_1334,N_1278);
xnor U1585 (N_1585,N_1249,N_1382);
and U1586 (N_1586,N_1205,N_1270);
nand U1587 (N_1587,N_1330,N_1238);
nand U1588 (N_1588,N_1267,N_1290);
nand U1589 (N_1589,N_1389,N_1293);
and U1590 (N_1590,N_1258,N_1285);
nor U1591 (N_1591,N_1291,N_1373);
or U1592 (N_1592,N_1381,N_1251);
nand U1593 (N_1593,N_1327,N_1231);
and U1594 (N_1594,N_1342,N_1254);
or U1595 (N_1595,N_1232,N_1397);
or U1596 (N_1596,N_1253,N_1262);
and U1597 (N_1597,N_1230,N_1226);
or U1598 (N_1598,N_1362,N_1327);
and U1599 (N_1599,N_1213,N_1204);
and U1600 (N_1600,N_1470,N_1559);
nor U1601 (N_1601,N_1407,N_1442);
nor U1602 (N_1602,N_1509,N_1441);
nor U1603 (N_1603,N_1539,N_1473);
and U1604 (N_1604,N_1452,N_1427);
or U1605 (N_1605,N_1483,N_1412);
or U1606 (N_1606,N_1578,N_1581);
or U1607 (N_1607,N_1534,N_1579);
nor U1608 (N_1608,N_1480,N_1421);
or U1609 (N_1609,N_1404,N_1532);
nand U1610 (N_1610,N_1454,N_1594);
and U1611 (N_1611,N_1546,N_1435);
or U1612 (N_1612,N_1455,N_1482);
nand U1613 (N_1613,N_1481,N_1597);
nand U1614 (N_1614,N_1447,N_1517);
nand U1615 (N_1615,N_1588,N_1484);
or U1616 (N_1616,N_1508,N_1566);
and U1617 (N_1617,N_1485,N_1431);
and U1618 (N_1618,N_1512,N_1541);
or U1619 (N_1619,N_1445,N_1433);
nor U1620 (N_1620,N_1565,N_1582);
nor U1621 (N_1621,N_1535,N_1558);
and U1622 (N_1622,N_1557,N_1591);
and U1623 (N_1623,N_1560,N_1564);
and U1624 (N_1624,N_1461,N_1444);
nor U1625 (N_1625,N_1448,N_1573);
and U1626 (N_1626,N_1527,N_1471);
nor U1627 (N_1627,N_1465,N_1569);
nand U1628 (N_1628,N_1443,N_1462);
nand U1629 (N_1629,N_1466,N_1576);
nand U1630 (N_1630,N_1515,N_1525);
nor U1631 (N_1631,N_1548,N_1472);
or U1632 (N_1632,N_1487,N_1419);
and U1633 (N_1633,N_1528,N_1577);
and U1634 (N_1634,N_1477,N_1598);
nand U1635 (N_1635,N_1493,N_1584);
nor U1636 (N_1636,N_1510,N_1556);
nor U1637 (N_1637,N_1511,N_1563);
and U1638 (N_1638,N_1550,N_1507);
or U1639 (N_1639,N_1537,N_1423);
and U1640 (N_1640,N_1592,N_1551);
and U1641 (N_1641,N_1467,N_1437);
and U1642 (N_1642,N_1439,N_1415);
or U1643 (N_1643,N_1552,N_1585);
nand U1644 (N_1644,N_1529,N_1432);
or U1645 (N_1645,N_1486,N_1418);
nand U1646 (N_1646,N_1492,N_1459);
or U1647 (N_1647,N_1436,N_1403);
and U1648 (N_1648,N_1568,N_1545);
nor U1649 (N_1649,N_1542,N_1497);
nand U1650 (N_1650,N_1434,N_1491);
and U1651 (N_1651,N_1420,N_1571);
nor U1652 (N_1652,N_1488,N_1475);
nand U1653 (N_1653,N_1496,N_1595);
and U1654 (N_1654,N_1408,N_1463);
nand U1655 (N_1655,N_1429,N_1424);
or U1656 (N_1656,N_1514,N_1458);
nor U1657 (N_1657,N_1446,N_1501);
nand U1658 (N_1658,N_1590,N_1464);
nand U1659 (N_1659,N_1468,N_1500);
nand U1660 (N_1660,N_1522,N_1416);
or U1661 (N_1661,N_1596,N_1599);
or U1662 (N_1662,N_1489,N_1479);
and U1663 (N_1663,N_1587,N_1456);
nand U1664 (N_1664,N_1440,N_1570);
nand U1665 (N_1665,N_1469,N_1575);
nand U1666 (N_1666,N_1478,N_1572);
and U1667 (N_1667,N_1502,N_1513);
or U1668 (N_1668,N_1554,N_1474);
or U1669 (N_1669,N_1521,N_1417);
nand U1670 (N_1670,N_1580,N_1504);
or U1671 (N_1671,N_1413,N_1518);
nor U1672 (N_1672,N_1505,N_1574);
and U1673 (N_1673,N_1499,N_1426);
and U1674 (N_1674,N_1457,N_1453);
or U1675 (N_1675,N_1516,N_1567);
and U1676 (N_1676,N_1506,N_1586);
or U1677 (N_1677,N_1549,N_1405);
nor U1678 (N_1678,N_1402,N_1533);
and U1679 (N_1679,N_1430,N_1410);
nand U1680 (N_1680,N_1593,N_1553);
or U1681 (N_1681,N_1526,N_1520);
nor U1682 (N_1682,N_1583,N_1409);
nor U1683 (N_1683,N_1460,N_1422);
xor U1684 (N_1684,N_1476,N_1519);
nor U1685 (N_1685,N_1530,N_1544);
or U1686 (N_1686,N_1438,N_1401);
nand U1687 (N_1687,N_1547,N_1451);
xor U1688 (N_1688,N_1494,N_1498);
or U1689 (N_1689,N_1543,N_1490);
nand U1690 (N_1690,N_1589,N_1400);
nand U1691 (N_1691,N_1428,N_1561);
or U1692 (N_1692,N_1555,N_1449);
or U1693 (N_1693,N_1524,N_1495);
nand U1694 (N_1694,N_1531,N_1536);
nand U1695 (N_1695,N_1411,N_1406);
nor U1696 (N_1696,N_1540,N_1562);
nor U1697 (N_1697,N_1538,N_1523);
nand U1698 (N_1698,N_1425,N_1503);
and U1699 (N_1699,N_1450,N_1414);
and U1700 (N_1700,N_1574,N_1577);
nand U1701 (N_1701,N_1489,N_1430);
and U1702 (N_1702,N_1589,N_1422);
and U1703 (N_1703,N_1410,N_1502);
or U1704 (N_1704,N_1554,N_1524);
and U1705 (N_1705,N_1523,N_1567);
or U1706 (N_1706,N_1533,N_1585);
and U1707 (N_1707,N_1476,N_1472);
nand U1708 (N_1708,N_1490,N_1576);
or U1709 (N_1709,N_1586,N_1418);
nor U1710 (N_1710,N_1533,N_1524);
and U1711 (N_1711,N_1441,N_1407);
or U1712 (N_1712,N_1596,N_1512);
and U1713 (N_1713,N_1568,N_1519);
nand U1714 (N_1714,N_1562,N_1505);
and U1715 (N_1715,N_1542,N_1597);
or U1716 (N_1716,N_1439,N_1591);
or U1717 (N_1717,N_1576,N_1552);
and U1718 (N_1718,N_1437,N_1531);
or U1719 (N_1719,N_1491,N_1578);
nand U1720 (N_1720,N_1455,N_1494);
xnor U1721 (N_1721,N_1531,N_1465);
nor U1722 (N_1722,N_1545,N_1453);
nor U1723 (N_1723,N_1488,N_1447);
and U1724 (N_1724,N_1462,N_1574);
xnor U1725 (N_1725,N_1410,N_1540);
nand U1726 (N_1726,N_1567,N_1556);
nor U1727 (N_1727,N_1476,N_1511);
nor U1728 (N_1728,N_1467,N_1495);
xnor U1729 (N_1729,N_1527,N_1599);
nor U1730 (N_1730,N_1596,N_1543);
and U1731 (N_1731,N_1486,N_1477);
nand U1732 (N_1732,N_1411,N_1541);
nor U1733 (N_1733,N_1531,N_1403);
nand U1734 (N_1734,N_1538,N_1550);
nor U1735 (N_1735,N_1520,N_1597);
nand U1736 (N_1736,N_1513,N_1499);
and U1737 (N_1737,N_1453,N_1558);
and U1738 (N_1738,N_1579,N_1423);
and U1739 (N_1739,N_1432,N_1578);
or U1740 (N_1740,N_1516,N_1419);
or U1741 (N_1741,N_1442,N_1536);
and U1742 (N_1742,N_1493,N_1583);
nor U1743 (N_1743,N_1427,N_1563);
or U1744 (N_1744,N_1558,N_1525);
and U1745 (N_1745,N_1437,N_1486);
or U1746 (N_1746,N_1491,N_1510);
nor U1747 (N_1747,N_1562,N_1545);
xor U1748 (N_1748,N_1599,N_1414);
xor U1749 (N_1749,N_1539,N_1597);
and U1750 (N_1750,N_1431,N_1453);
or U1751 (N_1751,N_1495,N_1442);
nand U1752 (N_1752,N_1551,N_1495);
or U1753 (N_1753,N_1409,N_1526);
or U1754 (N_1754,N_1597,N_1569);
or U1755 (N_1755,N_1502,N_1545);
or U1756 (N_1756,N_1423,N_1548);
nor U1757 (N_1757,N_1473,N_1577);
nor U1758 (N_1758,N_1465,N_1457);
xor U1759 (N_1759,N_1594,N_1463);
nand U1760 (N_1760,N_1519,N_1435);
and U1761 (N_1761,N_1520,N_1534);
nor U1762 (N_1762,N_1593,N_1497);
nor U1763 (N_1763,N_1485,N_1544);
nand U1764 (N_1764,N_1599,N_1490);
xor U1765 (N_1765,N_1451,N_1484);
nand U1766 (N_1766,N_1462,N_1429);
nand U1767 (N_1767,N_1452,N_1581);
or U1768 (N_1768,N_1453,N_1477);
and U1769 (N_1769,N_1576,N_1582);
nand U1770 (N_1770,N_1403,N_1570);
and U1771 (N_1771,N_1595,N_1540);
nor U1772 (N_1772,N_1401,N_1422);
nand U1773 (N_1773,N_1521,N_1511);
nor U1774 (N_1774,N_1519,N_1508);
or U1775 (N_1775,N_1591,N_1406);
xor U1776 (N_1776,N_1507,N_1594);
or U1777 (N_1777,N_1597,N_1550);
or U1778 (N_1778,N_1504,N_1506);
nor U1779 (N_1779,N_1517,N_1579);
nor U1780 (N_1780,N_1563,N_1404);
or U1781 (N_1781,N_1439,N_1563);
nand U1782 (N_1782,N_1425,N_1418);
nor U1783 (N_1783,N_1436,N_1483);
nand U1784 (N_1784,N_1577,N_1413);
nor U1785 (N_1785,N_1462,N_1585);
and U1786 (N_1786,N_1592,N_1508);
nand U1787 (N_1787,N_1516,N_1405);
or U1788 (N_1788,N_1419,N_1526);
nor U1789 (N_1789,N_1500,N_1566);
nand U1790 (N_1790,N_1406,N_1529);
nand U1791 (N_1791,N_1545,N_1506);
nor U1792 (N_1792,N_1528,N_1478);
or U1793 (N_1793,N_1527,N_1559);
or U1794 (N_1794,N_1555,N_1426);
or U1795 (N_1795,N_1514,N_1438);
nor U1796 (N_1796,N_1411,N_1529);
and U1797 (N_1797,N_1510,N_1558);
or U1798 (N_1798,N_1528,N_1594);
nor U1799 (N_1799,N_1576,N_1406);
and U1800 (N_1800,N_1748,N_1761);
nor U1801 (N_1801,N_1623,N_1646);
or U1802 (N_1802,N_1736,N_1638);
nor U1803 (N_1803,N_1744,N_1662);
nand U1804 (N_1804,N_1688,N_1661);
nand U1805 (N_1805,N_1706,N_1669);
nand U1806 (N_1806,N_1620,N_1626);
nor U1807 (N_1807,N_1765,N_1675);
nand U1808 (N_1808,N_1795,N_1619);
nand U1809 (N_1809,N_1693,N_1723);
nand U1810 (N_1810,N_1790,N_1618);
nand U1811 (N_1811,N_1622,N_1771);
or U1812 (N_1812,N_1658,N_1705);
nor U1813 (N_1813,N_1670,N_1787);
nand U1814 (N_1814,N_1682,N_1738);
nor U1815 (N_1815,N_1788,N_1684);
or U1816 (N_1816,N_1615,N_1660);
or U1817 (N_1817,N_1600,N_1668);
and U1818 (N_1818,N_1720,N_1613);
and U1819 (N_1819,N_1636,N_1632);
or U1820 (N_1820,N_1776,N_1757);
nand U1821 (N_1821,N_1641,N_1775);
nand U1822 (N_1822,N_1716,N_1633);
or U1823 (N_1823,N_1621,N_1731);
or U1824 (N_1824,N_1673,N_1697);
nor U1825 (N_1825,N_1650,N_1713);
nor U1826 (N_1826,N_1704,N_1778);
or U1827 (N_1827,N_1758,N_1654);
nand U1828 (N_1828,N_1612,N_1760);
nand U1829 (N_1829,N_1783,N_1610);
nand U1830 (N_1830,N_1728,N_1734);
nor U1831 (N_1831,N_1749,N_1674);
or U1832 (N_1832,N_1698,N_1784);
and U1833 (N_1833,N_1689,N_1742);
or U1834 (N_1834,N_1695,N_1782);
nand U1835 (N_1835,N_1602,N_1643);
xnor U1836 (N_1836,N_1656,N_1785);
xnor U1837 (N_1837,N_1665,N_1725);
or U1838 (N_1838,N_1666,N_1755);
nor U1839 (N_1839,N_1769,N_1735);
and U1840 (N_1840,N_1745,N_1730);
nor U1841 (N_1841,N_1694,N_1721);
nand U1842 (N_1842,N_1791,N_1649);
nor U1843 (N_1843,N_1768,N_1710);
nor U1844 (N_1844,N_1635,N_1604);
or U1845 (N_1845,N_1779,N_1740);
or U1846 (N_1846,N_1707,N_1762);
nor U1847 (N_1847,N_1630,N_1793);
and U1848 (N_1848,N_1789,N_1616);
or U1849 (N_1849,N_1756,N_1770);
and U1850 (N_1850,N_1709,N_1657);
nand U1851 (N_1851,N_1624,N_1629);
nor U1852 (N_1852,N_1644,N_1722);
nor U1853 (N_1853,N_1797,N_1772);
and U1854 (N_1854,N_1608,N_1799);
or U1855 (N_1855,N_1780,N_1691);
nor U1856 (N_1856,N_1699,N_1686);
nand U1857 (N_1857,N_1752,N_1711);
or U1858 (N_1858,N_1712,N_1690);
or U1859 (N_1859,N_1746,N_1763);
nor U1860 (N_1860,N_1727,N_1642);
or U1861 (N_1861,N_1667,N_1655);
or U1862 (N_1862,N_1733,N_1603);
nand U1863 (N_1863,N_1715,N_1634);
nand U1864 (N_1864,N_1659,N_1628);
or U1865 (N_1865,N_1743,N_1717);
nor U1866 (N_1866,N_1767,N_1773);
nand U1867 (N_1867,N_1753,N_1703);
nor U1868 (N_1868,N_1640,N_1609);
nor U1869 (N_1869,N_1648,N_1700);
nand U1870 (N_1870,N_1774,N_1671);
nand U1871 (N_1871,N_1701,N_1737);
nor U1872 (N_1872,N_1639,N_1759);
nand U1873 (N_1873,N_1677,N_1786);
nor U1874 (N_1874,N_1647,N_1676);
nor U1875 (N_1875,N_1754,N_1732);
and U1876 (N_1876,N_1702,N_1663);
or U1877 (N_1877,N_1653,N_1680);
and U1878 (N_1878,N_1781,N_1631);
nand U1879 (N_1879,N_1645,N_1714);
nand U1880 (N_1880,N_1679,N_1685);
and U1881 (N_1881,N_1692,N_1681);
or U1882 (N_1882,N_1708,N_1678);
or U1883 (N_1883,N_1696,N_1796);
and U1884 (N_1884,N_1764,N_1605);
nand U1885 (N_1885,N_1792,N_1617);
nor U1886 (N_1886,N_1687,N_1729);
nand U1887 (N_1887,N_1627,N_1672);
or U1888 (N_1888,N_1652,N_1766);
and U1889 (N_1889,N_1611,N_1637);
nor U1890 (N_1890,N_1751,N_1718);
nor U1891 (N_1891,N_1625,N_1724);
nand U1892 (N_1892,N_1651,N_1747);
nand U1893 (N_1893,N_1607,N_1794);
and U1894 (N_1894,N_1750,N_1726);
nand U1895 (N_1895,N_1741,N_1777);
and U1896 (N_1896,N_1601,N_1798);
and U1897 (N_1897,N_1683,N_1606);
or U1898 (N_1898,N_1664,N_1719);
and U1899 (N_1899,N_1614,N_1739);
nand U1900 (N_1900,N_1736,N_1646);
nor U1901 (N_1901,N_1607,N_1799);
and U1902 (N_1902,N_1657,N_1695);
and U1903 (N_1903,N_1760,N_1740);
or U1904 (N_1904,N_1617,N_1734);
and U1905 (N_1905,N_1739,N_1754);
nor U1906 (N_1906,N_1689,N_1622);
or U1907 (N_1907,N_1711,N_1703);
nand U1908 (N_1908,N_1692,N_1604);
or U1909 (N_1909,N_1625,N_1786);
and U1910 (N_1910,N_1651,N_1717);
and U1911 (N_1911,N_1734,N_1622);
nand U1912 (N_1912,N_1634,N_1638);
and U1913 (N_1913,N_1795,N_1693);
nand U1914 (N_1914,N_1788,N_1789);
and U1915 (N_1915,N_1648,N_1786);
and U1916 (N_1916,N_1629,N_1664);
or U1917 (N_1917,N_1694,N_1689);
and U1918 (N_1918,N_1680,N_1795);
nand U1919 (N_1919,N_1680,N_1764);
xor U1920 (N_1920,N_1632,N_1618);
xnor U1921 (N_1921,N_1685,N_1645);
nand U1922 (N_1922,N_1730,N_1769);
nor U1923 (N_1923,N_1716,N_1788);
and U1924 (N_1924,N_1666,N_1634);
nand U1925 (N_1925,N_1738,N_1763);
nand U1926 (N_1926,N_1714,N_1695);
xor U1927 (N_1927,N_1601,N_1674);
nand U1928 (N_1928,N_1629,N_1695);
nor U1929 (N_1929,N_1662,N_1658);
xnor U1930 (N_1930,N_1663,N_1665);
xnor U1931 (N_1931,N_1661,N_1603);
nor U1932 (N_1932,N_1659,N_1657);
nor U1933 (N_1933,N_1627,N_1699);
nand U1934 (N_1934,N_1738,N_1708);
and U1935 (N_1935,N_1612,N_1747);
xor U1936 (N_1936,N_1775,N_1771);
nand U1937 (N_1937,N_1652,N_1700);
nand U1938 (N_1938,N_1771,N_1708);
and U1939 (N_1939,N_1654,N_1796);
and U1940 (N_1940,N_1798,N_1785);
or U1941 (N_1941,N_1627,N_1670);
and U1942 (N_1942,N_1761,N_1772);
and U1943 (N_1943,N_1660,N_1709);
or U1944 (N_1944,N_1683,N_1708);
and U1945 (N_1945,N_1705,N_1641);
nand U1946 (N_1946,N_1637,N_1763);
and U1947 (N_1947,N_1669,N_1755);
and U1948 (N_1948,N_1671,N_1682);
nand U1949 (N_1949,N_1645,N_1773);
or U1950 (N_1950,N_1707,N_1795);
and U1951 (N_1951,N_1657,N_1728);
nand U1952 (N_1952,N_1747,N_1645);
nand U1953 (N_1953,N_1703,N_1616);
nor U1954 (N_1954,N_1727,N_1739);
or U1955 (N_1955,N_1618,N_1600);
nor U1956 (N_1956,N_1788,N_1625);
nor U1957 (N_1957,N_1695,N_1601);
nand U1958 (N_1958,N_1710,N_1746);
nand U1959 (N_1959,N_1795,N_1652);
or U1960 (N_1960,N_1727,N_1754);
nor U1961 (N_1961,N_1768,N_1714);
and U1962 (N_1962,N_1649,N_1737);
and U1963 (N_1963,N_1781,N_1687);
nand U1964 (N_1964,N_1774,N_1727);
nand U1965 (N_1965,N_1701,N_1774);
or U1966 (N_1966,N_1663,N_1619);
nor U1967 (N_1967,N_1700,N_1713);
and U1968 (N_1968,N_1611,N_1737);
or U1969 (N_1969,N_1683,N_1640);
or U1970 (N_1970,N_1758,N_1629);
and U1971 (N_1971,N_1683,N_1700);
or U1972 (N_1972,N_1601,N_1608);
and U1973 (N_1973,N_1726,N_1611);
and U1974 (N_1974,N_1641,N_1677);
or U1975 (N_1975,N_1624,N_1714);
or U1976 (N_1976,N_1727,N_1678);
nor U1977 (N_1977,N_1633,N_1710);
and U1978 (N_1978,N_1635,N_1640);
or U1979 (N_1979,N_1647,N_1734);
and U1980 (N_1980,N_1666,N_1609);
nor U1981 (N_1981,N_1656,N_1736);
nand U1982 (N_1982,N_1759,N_1680);
nand U1983 (N_1983,N_1719,N_1702);
nand U1984 (N_1984,N_1671,N_1673);
and U1985 (N_1985,N_1649,N_1799);
and U1986 (N_1986,N_1711,N_1604);
nor U1987 (N_1987,N_1731,N_1687);
or U1988 (N_1988,N_1617,N_1719);
or U1989 (N_1989,N_1660,N_1713);
nor U1990 (N_1990,N_1680,N_1602);
and U1991 (N_1991,N_1619,N_1742);
and U1992 (N_1992,N_1682,N_1673);
nand U1993 (N_1993,N_1694,N_1651);
or U1994 (N_1994,N_1627,N_1730);
xnor U1995 (N_1995,N_1755,N_1709);
or U1996 (N_1996,N_1788,N_1775);
nand U1997 (N_1997,N_1770,N_1758);
or U1998 (N_1998,N_1785,N_1720);
nand U1999 (N_1999,N_1643,N_1621);
nor U2000 (N_2000,N_1914,N_1801);
and U2001 (N_2001,N_1808,N_1951);
nand U2002 (N_2002,N_1950,N_1839);
nand U2003 (N_2003,N_1974,N_1867);
and U2004 (N_2004,N_1924,N_1966);
and U2005 (N_2005,N_1819,N_1946);
or U2006 (N_2006,N_1800,N_1932);
and U2007 (N_2007,N_1863,N_1810);
nor U2008 (N_2008,N_1864,N_1855);
nor U2009 (N_2009,N_1813,N_1910);
nor U2010 (N_2010,N_1917,N_1885);
nand U2011 (N_2011,N_1882,N_1991);
and U2012 (N_2012,N_1965,N_1986);
nor U2013 (N_2013,N_1967,N_1929);
nor U2014 (N_2014,N_1979,N_1846);
and U2015 (N_2015,N_1913,N_1835);
and U2016 (N_2016,N_1817,N_1812);
or U2017 (N_2017,N_1907,N_1814);
and U2018 (N_2018,N_1944,N_1978);
and U2019 (N_2019,N_1878,N_1933);
or U2020 (N_2020,N_1961,N_1927);
or U2021 (N_2021,N_1807,N_1862);
and U2022 (N_2022,N_1999,N_1942);
nand U2023 (N_2023,N_1922,N_1893);
nand U2024 (N_2024,N_1809,N_1827);
nor U2025 (N_2025,N_1925,N_1943);
nor U2026 (N_2026,N_1816,N_1840);
nor U2027 (N_2027,N_1897,N_1849);
or U2028 (N_2028,N_1815,N_1858);
nand U2029 (N_2029,N_1984,N_1805);
or U2030 (N_2030,N_1949,N_1930);
nand U2031 (N_2031,N_1877,N_1825);
nand U2032 (N_2032,N_1889,N_1952);
nand U2033 (N_2033,N_1923,N_1902);
or U2034 (N_2034,N_1912,N_1891);
and U2035 (N_2035,N_1853,N_1848);
nor U2036 (N_2036,N_1990,N_1995);
nor U2037 (N_2037,N_1982,N_1884);
nand U2038 (N_2038,N_1988,N_1935);
and U2039 (N_2039,N_1872,N_1981);
nor U2040 (N_2040,N_1919,N_1831);
or U2041 (N_2041,N_1941,N_1976);
nand U2042 (N_2042,N_1803,N_1939);
and U2043 (N_2043,N_1804,N_1994);
nand U2044 (N_2044,N_1842,N_1918);
or U2045 (N_2045,N_1873,N_1899);
nand U2046 (N_2046,N_1883,N_1880);
nor U2047 (N_2047,N_1868,N_1901);
and U2048 (N_2048,N_1894,N_1970);
nand U2049 (N_2049,N_1968,N_1953);
and U2050 (N_2050,N_1876,N_1909);
or U2051 (N_2051,N_1955,N_1983);
nand U2052 (N_2052,N_1888,N_1875);
and U2053 (N_2053,N_1911,N_1973);
nand U2054 (N_2054,N_1833,N_1856);
or U2055 (N_2055,N_1834,N_1963);
and U2056 (N_2056,N_1806,N_1900);
and U2057 (N_2057,N_1936,N_1823);
nor U2058 (N_2058,N_1860,N_1821);
nand U2059 (N_2059,N_1975,N_1904);
nand U2060 (N_2060,N_1956,N_1937);
nand U2061 (N_2061,N_1971,N_1903);
nand U2062 (N_2062,N_1836,N_1954);
and U2063 (N_2063,N_1938,N_1996);
nand U2064 (N_2064,N_1852,N_1820);
nor U2065 (N_2065,N_1920,N_1845);
xor U2066 (N_2066,N_1861,N_1998);
nand U2067 (N_2067,N_1850,N_1865);
nor U2068 (N_2068,N_1895,N_1881);
nand U2069 (N_2069,N_1972,N_1905);
or U2070 (N_2070,N_1843,N_1859);
nor U2071 (N_2071,N_1802,N_1841);
xnor U2072 (N_2072,N_1958,N_1824);
nor U2073 (N_2073,N_1989,N_1870);
nand U2074 (N_2074,N_1818,N_1811);
and U2075 (N_2075,N_1985,N_1916);
nand U2076 (N_2076,N_1987,N_1969);
or U2077 (N_2077,N_1959,N_1886);
or U2078 (N_2078,N_1945,N_1977);
or U2079 (N_2079,N_1832,N_1980);
or U2080 (N_2080,N_1993,N_1857);
or U2081 (N_2081,N_1890,N_1847);
nor U2082 (N_2082,N_1960,N_1931);
nor U2083 (N_2083,N_1915,N_1934);
nand U2084 (N_2084,N_1869,N_1822);
and U2085 (N_2085,N_1898,N_1871);
nor U2086 (N_2086,N_1948,N_1828);
nand U2087 (N_2087,N_1908,N_1892);
nor U2088 (N_2088,N_1887,N_1921);
nor U2089 (N_2089,N_1838,N_1947);
nor U2090 (N_2090,N_1992,N_1851);
nor U2091 (N_2091,N_1928,N_1957);
or U2092 (N_2092,N_1879,N_1940);
nand U2093 (N_2093,N_1964,N_1906);
and U2094 (N_2094,N_1854,N_1837);
and U2095 (N_2095,N_1926,N_1829);
nand U2096 (N_2096,N_1962,N_1896);
or U2097 (N_2097,N_1874,N_1997);
and U2098 (N_2098,N_1830,N_1844);
and U2099 (N_2099,N_1826,N_1866);
or U2100 (N_2100,N_1988,N_1817);
nor U2101 (N_2101,N_1882,N_1905);
xor U2102 (N_2102,N_1861,N_1855);
nor U2103 (N_2103,N_1872,N_1950);
nor U2104 (N_2104,N_1919,N_1813);
nor U2105 (N_2105,N_1818,N_1994);
and U2106 (N_2106,N_1829,N_1976);
nand U2107 (N_2107,N_1974,N_1939);
and U2108 (N_2108,N_1825,N_1961);
and U2109 (N_2109,N_1883,N_1825);
or U2110 (N_2110,N_1928,N_1803);
nand U2111 (N_2111,N_1845,N_1876);
and U2112 (N_2112,N_1877,N_1922);
nand U2113 (N_2113,N_1876,N_1839);
nor U2114 (N_2114,N_1884,N_1891);
and U2115 (N_2115,N_1943,N_1863);
and U2116 (N_2116,N_1917,N_1988);
and U2117 (N_2117,N_1957,N_1999);
nor U2118 (N_2118,N_1996,N_1879);
and U2119 (N_2119,N_1991,N_1822);
or U2120 (N_2120,N_1818,N_1827);
or U2121 (N_2121,N_1955,N_1925);
or U2122 (N_2122,N_1933,N_1815);
nand U2123 (N_2123,N_1922,N_1959);
or U2124 (N_2124,N_1809,N_1886);
or U2125 (N_2125,N_1878,N_1964);
or U2126 (N_2126,N_1922,N_1935);
and U2127 (N_2127,N_1991,N_1895);
nand U2128 (N_2128,N_1889,N_1894);
nand U2129 (N_2129,N_1853,N_1943);
nor U2130 (N_2130,N_1837,N_1956);
and U2131 (N_2131,N_1913,N_1863);
or U2132 (N_2132,N_1836,N_1927);
nand U2133 (N_2133,N_1816,N_1824);
nor U2134 (N_2134,N_1851,N_1980);
or U2135 (N_2135,N_1868,N_1872);
nor U2136 (N_2136,N_1887,N_1929);
nand U2137 (N_2137,N_1964,N_1991);
and U2138 (N_2138,N_1836,N_1951);
nor U2139 (N_2139,N_1956,N_1866);
and U2140 (N_2140,N_1804,N_1888);
or U2141 (N_2141,N_1948,N_1877);
nand U2142 (N_2142,N_1808,N_1905);
nand U2143 (N_2143,N_1978,N_1887);
nand U2144 (N_2144,N_1958,N_1820);
nor U2145 (N_2145,N_1874,N_1944);
or U2146 (N_2146,N_1947,N_1803);
and U2147 (N_2147,N_1806,N_1906);
or U2148 (N_2148,N_1930,N_1854);
and U2149 (N_2149,N_1908,N_1871);
and U2150 (N_2150,N_1912,N_1838);
nand U2151 (N_2151,N_1853,N_1924);
nor U2152 (N_2152,N_1990,N_1805);
nor U2153 (N_2153,N_1873,N_1875);
or U2154 (N_2154,N_1995,N_1959);
nand U2155 (N_2155,N_1826,N_1964);
and U2156 (N_2156,N_1838,N_1858);
nor U2157 (N_2157,N_1830,N_1911);
nand U2158 (N_2158,N_1978,N_1822);
nor U2159 (N_2159,N_1958,N_1910);
and U2160 (N_2160,N_1819,N_1926);
nand U2161 (N_2161,N_1989,N_1931);
nand U2162 (N_2162,N_1999,N_1890);
and U2163 (N_2163,N_1867,N_1874);
and U2164 (N_2164,N_1990,N_1851);
and U2165 (N_2165,N_1881,N_1934);
nor U2166 (N_2166,N_1956,N_1962);
or U2167 (N_2167,N_1802,N_1912);
nor U2168 (N_2168,N_1800,N_1804);
nand U2169 (N_2169,N_1979,N_1972);
xnor U2170 (N_2170,N_1834,N_1962);
or U2171 (N_2171,N_1825,N_1904);
and U2172 (N_2172,N_1811,N_1908);
and U2173 (N_2173,N_1913,N_1887);
and U2174 (N_2174,N_1947,N_1989);
and U2175 (N_2175,N_1988,N_1853);
or U2176 (N_2176,N_1921,N_1997);
or U2177 (N_2177,N_1983,N_1901);
nor U2178 (N_2178,N_1885,N_1854);
or U2179 (N_2179,N_1896,N_1937);
or U2180 (N_2180,N_1995,N_1950);
or U2181 (N_2181,N_1917,N_1870);
nor U2182 (N_2182,N_1979,N_1836);
and U2183 (N_2183,N_1922,N_1813);
nand U2184 (N_2184,N_1812,N_1990);
and U2185 (N_2185,N_1966,N_1981);
or U2186 (N_2186,N_1990,N_1973);
nor U2187 (N_2187,N_1982,N_1856);
nand U2188 (N_2188,N_1881,N_1856);
or U2189 (N_2189,N_1947,N_1827);
nor U2190 (N_2190,N_1854,N_1894);
nor U2191 (N_2191,N_1920,N_1853);
nor U2192 (N_2192,N_1992,N_1804);
nand U2193 (N_2193,N_1909,N_1966);
and U2194 (N_2194,N_1968,N_1827);
or U2195 (N_2195,N_1945,N_1821);
and U2196 (N_2196,N_1903,N_1981);
nor U2197 (N_2197,N_1989,N_1814);
nor U2198 (N_2198,N_1872,N_1955);
nand U2199 (N_2199,N_1860,N_1967);
or U2200 (N_2200,N_2155,N_2027);
nand U2201 (N_2201,N_2102,N_2164);
nor U2202 (N_2202,N_2199,N_2099);
nand U2203 (N_2203,N_2119,N_2136);
or U2204 (N_2204,N_2188,N_2032);
and U2205 (N_2205,N_2106,N_2041);
nand U2206 (N_2206,N_2069,N_2175);
or U2207 (N_2207,N_2170,N_2088);
nand U2208 (N_2208,N_2085,N_2153);
and U2209 (N_2209,N_2122,N_2114);
or U2210 (N_2210,N_2142,N_2100);
or U2211 (N_2211,N_2043,N_2059);
nand U2212 (N_2212,N_2079,N_2046);
or U2213 (N_2213,N_2190,N_2137);
nand U2214 (N_2214,N_2143,N_2076);
or U2215 (N_2215,N_2140,N_2149);
nand U2216 (N_2216,N_2061,N_2166);
nor U2217 (N_2217,N_2129,N_2078);
or U2218 (N_2218,N_2081,N_2019);
xor U2219 (N_2219,N_2003,N_2031);
nor U2220 (N_2220,N_2107,N_2150);
nor U2221 (N_2221,N_2048,N_2026);
nor U2222 (N_2222,N_2089,N_2171);
nor U2223 (N_2223,N_2033,N_2062);
nand U2224 (N_2224,N_2011,N_2192);
or U2225 (N_2225,N_2118,N_2006);
nor U2226 (N_2226,N_2072,N_2065);
nor U2227 (N_2227,N_2020,N_2074);
xor U2228 (N_2228,N_2034,N_2182);
nor U2229 (N_2229,N_2144,N_2185);
or U2230 (N_2230,N_2161,N_2145);
or U2231 (N_2231,N_2193,N_2198);
and U2232 (N_2232,N_2113,N_2179);
nor U2233 (N_2233,N_2060,N_2017);
or U2234 (N_2234,N_2025,N_2131);
nand U2235 (N_2235,N_2001,N_2028);
and U2236 (N_2236,N_2035,N_2053);
nand U2237 (N_2237,N_2167,N_2178);
or U2238 (N_2238,N_2047,N_2008);
nand U2239 (N_2239,N_2024,N_2052);
and U2240 (N_2240,N_2168,N_2067);
or U2241 (N_2241,N_2049,N_2058);
nand U2242 (N_2242,N_2196,N_2101);
or U2243 (N_2243,N_2176,N_2004);
nand U2244 (N_2244,N_2138,N_2181);
and U2245 (N_2245,N_2152,N_2187);
and U2246 (N_2246,N_2189,N_2117);
nor U2247 (N_2247,N_2197,N_2042);
nand U2248 (N_2248,N_2121,N_2158);
nand U2249 (N_2249,N_2183,N_2051);
nand U2250 (N_2250,N_2038,N_2000);
and U2251 (N_2251,N_2016,N_2098);
nor U2252 (N_2252,N_2056,N_2173);
nand U2253 (N_2253,N_2125,N_2172);
and U2254 (N_2254,N_2134,N_2133);
or U2255 (N_2255,N_2021,N_2063);
nand U2256 (N_2256,N_2156,N_2116);
nor U2257 (N_2257,N_2163,N_2130);
nor U2258 (N_2258,N_2139,N_2040);
nor U2259 (N_2259,N_2087,N_2112);
nand U2260 (N_2260,N_2068,N_2007);
nor U2261 (N_2261,N_2109,N_2036);
nand U2262 (N_2262,N_2093,N_2191);
or U2263 (N_2263,N_2110,N_2055);
nor U2264 (N_2264,N_2002,N_2115);
nor U2265 (N_2265,N_2180,N_2095);
or U2266 (N_2266,N_2169,N_2165);
nand U2267 (N_2267,N_2174,N_2091);
or U2268 (N_2268,N_2023,N_2012);
nand U2269 (N_2269,N_2097,N_2005);
nand U2270 (N_2270,N_2045,N_2111);
nor U2271 (N_2271,N_2075,N_2141);
nor U2272 (N_2272,N_2177,N_2108);
nand U2273 (N_2273,N_2057,N_2037);
nand U2274 (N_2274,N_2070,N_2127);
or U2275 (N_2275,N_2154,N_2084);
or U2276 (N_2276,N_2184,N_2126);
nand U2277 (N_2277,N_2013,N_2162);
nand U2278 (N_2278,N_2157,N_2066);
xor U2279 (N_2279,N_2105,N_2080);
and U2280 (N_2280,N_2077,N_2135);
and U2281 (N_2281,N_2195,N_2092);
nor U2282 (N_2282,N_2123,N_2018);
xor U2283 (N_2283,N_2015,N_2194);
or U2284 (N_2284,N_2159,N_2071);
or U2285 (N_2285,N_2160,N_2147);
nor U2286 (N_2286,N_2044,N_2103);
and U2287 (N_2287,N_2146,N_2010);
nor U2288 (N_2288,N_2094,N_2124);
nor U2289 (N_2289,N_2014,N_2086);
and U2290 (N_2290,N_2148,N_2029);
or U2291 (N_2291,N_2128,N_2186);
nor U2292 (N_2292,N_2096,N_2039);
or U2293 (N_2293,N_2009,N_2022);
nor U2294 (N_2294,N_2054,N_2132);
or U2295 (N_2295,N_2151,N_2050);
or U2296 (N_2296,N_2104,N_2090);
or U2297 (N_2297,N_2120,N_2064);
nor U2298 (N_2298,N_2082,N_2030);
nand U2299 (N_2299,N_2083,N_2073);
and U2300 (N_2300,N_2113,N_2144);
or U2301 (N_2301,N_2180,N_2189);
and U2302 (N_2302,N_2049,N_2193);
nor U2303 (N_2303,N_2148,N_2043);
or U2304 (N_2304,N_2039,N_2121);
nand U2305 (N_2305,N_2057,N_2039);
nand U2306 (N_2306,N_2017,N_2109);
and U2307 (N_2307,N_2166,N_2027);
nor U2308 (N_2308,N_2013,N_2016);
nand U2309 (N_2309,N_2151,N_2046);
or U2310 (N_2310,N_2140,N_2027);
or U2311 (N_2311,N_2178,N_2038);
nor U2312 (N_2312,N_2007,N_2136);
or U2313 (N_2313,N_2031,N_2134);
or U2314 (N_2314,N_2038,N_2164);
and U2315 (N_2315,N_2153,N_2015);
nor U2316 (N_2316,N_2082,N_2044);
nor U2317 (N_2317,N_2116,N_2063);
nand U2318 (N_2318,N_2186,N_2192);
or U2319 (N_2319,N_2012,N_2065);
nand U2320 (N_2320,N_2168,N_2022);
and U2321 (N_2321,N_2036,N_2073);
or U2322 (N_2322,N_2054,N_2079);
nand U2323 (N_2323,N_2032,N_2132);
and U2324 (N_2324,N_2176,N_2154);
nand U2325 (N_2325,N_2176,N_2118);
nand U2326 (N_2326,N_2048,N_2010);
nor U2327 (N_2327,N_2018,N_2085);
nand U2328 (N_2328,N_2179,N_2054);
nor U2329 (N_2329,N_2085,N_2058);
nand U2330 (N_2330,N_2066,N_2158);
and U2331 (N_2331,N_2104,N_2067);
nor U2332 (N_2332,N_2023,N_2169);
and U2333 (N_2333,N_2173,N_2047);
nand U2334 (N_2334,N_2071,N_2035);
nand U2335 (N_2335,N_2171,N_2043);
or U2336 (N_2336,N_2161,N_2088);
nor U2337 (N_2337,N_2110,N_2027);
nand U2338 (N_2338,N_2009,N_2177);
and U2339 (N_2339,N_2088,N_2165);
and U2340 (N_2340,N_2129,N_2125);
nor U2341 (N_2341,N_2180,N_2090);
and U2342 (N_2342,N_2005,N_2102);
nand U2343 (N_2343,N_2064,N_2096);
and U2344 (N_2344,N_2032,N_2041);
nor U2345 (N_2345,N_2081,N_2085);
or U2346 (N_2346,N_2175,N_2138);
and U2347 (N_2347,N_2071,N_2185);
nor U2348 (N_2348,N_2115,N_2189);
nor U2349 (N_2349,N_2082,N_2135);
nor U2350 (N_2350,N_2045,N_2035);
or U2351 (N_2351,N_2078,N_2049);
xor U2352 (N_2352,N_2171,N_2076);
nand U2353 (N_2353,N_2056,N_2032);
or U2354 (N_2354,N_2050,N_2143);
or U2355 (N_2355,N_2195,N_2003);
nand U2356 (N_2356,N_2014,N_2039);
or U2357 (N_2357,N_2099,N_2067);
or U2358 (N_2358,N_2056,N_2089);
or U2359 (N_2359,N_2034,N_2018);
nand U2360 (N_2360,N_2027,N_2163);
nor U2361 (N_2361,N_2139,N_2126);
and U2362 (N_2362,N_2169,N_2156);
and U2363 (N_2363,N_2185,N_2118);
nor U2364 (N_2364,N_2017,N_2070);
nand U2365 (N_2365,N_2016,N_2060);
nand U2366 (N_2366,N_2179,N_2020);
or U2367 (N_2367,N_2018,N_2033);
nor U2368 (N_2368,N_2160,N_2140);
or U2369 (N_2369,N_2135,N_2035);
nand U2370 (N_2370,N_2195,N_2127);
nor U2371 (N_2371,N_2094,N_2191);
nor U2372 (N_2372,N_2149,N_2043);
or U2373 (N_2373,N_2189,N_2041);
nor U2374 (N_2374,N_2007,N_2187);
and U2375 (N_2375,N_2175,N_2158);
and U2376 (N_2376,N_2193,N_2102);
and U2377 (N_2377,N_2128,N_2149);
nor U2378 (N_2378,N_2064,N_2013);
and U2379 (N_2379,N_2173,N_2064);
and U2380 (N_2380,N_2173,N_2068);
nor U2381 (N_2381,N_2036,N_2190);
and U2382 (N_2382,N_2079,N_2140);
nor U2383 (N_2383,N_2191,N_2091);
nor U2384 (N_2384,N_2171,N_2017);
or U2385 (N_2385,N_2028,N_2072);
or U2386 (N_2386,N_2108,N_2082);
or U2387 (N_2387,N_2174,N_2088);
or U2388 (N_2388,N_2111,N_2179);
or U2389 (N_2389,N_2116,N_2047);
or U2390 (N_2390,N_2020,N_2053);
and U2391 (N_2391,N_2114,N_2035);
nor U2392 (N_2392,N_2091,N_2101);
or U2393 (N_2393,N_2197,N_2023);
and U2394 (N_2394,N_2180,N_2093);
nor U2395 (N_2395,N_2043,N_2169);
nand U2396 (N_2396,N_2137,N_2140);
nand U2397 (N_2397,N_2133,N_2182);
and U2398 (N_2398,N_2044,N_2034);
or U2399 (N_2399,N_2082,N_2137);
and U2400 (N_2400,N_2200,N_2213);
nor U2401 (N_2401,N_2253,N_2382);
nor U2402 (N_2402,N_2259,N_2328);
or U2403 (N_2403,N_2327,N_2243);
nand U2404 (N_2404,N_2321,N_2278);
nand U2405 (N_2405,N_2335,N_2205);
and U2406 (N_2406,N_2202,N_2386);
or U2407 (N_2407,N_2367,N_2285);
nor U2408 (N_2408,N_2393,N_2322);
and U2409 (N_2409,N_2293,N_2223);
and U2410 (N_2410,N_2358,N_2201);
nor U2411 (N_2411,N_2303,N_2371);
and U2412 (N_2412,N_2354,N_2346);
and U2413 (N_2413,N_2390,N_2206);
or U2414 (N_2414,N_2214,N_2345);
nor U2415 (N_2415,N_2272,N_2313);
xnor U2416 (N_2416,N_2210,N_2376);
nor U2417 (N_2417,N_2352,N_2226);
nand U2418 (N_2418,N_2374,N_2363);
and U2419 (N_2419,N_2227,N_2276);
nand U2420 (N_2420,N_2217,N_2391);
nor U2421 (N_2421,N_2241,N_2248);
and U2422 (N_2422,N_2294,N_2366);
nand U2423 (N_2423,N_2373,N_2331);
nand U2424 (N_2424,N_2383,N_2256);
nor U2425 (N_2425,N_2362,N_2311);
nand U2426 (N_2426,N_2280,N_2349);
and U2427 (N_2427,N_2339,N_2399);
and U2428 (N_2428,N_2242,N_2379);
nor U2429 (N_2429,N_2368,N_2320);
and U2430 (N_2430,N_2221,N_2236);
nor U2431 (N_2431,N_2282,N_2292);
nand U2432 (N_2432,N_2343,N_2329);
nand U2433 (N_2433,N_2304,N_2245);
nor U2434 (N_2434,N_2317,N_2277);
or U2435 (N_2435,N_2237,N_2244);
and U2436 (N_2436,N_2216,N_2271);
nor U2437 (N_2437,N_2232,N_2398);
or U2438 (N_2438,N_2254,N_2336);
or U2439 (N_2439,N_2359,N_2283);
nor U2440 (N_2440,N_2234,N_2301);
or U2441 (N_2441,N_2314,N_2261);
nand U2442 (N_2442,N_2364,N_2264);
nor U2443 (N_2443,N_2218,N_2255);
nor U2444 (N_2444,N_2337,N_2340);
and U2445 (N_2445,N_2394,N_2208);
nand U2446 (N_2446,N_2222,N_2342);
nor U2447 (N_2447,N_2326,N_2308);
or U2448 (N_2448,N_2257,N_2385);
or U2449 (N_2449,N_2273,N_2250);
nand U2450 (N_2450,N_2333,N_2341);
nand U2451 (N_2451,N_2330,N_2387);
or U2452 (N_2452,N_2284,N_2384);
or U2453 (N_2453,N_2246,N_2262);
and U2454 (N_2454,N_2310,N_2224);
nor U2455 (N_2455,N_2323,N_2233);
or U2456 (N_2456,N_2252,N_2377);
or U2457 (N_2457,N_2268,N_2251);
or U2458 (N_2458,N_2392,N_2319);
and U2459 (N_2459,N_2309,N_2307);
nor U2460 (N_2460,N_2360,N_2220);
or U2461 (N_2461,N_2263,N_2380);
nor U2462 (N_2462,N_2375,N_2238);
or U2463 (N_2463,N_2239,N_2300);
nor U2464 (N_2464,N_2315,N_2356);
and U2465 (N_2465,N_2297,N_2369);
nand U2466 (N_2466,N_2247,N_2290);
nand U2467 (N_2467,N_2225,N_2334);
or U2468 (N_2468,N_2215,N_2231);
or U2469 (N_2469,N_2378,N_2302);
or U2470 (N_2470,N_2355,N_2325);
or U2471 (N_2471,N_2361,N_2316);
nor U2472 (N_2472,N_2260,N_2365);
and U2473 (N_2473,N_2332,N_2372);
nand U2474 (N_2474,N_2289,N_2240);
and U2475 (N_2475,N_2228,N_2353);
nor U2476 (N_2476,N_2389,N_2298);
and U2477 (N_2477,N_2324,N_2274);
nor U2478 (N_2478,N_2204,N_2203);
nand U2479 (N_2479,N_2312,N_2318);
or U2480 (N_2480,N_2265,N_2275);
or U2481 (N_2481,N_2299,N_2267);
and U2482 (N_2482,N_2212,N_2344);
nor U2483 (N_2483,N_2295,N_2351);
nand U2484 (N_2484,N_2306,N_2207);
and U2485 (N_2485,N_2270,N_2291);
and U2486 (N_2486,N_2348,N_2209);
nor U2487 (N_2487,N_2357,N_2288);
or U2488 (N_2488,N_2305,N_2229);
xor U2489 (N_2489,N_2235,N_2396);
nor U2490 (N_2490,N_2397,N_2395);
nand U2491 (N_2491,N_2281,N_2266);
nand U2492 (N_2492,N_2249,N_2269);
or U2493 (N_2493,N_2296,N_2388);
xnor U2494 (N_2494,N_2350,N_2211);
nor U2495 (N_2495,N_2347,N_2279);
nand U2496 (N_2496,N_2219,N_2286);
xnor U2497 (N_2497,N_2370,N_2230);
or U2498 (N_2498,N_2381,N_2338);
or U2499 (N_2499,N_2258,N_2287);
nor U2500 (N_2500,N_2231,N_2380);
nand U2501 (N_2501,N_2233,N_2387);
nor U2502 (N_2502,N_2254,N_2332);
and U2503 (N_2503,N_2222,N_2344);
and U2504 (N_2504,N_2248,N_2284);
nor U2505 (N_2505,N_2288,N_2286);
nor U2506 (N_2506,N_2271,N_2343);
or U2507 (N_2507,N_2341,N_2268);
nor U2508 (N_2508,N_2220,N_2251);
and U2509 (N_2509,N_2393,N_2335);
nor U2510 (N_2510,N_2220,N_2338);
or U2511 (N_2511,N_2263,N_2324);
nor U2512 (N_2512,N_2399,N_2272);
or U2513 (N_2513,N_2212,N_2330);
or U2514 (N_2514,N_2352,N_2248);
xnor U2515 (N_2515,N_2342,N_2214);
nor U2516 (N_2516,N_2234,N_2236);
nand U2517 (N_2517,N_2345,N_2306);
or U2518 (N_2518,N_2264,N_2269);
nor U2519 (N_2519,N_2318,N_2371);
and U2520 (N_2520,N_2293,N_2366);
nor U2521 (N_2521,N_2307,N_2275);
or U2522 (N_2522,N_2397,N_2364);
nand U2523 (N_2523,N_2256,N_2243);
or U2524 (N_2524,N_2278,N_2361);
or U2525 (N_2525,N_2393,N_2383);
nand U2526 (N_2526,N_2297,N_2210);
nand U2527 (N_2527,N_2295,N_2239);
or U2528 (N_2528,N_2352,N_2242);
or U2529 (N_2529,N_2371,N_2326);
nor U2530 (N_2530,N_2266,N_2307);
nand U2531 (N_2531,N_2286,N_2367);
or U2532 (N_2532,N_2203,N_2372);
xor U2533 (N_2533,N_2303,N_2395);
or U2534 (N_2534,N_2263,N_2312);
or U2535 (N_2535,N_2211,N_2337);
nand U2536 (N_2536,N_2330,N_2262);
or U2537 (N_2537,N_2353,N_2211);
and U2538 (N_2538,N_2269,N_2310);
nand U2539 (N_2539,N_2218,N_2357);
and U2540 (N_2540,N_2331,N_2285);
nand U2541 (N_2541,N_2235,N_2368);
nand U2542 (N_2542,N_2283,N_2318);
nor U2543 (N_2543,N_2285,N_2205);
or U2544 (N_2544,N_2203,N_2388);
and U2545 (N_2545,N_2248,N_2232);
nor U2546 (N_2546,N_2384,N_2361);
nand U2547 (N_2547,N_2259,N_2373);
and U2548 (N_2548,N_2288,N_2240);
and U2549 (N_2549,N_2312,N_2332);
nor U2550 (N_2550,N_2315,N_2220);
nor U2551 (N_2551,N_2377,N_2245);
nor U2552 (N_2552,N_2336,N_2381);
nand U2553 (N_2553,N_2249,N_2352);
nor U2554 (N_2554,N_2248,N_2254);
nor U2555 (N_2555,N_2289,N_2246);
or U2556 (N_2556,N_2385,N_2366);
nand U2557 (N_2557,N_2319,N_2393);
or U2558 (N_2558,N_2324,N_2280);
and U2559 (N_2559,N_2302,N_2386);
or U2560 (N_2560,N_2348,N_2240);
or U2561 (N_2561,N_2369,N_2208);
or U2562 (N_2562,N_2237,N_2362);
nor U2563 (N_2563,N_2315,N_2230);
or U2564 (N_2564,N_2360,N_2342);
nor U2565 (N_2565,N_2312,N_2237);
or U2566 (N_2566,N_2302,N_2244);
nand U2567 (N_2567,N_2368,N_2348);
nand U2568 (N_2568,N_2387,N_2399);
nor U2569 (N_2569,N_2387,N_2356);
and U2570 (N_2570,N_2205,N_2273);
nand U2571 (N_2571,N_2353,N_2345);
and U2572 (N_2572,N_2237,N_2276);
and U2573 (N_2573,N_2350,N_2212);
nor U2574 (N_2574,N_2224,N_2311);
or U2575 (N_2575,N_2366,N_2360);
nor U2576 (N_2576,N_2382,N_2385);
nand U2577 (N_2577,N_2355,N_2379);
and U2578 (N_2578,N_2200,N_2224);
and U2579 (N_2579,N_2222,N_2360);
and U2580 (N_2580,N_2353,N_2283);
nor U2581 (N_2581,N_2286,N_2223);
or U2582 (N_2582,N_2302,N_2246);
nor U2583 (N_2583,N_2321,N_2385);
nor U2584 (N_2584,N_2285,N_2269);
nand U2585 (N_2585,N_2227,N_2299);
or U2586 (N_2586,N_2264,N_2319);
nand U2587 (N_2587,N_2210,N_2354);
or U2588 (N_2588,N_2213,N_2262);
and U2589 (N_2589,N_2398,N_2385);
or U2590 (N_2590,N_2386,N_2211);
nor U2591 (N_2591,N_2347,N_2214);
nor U2592 (N_2592,N_2349,N_2296);
or U2593 (N_2593,N_2304,N_2380);
nor U2594 (N_2594,N_2362,N_2252);
nor U2595 (N_2595,N_2324,N_2226);
or U2596 (N_2596,N_2298,N_2278);
xor U2597 (N_2597,N_2378,N_2397);
nand U2598 (N_2598,N_2221,N_2258);
nand U2599 (N_2599,N_2278,N_2243);
nor U2600 (N_2600,N_2556,N_2434);
or U2601 (N_2601,N_2500,N_2430);
or U2602 (N_2602,N_2422,N_2426);
nand U2603 (N_2603,N_2541,N_2531);
and U2604 (N_2604,N_2550,N_2424);
nor U2605 (N_2605,N_2576,N_2544);
and U2606 (N_2606,N_2429,N_2418);
xor U2607 (N_2607,N_2560,N_2586);
or U2608 (N_2608,N_2527,N_2597);
nand U2609 (N_2609,N_2431,N_2583);
and U2610 (N_2610,N_2471,N_2573);
and U2611 (N_2611,N_2548,N_2417);
nor U2612 (N_2612,N_2523,N_2534);
nor U2613 (N_2613,N_2572,N_2520);
and U2614 (N_2614,N_2469,N_2462);
nor U2615 (N_2615,N_2467,N_2524);
nand U2616 (N_2616,N_2564,N_2447);
or U2617 (N_2617,N_2588,N_2511);
or U2618 (N_2618,N_2599,N_2449);
nor U2619 (N_2619,N_2575,N_2593);
or U2620 (N_2620,N_2540,N_2587);
nand U2621 (N_2621,N_2592,N_2551);
nor U2622 (N_2622,N_2538,N_2595);
nor U2623 (N_2623,N_2488,N_2501);
or U2624 (N_2624,N_2439,N_2400);
nand U2625 (N_2625,N_2533,N_2563);
nor U2626 (N_2626,N_2427,N_2553);
nand U2627 (N_2627,N_2459,N_2454);
nor U2628 (N_2628,N_2494,N_2547);
nor U2629 (N_2629,N_2489,N_2452);
or U2630 (N_2630,N_2464,N_2582);
and U2631 (N_2631,N_2561,N_2515);
nand U2632 (N_2632,N_2596,N_2451);
and U2633 (N_2633,N_2438,N_2528);
or U2634 (N_2634,N_2537,N_2519);
or U2635 (N_2635,N_2425,N_2437);
and U2636 (N_2636,N_2457,N_2455);
nor U2637 (N_2637,N_2420,N_2441);
and U2638 (N_2638,N_2559,N_2461);
nand U2639 (N_2639,N_2409,N_2529);
or U2640 (N_2640,N_2411,N_2498);
nand U2641 (N_2641,N_2522,N_2492);
and U2642 (N_2642,N_2594,N_2401);
and U2643 (N_2643,N_2435,N_2569);
or U2644 (N_2644,N_2490,N_2468);
nand U2645 (N_2645,N_2472,N_2482);
xor U2646 (N_2646,N_2562,N_2578);
or U2647 (N_2647,N_2443,N_2549);
nor U2648 (N_2648,N_2580,N_2480);
and U2649 (N_2649,N_2446,N_2554);
xnor U2650 (N_2650,N_2479,N_2558);
xor U2651 (N_2651,N_2581,N_2502);
nand U2652 (N_2652,N_2440,N_2445);
nand U2653 (N_2653,N_2516,N_2495);
nand U2654 (N_2654,N_2530,N_2466);
or U2655 (N_2655,N_2465,N_2532);
nand U2656 (N_2656,N_2407,N_2448);
nor U2657 (N_2657,N_2566,N_2470);
and U2658 (N_2658,N_2539,N_2496);
nor U2659 (N_2659,N_2460,N_2476);
and U2660 (N_2660,N_2535,N_2414);
and U2661 (N_2661,N_2584,N_2499);
or U2662 (N_2662,N_2518,N_2474);
nand U2663 (N_2663,N_2552,N_2433);
nor U2664 (N_2664,N_2481,N_2565);
nor U2665 (N_2665,N_2513,N_2497);
nand U2666 (N_2666,N_2483,N_2598);
or U2667 (N_2667,N_2557,N_2403);
or U2668 (N_2668,N_2484,N_2525);
xor U2669 (N_2669,N_2405,N_2444);
nor U2670 (N_2670,N_2577,N_2590);
or U2671 (N_2671,N_2510,N_2410);
or U2672 (N_2672,N_2402,N_2428);
nand U2673 (N_2673,N_2555,N_2442);
nand U2674 (N_2674,N_2574,N_2579);
or U2675 (N_2675,N_2477,N_2571);
or U2676 (N_2676,N_2521,N_2546);
nor U2677 (N_2677,N_2493,N_2491);
nor U2678 (N_2678,N_2487,N_2517);
or U2679 (N_2679,N_2406,N_2423);
or U2680 (N_2680,N_2463,N_2416);
or U2681 (N_2681,N_2475,N_2589);
or U2682 (N_2682,N_2512,N_2453);
nand U2683 (N_2683,N_2486,N_2508);
nor U2684 (N_2684,N_2505,N_2545);
nor U2685 (N_2685,N_2567,N_2450);
or U2686 (N_2686,N_2408,N_2570);
or U2687 (N_2687,N_2413,N_2404);
nand U2688 (N_2688,N_2436,N_2421);
or U2689 (N_2689,N_2543,N_2526);
nor U2690 (N_2690,N_2568,N_2514);
and U2691 (N_2691,N_2415,N_2503);
or U2692 (N_2692,N_2504,N_2485);
nor U2693 (N_2693,N_2542,N_2412);
nand U2694 (N_2694,N_2585,N_2536);
and U2695 (N_2695,N_2456,N_2432);
xnor U2696 (N_2696,N_2591,N_2507);
nand U2697 (N_2697,N_2506,N_2419);
and U2698 (N_2698,N_2473,N_2478);
and U2699 (N_2699,N_2458,N_2509);
nor U2700 (N_2700,N_2452,N_2404);
or U2701 (N_2701,N_2507,N_2582);
nand U2702 (N_2702,N_2472,N_2552);
or U2703 (N_2703,N_2487,N_2489);
or U2704 (N_2704,N_2583,N_2421);
or U2705 (N_2705,N_2441,N_2532);
nand U2706 (N_2706,N_2425,N_2556);
nor U2707 (N_2707,N_2488,N_2472);
and U2708 (N_2708,N_2437,N_2482);
and U2709 (N_2709,N_2543,N_2535);
nand U2710 (N_2710,N_2502,N_2524);
or U2711 (N_2711,N_2415,N_2547);
and U2712 (N_2712,N_2523,N_2421);
nand U2713 (N_2713,N_2504,N_2589);
nand U2714 (N_2714,N_2470,N_2433);
nand U2715 (N_2715,N_2427,N_2564);
nor U2716 (N_2716,N_2406,N_2564);
and U2717 (N_2717,N_2532,N_2563);
and U2718 (N_2718,N_2477,N_2508);
nand U2719 (N_2719,N_2513,N_2573);
nand U2720 (N_2720,N_2462,N_2504);
and U2721 (N_2721,N_2458,N_2405);
nand U2722 (N_2722,N_2423,N_2415);
nand U2723 (N_2723,N_2440,N_2560);
nor U2724 (N_2724,N_2534,N_2524);
or U2725 (N_2725,N_2483,N_2475);
or U2726 (N_2726,N_2531,N_2538);
nand U2727 (N_2727,N_2521,N_2518);
nand U2728 (N_2728,N_2548,N_2594);
nand U2729 (N_2729,N_2511,N_2534);
and U2730 (N_2730,N_2480,N_2403);
and U2731 (N_2731,N_2574,N_2555);
and U2732 (N_2732,N_2558,N_2562);
xnor U2733 (N_2733,N_2428,N_2418);
or U2734 (N_2734,N_2427,N_2408);
and U2735 (N_2735,N_2512,N_2598);
nor U2736 (N_2736,N_2408,N_2514);
or U2737 (N_2737,N_2473,N_2444);
nand U2738 (N_2738,N_2485,N_2571);
and U2739 (N_2739,N_2401,N_2543);
nor U2740 (N_2740,N_2429,N_2563);
nand U2741 (N_2741,N_2420,N_2400);
nand U2742 (N_2742,N_2533,N_2429);
or U2743 (N_2743,N_2494,N_2521);
nor U2744 (N_2744,N_2464,N_2536);
and U2745 (N_2745,N_2517,N_2510);
nand U2746 (N_2746,N_2467,N_2595);
or U2747 (N_2747,N_2594,N_2460);
nand U2748 (N_2748,N_2518,N_2544);
nand U2749 (N_2749,N_2473,N_2479);
or U2750 (N_2750,N_2504,N_2415);
nor U2751 (N_2751,N_2586,N_2413);
and U2752 (N_2752,N_2491,N_2433);
nor U2753 (N_2753,N_2541,N_2526);
or U2754 (N_2754,N_2586,N_2532);
nor U2755 (N_2755,N_2598,N_2450);
nor U2756 (N_2756,N_2519,N_2496);
nand U2757 (N_2757,N_2569,N_2564);
or U2758 (N_2758,N_2568,N_2545);
nor U2759 (N_2759,N_2508,N_2575);
nand U2760 (N_2760,N_2416,N_2477);
and U2761 (N_2761,N_2494,N_2413);
nor U2762 (N_2762,N_2484,N_2435);
nand U2763 (N_2763,N_2417,N_2590);
nand U2764 (N_2764,N_2559,N_2528);
and U2765 (N_2765,N_2487,N_2587);
and U2766 (N_2766,N_2556,N_2509);
or U2767 (N_2767,N_2461,N_2572);
and U2768 (N_2768,N_2434,N_2587);
nor U2769 (N_2769,N_2422,N_2406);
nor U2770 (N_2770,N_2481,N_2452);
nor U2771 (N_2771,N_2423,N_2510);
nand U2772 (N_2772,N_2558,N_2507);
xnor U2773 (N_2773,N_2513,N_2491);
nor U2774 (N_2774,N_2582,N_2414);
and U2775 (N_2775,N_2484,N_2477);
or U2776 (N_2776,N_2584,N_2445);
and U2777 (N_2777,N_2454,N_2591);
nand U2778 (N_2778,N_2514,N_2414);
nand U2779 (N_2779,N_2439,N_2554);
and U2780 (N_2780,N_2551,N_2489);
nor U2781 (N_2781,N_2472,N_2590);
or U2782 (N_2782,N_2547,N_2445);
or U2783 (N_2783,N_2406,N_2424);
and U2784 (N_2784,N_2569,N_2507);
nor U2785 (N_2785,N_2478,N_2598);
nand U2786 (N_2786,N_2505,N_2482);
or U2787 (N_2787,N_2437,N_2546);
and U2788 (N_2788,N_2531,N_2461);
or U2789 (N_2789,N_2422,N_2577);
and U2790 (N_2790,N_2590,N_2588);
nor U2791 (N_2791,N_2533,N_2463);
nand U2792 (N_2792,N_2435,N_2439);
and U2793 (N_2793,N_2571,N_2564);
or U2794 (N_2794,N_2544,N_2598);
nand U2795 (N_2795,N_2430,N_2569);
nor U2796 (N_2796,N_2592,N_2446);
and U2797 (N_2797,N_2534,N_2489);
and U2798 (N_2798,N_2496,N_2468);
nor U2799 (N_2799,N_2499,N_2471);
nand U2800 (N_2800,N_2672,N_2742);
or U2801 (N_2801,N_2780,N_2765);
or U2802 (N_2802,N_2653,N_2796);
and U2803 (N_2803,N_2723,N_2706);
nor U2804 (N_2804,N_2633,N_2603);
xor U2805 (N_2805,N_2762,N_2638);
nor U2806 (N_2806,N_2727,N_2641);
or U2807 (N_2807,N_2769,N_2629);
nor U2808 (N_2808,N_2715,N_2702);
nor U2809 (N_2809,N_2790,N_2787);
nor U2810 (N_2810,N_2660,N_2726);
and U2811 (N_2811,N_2754,N_2690);
and U2812 (N_2812,N_2652,N_2609);
nor U2813 (N_2813,N_2642,N_2650);
nand U2814 (N_2814,N_2788,N_2620);
or U2815 (N_2815,N_2774,N_2758);
nand U2816 (N_2816,N_2680,N_2608);
nor U2817 (N_2817,N_2734,N_2781);
nor U2818 (N_2818,N_2685,N_2744);
nor U2819 (N_2819,N_2622,N_2699);
or U2820 (N_2820,N_2729,N_2634);
and U2821 (N_2821,N_2683,N_2616);
or U2822 (N_2822,N_2659,N_2746);
nor U2823 (N_2823,N_2691,N_2631);
nand U2824 (N_2824,N_2752,N_2669);
or U2825 (N_2825,N_2719,N_2768);
nand U2826 (N_2826,N_2646,N_2736);
and U2827 (N_2827,N_2731,N_2645);
and U2828 (N_2828,N_2654,N_2604);
nor U2829 (N_2829,N_2751,N_2770);
xor U2830 (N_2830,N_2738,N_2610);
nand U2831 (N_2831,N_2735,N_2764);
nand U2832 (N_2832,N_2675,N_2643);
nand U2833 (N_2833,N_2743,N_2786);
nor U2834 (N_2834,N_2692,N_2748);
nand U2835 (N_2835,N_2623,N_2624);
nor U2836 (N_2836,N_2714,N_2625);
and U2837 (N_2837,N_2783,N_2655);
nand U2838 (N_2838,N_2741,N_2674);
and U2839 (N_2839,N_2637,N_2795);
and U2840 (N_2840,N_2640,N_2798);
or U2841 (N_2841,N_2757,N_2737);
nand U2842 (N_2842,N_2785,N_2662);
or U2843 (N_2843,N_2677,N_2724);
nand U2844 (N_2844,N_2772,N_2722);
nor U2845 (N_2845,N_2693,N_2750);
or U2846 (N_2846,N_2763,N_2687);
nand U2847 (N_2847,N_2618,N_2639);
and U2848 (N_2848,N_2688,N_2651);
nor U2849 (N_2849,N_2766,N_2767);
nand U2850 (N_2850,N_2739,N_2635);
nand U2851 (N_2851,N_2612,N_2728);
nor U2852 (N_2852,N_2730,N_2713);
or U2853 (N_2853,N_2761,N_2656);
nand U2854 (N_2854,N_2665,N_2601);
nor U2855 (N_2855,N_2753,N_2777);
nand U2856 (N_2856,N_2686,N_2708);
and U2857 (N_2857,N_2740,N_2789);
and U2858 (N_2858,N_2695,N_2689);
nor U2859 (N_2859,N_2681,N_2710);
or U2860 (N_2860,N_2626,N_2600);
and U2861 (N_2861,N_2602,N_2716);
nor U2862 (N_2862,N_2718,N_2791);
or U2863 (N_2863,N_2605,N_2663);
xor U2864 (N_2864,N_2679,N_2661);
and U2865 (N_2865,N_2648,N_2771);
nor U2866 (N_2866,N_2614,N_2676);
or U2867 (N_2867,N_2749,N_2696);
nand U2868 (N_2868,N_2760,N_2755);
and U2869 (N_2869,N_2632,N_2700);
nor U2870 (N_2870,N_2704,N_2621);
or U2871 (N_2871,N_2615,N_2712);
nor U2872 (N_2872,N_2636,N_2773);
xor U2873 (N_2873,N_2707,N_2611);
nor U2874 (N_2874,N_2792,N_2647);
nand U2875 (N_2875,N_2649,N_2720);
nand U2876 (N_2876,N_2698,N_2671);
nand U2877 (N_2877,N_2619,N_2617);
nor U2878 (N_2878,N_2779,N_2775);
or U2879 (N_2879,N_2799,N_2747);
nand U2880 (N_2880,N_2705,N_2670);
xor U2881 (N_2881,N_2782,N_2666);
nand U2882 (N_2882,N_2733,N_2756);
nand U2883 (N_2883,N_2664,N_2682);
or U2884 (N_2884,N_2776,N_2703);
or U2885 (N_2885,N_2709,N_2717);
and U2886 (N_2886,N_2667,N_2784);
and U2887 (N_2887,N_2628,N_2701);
nor U2888 (N_2888,N_2627,N_2797);
nor U2889 (N_2889,N_2711,N_2630);
and U2890 (N_2890,N_2606,N_2668);
xnor U2891 (N_2891,N_2673,N_2678);
nand U2892 (N_2892,N_2657,N_2793);
nor U2893 (N_2893,N_2697,N_2607);
nor U2894 (N_2894,N_2778,N_2658);
nand U2895 (N_2895,N_2644,N_2725);
nor U2896 (N_2896,N_2745,N_2684);
and U2897 (N_2897,N_2721,N_2732);
nor U2898 (N_2898,N_2759,N_2794);
nand U2899 (N_2899,N_2613,N_2694);
nor U2900 (N_2900,N_2700,N_2721);
nor U2901 (N_2901,N_2661,N_2639);
nand U2902 (N_2902,N_2647,N_2699);
nand U2903 (N_2903,N_2712,N_2693);
or U2904 (N_2904,N_2769,N_2603);
and U2905 (N_2905,N_2601,N_2796);
and U2906 (N_2906,N_2671,N_2626);
nand U2907 (N_2907,N_2708,N_2746);
or U2908 (N_2908,N_2697,N_2675);
or U2909 (N_2909,N_2702,N_2632);
nand U2910 (N_2910,N_2724,N_2750);
or U2911 (N_2911,N_2612,N_2719);
nor U2912 (N_2912,N_2708,N_2719);
nand U2913 (N_2913,N_2666,N_2691);
nor U2914 (N_2914,N_2747,N_2684);
and U2915 (N_2915,N_2602,N_2787);
and U2916 (N_2916,N_2699,N_2775);
and U2917 (N_2917,N_2619,N_2768);
nand U2918 (N_2918,N_2787,N_2726);
nor U2919 (N_2919,N_2702,N_2627);
nor U2920 (N_2920,N_2687,N_2674);
or U2921 (N_2921,N_2724,N_2774);
or U2922 (N_2922,N_2775,N_2722);
or U2923 (N_2923,N_2656,N_2615);
or U2924 (N_2924,N_2684,N_2754);
nand U2925 (N_2925,N_2659,N_2611);
nand U2926 (N_2926,N_2687,N_2622);
or U2927 (N_2927,N_2639,N_2671);
and U2928 (N_2928,N_2610,N_2605);
and U2929 (N_2929,N_2742,N_2629);
nand U2930 (N_2930,N_2764,N_2779);
nand U2931 (N_2931,N_2768,N_2631);
nand U2932 (N_2932,N_2672,N_2760);
nand U2933 (N_2933,N_2687,N_2659);
nand U2934 (N_2934,N_2604,N_2640);
nor U2935 (N_2935,N_2732,N_2786);
nand U2936 (N_2936,N_2791,N_2753);
nor U2937 (N_2937,N_2697,N_2677);
nor U2938 (N_2938,N_2693,N_2741);
nand U2939 (N_2939,N_2622,N_2728);
and U2940 (N_2940,N_2772,N_2715);
or U2941 (N_2941,N_2627,N_2694);
or U2942 (N_2942,N_2721,N_2657);
or U2943 (N_2943,N_2666,N_2628);
and U2944 (N_2944,N_2798,N_2679);
nor U2945 (N_2945,N_2710,N_2701);
or U2946 (N_2946,N_2788,N_2778);
or U2947 (N_2947,N_2682,N_2752);
or U2948 (N_2948,N_2793,N_2754);
or U2949 (N_2949,N_2772,N_2791);
nor U2950 (N_2950,N_2701,N_2754);
xnor U2951 (N_2951,N_2638,N_2777);
or U2952 (N_2952,N_2693,N_2767);
or U2953 (N_2953,N_2779,N_2681);
nor U2954 (N_2954,N_2623,N_2672);
nand U2955 (N_2955,N_2684,N_2691);
or U2956 (N_2956,N_2632,N_2623);
or U2957 (N_2957,N_2771,N_2755);
or U2958 (N_2958,N_2717,N_2726);
or U2959 (N_2959,N_2767,N_2607);
nand U2960 (N_2960,N_2798,N_2664);
or U2961 (N_2961,N_2638,N_2753);
nor U2962 (N_2962,N_2784,N_2651);
nor U2963 (N_2963,N_2669,N_2701);
nor U2964 (N_2964,N_2726,N_2714);
nor U2965 (N_2965,N_2706,N_2683);
nor U2966 (N_2966,N_2653,N_2652);
or U2967 (N_2967,N_2625,N_2671);
nor U2968 (N_2968,N_2702,N_2726);
and U2969 (N_2969,N_2666,N_2601);
or U2970 (N_2970,N_2604,N_2637);
or U2971 (N_2971,N_2730,N_2739);
nor U2972 (N_2972,N_2604,N_2765);
nor U2973 (N_2973,N_2620,N_2612);
or U2974 (N_2974,N_2736,N_2627);
xnor U2975 (N_2975,N_2608,N_2758);
and U2976 (N_2976,N_2715,N_2604);
nand U2977 (N_2977,N_2795,N_2658);
and U2978 (N_2978,N_2769,N_2602);
and U2979 (N_2979,N_2765,N_2692);
or U2980 (N_2980,N_2709,N_2767);
and U2981 (N_2981,N_2691,N_2603);
or U2982 (N_2982,N_2651,N_2661);
nor U2983 (N_2983,N_2743,N_2762);
and U2984 (N_2984,N_2769,N_2711);
nor U2985 (N_2985,N_2672,N_2605);
nand U2986 (N_2986,N_2676,N_2732);
nand U2987 (N_2987,N_2611,N_2603);
or U2988 (N_2988,N_2778,N_2708);
or U2989 (N_2989,N_2632,N_2728);
nand U2990 (N_2990,N_2702,N_2690);
or U2991 (N_2991,N_2662,N_2797);
or U2992 (N_2992,N_2795,N_2709);
nor U2993 (N_2993,N_2695,N_2781);
nand U2994 (N_2994,N_2661,N_2620);
or U2995 (N_2995,N_2636,N_2651);
nor U2996 (N_2996,N_2739,N_2648);
or U2997 (N_2997,N_2614,N_2765);
or U2998 (N_2998,N_2739,N_2777);
nor U2999 (N_2999,N_2603,N_2665);
nand U3000 (N_3000,N_2800,N_2854);
nor U3001 (N_3001,N_2868,N_2819);
or U3002 (N_3002,N_2812,N_2932);
nor U3003 (N_3003,N_2962,N_2897);
nor U3004 (N_3004,N_2990,N_2834);
nand U3005 (N_3005,N_2895,N_2810);
and U3006 (N_3006,N_2943,N_2956);
and U3007 (N_3007,N_2931,N_2978);
or U3008 (N_3008,N_2839,N_2910);
xor U3009 (N_3009,N_2824,N_2903);
and U3010 (N_3010,N_2808,N_2806);
nor U3011 (N_3011,N_2892,N_2933);
nand U3012 (N_3012,N_2885,N_2846);
nor U3013 (N_3013,N_2838,N_2882);
or U3014 (N_3014,N_2844,N_2878);
and U3015 (N_3015,N_2874,N_2862);
nand U3016 (N_3016,N_2803,N_2837);
xor U3017 (N_3017,N_2857,N_2909);
or U3018 (N_3018,N_2967,N_2983);
nor U3019 (N_3019,N_2993,N_2881);
nor U3020 (N_3020,N_2864,N_2900);
and U3021 (N_3021,N_2822,N_2984);
nand U3022 (N_3022,N_2826,N_2998);
nor U3023 (N_3023,N_2884,N_2996);
or U3024 (N_3024,N_2929,N_2893);
nand U3025 (N_3025,N_2814,N_2971);
and U3026 (N_3026,N_2977,N_2904);
and U3027 (N_3027,N_2914,N_2928);
nor U3028 (N_3028,N_2999,N_2825);
nor U3029 (N_3029,N_2924,N_2829);
nor U3030 (N_3030,N_2923,N_2994);
nand U3031 (N_3031,N_2859,N_2823);
and U3032 (N_3032,N_2852,N_2818);
nand U3033 (N_3033,N_2953,N_2888);
nand U3034 (N_3034,N_2902,N_2920);
and U3035 (N_3035,N_2847,N_2926);
and U3036 (N_3036,N_2957,N_2966);
nand U3037 (N_3037,N_2855,N_2841);
nor U3038 (N_3038,N_2991,N_2976);
nor U3039 (N_3039,N_2961,N_2916);
nand U3040 (N_3040,N_2908,N_2890);
nand U3041 (N_3041,N_2849,N_2905);
nor U3042 (N_3042,N_2913,N_2832);
nand U3043 (N_3043,N_2912,N_2907);
nor U3044 (N_3044,N_2981,N_2965);
nor U3045 (N_3045,N_2975,N_2873);
or U3046 (N_3046,N_2972,N_2937);
nor U3047 (N_3047,N_2860,N_2861);
or U3048 (N_3048,N_2948,N_2816);
nand U3049 (N_3049,N_2992,N_2987);
or U3050 (N_3050,N_2921,N_2807);
nor U3051 (N_3051,N_2946,N_2922);
and U3052 (N_3052,N_2830,N_2952);
nand U3053 (N_3053,N_2911,N_2982);
or U3054 (N_3054,N_2919,N_2872);
or U3055 (N_3055,N_2954,N_2896);
or U3056 (N_3056,N_2986,N_2968);
or U3057 (N_3057,N_2856,N_2809);
and U3058 (N_3058,N_2836,N_2831);
or U3059 (N_3059,N_2867,N_2970);
nand U3060 (N_3060,N_2886,N_2805);
nand U3061 (N_3061,N_2944,N_2883);
and U3062 (N_3062,N_2927,N_2955);
xor U3063 (N_3063,N_2817,N_2871);
or U3064 (N_3064,N_2821,N_2891);
xor U3065 (N_3065,N_2887,N_2945);
nand U3066 (N_3066,N_2877,N_2866);
and U3067 (N_3067,N_2833,N_2941);
nand U3068 (N_3068,N_2858,N_2845);
nand U3069 (N_3069,N_2827,N_2973);
xnor U3070 (N_3070,N_2942,N_2960);
nor U3071 (N_3071,N_2879,N_2876);
or U3072 (N_3072,N_2940,N_2917);
and U3073 (N_3073,N_2898,N_2947);
and U3074 (N_3074,N_2802,N_2915);
and U3075 (N_3075,N_2840,N_2951);
xor U3076 (N_3076,N_2801,N_2925);
or U3077 (N_3077,N_2848,N_2989);
nor U3078 (N_3078,N_2997,N_2930);
nand U3079 (N_3079,N_2901,N_2918);
nand U3080 (N_3080,N_2850,N_2851);
nand U3081 (N_3081,N_2985,N_2988);
or U3082 (N_3082,N_2980,N_2828);
nand U3083 (N_3083,N_2863,N_2870);
and U3084 (N_3084,N_2935,N_2969);
nand U3085 (N_3085,N_2815,N_2865);
nor U3086 (N_3086,N_2869,N_2889);
and U3087 (N_3087,N_2958,N_2842);
xnor U3088 (N_3088,N_2949,N_2995);
nor U3089 (N_3089,N_2899,N_2979);
nand U3090 (N_3090,N_2894,N_2880);
nand U3091 (N_3091,N_2875,N_2974);
xor U3092 (N_3092,N_2820,N_2938);
and U3093 (N_3093,N_2936,N_2963);
or U3094 (N_3094,N_2835,N_2964);
or U3095 (N_3095,N_2811,N_2959);
and U3096 (N_3096,N_2939,N_2934);
and U3097 (N_3097,N_2853,N_2906);
or U3098 (N_3098,N_2804,N_2813);
or U3099 (N_3099,N_2950,N_2843);
and U3100 (N_3100,N_2864,N_2920);
nand U3101 (N_3101,N_2944,N_2870);
nor U3102 (N_3102,N_2939,N_2991);
nand U3103 (N_3103,N_2853,N_2947);
nand U3104 (N_3104,N_2987,N_2806);
or U3105 (N_3105,N_2935,N_2922);
nand U3106 (N_3106,N_2867,N_2903);
nand U3107 (N_3107,N_2887,N_2991);
and U3108 (N_3108,N_2863,N_2878);
and U3109 (N_3109,N_2952,N_2818);
nor U3110 (N_3110,N_2805,N_2923);
nor U3111 (N_3111,N_2852,N_2841);
nor U3112 (N_3112,N_2963,N_2930);
and U3113 (N_3113,N_2819,N_2900);
nand U3114 (N_3114,N_2856,N_2824);
nor U3115 (N_3115,N_2934,N_2858);
nor U3116 (N_3116,N_2866,N_2833);
and U3117 (N_3117,N_2908,N_2954);
nor U3118 (N_3118,N_2820,N_2845);
nor U3119 (N_3119,N_2855,N_2920);
nand U3120 (N_3120,N_2831,N_2992);
or U3121 (N_3121,N_2994,N_2819);
nor U3122 (N_3122,N_2870,N_2820);
nand U3123 (N_3123,N_2992,N_2839);
nor U3124 (N_3124,N_2893,N_2978);
or U3125 (N_3125,N_2820,N_2918);
or U3126 (N_3126,N_2838,N_2962);
or U3127 (N_3127,N_2904,N_2829);
nand U3128 (N_3128,N_2853,N_2978);
or U3129 (N_3129,N_2817,N_2846);
and U3130 (N_3130,N_2907,N_2949);
or U3131 (N_3131,N_2807,N_2858);
nand U3132 (N_3132,N_2814,N_2975);
or U3133 (N_3133,N_2971,N_2939);
and U3134 (N_3134,N_2834,N_2937);
nand U3135 (N_3135,N_2815,N_2839);
nor U3136 (N_3136,N_2803,N_2978);
and U3137 (N_3137,N_2826,N_2952);
or U3138 (N_3138,N_2909,N_2918);
nor U3139 (N_3139,N_2804,N_2814);
or U3140 (N_3140,N_2826,N_2930);
nand U3141 (N_3141,N_2918,N_2900);
and U3142 (N_3142,N_2979,N_2964);
nor U3143 (N_3143,N_2903,N_2881);
nand U3144 (N_3144,N_2977,N_2802);
or U3145 (N_3145,N_2883,N_2956);
nand U3146 (N_3146,N_2945,N_2869);
nand U3147 (N_3147,N_2982,N_2976);
nand U3148 (N_3148,N_2862,N_2935);
nand U3149 (N_3149,N_2819,N_2917);
nand U3150 (N_3150,N_2910,N_2959);
nor U3151 (N_3151,N_2964,N_2865);
nor U3152 (N_3152,N_2983,N_2917);
nand U3153 (N_3153,N_2963,N_2851);
nor U3154 (N_3154,N_2882,N_2928);
nor U3155 (N_3155,N_2823,N_2990);
and U3156 (N_3156,N_2952,N_2814);
nand U3157 (N_3157,N_2814,N_2963);
or U3158 (N_3158,N_2841,N_2955);
and U3159 (N_3159,N_2966,N_2848);
and U3160 (N_3160,N_2957,N_2952);
nor U3161 (N_3161,N_2968,N_2823);
or U3162 (N_3162,N_2968,N_2992);
nand U3163 (N_3163,N_2883,N_2926);
and U3164 (N_3164,N_2933,N_2959);
nor U3165 (N_3165,N_2961,N_2912);
and U3166 (N_3166,N_2913,N_2930);
and U3167 (N_3167,N_2852,N_2942);
and U3168 (N_3168,N_2875,N_2827);
and U3169 (N_3169,N_2894,N_2914);
xor U3170 (N_3170,N_2829,N_2958);
and U3171 (N_3171,N_2802,N_2877);
nor U3172 (N_3172,N_2821,N_2881);
and U3173 (N_3173,N_2996,N_2861);
xor U3174 (N_3174,N_2830,N_2859);
and U3175 (N_3175,N_2978,N_2836);
or U3176 (N_3176,N_2846,N_2936);
nor U3177 (N_3177,N_2951,N_2847);
nand U3178 (N_3178,N_2881,N_2951);
and U3179 (N_3179,N_2942,N_2870);
nor U3180 (N_3180,N_2971,N_2934);
or U3181 (N_3181,N_2828,N_2956);
nor U3182 (N_3182,N_2846,N_2920);
nor U3183 (N_3183,N_2947,N_2966);
and U3184 (N_3184,N_2912,N_2891);
or U3185 (N_3185,N_2959,N_2940);
or U3186 (N_3186,N_2812,N_2909);
or U3187 (N_3187,N_2947,N_2857);
or U3188 (N_3188,N_2837,N_2925);
nand U3189 (N_3189,N_2842,N_2857);
nand U3190 (N_3190,N_2876,N_2944);
nor U3191 (N_3191,N_2931,N_2896);
or U3192 (N_3192,N_2978,N_2990);
and U3193 (N_3193,N_2927,N_2977);
and U3194 (N_3194,N_2854,N_2866);
and U3195 (N_3195,N_2897,N_2963);
and U3196 (N_3196,N_2808,N_2819);
and U3197 (N_3197,N_2900,N_2851);
and U3198 (N_3198,N_2954,N_2960);
nor U3199 (N_3199,N_2930,N_2848);
or U3200 (N_3200,N_3085,N_3158);
or U3201 (N_3201,N_3040,N_3015);
nor U3202 (N_3202,N_3136,N_3149);
and U3203 (N_3203,N_3076,N_3011);
and U3204 (N_3204,N_3027,N_3007);
and U3205 (N_3205,N_3053,N_3175);
nor U3206 (N_3206,N_3113,N_3020);
or U3207 (N_3207,N_3194,N_3168);
nand U3208 (N_3208,N_3097,N_3044);
or U3209 (N_3209,N_3024,N_3184);
or U3210 (N_3210,N_3073,N_3012);
nand U3211 (N_3211,N_3099,N_3045);
and U3212 (N_3212,N_3151,N_3019);
nor U3213 (N_3213,N_3051,N_3061);
nand U3214 (N_3214,N_3068,N_3057);
or U3215 (N_3215,N_3160,N_3058);
or U3216 (N_3216,N_3186,N_3060);
nand U3217 (N_3217,N_3088,N_3005);
nand U3218 (N_3218,N_3070,N_3188);
and U3219 (N_3219,N_3135,N_3112);
or U3220 (N_3220,N_3025,N_3154);
and U3221 (N_3221,N_3096,N_3091);
or U3222 (N_3222,N_3109,N_3187);
or U3223 (N_3223,N_3042,N_3167);
or U3224 (N_3224,N_3072,N_3115);
or U3225 (N_3225,N_3098,N_3043);
xnor U3226 (N_3226,N_3133,N_3089);
nor U3227 (N_3227,N_3153,N_3079);
nand U3228 (N_3228,N_3110,N_3146);
and U3229 (N_3229,N_3121,N_3004);
and U3230 (N_3230,N_3185,N_3084);
and U3231 (N_3231,N_3130,N_3124);
and U3232 (N_3232,N_3125,N_3148);
or U3233 (N_3233,N_3049,N_3018);
nor U3234 (N_3234,N_3196,N_3001);
or U3235 (N_3235,N_3156,N_3114);
and U3236 (N_3236,N_3122,N_3013);
xnor U3237 (N_3237,N_3180,N_3191);
nor U3238 (N_3238,N_3192,N_3034);
and U3239 (N_3239,N_3023,N_3086);
or U3240 (N_3240,N_3144,N_3128);
nand U3241 (N_3241,N_3108,N_3120);
and U3242 (N_3242,N_3172,N_3033);
nor U3243 (N_3243,N_3008,N_3032);
or U3244 (N_3244,N_3105,N_3095);
and U3245 (N_3245,N_3190,N_3164);
or U3246 (N_3246,N_3123,N_3117);
and U3247 (N_3247,N_3094,N_3028);
or U3248 (N_3248,N_3093,N_3181);
nor U3249 (N_3249,N_3179,N_3056);
or U3250 (N_3250,N_3141,N_3157);
nand U3251 (N_3251,N_3082,N_3118);
nand U3252 (N_3252,N_3116,N_3003);
nand U3253 (N_3253,N_3171,N_3131);
or U3254 (N_3254,N_3183,N_3074);
nand U3255 (N_3255,N_3195,N_3147);
or U3256 (N_3256,N_3126,N_3129);
nor U3257 (N_3257,N_3047,N_3170);
nand U3258 (N_3258,N_3055,N_3132);
xor U3259 (N_3259,N_3006,N_3162);
or U3260 (N_3260,N_3016,N_3002);
or U3261 (N_3261,N_3065,N_3026);
nor U3262 (N_3262,N_3041,N_3077);
or U3263 (N_3263,N_3182,N_3059);
nand U3264 (N_3264,N_3163,N_3197);
or U3265 (N_3265,N_3039,N_3062);
nor U3266 (N_3266,N_3067,N_3174);
nor U3267 (N_3267,N_3199,N_3021);
and U3268 (N_3268,N_3048,N_3176);
nand U3269 (N_3269,N_3193,N_3106);
and U3270 (N_3270,N_3038,N_3177);
nor U3271 (N_3271,N_3155,N_3165);
nand U3272 (N_3272,N_3143,N_3031);
or U3273 (N_3273,N_3142,N_3107);
or U3274 (N_3274,N_3104,N_3134);
nand U3275 (N_3275,N_3063,N_3101);
or U3276 (N_3276,N_3078,N_3102);
or U3277 (N_3277,N_3010,N_3198);
xor U3278 (N_3278,N_3046,N_3119);
nand U3279 (N_3279,N_3140,N_3111);
nor U3280 (N_3280,N_3050,N_3159);
nor U3281 (N_3281,N_3137,N_3000);
nand U3282 (N_3282,N_3087,N_3009);
or U3283 (N_3283,N_3090,N_3127);
and U3284 (N_3284,N_3081,N_3139);
and U3285 (N_3285,N_3083,N_3036);
or U3286 (N_3286,N_3075,N_3173);
and U3287 (N_3287,N_3150,N_3152);
nand U3288 (N_3288,N_3069,N_3052);
and U3289 (N_3289,N_3035,N_3022);
nand U3290 (N_3290,N_3166,N_3169);
and U3291 (N_3291,N_3066,N_3029);
nand U3292 (N_3292,N_3054,N_3138);
nor U3293 (N_3293,N_3189,N_3080);
or U3294 (N_3294,N_3071,N_3014);
nor U3295 (N_3295,N_3017,N_3161);
and U3296 (N_3296,N_3145,N_3092);
or U3297 (N_3297,N_3064,N_3030);
and U3298 (N_3298,N_3178,N_3100);
nand U3299 (N_3299,N_3103,N_3037);
nand U3300 (N_3300,N_3072,N_3055);
nand U3301 (N_3301,N_3076,N_3063);
or U3302 (N_3302,N_3063,N_3112);
nor U3303 (N_3303,N_3040,N_3001);
and U3304 (N_3304,N_3027,N_3195);
or U3305 (N_3305,N_3166,N_3177);
nor U3306 (N_3306,N_3133,N_3021);
and U3307 (N_3307,N_3195,N_3155);
and U3308 (N_3308,N_3169,N_3010);
or U3309 (N_3309,N_3082,N_3112);
and U3310 (N_3310,N_3024,N_3047);
or U3311 (N_3311,N_3157,N_3029);
nor U3312 (N_3312,N_3168,N_3020);
and U3313 (N_3313,N_3072,N_3060);
nor U3314 (N_3314,N_3155,N_3137);
and U3315 (N_3315,N_3002,N_3114);
nand U3316 (N_3316,N_3187,N_3146);
nor U3317 (N_3317,N_3161,N_3195);
and U3318 (N_3318,N_3060,N_3035);
and U3319 (N_3319,N_3121,N_3006);
nand U3320 (N_3320,N_3071,N_3199);
nor U3321 (N_3321,N_3114,N_3003);
nand U3322 (N_3322,N_3056,N_3082);
and U3323 (N_3323,N_3180,N_3006);
or U3324 (N_3324,N_3112,N_3111);
and U3325 (N_3325,N_3080,N_3156);
and U3326 (N_3326,N_3115,N_3103);
nor U3327 (N_3327,N_3037,N_3126);
and U3328 (N_3328,N_3149,N_3010);
nor U3329 (N_3329,N_3098,N_3069);
and U3330 (N_3330,N_3074,N_3086);
nand U3331 (N_3331,N_3012,N_3050);
nand U3332 (N_3332,N_3148,N_3181);
nand U3333 (N_3333,N_3039,N_3175);
or U3334 (N_3334,N_3130,N_3114);
nor U3335 (N_3335,N_3158,N_3155);
nand U3336 (N_3336,N_3006,N_3181);
or U3337 (N_3337,N_3052,N_3064);
or U3338 (N_3338,N_3007,N_3091);
or U3339 (N_3339,N_3041,N_3127);
or U3340 (N_3340,N_3035,N_3020);
or U3341 (N_3341,N_3168,N_3047);
and U3342 (N_3342,N_3075,N_3132);
nor U3343 (N_3343,N_3117,N_3084);
nor U3344 (N_3344,N_3086,N_3114);
or U3345 (N_3345,N_3092,N_3076);
nand U3346 (N_3346,N_3121,N_3051);
nand U3347 (N_3347,N_3014,N_3133);
and U3348 (N_3348,N_3045,N_3040);
or U3349 (N_3349,N_3045,N_3190);
or U3350 (N_3350,N_3193,N_3090);
or U3351 (N_3351,N_3133,N_3082);
nor U3352 (N_3352,N_3102,N_3070);
nand U3353 (N_3353,N_3026,N_3171);
nand U3354 (N_3354,N_3044,N_3100);
nor U3355 (N_3355,N_3067,N_3135);
nor U3356 (N_3356,N_3155,N_3045);
nand U3357 (N_3357,N_3021,N_3093);
nor U3358 (N_3358,N_3073,N_3122);
and U3359 (N_3359,N_3135,N_3097);
or U3360 (N_3360,N_3078,N_3117);
nand U3361 (N_3361,N_3014,N_3162);
nor U3362 (N_3362,N_3075,N_3083);
nand U3363 (N_3363,N_3133,N_3137);
and U3364 (N_3364,N_3035,N_3151);
and U3365 (N_3365,N_3158,N_3172);
or U3366 (N_3366,N_3124,N_3051);
or U3367 (N_3367,N_3063,N_3092);
or U3368 (N_3368,N_3068,N_3188);
nand U3369 (N_3369,N_3147,N_3114);
nand U3370 (N_3370,N_3024,N_3100);
and U3371 (N_3371,N_3155,N_3199);
and U3372 (N_3372,N_3148,N_3011);
nand U3373 (N_3373,N_3067,N_3171);
nor U3374 (N_3374,N_3137,N_3080);
nor U3375 (N_3375,N_3164,N_3107);
xor U3376 (N_3376,N_3114,N_3199);
or U3377 (N_3377,N_3065,N_3111);
nand U3378 (N_3378,N_3090,N_3047);
and U3379 (N_3379,N_3124,N_3040);
or U3380 (N_3380,N_3036,N_3016);
xor U3381 (N_3381,N_3095,N_3121);
nor U3382 (N_3382,N_3004,N_3192);
nor U3383 (N_3383,N_3045,N_3197);
or U3384 (N_3384,N_3061,N_3094);
and U3385 (N_3385,N_3062,N_3000);
and U3386 (N_3386,N_3129,N_3120);
and U3387 (N_3387,N_3084,N_3100);
and U3388 (N_3388,N_3075,N_3095);
nand U3389 (N_3389,N_3107,N_3175);
xnor U3390 (N_3390,N_3104,N_3103);
nand U3391 (N_3391,N_3029,N_3114);
nor U3392 (N_3392,N_3033,N_3015);
or U3393 (N_3393,N_3133,N_3062);
or U3394 (N_3394,N_3046,N_3042);
or U3395 (N_3395,N_3005,N_3182);
nand U3396 (N_3396,N_3021,N_3103);
nand U3397 (N_3397,N_3062,N_3090);
or U3398 (N_3398,N_3011,N_3123);
nor U3399 (N_3399,N_3036,N_3140);
and U3400 (N_3400,N_3371,N_3347);
or U3401 (N_3401,N_3291,N_3246);
or U3402 (N_3402,N_3212,N_3234);
nor U3403 (N_3403,N_3351,N_3383);
nor U3404 (N_3404,N_3217,N_3397);
and U3405 (N_3405,N_3261,N_3337);
or U3406 (N_3406,N_3319,N_3238);
nand U3407 (N_3407,N_3381,N_3267);
nand U3408 (N_3408,N_3262,N_3331);
or U3409 (N_3409,N_3244,N_3318);
nand U3410 (N_3410,N_3227,N_3209);
or U3411 (N_3411,N_3226,N_3256);
nor U3412 (N_3412,N_3210,N_3270);
nand U3413 (N_3413,N_3392,N_3286);
and U3414 (N_3414,N_3251,N_3295);
and U3415 (N_3415,N_3394,N_3367);
xnor U3416 (N_3416,N_3354,N_3340);
nor U3417 (N_3417,N_3206,N_3399);
and U3418 (N_3418,N_3384,N_3203);
or U3419 (N_3419,N_3249,N_3366);
or U3420 (N_3420,N_3283,N_3219);
or U3421 (N_3421,N_3271,N_3306);
or U3422 (N_3422,N_3250,N_3382);
nand U3423 (N_3423,N_3326,N_3221);
nor U3424 (N_3424,N_3360,N_3298);
or U3425 (N_3425,N_3229,N_3235);
or U3426 (N_3426,N_3315,N_3330);
or U3427 (N_3427,N_3390,N_3302);
or U3428 (N_3428,N_3204,N_3387);
nand U3429 (N_3429,N_3274,N_3389);
nor U3430 (N_3430,N_3328,N_3355);
nor U3431 (N_3431,N_3290,N_3338);
and U3432 (N_3432,N_3325,N_3341);
or U3433 (N_3433,N_3281,N_3211);
and U3434 (N_3434,N_3259,N_3314);
nor U3435 (N_3435,N_3264,N_3329);
and U3436 (N_3436,N_3357,N_3300);
and U3437 (N_3437,N_3398,N_3254);
and U3438 (N_3438,N_3363,N_3265);
xor U3439 (N_3439,N_3385,N_3202);
nor U3440 (N_3440,N_3359,N_3245);
nand U3441 (N_3441,N_3370,N_3232);
and U3442 (N_3442,N_3241,N_3247);
and U3443 (N_3443,N_3278,N_3207);
or U3444 (N_3444,N_3258,N_3374);
nor U3445 (N_3445,N_3335,N_3368);
nor U3446 (N_3446,N_3301,N_3252);
nor U3447 (N_3447,N_3242,N_3350);
nand U3448 (N_3448,N_3375,N_3324);
nand U3449 (N_3449,N_3343,N_3276);
nor U3450 (N_3450,N_3280,N_3218);
nand U3451 (N_3451,N_3275,N_3396);
or U3452 (N_3452,N_3386,N_3236);
and U3453 (N_3453,N_3346,N_3378);
or U3454 (N_3454,N_3200,N_3353);
nor U3455 (N_3455,N_3284,N_3323);
nor U3456 (N_3456,N_3316,N_3214);
and U3457 (N_3457,N_3327,N_3379);
nand U3458 (N_3458,N_3289,N_3208);
or U3459 (N_3459,N_3233,N_3294);
nand U3460 (N_3460,N_3313,N_3395);
and U3461 (N_3461,N_3239,N_3213);
and U3462 (N_3462,N_3305,N_3272);
nand U3463 (N_3463,N_3237,N_3266);
and U3464 (N_3464,N_3255,N_3260);
and U3465 (N_3465,N_3348,N_3273);
nand U3466 (N_3466,N_3321,N_3356);
nand U3467 (N_3467,N_3344,N_3352);
and U3468 (N_3468,N_3308,N_3339);
nor U3469 (N_3469,N_3287,N_3393);
and U3470 (N_3470,N_3345,N_3228);
and U3471 (N_3471,N_3230,N_3277);
or U3472 (N_3472,N_3342,N_3248);
nand U3473 (N_3473,N_3369,N_3225);
xnor U3474 (N_3474,N_3320,N_3380);
or U3475 (N_3475,N_3268,N_3332);
or U3476 (N_3476,N_3373,N_3358);
or U3477 (N_3477,N_3365,N_3362);
nand U3478 (N_3478,N_3224,N_3307);
xor U3479 (N_3479,N_3322,N_3388);
and U3480 (N_3480,N_3288,N_3223);
nand U3481 (N_3481,N_3377,N_3310);
and U3482 (N_3482,N_3304,N_3231);
nor U3483 (N_3483,N_3296,N_3372);
nor U3484 (N_3484,N_3349,N_3333);
nor U3485 (N_3485,N_3336,N_3312);
or U3486 (N_3486,N_3303,N_3269);
or U3487 (N_3487,N_3334,N_3257);
and U3488 (N_3488,N_3222,N_3285);
nor U3489 (N_3489,N_3279,N_3361);
or U3490 (N_3490,N_3253,N_3216);
or U3491 (N_3491,N_3220,N_3243);
or U3492 (N_3492,N_3311,N_3263);
nor U3493 (N_3493,N_3317,N_3205);
and U3494 (N_3494,N_3309,N_3376);
nor U3495 (N_3495,N_3240,N_3293);
or U3496 (N_3496,N_3282,N_3364);
or U3497 (N_3497,N_3299,N_3292);
or U3498 (N_3498,N_3215,N_3391);
and U3499 (N_3499,N_3297,N_3201);
and U3500 (N_3500,N_3238,N_3292);
nand U3501 (N_3501,N_3311,N_3307);
and U3502 (N_3502,N_3383,N_3326);
or U3503 (N_3503,N_3331,N_3265);
or U3504 (N_3504,N_3214,N_3259);
nand U3505 (N_3505,N_3398,N_3315);
nor U3506 (N_3506,N_3263,N_3275);
or U3507 (N_3507,N_3295,N_3377);
and U3508 (N_3508,N_3300,N_3289);
and U3509 (N_3509,N_3307,N_3329);
nor U3510 (N_3510,N_3279,N_3357);
nor U3511 (N_3511,N_3243,N_3380);
nand U3512 (N_3512,N_3246,N_3335);
nand U3513 (N_3513,N_3229,N_3236);
nand U3514 (N_3514,N_3282,N_3369);
nor U3515 (N_3515,N_3351,N_3371);
nor U3516 (N_3516,N_3244,N_3307);
or U3517 (N_3517,N_3201,N_3396);
or U3518 (N_3518,N_3343,N_3285);
nand U3519 (N_3519,N_3222,N_3388);
or U3520 (N_3520,N_3265,N_3234);
nor U3521 (N_3521,N_3363,N_3213);
nand U3522 (N_3522,N_3368,N_3339);
or U3523 (N_3523,N_3294,N_3246);
nand U3524 (N_3524,N_3235,N_3336);
nand U3525 (N_3525,N_3255,N_3380);
nand U3526 (N_3526,N_3322,N_3344);
or U3527 (N_3527,N_3324,N_3281);
and U3528 (N_3528,N_3209,N_3340);
xor U3529 (N_3529,N_3218,N_3328);
nand U3530 (N_3530,N_3290,N_3336);
and U3531 (N_3531,N_3216,N_3245);
nand U3532 (N_3532,N_3276,N_3365);
nand U3533 (N_3533,N_3220,N_3344);
nand U3534 (N_3534,N_3300,N_3200);
nor U3535 (N_3535,N_3249,N_3374);
nand U3536 (N_3536,N_3200,N_3294);
nor U3537 (N_3537,N_3267,N_3373);
or U3538 (N_3538,N_3331,N_3297);
nand U3539 (N_3539,N_3393,N_3318);
and U3540 (N_3540,N_3227,N_3330);
or U3541 (N_3541,N_3241,N_3220);
nor U3542 (N_3542,N_3234,N_3336);
and U3543 (N_3543,N_3329,N_3388);
or U3544 (N_3544,N_3343,N_3338);
nor U3545 (N_3545,N_3228,N_3391);
nand U3546 (N_3546,N_3290,N_3348);
and U3547 (N_3547,N_3290,N_3240);
and U3548 (N_3548,N_3337,N_3363);
or U3549 (N_3549,N_3383,N_3250);
or U3550 (N_3550,N_3365,N_3311);
and U3551 (N_3551,N_3290,N_3215);
and U3552 (N_3552,N_3389,N_3369);
and U3553 (N_3553,N_3218,N_3376);
and U3554 (N_3554,N_3395,N_3275);
nor U3555 (N_3555,N_3363,N_3350);
or U3556 (N_3556,N_3344,N_3251);
nand U3557 (N_3557,N_3210,N_3297);
or U3558 (N_3558,N_3308,N_3338);
or U3559 (N_3559,N_3287,N_3300);
nand U3560 (N_3560,N_3367,N_3264);
and U3561 (N_3561,N_3250,N_3374);
and U3562 (N_3562,N_3205,N_3251);
nor U3563 (N_3563,N_3314,N_3388);
nor U3564 (N_3564,N_3360,N_3304);
nand U3565 (N_3565,N_3208,N_3358);
nand U3566 (N_3566,N_3384,N_3392);
and U3567 (N_3567,N_3308,N_3270);
nand U3568 (N_3568,N_3238,N_3353);
nor U3569 (N_3569,N_3339,N_3372);
or U3570 (N_3570,N_3230,N_3360);
nor U3571 (N_3571,N_3338,N_3332);
nor U3572 (N_3572,N_3296,N_3266);
or U3573 (N_3573,N_3249,N_3312);
or U3574 (N_3574,N_3370,N_3218);
or U3575 (N_3575,N_3289,N_3266);
and U3576 (N_3576,N_3230,N_3383);
or U3577 (N_3577,N_3264,N_3363);
xnor U3578 (N_3578,N_3280,N_3345);
nand U3579 (N_3579,N_3313,N_3251);
and U3580 (N_3580,N_3243,N_3244);
and U3581 (N_3581,N_3381,N_3295);
nand U3582 (N_3582,N_3214,N_3343);
nor U3583 (N_3583,N_3368,N_3312);
nor U3584 (N_3584,N_3256,N_3286);
nor U3585 (N_3585,N_3287,N_3357);
and U3586 (N_3586,N_3350,N_3348);
or U3587 (N_3587,N_3276,N_3312);
or U3588 (N_3588,N_3223,N_3209);
or U3589 (N_3589,N_3390,N_3292);
nand U3590 (N_3590,N_3226,N_3284);
nand U3591 (N_3591,N_3329,N_3311);
nand U3592 (N_3592,N_3368,N_3230);
and U3593 (N_3593,N_3290,N_3325);
or U3594 (N_3594,N_3377,N_3370);
nand U3595 (N_3595,N_3395,N_3316);
or U3596 (N_3596,N_3331,N_3216);
and U3597 (N_3597,N_3251,N_3353);
and U3598 (N_3598,N_3297,N_3225);
and U3599 (N_3599,N_3350,N_3281);
or U3600 (N_3600,N_3574,N_3590);
and U3601 (N_3601,N_3508,N_3511);
and U3602 (N_3602,N_3460,N_3415);
nand U3603 (N_3603,N_3483,N_3421);
and U3604 (N_3604,N_3403,N_3571);
or U3605 (N_3605,N_3587,N_3413);
nor U3606 (N_3606,N_3546,N_3539);
and U3607 (N_3607,N_3527,N_3420);
nand U3608 (N_3608,N_3585,N_3406);
xnor U3609 (N_3609,N_3432,N_3576);
xor U3610 (N_3610,N_3427,N_3561);
nor U3611 (N_3611,N_3497,N_3567);
or U3612 (N_3612,N_3437,N_3500);
nor U3613 (N_3613,N_3407,N_3534);
or U3614 (N_3614,N_3519,N_3402);
nor U3615 (N_3615,N_3468,N_3565);
nor U3616 (N_3616,N_3541,N_3502);
nor U3617 (N_3617,N_3471,N_3465);
and U3618 (N_3618,N_3419,N_3531);
nand U3619 (N_3619,N_3449,N_3487);
nand U3620 (N_3620,N_3481,N_3470);
nor U3621 (N_3621,N_3505,N_3532);
xor U3622 (N_3622,N_3488,N_3552);
nand U3623 (N_3623,N_3446,N_3447);
nand U3624 (N_3624,N_3451,N_3504);
nand U3625 (N_3625,N_3591,N_3463);
nand U3626 (N_3626,N_3443,N_3431);
nor U3627 (N_3627,N_3557,N_3551);
or U3628 (N_3628,N_3485,N_3526);
nor U3629 (N_3629,N_3475,N_3422);
or U3630 (N_3630,N_3401,N_3434);
or U3631 (N_3631,N_3423,N_3499);
xor U3632 (N_3632,N_3512,N_3575);
or U3633 (N_3633,N_3491,N_3582);
nor U3634 (N_3634,N_3495,N_3428);
nor U3635 (N_3635,N_3510,N_3518);
and U3636 (N_3636,N_3404,N_3572);
nand U3637 (N_3637,N_3472,N_3598);
and U3638 (N_3638,N_3545,N_3548);
and U3639 (N_3639,N_3515,N_3599);
nor U3640 (N_3640,N_3584,N_3452);
nor U3641 (N_3641,N_3445,N_3562);
and U3642 (N_3642,N_3412,N_3597);
or U3643 (N_3643,N_3558,N_3596);
nor U3644 (N_3644,N_3478,N_3528);
and U3645 (N_3645,N_3520,N_3569);
nor U3646 (N_3646,N_3408,N_3524);
nand U3647 (N_3647,N_3581,N_3442);
and U3648 (N_3648,N_3530,N_3554);
nor U3649 (N_3649,N_3486,N_3489);
and U3650 (N_3650,N_3564,N_3513);
or U3651 (N_3651,N_3514,N_3560);
or U3652 (N_3652,N_3456,N_3559);
and U3653 (N_3653,N_3547,N_3568);
and U3654 (N_3654,N_3540,N_3426);
or U3655 (N_3655,N_3493,N_3474);
or U3656 (N_3656,N_3523,N_3516);
nand U3657 (N_3657,N_3577,N_3461);
nand U3658 (N_3658,N_3553,N_3436);
xnor U3659 (N_3659,N_3570,N_3555);
and U3660 (N_3660,N_3424,N_3417);
nand U3661 (N_3661,N_3578,N_3476);
nand U3662 (N_3662,N_3464,N_3425);
and U3663 (N_3663,N_3457,N_3494);
or U3664 (N_3664,N_3498,N_3459);
nand U3665 (N_3665,N_3440,N_3586);
and U3666 (N_3666,N_3563,N_3537);
and U3667 (N_3667,N_3454,N_3579);
nor U3668 (N_3668,N_3430,N_3429);
nor U3669 (N_3669,N_3521,N_3550);
nor U3670 (N_3670,N_3477,N_3450);
nor U3671 (N_3671,N_3506,N_3593);
or U3672 (N_3672,N_3595,N_3544);
or U3673 (N_3673,N_3525,N_3543);
nor U3674 (N_3674,N_3411,N_3580);
and U3675 (N_3675,N_3480,N_3473);
or U3676 (N_3676,N_3503,N_3549);
xor U3677 (N_3677,N_3566,N_3400);
and U3678 (N_3678,N_3405,N_3509);
nor U3679 (N_3679,N_3453,N_3536);
nand U3680 (N_3680,N_3492,N_3441);
or U3681 (N_3681,N_3490,N_3458);
nand U3682 (N_3682,N_3588,N_3414);
and U3683 (N_3683,N_3529,N_3589);
nor U3684 (N_3684,N_3466,N_3416);
nand U3685 (N_3685,N_3467,N_3496);
and U3686 (N_3686,N_3583,N_3594);
or U3687 (N_3687,N_3517,N_3482);
nand U3688 (N_3688,N_3592,N_3439);
nor U3689 (N_3689,N_3479,N_3535);
nor U3690 (N_3690,N_3448,N_3507);
nor U3691 (N_3691,N_3435,N_3455);
or U3692 (N_3692,N_3501,N_3522);
and U3693 (N_3693,N_3484,N_3538);
nand U3694 (N_3694,N_3573,N_3469);
or U3695 (N_3695,N_3410,N_3556);
or U3696 (N_3696,N_3418,N_3438);
nand U3697 (N_3697,N_3462,N_3542);
or U3698 (N_3698,N_3533,N_3433);
nor U3699 (N_3699,N_3444,N_3409);
and U3700 (N_3700,N_3469,N_3594);
or U3701 (N_3701,N_3425,N_3514);
nand U3702 (N_3702,N_3541,N_3555);
and U3703 (N_3703,N_3462,N_3546);
nor U3704 (N_3704,N_3540,N_3579);
and U3705 (N_3705,N_3493,N_3447);
and U3706 (N_3706,N_3583,N_3587);
nor U3707 (N_3707,N_3483,N_3514);
and U3708 (N_3708,N_3426,N_3441);
nor U3709 (N_3709,N_3565,N_3431);
nor U3710 (N_3710,N_3442,N_3489);
nor U3711 (N_3711,N_3561,N_3581);
and U3712 (N_3712,N_3442,N_3476);
and U3713 (N_3713,N_3453,N_3532);
nand U3714 (N_3714,N_3505,N_3403);
or U3715 (N_3715,N_3513,N_3502);
and U3716 (N_3716,N_3496,N_3524);
and U3717 (N_3717,N_3472,N_3585);
and U3718 (N_3718,N_3458,N_3460);
or U3719 (N_3719,N_3591,N_3462);
or U3720 (N_3720,N_3464,N_3457);
xor U3721 (N_3721,N_3551,N_3585);
nor U3722 (N_3722,N_3557,N_3432);
nand U3723 (N_3723,N_3537,N_3531);
or U3724 (N_3724,N_3541,N_3532);
nand U3725 (N_3725,N_3529,N_3590);
or U3726 (N_3726,N_3576,N_3423);
nor U3727 (N_3727,N_3458,N_3594);
nor U3728 (N_3728,N_3509,N_3500);
and U3729 (N_3729,N_3581,N_3543);
nor U3730 (N_3730,N_3456,N_3479);
nand U3731 (N_3731,N_3500,N_3461);
nand U3732 (N_3732,N_3586,N_3507);
nand U3733 (N_3733,N_3521,N_3494);
and U3734 (N_3734,N_3418,N_3581);
nand U3735 (N_3735,N_3466,N_3595);
or U3736 (N_3736,N_3432,N_3595);
and U3737 (N_3737,N_3561,N_3573);
or U3738 (N_3738,N_3571,N_3547);
nor U3739 (N_3739,N_3592,N_3515);
and U3740 (N_3740,N_3411,N_3448);
nand U3741 (N_3741,N_3488,N_3417);
or U3742 (N_3742,N_3413,N_3518);
nand U3743 (N_3743,N_3530,N_3433);
nand U3744 (N_3744,N_3402,N_3468);
nand U3745 (N_3745,N_3514,N_3497);
or U3746 (N_3746,N_3575,N_3540);
or U3747 (N_3747,N_3518,N_3410);
and U3748 (N_3748,N_3538,N_3576);
or U3749 (N_3749,N_3574,N_3429);
nor U3750 (N_3750,N_3452,N_3577);
nand U3751 (N_3751,N_3497,N_3449);
nand U3752 (N_3752,N_3426,N_3566);
and U3753 (N_3753,N_3433,N_3540);
or U3754 (N_3754,N_3580,N_3414);
nor U3755 (N_3755,N_3478,N_3594);
nor U3756 (N_3756,N_3444,N_3453);
nor U3757 (N_3757,N_3480,N_3488);
nand U3758 (N_3758,N_3558,N_3584);
or U3759 (N_3759,N_3417,N_3588);
nor U3760 (N_3760,N_3400,N_3545);
and U3761 (N_3761,N_3482,N_3596);
and U3762 (N_3762,N_3534,N_3433);
nand U3763 (N_3763,N_3473,N_3582);
nor U3764 (N_3764,N_3499,N_3476);
nor U3765 (N_3765,N_3529,N_3472);
xor U3766 (N_3766,N_3405,N_3505);
nand U3767 (N_3767,N_3525,N_3470);
nor U3768 (N_3768,N_3428,N_3510);
nand U3769 (N_3769,N_3520,N_3413);
nor U3770 (N_3770,N_3501,N_3592);
or U3771 (N_3771,N_3443,N_3500);
and U3772 (N_3772,N_3509,N_3488);
xor U3773 (N_3773,N_3431,N_3464);
nor U3774 (N_3774,N_3437,N_3476);
nor U3775 (N_3775,N_3467,N_3465);
or U3776 (N_3776,N_3491,N_3520);
and U3777 (N_3777,N_3516,N_3519);
and U3778 (N_3778,N_3491,N_3457);
nor U3779 (N_3779,N_3461,N_3589);
nor U3780 (N_3780,N_3591,N_3465);
and U3781 (N_3781,N_3581,N_3556);
nand U3782 (N_3782,N_3451,N_3524);
nor U3783 (N_3783,N_3405,N_3569);
nand U3784 (N_3784,N_3542,N_3526);
and U3785 (N_3785,N_3441,N_3494);
nand U3786 (N_3786,N_3498,N_3509);
nand U3787 (N_3787,N_3426,N_3461);
or U3788 (N_3788,N_3417,N_3559);
and U3789 (N_3789,N_3506,N_3550);
and U3790 (N_3790,N_3484,N_3431);
and U3791 (N_3791,N_3471,N_3527);
or U3792 (N_3792,N_3565,N_3452);
and U3793 (N_3793,N_3587,N_3432);
nor U3794 (N_3794,N_3579,N_3510);
nand U3795 (N_3795,N_3445,N_3493);
nand U3796 (N_3796,N_3485,N_3511);
nor U3797 (N_3797,N_3531,N_3475);
or U3798 (N_3798,N_3570,N_3476);
nand U3799 (N_3799,N_3515,N_3554);
nor U3800 (N_3800,N_3696,N_3652);
nand U3801 (N_3801,N_3659,N_3779);
nand U3802 (N_3802,N_3604,N_3637);
or U3803 (N_3803,N_3754,N_3661);
or U3804 (N_3804,N_3697,N_3737);
or U3805 (N_3805,N_3683,N_3686);
or U3806 (N_3806,N_3681,N_3702);
and U3807 (N_3807,N_3773,N_3674);
xnor U3808 (N_3808,N_3717,N_3694);
nand U3809 (N_3809,N_3690,N_3768);
nand U3810 (N_3810,N_3763,N_3756);
or U3811 (N_3811,N_3735,N_3676);
nand U3812 (N_3812,N_3767,N_3720);
nand U3813 (N_3813,N_3700,N_3678);
or U3814 (N_3814,N_3682,N_3641);
nor U3815 (N_3815,N_3771,N_3626);
nor U3816 (N_3816,N_3660,N_3797);
nor U3817 (N_3817,N_3792,N_3786);
nand U3818 (N_3818,N_3671,N_3615);
or U3819 (N_3819,N_3772,N_3755);
nand U3820 (N_3820,N_3691,N_3625);
nor U3821 (N_3821,N_3669,N_3651);
or U3822 (N_3822,N_3627,N_3715);
nand U3823 (N_3823,N_3747,N_3736);
or U3824 (N_3824,N_3619,N_3733);
and U3825 (N_3825,N_3648,N_3611);
or U3826 (N_3826,N_3609,N_3710);
and U3827 (N_3827,N_3738,N_3628);
and U3828 (N_3828,N_3680,N_3643);
nand U3829 (N_3829,N_3750,N_3712);
or U3830 (N_3830,N_3752,N_3782);
or U3831 (N_3831,N_3788,N_3751);
nor U3832 (N_3832,N_3721,N_3638);
nand U3833 (N_3833,N_3618,N_3608);
nor U3834 (N_3834,N_3706,N_3603);
nand U3835 (N_3835,N_3708,N_3605);
and U3836 (N_3836,N_3718,N_3701);
and U3837 (N_3837,N_3666,N_3798);
nand U3838 (N_3838,N_3653,N_3724);
and U3839 (N_3839,N_3760,N_3654);
nor U3840 (N_3840,N_3732,N_3699);
and U3841 (N_3841,N_3663,N_3765);
and U3842 (N_3842,N_3727,N_3789);
nor U3843 (N_3843,N_3784,N_3650);
and U3844 (N_3844,N_3730,N_3734);
nor U3845 (N_3845,N_3793,N_3723);
and U3846 (N_3846,N_3725,N_3606);
or U3847 (N_3847,N_3799,N_3623);
nor U3848 (N_3848,N_3693,N_3631);
and U3849 (N_3849,N_3749,N_3764);
or U3850 (N_3850,N_3685,N_3649);
or U3851 (N_3851,N_3675,N_3688);
or U3852 (N_3852,N_3743,N_3741);
nand U3853 (N_3853,N_3729,N_3658);
nand U3854 (N_3854,N_3709,N_3769);
or U3855 (N_3855,N_3679,N_3778);
nor U3856 (N_3856,N_3642,N_3629);
nor U3857 (N_3857,N_3766,N_3672);
and U3858 (N_3858,N_3634,N_3647);
nand U3859 (N_3859,N_3639,N_3762);
nor U3860 (N_3860,N_3602,N_3600);
nor U3861 (N_3861,N_3781,N_3776);
nand U3862 (N_3862,N_3745,N_3705);
nand U3863 (N_3863,N_3746,N_3613);
and U3864 (N_3864,N_3722,N_3630);
and U3865 (N_3865,N_3795,N_3783);
or U3866 (N_3866,N_3757,N_3614);
nand U3867 (N_3867,N_3728,N_3684);
nor U3868 (N_3868,N_3713,N_3759);
nor U3869 (N_3869,N_3633,N_3689);
or U3870 (N_3870,N_3707,N_3644);
or U3871 (N_3871,N_3662,N_3753);
and U3872 (N_3872,N_3656,N_3677);
or U3873 (N_3873,N_3770,N_3740);
or U3874 (N_3874,N_3719,N_3714);
and U3875 (N_3875,N_3635,N_3610);
nor U3876 (N_3876,N_3617,N_3620);
nand U3877 (N_3877,N_3664,N_3731);
or U3878 (N_3878,N_3790,N_3687);
nand U3879 (N_3879,N_3622,N_3607);
and U3880 (N_3880,N_3621,N_3657);
and U3881 (N_3881,N_3796,N_3668);
nor U3882 (N_3882,N_3758,N_3698);
or U3883 (N_3883,N_3744,N_3670);
and U3884 (N_3884,N_3645,N_3640);
xnor U3885 (N_3885,N_3695,N_3791);
nor U3886 (N_3886,N_3612,N_3601);
nor U3887 (N_3887,N_3692,N_3726);
nor U3888 (N_3888,N_3716,N_3785);
nand U3889 (N_3889,N_3777,N_3632);
xnor U3890 (N_3890,N_3748,N_3761);
and U3891 (N_3891,N_3667,N_3616);
or U3892 (N_3892,N_3624,N_3646);
and U3893 (N_3893,N_3704,N_3636);
nor U3894 (N_3894,N_3787,N_3780);
and U3895 (N_3895,N_3711,N_3794);
or U3896 (N_3896,N_3739,N_3673);
or U3897 (N_3897,N_3742,N_3775);
nand U3898 (N_3898,N_3703,N_3665);
and U3899 (N_3899,N_3655,N_3774);
and U3900 (N_3900,N_3773,N_3648);
nor U3901 (N_3901,N_3622,N_3604);
and U3902 (N_3902,N_3626,N_3789);
or U3903 (N_3903,N_3797,N_3698);
or U3904 (N_3904,N_3657,N_3730);
nor U3905 (N_3905,N_3639,N_3758);
and U3906 (N_3906,N_3675,N_3782);
nand U3907 (N_3907,N_3670,N_3695);
and U3908 (N_3908,N_3777,N_3639);
nand U3909 (N_3909,N_3617,N_3602);
nand U3910 (N_3910,N_3655,N_3790);
and U3911 (N_3911,N_3778,N_3685);
nand U3912 (N_3912,N_3693,N_3633);
and U3913 (N_3913,N_3781,N_3719);
and U3914 (N_3914,N_3704,N_3627);
nand U3915 (N_3915,N_3734,N_3713);
and U3916 (N_3916,N_3630,N_3684);
nand U3917 (N_3917,N_3664,N_3699);
xor U3918 (N_3918,N_3627,N_3651);
nor U3919 (N_3919,N_3659,N_3604);
nor U3920 (N_3920,N_3796,N_3617);
and U3921 (N_3921,N_3609,N_3646);
nor U3922 (N_3922,N_3617,N_3708);
or U3923 (N_3923,N_3739,N_3714);
nor U3924 (N_3924,N_3667,N_3724);
nor U3925 (N_3925,N_3778,N_3654);
nor U3926 (N_3926,N_3675,N_3780);
or U3927 (N_3927,N_3773,N_3721);
and U3928 (N_3928,N_3638,N_3736);
or U3929 (N_3929,N_3706,N_3646);
nor U3930 (N_3930,N_3625,N_3637);
or U3931 (N_3931,N_3606,N_3788);
or U3932 (N_3932,N_3757,N_3691);
nor U3933 (N_3933,N_3660,N_3615);
nor U3934 (N_3934,N_3641,N_3760);
or U3935 (N_3935,N_3658,N_3770);
nor U3936 (N_3936,N_3656,N_3787);
nand U3937 (N_3937,N_3716,N_3735);
nand U3938 (N_3938,N_3727,N_3641);
nand U3939 (N_3939,N_3786,N_3649);
or U3940 (N_3940,N_3632,N_3676);
nor U3941 (N_3941,N_3732,N_3667);
nand U3942 (N_3942,N_3783,N_3799);
nor U3943 (N_3943,N_3750,N_3643);
and U3944 (N_3944,N_3759,N_3675);
or U3945 (N_3945,N_3633,N_3684);
nor U3946 (N_3946,N_3790,N_3724);
or U3947 (N_3947,N_3700,N_3630);
and U3948 (N_3948,N_3600,N_3781);
nand U3949 (N_3949,N_3739,N_3608);
and U3950 (N_3950,N_3689,N_3722);
or U3951 (N_3951,N_3620,N_3730);
and U3952 (N_3952,N_3612,N_3780);
and U3953 (N_3953,N_3730,N_3628);
nor U3954 (N_3954,N_3613,N_3676);
nand U3955 (N_3955,N_3730,N_3644);
nand U3956 (N_3956,N_3687,N_3757);
and U3957 (N_3957,N_3781,N_3724);
and U3958 (N_3958,N_3620,N_3774);
and U3959 (N_3959,N_3701,N_3767);
nor U3960 (N_3960,N_3616,N_3751);
xnor U3961 (N_3961,N_3791,N_3767);
nor U3962 (N_3962,N_3708,N_3719);
and U3963 (N_3963,N_3653,N_3716);
nor U3964 (N_3964,N_3679,N_3648);
nand U3965 (N_3965,N_3753,N_3724);
nand U3966 (N_3966,N_3626,N_3777);
and U3967 (N_3967,N_3682,N_3697);
nand U3968 (N_3968,N_3633,N_3793);
nor U3969 (N_3969,N_3658,N_3651);
or U3970 (N_3970,N_3677,N_3766);
nand U3971 (N_3971,N_3671,N_3707);
and U3972 (N_3972,N_3615,N_3611);
or U3973 (N_3973,N_3761,N_3626);
or U3974 (N_3974,N_3727,N_3665);
or U3975 (N_3975,N_3625,N_3653);
nor U3976 (N_3976,N_3711,N_3658);
nor U3977 (N_3977,N_3769,N_3787);
and U3978 (N_3978,N_3736,N_3689);
nor U3979 (N_3979,N_3713,N_3725);
and U3980 (N_3980,N_3694,N_3676);
nand U3981 (N_3981,N_3730,N_3615);
or U3982 (N_3982,N_3661,N_3629);
xor U3983 (N_3983,N_3609,N_3688);
nand U3984 (N_3984,N_3780,N_3757);
nor U3985 (N_3985,N_3761,N_3683);
and U3986 (N_3986,N_3628,N_3605);
or U3987 (N_3987,N_3695,N_3714);
and U3988 (N_3988,N_3660,N_3719);
nor U3989 (N_3989,N_3764,N_3760);
and U3990 (N_3990,N_3611,N_3654);
nor U3991 (N_3991,N_3793,N_3783);
or U3992 (N_3992,N_3735,N_3650);
or U3993 (N_3993,N_3628,N_3611);
nor U3994 (N_3994,N_3673,N_3769);
or U3995 (N_3995,N_3738,N_3705);
nand U3996 (N_3996,N_3613,N_3783);
nand U3997 (N_3997,N_3611,N_3797);
or U3998 (N_3998,N_3684,N_3629);
and U3999 (N_3999,N_3730,N_3774);
nand U4000 (N_4000,N_3948,N_3802);
or U4001 (N_4001,N_3929,N_3821);
or U4002 (N_4002,N_3898,N_3878);
nor U4003 (N_4003,N_3819,N_3840);
and U4004 (N_4004,N_3993,N_3826);
and U4005 (N_4005,N_3851,N_3931);
and U4006 (N_4006,N_3978,N_3964);
and U4007 (N_4007,N_3858,N_3904);
or U4008 (N_4008,N_3801,N_3998);
nand U4009 (N_4009,N_3943,N_3930);
and U4010 (N_4010,N_3982,N_3823);
nand U4011 (N_4011,N_3979,N_3808);
and U4012 (N_4012,N_3945,N_3951);
nand U4013 (N_4013,N_3970,N_3852);
or U4014 (N_4014,N_3975,N_3902);
nor U4015 (N_4015,N_3992,N_3994);
nand U4016 (N_4016,N_3845,N_3919);
and U4017 (N_4017,N_3922,N_3844);
or U4018 (N_4018,N_3894,N_3969);
nand U4019 (N_4019,N_3838,N_3933);
nand U4020 (N_4020,N_3984,N_3952);
nand U4021 (N_4021,N_3804,N_3927);
nor U4022 (N_4022,N_3849,N_3842);
and U4023 (N_4023,N_3918,N_3863);
nand U4024 (N_4024,N_3911,N_3907);
nand U4025 (N_4025,N_3806,N_3879);
nand U4026 (N_4026,N_3910,N_3967);
and U4027 (N_4027,N_3854,N_3833);
nand U4028 (N_4028,N_3864,N_3848);
and U4029 (N_4029,N_3890,N_3835);
and U4030 (N_4030,N_3891,N_3853);
nor U4031 (N_4031,N_3991,N_3820);
and U4032 (N_4032,N_3814,N_3980);
or U4033 (N_4033,N_3981,N_3834);
nor U4034 (N_4034,N_3875,N_3824);
xnor U4035 (N_4035,N_3822,N_3995);
nor U4036 (N_4036,N_3810,N_3869);
nor U4037 (N_4037,N_3850,N_3928);
nand U4038 (N_4038,N_3989,N_3867);
nor U4039 (N_4039,N_3974,N_3997);
and U4040 (N_4040,N_3914,N_3971);
nor U4041 (N_4041,N_3966,N_3962);
nor U4042 (N_4042,N_3959,N_3940);
and U4043 (N_4043,N_3990,N_3908);
nand U4044 (N_4044,N_3901,N_3868);
or U4045 (N_4045,N_3946,N_3924);
nand U4046 (N_4046,N_3889,N_3950);
nor U4047 (N_4047,N_3941,N_3818);
and U4048 (N_4048,N_3957,N_3986);
nor U4049 (N_4049,N_3881,N_3866);
or U4050 (N_4050,N_3988,N_3809);
nand U4051 (N_4051,N_3909,N_3903);
nor U4052 (N_4052,N_3953,N_3856);
nor U4053 (N_4053,N_3841,N_3800);
nand U4054 (N_4054,N_3843,N_3917);
or U4055 (N_4055,N_3973,N_3932);
or U4056 (N_4056,N_3985,N_3883);
or U4057 (N_4057,N_3897,N_3949);
nand U4058 (N_4058,N_3939,N_3965);
and U4059 (N_4059,N_3885,N_3923);
nand U4060 (N_4060,N_3895,N_3862);
nand U4061 (N_4061,N_3831,N_3815);
nand U4062 (N_4062,N_3837,N_3871);
nand U4063 (N_4063,N_3812,N_3916);
or U4064 (N_4064,N_3884,N_3926);
nor U4065 (N_4065,N_3873,N_3920);
nand U4066 (N_4066,N_3807,N_3936);
nor U4067 (N_4067,N_3861,N_3934);
or U4068 (N_4068,N_3961,N_3882);
nor U4069 (N_4069,N_3976,N_3983);
xnor U4070 (N_4070,N_3960,N_3888);
nand U4071 (N_4071,N_3832,N_3905);
and U4072 (N_4072,N_3938,N_3996);
nand U4073 (N_4073,N_3999,N_3937);
nor U4074 (N_4074,N_3830,N_3987);
nand U4075 (N_4075,N_3935,N_3865);
or U4076 (N_4076,N_3921,N_3860);
or U4077 (N_4077,N_3906,N_3968);
and U4078 (N_4078,N_3956,N_3803);
or U4079 (N_4079,N_3886,N_3913);
nor U4080 (N_4080,N_3925,N_3829);
or U4081 (N_4081,N_3877,N_3972);
nand U4082 (N_4082,N_3947,N_3912);
or U4083 (N_4083,N_3880,N_3899);
nor U4084 (N_4084,N_3811,N_3963);
nor U4085 (N_4085,N_3855,N_3900);
nor U4086 (N_4086,N_3805,N_3954);
or U4087 (N_4087,N_3887,N_3859);
nand U4088 (N_4088,N_3874,N_3817);
and U4089 (N_4089,N_3892,N_3825);
nor U4090 (N_4090,N_3813,N_3816);
or U4091 (N_4091,N_3915,N_3955);
or U4092 (N_4092,N_3896,N_3839);
and U4093 (N_4093,N_3846,N_3836);
and U4094 (N_4094,N_3827,N_3942);
and U4095 (N_4095,N_3958,N_3977);
nor U4096 (N_4096,N_3870,N_3872);
or U4097 (N_4097,N_3828,N_3876);
or U4098 (N_4098,N_3893,N_3847);
nand U4099 (N_4099,N_3944,N_3857);
and U4100 (N_4100,N_3995,N_3929);
and U4101 (N_4101,N_3851,N_3989);
nor U4102 (N_4102,N_3855,N_3992);
nand U4103 (N_4103,N_3842,N_3837);
and U4104 (N_4104,N_3817,N_3984);
and U4105 (N_4105,N_3812,N_3954);
nor U4106 (N_4106,N_3972,N_3921);
and U4107 (N_4107,N_3906,N_3853);
or U4108 (N_4108,N_3823,N_3922);
or U4109 (N_4109,N_3811,N_3982);
and U4110 (N_4110,N_3983,N_3831);
and U4111 (N_4111,N_3990,N_3859);
and U4112 (N_4112,N_3942,N_3957);
and U4113 (N_4113,N_3929,N_3815);
nor U4114 (N_4114,N_3984,N_3853);
or U4115 (N_4115,N_3881,N_3983);
nor U4116 (N_4116,N_3987,N_3928);
nand U4117 (N_4117,N_3923,N_3963);
or U4118 (N_4118,N_3867,N_3871);
nand U4119 (N_4119,N_3829,N_3886);
nand U4120 (N_4120,N_3892,N_3815);
and U4121 (N_4121,N_3813,N_3823);
and U4122 (N_4122,N_3935,N_3973);
nor U4123 (N_4123,N_3829,N_3876);
nand U4124 (N_4124,N_3843,N_3807);
and U4125 (N_4125,N_3823,N_3897);
xnor U4126 (N_4126,N_3991,N_3982);
nand U4127 (N_4127,N_3870,N_3910);
or U4128 (N_4128,N_3879,N_3841);
and U4129 (N_4129,N_3885,N_3909);
nor U4130 (N_4130,N_3954,N_3876);
or U4131 (N_4131,N_3878,N_3836);
and U4132 (N_4132,N_3828,N_3801);
nor U4133 (N_4133,N_3876,N_3870);
and U4134 (N_4134,N_3989,N_3931);
nor U4135 (N_4135,N_3929,N_3868);
nor U4136 (N_4136,N_3873,N_3866);
or U4137 (N_4137,N_3854,N_3873);
nor U4138 (N_4138,N_3967,N_3969);
and U4139 (N_4139,N_3903,N_3800);
or U4140 (N_4140,N_3978,N_3832);
nor U4141 (N_4141,N_3901,N_3803);
nor U4142 (N_4142,N_3887,N_3860);
or U4143 (N_4143,N_3884,N_3980);
nand U4144 (N_4144,N_3860,N_3927);
nor U4145 (N_4145,N_3871,N_3954);
and U4146 (N_4146,N_3955,N_3800);
and U4147 (N_4147,N_3971,N_3806);
nand U4148 (N_4148,N_3910,N_3882);
nand U4149 (N_4149,N_3854,N_3982);
or U4150 (N_4150,N_3970,N_3839);
and U4151 (N_4151,N_3831,N_3944);
and U4152 (N_4152,N_3943,N_3890);
and U4153 (N_4153,N_3957,N_3814);
and U4154 (N_4154,N_3936,N_3998);
nor U4155 (N_4155,N_3971,N_3807);
or U4156 (N_4156,N_3849,N_3835);
nand U4157 (N_4157,N_3996,N_3933);
nand U4158 (N_4158,N_3970,N_3834);
nor U4159 (N_4159,N_3899,N_3970);
nor U4160 (N_4160,N_3881,N_3962);
nand U4161 (N_4161,N_3926,N_3885);
nor U4162 (N_4162,N_3892,N_3955);
or U4163 (N_4163,N_3910,N_3908);
or U4164 (N_4164,N_3833,N_3991);
xnor U4165 (N_4165,N_3883,N_3938);
and U4166 (N_4166,N_3906,N_3964);
nor U4167 (N_4167,N_3888,N_3985);
and U4168 (N_4168,N_3994,N_3924);
nor U4169 (N_4169,N_3835,N_3858);
nand U4170 (N_4170,N_3878,N_3889);
or U4171 (N_4171,N_3872,N_3980);
nand U4172 (N_4172,N_3955,N_3855);
nand U4173 (N_4173,N_3801,N_3866);
or U4174 (N_4174,N_3943,N_3834);
nor U4175 (N_4175,N_3998,N_3827);
xor U4176 (N_4176,N_3859,N_3809);
nor U4177 (N_4177,N_3949,N_3992);
nand U4178 (N_4178,N_3955,N_3805);
nor U4179 (N_4179,N_3857,N_3931);
nand U4180 (N_4180,N_3945,N_3856);
and U4181 (N_4181,N_3895,N_3805);
nand U4182 (N_4182,N_3956,N_3860);
or U4183 (N_4183,N_3922,N_3978);
or U4184 (N_4184,N_3860,N_3967);
and U4185 (N_4185,N_3895,N_3972);
and U4186 (N_4186,N_3944,N_3917);
nand U4187 (N_4187,N_3900,N_3897);
or U4188 (N_4188,N_3875,N_3841);
nor U4189 (N_4189,N_3966,N_3890);
and U4190 (N_4190,N_3954,N_3907);
nand U4191 (N_4191,N_3872,N_3984);
nand U4192 (N_4192,N_3910,N_3865);
nand U4193 (N_4193,N_3877,N_3832);
nand U4194 (N_4194,N_3921,N_3918);
nor U4195 (N_4195,N_3824,N_3929);
nand U4196 (N_4196,N_3838,N_3808);
nand U4197 (N_4197,N_3953,N_3849);
nor U4198 (N_4198,N_3943,N_3900);
or U4199 (N_4199,N_3803,N_3962);
nor U4200 (N_4200,N_4095,N_4004);
or U4201 (N_4201,N_4154,N_4081);
or U4202 (N_4202,N_4120,N_4187);
or U4203 (N_4203,N_4012,N_4073);
nand U4204 (N_4204,N_4186,N_4178);
or U4205 (N_4205,N_4123,N_4116);
nand U4206 (N_4206,N_4079,N_4151);
and U4207 (N_4207,N_4113,N_4170);
and U4208 (N_4208,N_4133,N_4054);
nor U4209 (N_4209,N_4105,N_4180);
or U4210 (N_4210,N_4162,N_4124);
or U4211 (N_4211,N_4036,N_4099);
and U4212 (N_4212,N_4145,N_4006);
nor U4213 (N_4213,N_4074,N_4059);
and U4214 (N_4214,N_4017,N_4129);
nor U4215 (N_4215,N_4098,N_4007);
nand U4216 (N_4216,N_4009,N_4111);
nand U4217 (N_4217,N_4114,N_4031);
and U4218 (N_4218,N_4008,N_4048);
and U4219 (N_4219,N_4002,N_4148);
or U4220 (N_4220,N_4166,N_4051);
or U4221 (N_4221,N_4100,N_4084);
or U4222 (N_4222,N_4069,N_4027);
nor U4223 (N_4223,N_4102,N_4164);
nand U4224 (N_4224,N_4091,N_4001);
and U4225 (N_4225,N_4039,N_4088);
or U4226 (N_4226,N_4107,N_4126);
and U4227 (N_4227,N_4143,N_4174);
nand U4228 (N_4228,N_4147,N_4066);
or U4229 (N_4229,N_4153,N_4061);
and U4230 (N_4230,N_4045,N_4135);
nand U4231 (N_4231,N_4130,N_4092);
nand U4232 (N_4232,N_4060,N_4190);
or U4233 (N_4233,N_4196,N_4049);
and U4234 (N_4234,N_4015,N_4159);
or U4235 (N_4235,N_4115,N_4118);
and U4236 (N_4236,N_4128,N_4056);
nand U4237 (N_4237,N_4044,N_4005);
or U4238 (N_4238,N_4168,N_4052);
or U4239 (N_4239,N_4037,N_4150);
nor U4240 (N_4240,N_4139,N_4000);
or U4241 (N_4241,N_4110,N_4167);
or U4242 (N_4242,N_4109,N_4199);
and U4243 (N_4243,N_4131,N_4137);
or U4244 (N_4244,N_4158,N_4185);
nor U4245 (N_4245,N_4097,N_4014);
nor U4246 (N_4246,N_4046,N_4020);
or U4247 (N_4247,N_4197,N_4138);
or U4248 (N_4248,N_4163,N_4101);
xor U4249 (N_4249,N_4025,N_4161);
nor U4250 (N_4250,N_4089,N_4112);
or U4251 (N_4251,N_4042,N_4171);
and U4252 (N_4252,N_4157,N_4043);
or U4253 (N_4253,N_4075,N_4077);
xnor U4254 (N_4254,N_4189,N_4010);
or U4255 (N_4255,N_4125,N_4177);
nor U4256 (N_4256,N_4041,N_4016);
or U4257 (N_4257,N_4179,N_4030);
nor U4258 (N_4258,N_4011,N_4176);
nor U4259 (N_4259,N_4033,N_4076);
and U4260 (N_4260,N_4122,N_4188);
or U4261 (N_4261,N_4144,N_4195);
nand U4262 (N_4262,N_4050,N_4149);
nor U4263 (N_4263,N_4182,N_4018);
nor U4264 (N_4264,N_4071,N_4136);
nand U4265 (N_4265,N_4085,N_4019);
nand U4266 (N_4266,N_4198,N_4181);
or U4267 (N_4267,N_4024,N_4169);
nor U4268 (N_4268,N_4068,N_4029);
and U4269 (N_4269,N_4086,N_4175);
and U4270 (N_4270,N_4140,N_4155);
nor U4271 (N_4271,N_4106,N_4152);
nor U4272 (N_4272,N_4032,N_4119);
or U4273 (N_4273,N_4034,N_4090);
nor U4274 (N_4274,N_4062,N_4165);
nand U4275 (N_4275,N_4047,N_4193);
and U4276 (N_4276,N_4184,N_4087);
and U4277 (N_4277,N_4093,N_4078);
or U4278 (N_4278,N_4083,N_4121);
nor U4279 (N_4279,N_4064,N_4172);
and U4280 (N_4280,N_4173,N_4058);
nand U4281 (N_4281,N_4082,N_4194);
nand U4282 (N_4282,N_4053,N_4022);
nand U4283 (N_4283,N_4142,N_4003);
nor U4284 (N_4284,N_4127,N_4013);
and U4285 (N_4285,N_4096,N_4117);
or U4286 (N_4286,N_4104,N_4028);
nand U4287 (N_4287,N_4103,N_4141);
nor U4288 (N_4288,N_4156,N_4134);
and U4289 (N_4289,N_4035,N_4072);
nor U4290 (N_4290,N_4055,N_4191);
or U4291 (N_4291,N_4192,N_4094);
nand U4292 (N_4292,N_4038,N_4070);
nor U4293 (N_4293,N_4021,N_4132);
nand U4294 (N_4294,N_4160,N_4023);
and U4295 (N_4295,N_4057,N_4146);
nor U4296 (N_4296,N_4080,N_4183);
or U4297 (N_4297,N_4108,N_4026);
and U4298 (N_4298,N_4063,N_4067);
or U4299 (N_4299,N_4040,N_4065);
nand U4300 (N_4300,N_4133,N_4117);
nand U4301 (N_4301,N_4135,N_4065);
nor U4302 (N_4302,N_4024,N_4193);
and U4303 (N_4303,N_4060,N_4010);
nand U4304 (N_4304,N_4198,N_4152);
and U4305 (N_4305,N_4181,N_4142);
and U4306 (N_4306,N_4056,N_4156);
nand U4307 (N_4307,N_4061,N_4106);
and U4308 (N_4308,N_4142,N_4054);
or U4309 (N_4309,N_4059,N_4096);
nor U4310 (N_4310,N_4066,N_4095);
or U4311 (N_4311,N_4173,N_4001);
and U4312 (N_4312,N_4130,N_4062);
nand U4313 (N_4313,N_4084,N_4073);
and U4314 (N_4314,N_4039,N_4104);
nand U4315 (N_4315,N_4025,N_4183);
nor U4316 (N_4316,N_4089,N_4100);
nand U4317 (N_4317,N_4044,N_4168);
or U4318 (N_4318,N_4140,N_4117);
nor U4319 (N_4319,N_4057,N_4153);
xnor U4320 (N_4320,N_4035,N_4009);
nor U4321 (N_4321,N_4092,N_4137);
nand U4322 (N_4322,N_4171,N_4138);
nand U4323 (N_4323,N_4002,N_4064);
nand U4324 (N_4324,N_4168,N_4075);
and U4325 (N_4325,N_4047,N_4167);
nand U4326 (N_4326,N_4178,N_4031);
nand U4327 (N_4327,N_4049,N_4067);
or U4328 (N_4328,N_4132,N_4167);
and U4329 (N_4329,N_4118,N_4165);
and U4330 (N_4330,N_4136,N_4085);
nand U4331 (N_4331,N_4083,N_4050);
nand U4332 (N_4332,N_4118,N_4117);
nand U4333 (N_4333,N_4164,N_4059);
and U4334 (N_4334,N_4101,N_4114);
and U4335 (N_4335,N_4100,N_4060);
xnor U4336 (N_4336,N_4158,N_4146);
and U4337 (N_4337,N_4019,N_4153);
nand U4338 (N_4338,N_4115,N_4001);
or U4339 (N_4339,N_4062,N_4057);
nor U4340 (N_4340,N_4184,N_4066);
xor U4341 (N_4341,N_4036,N_4101);
nand U4342 (N_4342,N_4111,N_4137);
nor U4343 (N_4343,N_4132,N_4080);
nor U4344 (N_4344,N_4196,N_4095);
nand U4345 (N_4345,N_4008,N_4117);
or U4346 (N_4346,N_4139,N_4162);
nand U4347 (N_4347,N_4057,N_4049);
or U4348 (N_4348,N_4143,N_4009);
xor U4349 (N_4349,N_4098,N_4119);
nand U4350 (N_4350,N_4018,N_4128);
and U4351 (N_4351,N_4108,N_4020);
and U4352 (N_4352,N_4158,N_4090);
and U4353 (N_4353,N_4022,N_4051);
or U4354 (N_4354,N_4040,N_4093);
nand U4355 (N_4355,N_4050,N_4136);
nand U4356 (N_4356,N_4095,N_4016);
and U4357 (N_4357,N_4054,N_4049);
nor U4358 (N_4358,N_4150,N_4128);
nand U4359 (N_4359,N_4006,N_4126);
or U4360 (N_4360,N_4184,N_4127);
nor U4361 (N_4361,N_4152,N_4172);
or U4362 (N_4362,N_4167,N_4184);
and U4363 (N_4363,N_4110,N_4045);
and U4364 (N_4364,N_4065,N_4024);
nor U4365 (N_4365,N_4005,N_4021);
nor U4366 (N_4366,N_4097,N_4062);
nand U4367 (N_4367,N_4176,N_4040);
nand U4368 (N_4368,N_4042,N_4059);
and U4369 (N_4369,N_4066,N_4030);
and U4370 (N_4370,N_4032,N_4152);
and U4371 (N_4371,N_4056,N_4180);
and U4372 (N_4372,N_4013,N_4063);
or U4373 (N_4373,N_4050,N_4169);
and U4374 (N_4374,N_4123,N_4010);
nor U4375 (N_4375,N_4073,N_4005);
and U4376 (N_4376,N_4112,N_4063);
and U4377 (N_4377,N_4002,N_4155);
and U4378 (N_4378,N_4186,N_4160);
nand U4379 (N_4379,N_4111,N_4002);
nand U4380 (N_4380,N_4134,N_4098);
nor U4381 (N_4381,N_4146,N_4135);
nor U4382 (N_4382,N_4100,N_4005);
or U4383 (N_4383,N_4032,N_4093);
nand U4384 (N_4384,N_4017,N_4088);
nand U4385 (N_4385,N_4146,N_4003);
or U4386 (N_4386,N_4154,N_4173);
and U4387 (N_4387,N_4029,N_4174);
and U4388 (N_4388,N_4041,N_4085);
nand U4389 (N_4389,N_4027,N_4182);
or U4390 (N_4390,N_4181,N_4018);
nor U4391 (N_4391,N_4063,N_4031);
and U4392 (N_4392,N_4013,N_4095);
and U4393 (N_4393,N_4005,N_4069);
or U4394 (N_4394,N_4037,N_4125);
nor U4395 (N_4395,N_4051,N_4005);
nor U4396 (N_4396,N_4052,N_4036);
and U4397 (N_4397,N_4192,N_4012);
and U4398 (N_4398,N_4153,N_4113);
nand U4399 (N_4399,N_4132,N_4184);
and U4400 (N_4400,N_4250,N_4245);
and U4401 (N_4401,N_4322,N_4312);
nand U4402 (N_4402,N_4348,N_4267);
and U4403 (N_4403,N_4328,N_4356);
and U4404 (N_4404,N_4284,N_4384);
or U4405 (N_4405,N_4238,N_4352);
nor U4406 (N_4406,N_4357,N_4371);
nand U4407 (N_4407,N_4265,N_4351);
nand U4408 (N_4408,N_4343,N_4239);
nor U4409 (N_4409,N_4347,N_4386);
or U4410 (N_4410,N_4337,N_4314);
and U4411 (N_4411,N_4358,N_4307);
nand U4412 (N_4412,N_4233,N_4216);
nor U4413 (N_4413,N_4393,N_4395);
or U4414 (N_4414,N_4211,N_4361);
or U4415 (N_4415,N_4215,N_4375);
nor U4416 (N_4416,N_4226,N_4303);
nor U4417 (N_4417,N_4300,N_4364);
or U4418 (N_4418,N_4212,N_4362);
nor U4419 (N_4419,N_4349,N_4323);
nor U4420 (N_4420,N_4268,N_4333);
nand U4421 (N_4421,N_4370,N_4329);
or U4422 (N_4422,N_4260,N_4276);
or U4423 (N_4423,N_4293,N_4301);
or U4424 (N_4424,N_4382,N_4278);
nand U4425 (N_4425,N_4374,N_4202);
and U4426 (N_4426,N_4366,N_4200);
or U4427 (N_4427,N_4282,N_4299);
nor U4428 (N_4428,N_4380,N_4230);
or U4429 (N_4429,N_4368,N_4372);
nand U4430 (N_4430,N_4206,N_4399);
nor U4431 (N_4431,N_4221,N_4365);
and U4432 (N_4432,N_4305,N_4255);
and U4433 (N_4433,N_4251,N_4252);
or U4434 (N_4434,N_4376,N_4218);
and U4435 (N_4435,N_4344,N_4317);
nor U4436 (N_4436,N_4290,N_4394);
or U4437 (N_4437,N_4346,N_4367);
and U4438 (N_4438,N_4275,N_4355);
nand U4439 (N_4439,N_4208,N_4283);
nand U4440 (N_4440,N_4389,N_4330);
nor U4441 (N_4441,N_4280,N_4273);
nand U4442 (N_4442,N_4397,N_4227);
or U4443 (N_4443,N_4246,N_4334);
and U4444 (N_4444,N_4306,N_4225);
nand U4445 (N_4445,N_4277,N_4271);
nand U4446 (N_4446,N_4237,N_4287);
and U4447 (N_4447,N_4315,N_4220);
and U4448 (N_4448,N_4342,N_4304);
and U4449 (N_4449,N_4338,N_4207);
nand U4450 (N_4450,N_4257,N_4231);
or U4451 (N_4451,N_4224,N_4331);
and U4452 (N_4452,N_4345,N_4219);
nand U4453 (N_4453,N_4209,N_4248);
or U4454 (N_4454,N_4388,N_4340);
nand U4455 (N_4455,N_4288,N_4321);
or U4456 (N_4456,N_4373,N_4274);
nand U4457 (N_4457,N_4232,N_4359);
or U4458 (N_4458,N_4327,N_4201);
and U4459 (N_4459,N_4294,N_4295);
nand U4460 (N_4460,N_4217,N_4378);
nand U4461 (N_4461,N_4286,N_4297);
xor U4462 (N_4462,N_4289,N_4236);
and U4463 (N_4463,N_4360,N_4387);
or U4464 (N_4464,N_4244,N_4223);
nor U4465 (N_4465,N_4249,N_4264);
and U4466 (N_4466,N_4256,N_4354);
and U4467 (N_4467,N_4204,N_4279);
nor U4468 (N_4468,N_4261,N_4324);
nand U4469 (N_4469,N_4332,N_4222);
xor U4470 (N_4470,N_4292,N_4377);
or U4471 (N_4471,N_4214,N_4398);
or U4472 (N_4472,N_4363,N_4205);
or U4473 (N_4473,N_4241,N_4341);
or U4474 (N_4474,N_4259,N_4254);
nor U4475 (N_4475,N_4298,N_4291);
nor U4476 (N_4476,N_4381,N_4313);
and U4477 (N_4477,N_4318,N_4281);
and U4478 (N_4478,N_4369,N_4272);
or U4479 (N_4479,N_4336,N_4319);
nor U4480 (N_4480,N_4390,N_4309);
and U4481 (N_4481,N_4213,N_4229);
nand U4482 (N_4482,N_4262,N_4326);
or U4483 (N_4483,N_4383,N_4263);
nor U4484 (N_4484,N_4379,N_4253);
nand U4485 (N_4485,N_4266,N_4335);
nor U4486 (N_4486,N_4269,N_4311);
nor U4487 (N_4487,N_4235,N_4391);
or U4488 (N_4488,N_4385,N_4247);
nor U4489 (N_4489,N_4350,N_4243);
or U4490 (N_4490,N_4210,N_4240);
nor U4491 (N_4491,N_4320,N_4339);
nor U4492 (N_4492,N_4270,N_4392);
nand U4493 (N_4493,N_4228,N_4396);
nor U4494 (N_4494,N_4308,N_4296);
or U4495 (N_4495,N_4310,N_4325);
nor U4496 (N_4496,N_4234,N_4285);
nand U4497 (N_4497,N_4203,N_4302);
nor U4498 (N_4498,N_4242,N_4258);
and U4499 (N_4499,N_4316,N_4353);
or U4500 (N_4500,N_4205,N_4395);
nor U4501 (N_4501,N_4365,N_4235);
and U4502 (N_4502,N_4304,N_4293);
and U4503 (N_4503,N_4336,N_4321);
or U4504 (N_4504,N_4323,N_4385);
nor U4505 (N_4505,N_4256,N_4304);
or U4506 (N_4506,N_4252,N_4244);
or U4507 (N_4507,N_4239,N_4269);
or U4508 (N_4508,N_4393,N_4347);
nand U4509 (N_4509,N_4321,N_4302);
or U4510 (N_4510,N_4215,N_4297);
nor U4511 (N_4511,N_4377,N_4391);
and U4512 (N_4512,N_4325,N_4344);
nand U4513 (N_4513,N_4256,N_4208);
or U4514 (N_4514,N_4317,N_4223);
or U4515 (N_4515,N_4326,N_4373);
nand U4516 (N_4516,N_4358,N_4204);
and U4517 (N_4517,N_4357,N_4315);
nor U4518 (N_4518,N_4341,N_4205);
nor U4519 (N_4519,N_4347,N_4369);
nand U4520 (N_4520,N_4258,N_4214);
nor U4521 (N_4521,N_4235,N_4314);
nand U4522 (N_4522,N_4377,N_4212);
and U4523 (N_4523,N_4369,N_4368);
nor U4524 (N_4524,N_4352,N_4340);
nor U4525 (N_4525,N_4295,N_4364);
nand U4526 (N_4526,N_4382,N_4388);
and U4527 (N_4527,N_4340,N_4353);
nor U4528 (N_4528,N_4313,N_4273);
or U4529 (N_4529,N_4303,N_4245);
xor U4530 (N_4530,N_4334,N_4258);
nor U4531 (N_4531,N_4284,N_4256);
and U4532 (N_4532,N_4379,N_4317);
and U4533 (N_4533,N_4254,N_4297);
or U4534 (N_4534,N_4252,N_4220);
nand U4535 (N_4535,N_4258,N_4207);
and U4536 (N_4536,N_4375,N_4322);
or U4537 (N_4537,N_4228,N_4321);
and U4538 (N_4538,N_4385,N_4304);
nor U4539 (N_4539,N_4201,N_4356);
nor U4540 (N_4540,N_4381,N_4315);
or U4541 (N_4541,N_4247,N_4389);
nor U4542 (N_4542,N_4372,N_4324);
nor U4543 (N_4543,N_4278,N_4379);
or U4544 (N_4544,N_4237,N_4221);
nand U4545 (N_4545,N_4203,N_4202);
or U4546 (N_4546,N_4362,N_4203);
or U4547 (N_4547,N_4375,N_4216);
nand U4548 (N_4548,N_4331,N_4354);
nor U4549 (N_4549,N_4269,N_4260);
nand U4550 (N_4550,N_4373,N_4350);
nand U4551 (N_4551,N_4348,N_4217);
or U4552 (N_4552,N_4314,N_4277);
nor U4553 (N_4553,N_4341,N_4313);
nand U4554 (N_4554,N_4329,N_4203);
and U4555 (N_4555,N_4320,N_4293);
and U4556 (N_4556,N_4208,N_4338);
nor U4557 (N_4557,N_4385,N_4368);
nor U4558 (N_4558,N_4389,N_4366);
xnor U4559 (N_4559,N_4371,N_4391);
nor U4560 (N_4560,N_4203,N_4357);
or U4561 (N_4561,N_4394,N_4278);
and U4562 (N_4562,N_4234,N_4376);
nand U4563 (N_4563,N_4276,N_4258);
nor U4564 (N_4564,N_4223,N_4251);
and U4565 (N_4565,N_4370,N_4340);
nor U4566 (N_4566,N_4265,N_4378);
nand U4567 (N_4567,N_4280,N_4236);
and U4568 (N_4568,N_4250,N_4349);
or U4569 (N_4569,N_4281,N_4223);
nor U4570 (N_4570,N_4305,N_4370);
or U4571 (N_4571,N_4293,N_4340);
nor U4572 (N_4572,N_4382,N_4237);
nand U4573 (N_4573,N_4393,N_4235);
and U4574 (N_4574,N_4300,N_4297);
or U4575 (N_4575,N_4358,N_4251);
and U4576 (N_4576,N_4382,N_4267);
nor U4577 (N_4577,N_4259,N_4272);
or U4578 (N_4578,N_4233,N_4207);
and U4579 (N_4579,N_4236,N_4340);
and U4580 (N_4580,N_4214,N_4368);
xor U4581 (N_4581,N_4279,N_4291);
nand U4582 (N_4582,N_4217,N_4259);
or U4583 (N_4583,N_4243,N_4261);
and U4584 (N_4584,N_4238,N_4345);
nand U4585 (N_4585,N_4301,N_4240);
and U4586 (N_4586,N_4256,N_4337);
nor U4587 (N_4587,N_4291,N_4356);
and U4588 (N_4588,N_4237,N_4316);
nor U4589 (N_4589,N_4273,N_4211);
and U4590 (N_4590,N_4375,N_4396);
nor U4591 (N_4591,N_4338,N_4322);
or U4592 (N_4592,N_4214,N_4213);
or U4593 (N_4593,N_4352,N_4390);
or U4594 (N_4594,N_4379,N_4337);
and U4595 (N_4595,N_4368,N_4209);
nor U4596 (N_4596,N_4244,N_4301);
nand U4597 (N_4597,N_4285,N_4368);
nor U4598 (N_4598,N_4397,N_4223);
and U4599 (N_4599,N_4271,N_4274);
nor U4600 (N_4600,N_4435,N_4591);
or U4601 (N_4601,N_4489,N_4565);
nand U4602 (N_4602,N_4443,N_4549);
nor U4603 (N_4603,N_4590,N_4563);
and U4604 (N_4604,N_4496,N_4556);
or U4605 (N_4605,N_4525,N_4479);
and U4606 (N_4606,N_4481,N_4430);
or U4607 (N_4607,N_4582,N_4548);
and U4608 (N_4608,N_4573,N_4567);
nor U4609 (N_4609,N_4533,N_4453);
or U4610 (N_4610,N_4597,N_4423);
nand U4611 (N_4611,N_4519,N_4522);
and U4612 (N_4612,N_4578,N_4595);
and U4613 (N_4613,N_4583,N_4586);
nand U4614 (N_4614,N_4524,N_4551);
or U4615 (N_4615,N_4436,N_4521);
nor U4616 (N_4616,N_4514,N_4469);
nand U4617 (N_4617,N_4598,N_4488);
nor U4618 (N_4618,N_4425,N_4542);
and U4619 (N_4619,N_4486,N_4570);
nor U4620 (N_4620,N_4465,N_4404);
and U4621 (N_4621,N_4528,N_4501);
nand U4622 (N_4622,N_4456,N_4449);
or U4623 (N_4623,N_4500,N_4434);
or U4624 (N_4624,N_4530,N_4566);
and U4625 (N_4625,N_4596,N_4510);
nor U4626 (N_4626,N_4538,N_4473);
and U4627 (N_4627,N_4448,N_4568);
nand U4628 (N_4628,N_4499,N_4503);
nand U4629 (N_4629,N_4403,N_4508);
nand U4630 (N_4630,N_4461,N_4491);
and U4631 (N_4631,N_4547,N_4516);
or U4632 (N_4632,N_4402,N_4438);
nor U4633 (N_4633,N_4541,N_4559);
nand U4634 (N_4634,N_4405,N_4526);
nor U4635 (N_4635,N_4484,N_4564);
nand U4636 (N_4636,N_4544,N_4589);
nand U4637 (N_4637,N_4447,N_4537);
nand U4638 (N_4638,N_4413,N_4477);
or U4639 (N_4639,N_4409,N_4463);
and U4640 (N_4640,N_4459,N_4588);
nand U4641 (N_4641,N_4444,N_4407);
nor U4642 (N_4642,N_4460,N_4527);
nand U4643 (N_4643,N_4467,N_4552);
or U4644 (N_4644,N_4575,N_4584);
nand U4645 (N_4645,N_4506,N_4440);
or U4646 (N_4646,N_4464,N_4441);
or U4647 (N_4647,N_4452,N_4468);
or U4648 (N_4648,N_4458,N_4412);
and U4649 (N_4649,N_4502,N_4482);
nor U4650 (N_4650,N_4437,N_4408);
nand U4651 (N_4651,N_4487,N_4427);
and U4652 (N_4652,N_4572,N_4555);
nor U4653 (N_4653,N_4536,N_4557);
or U4654 (N_4654,N_4561,N_4517);
and U4655 (N_4655,N_4462,N_4497);
nand U4656 (N_4656,N_4580,N_4439);
or U4657 (N_4657,N_4422,N_4543);
nand U4658 (N_4658,N_4470,N_4478);
nand U4659 (N_4659,N_4535,N_4593);
or U4660 (N_4660,N_4581,N_4546);
and U4661 (N_4661,N_4431,N_4429);
nand U4662 (N_4662,N_4445,N_4520);
nor U4663 (N_4663,N_4594,N_4466);
nand U4664 (N_4664,N_4529,N_4498);
and U4665 (N_4665,N_4454,N_4476);
and U4666 (N_4666,N_4419,N_4442);
nor U4667 (N_4667,N_4574,N_4550);
nor U4668 (N_4668,N_4505,N_4599);
and U4669 (N_4669,N_4421,N_4490);
or U4670 (N_4670,N_4426,N_4457);
and U4671 (N_4671,N_4553,N_4579);
nand U4672 (N_4672,N_4523,N_4592);
and U4673 (N_4673,N_4455,N_4446);
nor U4674 (N_4674,N_4577,N_4415);
or U4675 (N_4675,N_4512,N_4451);
nand U4676 (N_4676,N_4401,N_4513);
nor U4677 (N_4677,N_4532,N_4545);
and U4678 (N_4678,N_4420,N_4587);
nor U4679 (N_4679,N_4400,N_4417);
nor U4680 (N_4680,N_4494,N_4433);
nand U4681 (N_4681,N_4492,N_4507);
nor U4682 (N_4682,N_4540,N_4539);
or U4683 (N_4683,N_4406,N_4428);
nand U4684 (N_4684,N_4554,N_4560);
or U4685 (N_4685,N_4418,N_4474);
and U4686 (N_4686,N_4511,N_4518);
or U4687 (N_4687,N_4472,N_4495);
nor U4688 (N_4688,N_4509,N_4414);
or U4689 (N_4689,N_4485,N_4410);
nand U4690 (N_4690,N_4534,N_4569);
nor U4691 (N_4691,N_4416,N_4483);
and U4692 (N_4692,N_4562,N_4450);
nor U4693 (N_4693,N_4571,N_4471);
nor U4694 (N_4694,N_4475,N_4576);
or U4695 (N_4695,N_4585,N_4531);
nor U4696 (N_4696,N_4493,N_4424);
nand U4697 (N_4697,N_4480,N_4411);
nor U4698 (N_4698,N_4558,N_4504);
nand U4699 (N_4699,N_4515,N_4432);
or U4700 (N_4700,N_4490,N_4594);
and U4701 (N_4701,N_4438,N_4411);
and U4702 (N_4702,N_4411,N_4531);
or U4703 (N_4703,N_4587,N_4546);
nor U4704 (N_4704,N_4483,N_4511);
and U4705 (N_4705,N_4483,N_4512);
or U4706 (N_4706,N_4450,N_4401);
or U4707 (N_4707,N_4480,N_4416);
nor U4708 (N_4708,N_4509,N_4486);
and U4709 (N_4709,N_4594,N_4512);
nand U4710 (N_4710,N_4401,N_4417);
nand U4711 (N_4711,N_4411,N_4446);
nand U4712 (N_4712,N_4438,N_4443);
nor U4713 (N_4713,N_4593,N_4439);
nand U4714 (N_4714,N_4464,N_4494);
and U4715 (N_4715,N_4424,N_4555);
nand U4716 (N_4716,N_4559,N_4427);
and U4717 (N_4717,N_4432,N_4423);
and U4718 (N_4718,N_4537,N_4430);
nor U4719 (N_4719,N_4573,N_4563);
nor U4720 (N_4720,N_4436,N_4502);
nor U4721 (N_4721,N_4547,N_4544);
nor U4722 (N_4722,N_4437,N_4464);
or U4723 (N_4723,N_4450,N_4507);
and U4724 (N_4724,N_4483,N_4599);
and U4725 (N_4725,N_4472,N_4418);
nand U4726 (N_4726,N_4429,N_4438);
and U4727 (N_4727,N_4587,N_4567);
or U4728 (N_4728,N_4515,N_4559);
xor U4729 (N_4729,N_4548,N_4596);
and U4730 (N_4730,N_4519,N_4456);
or U4731 (N_4731,N_4445,N_4411);
and U4732 (N_4732,N_4495,N_4543);
or U4733 (N_4733,N_4442,N_4446);
nand U4734 (N_4734,N_4542,N_4508);
and U4735 (N_4735,N_4525,N_4512);
nor U4736 (N_4736,N_4400,N_4425);
nand U4737 (N_4737,N_4426,N_4540);
nor U4738 (N_4738,N_4482,N_4554);
nor U4739 (N_4739,N_4565,N_4473);
nand U4740 (N_4740,N_4523,N_4443);
nand U4741 (N_4741,N_4563,N_4597);
nor U4742 (N_4742,N_4418,N_4516);
nor U4743 (N_4743,N_4505,N_4405);
or U4744 (N_4744,N_4557,N_4413);
nor U4745 (N_4745,N_4568,N_4549);
and U4746 (N_4746,N_4492,N_4403);
or U4747 (N_4747,N_4409,N_4594);
or U4748 (N_4748,N_4599,N_4536);
and U4749 (N_4749,N_4450,N_4522);
or U4750 (N_4750,N_4400,N_4456);
and U4751 (N_4751,N_4450,N_4405);
and U4752 (N_4752,N_4531,N_4534);
and U4753 (N_4753,N_4509,N_4493);
or U4754 (N_4754,N_4583,N_4553);
nor U4755 (N_4755,N_4538,N_4509);
nand U4756 (N_4756,N_4457,N_4401);
and U4757 (N_4757,N_4464,N_4483);
nor U4758 (N_4758,N_4457,N_4545);
nor U4759 (N_4759,N_4465,N_4452);
nor U4760 (N_4760,N_4589,N_4412);
or U4761 (N_4761,N_4434,N_4419);
or U4762 (N_4762,N_4444,N_4493);
or U4763 (N_4763,N_4497,N_4539);
nor U4764 (N_4764,N_4595,N_4401);
nand U4765 (N_4765,N_4447,N_4544);
and U4766 (N_4766,N_4574,N_4487);
nor U4767 (N_4767,N_4498,N_4515);
nand U4768 (N_4768,N_4414,N_4493);
nor U4769 (N_4769,N_4512,N_4492);
or U4770 (N_4770,N_4584,N_4435);
nand U4771 (N_4771,N_4571,N_4424);
or U4772 (N_4772,N_4531,N_4527);
nor U4773 (N_4773,N_4507,N_4414);
or U4774 (N_4774,N_4416,N_4430);
nor U4775 (N_4775,N_4588,N_4472);
nand U4776 (N_4776,N_4488,N_4458);
and U4777 (N_4777,N_4448,N_4466);
or U4778 (N_4778,N_4517,N_4443);
nand U4779 (N_4779,N_4526,N_4437);
and U4780 (N_4780,N_4401,N_4552);
nor U4781 (N_4781,N_4561,N_4489);
nor U4782 (N_4782,N_4440,N_4424);
nand U4783 (N_4783,N_4407,N_4517);
and U4784 (N_4784,N_4442,N_4595);
nor U4785 (N_4785,N_4511,N_4463);
nor U4786 (N_4786,N_4570,N_4499);
or U4787 (N_4787,N_4566,N_4416);
and U4788 (N_4788,N_4582,N_4468);
and U4789 (N_4789,N_4499,N_4547);
nand U4790 (N_4790,N_4524,N_4418);
nand U4791 (N_4791,N_4522,N_4464);
nor U4792 (N_4792,N_4512,N_4597);
and U4793 (N_4793,N_4417,N_4449);
and U4794 (N_4794,N_4571,N_4512);
or U4795 (N_4795,N_4535,N_4582);
nand U4796 (N_4796,N_4517,N_4429);
and U4797 (N_4797,N_4476,N_4466);
nor U4798 (N_4798,N_4586,N_4520);
and U4799 (N_4799,N_4547,N_4480);
nor U4800 (N_4800,N_4668,N_4625);
and U4801 (N_4801,N_4600,N_4611);
or U4802 (N_4802,N_4710,N_4716);
and U4803 (N_4803,N_4749,N_4689);
and U4804 (N_4804,N_4660,N_4702);
xnor U4805 (N_4805,N_4667,N_4721);
nand U4806 (N_4806,N_4651,N_4615);
nor U4807 (N_4807,N_4727,N_4766);
nor U4808 (N_4808,N_4735,N_4671);
and U4809 (N_4809,N_4670,N_4736);
nand U4810 (N_4810,N_4718,N_4664);
and U4811 (N_4811,N_4786,N_4753);
and U4812 (N_4812,N_4764,N_4769);
or U4813 (N_4813,N_4709,N_4791);
and U4814 (N_4814,N_4708,N_4799);
or U4815 (N_4815,N_4606,N_4740);
and U4816 (N_4816,N_4657,N_4618);
or U4817 (N_4817,N_4647,N_4772);
nor U4818 (N_4818,N_4674,N_4713);
or U4819 (N_4819,N_4744,N_4682);
or U4820 (N_4820,N_4707,N_4739);
and U4821 (N_4821,N_4691,N_4617);
nand U4822 (N_4822,N_4788,N_4763);
nand U4823 (N_4823,N_4659,N_4728);
or U4824 (N_4824,N_4720,N_4774);
and U4825 (N_4825,N_4726,N_4692);
and U4826 (N_4826,N_4782,N_4656);
and U4827 (N_4827,N_4648,N_4759);
and U4828 (N_4828,N_4601,N_4655);
nand U4829 (N_4829,N_4737,N_4604);
nor U4830 (N_4830,N_4704,N_4662);
and U4831 (N_4831,N_4738,N_4676);
nor U4832 (N_4832,N_4645,N_4694);
nor U4833 (N_4833,N_4652,N_4781);
or U4834 (N_4834,N_4747,N_4731);
nand U4835 (N_4835,N_4658,N_4722);
or U4836 (N_4836,N_4609,N_4614);
nor U4837 (N_4837,N_4665,N_4733);
nand U4838 (N_4838,N_4717,N_4608);
xnor U4839 (N_4839,N_4777,N_4603);
nor U4840 (N_4840,N_4767,N_4790);
nand U4841 (N_4841,N_4765,N_4621);
and U4842 (N_4842,N_4636,N_4612);
nand U4843 (N_4843,N_4632,N_4687);
and U4844 (N_4844,N_4783,N_4785);
nand U4845 (N_4845,N_4638,N_4698);
or U4846 (N_4846,N_4754,N_4641);
nor U4847 (N_4847,N_4684,N_4616);
or U4848 (N_4848,N_4789,N_4607);
nor U4849 (N_4849,N_4680,N_4643);
nor U4850 (N_4850,N_4771,N_4624);
nand U4851 (N_4851,N_4755,N_4743);
and U4852 (N_4852,N_4703,N_4635);
and U4853 (N_4853,N_4768,N_4773);
nand U4854 (N_4854,N_4775,N_4639);
nand U4855 (N_4855,N_4634,N_4675);
and U4856 (N_4856,N_4795,N_4619);
nand U4857 (N_4857,N_4719,N_4792);
or U4858 (N_4858,N_4760,N_4650);
or U4859 (N_4859,N_4693,N_4796);
or U4860 (N_4860,N_4734,N_4688);
or U4861 (N_4861,N_4752,N_4715);
nand U4862 (N_4862,N_4701,N_4654);
nand U4863 (N_4863,N_4623,N_4745);
nand U4864 (N_4864,N_4613,N_4685);
or U4865 (N_4865,N_4661,N_4673);
and U4866 (N_4866,N_4602,N_4798);
nor U4867 (N_4867,N_4669,N_4620);
nor U4868 (N_4868,N_4725,N_4761);
nand U4869 (N_4869,N_4683,N_4678);
and U4870 (N_4870,N_4646,N_4712);
and U4871 (N_4871,N_4756,N_4714);
and U4872 (N_4872,N_4695,N_4750);
and U4873 (N_4873,N_4776,N_4778);
or U4874 (N_4874,N_4622,N_4681);
nor U4875 (N_4875,N_4644,N_4653);
nand U4876 (N_4876,N_4631,N_4751);
and U4877 (N_4877,N_4780,N_4706);
nor U4878 (N_4878,N_4627,N_4672);
and U4879 (N_4879,N_4758,N_4730);
nor U4880 (N_4880,N_4629,N_4679);
or U4881 (N_4881,N_4762,N_4610);
or U4882 (N_4882,N_4723,N_4697);
nor U4883 (N_4883,N_4605,N_4677);
nand U4884 (N_4884,N_4699,N_4640);
nor U4885 (N_4885,N_4630,N_4700);
xnor U4886 (N_4886,N_4686,N_4637);
nand U4887 (N_4887,N_4729,N_4705);
and U4888 (N_4888,N_4649,N_4794);
and U4889 (N_4889,N_4724,N_4741);
or U4890 (N_4890,N_4633,N_4779);
and U4891 (N_4891,N_4787,N_4746);
or U4892 (N_4892,N_4797,N_4628);
nor U4893 (N_4893,N_4663,N_4732);
or U4894 (N_4894,N_4770,N_4793);
and U4895 (N_4895,N_4711,N_4666);
or U4896 (N_4896,N_4690,N_4742);
xnor U4897 (N_4897,N_4626,N_4748);
nor U4898 (N_4898,N_4642,N_4757);
nor U4899 (N_4899,N_4696,N_4784);
nor U4900 (N_4900,N_4724,N_4608);
or U4901 (N_4901,N_4609,N_4664);
or U4902 (N_4902,N_4729,N_4784);
or U4903 (N_4903,N_4614,N_4788);
or U4904 (N_4904,N_4656,N_4648);
and U4905 (N_4905,N_4638,N_4711);
nand U4906 (N_4906,N_4739,N_4696);
or U4907 (N_4907,N_4785,N_4708);
xor U4908 (N_4908,N_4638,N_4660);
xnor U4909 (N_4909,N_4702,N_4666);
or U4910 (N_4910,N_4603,N_4735);
nor U4911 (N_4911,N_4784,N_4644);
nand U4912 (N_4912,N_4646,N_4773);
or U4913 (N_4913,N_4789,N_4623);
xnor U4914 (N_4914,N_4628,N_4697);
nor U4915 (N_4915,N_4763,N_4756);
or U4916 (N_4916,N_4783,N_4788);
nor U4917 (N_4917,N_4691,N_4633);
and U4918 (N_4918,N_4637,N_4749);
and U4919 (N_4919,N_4683,N_4619);
and U4920 (N_4920,N_4677,N_4707);
or U4921 (N_4921,N_4789,N_4712);
nand U4922 (N_4922,N_4757,N_4729);
and U4923 (N_4923,N_4724,N_4709);
and U4924 (N_4924,N_4669,N_4656);
or U4925 (N_4925,N_4721,N_4614);
nand U4926 (N_4926,N_4788,N_4754);
nor U4927 (N_4927,N_4650,N_4624);
or U4928 (N_4928,N_4635,N_4797);
or U4929 (N_4929,N_4744,N_4679);
or U4930 (N_4930,N_4660,N_4776);
nor U4931 (N_4931,N_4623,N_4797);
or U4932 (N_4932,N_4733,N_4707);
xnor U4933 (N_4933,N_4741,N_4624);
nand U4934 (N_4934,N_4765,N_4712);
and U4935 (N_4935,N_4741,N_4709);
and U4936 (N_4936,N_4715,N_4792);
or U4937 (N_4937,N_4783,N_4726);
or U4938 (N_4938,N_4769,N_4656);
nand U4939 (N_4939,N_4766,N_4752);
and U4940 (N_4940,N_4666,N_4795);
and U4941 (N_4941,N_4766,N_4735);
nand U4942 (N_4942,N_4617,N_4683);
or U4943 (N_4943,N_4664,N_4777);
nor U4944 (N_4944,N_4699,N_4676);
or U4945 (N_4945,N_4694,N_4797);
or U4946 (N_4946,N_4625,N_4649);
or U4947 (N_4947,N_4787,N_4764);
and U4948 (N_4948,N_4735,N_4632);
and U4949 (N_4949,N_4752,N_4723);
nand U4950 (N_4950,N_4732,N_4662);
nor U4951 (N_4951,N_4606,N_4707);
nand U4952 (N_4952,N_4727,N_4645);
and U4953 (N_4953,N_4604,N_4623);
nand U4954 (N_4954,N_4722,N_4712);
and U4955 (N_4955,N_4680,N_4608);
nand U4956 (N_4956,N_4703,N_4728);
nand U4957 (N_4957,N_4691,N_4746);
and U4958 (N_4958,N_4782,N_4752);
and U4959 (N_4959,N_4739,N_4624);
nor U4960 (N_4960,N_4662,N_4791);
and U4961 (N_4961,N_4681,N_4656);
and U4962 (N_4962,N_4750,N_4628);
and U4963 (N_4963,N_4757,N_4690);
nor U4964 (N_4964,N_4783,N_4648);
and U4965 (N_4965,N_4713,N_4601);
or U4966 (N_4966,N_4735,N_4691);
or U4967 (N_4967,N_4679,N_4695);
nand U4968 (N_4968,N_4661,N_4720);
and U4969 (N_4969,N_4656,N_4731);
nand U4970 (N_4970,N_4689,N_4627);
or U4971 (N_4971,N_4618,N_4648);
nand U4972 (N_4972,N_4616,N_4677);
nand U4973 (N_4973,N_4706,N_4665);
nand U4974 (N_4974,N_4777,N_4785);
and U4975 (N_4975,N_4683,N_4718);
or U4976 (N_4976,N_4707,N_4756);
and U4977 (N_4977,N_4723,N_4732);
nand U4978 (N_4978,N_4631,N_4610);
nor U4979 (N_4979,N_4758,N_4669);
nand U4980 (N_4980,N_4761,N_4710);
nor U4981 (N_4981,N_4632,N_4648);
nand U4982 (N_4982,N_4624,N_4615);
nor U4983 (N_4983,N_4646,N_4752);
or U4984 (N_4984,N_4692,N_4725);
nand U4985 (N_4985,N_4695,N_4722);
and U4986 (N_4986,N_4616,N_4777);
xnor U4987 (N_4987,N_4765,N_4611);
and U4988 (N_4988,N_4727,N_4606);
and U4989 (N_4989,N_4726,N_4655);
nor U4990 (N_4990,N_4696,N_4659);
or U4991 (N_4991,N_4775,N_4751);
or U4992 (N_4992,N_4620,N_4711);
nor U4993 (N_4993,N_4704,N_4724);
nor U4994 (N_4994,N_4635,N_4746);
and U4995 (N_4995,N_4633,N_4600);
or U4996 (N_4996,N_4751,N_4624);
nor U4997 (N_4997,N_4798,N_4731);
nand U4998 (N_4998,N_4647,N_4765);
or U4999 (N_4999,N_4768,N_4656);
and UO_0 (O_0,N_4855,N_4889);
or UO_1 (O_1,N_4993,N_4965);
or UO_2 (O_2,N_4847,N_4968);
and UO_3 (O_3,N_4918,N_4950);
nor UO_4 (O_4,N_4819,N_4902);
or UO_5 (O_5,N_4881,N_4865);
or UO_6 (O_6,N_4888,N_4990);
nand UO_7 (O_7,N_4953,N_4824);
and UO_8 (O_8,N_4930,N_4982);
and UO_9 (O_9,N_4810,N_4923);
nand UO_10 (O_10,N_4894,N_4941);
nor UO_11 (O_11,N_4801,N_4830);
or UO_12 (O_12,N_4875,N_4975);
nand UO_13 (O_13,N_4986,N_4859);
or UO_14 (O_14,N_4878,N_4814);
and UO_15 (O_15,N_4959,N_4999);
and UO_16 (O_16,N_4840,N_4914);
or UO_17 (O_17,N_4987,N_4880);
or UO_18 (O_18,N_4850,N_4940);
nand UO_19 (O_19,N_4861,N_4843);
nand UO_20 (O_20,N_4837,N_4925);
nand UO_21 (O_21,N_4816,N_4802);
and UO_22 (O_22,N_4826,N_4946);
or UO_23 (O_23,N_4863,N_4919);
and UO_24 (O_24,N_4917,N_4967);
and UO_25 (O_25,N_4945,N_4876);
or UO_26 (O_26,N_4927,N_4877);
or UO_27 (O_27,N_4951,N_4901);
xnor UO_28 (O_28,N_4885,N_4961);
or UO_29 (O_29,N_4898,N_4866);
nor UO_30 (O_30,N_4886,N_4872);
nor UO_31 (O_31,N_4893,N_4972);
and UO_32 (O_32,N_4812,N_4883);
nand UO_33 (O_33,N_4807,N_4831);
nand UO_34 (O_34,N_4960,N_4958);
nand UO_35 (O_35,N_4904,N_4813);
and UO_36 (O_36,N_4842,N_4922);
nand UO_37 (O_37,N_4938,N_4935);
nor UO_38 (O_38,N_4803,N_4948);
or UO_39 (O_39,N_4974,N_4949);
nor UO_40 (O_40,N_4907,N_4832);
nand UO_41 (O_41,N_4976,N_4884);
or UO_42 (O_42,N_4827,N_4873);
nand UO_43 (O_43,N_4952,N_4800);
nor UO_44 (O_44,N_4864,N_4882);
and UO_45 (O_45,N_4811,N_4985);
or UO_46 (O_46,N_4834,N_4853);
or UO_47 (O_47,N_4858,N_4908);
or UO_48 (O_48,N_4833,N_4829);
nand UO_49 (O_49,N_4848,N_4869);
nand UO_50 (O_50,N_4804,N_4926);
nand UO_51 (O_51,N_4929,N_4977);
and UO_52 (O_52,N_4969,N_4856);
or UO_53 (O_53,N_4809,N_4934);
nand UO_54 (O_54,N_4921,N_4964);
nor UO_55 (O_55,N_4887,N_4947);
and UO_56 (O_56,N_4933,N_4903);
and UO_57 (O_57,N_4870,N_4896);
nor UO_58 (O_58,N_4944,N_4818);
nand UO_59 (O_59,N_4931,N_4906);
nor UO_60 (O_60,N_4897,N_4808);
and UO_61 (O_61,N_4857,N_4932);
or UO_62 (O_62,N_4900,N_4992);
nand UO_63 (O_63,N_4989,N_4971);
nand UO_64 (O_64,N_4899,N_4913);
nand UO_65 (O_65,N_4956,N_4996);
or UO_66 (O_66,N_4806,N_4963);
or UO_67 (O_67,N_4928,N_4852);
nand UO_68 (O_68,N_4890,N_4871);
nand UO_69 (O_69,N_4912,N_4915);
nand UO_70 (O_70,N_4984,N_4916);
nand UO_71 (O_71,N_4955,N_4942);
or UO_72 (O_72,N_4879,N_4991);
nor UO_73 (O_73,N_4936,N_4980);
and UO_74 (O_74,N_4978,N_4981);
nor UO_75 (O_75,N_4860,N_4805);
nand UO_76 (O_76,N_4892,N_4821);
nand UO_77 (O_77,N_4868,N_4846);
nor UO_78 (O_78,N_4939,N_4994);
nand UO_79 (O_79,N_4844,N_4838);
nor UO_80 (O_80,N_4845,N_4937);
nor UO_81 (O_81,N_4867,N_4943);
nand UO_82 (O_82,N_4995,N_4841);
nor UO_83 (O_83,N_4970,N_4874);
or UO_84 (O_84,N_4839,N_4825);
or UO_85 (O_85,N_4920,N_4905);
nand UO_86 (O_86,N_4998,N_4909);
or UO_87 (O_87,N_4954,N_4822);
nor UO_88 (O_88,N_4817,N_4962);
and UO_89 (O_89,N_4988,N_4895);
nor UO_90 (O_90,N_4966,N_4835);
and UO_91 (O_91,N_4836,N_4891);
nor UO_92 (O_92,N_4849,N_4973);
and UO_93 (O_93,N_4997,N_4823);
nand UO_94 (O_94,N_4862,N_4957);
nand UO_95 (O_95,N_4983,N_4820);
or UO_96 (O_96,N_4924,N_4851);
nand UO_97 (O_97,N_4815,N_4828);
nor UO_98 (O_98,N_4979,N_4911);
nand UO_99 (O_99,N_4854,N_4910);
and UO_100 (O_100,N_4822,N_4945);
and UO_101 (O_101,N_4955,N_4862);
and UO_102 (O_102,N_4916,N_4826);
nand UO_103 (O_103,N_4897,N_4947);
nor UO_104 (O_104,N_4848,N_4824);
or UO_105 (O_105,N_4953,N_4854);
nor UO_106 (O_106,N_4861,N_4840);
and UO_107 (O_107,N_4817,N_4890);
nand UO_108 (O_108,N_4994,N_4864);
nand UO_109 (O_109,N_4961,N_4952);
nor UO_110 (O_110,N_4905,N_4810);
and UO_111 (O_111,N_4933,N_4948);
nor UO_112 (O_112,N_4880,N_4985);
and UO_113 (O_113,N_4881,N_4965);
or UO_114 (O_114,N_4865,N_4800);
and UO_115 (O_115,N_4866,N_4808);
and UO_116 (O_116,N_4898,N_4920);
nand UO_117 (O_117,N_4838,N_4924);
or UO_118 (O_118,N_4819,N_4944);
and UO_119 (O_119,N_4983,N_4962);
and UO_120 (O_120,N_4836,N_4817);
or UO_121 (O_121,N_4812,N_4900);
or UO_122 (O_122,N_4959,N_4816);
nor UO_123 (O_123,N_4843,N_4823);
and UO_124 (O_124,N_4937,N_4859);
or UO_125 (O_125,N_4884,N_4896);
nand UO_126 (O_126,N_4910,N_4944);
and UO_127 (O_127,N_4956,N_4872);
nor UO_128 (O_128,N_4945,N_4932);
and UO_129 (O_129,N_4995,N_4828);
nor UO_130 (O_130,N_4890,N_4832);
nand UO_131 (O_131,N_4923,N_4803);
or UO_132 (O_132,N_4837,N_4955);
nand UO_133 (O_133,N_4849,N_4946);
and UO_134 (O_134,N_4834,N_4975);
nor UO_135 (O_135,N_4880,N_4819);
nand UO_136 (O_136,N_4809,N_4854);
or UO_137 (O_137,N_4865,N_4884);
and UO_138 (O_138,N_4960,N_4979);
or UO_139 (O_139,N_4885,N_4988);
or UO_140 (O_140,N_4941,N_4949);
nor UO_141 (O_141,N_4854,N_4897);
or UO_142 (O_142,N_4869,N_4871);
nor UO_143 (O_143,N_4887,N_4993);
and UO_144 (O_144,N_4948,N_4942);
or UO_145 (O_145,N_4815,N_4810);
nor UO_146 (O_146,N_4888,N_4996);
xnor UO_147 (O_147,N_4984,N_4895);
nor UO_148 (O_148,N_4928,N_4836);
nor UO_149 (O_149,N_4838,N_4853);
nand UO_150 (O_150,N_4913,N_4855);
nor UO_151 (O_151,N_4913,N_4892);
nand UO_152 (O_152,N_4841,N_4891);
or UO_153 (O_153,N_4875,N_4919);
and UO_154 (O_154,N_4959,N_4928);
and UO_155 (O_155,N_4804,N_4961);
and UO_156 (O_156,N_4911,N_4984);
nand UO_157 (O_157,N_4899,N_4992);
nand UO_158 (O_158,N_4868,N_4851);
and UO_159 (O_159,N_4948,N_4970);
xor UO_160 (O_160,N_4912,N_4844);
nand UO_161 (O_161,N_4886,N_4879);
and UO_162 (O_162,N_4985,N_4944);
nand UO_163 (O_163,N_4955,N_4981);
nor UO_164 (O_164,N_4994,N_4855);
and UO_165 (O_165,N_4933,N_4954);
and UO_166 (O_166,N_4934,N_4829);
nor UO_167 (O_167,N_4978,N_4994);
or UO_168 (O_168,N_4888,N_4964);
nand UO_169 (O_169,N_4905,N_4830);
and UO_170 (O_170,N_4879,N_4865);
nor UO_171 (O_171,N_4993,N_4996);
nand UO_172 (O_172,N_4968,N_4809);
nand UO_173 (O_173,N_4976,N_4880);
nand UO_174 (O_174,N_4935,N_4912);
nor UO_175 (O_175,N_4812,N_4859);
or UO_176 (O_176,N_4990,N_4962);
or UO_177 (O_177,N_4881,N_4960);
and UO_178 (O_178,N_4858,N_4818);
and UO_179 (O_179,N_4925,N_4905);
nand UO_180 (O_180,N_4999,N_4853);
nand UO_181 (O_181,N_4844,N_4862);
xor UO_182 (O_182,N_4905,N_4864);
nor UO_183 (O_183,N_4802,N_4998);
nand UO_184 (O_184,N_4848,N_4809);
or UO_185 (O_185,N_4962,N_4934);
and UO_186 (O_186,N_4835,N_4962);
or UO_187 (O_187,N_4921,N_4967);
and UO_188 (O_188,N_4855,N_4961);
and UO_189 (O_189,N_4831,N_4817);
nand UO_190 (O_190,N_4929,N_4988);
or UO_191 (O_191,N_4903,N_4821);
nand UO_192 (O_192,N_4812,N_4930);
nand UO_193 (O_193,N_4821,N_4873);
or UO_194 (O_194,N_4970,N_4957);
or UO_195 (O_195,N_4897,N_4823);
xnor UO_196 (O_196,N_4929,N_4831);
and UO_197 (O_197,N_4975,N_4918);
or UO_198 (O_198,N_4919,N_4981);
or UO_199 (O_199,N_4951,N_4850);
or UO_200 (O_200,N_4931,N_4947);
nand UO_201 (O_201,N_4891,N_4929);
and UO_202 (O_202,N_4849,N_4824);
and UO_203 (O_203,N_4887,N_4841);
and UO_204 (O_204,N_4912,N_4976);
and UO_205 (O_205,N_4880,N_4846);
xor UO_206 (O_206,N_4845,N_4951);
nand UO_207 (O_207,N_4863,N_4916);
nand UO_208 (O_208,N_4954,N_4951);
nand UO_209 (O_209,N_4873,N_4972);
nand UO_210 (O_210,N_4882,N_4973);
and UO_211 (O_211,N_4845,N_4865);
and UO_212 (O_212,N_4925,N_4895);
nand UO_213 (O_213,N_4864,N_4855);
and UO_214 (O_214,N_4892,N_4830);
nor UO_215 (O_215,N_4919,N_4971);
nor UO_216 (O_216,N_4925,N_4958);
nor UO_217 (O_217,N_4997,N_4836);
nor UO_218 (O_218,N_4872,N_4806);
nor UO_219 (O_219,N_4802,N_4918);
nand UO_220 (O_220,N_4833,N_4931);
nand UO_221 (O_221,N_4889,N_4870);
or UO_222 (O_222,N_4801,N_4814);
nor UO_223 (O_223,N_4973,N_4906);
nor UO_224 (O_224,N_4899,N_4830);
or UO_225 (O_225,N_4840,N_4855);
and UO_226 (O_226,N_4917,N_4929);
nand UO_227 (O_227,N_4955,N_4991);
and UO_228 (O_228,N_4882,N_4814);
or UO_229 (O_229,N_4924,N_4932);
xor UO_230 (O_230,N_4859,N_4964);
nor UO_231 (O_231,N_4815,N_4872);
nor UO_232 (O_232,N_4816,N_4860);
nor UO_233 (O_233,N_4847,N_4959);
and UO_234 (O_234,N_4926,N_4924);
nor UO_235 (O_235,N_4961,N_4933);
or UO_236 (O_236,N_4909,N_4851);
nor UO_237 (O_237,N_4975,N_4950);
xnor UO_238 (O_238,N_4956,N_4846);
nor UO_239 (O_239,N_4875,N_4889);
and UO_240 (O_240,N_4868,N_4871);
nor UO_241 (O_241,N_4836,N_4951);
nor UO_242 (O_242,N_4921,N_4914);
or UO_243 (O_243,N_4879,N_4952);
or UO_244 (O_244,N_4973,N_4805);
and UO_245 (O_245,N_4875,N_4819);
nor UO_246 (O_246,N_4943,N_4835);
or UO_247 (O_247,N_4994,N_4875);
nand UO_248 (O_248,N_4886,N_4983);
and UO_249 (O_249,N_4840,N_4823);
nor UO_250 (O_250,N_4854,N_4988);
xnor UO_251 (O_251,N_4802,N_4838);
nor UO_252 (O_252,N_4834,N_4991);
or UO_253 (O_253,N_4856,N_4911);
nor UO_254 (O_254,N_4807,N_4941);
or UO_255 (O_255,N_4822,N_4868);
or UO_256 (O_256,N_4831,N_4952);
nor UO_257 (O_257,N_4834,N_4949);
nand UO_258 (O_258,N_4861,N_4996);
nand UO_259 (O_259,N_4970,N_4812);
or UO_260 (O_260,N_4955,N_4938);
nor UO_261 (O_261,N_4955,N_4860);
or UO_262 (O_262,N_4991,N_4880);
nor UO_263 (O_263,N_4960,N_4948);
nor UO_264 (O_264,N_4900,N_4980);
and UO_265 (O_265,N_4894,N_4825);
nor UO_266 (O_266,N_4948,N_4843);
nor UO_267 (O_267,N_4995,N_4925);
or UO_268 (O_268,N_4960,N_4965);
nor UO_269 (O_269,N_4817,N_4984);
or UO_270 (O_270,N_4982,N_4991);
nor UO_271 (O_271,N_4959,N_4865);
or UO_272 (O_272,N_4943,N_4884);
nor UO_273 (O_273,N_4850,N_4870);
nand UO_274 (O_274,N_4870,N_4946);
nand UO_275 (O_275,N_4978,N_4953);
and UO_276 (O_276,N_4873,N_4863);
or UO_277 (O_277,N_4895,N_4959);
nand UO_278 (O_278,N_4950,N_4844);
and UO_279 (O_279,N_4903,N_4947);
nand UO_280 (O_280,N_4867,N_4894);
nor UO_281 (O_281,N_4861,N_4991);
nand UO_282 (O_282,N_4955,N_4863);
and UO_283 (O_283,N_4841,N_4881);
and UO_284 (O_284,N_4932,N_4931);
and UO_285 (O_285,N_4829,N_4991);
or UO_286 (O_286,N_4977,N_4837);
and UO_287 (O_287,N_4884,N_4859);
or UO_288 (O_288,N_4966,N_4920);
nand UO_289 (O_289,N_4888,N_4953);
nor UO_290 (O_290,N_4845,N_4936);
nor UO_291 (O_291,N_4886,N_4887);
or UO_292 (O_292,N_4848,N_4852);
and UO_293 (O_293,N_4837,N_4828);
nand UO_294 (O_294,N_4847,N_4803);
nor UO_295 (O_295,N_4847,N_4815);
nand UO_296 (O_296,N_4875,N_4849);
and UO_297 (O_297,N_4980,N_4967);
and UO_298 (O_298,N_4840,N_4900);
and UO_299 (O_299,N_4856,N_4934);
nand UO_300 (O_300,N_4931,N_4846);
nand UO_301 (O_301,N_4895,N_4831);
nor UO_302 (O_302,N_4978,N_4817);
nand UO_303 (O_303,N_4988,N_4956);
nor UO_304 (O_304,N_4886,N_4889);
or UO_305 (O_305,N_4947,N_4921);
xnor UO_306 (O_306,N_4958,N_4919);
nand UO_307 (O_307,N_4978,N_4833);
nor UO_308 (O_308,N_4850,N_4943);
or UO_309 (O_309,N_4804,N_4824);
nor UO_310 (O_310,N_4986,N_4987);
nor UO_311 (O_311,N_4972,N_4919);
nand UO_312 (O_312,N_4912,N_4885);
nand UO_313 (O_313,N_4854,N_4841);
nand UO_314 (O_314,N_4869,N_4944);
nor UO_315 (O_315,N_4885,N_4994);
or UO_316 (O_316,N_4803,N_4914);
nand UO_317 (O_317,N_4977,N_4830);
nor UO_318 (O_318,N_4971,N_4886);
or UO_319 (O_319,N_4800,N_4936);
nand UO_320 (O_320,N_4940,N_4913);
or UO_321 (O_321,N_4986,N_4808);
nand UO_322 (O_322,N_4886,N_4934);
and UO_323 (O_323,N_4934,N_4854);
nand UO_324 (O_324,N_4820,N_4898);
and UO_325 (O_325,N_4894,N_4818);
nor UO_326 (O_326,N_4835,N_4808);
nor UO_327 (O_327,N_4855,N_4827);
and UO_328 (O_328,N_4975,N_4893);
nor UO_329 (O_329,N_4941,N_4994);
nor UO_330 (O_330,N_4945,N_4819);
nand UO_331 (O_331,N_4927,N_4936);
and UO_332 (O_332,N_4910,N_4975);
nor UO_333 (O_333,N_4921,N_4884);
and UO_334 (O_334,N_4867,N_4883);
nand UO_335 (O_335,N_4936,N_4902);
or UO_336 (O_336,N_4971,N_4819);
nor UO_337 (O_337,N_4951,N_4990);
or UO_338 (O_338,N_4989,N_4985);
nand UO_339 (O_339,N_4997,N_4982);
and UO_340 (O_340,N_4899,N_4911);
or UO_341 (O_341,N_4892,N_4801);
nand UO_342 (O_342,N_4971,N_4951);
or UO_343 (O_343,N_4890,N_4962);
nor UO_344 (O_344,N_4945,N_4866);
and UO_345 (O_345,N_4808,N_4862);
or UO_346 (O_346,N_4841,N_4839);
and UO_347 (O_347,N_4916,N_4950);
nand UO_348 (O_348,N_4982,N_4847);
nand UO_349 (O_349,N_4905,N_4869);
nand UO_350 (O_350,N_4979,N_4889);
nand UO_351 (O_351,N_4908,N_4876);
or UO_352 (O_352,N_4891,N_4914);
or UO_353 (O_353,N_4913,N_4843);
and UO_354 (O_354,N_4815,N_4879);
nand UO_355 (O_355,N_4942,N_4891);
nor UO_356 (O_356,N_4839,N_4808);
nor UO_357 (O_357,N_4834,N_4960);
nor UO_358 (O_358,N_4907,N_4914);
and UO_359 (O_359,N_4988,N_4871);
or UO_360 (O_360,N_4898,N_4899);
nand UO_361 (O_361,N_4817,N_4977);
and UO_362 (O_362,N_4978,N_4898);
or UO_363 (O_363,N_4870,N_4881);
nor UO_364 (O_364,N_4961,N_4957);
and UO_365 (O_365,N_4974,N_4991);
and UO_366 (O_366,N_4938,N_4902);
and UO_367 (O_367,N_4869,N_4971);
or UO_368 (O_368,N_4874,N_4869);
nand UO_369 (O_369,N_4805,N_4835);
nor UO_370 (O_370,N_4989,N_4910);
nor UO_371 (O_371,N_4948,N_4854);
and UO_372 (O_372,N_4868,N_4949);
nand UO_373 (O_373,N_4809,N_4941);
nand UO_374 (O_374,N_4986,N_4800);
nand UO_375 (O_375,N_4866,N_4910);
and UO_376 (O_376,N_4879,N_4945);
nand UO_377 (O_377,N_4905,N_4842);
or UO_378 (O_378,N_4947,N_4806);
nor UO_379 (O_379,N_4850,N_4835);
and UO_380 (O_380,N_4973,N_4812);
or UO_381 (O_381,N_4890,N_4827);
or UO_382 (O_382,N_4940,N_4906);
nor UO_383 (O_383,N_4815,N_4980);
nor UO_384 (O_384,N_4982,N_4910);
nand UO_385 (O_385,N_4831,N_4838);
or UO_386 (O_386,N_4979,N_4806);
nor UO_387 (O_387,N_4836,N_4973);
and UO_388 (O_388,N_4921,N_4990);
or UO_389 (O_389,N_4979,N_4871);
and UO_390 (O_390,N_4943,N_4921);
or UO_391 (O_391,N_4927,N_4845);
nand UO_392 (O_392,N_4928,N_4872);
or UO_393 (O_393,N_4822,N_4890);
nor UO_394 (O_394,N_4936,N_4868);
or UO_395 (O_395,N_4812,N_4995);
nor UO_396 (O_396,N_4825,N_4941);
or UO_397 (O_397,N_4831,N_4933);
nand UO_398 (O_398,N_4950,N_4945);
nand UO_399 (O_399,N_4991,N_4996);
and UO_400 (O_400,N_4944,N_4857);
and UO_401 (O_401,N_4928,N_4939);
and UO_402 (O_402,N_4949,N_4814);
and UO_403 (O_403,N_4807,N_4977);
and UO_404 (O_404,N_4882,N_4808);
or UO_405 (O_405,N_4964,N_4829);
or UO_406 (O_406,N_4884,N_4922);
nand UO_407 (O_407,N_4893,N_4832);
or UO_408 (O_408,N_4843,N_4972);
and UO_409 (O_409,N_4938,N_4956);
nand UO_410 (O_410,N_4945,N_4906);
and UO_411 (O_411,N_4994,N_4956);
and UO_412 (O_412,N_4942,N_4833);
or UO_413 (O_413,N_4966,N_4820);
or UO_414 (O_414,N_4820,N_4865);
or UO_415 (O_415,N_4815,N_4808);
nand UO_416 (O_416,N_4807,N_4935);
nand UO_417 (O_417,N_4885,N_4967);
nor UO_418 (O_418,N_4889,N_4967);
or UO_419 (O_419,N_4896,N_4813);
nand UO_420 (O_420,N_4808,N_4956);
xnor UO_421 (O_421,N_4886,N_4892);
or UO_422 (O_422,N_4910,N_4977);
and UO_423 (O_423,N_4890,N_4915);
and UO_424 (O_424,N_4838,N_4934);
or UO_425 (O_425,N_4862,N_4998);
or UO_426 (O_426,N_4929,N_4822);
nor UO_427 (O_427,N_4887,N_4849);
or UO_428 (O_428,N_4866,N_4823);
and UO_429 (O_429,N_4882,N_4899);
or UO_430 (O_430,N_4855,N_4979);
or UO_431 (O_431,N_4964,N_4896);
nor UO_432 (O_432,N_4927,N_4861);
or UO_433 (O_433,N_4866,N_4939);
or UO_434 (O_434,N_4902,N_4909);
nor UO_435 (O_435,N_4830,N_4822);
nand UO_436 (O_436,N_4887,N_4813);
nor UO_437 (O_437,N_4966,N_4977);
or UO_438 (O_438,N_4835,N_4979);
nand UO_439 (O_439,N_4870,N_4908);
nand UO_440 (O_440,N_4841,N_4981);
xnor UO_441 (O_441,N_4820,N_4887);
or UO_442 (O_442,N_4852,N_4866);
nor UO_443 (O_443,N_4922,N_4872);
and UO_444 (O_444,N_4973,N_4861);
and UO_445 (O_445,N_4916,N_4856);
or UO_446 (O_446,N_4842,N_4843);
and UO_447 (O_447,N_4842,N_4867);
or UO_448 (O_448,N_4819,N_4986);
or UO_449 (O_449,N_4921,N_4984);
and UO_450 (O_450,N_4828,N_4961);
nor UO_451 (O_451,N_4980,N_4866);
and UO_452 (O_452,N_4880,N_4872);
nor UO_453 (O_453,N_4883,N_4837);
nand UO_454 (O_454,N_4815,N_4970);
or UO_455 (O_455,N_4937,N_4919);
nor UO_456 (O_456,N_4898,N_4810);
and UO_457 (O_457,N_4959,N_4962);
nor UO_458 (O_458,N_4900,N_4833);
and UO_459 (O_459,N_4916,N_4913);
nand UO_460 (O_460,N_4907,N_4928);
nand UO_461 (O_461,N_4980,N_4928);
or UO_462 (O_462,N_4800,N_4966);
nand UO_463 (O_463,N_4986,N_4810);
or UO_464 (O_464,N_4855,N_4890);
and UO_465 (O_465,N_4883,N_4819);
nand UO_466 (O_466,N_4952,N_4818);
nor UO_467 (O_467,N_4892,N_4800);
nand UO_468 (O_468,N_4928,N_4869);
or UO_469 (O_469,N_4923,N_4834);
and UO_470 (O_470,N_4849,N_4929);
or UO_471 (O_471,N_4816,N_4853);
nor UO_472 (O_472,N_4961,N_4872);
nor UO_473 (O_473,N_4997,N_4834);
or UO_474 (O_474,N_4844,N_4814);
nor UO_475 (O_475,N_4846,N_4863);
and UO_476 (O_476,N_4971,N_4820);
and UO_477 (O_477,N_4997,N_4852);
or UO_478 (O_478,N_4939,N_4892);
nand UO_479 (O_479,N_4992,N_4912);
and UO_480 (O_480,N_4950,N_4818);
nand UO_481 (O_481,N_4980,N_4998);
and UO_482 (O_482,N_4818,N_4903);
or UO_483 (O_483,N_4906,N_4859);
nor UO_484 (O_484,N_4894,N_4996);
and UO_485 (O_485,N_4973,N_4904);
nor UO_486 (O_486,N_4806,N_4902);
nand UO_487 (O_487,N_4973,N_4991);
nor UO_488 (O_488,N_4915,N_4808);
nor UO_489 (O_489,N_4996,N_4887);
nand UO_490 (O_490,N_4865,N_4919);
or UO_491 (O_491,N_4875,N_4878);
nand UO_492 (O_492,N_4921,N_4920);
and UO_493 (O_493,N_4835,N_4846);
and UO_494 (O_494,N_4818,N_4875);
nor UO_495 (O_495,N_4981,N_4838);
or UO_496 (O_496,N_4832,N_4833);
nor UO_497 (O_497,N_4894,N_4960);
and UO_498 (O_498,N_4903,N_4922);
or UO_499 (O_499,N_4978,N_4931);
or UO_500 (O_500,N_4902,N_4997);
nor UO_501 (O_501,N_4928,N_4997);
or UO_502 (O_502,N_4909,N_4951);
or UO_503 (O_503,N_4905,N_4848);
and UO_504 (O_504,N_4873,N_4881);
nor UO_505 (O_505,N_4968,N_4951);
and UO_506 (O_506,N_4945,N_4953);
and UO_507 (O_507,N_4972,N_4882);
and UO_508 (O_508,N_4953,N_4837);
nor UO_509 (O_509,N_4866,N_4807);
and UO_510 (O_510,N_4948,N_4861);
and UO_511 (O_511,N_4896,N_4887);
and UO_512 (O_512,N_4869,N_4875);
nor UO_513 (O_513,N_4969,N_4814);
or UO_514 (O_514,N_4932,N_4843);
and UO_515 (O_515,N_4945,N_4816);
and UO_516 (O_516,N_4834,N_4940);
nor UO_517 (O_517,N_4818,N_4812);
nor UO_518 (O_518,N_4950,N_4928);
nand UO_519 (O_519,N_4817,N_4931);
nor UO_520 (O_520,N_4978,N_4846);
nand UO_521 (O_521,N_4841,N_4884);
nand UO_522 (O_522,N_4938,N_4996);
nor UO_523 (O_523,N_4982,N_4813);
and UO_524 (O_524,N_4959,N_4844);
and UO_525 (O_525,N_4843,N_4820);
nor UO_526 (O_526,N_4973,N_4985);
or UO_527 (O_527,N_4853,N_4940);
and UO_528 (O_528,N_4800,N_4914);
and UO_529 (O_529,N_4839,N_4906);
or UO_530 (O_530,N_4919,N_4846);
nor UO_531 (O_531,N_4929,N_4926);
and UO_532 (O_532,N_4935,N_4861);
or UO_533 (O_533,N_4822,N_4978);
nand UO_534 (O_534,N_4918,N_4824);
or UO_535 (O_535,N_4920,N_4886);
nand UO_536 (O_536,N_4978,N_4811);
nor UO_537 (O_537,N_4958,N_4927);
and UO_538 (O_538,N_4949,N_4815);
xnor UO_539 (O_539,N_4892,N_4955);
nor UO_540 (O_540,N_4907,N_4967);
nand UO_541 (O_541,N_4882,N_4836);
and UO_542 (O_542,N_4989,N_4953);
nand UO_543 (O_543,N_4947,N_4807);
nor UO_544 (O_544,N_4936,N_4813);
and UO_545 (O_545,N_4819,N_4829);
nand UO_546 (O_546,N_4949,N_4936);
nor UO_547 (O_547,N_4948,N_4846);
nor UO_548 (O_548,N_4809,N_4920);
or UO_549 (O_549,N_4971,N_4953);
or UO_550 (O_550,N_4883,N_4829);
nand UO_551 (O_551,N_4964,N_4833);
and UO_552 (O_552,N_4840,N_4853);
and UO_553 (O_553,N_4997,N_4866);
or UO_554 (O_554,N_4863,N_4901);
and UO_555 (O_555,N_4981,N_4974);
nand UO_556 (O_556,N_4942,N_4940);
nand UO_557 (O_557,N_4945,N_4878);
xor UO_558 (O_558,N_4869,N_4926);
and UO_559 (O_559,N_4886,N_4996);
and UO_560 (O_560,N_4854,N_4922);
nor UO_561 (O_561,N_4841,N_4821);
xor UO_562 (O_562,N_4917,N_4956);
or UO_563 (O_563,N_4906,N_4820);
nand UO_564 (O_564,N_4882,N_4893);
and UO_565 (O_565,N_4992,N_4930);
xnor UO_566 (O_566,N_4821,N_4869);
nor UO_567 (O_567,N_4966,N_4830);
and UO_568 (O_568,N_4830,N_4843);
nor UO_569 (O_569,N_4926,N_4856);
and UO_570 (O_570,N_4990,N_4960);
nor UO_571 (O_571,N_4948,N_4926);
and UO_572 (O_572,N_4974,N_4805);
nand UO_573 (O_573,N_4970,N_4859);
nor UO_574 (O_574,N_4813,N_4808);
or UO_575 (O_575,N_4808,N_4887);
nor UO_576 (O_576,N_4870,N_4864);
nor UO_577 (O_577,N_4848,N_4920);
or UO_578 (O_578,N_4899,N_4960);
and UO_579 (O_579,N_4868,N_4844);
and UO_580 (O_580,N_4818,N_4962);
and UO_581 (O_581,N_4912,N_4902);
nand UO_582 (O_582,N_4972,N_4945);
and UO_583 (O_583,N_4879,N_4841);
or UO_584 (O_584,N_4995,N_4857);
nand UO_585 (O_585,N_4957,N_4885);
or UO_586 (O_586,N_4923,N_4947);
xor UO_587 (O_587,N_4890,N_4807);
nor UO_588 (O_588,N_4906,N_4966);
nor UO_589 (O_589,N_4983,N_4865);
nand UO_590 (O_590,N_4900,N_4835);
xor UO_591 (O_591,N_4810,N_4933);
nand UO_592 (O_592,N_4811,N_4980);
and UO_593 (O_593,N_4996,N_4962);
nor UO_594 (O_594,N_4911,N_4884);
nand UO_595 (O_595,N_4990,N_4873);
and UO_596 (O_596,N_4935,N_4867);
or UO_597 (O_597,N_4998,N_4825);
and UO_598 (O_598,N_4912,N_4947);
nand UO_599 (O_599,N_4859,N_4803);
or UO_600 (O_600,N_4959,N_4822);
nand UO_601 (O_601,N_4950,N_4843);
nand UO_602 (O_602,N_4839,N_4838);
nand UO_603 (O_603,N_4844,N_4923);
nand UO_604 (O_604,N_4836,N_4909);
nor UO_605 (O_605,N_4989,N_4904);
nand UO_606 (O_606,N_4809,N_4963);
and UO_607 (O_607,N_4999,N_4872);
nor UO_608 (O_608,N_4953,N_4821);
nor UO_609 (O_609,N_4978,N_4977);
or UO_610 (O_610,N_4848,N_4966);
or UO_611 (O_611,N_4837,N_4808);
nand UO_612 (O_612,N_4903,N_4987);
nand UO_613 (O_613,N_4955,N_4957);
and UO_614 (O_614,N_4950,N_4805);
and UO_615 (O_615,N_4876,N_4934);
and UO_616 (O_616,N_4972,N_4952);
and UO_617 (O_617,N_4839,N_4820);
or UO_618 (O_618,N_4980,N_4897);
xnor UO_619 (O_619,N_4899,N_4977);
nor UO_620 (O_620,N_4941,N_4987);
or UO_621 (O_621,N_4880,N_4958);
and UO_622 (O_622,N_4866,N_4877);
nor UO_623 (O_623,N_4826,N_4967);
nor UO_624 (O_624,N_4973,N_4824);
nor UO_625 (O_625,N_4866,N_4893);
and UO_626 (O_626,N_4894,N_4834);
xnor UO_627 (O_627,N_4824,N_4811);
and UO_628 (O_628,N_4979,N_4867);
or UO_629 (O_629,N_4905,N_4961);
or UO_630 (O_630,N_4920,N_4934);
nand UO_631 (O_631,N_4884,N_4993);
nand UO_632 (O_632,N_4979,N_4987);
nand UO_633 (O_633,N_4815,N_4862);
nand UO_634 (O_634,N_4941,N_4958);
nor UO_635 (O_635,N_4900,N_4908);
nand UO_636 (O_636,N_4907,N_4837);
or UO_637 (O_637,N_4856,N_4889);
and UO_638 (O_638,N_4963,N_4830);
or UO_639 (O_639,N_4974,N_4975);
nor UO_640 (O_640,N_4992,N_4988);
or UO_641 (O_641,N_4886,N_4919);
nand UO_642 (O_642,N_4811,N_4838);
and UO_643 (O_643,N_4954,N_4961);
and UO_644 (O_644,N_4809,N_4865);
nor UO_645 (O_645,N_4908,N_4910);
and UO_646 (O_646,N_4953,N_4999);
nand UO_647 (O_647,N_4924,N_4894);
or UO_648 (O_648,N_4965,N_4901);
or UO_649 (O_649,N_4954,N_4967);
or UO_650 (O_650,N_4834,N_4941);
nor UO_651 (O_651,N_4887,N_4899);
or UO_652 (O_652,N_4993,N_4816);
and UO_653 (O_653,N_4822,N_4851);
nand UO_654 (O_654,N_4830,N_4850);
and UO_655 (O_655,N_4828,N_4980);
nor UO_656 (O_656,N_4826,N_4888);
nand UO_657 (O_657,N_4955,N_4811);
or UO_658 (O_658,N_4926,N_4992);
nand UO_659 (O_659,N_4891,N_4973);
nor UO_660 (O_660,N_4979,N_4879);
or UO_661 (O_661,N_4920,N_4813);
nor UO_662 (O_662,N_4844,N_4807);
nor UO_663 (O_663,N_4802,N_4972);
nor UO_664 (O_664,N_4895,N_4888);
nor UO_665 (O_665,N_4881,N_4885);
and UO_666 (O_666,N_4882,N_4834);
and UO_667 (O_667,N_4829,N_4860);
and UO_668 (O_668,N_4926,N_4946);
nor UO_669 (O_669,N_4956,N_4948);
nand UO_670 (O_670,N_4916,N_4876);
nor UO_671 (O_671,N_4911,N_4880);
nand UO_672 (O_672,N_4816,N_4820);
and UO_673 (O_673,N_4928,N_4876);
or UO_674 (O_674,N_4831,N_4908);
or UO_675 (O_675,N_4958,N_4837);
and UO_676 (O_676,N_4971,N_4899);
and UO_677 (O_677,N_4989,N_4837);
and UO_678 (O_678,N_4906,N_4900);
or UO_679 (O_679,N_4975,N_4958);
nor UO_680 (O_680,N_4830,N_4970);
and UO_681 (O_681,N_4867,N_4940);
nand UO_682 (O_682,N_4903,N_4904);
nand UO_683 (O_683,N_4931,N_4900);
and UO_684 (O_684,N_4807,N_4812);
nand UO_685 (O_685,N_4828,N_4846);
nor UO_686 (O_686,N_4941,N_4824);
or UO_687 (O_687,N_4986,N_4897);
and UO_688 (O_688,N_4800,N_4838);
or UO_689 (O_689,N_4815,N_4841);
nand UO_690 (O_690,N_4896,N_4986);
nor UO_691 (O_691,N_4957,N_4801);
and UO_692 (O_692,N_4892,N_4954);
nand UO_693 (O_693,N_4941,N_4983);
and UO_694 (O_694,N_4808,N_4852);
nor UO_695 (O_695,N_4957,N_4809);
or UO_696 (O_696,N_4870,N_4950);
nor UO_697 (O_697,N_4977,N_4847);
and UO_698 (O_698,N_4894,N_4808);
or UO_699 (O_699,N_4959,N_4883);
or UO_700 (O_700,N_4804,N_4848);
nor UO_701 (O_701,N_4989,N_4968);
or UO_702 (O_702,N_4812,N_4879);
or UO_703 (O_703,N_4896,N_4906);
and UO_704 (O_704,N_4852,N_4938);
nor UO_705 (O_705,N_4821,N_4833);
nor UO_706 (O_706,N_4972,N_4879);
nand UO_707 (O_707,N_4836,N_4806);
or UO_708 (O_708,N_4813,N_4939);
or UO_709 (O_709,N_4912,N_4920);
nand UO_710 (O_710,N_4960,N_4967);
nor UO_711 (O_711,N_4978,N_4839);
and UO_712 (O_712,N_4830,N_4813);
or UO_713 (O_713,N_4814,N_4921);
and UO_714 (O_714,N_4924,N_4995);
and UO_715 (O_715,N_4909,N_4922);
and UO_716 (O_716,N_4918,N_4925);
and UO_717 (O_717,N_4975,N_4968);
nand UO_718 (O_718,N_4998,N_4822);
or UO_719 (O_719,N_4885,N_4889);
nor UO_720 (O_720,N_4826,N_4840);
nor UO_721 (O_721,N_4847,N_4886);
or UO_722 (O_722,N_4993,N_4925);
nand UO_723 (O_723,N_4940,N_4960);
or UO_724 (O_724,N_4832,N_4808);
nand UO_725 (O_725,N_4834,N_4896);
nand UO_726 (O_726,N_4954,N_4920);
nor UO_727 (O_727,N_4966,N_4869);
and UO_728 (O_728,N_4827,N_4809);
or UO_729 (O_729,N_4987,N_4815);
nand UO_730 (O_730,N_4960,N_4849);
or UO_731 (O_731,N_4951,N_4840);
xor UO_732 (O_732,N_4949,N_4914);
or UO_733 (O_733,N_4832,N_4996);
and UO_734 (O_734,N_4935,N_4992);
nand UO_735 (O_735,N_4838,N_4861);
nand UO_736 (O_736,N_4939,N_4969);
and UO_737 (O_737,N_4862,N_4893);
nor UO_738 (O_738,N_4816,N_4893);
nor UO_739 (O_739,N_4966,N_4839);
or UO_740 (O_740,N_4891,N_4964);
and UO_741 (O_741,N_4937,N_4821);
nand UO_742 (O_742,N_4849,N_4977);
nor UO_743 (O_743,N_4891,N_4866);
nand UO_744 (O_744,N_4974,N_4927);
nand UO_745 (O_745,N_4957,N_4889);
or UO_746 (O_746,N_4958,N_4910);
or UO_747 (O_747,N_4827,N_4936);
or UO_748 (O_748,N_4878,N_4957);
nor UO_749 (O_749,N_4873,N_4801);
or UO_750 (O_750,N_4875,N_4811);
or UO_751 (O_751,N_4814,N_4970);
nor UO_752 (O_752,N_4985,N_4822);
and UO_753 (O_753,N_4868,N_4903);
and UO_754 (O_754,N_4901,N_4957);
and UO_755 (O_755,N_4838,N_4945);
and UO_756 (O_756,N_4918,N_4806);
and UO_757 (O_757,N_4935,N_4983);
and UO_758 (O_758,N_4951,N_4979);
and UO_759 (O_759,N_4835,N_4961);
or UO_760 (O_760,N_4911,N_4956);
and UO_761 (O_761,N_4849,N_4831);
and UO_762 (O_762,N_4978,N_4951);
and UO_763 (O_763,N_4937,N_4817);
or UO_764 (O_764,N_4952,N_4856);
nor UO_765 (O_765,N_4958,N_4883);
and UO_766 (O_766,N_4848,N_4896);
and UO_767 (O_767,N_4908,N_4907);
and UO_768 (O_768,N_4826,N_4951);
nor UO_769 (O_769,N_4903,N_4996);
and UO_770 (O_770,N_4883,N_4912);
nand UO_771 (O_771,N_4852,N_4967);
or UO_772 (O_772,N_4944,N_4826);
nor UO_773 (O_773,N_4986,N_4829);
or UO_774 (O_774,N_4952,N_4845);
or UO_775 (O_775,N_4991,N_4891);
nor UO_776 (O_776,N_4929,N_4997);
or UO_777 (O_777,N_4817,N_4905);
or UO_778 (O_778,N_4856,N_4903);
or UO_779 (O_779,N_4990,N_4837);
nand UO_780 (O_780,N_4970,N_4845);
nand UO_781 (O_781,N_4911,N_4813);
nor UO_782 (O_782,N_4937,N_4938);
or UO_783 (O_783,N_4839,N_4947);
nor UO_784 (O_784,N_4920,N_4950);
or UO_785 (O_785,N_4975,N_4936);
and UO_786 (O_786,N_4976,N_4902);
or UO_787 (O_787,N_4947,N_4812);
nand UO_788 (O_788,N_4812,N_4835);
or UO_789 (O_789,N_4915,N_4979);
nor UO_790 (O_790,N_4908,N_4812);
nand UO_791 (O_791,N_4955,N_4903);
nor UO_792 (O_792,N_4854,N_4923);
nor UO_793 (O_793,N_4937,N_4861);
and UO_794 (O_794,N_4914,N_4819);
or UO_795 (O_795,N_4889,N_4912);
nor UO_796 (O_796,N_4871,N_4831);
nand UO_797 (O_797,N_4970,N_4846);
nand UO_798 (O_798,N_4863,N_4903);
or UO_799 (O_799,N_4833,N_4839);
nand UO_800 (O_800,N_4898,N_4993);
or UO_801 (O_801,N_4877,N_4880);
or UO_802 (O_802,N_4928,N_4908);
nand UO_803 (O_803,N_4968,N_4811);
or UO_804 (O_804,N_4938,N_4839);
nor UO_805 (O_805,N_4811,N_4823);
nor UO_806 (O_806,N_4858,N_4884);
nor UO_807 (O_807,N_4907,N_4965);
nand UO_808 (O_808,N_4860,N_4971);
or UO_809 (O_809,N_4834,N_4867);
nand UO_810 (O_810,N_4838,N_4840);
or UO_811 (O_811,N_4840,N_4865);
xnor UO_812 (O_812,N_4901,N_4882);
nand UO_813 (O_813,N_4827,N_4989);
nor UO_814 (O_814,N_4902,N_4832);
or UO_815 (O_815,N_4945,N_4883);
and UO_816 (O_816,N_4819,N_4923);
and UO_817 (O_817,N_4933,N_4847);
nor UO_818 (O_818,N_4940,N_4985);
or UO_819 (O_819,N_4835,N_4911);
and UO_820 (O_820,N_4973,N_4948);
nor UO_821 (O_821,N_4989,N_4800);
and UO_822 (O_822,N_4869,N_4910);
xor UO_823 (O_823,N_4921,N_4833);
nand UO_824 (O_824,N_4938,N_4993);
or UO_825 (O_825,N_4805,N_4801);
and UO_826 (O_826,N_4896,N_4927);
nand UO_827 (O_827,N_4809,N_4978);
nand UO_828 (O_828,N_4993,N_4859);
nand UO_829 (O_829,N_4909,N_4840);
nor UO_830 (O_830,N_4952,N_4911);
or UO_831 (O_831,N_4821,N_4850);
or UO_832 (O_832,N_4813,N_4811);
or UO_833 (O_833,N_4833,N_4819);
nand UO_834 (O_834,N_4888,N_4907);
nor UO_835 (O_835,N_4881,N_4980);
nor UO_836 (O_836,N_4911,N_4977);
or UO_837 (O_837,N_4835,N_4928);
nor UO_838 (O_838,N_4817,N_4822);
and UO_839 (O_839,N_4996,N_4896);
and UO_840 (O_840,N_4937,N_4822);
nor UO_841 (O_841,N_4979,N_4949);
nand UO_842 (O_842,N_4930,N_4987);
and UO_843 (O_843,N_4830,N_4964);
nand UO_844 (O_844,N_4972,N_4866);
nor UO_845 (O_845,N_4884,N_4995);
or UO_846 (O_846,N_4935,N_4864);
xnor UO_847 (O_847,N_4985,N_4807);
nand UO_848 (O_848,N_4826,N_4958);
nand UO_849 (O_849,N_4937,N_4904);
nand UO_850 (O_850,N_4920,N_4973);
nor UO_851 (O_851,N_4974,N_4875);
nand UO_852 (O_852,N_4914,N_4918);
nor UO_853 (O_853,N_4823,N_4955);
xor UO_854 (O_854,N_4891,N_4875);
or UO_855 (O_855,N_4887,N_4822);
nor UO_856 (O_856,N_4815,N_4889);
nor UO_857 (O_857,N_4836,N_4981);
and UO_858 (O_858,N_4801,N_4966);
xor UO_859 (O_859,N_4972,N_4969);
or UO_860 (O_860,N_4944,N_4845);
and UO_861 (O_861,N_4914,N_4815);
nand UO_862 (O_862,N_4996,N_4807);
nand UO_863 (O_863,N_4910,N_4852);
or UO_864 (O_864,N_4979,N_4810);
nand UO_865 (O_865,N_4904,N_4990);
and UO_866 (O_866,N_4872,N_4855);
nand UO_867 (O_867,N_4803,N_4990);
or UO_868 (O_868,N_4803,N_4904);
or UO_869 (O_869,N_4945,N_4835);
or UO_870 (O_870,N_4977,N_4879);
nor UO_871 (O_871,N_4947,N_4964);
or UO_872 (O_872,N_4972,N_4921);
nor UO_873 (O_873,N_4921,N_4980);
nor UO_874 (O_874,N_4985,N_4848);
and UO_875 (O_875,N_4923,N_4870);
nand UO_876 (O_876,N_4927,N_4852);
nor UO_877 (O_877,N_4817,N_4998);
nand UO_878 (O_878,N_4926,N_4985);
or UO_879 (O_879,N_4857,N_4937);
xor UO_880 (O_880,N_4861,N_4862);
nand UO_881 (O_881,N_4986,N_4849);
nor UO_882 (O_882,N_4938,N_4995);
or UO_883 (O_883,N_4825,N_4952);
nor UO_884 (O_884,N_4884,N_4989);
or UO_885 (O_885,N_4882,N_4846);
and UO_886 (O_886,N_4857,N_4955);
and UO_887 (O_887,N_4938,N_4985);
or UO_888 (O_888,N_4998,N_4948);
nor UO_889 (O_889,N_4871,N_4963);
or UO_890 (O_890,N_4897,N_4853);
and UO_891 (O_891,N_4825,N_4830);
or UO_892 (O_892,N_4931,N_4869);
or UO_893 (O_893,N_4917,N_4941);
or UO_894 (O_894,N_4959,N_4837);
nor UO_895 (O_895,N_4899,N_4815);
nor UO_896 (O_896,N_4914,N_4829);
nor UO_897 (O_897,N_4973,N_4876);
nand UO_898 (O_898,N_4921,N_4844);
or UO_899 (O_899,N_4942,N_4910);
and UO_900 (O_900,N_4806,N_4851);
or UO_901 (O_901,N_4921,N_4904);
nor UO_902 (O_902,N_4826,N_4816);
nor UO_903 (O_903,N_4826,N_4857);
nor UO_904 (O_904,N_4986,N_4970);
nand UO_905 (O_905,N_4817,N_4832);
nor UO_906 (O_906,N_4950,N_4882);
and UO_907 (O_907,N_4973,N_4809);
nand UO_908 (O_908,N_4893,N_4835);
nor UO_909 (O_909,N_4859,N_4874);
or UO_910 (O_910,N_4843,N_4921);
nand UO_911 (O_911,N_4867,N_4874);
or UO_912 (O_912,N_4967,N_4872);
or UO_913 (O_913,N_4993,N_4948);
nor UO_914 (O_914,N_4850,N_4814);
and UO_915 (O_915,N_4834,N_4982);
and UO_916 (O_916,N_4840,N_4920);
nor UO_917 (O_917,N_4997,N_4819);
nand UO_918 (O_918,N_4935,N_4846);
nand UO_919 (O_919,N_4939,N_4997);
nand UO_920 (O_920,N_4822,N_4867);
or UO_921 (O_921,N_4943,N_4864);
or UO_922 (O_922,N_4825,N_4854);
nand UO_923 (O_923,N_4978,N_4941);
nor UO_924 (O_924,N_4898,N_4880);
nand UO_925 (O_925,N_4832,N_4879);
xor UO_926 (O_926,N_4956,N_4970);
nand UO_927 (O_927,N_4834,N_4954);
and UO_928 (O_928,N_4959,N_4916);
and UO_929 (O_929,N_4929,N_4833);
nor UO_930 (O_930,N_4919,N_4965);
nor UO_931 (O_931,N_4805,N_4845);
nand UO_932 (O_932,N_4970,N_4932);
nand UO_933 (O_933,N_4878,N_4829);
nor UO_934 (O_934,N_4928,N_4860);
or UO_935 (O_935,N_4867,N_4944);
and UO_936 (O_936,N_4868,N_4985);
nand UO_937 (O_937,N_4897,N_4951);
nor UO_938 (O_938,N_4985,N_4945);
nand UO_939 (O_939,N_4880,N_4971);
or UO_940 (O_940,N_4903,N_4852);
nor UO_941 (O_941,N_4973,N_4845);
nand UO_942 (O_942,N_4965,N_4808);
nor UO_943 (O_943,N_4830,N_4823);
or UO_944 (O_944,N_4894,N_4899);
nor UO_945 (O_945,N_4956,N_4876);
or UO_946 (O_946,N_4828,N_4992);
and UO_947 (O_947,N_4827,N_4937);
and UO_948 (O_948,N_4801,N_4930);
nand UO_949 (O_949,N_4930,N_4902);
xnor UO_950 (O_950,N_4987,N_4804);
nand UO_951 (O_951,N_4832,N_4804);
or UO_952 (O_952,N_4947,N_4873);
or UO_953 (O_953,N_4918,N_4810);
nand UO_954 (O_954,N_4831,N_4890);
nor UO_955 (O_955,N_4955,N_4949);
nor UO_956 (O_956,N_4965,N_4922);
or UO_957 (O_957,N_4975,N_4924);
or UO_958 (O_958,N_4848,N_4901);
or UO_959 (O_959,N_4929,N_4847);
nand UO_960 (O_960,N_4939,N_4982);
nand UO_961 (O_961,N_4856,N_4979);
or UO_962 (O_962,N_4843,N_4879);
nor UO_963 (O_963,N_4927,N_4933);
or UO_964 (O_964,N_4828,N_4889);
and UO_965 (O_965,N_4964,N_4816);
nand UO_966 (O_966,N_4983,N_4986);
and UO_967 (O_967,N_4990,N_4868);
and UO_968 (O_968,N_4838,N_4925);
nand UO_969 (O_969,N_4851,N_4918);
nand UO_970 (O_970,N_4843,N_4978);
or UO_971 (O_971,N_4843,N_4817);
or UO_972 (O_972,N_4895,N_4825);
or UO_973 (O_973,N_4812,N_4841);
nor UO_974 (O_974,N_4823,N_4930);
nor UO_975 (O_975,N_4966,N_4858);
and UO_976 (O_976,N_4888,N_4812);
nand UO_977 (O_977,N_4966,N_4909);
nor UO_978 (O_978,N_4972,N_4869);
nand UO_979 (O_979,N_4974,N_4862);
nor UO_980 (O_980,N_4929,N_4956);
or UO_981 (O_981,N_4891,N_4919);
and UO_982 (O_982,N_4913,N_4995);
nor UO_983 (O_983,N_4930,N_4914);
nand UO_984 (O_984,N_4874,N_4999);
or UO_985 (O_985,N_4901,N_4888);
and UO_986 (O_986,N_4849,N_4925);
or UO_987 (O_987,N_4968,N_4867);
nand UO_988 (O_988,N_4999,N_4936);
nand UO_989 (O_989,N_4852,N_4893);
or UO_990 (O_990,N_4953,N_4810);
nand UO_991 (O_991,N_4948,N_4896);
nand UO_992 (O_992,N_4857,N_4962);
nor UO_993 (O_993,N_4837,N_4949);
nand UO_994 (O_994,N_4953,N_4816);
and UO_995 (O_995,N_4890,N_4901);
xor UO_996 (O_996,N_4855,N_4925);
nand UO_997 (O_997,N_4879,N_4861);
nand UO_998 (O_998,N_4919,N_4918);
xnor UO_999 (O_999,N_4882,N_4991);
endmodule