module basic_2500_25000_3000_100_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_131,In_599);
and U1 (N_1,In_1247,In_445);
or U2 (N_2,In_2323,In_1615);
xor U3 (N_3,In_184,In_1179);
xnor U4 (N_4,In_2361,In_1498);
nor U5 (N_5,In_2006,In_820);
and U6 (N_6,In_2457,In_1654);
and U7 (N_7,In_240,In_1770);
nor U8 (N_8,In_323,In_2077);
nand U9 (N_9,In_2037,In_41);
or U10 (N_10,In_1979,In_174);
or U11 (N_11,In_1273,In_2447);
xor U12 (N_12,In_1111,In_2452);
xor U13 (N_13,In_2218,In_1637);
or U14 (N_14,In_814,In_892);
or U15 (N_15,In_865,In_17);
and U16 (N_16,In_616,In_2263);
and U17 (N_17,In_2220,In_2003);
or U18 (N_18,In_1538,In_2126);
and U19 (N_19,In_1905,In_2360);
xnor U20 (N_20,In_791,In_2418);
nand U21 (N_21,In_662,In_2476);
nor U22 (N_22,In_263,In_1885);
nand U23 (N_23,In_2048,In_919);
xnor U24 (N_24,In_2245,In_154);
xor U25 (N_25,In_459,In_2058);
or U26 (N_26,In_1049,In_710);
nand U27 (N_27,In_54,In_1570);
and U28 (N_28,In_1258,In_187);
and U29 (N_29,In_49,In_1406);
nand U30 (N_30,In_2273,In_1157);
nand U31 (N_31,In_731,In_1205);
nand U32 (N_32,In_2009,In_2300);
nand U33 (N_33,In_626,In_787);
nor U34 (N_34,In_2364,In_816);
xnor U35 (N_35,In_1360,In_166);
or U36 (N_36,In_1963,In_2270);
xor U37 (N_37,In_1248,In_128);
nand U38 (N_38,In_124,In_754);
nand U39 (N_39,In_1984,In_117);
nor U40 (N_40,In_1310,In_1344);
or U41 (N_41,In_1565,In_717);
nor U42 (N_42,In_1268,In_2340);
and U43 (N_43,In_903,In_2297);
and U44 (N_44,In_56,In_1337);
or U45 (N_45,In_1354,In_2331);
nor U46 (N_46,In_123,In_1171);
xor U47 (N_47,In_2293,In_2413);
nor U48 (N_48,In_2326,In_2443);
or U49 (N_49,In_1071,In_1782);
xnor U50 (N_50,In_947,In_1780);
or U51 (N_51,In_2493,In_1038);
and U52 (N_52,In_673,In_525);
or U53 (N_53,In_2351,In_2159);
nor U54 (N_54,In_2176,In_278);
xnor U55 (N_55,In_427,In_2061);
or U56 (N_56,In_2164,In_2213);
nor U57 (N_57,In_2154,In_1808);
xor U58 (N_58,In_2316,In_946);
and U59 (N_59,In_970,In_850);
and U60 (N_60,In_1469,In_2483);
or U61 (N_61,In_1165,In_2199);
nand U62 (N_62,In_1145,In_640);
xor U63 (N_63,In_2389,In_1426);
nand U64 (N_64,In_1900,In_341);
xnor U65 (N_65,In_1773,In_2022);
or U66 (N_66,In_2466,In_1217);
xor U67 (N_67,In_678,In_1919);
or U68 (N_68,In_1184,In_189);
or U69 (N_69,In_1794,In_473);
nand U70 (N_70,In_193,In_1875);
and U71 (N_71,In_1699,In_2454);
nor U72 (N_72,In_1456,In_311);
xnor U73 (N_73,In_37,In_1209);
nor U74 (N_74,In_1660,In_160);
and U75 (N_75,In_923,In_1430);
xnor U76 (N_76,In_1580,In_556);
or U77 (N_77,In_543,In_752);
nor U78 (N_78,In_2070,In_1853);
xnor U79 (N_79,In_1126,In_243);
nor U80 (N_80,In_1192,In_1723);
xnor U81 (N_81,In_637,In_1581);
or U82 (N_82,In_294,In_1446);
or U83 (N_83,In_446,In_748);
nand U84 (N_84,In_1471,In_2183);
nor U85 (N_85,In_35,In_1944);
nor U86 (N_86,In_1010,In_1492);
nand U87 (N_87,In_1864,In_1137);
nor U88 (N_88,In_1345,In_1898);
and U89 (N_89,In_547,In_1130);
nand U90 (N_90,In_1241,In_338);
or U91 (N_91,In_310,In_1429);
nand U92 (N_92,In_1549,In_284);
nor U93 (N_93,In_2371,In_1801);
nor U94 (N_94,In_438,In_2414);
and U95 (N_95,In_2083,In_2259);
nand U96 (N_96,In_1792,In_262);
nand U97 (N_97,In_1428,In_1011);
nand U98 (N_98,In_139,In_1735);
nor U99 (N_99,In_343,In_272);
nor U100 (N_100,In_623,In_1304);
nand U101 (N_101,In_258,In_1215);
nor U102 (N_102,In_1749,In_855);
nand U103 (N_103,In_1854,In_1674);
nor U104 (N_104,In_1131,In_2444);
nand U105 (N_105,In_1954,In_712);
or U106 (N_106,In_1845,In_213);
nand U107 (N_107,In_967,In_1932);
or U108 (N_108,In_2288,In_1659);
nand U109 (N_109,In_1311,In_1933);
nor U110 (N_110,In_1265,In_212);
nand U111 (N_111,In_1557,In_1007);
or U112 (N_112,In_274,In_1783);
and U113 (N_113,In_1180,In_2087);
and U114 (N_114,In_1608,In_2084);
and U115 (N_115,In_186,In_1865);
or U116 (N_116,In_839,In_122);
or U117 (N_117,In_1104,In_1534);
xnor U118 (N_118,In_1462,In_380);
nor U119 (N_119,In_2461,In_1275);
xnor U120 (N_120,In_2252,In_289);
or U121 (N_121,In_998,In_760);
and U122 (N_122,In_2395,In_1561);
nor U123 (N_123,In_2404,In_2327);
or U124 (N_124,In_236,In_396);
xnor U125 (N_125,In_1347,In_144);
or U126 (N_126,In_422,In_2460);
and U127 (N_127,In_636,In_1294);
and U128 (N_128,In_251,In_1955);
xor U129 (N_129,In_237,In_1411);
nor U130 (N_130,In_141,In_2482);
nand U131 (N_131,In_235,In_142);
xor U132 (N_132,In_1587,In_2317);
or U133 (N_133,In_1826,In_1260);
nor U134 (N_134,In_29,In_1645);
nor U135 (N_135,In_127,In_1724);
nand U136 (N_136,In_1213,In_1834);
nand U137 (N_137,In_2028,In_1786);
nand U138 (N_138,In_1006,In_2489);
xor U139 (N_139,In_366,In_2302);
nand U140 (N_140,In_1523,In_324);
or U141 (N_141,In_1230,In_2335);
and U142 (N_142,In_518,In_978);
nand U143 (N_143,In_1370,In_625);
or U144 (N_144,In_1761,In_620);
and U145 (N_145,In_936,In_671);
nor U146 (N_146,In_2142,In_2093);
nor U147 (N_147,In_2255,In_1291);
or U148 (N_148,In_1282,In_904);
or U149 (N_149,In_1828,In_680);
nand U150 (N_150,In_440,In_780);
nor U151 (N_151,In_1218,In_1142);
nand U152 (N_152,In_1470,In_1402);
or U153 (N_153,In_1415,In_8);
nand U154 (N_154,In_1056,In_1926);
xor U155 (N_155,In_431,In_293);
nor U156 (N_156,In_639,In_1817);
and U157 (N_157,In_521,In_1095);
or U158 (N_158,In_701,In_1895);
or U159 (N_159,In_1434,In_1738);
nor U160 (N_160,In_1520,In_1222);
nor U161 (N_161,In_206,In_1316);
and U162 (N_162,In_38,In_2200);
nor U163 (N_163,In_511,In_1298);
or U164 (N_164,In_484,In_2248);
xnor U165 (N_165,In_485,In_1063);
and U166 (N_166,In_2422,In_171);
nor U167 (N_167,In_708,In_1403);
and U168 (N_168,In_617,In_67);
or U169 (N_169,In_58,In_574);
and U170 (N_170,In_2212,In_2014);
or U171 (N_171,In_1968,In_1270);
xnor U172 (N_172,In_1663,In_857);
nor U173 (N_173,In_1119,In_1053);
and U174 (N_174,In_98,In_1026);
and U175 (N_175,In_1886,In_1485);
or U176 (N_176,In_702,In_515);
and U177 (N_177,In_798,In_394);
xnor U178 (N_178,In_1941,In_503);
or U179 (N_179,In_2057,In_1);
nor U180 (N_180,In_88,In_492);
or U181 (N_181,In_704,In_1301);
xor U182 (N_182,In_1141,In_893);
xor U183 (N_183,In_1863,In_1443);
nand U184 (N_184,In_2221,In_1516);
nor U185 (N_185,In_2049,In_1057);
xor U186 (N_186,In_1987,In_1913);
nor U187 (N_187,In_1669,In_1767);
and U188 (N_188,In_42,In_887);
nor U189 (N_189,In_447,In_937);
and U190 (N_190,In_1021,In_1093);
or U191 (N_191,In_1398,In_1476);
nand U192 (N_192,In_2148,In_2353);
nand U193 (N_193,In_1855,In_1951);
nor U194 (N_194,In_1902,In_968);
and U195 (N_195,In_333,In_1986);
or U196 (N_196,In_2090,In_2105);
nand U197 (N_197,In_1159,In_2125);
nor U198 (N_198,In_1607,In_1810);
nor U199 (N_199,In_2226,In_2133);
xnor U200 (N_200,In_2031,In_1843);
xor U201 (N_201,In_1251,In_573);
xor U202 (N_202,In_1976,In_513);
nand U203 (N_203,In_416,In_992);
xor U204 (N_204,In_1064,In_2102);
or U205 (N_205,In_2394,In_1766);
xor U206 (N_206,In_175,In_581);
or U207 (N_207,In_552,In_303);
or U208 (N_208,In_1259,In_1558);
nand U209 (N_209,In_2195,In_2425);
nor U210 (N_210,In_533,In_849);
nand U211 (N_211,In_1803,In_241);
nor U212 (N_212,In_1500,In_351);
or U213 (N_213,In_2411,In_2118);
xnor U214 (N_214,In_1728,In_995);
or U215 (N_215,In_1466,In_1715);
xnor U216 (N_216,In_593,In_1975);
nor U217 (N_217,In_1383,In_390);
nand U218 (N_218,In_2309,In_907);
nor U219 (N_219,In_2408,In_1676);
nand U220 (N_220,In_1228,In_1689);
or U221 (N_221,In_1395,In_1278);
or U222 (N_222,In_1593,In_2069);
xnor U223 (N_223,In_1582,In_1318);
nand U224 (N_224,In_2374,In_860);
xnor U225 (N_225,In_2065,In_2169);
nand U226 (N_226,In_945,In_786);
nand U227 (N_227,In_1404,In_1363);
nand U228 (N_228,In_1477,In_455);
and U229 (N_229,In_340,In_544);
and U230 (N_230,In_826,In_761);
or U231 (N_231,In_1336,In_570);
nand U232 (N_232,In_1326,In_1991);
and U233 (N_233,In_2187,In_107);
nor U234 (N_234,In_1096,In_328);
nand U235 (N_235,In_2315,In_1977);
and U236 (N_236,In_1529,In_2388);
nand U237 (N_237,In_990,In_707);
nor U238 (N_238,In_2188,In_932);
xnor U239 (N_239,In_1331,In_225);
nor U240 (N_240,In_2209,In_987);
or U241 (N_241,In_999,In_1559);
or U242 (N_242,In_1505,In_253);
or U243 (N_243,In_1914,In_822);
nand U244 (N_244,In_153,In_762);
xor U245 (N_245,In_800,In_2429);
nand U246 (N_246,In_1619,In_1702);
and U247 (N_247,In_2344,In_2310);
xor U248 (N_248,In_993,In_2092);
xor U249 (N_249,In_629,In_2358);
xnor U250 (N_250,In_631,In_2107);
nand U251 (N_251,In_137,In_306);
nor U252 (N_252,In_775,In_506);
xnor U253 (N_253,In_1579,In_1254);
or U254 (N_254,In_1765,In_1138);
and U255 (N_255,In_989,In_1566);
nand U256 (N_256,In_2324,In_668);
nor U257 (N_257,In_1051,N_100);
or U258 (N_258,In_75,In_1210);
nand U259 (N_259,In_345,N_217);
xnor U260 (N_260,In_1473,In_2046);
nand U261 (N_261,N_188,In_1405);
nand U262 (N_262,In_1849,In_1460);
and U263 (N_263,In_742,In_654);
and U264 (N_264,In_2285,N_94);
nand U265 (N_265,In_650,In_528);
or U266 (N_266,In_612,In_1638);
nand U267 (N_267,In_2428,In_1758);
xnor U268 (N_268,In_143,In_1322);
xor U269 (N_269,In_1151,In_1467);
and U270 (N_270,In_2250,In_1644);
nand U271 (N_271,In_304,In_2455);
or U272 (N_272,In_1504,In_1734);
xor U273 (N_273,In_818,In_1465);
or U274 (N_274,In_1160,In_804);
nand U275 (N_275,N_208,N_237);
nand U276 (N_276,In_2217,In_1245);
xor U277 (N_277,In_981,In_2000);
xor U278 (N_278,In_5,In_1974);
or U279 (N_279,In_530,In_1704);
and U280 (N_280,In_494,In_1379);
xnor U281 (N_281,In_2086,In_1733);
xnor U282 (N_282,In_1501,In_1166);
or U283 (N_283,In_1385,N_216);
nand U284 (N_284,In_935,In_2264);
and U285 (N_285,In_2433,In_2230);
xor U286 (N_286,In_2030,In_1631);
and U287 (N_287,In_412,In_2227);
nand U288 (N_288,In_920,In_2321);
or U289 (N_289,In_778,In_1277);
nor U290 (N_290,In_1391,In_1475);
or U291 (N_291,In_413,In_1329);
xor U292 (N_292,In_1703,In_2190);
nor U293 (N_293,In_1949,N_242);
nand U294 (N_294,In_1811,In_1121);
and U295 (N_295,In_1636,In_2400);
nor U296 (N_296,In_550,In_635);
nand U297 (N_297,In_2244,In_886);
xor U298 (N_298,In_1693,In_2269);
nand U299 (N_299,N_179,In_1651);
or U300 (N_300,In_2062,N_66);
or U301 (N_301,In_2258,In_1113);
nand U302 (N_302,In_2256,In_1726);
xor U303 (N_303,In_238,In_1697);
and U304 (N_304,In_176,In_1981);
nor U305 (N_305,In_1164,In_890);
xnor U306 (N_306,In_1400,In_1450);
and U307 (N_307,In_103,In_147);
nor U308 (N_308,In_1355,In_2041);
xor U309 (N_309,In_2091,In_1356);
or U310 (N_310,In_1483,In_1237);
and U311 (N_311,In_1934,In_2468);
nand U312 (N_312,N_138,In_519);
nor U313 (N_313,In_386,In_2392);
nand U314 (N_314,In_1199,In_2238);
and U315 (N_315,In_1317,In_2306);
nand U316 (N_316,In_827,In_1369);
or U317 (N_317,In_1343,In_472);
and U318 (N_318,In_256,In_2410);
nor U319 (N_319,In_2026,In_876);
xor U320 (N_320,In_1267,In_1745);
xor U321 (N_321,In_493,In_885);
and U322 (N_322,In_1805,In_705);
xnor U323 (N_323,In_2241,In_470);
or U324 (N_324,In_1929,In_882);
and U325 (N_325,In_2224,In_1838);
or U326 (N_326,In_2137,In_1844);
and U327 (N_327,N_235,In_715);
xnor U328 (N_328,In_833,In_1796);
xor U329 (N_329,In_1410,In_2004);
xnor U330 (N_330,In_1208,In_2391);
nand U331 (N_331,In_1711,In_220);
nand U332 (N_332,In_1156,In_2231);
or U333 (N_333,In_168,In_1731);
nand U334 (N_334,In_1576,In_618);
xnor U335 (N_335,In_410,In_105);
or U336 (N_336,In_401,In_1445);
xnor U337 (N_337,In_2072,In_2446);
nand U338 (N_338,N_122,In_1563);
or U339 (N_339,In_239,In_1246);
or U340 (N_340,In_1435,In_1081);
or U341 (N_341,In_834,In_387);
or U342 (N_342,In_93,N_219);
nand U343 (N_343,In_1721,In_1964);
xnor U344 (N_344,In_1662,In_486);
xor U345 (N_345,In_1220,In_167);
or U346 (N_346,N_32,In_1824);
and U347 (N_347,In_1709,In_2112);
nand U348 (N_348,In_592,In_178);
or U349 (N_349,N_245,In_2172);
or U350 (N_350,N_205,In_465);
and U351 (N_351,In_703,In_1312);
and U352 (N_352,N_226,In_698);
nor U353 (N_353,N_55,In_2120);
xnor U354 (N_354,In_2016,In_1630);
nor U355 (N_355,N_62,In_955);
xnor U356 (N_356,In_79,In_1596);
or U357 (N_357,In_2354,In_1008);
nor U358 (N_358,In_463,In_2098);
and U359 (N_359,In_594,In_145);
nor U360 (N_360,In_1859,In_769);
nor U361 (N_361,N_224,In_1269);
nand U362 (N_362,In_2456,In_2445);
or U363 (N_363,N_29,In_1441);
and U364 (N_364,In_824,In_2267);
and U365 (N_365,In_1306,In_576);
xor U366 (N_366,In_790,In_548);
or U367 (N_367,In_542,In_260);
and U368 (N_368,In_1906,In_27);
xnor U369 (N_369,In_1725,In_1299);
and U370 (N_370,In_182,In_1302);
xor U371 (N_371,In_223,In_1629);
and U372 (N_372,In_2407,In_645);
or U373 (N_373,N_181,In_1670);
and U374 (N_374,In_23,In_524);
or U375 (N_375,In_723,In_746);
nand U376 (N_376,In_1396,In_2451);
and U377 (N_377,In_1169,In_807);
or U378 (N_378,In_481,In_1996);
xnor U379 (N_379,In_873,In_916);
nand U380 (N_380,N_136,In_10);
and U381 (N_381,In_1793,In_1648);
nor U382 (N_382,In_951,In_693);
nor U383 (N_383,In_2420,In_1188);
or U384 (N_384,In_403,In_765);
and U385 (N_385,In_2140,In_1283);
or U386 (N_386,In_901,N_192);
and U387 (N_387,In_36,N_75);
nand U388 (N_388,In_1155,N_137);
and U389 (N_389,In_1797,In_1789);
and U390 (N_390,In_2033,In_1285);
or U391 (N_391,N_81,In_1862);
or U392 (N_392,N_215,In_852);
or U393 (N_393,In_2472,In_1778);
or U394 (N_394,In_1571,N_31);
or U395 (N_395,In_1102,N_153);
or U396 (N_396,In_1392,In_218);
nor U397 (N_397,In_2431,In_442);
nor U398 (N_398,In_1531,In_1556);
and U399 (N_399,In_1055,In_719);
and U400 (N_400,In_1948,N_218);
and U401 (N_401,In_376,N_180);
nand U402 (N_402,In_1146,In_2415);
xnor U403 (N_403,N_107,In_2257);
or U404 (N_404,N_220,In_732);
and U405 (N_405,In_562,In_2134);
xnor U406 (N_406,N_162,In_32);
and U407 (N_407,In_1583,In_577);
nand U408 (N_408,N_108,In_25);
nand U409 (N_409,In_1816,In_2254);
or U410 (N_410,In_20,N_11);
or U411 (N_411,In_1009,In_1280);
and U412 (N_412,In_2100,In_538);
nor U413 (N_413,In_2122,In_259);
and U414 (N_414,In_50,N_123);
nor U415 (N_415,N_155,In_974);
xor U416 (N_416,In_914,In_764);
or U417 (N_417,In_1564,N_130);
nor U418 (N_418,In_1378,In_1321);
nor U419 (N_419,In_1958,In_1459);
xor U420 (N_420,In_1050,In_1062);
or U421 (N_421,In_1233,In_1152);
nand U422 (N_422,In_169,In_332);
nor U423 (N_423,In_733,In_450);
or U424 (N_424,In_1992,In_467);
nor U425 (N_425,In_686,In_221);
nand U426 (N_426,In_1324,In_1120);
and U427 (N_427,In_423,In_1706);
or U428 (N_428,In_871,N_232);
xor U429 (N_429,In_2329,In_2047);
or U430 (N_430,In_1373,In_1536);
and U431 (N_431,N_70,In_1621);
xnor U432 (N_432,In_2002,In_582);
nand U433 (N_433,In_2253,In_1072);
and U434 (N_434,In_110,In_1397);
and U435 (N_435,In_209,In_1628);
xor U436 (N_436,N_204,In_452);
nand U437 (N_437,In_2146,In_0);
nor U438 (N_438,In_1533,In_555);
nor U439 (N_439,In_1181,In_1463);
and U440 (N_440,In_2399,In_1236);
and U441 (N_441,In_104,N_102);
and U442 (N_442,N_167,In_1161);
nor U443 (N_443,In_2390,In_2325);
or U444 (N_444,In_1425,In_121);
nand U445 (N_445,In_299,In_198);
or U446 (N_446,In_801,In_1802);
and U447 (N_447,In_350,In_1227);
nor U448 (N_448,In_1114,In_1399);
or U449 (N_449,In_2382,In_2368);
and U450 (N_450,In_1436,In_540);
nor U451 (N_451,N_190,In_1655);
or U452 (N_452,In_1994,In_808);
xnor U453 (N_453,In_2330,N_12);
nor U454 (N_454,In_290,In_1718);
and U455 (N_455,In_1387,In_1315);
and U456 (N_456,In_233,In_1742);
xor U457 (N_457,In_2423,In_2369);
xor U458 (N_458,In_656,In_2470);
xnor U459 (N_459,In_1195,In_1671);
nand U460 (N_460,In_96,In_211);
and U461 (N_461,In_1874,In_357);
and U462 (N_462,In_614,In_1950);
and U463 (N_463,In_449,In_848);
xnor U464 (N_464,In_402,In_2158);
or U465 (N_465,In_1978,In_1769);
nand U466 (N_466,N_223,N_248);
xor U467 (N_467,In_2492,In_565);
nor U468 (N_468,In_47,In_553);
nand U469 (N_469,In_1692,In_1668);
nor U470 (N_470,In_2484,In_215);
or U471 (N_471,In_1752,N_79);
xnor U472 (N_472,In_983,In_1681);
nor U473 (N_473,N_202,In_2471);
or U474 (N_474,In_330,In_1686);
and U475 (N_475,In_690,In_1930);
or U476 (N_476,In_1879,In_2294);
nor U477 (N_477,In_858,In_609);
nand U478 (N_478,In_111,In_320);
xnor U479 (N_479,In_1719,In_1257);
xor U480 (N_480,In_2333,In_2442);
and U481 (N_481,In_292,In_1086);
and U482 (N_482,In_1376,In_2063);
and U483 (N_483,In_1335,N_97);
xnor U484 (N_484,In_1226,In_984);
nor U485 (N_485,In_1781,In_1545);
nor U486 (N_486,In_1133,In_1649);
and U487 (N_487,In_1232,In_52);
nand U488 (N_488,In_1212,In_78);
or U489 (N_489,In_1904,In_2064);
nor U490 (N_490,In_2071,In_1044);
or U491 (N_491,In_2332,In_1235);
nor U492 (N_492,In_1082,In_480);
or U493 (N_493,In_2201,In_2210);
xor U494 (N_494,In_2149,In_1183);
and U495 (N_495,In_2345,In_600);
or U496 (N_496,In_2163,In_1988);
or U497 (N_497,In_2338,In_1490);
or U498 (N_498,In_1320,In_1388);
nand U499 (N_499,In_150,In_348);
nand U500 (N_500,N_486,In_1650);
nand U501 (N_501,In_862,In_931);
or U502 (N_502,In_45,In_81);
xor U503 (N_503,In_1309,In_1330);
nand U504 (N_504,In_1153,In_1727);
and U505 (N_505,In_2491,In_432);
xnor U506 (N_506,N_424,N_358);
nor U507 (N_507,In_1461,In_2008);
xor U508 (N_508,In_792,In_1846);
and U509 (N_509,N_93,In_739);
or U510 (N_510,In_1069,N_326);
or U511 (N_511,In_1271,In_926);
xor U512 (N_512,N_306,In_2029);
xor U513 (N_513,In_2450,In_371);
xnor U514 (N_514,In_1013,In_326);
or U515 (N_515,N_57,In_2295);
and U516 (N_516,In_1274,N_90);
nor U517 (N_517,In_1829,In_691);
and U518 (N_518,In_1468,In_2211);
nor U519 (N_519,In_880,In_1019);
nor U520 (N_520,In_924,In_1548);
and U521 (N_521,In_331,N_293);
nor U522 (N_522,In_2075,In_720);
nand U523 (N_523,In_1041,In_2039);
nor U524 (N_524,In_242,In_19);
or U525 (N_525,In_2116,In_2150);
nor U526 (N_526,In_419,In_1117);
nand U527 (N_527,In_859,N_83);
nand U528 (N_528,In_1876,In_1384);
nor U529 (N_529,In_1207,In_2469);
and U530 (N_530,In_1641,In_1850);
and U531 (N_531,In_2373,In_1807);
and U532 (N_532,N_89,In_1386);
or U533 (N_533,In_33,N_114);
nand U534 (N_534,In_1746,In_1047);
and U535 (N_535,In_688,N_115);
and U536 (N_536,In_782,In_317);
nor U537 (N_537,N_272,In_1952);
or U538 (N_538,N_36,In_641);
and U539 (N_539,N_408,In_1956);
xnor U540 (N_540,N_48,In_309);
nor U541 (N_541,In_382,In_539);
xnor U542 (N_542,In_1763,In_2082);
xor U543 (N_543,In_1589,In_2370);
nor U544 (N_544,In_395,In_568);
xnor U545 (N_545,In_232,In_785);
and U546 (N_546,N_172,In_159);
or U547 (N_547,In_1967,In_551);
xor U548 (N_548,In_2222,In_1349);
xnor U549 (N_549,N_262,N_34);
nand U550 (N_550,In_583,In_1931);
nand U551 (N_551,In_510,In_1586);
and U552 (N_552,N_243,In_483);
or U553 (N_553,In_2307,In_1424);
xor U554 (N_554,In_1626,In_763);
and U555 (N_555,In_1661,In_2464);
xor U556 (N_556,In_72,In_230);
nor U557 (N_557,In_1600,In_2053);
or U558 (N_558,In_1541,In_12);
and U559 (N_559,In_185,N_234);
nor U560 (N_560,In_725,In_580);
and U561 (N_561,In_900,In_1393);
xnor U562 (N_562,In_361,In_1432);
nor U563 (N_563,N_105,N_295);
xor U564 (N_564,In_1224,In_2203);
or U565 (N_565,In_943,In_2152);
nor U566 (N_566,N_318,In_1412);
nor U567 (N_567,In_458,In_1078);
and U568 (N_568,In_421,N_431);
nor U569 (N_569,In_889,In_116);
xnor U570 (N_570,In_2108,N_440);
or U571 (N_571,In_2465,In_1239);
and U572 (N_572,In_921,In_273);
nor U573 (N_573,In_985,In_1613);
or U574 (N_574,N_384,N_189);
nor U575 (N_575,N_296,In_268);
xor U576 (N_576,In_196,N_46);
nand U577 (N_577,In_1890,In_1634);
xor U578 (N_578,In_779,In_1149);
and U579 (N_579,In_2156,In_2161);
or U580 (N_580,In_2129,N_314);
xnor U581 (N_581,In_318,N_365);
and U582 (N_582,In_870,In_1073);
nor U583 (N_583,N_64,In_1922);
nand U584 (N_584,In_1418,In_2430);
nand U585 (N_585,In_280,In_94);
nand U586 (N_586,In_1687,In_496);
nor U587 (N_587,In_1325,In_692);
and U588 (N_588,N_464,In_255);
and U589 (N_589,In_918,In_2229);
nor U590 (N_590,N_156,In_31);
xnor U591 (N_591,In_2490,In_1666);
or U592 (N_592,In_2113,In_468);
or U593 (N_593,In_1908,In_1037);
nor U594 (N_594,In_1106,In_89);
and U595 (N_595,In_1677,In_1889);
and U596 (N_596,N_28,N_310);
nor U597 (N_597,In_1771,In_2167);
xnor U598 (N_598,In_638,In_1109);
nor U599 (N_599,In_214,In_1525);
or U600 (N_600,In_172,In_2346);
or U601 (N_601,In_234,In_1389);
and U602 (N_602,N_392,In_1775);
nor U603 (N_603,In_1526,In_1888);
xnor U604 (N_604,In_1023,In_1296);
or U605 (N_605,In_2143,In_884);
and U606 (N_606,In_1417,In_986);
nand U607 (N_607,In_768,In_597);
nand U608 (N_608,In_794,N_485);
or U609 (N_609,In_2103,In_2165);
nor U610 (N_610,In_1288,In_647);
nand U611 (N_611,In_805,In_1835);
or U612 (N_612,In_1036,N_164);
nor U613 (N_613,N_203,In_819);
nand U614 (N_614,In_2085,N_428);
and U615 (N_615,In_60,In_2130);
xor U616 (N_616,In_1907,In_1174);
xor U617 (N_617,In_770,In_1016);
nor U618 (N_618,In_602,In_2271);
nor U619 (N_619,In_1680,In_1831);
and U620 (N_620,In_1891,In_210);
and U621 (N_621,In_1502,N_273);
xnor U622 (N_622,In_1925,In_397);
and U623 (N_623,N_16,In_1487);
xnor U624 (N_624,In_1266,N_341);
nor U625 (N_625,In_1422,In_1867);
and U626 (N_626,In_917,In_114);
nand U627 (N_627,In_1936,In_389);
nor U628 (N_628,In_1966,In_1458);
xnor U629 (N_629,In_420,In_475);
or U630 (N_630,In_1927,N_268);
and U631 (N_631,In_2379,In_1452);
and U632 (N_632,N_227,In_398);
nand U633 (N_633,In_1453,In_2228);
or U634 (N_634,In_1442,In_1140);
and U635 (N_635,In_689,In_1756);
xnor U636 (N_636,In_2318,In_1042);
nor U637 (N_637,In_1000,In_257);
nor U638 (N_638,In_961,In_2193);
nand U639 (N_639,In_2479,In_1127);
xnor U640 (N_640,In_1032,N_54);
and U641 (N_641,In_2043,N_421);
nand U642 (N_642,In_85,In_2025);
or U643 (N_643,In_2434,In_608);
nand U644 (N_644,In_632,N_148);
nor U645 (N_645,In_1736,In_959);
nand U646 (N_646,In_322,N_336);
xor U647 (N_647,In_1918,In_501);
nand U648 (N_648,In_2498,In_1408);
nand U649 (N_649,N_276,In_1851);
nand U650 (N_650,N_413,In_228);
nand U651 (N_651,In_349,N_150);
nor U652 (N_652,In_2066,N_140);
or U653 (N_653,In_996,In_1488);
or U654 (N_654,In_1646,In_1800);
xnor U655 (N_655,In_972,In_812);
xnor U656 (N_656,N_359,In_759);
xnor U657 (N_657,In_2198,In_2322);
or U658 (N_658,In_249,In_1601);
nor U659 (N_659,In_534,In_453);
nand U660 (N_660,In_505,In_1937);
or U661 (N_661,In_512,N_68);
and U662 (N_662,N_454,In_1658);
and U663 (N_663,N_72,In_744);
nor U664 (N_664,In_1688,N_321);
xnor U665 (N_665,In_912,N_283);
or U666 (N_666,N_438,In_405);
or U667 (N_667,In_2119,In_136);
nor U668 (N_668,In_92,N_19);
and U669 (N_669,In_897,N_374);
nor U670 (N_670,N_33,In_1705);
xnor U671 (N_671,In_277,In_352);
xnor U672 (N_672,In_430,In_1544);
or U673 (N_673,In_1560,N_448);
xnor U674 (N_674,In_1740,In_2151);
nor U675 (N_675,N_400,In_300);
or U676 (N_676,In_1058,In_1314);
and U677 (N_677,In_97,In_1061);
and U678 (N_678,N_354,In_90);
and U679 (N_679,N_261,In_1760);
xor U680 (N_680,N_65,In_606);
nand U681 (N_681,In_1656,In_526);
and U682 (N_682,N_24,In_16);
or U683 (N_683,In_265,In_302);
nand U684 (N_684,In_109,N_13);
xor U685 (N_685,In_2180,In_1381);
or U686 (N_686,In_180,In_694);
and U687 (N_687,In_1935,In_745);
xor U688 (N_688,In_2184,In_520);
nor U689 (N_689,In_1748,N_2);
nor U690 (N_690,In_404,In_1015);
nand U691 (N_691,N_125,N_161);
nor U692 (N_692,N_129,N_27);
nand U693 (N_693,In_1107,In_1897);
and U694 (N_694,In_584,In_155);
or U695 (N_695,In_2398,In_913);
xnor U696 (N_696,In_1540,In_1448);
nand U697 (N_697,In_1539,In_2242);
nand U698 (N_698,N_78,In_2234);
and U699 (N_699,In_1852,In_2136);
or U700 (N_700,In_2298,N_106);
nand U701 (N_701,In_385,In_478);
or U702 (N_702,In_202,In_364);
or U703 (N_703,In_558,N_92);
xnor U704 (N_704,N_38,In_2376);
nor U705 (N_705,In_535,In_2020);
or U706 (N_706,In_2453,N_35);
and U707 (N_707,N_355,In_1962);
and U708 (N_708,N_56,N_456);
nor U709 (N_709,In_1413,N_493);
and U710 (N_710,In_1364,In_298);
nor U711 (N_711,N_451,In_73);
xnor U712 (N_712,In_2074,In_488);
and U713 (N_713,In_767,N_370);
and U714 (N_714,In_164,In_1917);
xnor U715 (N_715,N_256,In_2280);
and U716 (N_716,In_1840,In_590);
or U717 (N_717,In_1550,In_2067);
and U718 (N_718,N_91,In_1856);
nor U719 (N_719,In_2287,In_1489);
and U720 (N_720,In_30,N_414);
or U721 (N_721,In_1033,In_1791);
and U722 (N_722,N_435,In_1454);
nor U723 (N_723,In_682,In_1372);
or U724 (N_724,In_541,N_174);
or U725 (N_725,N_308,In_2);
nand U726 (N_726,In_365,In_734);
nor U727 (N_727,N_327,N_152);
xnor U728 (N_728,In_227,In_979);
or U729 (N_729,N_353,In_1039);
nand U730 (N_730,N_285,In_2115);
nor U731 (N_731,In_1264,In_1018);
xnor U732 (N_732,In_222,In_1262);
and U733 (N_733,N_317,N_479);
and U734 (N_734,In_928,In_2435);
nand U735 (N_735,In_711,In_1499);
or U736 (N_736,In_205,In_958);
or U737 (N_737,In_1795,N_103);
nand U738 (N_738,In_1640,In_1880);
nor U739 (N_739,N_7,N_313);
or U740 (N_740,N_42,In_471);
nand U741 (N_741,In_2153,In_1598);
nor U742 (N_742,In_1043,N_426);
xor U743 (N_743,In_291,N_364);
xor U744 (N_744,N_98,In_1122);
nand U745 (N_745,In_836,In_1998);
xor U746 (N_746,N_447,In_2265);
or U747 (N_747,In_596,In_630);
nor U748 (N_748,In_709,In_2088);
nor U749 (N_749,In_1197,N_96);
nor U750 (N_750,In_700,N_573);
and U751 (N_751,In_1060,N_241);
nor U752 (N_752,In_40,N_533);
nor U753 (N_753,N_281,In_14);
and U754 (N_754,N_270,N_737);
nor U755 (N_755,N_391,N_213);
and U756 (N_756,In_1186,In_2186);
or U757 (N_757,In_2268,In_1377);
nor U758 (N_758,In_1067,In_1762);
or U759 (N_759,In_2282,In_813);
xnor U760 (N_760,N_658,In_627);
or U761 (N_761,N_342,In_1070);
xor U762 (N_762,In_2432,In_669);
or U763 (N_763,N_386,N_104);
nand U764 (N_764,In_2060,N_187);
nor U765 (N_765,N_372,In_68);
xor U766 (N_766,In_1739,In_2372);
and U767 (N_767,In_2243,N_290);
nor U768 (N_768,In_1240,N_228);
or U769 (N_769,In_1170,N_373);
xor U770 (N_770,In_1915,N_510);
nand U771 (N_771,N_524,In_1877);
and U772 (N_772,In_1367,In_1616);
or U773 (N_773,In_129,N_649);
and U774 (N_774,In_585,In_368);
and U775 (N_775,In_1286,N_47);
nor U776 (N_776,In_2286,N_334);
and U777 (N_777,In_1361,In_1255);
nand U778 (N_778,In_624,In_2144);
xor U779 (N_779,In_1785,N_168);
or U780 (N_780,In_716,In_2235);
xor U781 (N_781,In_406,In_1177);
xnor U782 (N_782,In_2251,N_282);
and U783 (N_783,In_1971,In_956);
and U784 (N_784,N_498,N_51);
nor U785 (N_785,In_676,In_1014);
nand U786 (N_786,In_648,N_585);
nand U787 (N_787,N_646,N_288);
nor U788 (N_788,N_49,In_199);
nor U789 (N_789,In_971,In_1481);
xor U790 (N_790,N_247,N_291);
nand U791 (N_791,In_1374,In_1591);
nand U792 (N_792,In_685,N_73);
nand U793 (N_793,In_2266,In_4);
or U794 (N_794,N_597,In_83);
nand U795 (N_795,In_1820,In_2089);
xor U796 (N_796,In_657,N_722);
nand U797 (N_797,In_1696,N_144);
nor U798 (N_798,In_106,In_777);
nor U799 (N_799,In_1457,In_15);
nand U800 (N_800,In_898,In_254);
or U801 (N_801,In_435,In_667);
and U802 (N_802,N_340,In_699);
and U803 (N_803,In_1744,N_742);
or U804 (N_804,N_0,In_1287);
nand U805 (N_805,N_407,In_119);
and U806 (N_806,In_2059,In_532);
or U807 (N_807,In_1508,In_477);
nand U808 (N_808,In_1401,In_1219);
nor U809 (N_809,N_668,In_674);
xnor U810 (N_810,N_363,N_176);
nand U811 (N_811,In_1804,In_2094);
nand U812 (N_812,In_566,In_2378);
nand U813 (N_813,In_1125,In_1577);
xor U814 (N_814,In_2359,In_1819);
nor U815 (N_815,In_1144,In_1923);
nand U816 (N_816,N_543,N_4);
or U817 (N_817,N_650,In_2367);
xnor U818 (N_818,In_864,N_133);
nand U819 (N_819,N_548,N_519);
xnor U820 (N_820,N_483,N_319);
and U821 (N_821,N_606,N_542);
nand U822 (N_822,N_662,In_2343);
xnor U823 (N_823,N_655,In_1517);
nor U824 (N_824,In_2032,In_1784);
xor U825 (N_825,In_1390,N_732);
nor U826 (N_826,In_1162,In_1204);
and U827 (N_827,N_729,N_324);
or U828 (N_828,N_579,In_34);
xor U829 (N_829,N_134,In_1633);
and U830 (N_830,In_1341,In_830);
nand U831 (N_831,N_690,N_111);
nor U832 (N_832,In_1868,In_508);
or U833 (N_833,N_323,In_201);
xnor U834 (N_834,In_347,N_528);
xnor U835 (N_835,In_2249,In_1185);
nand U836 (N_836,In_910,In_1029);
xor U837 (N_837,N_577,In_113);
nand U838 (N_838,N_501,N_626);
or U839 (N_839,N_378,N_664);
nand U840 (N_840,N_613,In_842);
xor U841 (N_841,N_605,In_753);
or U842 (N_842,In_724,N_499);
or U843 (N_843,N_651,In_2175);
or U844 (N_844,N_286,In_1005);
nor U845 (N_845,N_320,N_629);
nand U846 (N_846,In_1882,In_1150);
nor U847 (N_847,N_446,N_8);
nor U848 (N_848,In_851,In_57);
xnor U849 (N_849,In_1289,In_2419);
xor U850 (N_850,In_2274,In_51);
or U851 (N_851,In_1892,In_425);
and U852 (N_852,In_1861,In_817);
nand U853 (N_853,In_1173,N_165);
nand U854 (N_854,N_297,N_581);
or U855 (N_855,N_44,N_462);
nand U856 (N_856,In_658,N_538);
and U857 (N_857,N_21,In_1158);
nand U858 (N_858,N_22,N_246);
nor U859 (N_859,In_2401,In_183);
or U860 (N_860,N_686,In_118);
nor U861 (N_861,In_2178,In_1916);
nand U862 (N_862,In_1753,N_653);
nor U863 (N_863,In_1546,In_684);
xnor U864 (N_864,In_905,In_285);
xnor U865 (N_865,N_625,In_1167);
xnor U866 (N_866,In_2124,In_1211);
xnor U867 (N_867,N_275,In_1690);
and U868 (N_868,In_1261,In_3);
or U869 (N_869,In_1827,In_982);
nor U870 (N_870,N_708,In_706);
and U871 (N_871,In_829,In_1099);
xor U872 (N_872,In_578,In_489);
and U873 (N_873,In_1836,In_1447);
nor U874 (N_874,N_410,In_743);
and U875 (N_875,In_908,N_482);
nor U876 (N_876,In_2170,N_560);
nand U877 (N_877,In_1695,N_411);
nor U878 (N_878,In_429,In_9);
xnor U879 (N_879,In_1813,In_2342);
xnor U880 (N_880,In_495,In_784);
or U881 (N_881,In_595,In_1416);
nor U882 (N_882,In_1419,In_1045);
or U883 (N_883,In_1365,In_911);
nand U884 (N_884,N_595,In_76);
nand U885 (N_885,N_600,In_735);
and U886 (N_886,N_312,In_152);
nor U887 (N_887,In_1957,N_344);
nor U888 (N_888,In_756,In_665);
or U889 (N_889,In_2311,In_1894);
nand U890 (N_890,In_163,In_1143);
or U891 (N_891,In_1682,In_2132);
nor U892 (N_892,N_266,In_844);
and U893 (N_893,N_26,In_126);
nor U894 (N_894,In_1527,In_462);
and U895 (N_895,In_2279,N_436);
xnor U896 (N_896,In_1148,In_537);
or U897 (N_897,N_667,In_400);
or U898 (N_898,N_615,In_335);
or U899 (N_899,In_53,In_2352);
and U900 (N_900,In_1420,N_199);
nand U901 (N_901,N_294,In_1945);
nand U902 (N_902,In_266,N_720);
nand U903 (N_903,In_1472,In_80);
xnor U904 (N_904,In_1079,In_1368);
nor U905 (N_905,In_563,In_687);
and U906 (N_906,In_934,In_696);
nand U907 (N_907,N_660,In_1409);
nand U908 (N_908,N_20,N_559);
nand U909 (N_909,In_1124,In_448);
nand U910 (N_910,N_504,In_730);
and U911 (N_911,N_361,In_1059);
xor U912 (N_912,In_454,In_1920);
xor U913 (N_913,In_1136,In_250);
nand U914 (N_914,N_683,In_342);
nor U915 (N_915,In_130,In_1672);
xor U916 (N_916,In_2042,N_561);
xnor U917 (N_917,N_500,N_126);
and U918 (N_918,In_869,In_1909);
xor U919 (N_919,In_2437,In_2494);
nor U920 (N_920,N_691,N_390);
nand U921 (N_921,In_1242,In_1348);
nand U922 (N_922,N_682,In_1098);
nand U923 (N_923,In_1089,In_443);
or U924 (N_924,In_938,N_592);
and U925 (N_925,In_270,In_1764);
xor U926 (N_926,In_2350,In_1684);
xnor U927 (N_927,In_2424,N_131);
xor U928 (N_928,In_2405,In_2051);
xor U929 (N_929,In_1444,In_2179);
xnor U930 (N_930,N_419,N_149);
nand U931 (N_931,In_517,In_878);
and U932 (N_932,N_117,In_2397);
xor U933 (N_933,N_250,In_933);
nor U934 (N_934,In_843,In_61);
nand U935 (N_935,In_1606,In_1940);
nor U936 (N_936,N_659,In_1642);
nand U937 (N_937,N_145,N_120);
nand U938 (N_938,N_636,In_2012);
or U939 (N_939,N_170,In_1653);
nor U940 (N_940,N_596,In_408);
and U941 (N_941,In_988,N_680);
and U942 (N_942,In_514,N_240);
and U943 (N_943,In_1074,N_439);
nor U944 (N_944,N_271,N_707);
or U945 (N_945,In_1478,N_470);
nor U946 (N_946,N_638,In_2487);
and U947 (N_947,N_478,N_401);
or U948 (N_948,N_745,In_589);
and U949 (N_949,In_622,N_331);
xnor U950 (N_950,In_1713,In_2219);
nor U951 (N_951,In_1479,In_296);
nor U952 (N_952,In_388,In_1537);
nor U953 (N_953,In_194,In_729);
nand U954 (N_954,In_1722,In_2341);
or U955 (N_955,N_522,In_906);
nor U956 (N_956,In_611,In_1573);
nor U957 (N_957,In_1747,In_1757);
and U958 (N_958,N_545,N_724);
or U959 (N_959,In_1253,In_1382);
or U960 (N_960,In_888,In_726);
and U961 (N_961,N_603,In_776);
nand U962 (N_962,In_1612,N_617);
nor U963 (N_963,N_621,In_1027);
nand U964 (N_964,N_425,In_2357);
or U965 (N_965,In_1519,N_77);
and U966 (N_966,In_1632,N_555);
xor U967 (N_967,N_347,In_1667);
or U968 (N_968,In_1961,In_523);
nand U969 (N_969,In_140,In_683);
or U970 (N_970,In_1080,In_621);
nor U971 (N_971,N_387,N_458);
xor U972 (N_972,N_739,In_2276);
and U973 (N_973,In_736,In_1720);
nand U974 (N_974,N_574,N_142);
or U975 (N_975,In_2168,N_568);
nor U976 (N_976,In_195,In_207);
and U977 (N_977,In_219,N_488);
xnor U978 (N_978,N_610,N_301);
xor U979 (N_979,In_1912,In_1290);
nor U980 (N_980,N_415,N_688);
or U981 (N_981,N_637,In_1407);
nand U982 (N_982,N_703,N_481);
nand U983 (N_983,N_672,N_643);
or U984 (N_984,In_1342,In_456);
or U985 (N_985,In_1928,In_2097);
nand U986 (N_986,In_1750,In_902);
nand U987 (N_987,N_292,N_450);
xnor U988 (N_988,N_551,In_2356);
and U989 (N_989,N_728,N_715);
nor U990 (N_990,In_2278,In_2308);
nand U991 (N_991,In_2362,In_866);
nor U992 (N_992,N_339,In_1252);
xor U993 (N_993,N_469,N_652);
and U994 (N_994,In_1694,In_1679);
and U995 (N_995,N_445,In_1620);
or U996 (N_996,N_267,N_571);
or U997 (N_997,N_702,In_2206);
and U998 (N_998,N_116,N_206);
nand U999 (N_999,In_1657,In_1433);
nor U1000 (N_1000,N_200,In_1960);
or U1001 (N_1001,N_848,In_246);
or U1002 (N_1002,In_2117,N_429);
xor U1003 (N_1003,N_565,In_1048);
or U1004 (N_1004,In_1946,N_527);
nor U1005 (N_1005,N_278,N_566);
xnor U1006 (N_1006,In_1611,N_80);
nor U1007 (N_1007,In_941,In_91);
or U1008 (N_1008,In_377,N_891);
xnor U1009 (N_1009,In_663,In_1618);
xor U1010 (N_1010,In_1614,In_980);
xor U1011 (N_1011,In_1602,In_1297);
nand U1012 (N_1012,N_112,In_1691);
and U1013 (N_1013,N_681,In_264);
and U1014 (N_1014,N_888,In_1509);
nor U1015 (N_1015,N_974,In_339);
nand U1016 (N_1016,In_362,N_736);
nor U1017 (N_1017,In_670,N_723);
or U1018 (N_1018,In_1484,In_1154);
nand U1019 (N_1019,N_804,N_754);
nand U1020 (N_1020,In_355,N_734);
xnor U1021 (N_1021,In_316,In_721);
nand U1022 (N_1022,N_946,In_1293);
or U1023 (N_1023,In_1883,In_279);
xor U1024 (N_1024,N_397,In_991);
nand U1025 (N_1025,In_846,N_497);
and U1026 (N_1026,N_74,In_1772);
nand U1027 (N_1027,N_514,In_2384);
xnor U1028 (N_1028,N_694,N_823);
xor U1029 (N_1029,In_2478,N_222);
nor U1030 (N_1030,In_1832,N_714);
and U1031 (N_1031,In_940,In_809);
or U1032 (N_1032,N_532,In_65);
nor U1033 (N_1033,N_997,N_850);
and U1034 (N_1034,N_158,N_837);
nor U1035 (N_1035,In_997,N_182);
xor U1036 (N_1036,N_132,In_2355);
or U1037 (N_1037,In_2078,In_1380);
nor U1038 (N_1038,In_1881,N_303);
nand U1039 (N_1039,N_396,In_875);
xnor U1040 (N_1040,In_1231,In_675);
and U1041 (N_1041,N_692,In_372);
and U1042 (N_1042,N_367,In_151);
xor U1043 (N_1043,In_1474,N_788);
and U1044 (N_1044,In_531,In_1592);
and U1045 (N_1045,In_976,N_991);
nand U1046 (N_1046,N_371,In_1346);
or U1047 (N_1047,In_655,N_857);
nand U1048 (N_1048,N_183,N_738);
nand U1049 (N_1049,In_2160,N_151);
and U1050 (N_1050,N_377,In_433);
and U1051 (N_1051,N_385,In_1332);
or U1052 (N_1052,In_460,N_958);
and U1053 (N_1053,In_1959,In_444);
xor U1054 (N_1054,N_757,In_2381);
xnor U1055 (N_1055,In_837,N_356);
nor U1056 (N_1056,N_789,In_965);
or U1057 (N_1057,In_977,In_281);
and U1058 (N_1058,N_460,N_821);
nor U1059 (N_1059,In_2339,N_726);
or U1060 (N_1060,N_871,In_1340);
xnor U1061 (N_1061,In_1938,In_2204);
nand U1062 (N_1062,N_910,In_1751);
nand U1063 (N_1063,In_482,N_874);
nor U1064 (N_1064,In_795,In_1604);
and U1065 (N_1065,In_1787,In_1223);
and U1066 (N_1066,In_758,In_1698);
or U1067 (N_1067,In_44,In_766);
nand U1068 (N_1068,In_1841,In_1308);
xnor U1069 (N_1069,In_561,In_2095);
and U1070 (N_1070,In_245,In_1754);
nor U1071 (N_1071,In_2121,In_2237);
or U1072 (N_1072,N_803,In_62);
and U1073 (N_1073,In_527,In_498);
or U1074 (N_1074,In_267,N_302);
nor U1075 (N_1075,In_2123,N_762);
xor U1076 (N_1076,In_1575,In_1350);
or U1077 (N_1077,In_1741,N_350);
and U1078 (N_1078,In_781,In_1200);
or U1079 (N_1079,N_858,N_774);
and U1080 (N_1080,N_260,N_379);
nand U1081 (N_1081,In_619,In_1123);
nand U1082 (N_1082,In_1623,In_286);
nor U1083 (N_1083,In_1092,In_1191);
or U1084 (N_1084,N_719,In_1528);
nor U1085 (N_1085,In_2010,In_1464);
nand U1086 (N_1086,In_2305,In_179);
nor U1087 (N_1087,In_2202,N_399);
nand U1088 (N_1088,In_2207,In_942);
nor U1089 (N_1089,In_457,In_2017);
or U1090 (N_1090,N_198,In_1094);
or U1091 (N_1091,In_579,N_817);
xor U1092 (N_1092,N_520,N_572);
or U1093 (N_1093,N_337,In_1238);
nand U1094 (N_1094,In_1617,N_859);
nand U1095 (N_1095,N_725,In_1182);
and U1096 (N_1096,In_1075,N_900);
nor U1097 (N_1097,In_835,N_645);
and U1098 (N_1098,In_797,N_423);
nand U1099 (N_1099,In_522,In_1901);
and U1100 (N_1100,In_1002,In_158);
or U1101 (N_1101,In_1338,In_1134);
or U1102 (N_1102,In_772,In_82);
xnor U1103 (N_1103,In_2191,N_845);
and U1104 (N_1104,In_2080,N_214);
nand U1105 (N_1105,N_343,In_354);
or U1106 (N_1106,In_2054,In_877);
xnor U1107 (N_1107,In_881,N_921);
nor U1108 (N_1108,N_811,N_18);
nor U1109 (N_1109,N_790,In_248);
xnor U1110 (N_1110,N_146,N_966);
nor U1111 (N_1111,N_578,N_780);
xnor U1112 (N_1112,In_651,N_750);
nor U1113 (N_1113,In_63,In_231);
and U1114 (N_1114,N_135,In_2375);
xor U1115 (N_1115,N_979,In_586);
or U1116 (N_1116,N_39,N_633);
or U1117 (N_1117,In_1358,In_1590);
nand U1118 (N_1118,N_870,In_1652);
nor U1119 (N_1119,N_984,N_76);
and U1120 (N_1120,In_828,N_710);
and U1121 (N_1121,In_1594,In_261);
nand U1122 (N_1122,N_711,In_783);
and U1123 (N_1123,N_284,In_69);
xor U1124 (N_1124,N_229,N_484);
xor U1125 (N_1125,In_1307,N_935);
nor U1126 (N_1126,N_824,In_46);
or U1127 (N_1127,In_960,N_644);
nand U1128 (N_1128,N_67,In_509);
xnor U1129 (N_1129,In_1030,N_163);
nand U1130 (N_1130,N_620,In_216);
nand U1131 (N_1131,In_841,In_2440);
and U1132 (N_1132,N_444,N_700);
nor U1133 (N_1133,In_399,N_657);
nor U1134 (N_1134,In_1507,In_2197);
xor U1135 (N_1135,In_346,N_434);
or U1136 (N_1136,In_1712,In_810);
xnor U1137 (N_1137,In_2328,N_523);
nand U1138 (N_1138,In_1486,N_207);
xnor U1139 (N_1139,In_275,N_143);
nor U1140 (N_1140,N_328,In_500);
nand U1141 (N_1141,In_879,In_1866);
xnor U1142 (N_1142,N_994,In_1451);
and U1143 (N_1143,In_939,N_590);
nor U1144 (N_1144,N_922,N_701);
and U1145 (N_1145,N_630,N_244);
and U1146 (N_1146,N_976,In_1168);
or U1147 (N_1147,In_1777,In_2155);
nor U1148 (N_1148,In_1139,In_1524);
and U1149 (N_1149,N_964,In_1858);
and U1150 (N_1150,In_99,In_1353);
xor U1151 (N_1151,N_552,In_1362);
xnor U1152 (N_1152,N_480,In_1647);
or U1153 (N_1153,N_882,In_1983);
and U1154 (N_1154,N_84,In_1806);
nand U1155 (N_1155,In_6,N_775);
and U1156 (N_1156,In_1799,In_1921);
nand U1157 (N_1157,N_920,In_360);
xnor U1158 (N_1158,N_608,N_127);
nand U1159 (N_1159,N_259,In_344);
nor U1160 (N_1160,N_557,In_192);
and U1161 (N_1161,N_805,N_395);
or U1162 (N_1162,In_2260,In_1993);
nand U1163 (N_1163,In_2055,In_108);
nor U1164 (N_1164,In_664,In_24);
and U1165 (N_1165,In_1535,In_1815);
and U1166 (N_1166,In_2021,In_1214);
nor U1167 (N_1167,N_69,In_411);
and U1168 (N_1168,In_149,In_191);
or U1169 (N_1169,In_1319,In_601);
xor U1170 (N_1170,In_2145,In_1562);
nor U1171 (N_1171,N_191,N_536);
and U1172 (N_1172,In_204,In_714);
xor U1173 (N_1173,In_2336,In_2147);
and U1174 (N_1174,In_2019,N_264);
xor U1175 (N_1175,In_190,N_554);
nor U1176 (N_1176,In_1788,In_1371);
or U1177 (N_1177,N_912,N_800);
xnor U1178 (N_1178,In_203,N_389);
nor U1179 (N_1179,N_795,In_1737);
xor U1180 (N_1180,In_43,In_1768);
or U1181 (N_1181,In_2393,In_2458);
or U1182 (N_1182,N_902,N_853);
and U1183 (N_1183,N_558,N_466);
xor U1184 (N_1184,In_1076,In_1542);
or U1185 (N_1185,N_836,N_587);
or U1186 (N_1186,N_40,In_1790);
xnor U1187 (N_1187,N_985,In_2171);
or U1188 (N_1188,In_679,In_738);
or U1189 (N_1189,In_181,N_956);
or U1190 (N_1190,In_1584,In_2386);
nand U1191 (N_1191,N_254,In_491);
nand U1192 (N_1192,N_872,In_894);
nor U1193 (N_1193,In_1077,N_895);
nor U1194 (N_1194,N_901,In_1574);
xnor U1195 (N_1195,N_211,N_87);
xor U1196 (N_1196,In_208,In_1066);
nand U1197 (N_1197,In_1194,N_416);
or U1198 (N_1198,In_1701,In_2291);
or U1199 (N_1199,N_186,N_733);
xnor U1200 (N_1200,N_796,N_851);
nor U1201 (N_1201,N_599,In_2402);
xor U1202 (N_1202,N_713,In_575);
nand U1203 (N_1203,N_842,N_210);
nand U1204 (N_1204,N_453,N_860);
nor U1205 (N_1205,N_381,In_1284);
and U1206 (N_1206,In_2127,In_84);
nor U1207 (N_1207,N_516,In_1328);
and U1208 (N_1208,In_2403,In_135);
or U1209 (N_1209,In_1743,N_584);
and U1210 (N_1210,N_157,N_990);
xnor U1211 (N_1211,N_304,N_169);
and U1212 (N_1212,In_7,N_71);
nor U1213 (N_1213,In_2296,In_1054);
nand U1214 (N_1214,In_1101,N_300);
nand U1215 (N_1215,N_496,In_2101);
nor U1216 (N_1216,N_685,In_2284);
and U1217 (N_1217,In_271,In_713);
or U1218 (N_1218,In_1515,In_2366);
xor U1219 (N_1219,N_433,In_2495);
or U1220 (N_1220,In_646,N_556);
and U1221 (N_1221,In_610,In_1202);
nor U1222 (N_1222,N_154,In_1871);
or U1223 (N_1223,In_1953,N_813);
and U1224 (N_1224,In_276,In_464);
xor U1225 (N_1225,In_854,N_751);
nand U1226 (N_1226,N_109,N_325);
nor U1227 (N_1227,In_374,In_1512);
nand U1228 (N_1228,N_139,In_872);
nand U1229 (N_1229,In_516,In_831);
and U1230 (N_1230,In_644,N_611);
xor U1231 (N_1231,In_157,N_676);
and U1232 (N_1232,In_895,N_521);
and U1233 (N_1233,In_120,In_1635);
nand U1234 (N_1234,In_2131,N_564);
xnor U1235 (N_1235,N_263,In_1730);
nand U1236 (N_1236,N_329,N_883);
xnor U1237 (N_1237,In_793,N_945);
or U1238 (N_1238,N_586,In_1198);
or U1239 (N_1239,In_2018,N_778);
xnor U1240 (N_1240,In_1990,N_333);
nor U1241 (N_1241,In_64,In_949);
xor U1242 (N_1242,In_479,In_1774);
nor U1243 (N_1243,In_507,In_2449);
xnor U1244 (N_1244,N_406,N_593);
nand U1245 (N_1245,N_787,N_529);
nand U1246 (N_1246,N_934,In_1414);
nand U1247 (N_1247,N_838,N_345);
or U1248 (N_1248,In_353,In_1281);
and U1249 (N_1249,In_1193,N_918);
and U1250 (N_1250,In_2448,In_1521);
or U1251 (N_1251,N_1196,N_712);
or U1252 (N_1252,In_1664,In_727);
xor U1253 (N_1253,N_889,In_899);
xor U1254 (N_1254,In_660,In_305);
xor U1255 (N_1255,N_886,N_258);
and U1256 (N_1256,N_1016,N_357);
or U1257 (N_1257,In_409,In_418);
or U1258 (N_1258,N_1110,N_398);
or U1259 (N_1259,In_815,N_1148);
or U1260 (N_1260,In_874,In_1256);
nor U1261 (N_1261,N_786,N_943);
nand U1262 (N_1262,In_2182,N_1041);
nor U1263 (N_1263,N_830,N_476);
nor U1264 (N_1264,In_751,In_806);
or U1265 (N_1265,N_1235,In_948);
or U1266 (N_1266,In_1710,N_1084);
and U1267 (N_1267,N_1071,In_451);
nand U1268 (N_1268,N_826,In_1675);
and U1269 (N_1269,In_2215,In_321);
nand U1270 (N_1270,In_1295,N_833);
and U1271 (N_1271,N_147,In_1455);
and U1272 (N_1272,N_1143,N_1161);
and U1273 (N_1273,In_1012,N_770);
xor U1274 (N_1274,In_1439,In_957);
or U1275 (N_1275,In_741,In_1105);
xnor U1276 (N_1276,In_554,N_1028);
or U1277 (N_1277,In_1091,In_2173);
and U1278 (N_1278,N_1173,N_898);
nor U1279 (N_1279,In_2473,N_468);
and U1280 (N_1280,In_1449,In_1842);
or U1281 (N_1281,In_161,In_1083);
nand U1282 (N_1282,N_6,N_1170);
and U1283 (N_1283,N_1103,In_1857);
nand U1284 (N_1284,N_1099,In_434);
xnor U1285 (N_1285,In_2426,N_972);
nand U1286 (N_1286,In_1673,In_845);
and U1287 (N_1287,N_876,In_2314);
or U1288 (N_1288,In_11,In_2023);
nor U1289 (N_1289,In_1031,In_2099);
and U1290 (N_1290,In_749,In_545);
or U1291 (N_1291,In_2076,In_1823);
xnor U1292 (N_1292,N_201,N_509);
and U1293 (N_1293,N_1091,N_1021);
nor U1294 (N_1294,In_1514,In_633);
nor U1295 (N_1295,In_2488,N_1083);
nor U1296 (N_1296,N_463,N_783);
or U1297 (N_1297,N_828,In_1776);
or U1298 (N_1298,In_1244,N_846);
and U1299 (N_1299,N_944,N_335);
and U1300 (N_1300,In_963,In_1605);
xor U1301 (N_1301,N_1152,In_2081);
xor U1302 (N_1302,N_1125,N_767);
xor U1303 (N_1303,N_178,In_915);
xnor U1304 (N_1304,In_2334,In_1513);
nor U1305 (N_1305,N_525,In_677);
and U1306 (N_1306,In_969,In_188);
nand U1307 (N_1307,In_74,N_59);
or U1308 (N_1308,N_1195,In_393);
xnor U1309 (N_1309,In_774,N_221);
nand U1310 (N_1310,N_699,N_1105);
or U1311 (N_1311,In_1438,N_793);
nand U1312 (N_1312,In_1203,N_1027);
or U1313 (N_1313,N_1214,N_531);
xor U1314 (N_1314,N_1158,In_2301);
and U1315 (N_1315,In_1351,In_722);
xnor U1316 (N_1316,In_1333,In_18);
and U1317 (N_1317,N_1060,N_280);
or U1318 (N_1318,In_1510,N_17);
or U1319 (N_1319,N_963,N_973);
or U1320 (N_1320,N_360,In_2474);
and U1321 (N_1321,N_905,N_1127);
and U1322 (N_1322,In_649,N_756);
nor U1323 (N_1323,N_735,In_1554);
nand U1324 (N_1324,N_806,N_277);
and U1325 (N_1325,In_2141,N_1096);
nand U1326 (N_1326,N_307,N_1058);
or U1327 (N_1327,N_305,In_312);
nand U1328 (N_1328,N_1093,N_1070);
or U1329 (N_1329,N_998,N_971);
and U1330 (N_1330,N_760,N_960);
or U1331 (N_1331,N_1039,In_2034);
or U1332 (N_1332,N_752,N_30);
or U1333 (N_1333,In_757,In_1552);
nand U1334 (N_1334,N_1151,In_2481);
nor U1335 (N_1335,In_2380,In_2462);
or U1336 (N_1336,N_230,N_576);
or U1337 (N_1337,N_352,N_1085);
nor U1338 (N_1338,N_1216,N_212);
nor U1339 (N_1339,In_378,N_949);
nor U1340 (N_1340,In_1052,N_113);
or U1341 (N_1341,N_588,N_666);
or U1342 (N_1342,In_379,In_252);
and U1343 (N_1343,In_2216,N_822);
and U1344 (N_1344,N_948,N_1063);
or U1345 (N_1345,N_977,In_287);
nor U1346 (N_1346,N_589,In_26);
and U1347 (N_1347,In_2383,N_1220);
and U1348 (N_1348,In_2385,N_1086);
xor U1349 (N_1349,In_930,In_86);
or U1350 (N_1350,N_23,N_880);
nor U1351 (N_1351,N_799,N_1182);
and U1352 (N_1352,N_9,In_1965);
nand U1353 (N_1353,In_2223,N_5);
nor U1354 (N_1354,N_316,In_2377);
nor U1355 (N_1355,In_2189,N_635);
and U1356 (N_1356,N_1053,N_507);
and U1357 (N_1357,N_298,In_134);
nand U1358 (N_1358,In_1553,N_159);
and U1359 (N_1359,In_415,In_504);
and U1360 (N_1360,In_2239,N_947);
xor U1361 (N_1361,N_1040,N_1019);
nor U1362 (N_1362,N_1238,N_849);
and U1363 (N_1363,N_121,N_1030);
or U1364 (N_1364,N_791,In_1825);
or U1365 (N_1365,In_1147,N_380);
xnor U1366 (N_1366,N_1192,In_994);
xnor U1367 (N_1367,N_1226,N_1012);
nor U1368 (N_1368,N_128,In_1421);
or U1369 (N_1369,In_2337,N_969);
xor U1370 (N_1370,In_549,N_1094);
nand U1371 (N_1371,N_1136,In_2177);
xor U1372 (N_1372,In_101,In_572);
or U1373 (N_1373,N_996,In_1493);
or U1374 (N_1374,N_687,N_101);
or U1375 (N_1375,N_684,N_1133);
and U1376 (N_1376,N_907,N_640);
and U1377 (N_1377,N_1176,N_717);
nor U1378 (N_1378,In_737,N_14);
or U1379 (N_1379,N_1097,In_162);
nor U1380 (N_1380,In_2106,N_814);
or U1381 (N_1381,In_2011,N_249);
nor U1382 (N_1382,N_506,In_1973);
and U1383 (N_1383,In_560,In_1818);
and U1384 (N_1384,N_409,In_2205);
xnor U1385 (N_1385,In_1339,In_883);
nor U1386 (N_1386,N_868,In_384);
nor U1387 (N_1387,In_1305,In_2104);
xnor U1388 (N_1388,In_1300,In_1216);
xnor U1389 (N_1389,In_615,N_541);
or U1390 (N_1390,In_177,In_750);
and U1391 (N_1391,N_591,In_1085);
nor U1392 (N_1392,N_1034,In_628);
xnor U1393 (N_1393,N_1159,In_2073);
and U1394 (N_1394,In_2497,In_1132);
or U1395 (N_1395,N_518,N_706);
xnor U1396 (N_1396,In_2320,In_1263);
and U1397 (N_1397,In_925,N_797);
or U1398 (N_1398,N_1044,N_878);
nor U1399 (N_1399,N_1171,N_854);
or U1400 (N_1400,N_10,In_1997);
or U1401 (N_1401,N_965,In_1494);
nand U1402 (N_1402,N_818,N_441);
nor U1403 (N_1403,In_1118,N_890);
and U1404 (N_1404,N_491,N_257);
or U1405 (N_1405,N_311,In_789);
and U1406 (N_1406,N_1209,N_437);
xor U1407 (N_1407,In_2480,In_1873);
xor U1408 (N_1408,N_1140,In_1969);
nand U1409 (N_1409,In_1821,In_587);
and U1410 (N_1410,In_728,N_741);
or U1411 (N_1411,In_697,In_1622);
xor U1412 (N_1412,In_2024,In_2313);
nand U1413 (N_1413,N_1199,In_70);
xnor U1414 (N_1414,In_567,N_1179);
and U1415 (N_1415,N_1198,N_1010);
nand U1416 (N_1416,In_811,N_1211);
nor U1417 (N_1417,N_1227,N_1123);
or U1418 (N_1418,In_2406,In_200);
xnor U1419 (N_1419,In_1532,N_457);
xor U1420 (N_1420,N_829,In_2496);
or U1421 (N_1421,N_185,In_1995);
and U1422 (N_1422,N_376,N_906);
or U1423 (N_1423,In_229,N_1088);
or U1424 (N_1424,In_132,N_697);
and U1425 (N_1425,N_1218,N_746);
nand U1426 (N_1426,N_899,In_2363);
or U1427 (N_1427,In_1530,N_1118);
and U1428 (N_1428,N_1124,N_544);
nor U1429 (N_1429,N_274,N_362);
nand U1430 (N_1430,In_414,In_2040);
nand U1431 (N_1431,N_171,N_1001);
xor U1432 (N_1432,N_675,In_356);
and U1433 (N_1433,In_1779,N_825);
nor U1434 (N_1434,N_1121,In_499);
nand U1435 (N_1435,In_2475,In_1040);
xnor U1436 (N_1436,In_2194,N_1128);
and U1437 (N_1437,In_1833,N_330);
and U1438 (N_1438,N_929,N_269);
and U1439 (N_1439,N_856,In_369);
and U1440 (N_1440,N_908,N_513);
or U1441 (N_1441,N_534,In_868);
nand U1442 (N_1442,N_884,In_718);
nand U1443 (N_1443,N_1200,In_1578);
xor U1444 (N_1444,N_616,N_819);
nand U1445 (N_1445,N_932,N_1059);
xor U1446 (N_1446,N_916,N_771);
nor U1447 (N_1447,In_391,In_653);
and U1448 (N_1448,N_1102,N_1106);
or U1449 (N_1449,N_1082,N_598);
nor U1450 (N_1450,N_749,In_437);
nor U1451 (N_1451,In_2196,N_1022);
and U1452 (N_1452,In_944,In_297);
and U1453 (N_1453,In_48,N_1080);
and U1454 (N_1454,N_1073,In_424);
xnor U1455 (N_1455,In_13,In_1279);
nor U1456 (N_1456,In_2157,In_1366);
nor U1457 (N_1457,In_1610,In_922);
and U1458 (N_1458,N_631,In_125);
xnor U1459 (N_1459,N_975,In_975);
or U1460 (N_1460,N_1210,In_605);
nor U1461 (N_1461,N_1150,In_788);
nor U1462 (N_1462,N_915,In_1068);
xor U1463 (N_1463,N_512,In_799);
nand U1464 (N_1464,N_832,N_928);
or U1465 (N_1465,N_193,In_497);
nand U1466 (N_1466,N_1206,N_383);
nand U1467 (N_1467,In_358,In_439);
xnor U1468 (N_1468,N_855,N_1248);
and U1469 (N_1469,N_1122,N_1077);
nand U1470 (N_1470,N_405,N_487);
or U1471 (N_1471,N_801,In_115);
nand U1472 (N_1472,N_954,In_1707);
nand U1473 (N_1473,N_1228,N_1219);
xor U1474 (N_1474,N_1202,N_747);
or U1475 (N_1475,N_1147,N_993);
nand U1476 (N_1476,In_1685,N_923);
or U1477 (N_1477,In_1103,N_1184);
nor U1478 (N_1478,N_1240,N_1190);
nor U1479 (N_1479,N_160,In_598);
or U1480 (N_1480,In_1025,In_1872);
nand U1481 (N_1481,N_709,In_1522);
nand U1482 (N_1482,In_747,N_769);
and U1483 (N_1483,In_1187,In_840);
xor U1484 (N_1484,N_63,In_821);
and U1485 (N_1485,N_1007,In_755);
xnor U1486 (N_1486,N_1052,N_1108);
nor U1487 (N_1487,N_197,In_2272);
or U1488 (N_1488,N_785,In_2303);
nand U1489 (N_1489,N_671,N_1186);
nor U1490 (N_1490,N_1113,N_1006);
and U1491 (N_1491,In_1065,In_613);
or U1492 (N_1492,N_61,In_1878);
and U1493 (N_1493,In_1024,In_1567);
nand U1494 (N_1494,N_99,In_1176);
xnor U1495 (N_1495,N_1089,In_39);
nand U1496 (N_1496,In_2421,In_1327);
and U1497 (N_1497,In_2052,In_863);
nor U1498 (N_1498,N_402,In_1798);
xor U1499 (N_1499,N_1130,In_2441);
nor U1500 (N_1500,N_744,N_816);
and U1501 (N_1501,N_1051,N_1243);
and U1502 (N_1502,N_642,N_1245);
xor U1503 (N_1503,N_1185,N_452);
xnor U1504 (N_1504,N_1055,N_1275);
or U1505 (N_1505,N_1323,N_1388);
and U1506 (N_1506,In_1046,N_1359);
or U1507 (N_1507,In_1087,In_1830);
and U1508 (N_1508,N_1075,In_546);
nand U1509 (N_1509,N_1347,N_1327);
nor U1510 (N_1510,In_170,N_1046);
nand U1511 (N_1511,N_86,N_1419);
or U1512 (N_1512,N_1333,N_1242);
xnor U1513 (N_1513,In_428,In_695);
nand U1514 (N_1514,N_1467,In_1555);
nand U1515 (N_1515,In_301,N_718);
and U1516 (N_1516,N_1390,N_863);
and U1517 (N_1517,In_1683,N_332);
nand U1518 (N_1518,N_1222,In_2477);
xor U1519 (N_1519,In_1423,N_1104);
and U1520 (N_1520,N_60,In_603);
and U1521 (N_1521,N_1068,N_677);
or U1522 (N_1522,N_1404,In_832);
or U1523 (N_1523,N_1141,N_867);
or U1524 (N_1524,N_716,N_1290);
xnor U1525 (N_1525,In_2240,In_1511);
nand U1526 (N_1526,N_1295,In_138);
and U1527 (N_1527,In_672,In_392);
and U1528 (N_1528,In_823,N_1344);
and U1529 (N_1529,N_1278,In_1595);
nand U1530 (N_1530,N_740,N_619);
nor U1531 (N_1531,N_1294,N_913);
nand U1532 (N_1532,N_309,In_327);
nor U1533 (N_1533,N_1066,In_2185);
or U1534 (N_1534,In_1323,In_1090);
and U1535 (N_1535,N_1334,In_1708);
nor U1536 (N_1536,In_867,N_1225);
xnor U1537 (N_1537,In_66,N_95);
nor U1538 (N_1538,N_539,In_315);
nor U1539 (N_1539,N_1301,N_970);
nand U1540 (N_1540,N_1336,In_1172);
nand U1541 (N_1541,N_1326,In_197);
or U1542 (N_1542,N_1135,N_194);
nor U1543 (N_1543,N_961,N_1385);
and U1544 (N_1544,N_299,N_184);
xor U1545 (N_1545,N_1191,N_897);
and U1546 (N_1546,In_336,N_1160);
nand U1547 (N_1547,N_53,N_670);
nor U1548 (N_1548,In_953,N_1455);
nor U1549 (N_1549,N_705,In_1943);
xnor U1550 (N_1550,In_642,In_2166);
nand U1551 (N_1551,In_77,In_490);
nand U1552 (N_1552,N_1298,In_474);
and U1553 (N_1553,N_1405,N_1236);
and U1554 (N_1554,N_1485,N_776);
and U1555 (N_1555,In_244,N_1484);
and U1556 (N_1556,N_1306,In_1440);
nor U1557 (N_1557,N_1213,N_1069);
nor U1558 (N_1558,N_1436,N_843);
xnor U1559 (N_1559,In_2214,N_1024);
or U1560 (N_1560,In_1568,In_148);
and U1561 (N_1561,N_1346,N_1362);
nand U1562 (N_1562,N_1233,N_1407);
nand U1563 (N_1563,In_1839,In_1911);
or U1564 (N_1564,N_1036,N_607);
and U1565 (N_1565,N_995,N_375);
or U1566 (N_1566,In_2038,N_1338);
or U1567 (N_1567,N_1189,N_1394);
and U1568 (N_1568,N_1343,N_885);
nand U1569 (N_1569,N_1215,N_1074);
xor U1570 (N_1570,N_879,N_865);
or U1571 (N_1571,N_1244,N_982);
or U1572 (N_1572,N_238,In_1292);
or U1573 (N_1573,N_1307,N_394);
nor U1574 (N_1574,N_1495,N_349);
nand U1575 (N_1575,In_1116,In_2174);
nor U1576 (N_1576,N_758,N_403);
nor U1577 (N_1577,N_904,N_1029);
or U1578 (N_1578,In_2427,N_1247);
or U1579 (N_1579,In_2289,N_1462);
or U1580 (N_1580,N_1329,In_950);
nor U1581 (N_1581,N_933,N_1156);
nor U1582 (N_1582,In_1431,In_1989);
and U1583 (N_1583,In_373,N_1285);
and U1584 (N_1584,N_647,N_82);
nor U1585 (N_1585,N_1061,N_1175);
nor U1586 (N_1586,N_124,N_1350);
xnor U1587 (N_1587,In_2463,N_37);
nand U1588 (N_1588,N_1435,In_891);
nand U1589 (N_1589,N_1239,In_22);
or U1590 (N_1590,N_1486,N_465);
nor U1591 (N_1591,N_1157,N_88);
nor U1592 (N_1592,N_937,In_1088);
nor U1593 (N_1593,N_388,In_1250);
nor U1594 (N_1594,In_773,N_1270);
and U1595 (N_1595,In_2027,N_1470);
and U1596 (N_1596,N_981,In_1352);
or U1597 (N_1597,In_2396,In_1480);
xor U1598 (N_1598,N_1360,In_954);
nand U1599 (N_1599,N_495,In_1272);
or U1600 (N_1600,N_1457,In_2110);
nand U1601 (N_1601,N_917,In_802);
or U1602 (N_1602,N_41,In_2139);
or U1603 (N_1603,N_1138,In_659);
or U1604 (N_1604,In_2365,In_55);
or U1605 (N_1605,N_251,N_196);
and U1606 (N_1606,In_2349,In_1115);
nor U1607 (N_1607,N_477,N_1000);
or U1608 (N_1608,N_1383,N_472);
xor U1609 (N_1609,N_1255,N_881);
xor U1610 (N_1610,In_1234,N_1365);
nand U1611 (N_1611,N_1440,N_1273);
nor U1612 (N_1612,In_2045,In_21);
or U1613 (N_1613,N_1471,N_1288);
nor U1614 (N_1614,N_808,N_1309);
xnor U1615 (N_1615,N_474,N_731);
xor U1616 (N_1616,In_666,N_1048);
xor U1617 (N_1617,In_1543,N_1092);
xnor U1618 (N_1618,N_1208,In_929);
nor U1619 (N_1619,N_1487,N_1087);
nor U1620 (N_1620,N_1392,N_1476);
or U1621 (N_1621,In_2013,In_952);
and U1622 (N_1622,N_779,N_45);
nor U1623 (N_1623,N_748,N_798);
nand U1624 (N_1624,In_1427,N_1237);
xnor U1625 (N_1625,N_1480,N_346);
and U1626 (N_1626,In_173,N_1400);
or U1627 (N_1627,N_1032,N_1090);
xor U1628 (N_1628,N_1361,In_847);
nor U1629 (N_1629,N_1406,In_2438);
nor U1630 (N_1630,N_489,N_766);
xor U1631 (N_1631,In_2135,In_1678);
xor U1632 (N_1632,In_1375,N_1076);
xor U1633 (N_1633,N_810,N_537);
nand U1634 (N_1634,N_1109,N_1339);
xnor U1635 (N_1635,In_2409,In_962);
or U1636 (N_1636,N_287,N_602);
and U1637 (N_1637,N_1315,N_1155);
nand U1638 (N_1638,N_931,N_841);
or U1639 (N_1639,N_1493,N_505);
and U1640 (N_1640,In_2247,N_1217);
xnor U1641 (N_1641,In_417,N_1351);
or U1642 (N_1642,N_1421,N_1296);
or U1643 (N_1643,N_978,In_1884);
nor U1644 (N_1644,N_25,N_794);
xor U1645 (N_1645,N_1310,N_1448);
or U1646 (N_1646,In_1229,N_1107);
nand U1647 (N_1647,N_1356,N_473);
xnor U1648 (N_1648,In_2225,N_1477);
nand U1649 (N_1649,In_1572,N_1037);
xnor U1650 (N_1650,N_1165,N_689);
xor U1651 (N_1651,N_567,N_1129);
or U1652 (N_1652,N_1414,N_1302);
and U1653 (N_1653,N_553,N_1300);
xnor U1654 (N_1654,N_1095,N_951);
and U1655 (N_1655,N_1342,In_2275);
or U1656 (N_1656,N_1119,In_283);
xnor U1657 (N_1657,N_580,N_892);
xnor U1658 (N_1658,In_461,N_663);
nor U1659 (N_1659,N_1317,In_2281);
nor U1660 (N_1660,N_656,N_1320);
nand U1661 (N_1661,N_761,In_1729);
or U1662 (N_1662,In_247,In_2005);
and U1663 (N_1663,N_614,N_1374);
nor U1664 (N_1664,N_1035,In_307);
and U1665 (N_1665,N_1429,In_95);
or U1666 (N_1666,N_1411,N_1201);
nand U1667 (N_1667,N_459,N_1100);
xor U1668 (N_1668,N_1271,N_930);
nor U1669 (N_1669,In_2035,N_1494);
xor U1670 (N_1670,N_743,N_1398);
nand U1671 (N_1671,N_847,N_893);
or U1672 (N_1672,In_407,In_469);
xnor U1673 (N_1673,In_133,In_1716);
and U1674 (N_1674,In_367,N_1177);
nor U1675 (N_1675,N_1376,In_226);
or U1676 (N_1676,N_809,N_1409);
nand U1677 (N_1677,In_436,N_831);
or U1678 (N_1678,In_375,N_1331);
xnor U1679 (N_1679,N_1131,N_1410);
or U1680 (N_1680,N_348,In_1206);
xnor U1681 (N_1681,N_1266,N_1451);
nand U1682 (N_1682,N_869,In_295);
or U1683 (N_1683,N_562,In_2348);
nor U1684 (N_1684,In_102,N_1162);
xor U1685 (N_1685,In_363,In_2050);
nor U1686 (N_1686,N_549,N_1038);
nand U1687 (N_1687,In_1357,In_803);
nor U1688 (N_1688,N_1305,N_1241);
nand U1689 (N_1689,N_515,In_2304);
and U1690 (N_1690,N_938,N_988);
or U1691 (N_1691,N_1281,N_1496);
nor U1692 (N_1692,N_502,N_693);
and U1693 (N_1693,In_71,In_2036);
and U1694 (N_1694,N_430,In_2417);
nand U1695 (N_1695,In_282,N_1437);
and U1696 (N_1696,N_1422,N_1205);
or U1697 (N_1697,N_1252,N_628);
and U1698 (N_1698,N_987,In_1110);
or U1699 (N_1699,N_1489,N_141);
nand U1700 (N_1700,N_781,In_1201);
nor U1701 (N_1701,In_740,N_1375);
xor U1702 (N_1702,N_1464,In_2499);
nor U1703 (N_1703,N_807,N_1491);
xnor U1704 (N_1704,N_583,N_894);
nor U1705 (N_1705,N_1004,N_1445);
xnor U1706 (N_1706,N_1279,In_476);
xnor U1707 (N_1707,In_559,In_861);
nand U1708 (N_1708,N_1438,N_1416);
nor U1709 (N_1709,N_1426,In_28);
xor U1710 (N_1710,N_1337,N_1452);
nor U1711 (N_1711,N_508,In_1225);
or U1712 (N_1712,In_1028,In_1394);
and U1713 (N_1713,N_903,N_503);
and U1714 (N_1714,In_1503,N_1231);
xnor U1715 (N_1715,N_289,N_1137);
nand U1716 (N_1716,N_492,N_1254);
xnor U1717 (N_1717,In_2439,N_759);
nor U1718 (N_1718,In_1980,N_547);
or U1719 (N_1719,In_973,N_517);
or U1720 (N_1720,N_239,N_1458);
and U1721 (N_1721,In_2299,N_315);
nand U1722 (N_1722,N_1292,N_1002);
nand U1723 (N_1723,N_925,N_624);
xnor U1724 (N_1724,N_840,N_835);
nor U1725 (N_1725,N_777,In_1599);
or U1726 (N_1726,In_634,N_1319);
xor U1727 (N_1727,N_1149,In_1034);
or U1728 (N_1728,N_1293,N_1072);
and U1729 (N_1729,N_1197,In_1022);
nand U1730 (N_1730,N_1047,N_623);
nand U1731 (N_1731,In_2416,N_1322);
or U1732 (N_1732,In_1627,In_156);
nor U1733 (N_1733,N_968,N_896);
nor U1734 (N_1734,N_1482,N_844);
nor U1735 (N_1735,N_955,In_288);
or U1736 (N_1736,N_604,N_1018);
nand U1737 (N_1737,N_612,N_980);
nand U1738 (N_1738,N_1490,N_1427);
xor U1739 (N_1739,In_1001,N_546);
and U1740 (N_1740,N_753,In_1497);
nand U1741 (N_1741,In_2486,In_1910);
nor U1742 (N_1742,N_1304,N_1297);
nand U1743 (N_1743,In_2246,N_704);
nand U1744 (N_1744,In_681,In_1822);
or U1745 (N_1745,N_368,In_1870);
nand U1746 (N_1746,N_1269,In_2001);
nand U1747 (N_1747,N_1370,In_2262);
and U1748 (N_1748,N_679,In_1276);
nand U1749 (N_1749,N_941,N_177);
nor U1750 (N_1750,N_1276,N_1634);
and U1751 (N_1751,N_1511,N_1594);
nand U1752 (N_1752,N_1614,N_1335);
nor U1753 (N_1753,N_1629,In_441);
and U1754 (N_1754,N_1067,N_1396);
and U1755 (N_1755,N_1504,N_1503);
or U1756 (N_1756,N_1580,N_1677);
nor U1757 (N_1757,N_1586,In_2467);
nand U1758 (N_1758,N_1249,N_575);
or U1759 (N_1759,In_1985,In_1128);
and U1760 (N_1760,N_962,N_1715);
nand U1761 (N_1761,N_1683,N_1613);
and U1762 (N_1762,N_926,N_1546);
nor U1763 (N_1763,In_1903,N_986);
nand U1764 (N_1764,N_1747,In_2109);
and U1765 (N_1765,N_530,N_1609);
or U1766 (N_1766,N_1741,N_1732);
or U1767 (N_1767,N_1532,N_1558);
and U1768 (N_1768,N_1686,N_983);
and U1769 (N_1769,In_1812,In_2068);
nand U1770 (N_1770,N_1508,N_1043);
xnor U1771 (N_1771,N_1193,In_588);
or U1772 (N_1772,In_2181,In_1942);
or U1773 (N_1773,N_1563,N_1519);
nor U1774 (N_1774,N_1665,In_1437);
and U1775 (N_1775,N_1497,N_1540);
xor U1776 (N_1776,N_1,In_856);
nand U1777 (N_1777,N_1251,N_1737);
xor U1778 (N_1778,N_1703,N_1627);
and U1779 (N_1779,N_1167,In_2079);
or U1780 (N_1780,N_1569,N_1013);
and U1781 (N_1781,N_418,N_695);
nor U1782 (N_1782,N_1535,In_607);
nor U1783 (N_1783,N_1657,N_1740);
or U1784 (N_1784,N_1723,N_1433);
xor U1785 (N_1785,N_763,In_1359);
or U1786 (N_1786,In_1100,N_1221);
nand U1787 (N_1787,In_2096,N_1020);
nor U1788 (N_1788,N_511,N_1551);
nor U1789 (N_1789,N_1314,In_536);
and U1790 (N_1790,N_1585,N_1264);
and U1791 (N_1791,N_1364,N_1605);
nand U1792 (N_1792,N_1229,N_1660);
xor U1793 (N_1793,N_1166,N_563);
xor U1794 (N_1794,N_1262,N_1702);
and U1795 (N_1795,N_1547,N_1461);
nand U1796 (N_1796,N_1472,N_1636);
and U1797 (N_1797,N_1582,In_2412);
or U1798 (N_1798,N_1291,N_1111);
nand U1799 (N_1799,In_2236,N_1724);
nor U1800 (N_1800,In_1982,N_427);
or U1801 (N_1801,N_1510,N_1670);
or U1802 (N_1802,N_432,N_914);
and U1803 (N_1803,N_1420,N_85);
or U1804 (N_1804,N_1379,N_1666);
xor U1805 (N_1805,N_1134,N_366);
nor U1806 (N_1806,N_924,N_1712);
and U1807 (N_1807,N_936,In_146);
or U1808 (N_1808,N_110,In_2261);
and U1809 (N_1809,N_1126,N_404);
nor U1810 (N_1810,N_1194,N_1685);
and U1811 (N_1811,N_665,N_1009);
or U1812 (N_1812,N_1548,N_641);
and U1813 (N_1813,N_1742,N_1710);
nor U1814 (N_1814,N_1498,In_2208);
nor U1815 (N_1815,In_2277,In_1588);
nand U1816 (N_1816,N_1473,N_1526);
or U1817 (N_1817,N_1469,In_1714);
nor U1818 (N_1818,In_112,N_1353);
and U1819 (N_1819,In_1597,N_461);
and U1820 (N_1820,N_1349,N_764);
xor U1821 (N_1821,In_1482,N_1223);
xor U1822 (N_1822,In_1665,N_1735);
or U1823 (N_1823,N_1524,N_535);
xor U1824 (N_1824,N_1687,N_1705);
or U1825 (N_1825,N_1050,N_1543);
and U1826 (N_1826,N_1624,N_1465);
nor U1827 (N_1827,In_1569,N_1054);
or U1828 (N_1828,In_1837,N_1516);
nand U1829 (N_1829,N_1397,N_1224);
nand U1830 (N_1830,N_1651,N_1599);
xnor U1831 (N_1831,In_569,N_1232);
xor U1832 (N_1832,N_1479,N_1549);
and U1833 (N_1833,N_1533,In_2007);
and U1834 (N_1834,N_1014,N_1286);
xor U1835 (N_1835,N_1324,In_1547);
and U1836 (N_1836,N_661,N_231);
xnor U1837 (N_1837,N_1691,N_1707);
or U1838 (N_1838,N_967,N_1234);
nand U1839 (N_1839,N_1261,N_989);
and U1840 (N_1840,In_1313,N_351);
nor U1841 (N_1841,N_1632,N_1415);
xor U1842 (N_1842,N_634,N_839);
and U1843 (N_1843,N_279,N_1428);
or U1844 (N_1844,In_334,N_768);
nand U1845 (N_1845,In_1860,N_1449);
or U1846 (N_1846,In_1700,N_1562);
nand U1847 (N_1847,N_609,N_1635);
and U1848 (N_1848,N_1537,N_1717);
or U1849 (N_1849,N_1507,N_1023);
or U1850 (N_1850,N_1572,N_654);
nor U1851 (N_1851,N_1432,N_1530);
or U1852 (N_1852,N_15,N_118);
nand U1853 (N_1853,N_1492,N_475);
nor U1854 (N_1854,N_1719,N_1697);
nor U1855 (N_1855,N_1584,N_1423);
nor U1856 (N_1856,In_314,N_1610);
nand U1857 (N_1857,N_1725,N_1675);
xor U1858 (N_1858,N_1611,In_1732);
and U1859 (N_1859,N_1008,In_1639);
nand U1860 (N_1860,N_940,N_1153);
nand U1861 (N_1861,N_1713,N_1721);
or U1862 (N_1862,N_1738,N_1711);
nor U1863 (N_1863,N_1373,N_1728);
xnor U1864 (N_1864,N_1591,In_1947);
xor U1865 (N_1865,N_1655,In_1035);
nand U1866 (N_1866,N_119,In_1221);
nor U1867 (N_1867,N_1284,N_1430);
xnor U1868 (N_1868,N_1522,N_1576);
nand U1869 (N_1869,In_1112,N_772);
and U1870 (N_1870,N_1637,In_1551);
or U1871 (N_1871,N_1267,N_1425);
nand U1872 (N_1872,N_1056,N_1345);
and U1873 (N_1873,N_1328,N_873);
and U1874 (N_1874,N_1488,In_217);
or U1875 (N_1875,N_233,N_338);
and U1876 (N_1876,N_1617,N_1690);
and U1877 (N_1877,N_1631,N_1207);
and U1878 (N_1878,In_1887,N_1268);
and U1879 (N_1879,N_1653,N_1623);
nor U1880 (N_1880,N_1662,N_1378);
or U1881 (N_1881,N_52,N_1694);
or U1882 (N_1882,N_1699,In_1004);
nand U1883 (N_1883,N_1188,N_696);
and U1884 (N_1884,N_1557,N_1589);
nor U1885 (N_1885,N_1528,N_1340);
nand U1886 (N_1886,N_782,N_1669);
nand U1887 (N_1887,N_1253,N_1645);
nand U1888 (N_1888,N_911,N_1658);
xor U1889 (N_1889,N_1668,N_550);
and U1890 (N_1890,N_755,In_383);
xor U1891 (N_1891,N_861,N_1706);
xnor U1892 (N_1892,N_1117,N_422);
and U1893 (N_1893,In_2319,N_1402);
xnor U1894 (N_1894,N_875,N_1263);
or U1895 (N_1895,In_1893,N_43);
nor U1896 (N_1896,In_2015,N_1698);
or U1897 (N_1897,N_1597,N_1633);
nand U1898 (N_1898,N_1680,N_648);
nand U1899 (N_1899,N_1506,N_1746);
or U1900 (N_1900,N_382,In_359);
xnor U1901 (N_1901,N_1716,In_426);
or U1902 (N_1902,N_1114,N_939);
or U1903 (N_1903,N_1120,N_1602);
nand U1904 (N_1904,N_1619,In_1585);
xnor U1905 (N_1905,N_1544,In_1003);
or U1906 (N_1906,N_1139,N_1689);
or U1907 (N_1907,N_1643,N_1444);
nor U1908 (N_1908,N_1318,N_175);
and U1909 (N_1909,N_1062,N_1590);
nand U1910 (N_1910,In_661,In_1334);
xnor U1911 (N_1911,N_1517,N_1441);
or U1912 (N_1912,N_952,In_927);
nor U1913 (N_1913,N_1033,N_1595);
and U1914 (N_1914,N_1174,N_1749);
nor U1915 (N_1915,N_1621,N_1638);
nand U1916 (N_1916,N_1098,N_1389);
xnor U1917 (N_1917,N_1384,N_950);
nor U1918 (N_1918,N_1681,N_1622);
nand U1919 (N_1919,N_1671,N_1368);
or U1920 (N_1920,N_1570,N_1412);
nand U1921 (N_1921,In_2387,N_1354);
nor U1922 (N_1922,N_1654,In_1190);
or U1923 (N_1923,In_571,N_622);
or U1924 (N_1924,N_1311,In_466);
or U1925 (N_1925,N_1729,N_864);
nor U1926 (N_1926,In_165,In_591);
nand U1927 (N_1927,N_1501,In_59);
or U1928 (N_1928,N_58,N_1369);
or U1929 (N_1929,N_1178,In_1717);
nor U1930 (N_1930,In_1869,N_494);
nand U1931 (N_1931,N_866,N_393);
nand U1932 (N_1932,N_1169,N_1628);
or U1933 (N_1933,N_1142,In_2459);
and U1934 (N_1934,In_1643,N_1481);
or U1935 (N_1935,N_1647,N_727);
or U1936 (N_1936,In_308,N_1413);
and U1937 (N_1937,N_627,N_1652);
nand U1938 (N_1938,N_252,N_959);
nand U1939 (N_1939,N_957,N_820);
nand U1940 (N_1940,N_1112,In_966);
nor U1941 (N_1941,In_1603,N_1168);
nand U1942 (N_1942,In_1017,N_1556);
nand U1943 (N_1943,N_1395,In_1178);
nand U1944 (N_1944,N_1164,N_1355);
xor U1945 (N_1945,N_1720,N_1531);
xnor U1946 (N_1946,N_1553,N_1308);
nand U1947 (N_1947,N_1316,N_1640);
xor U1948 (N_1948,N_887,N_1583);
xor U1949 (N_1949,N_1559,In_1759);
or U1950 (N_1950,In_604,In_1939);
nand U1951 (N_1951,N_1674,N_1539);
nand U1952 (N_1952,N_1521,N_1550);
or U1953 (N_1953,N_1144,N_1443);
and U1954 (N_1954,N_594,N_1442);
xnor U1955 (N_1955,In_2232,N_1439);
xor U1956 (N_1956,In_2128,N_1003);
or U1957 (N_1957,N_1341,N_1600);
xnor U1958 (N_1958,N_1483,N_1575);
nor U1959 (N_1959,In_329,N_1250);
or U1960 (N_1960,N_1387,In_796);
xor U1961 (N_1961,N_1132,N_678);
nor U1962 (N_1962,In_825,N_1450);
xnor U1963 (N_1963,N_1672,In_652);
and U1964 (N_1964,N_1154,N_1274);
xor U1965 (N_1965,N_1203,In_370);
or U1966 (N_1966,N_1648,N_1649);
nor U1967 (N_1967,N_1541,N_1667);
nor U1968 (N_1968,N_236,N_1518);
xnor U1969 (N_1969,N_1722,N_1399);
nor U1970 (N_1970,N_1515,N_815);
nand U1971 (N_1971,N_417,N_1513);
nor U1972 (N_1972,N_1081,N_1708);
nor U1973 (N_1973,N_582,N_1603);
nand U1974 (N_1974,In_1899,In_529);
or U1975 (N_1975,In_2290,N_1692);
or U1976 (N_1976,N_1574,In_1243);
nor U1977 (N_1977,N_1688,N_412);
nor U1978 (N_1978,In_1097,N_443);
and U1979 (N_1979,N_1571,In_1755);
nor U1980 (N_1980,N_1568,In_1189);
xor U1981 (N_1981,N_1608,N_1348);
or U1982 (N_1982,N_812,N_669);
or U1983 (N_1983,N_322,N_265);
nor U1984 (N_1984,In_1163,N_225);
or U1985 (N_1985,N_1695,N_1731);
nand U1986 (N_1986,N_540,In_1108);
or U1987 (N_1987,N_1078,N_1499);
nor U1988 (N_1988,In_224,N_1418);
and U1989 (N_1989,N_601,In_487);
or U1990 (N_1990,N_1523,In_1249);
and U1991 (N_1991,N_1466,N_1545);
and U1992 (N_1992,In_2312,N_1408);
nor U1993 (N_1993,N_1145,In_771);
nand U1994 (N_1994,In_2233,N_877);
nand U1995 (N_1995,N_1745,N_1514);
nor U1996 (N_1996,In_1129,N_639);
xnor U1997 (N_1997,N_1280,N_1704);
nor U1998 (N_1998,In_337,N_1678);
and U1999 (N_1999,N_784,N_673);
nand U2000 (N_2000,N_1393,N_1701);
xor U2001 (N_2001,N_1951,N_1612);
or U2002 (N_2002,N_1116,In_502);
or U2003 (N_2003,N_698,N_1790);
nor U2004 (N_2004,In_1972,In_269);
nor U2005 (N_2005,N_1979,N_1851);
xor U2006 (N_2006,N_1256,N_369);
xnor U2007 (N_2007,N_730,N_1718);
nand U2008 (N_2008,N_1259,N_1750);
xor U2009 (N_2009,N_1963,In_1624);
nor U2010 (N_2010,N_1726,N_1764);
nand U2011 (N_2011,N_1567,N_1774);
nand U2012 (N_2012,N_1332,N_1981);
nand U2013 (N_2013,In_1020,N_1793);
and U2014 (N_2014,N_1604,N_1770);
xnor U2015 (N_2015,N_765,N_1855);
or U2016 (N_2016,N_1313,N_1596);
xor U2017 (N_2017,N_1456,N_1900);
and U2018 (N_2018,N_1552,In_964);
or U2019 (N_2019,N_1468,N_1944);
or U2020 (N_2020,N_1791,N_1630);
xor U2021 (N_2021,N_1928,N_1709);
or U2022 (N_2022,N_253,N_1277);
or U2023 (N_2023,N_1919,N_1898);
or U2024 (N_2024,N_1788,N_1795);
nor U2025 (N_2025,N_1767,N_1593);
nor U2026 (N_2026,N_1842,N_1357);
nor U2027 (N_2027,N_471,N_1371);
and U2028 (N_2028,N_1743,N_1835);
nor U2029 (N_2029,N_1696,In_1518);
or U2030 (N_2030,N_1930,N_1852);
nor U2031 (N_2031,In_2292,N_1830);
nor U2032 (N_2032,N_1969,N_1753);
nand U2033 (N_2033,N_1973,N_1932);
xor U2034 (N_2034,N_1839,N_919);
nor U2035 (N_2035,N_1936,In_2485);
xor U2036 (N_2036,N_1999,N_1592);
or U2037 (N_2037,N_1769,N_166);
xor U2038 (N_2038,N_1854,N_1922);
and U2039 (N_2039,N_1841,N_1967);
or U2040 (N_2040,N_1042,N_526);
and U2041 (N_2041,N_1891,N_1893);
nor U2042 (N_2042,N_1049,N_1934);
xor U2043 (N_2043,N_1798,N_1011);
or U2044 (N_2044,N_1434,N_1025);
xor U2045 (N_2045,In_896,N_1079);
xor U2046 (N_2046,N_1401,N_1330);
nor U2047 (N_2047,N_1938,N_1914);
and U2048 (N_2048,In_319,N_1751);
and U2049 (N_2049,N_1915,N_1831);
nor U2050 (N_2050,N_1756,N_1864);
nand U2051 (N_2051,N_1380,N_1403);
xnor U2052 (N_2052,N_1878,N_1644);
nand U2053 (N_2053,N_1417,N_1664);
nand U2054 (N_2054,N_1739,N_1799);
nand U2055 (N_2055,In_1084,N_1529);
xor U2056 (N_2056,N_1475,N_1312);
nand U2057 (N_2057,In_1609,N_1843);
and U2058 (N_2058,N_1760,N_1984);
or U2059 (N_2059,N_992,N_1912);
and U2060 (N_2060,N_1714,N_1618);
nand U2061 (N_2061,N_1772,N_1031);
nor U2062 (N_2062,N_1931,N_1943);
and U2063 (N_2063,N_1386,N_1890);
or U2064 (N_2064,N_1065,N_1146);
nor U2065 (N_2065,N_1446,In_2044);
or U2066 (N_2066,N_1727,N_1650);
and U2067 (N_2067,N_1820,N_1287);
xor U2068 (N_2068,N_1026,N_999);
or U2069 (N_2069,N_1454,N_1564);
nor U2070 (N_2070,N_909,N_1555);
nand U2071 (N_2071,N_1800,N_1869);
and U2072 (N_2072,N_1862,N_1787);
and U2073 (N_2073,N_1607,N_1858);
nand U2074 (N_2074,In_325,N_1172);
xor U2075 (N_2075,N_50,N_1474);
and U2076 (N_2076,N_1780,N_1982);
nand U2077 (N_2077,N_1974,N_1246);
or U2078 (N_2078,In_1625,N_570);
and U2079 (N_2079,N_1786,N_1847);
or U2080 (N_2080,N_1865,N_173);
and U2081 (N_2081,N_1525,N_1453);
and U2082 (N_2082,N_1956,In_2056);
nand U2083 (N_2083,N_1775,N_1926);
nand U2084 (N_2084,In_1847,N_1777);
xor U2085 (N_2085,N_1299,N_1971);
and U2086 (N_2086,N_1902,N_1762);
or U2087 (N_2087,N_1832,N_1005);
or U2088 (N_2088,N_834,N_209);
or U2089 (N_2089,In_1175,N_1757);
nor U2090 (N_2090,N_1837,N_1966);
and U2091 (N_2091,N_1916,N_1868);
and U2092 (N_2092,N_1500,N_1904);
xnor U2093 (N_2093,In_100,N_1994);
nor U2094 (N_2094,N_1230,N_1283);
nand U2095 (N_2095,N_1935,N_1017);
nor U2096 (N_2096,N_1889,N_1807);
xnor U2097 (N_2097,N_1846,N_1748);
nor U2098 (N_2098,N_1759,N_1573);
and U2099 (N_2099,N_1988,N_1661);
and U2100 (N_2100,N_1987,N_1899);
xnor U2101 (N_2101,N_1870,N_1765);
nand U2102 (N_2102,N_1954,N_1792);
xor U2103 (N_2103,N_1905,N_1431);
nor U2104 (N_2104,N_1998,N_1819);
or U2105 (N_2105,N_1700,N_1684);
nor U2106 (N_2106,N_1561,N_1975);
xor U2107 (N_2107,N_1520,N_1833);
and U2108 (N_2108,N_1925,N_1803);
and U2109 (N_2109,N_1964,N_1921);
nand U2110 (N_2110,N_927,N_1826);
or U2111 (N_2111,In_643,N_1989);
nand U2112 (N_2112,N_1886,N_1463);
nor U2113 (N_2113,N_1913,N_1258);
or U2114 (N_2114,N_1783,N_942);
and U2115 (N_2115,N_1953,N_1952);
and U2116 (N_2116,N_953,N_1882);
or U2117 (N_2117,N_455,N_1796);
nor U2118 (N_2118,N_1785,N_1942);
nand U2119 (N_2119,N_1372,N_1863);
nor U2120 (N_2120,N_1901,N_1840);
and U2121 (N_2121,N_1771,N_1888);
nand U2122 (N_2122,N_1781,N_1616);
and U2123 (N_2123,N_1587,In_2162);
nand U2124 (N_2124,N_1908,N_1879);
nor U2125 (N_2125,N_1949,In_838);
and U2126 (N_2126,N_1755,N_1829);
nor U2127 (N_2127,N_1779,N_1945);
and U2128 (N_2128,N_1358,N_1502);
or U2129 (N_2129,N_1693,N_1181);
or U2130 (N_2130,N_1761,N_1923);
and U2131 (N_2131,N_1993,In_2138);
or U2132 (N_2132,In_1999,N_1560);
nand U2133 (N_2133,N_1057,N_1825);
and U2134 (N_2134,N_1730,N_1736);
and U2135 (N_2135,N_1289,N_420);
and U2136 (N_2136,N_862,N_1542);
nand U2137 (N_2137,N_1381,N_1968);
xnor U2138 (N_2138,N_1615,N_1804);
xor U2139 (N_2139,N_1903,In_2114);
and U2140 (N_2140,In_381,N_1814);
or U2141 (N_2141,N_1794,N_1857);
or U2142 (N_2142,N_1763,In_1495);
nand U2143 (N_2143,N_1887,N_1929);
xor U2144 (N_2144,N_1536,In_1506);
xnor U2145 (N_2145,N_1766,In_1496);
nand U2146 (N_2146,N_1606,N_1872);
nand U2147 (N_2147,N_3,N_1797);
and U2148 (N_2148,N_1961,In_1809);
nor U2149 (N_2149,N_1828,N_1015);
xnor U2150 (N_2150,N_1896,N_1970);
xnor U2151 (N_2151,N_1946,N_1990);
xnor U2152 (N_2152,N_1566,N_1554);
nand U2153 (N_2153,N_1758,N_802);
and U2154 (N_2154,N_467,N_1906);
or U2155 (N_2155,N_1064,N_1850);
nand U2156 (N_2156,N_1883,N_1808);
and U2157 (N_2157,N_1512,N_632);
xor U2158 (N_2158,N_1867,N_1958);
nand U2159 (N_2159,N_1844,N_1382);
or U2160 (N_2160,N_1941,N_1897);
nand U2161 (N_2161,N_1991,N_1625);
nor U2162 (N_2162,In_2111,N_1180);
xor U2163 (N_2163,N_1866,N_1810);
or U2164 (N_2164,N_1754,N_1183);
and U2165 (N_2165,In_1303,N_1367);
xor U2166 (N_2166,N_1656,N_1101);
nand U2167 (N_2167,N_1115,N_1641);
xnor U2168 (N_2168,N_1773,N_1873);
nor U2169 (N_2169,In_1924,N_1626);
or U2170 (N_2170,N_569,N_827);
nor U2171 (N_2171,N_1895,N_1588);
and U2172 (N_2172,N_1538,N_1909);
nand U2173 (N_2173,N_1976,N_1924);
nand U2174 (N_2174,N_1874,N_1257);
or U2175 (N_2175,N_1983,In_557);
xnor U2176 (N_2176,N_1995,N_1860);
xnor U2177 (N_2177,N_1816,In_313);
or U2178 (N_2178,N_1577,N_1424);
or U2179 (N_2179,N_1163,N_1940);
or U2180 (N_2180,N_1673,N_1282);
xnor U2181 (N_2181,N_490,N_1950);
xor U2182 (N_2182,N_1639,N_1447);
or U2183 (N_2183,N_1620,In_1491);
nand U2184 (N_2184,N_1823,N_1789);
or U2185 (N_2185,N_1204,N_674);
xor U2186 (N_2186,N_1460,N_1752);
or U2187 (N_2187,N_1996,N_1734);
or U2188 (N_2188,N_1776,N_1965);
xnor U2189 (N_2189,N_1676,N_1811);
xnor U2190 (N_2190,In_2347,N_1955);
nor U2191 (N_2191,N_1892,N_1962);
xnor U2192 (N_2192,N_1907,N_1849);
xnor U2193 (N_2193,N_1937,In_2192);
nand U2194 (N_2194,N_1805,N_1972);
or U2195 (N_2195,N_1784,N_1861);
nand U2196 (N_2196,N_1806,N_792);
xnor U2197 (N_2197,N_1212,N_1778);
xor U2198 (N_2198,N_1598,N_618);
and U2199 (N_2199,N_1768,N_1659);
or U2200 (N_2200,N_442,N_773);
nor U2201 (N_2201,N_1272,N_852);
nor U2202 (N_2202,N_1679,N_1352);
or U2203 (N_2203,N_1917,N_1848);
nor U2204 (N_2204,N_1534,N_1910);
and U2205 (N_2205,N_1377,N_1642);
nor U2206 (N_2206,N_1845,N_1321);
xnor U2207 (N_2207,N_195,N_1918);
and U2208 (N_2208,N_1809,N_1997);
nand U2209 (N_2209,N_1817,N_449);
or U2210 (N_2210,N_1859,N_1960);
and U2211 (N_2211,N_1744,In_1135);
and U2212 (N_2212,N_1363,N_1877);
and U2213 (N_2213,N_1920,N_1601);
nor U2214 (N_2214,In_2283,In_1970);
and U2215 (N_2215,N_1646,N_1325);
nor U2216 (N_2216,N_1836,N_1894);
nand U2217 (N_2217,N_1459,N_1980);
and U2218 (N_2218,N_1871,N_1801);
and U2219 (N_2219,N_1812,In_1814);
or U2220 (N_2220,N_1838,N_1366);
or U2221 (N_2221,N_1876,N_1827);
and U2222 (N_2222,N_1948,N_1578);
xnor U2223 (N_2223,N_1992,N_1802);
nand U2224 (N_2224,N_1303,N_255);
and U2225 (N_2225,N_1875,N_1821);
and U2226 (N_2226,N_1933,N_1939);
or U2227 (N_2227,N_1884,In_1196);
xor U2228 (N_2228,N_1815,N_1527);
xnor U2229 (N_2229,N_1581,N_1985);
or U2230 (N_2230,N_1045,N_1391);
nand U2231 (N_2231,N_1505,N_1663);
and U2232 (N_2232,N_1682,In_2436);
nor U2233 (N_2233,In_87,N_1187);
or U2234 (N_2234,N_1927,N_1959);
or U2235 (N_2235,N_1957,In_909);
or U2236 (N_2236,N_1822,N_1856);
xnor U2237 (N_2237,N_1478,N_1911);
nor U2238 (N_2238,In_1896,N_1880);
or U2239 (N_2239,N_1986,N_1509);
nand U2240 (N_2240,N_1782,N_1565);
or U2241 (N_2241,N_1885,N_1834);
xor U2242 (N_2242,In_564,N_1818);
and U2243 (N_2243,N_1265,N_1813);
nand U2244 (N_2244,N_1853,N_721);
nor U2245 (N_2245,In_853,N_1947);
and U2246 (N_2246,N_1579,N_1978);
nand U2247 (N_2247,N_1977,N_1733);
or U2248 (N_2248,N_1260,In_1848);
nand U2249 (N_2249,N_1824,N_1881);
or U2250 (N_2250,N_2205,N_2219);
xor U2251 (N_2251,N_2193,N_2047);
nand U2252 (N_2252,N_2177,N_2033);
nand U2253 (N_2253,N_2059,N_2171);
xnor U2254 (N_2254,N_2133,N_2196);
nand U2255 (N_2255,N_2165,N_2118);
and U2256 (N_2256,N_2107,N_2216);
nor U2257 (N_2257,N_2231,N_2218);
and U2258 (N_2258,N_2140,N_2122);
xor U2259 (N_2259,N_2138,N_2108);
nor U2260 (N_2260,N_2224,N_2173);
nand U2261 (N_2261,N_2227,N_2199);
nand U2262 (N_2262,N_2155,N_2065);
and U2263 (N_2263,N_2030,N_2192);
xnor U2264 (N_2264,N_2167,N_2111);
nor U2265 (N_2265,N_2249,N_2142);
or U2266 (N_2266,N_2197,N_2166);
xnor U2267 (N_2267,N_2057,N_2044);
and U2268 (N_2268,N_2037,N_2087);
xnor U2269 (N_2269,N_2116,N_2055);
or U2270 (N_2270,N_2103,N_2201);
xor U2271 (N_2271,N_2072,N_2094);
or U2272 (N_2272,N_2035,N_2176);
and U2273 (N_2273,N_2150,N_2169);
xor U2274 (N_2274,N_2245,N_2164);
and U2275 (N_2275,N_2183,N_2151);
nand U2276 (N_2276,N_2112,N_2115);
nor U2277 (N_2277,N_2212,N_2110);
nor U2278 (N_2278,N_2002,N_2010);
and U2279 (N_2279,N_2052,N_2060);
xnor U2280 (N_2280,N_2195,N_2147);
xor U2281 (N_2281,N_2001,N_2004);
nand U2282 (N_2282,N_2029,N_2109);
nor U2283 (N_2283,N_2117,N_2238);
nand U2284 (N_2284,N_2056,N_2102);
and U2285 (N_2285,N_2200,N_2185);
and U2286 (N_2286,N_2003,N_2043);
nor U2287 (N_2287,N_2092,N_2069);
and U2288 (N_2288,N_2208,N_2038);
nand U2289 (N_2289,N_2246,N_2143);
nor U2290 (N_2290,N_2214,N_2141);
and U2291 (N_2291,N_2063,N_2130);
nand U2292 (N_2292,N_2040,N_2244);
nand U2293 (N_2293,N_2194,N_2210);
xor U2294 (N_2294,N_2049,N_2139);
xnor U2295 (N_2295,N_2021,N_2084);
nand U2296 (N_2296,N_2067,N_2154);
and U2297 (N_2297,N_2051,N_2162);
or U2298 (N_2298,N_2163,N_2221);
nor U2299 (N_2299,N_2024,N_2160);
or U2300 (N_2300,N_2120,N_2175);
nand U2301 (N_2301,N_2093,N_2054);
xnor U2302 (N_2302,N_2188,N_2020);
nand U2303 (N_2303,N_2158,N_2011);
or U2304 (N_2304,N_2028,N_2036);
or U2305 (N_2305,N_2000,N_2228);
and U2306 (N_2306,N_2085,N_2106);
and U2307 (N_2307,N_2039,N_2025);
or U2308 (N_2308,N_2125,N_2089);
and U2309 (N_2309,N_2204,N_2009);
and U2310 (N_2310,N_2136,N_2068);
or U2311 (N_2311,N_2174,N_2235);
xor U2312 (N_2312,N_2058,N_2070);
nor U2313 (N_2313,N_2086,N_2189);
or U2314 (N_2314,N_2064,N_2017);
or U2315 (N_2315,N_2157,N_2159);
nor U2316 (N_2316,N_2191,N_2023);
and U2317 (N_2317,N_2016,N_2124);
nor U2318 (N_2318,N_2222,N_2091);
nand U2319 (N_2319,N_2234,N_2226);
nand U2320 (N_2320,N_2248,N_2146);
and U2321 (N_2321,N_2145,N_2180);
and U2322 (N_2322,N_2129,N_2123);
or U2323 (N_2323,N_2223,N_2076);
xnor U2324 (N_2324,N_2104,N_2137);
nand U2325 (N_2325,N_2131,N_2209);
nor U2326 (N_2326,N_2041,N_2190);
and U2327 (N_2327,N_2127,N_2097);
xnor U2328 (N_2328,N_2083,N_2132);
nand U2329 (N_2329,N_2178,N_2082);
and U2330 (N_2330,N_2042,N_2031);
or U2331 (N_2331,N_2046,N_2012);
nand U2332 (N_2332,N_2217,N_2186);
xnor U2333 (N_2333,N_2095,N_2101);
and U2334 (N_2334,N_2061,N_2081);
nand U2335 (N_2335,N_2078,N_2013);
nor U2336 (N_2336,N_2242,N_2098);
nand U2337 (N_2337,N_2247,N_2005);
nand U2338 (N_2338,N_2113,N_2229);
and U2339 (N_2339,N_2207,N_2014);
and U2340 (N_2340,N_2080,N_2032);
xor U2341 (N_2341,N_2187,N_2114);
xor U2342 (N_2342,N_2119,N_2230);
xnor U2343 (N_2343,N_2156,N_2053);
or U2344 (N_2344,N_2240,N_2045);
nor U2345 (N_2345,N_2148,N_2026);
nand U2346 (N_2346,N_2050,N_2203);
and U2347 (N_2347,N_2168,N_2179);
and U2348 (N_2348,N_2126,N_2019);
and U2349 (N_2349,N_2048,N_2077);
xnor U2350 (N_2350,N_2233,N_2096);
or U2351 (N_2351,N_2088,N_2007);
xor U2352 (N_2352,N_2034,N_2066);
and U2353 (N_2353,N_2022,N_2018);
and U2354 (N_2354,N_2121,N_2071);
xnor U2355 (N_2355,N_2079,N_2153);
nand U2356 (N_2356,N_2170,N_2239);
nor U2357 (N_2357,N_2008,N_2202);
or U2358 (N_2358,N_2090,N_2006);
nand U2359 (N_2359,N_2198,N_2135);
and U2360 (N_2360,N_2236,N_2149);
or U2361 (N_2361,N_2237,N_2215);
xnor U2362 (N_2362,N_2225,N_2100);
or U2363 (N_2363,N_2220,N_2182);
nor U2364 (N_2364,N_2241,N_2099);
xor U2365 (N_2365,N_2206,N_2074);
nand U2366 (N_2366,N_2232,N_2015);
and U2367 (N_2367,N_2211,N_2105);
or U2368 (N_2368,N_2172,N_2134);
nor U2369 (N_2369,N_2027,N_2075);
and U2370 (N_2370,N_2152,N_2243);
and U2371 (N_2371,N_2062,N_2144);
nand U2372 (N_2372,N_2073,N_2213);
nor U2373 (N_2373,N_2161,N_2184);
nor U2374 (N_2374,N_2128,N_2181);
and U2375 (N_2375,N_2148,N_2176);
and U2376 (N_2376,N_2225,N_2134);
xnor U2377 (N_2377,N_2059,N_2101);
xnor U2378 (N_2378,N_2132,N_2031);
xnor U2379 (N_2379,N_2021,N_2067);
nor U2380 (N_2380,N_2157,N_2021);
or U2381 (N_2381,N_2206,N_2248);
xor U2382 (N_2382,N_2090,N_2059);
nor U2383 (N_2383,N_2135,N_2019);
xnor U2384 (N_2384,N_2217,N_2042);
nor U2385 (N_2385,N_2220,N_2053);
xnor U2386 (N_2386,N_2233,N_2058);
or U2387 (N_2387,N_2207,N_2029);
nor U2388 (N_2388,N_2069,N_2114);
nand U2389 (N_2389,N_2084,N_2236);
and U2390 (N_2390,N_2234,N_2070);
or U2391 (N_2391,N_2226,N_2027);
and U2392 (N_2392,N_2140,N_2155);
and U2393 (N_2393,N_2174,N_2110);
nand U2394 (N_2394,N_2030,N_2040);
or U2395 (N_2395,N_2037,N_2000);
or U2396 (N_2396,N_2047,N_2233);
and U2397 (N_2397,N_2205,N_2216);
or U2398 (N_2398,N_2100,N_2088);
and U2399 (N_2399,N_2118,N_2031);
or U2400 (N_2400,N_2132,N_2130);
xnor U2401 (N_2401,N_2109,N_2015);
nor U2402 (N_2402,N_2058,N_2205);
xor U2403 (N_2403,N_2148,N_2076);
and U2404 (N_2404,N_2104,N_2114);
xor U2405 (N_2405,N_2095,N_2074);
xnor U2406 (N_2406,N_2208,N_2194);
nor U2407 (N_2407,N_2192,N_2110);
xnor U2408 (N_2408,N_2214,N_2145);
nand U2409 (N_2409,N_2021,N_2020);
xnor U2410 (N_2410,N_2134,N_2074);
nand U2411 (N_2411,N_2057,N_2007);
nor U2412 (N_2412,N_2120,N_2102);
nor U2413 (N_2413,N_2068,N_2160);
xnor U2414 (N_2414,N_2112,N_2200);
nand U2415 (N_2415,N_2071,N_2062);
xor U2416 (N_2416,N_2125,N_2168);
nand U2417 (N_2417,N_2235,N_2180);
and U2418 (N_2418,N_2041,N_2098);
or U2419 (N_2419,N_2051,N_2194);
nor U2420 (N_2420,N_2246,N_2211);
xor U2421 (N_2421,N_2092,N_2204);
nand U2422 (N_2422,N_2004,N_2049);
xor U2423 (N_2423,N_2060,N_2119);
xor U2424 (N_2424,N_2200,N_2106);
nor U2425 (N_2425,N_2200,N_2116);
nand U2426 (N_2426,N_2059,N_2098);
nand U2427 (N_2427,N_2166,N_2000);
nand U2428 (N_2428,N_2195,N_2228);
and U2429 (N_2429,N_2187,N_2141);
nor U2430 (N_2430,N_2025,N_2129);
or U2431 (N_2431,N_2136,N_2045);
and U2432 (N_2432,N_2094,N_2108);
xor U2433 (N_2433,N_2007,N_2034);
nor U2434 (N_2434,N_2143,N_2102);
nand U2435 (N_2435,N_2195,N_2238);
nand U2436 (N_2436,N_2077,N_2014);
xor U2437 (N_2437,N_2154,N_2137);
and U2438 (N_2438,N_2007,N_2216);
nor U2439 (N_2439,N_2053,N_2180);
nand U2440 (N_2440,N_2140,N_2171);
nor U2441 (N_2441,N_2099,N_2060);
xor U2442 (N_2442,N_2147,N_2172);
or U2443 (N_2443,N_2247,N_2060);
and U2444 (N_2444,N_2045,N_2229);
and U2445 (N_2445,N_2106,N_2160);
or U2446 (N_2446,N_2136,N_2241);
xor U2447 (N_2447,N_2032,N_2079);
or U2448 (N_2448,N_2181,N_2230);
and U2449 (N_2449,N_2170,N_2191);
and U2450 (N_2450,N_2215,N_2236);
nor U2451 (N_2451,N_2170,N_2156);
and U2452 (N_2452,N_2173,N_2101);
or U2453 (N_2453,N_2158,N_2031);
or U2454 (N_2454,N_2203,N_2104);
and U2455 (N_2455,N_2020,N_2192);
xor U2456 (N_2456,N_2211,N_2232);
nor U2457 (N_2457,N_2161,N_2104);
and U2458 (N_2458,N_2113,N_2221);
and U2459 (N_2459,N_2129,N_2153);
xor U2460 (N_2460,N_2104,N_2215);
nor U2461 (N_2461,N_2134,N_2037);
or U2462 (N_2462,N_2037,N_2135);
nand U2463 (N_2463,N_2033,N_2231);
or U2464 (N_2464,N_2154,N_2212);
xor U2465 (N_2465,N_2043,N_2077);
nand U2466 (N_2466,N_2032,N_2100);
or U2467 (N_2467,N_2230,N_2064);
nand U2468 (N_2468,N_2091,N_2057);
xor U2469 (N_2469,N_2014,N_2244);
or U2470 (N_2470,N_2194,N_2205);
xnor U2471 (N_2471,N_2139,N_2009);
nand U2472 (N_2472,N_2120,N_2217);
xor U2473 (N_2473,N_2176,N_2212);
or U2474 (N_2474,N_2109,N_2085);
nand U2475 (N_2475,N_2031,N_2046);
nor U2476 (N_2476,N_2143,N_2022);
or U2477 (N_2477,N_2005,N_2157);
or U2478 (N_2478,N_2039,N_2159);
xnor U2479 (N_2479,N_2136,N_2249);
nor U2480 (N_2480,N_2040,N_2032);
xor U2481 (N_2481,N_2123,N_2167);
or U2482 (N_2482,N_2137,N_2162);
xnor U2483 (N_2483,N_2100,N_2019);
and U2484 (N_2484,N_2221,N_2038);
and U2485 (N_2485,N_2095,N_2206);
nand U2486 (N_2486,N_2224,N_2244);
and U2487 (N_2487,N_2185,N_2191);
or U2488 (N_2488,N_2231,N_2119);
or U2489 (N_2489,N_2111,N_2163);
nor U2490 (N_2490,N_2156,N_2228);
nand U2491 (N_2491,N_2143,N_2133);
or U2492 (N_2492,N_2193,N_2036);
and U2493 (N_2493,N_2001,N_2020);
xnor U2494 (N_2494,N_2049,N_2050);
nor U2495 (N_2495,N_2179,N_2232);
nand U2496 (N_2496,N_2111,N_2065);
and U2497 (N_2497,N_2094,N_2128);
or U2498 (N_2498,N_2181,N_2074);
nand U2499 (N_2499,N_2011,N_2185);
xor U2500 (N_2500,N_2378,N_2301);
nor U2501 (N_2501,N_2264,N_2275);
nand U2502 (N_2502,N_2306,N_2458);
nor U2503 (N_2503,N_2416,N_2476);
xor U2504 (N_2504,N_2493,N_2252);
nand U2505 (N_2505,N_2345,N_2388);
nand U2506 (N_2506,N_2364,N_2270);
nand U2507 (N_2507,N_2420,N_2479);
xnor U2508 (N_2508,N_2439,N_2438);
nor U2509 (N_2509,N_2347,N_2279);
and U2510 (N_2510,N_2392,N_2253);
and U2511 (N_2511,N_2498,N_2339);
xor U2512 (N_2512,N_2332,N_2318);
xnor U2513 (N_2513,N_2419,N_2446);
or U2514 (N_2514,N_2311,N_2471);
nand U2515 (N_2515,N_2467,N_2254);
nand U2516 (N_2516,N_2278,N_2309);
or U2517 (N_2517,N_2369,N_2346);
and U2518 (N_2518,N_2292,N_2331);
or U2519 (N_2519,N_2360,N_2308);
and U2520 (N_2520,N_2461,N_2468);
nor U2521 (N_2521,N_2299,N_2336);
and U2522 (N_2522,N_2302,N_2286);
xnor U2523 (N_2523,N_2442,N_2291);
and U2524 (N_2524,N_2402,N_2435);
xor U2525 (N_2525,N_2454,N_2460);
and U2526 (N_2526,N_2405,N_2449);
nand U2527 (N_2527,N_2317,N_2492);
nand U2528 (N_2528,N_2355,N_2422);
and U2529 (N_2529,N_2394,N_2362);
nor U2530 (N_2530,N_2404,N_2289);
and U2531 (N_2531,N_2497,N_2398);
nor U2532 (N_2532,N_2379,N_2418);
nand U2533 (N_2533,N_2256,N_2396);
and U2534 (N_2534,N_2353,N_2282);
xnor U2535 (N_2535,N_2411,N_2348);
nand U2536 (N_2536,N_2349,N_2257);
nand U2537 (N_2537,N_2481,N_2295);
nor U2538 (N_2538,N_2459,N_2401);
xnor U2539 (N_2539,N_2304,N_2277);
or U2540 (N_2540,N_2451,N_2274);
or U2541 (N_2541,N_2276,N_2395);
or U2542 (N_2542,N_2478,N_2310);
and U2543 (N_2543,N_2367,N_2477);
nand U2544 (N_2544,N_2259,N_2445);
nor U2545 (N_2545,N_2415,N_2487);
xnor U2546 (N_2546,N_2366,N_2485);
xnor U2547 (N_2547,N_2327,N_2303);
nand U2548 (N_2548,N_2456,N_2316);
or U2549 (N_2549,N_2329,N_2272);
and U2550 (N_2550,N_2465,N_2382);
nand U2551 (N_2551,N_2389,N_2338);
and U2552 (N_2552,N_2473,N_2281);
nor U2553 (N_2553,N_2262,N_2384);
or U2554 (N_2554,N_2255,N_2258);
or U2555 (N_2555,N_2437,N_2436);
and U2556 (N_2556,N_2261,N_2483);
nor U2557 (N_2557,N_2496,N_2328);
and U2558 (N_2558,N_2495,N_2283);
xor U2559 (N_2559,N_2391,N_2410);
xnor U2560 (N_2560,N_2285,N_2490);
and U2561 (N_2561,N_2335,N_2350);
and U2562 (N_2562,N_2361,N_2374);
and U2563 (N_2563,N_2466,N_2406);
or U2564 (N_2564,N_2486,N_2413);
or U2565 (N_2565,N_2408,N_2489);
nand U2566 (N_2566,N_2273,N_2429);
and U2567 (N_2567,N_2323,N_2450);
xor U2568 (N_2568,N_2342,N_2298);
and U2569 (N_2569,N_2284,N_2421);
or U2570 (N_2570,N_2475,N_2368);
nand U2571 (N_2571,N_2463,N_2387);
xor U2572 (N_2572,N_2484,N_2337);
nor U2573 (N_2573,N_2455,N_2397);
xor U2574 (N_2574,N_2354,N_2357);
xnor U2575 (N_2575,N_2326,N_2296);
nand U2576 (N_2576,N_2430,N_2433);
xnor U2577 (N_2577,N_2321,N_2322);
or U2578 (N_2578,N_2359,N_2363);
nor U2579 (N_2579,N_2365,N_2440);
xnor U2580 (N_2580,N_2325,N_2474);
and U2581 (N_2581,N_2417,N_2351);
and U2582 (N_2582,N_2324,N_2453);
xor U2583 (N_2583,N_2305,N_2290);
xnor U2584 (N_2584,N_2432,N_2424);
xor U2585 (N_2585,N_2425,N_2383);
nor U2586 (N_2586,N_2314,N_2315);
or U2587 (N_2587,N_2400,N_2431);
or U2588 (N_2588,N_2293,N_2482);
nor U2589 (N_2589,N_2414,N_2447);
or U2590 (N_2590,N_2263,N_2499);
xnor U2591 (N_2591,N_2470,N_2494);
and U2592 (N_2592,N_2251,N_2268);
nand U2593 (N_2593,N_2333,N_2480);
xor U2594 (N_2594,N_2267,N_2265);
xnor U2595 (N_2595,N_2358,N_2330);
or U2596 (N_2596,N_2297,N_2260);
nor U2597 (N_2597,N_2491,N_2462);
nand U2598 (N_2598,N_2423,N_2386);
nand U2599 (N_2599,N_2287,N_2393);
xnor U2600 (N_2600,N_2266,N_2312);
nor U2601 (N_2601,N_2313,N_2434);
and U2602 (N_2602,N_2426,N_2448);
nand U2603 (N_2603,N_2385,N_2344);
and U2604 (N_2604,N_2372,N_2428);
xnor U2605 (N_2605,N_2376,N_2452);
and U2606 (N_2606,N_2343,N_2469);
nor U2607 (N_2607,N_2250,N_2288);
nor U2608 (N_2608,N_2399,N_2380);
or U2609 (N_2609,N_2427,N_2390);
nand U2610 (N_2610,N_2464,N_2269);
nor U2611 (N_2611,N_2352,N_2356);
nand U2612 (N_2612,N_2381,N_2319);
xor U2613 (N_2613,N_2409,N_2407);
or U2614 (N_2614,N_2488,N_2443);
nand U2615 (N_2615,N_2271,N_2444);
nor U2616 (N_2616,N_2412,N_2307);
and U2617 (N_2617,N_2377,N_2334);
nand U2618 (N_2618,N_2375,N_2371);
or U2619 (N_2619,N_2403,N_2300);
and U2620 (N_2620,N_2441,N_2472);
xnor U2621 (N_2621,N_2280,N_2457);
nand U2622 (N_2622,N_2373,N_2320);
nor U2623 (N_2623,N_2370,N_2294);
nor U2624 (N_2624,N_2341,N_2340);
nand U2625 (N_2625,N_2270,N_2437);
or U2626 (N_2626,N_2498,N_2492);
and U2627 (N_2627,N_2381,N_2331);
or U2628 (N_2628,N_2495,N_2449);
xnor U2629 (N_2629,N_2303,N_2282);
or U2630 (N_2630,N_2338,N_2452);
and U2631 (N_2631,N_2345,N_2374);
or U2632 (N_2632,N_2404,N_2272);
and U2633 (N_2633,N_2379,N_2304);
nand U2634 (N_2634,N_2284,N_2326);
nand U2635 (N_2635,N_2395,N_2365);
or U2636 (N_2636,N_2307,N_2292);
nor U2637 (N_2637,N_2267,N_2479);
nor U2638 (N_2638,N_2479,N_2416);
nand U2639 (N_2639,N_2441,N_2494);
xor U2640 (N_2640,N_2454,N_2287);
nand U2641 (N_2641,N_2352,N_2392);
and U2642 (N_2642,N_2417,N_2409);
or U2643 (N_2643,N_2311,N_2288);
nand U2644 (N_2644,N_2309,N_2440);
or U2645 (N_2645,N_2250,N_2353);
nand U2646 (N_2646,N_2391,N_2319);
nor U2647 (N_2647,N_2427,N_2355);
and U2648 (N_2648,N_2283,N_2266);
and U2649 (N_2649,N_2293,N_2317);
and U2650 (N_2650,N_2324,N_2256);
xor U2651 (N_2651,N_2468,N_2295);
and U2652 (N_2652,N_2327,N_2444);
xor U2653 (N_2653,N_2444,N_2342);
nand U2654 (N_2654,N_2493,N_2445);
or U2655 (N_2655,N_2402,N_2258);
nor U2656 (N_2656,N_2423,N_2315);
xnor U2657 (N_2657,N_2469,N_2455);
xnor U2658 (N_2658,N_2460,N_2453);
xnor U2659 (N_2659,N_2436,N_2343);
nor U2660 (N_2660,N_2448,N_2455);
nand U2661 (N_2661,N_2479,N_2398);
nor U2662 (N_2662,N_2426,N_2256);
xnor U2663 (N_2663,N_2450,N_2456);
xnor U2664 (N_2664,N_2400,N_2311);
nand U2665 (N_2665,N_2415,N_2384);
and U2666 (N_2666,N_2431,N_2309);
or U2667 (N_2667,N_2364,N_2471);
nor U2668 (N_2668,N_2457,N_2399);
and U2669 (N_2669,N_2295,N_2425);
nand U2670 (N_2670,N_2356,N_2456);
nor U2671 (N_2671,N_2250,N_2361);
and U2672 (N_2672,N_2404,N_2277);
nor U2673 (N_2673,N_2289,N_2417);
and U2674 (N_2674,N_2271,N_2472);
or U2675 (N_2675,N_2253,N_2412);
and U2676 (N_2676,N_2299,N_2443);
and U2677 (N_2677,N_2301,N_2413);
or U2678 (N_2678,N_2279,N_2322);
nand U2679 (N_2679,N_2402,N_2280);
nor U2680 (N_2680,N_2457,N_2498);
nand U2681 (N_2681,N_2284,N_2277);
and U2682 (N_2682,N_2419,N_2409);
nor U2683 (N_2683,N_2357,N_2496);
and U2684 (N_2684,N_2387,N_2462);
nor U2685 (N_2685,N_2380,N_2306);
or U2686 (N_2686,N_2334,N_2333);
nand U2687 (N_2687,N_2402,N_2265);
nor U2688 (N_2688,N_2488,N_2461);
or U2689 (N_2689,N_2370,N_2254);
or U2690 (N_2690,N_2479,N_2424);
or U2691 (N_2691,N_2270,N_2295);
or U2692 (N_2692,N_2359,N_2464);
or U2693 (N_2693,N_2303,N_2345);
or U2694 (N_2694,N_2334,N_2482);
and U2695 (N_2695,N_2340,N_2474);
nand U2696 (N_2696,N_2383,N_2334);
xnor U2697 (N_2697,N_2427,N_2295);
xor U2698 (N_2698,N_2339,N_2433);
xnor U2699 (N_2699,N_2456,N_2490);
xnor U2700 (N_2700,N_2376,N_2307);
nor U2701 (N_2701,N_2273,N_2417);
and U2702 (N_2702,N_2426,N_2439);
or U2703 (N_2703,N_2302,N_2292);
and U2704 (N_2704,N_2394,N_2371);
xnor U2705 (N_2705,N_2317,N_2439);
nand U2706 (N_2706,N_2323,N_2405);
nand U2707 (N_2707,N_2293,N_2308);
and U2708 (N_2708,N_2325,N_2460);
and U2709 (N_2709,N_2432,N_2279);
or U2710 (N_2710,N_2438,N_2479);
nand U2711 (N_2711,N_2484,N_2273);
nand U2712 (N_2712,N_2323,N_2319);
nor U2713 (N_2713,N_2467,N_2369);
xnor U2714 (N_2714,N_2448,N_2442);
xor U2715 (N_2715,N_2251,N_2308);
nand U2716 (N_2716,N_2284,N_2283);
nor U2717 (N_2717,N_2402,N_2331);
nor U2718 (N_2718,N_2308,N_2447);
nand U2719 (N_2719,N_2480,N_2445);
xnor U2720 (N_2720,N_2476,N_2481);
xor U2721 (N_2721,N_2480,N_2337);
or U2722 (N_2722,N_2430,N_2313);
or U2723 (N_2723,N_2384,N_2430);
and U2724 (N_2724,N_2460,N_2375);
and U2725 (N_2725,N_2282,N_2267);
and U2726 (N_2726,N_2281,N_2435);
xnor U2727 (N_2727,N_2426,N_2491);
and U2728 (N_2728,N_2381,N_2487);
or U2729 (N_2729,N_2291,N_2270);
xnor U2730 (N_2730,N_2471,N_2282);
or U2731 (N_2731,N_2278,N_2464);
or U2732 (N_2732,N_2380,N_2371);
xor U2733 (N_2733,N_2397,N_2255);
or U2734 (N_2734,N_2455,N_2384);
or U2735 (N_2735,N_2291,N_2472);
nand U2736 (N_2736,N_2341,N_2262);
nor U2737 (N_2737,N_2458,N_2367);
nor U2738 (N_2738,N_2250,N_2357);
nor U2739 (N_2739,N_2305,N_2497);
xnor U2740 (N_2740,N_2370,N_2259);
xnor U2741 (N_2741,N_2457,N_2363);
nor U2742 (N_2742,N_2254,N_2302);
and U2743 (N_2743,N_2472,N_2410);
nand U2744 (N_2744,N_2462,N_2379);
nand U2745 (N_2745,N_2478,N_2343);
or U2746 (N_2746,N_2435,N_2409);
nand U2747 (N_2747,N_2335,N_2357);
and U2748 (N_2748,N_2332,N_2311);
and U2749 (N_2749,N_2293,N_2415);
or U2750 (N_2750,N_2551,N_2730);
and U2751 (N_2751,N_2691,N_2686);
or U2752 (N_2752,N_2571,N_2631);
and U2753 (N_2753,N_2707,N_2549);
xnor U2754 (N_2754,N_2722,N_2633);
nand U2755 (N_2755,N_2718,N_2527);
and U2756 (N_2756,N_2617,N_2674);
nand U2757 (N_2757,N_2590,N_2662);
or U2758 (N_2758,N_2698,N_2605);
nor U2759 (N_2759,N_2550,N_2664);
or U2760 (N_2760,N_2723,N_2608);
nor U2761 (N_2761,N_2545,N_2560);
nor U2762 (N_2762,N_2610,N_2502);
or U2763 (N_2763,N_2602,N_2531);
or U2764 (N_2764,N_2629,N_2692);
or U2765 (N_2765,N_2626,N_2713);
xnor U2766 (N_2766,N_2657,N_2574);
or U2767 (N_2767,N_2620,N_2685);
and U2768 (N_2768,N_2632,N_2697);
nor U2769 (N_2769,N_2640,N_2643);
nor U2770 (N_2770,N_2743,N_2727);
xnor U2771 (N_2771,N_2612,N_2699);
or U2772 (N_2772,N_2503,N_2696);
or U2773 (N_2773,N_2592,N_2706);
or U2774 (N_2774,N_2519,N_2580);
and U2775 (N_2775,N_2599,N_2651);
xnor U2776 (N_2776,N_2573,N_2583);
nor U2777 (N_2777,N_2601,N_2703);
or U2778 (N_2778,N_2719,N_2581);
nand U2779 (N_2779,N_2740,N_2732);
xor U2780 (N_2780,N_2660,N_2704);
and U2781 (N_2781,N_2589,N_2665);
nor U2782 (N_2782,N_2563,N_2734);
and U2783 (N_2783,N_2544,N_2611);
nand U2784 (N_2784,N_2733,N_2509);
and U2785 (N_2785,N_2619,N_2736);
and U2786 (N_2786,N_2600,N_2546);
xnor U2787 (N_2787,N_2711,N_2562);
nand U2788 (N_2788,N_2523,N_2529);
and U2789 (N_2789,N_2705,N_2615);
xor U2790 (N_2790,N_2624,N_2582);
xor U2791 (N_2791,N_2678,N_2726);
and U2792 (N_2792,N_2561,N_2683);
nand U2793 (N_2793,N_2653,N_2625);
xnor U2794 (N_2794,N_2663,N_2712);
and U2795 (N_2795,N_2717,N_2675);
nor U2796 (N_2796,N_2649,N_2558);
nor U2797 (N_2797,N_2721,N_2587);
xnor U2798 (N_2798,N_2634,N_2618);
nand U2799 (N_2799,N_2532,N_2728);
xnor U2800 (N_2800,N_2689,N_2627);
or U2801 (N_2801,N_2747,N_2729);
or U2802 (N_2802,N_2507,N_2506);
nor U2803 (N_2803,N_2654,N_2742);
nor U2804 (N_2804,N_2623,N_2630);
nor U2805 (N_2805,N_2701,N_2700);
nor U2806 (N_2806,N_2598,N_2510);
and U2807 (N_2807,N_2534,N_2593);
and U2808 (N_2808,N_2744,N_2512);
and U2809 (N_2809,N_2525,N_2679);
nand U2810 (N_2810,N_2749,N_2690);
xnor U2811 (N_2811,N_2738,N_2748);
nor U2812 (N_2812,N_2637,N_2709);
or U2813 (N_2813,N_2737,N_2745);
nor U2814 (N_2814,N_2672,N_2500);
or U2815 (N_2815,N_2676,N_2661);
and U2816 (N_2816,N_2597,N_2693);
nor U2817 (N_2817,N_2528,N_2609);
and U2818 (N_2818,N_2715,N_2584);
or U2819 (N_2819,N_2644,N_2659);
and U2820 (N_2820,N_2702,N_2658);
xnor U2821 (N_2821,N_2667,N_2518);
xnor U2822 (N_2822,N_2710,N_2638);
and U2823 (N_2823,N_2616,N_2541);
nor U2824 (N_2824,N_2552,N_2514);
or U2825 (N_2825,N_2588,N_2668);
nand U2826 (N_2826,N_2714,N_2570);
nor U2827 (N_2827,N_2606,N_2547);
nor U2828 (N_2828,N_2669,N_2575);
and U2829 (N_2829,N_2542,N_2622);
xnor U2830 (N_2830,N_2567,N_2670);
or U2831 (N_2831,N_2564,N_2595);
and U2832 (N_2832,N_2526,N_2524);
nand U2833 (N_2833,N_2533,N_2555);
or U2834 (N_2834,N_2586,N_2577);
nor U2835 (N_2835,N_2565,N_2716);
or U2836 (N_2836,N_2677,N_2596);
nor U2837 (N_2837,N_2604,N_2641);
nand U2838 (N_2838,N_2687,N_2513);
and U2839 (N_2839,N_2538,N_2539);
xnor U2840 (N_2840,N_2746,N_2594);
xor U2841 (N_2841,N_2739,N_2725);
xor U2842 (N_2842,N_2621,N_2603);
and U2843 (N_2843,N_2642,N_2585);
nand U2844 (N_2844,N_2522,N_2501);
nor U2845 (N_2845,N_2694,N_2548);
and U2846 (N_2846,N_2557,N_2568);
xnor U2847 (N_2847,N_2614,N_2579);
nor U2848 (N_2848,N_2735,N_2566);
and U2849 (N_2849,N_2505,N_2671);
nor U2850 (N_2850,N_2647,N_2559);
nand U2851 (N_2851,N_2536,N_2655);
and U2852 (N_2852,N_2521,N_2639);
xor U2853 (N_2853,N_2682,N_2652);
xnor U2854 (N_2854,N_2724,N_2572);
nor U2855 (N_2855,N_2517,N_2516);
nand U2856 (N_2856,N_2553,N_2628);
or U2857 (N_2857,N_2648,N_2650);
nand U2858 (N_2858,N_2646,N_2504);
nand U2859 (N_2859,N_2673,N_2680);
and U2860 (N_2860,N_2720,N_2520);
or U2861 (N_2861,N_2656,N_2569);
nor U2862 (N_2862,N_2695,N_2636);
or U2863 (N_2863,N_2515,N_2708);
xnor U2864 (N_2864,N_2635,N_2530);
xnor U2865 (N_2865,N_2607,N_2576);
nor U2866 (N_2866,N_2591,N_2543);
and U2867 (N_2867,N_2540,N_2554);
xor U2868 (N_2868,N_2556,N_2681);
nor U2869 (N_2869,N_2508,N_2741);
and U2870 (N_2870,N_2535,N_2537);
or U2871 (N_2871,N_2645,N_2688);
xnor U2872 (N_2872,N_2511,N_2666);
nand U2873 (N_2873,N_2684,N_2731);
or U2874 (N_2874,N_2578,N_2613);
or U2875 (N_2875,N_2548,N_2545);
nor U2876 (N_2876,N_2728,N_2596);
nor U2877 (N_2877,N_2562,N_2730);
xor U2878 (N_2878,N_2530,N_2521);
nor U2879 (N_2879,N_2573,N_2510);
nor U2880 (N_2880,N_2664,N_2700);
xor U2881 (N_2881,N_2715,N_2624);
or U2882 (N_2882,N_2689,N_2595);
nor U2883 (N_2883,N_2706,N_2673);
or U2884 (N_2884,N_2680,N_2654);
or U2885 (N_2885,N_2522,N_2687);
nand U2886 (N_2886,N_2579,N_2664);
xnor U2887 (N_2887,N_2689,N_2686);
nand U2888 (N_2888,N_2516,N_2555);
nand U2889 (N_2889,N_2546,N_2623);
and U2890 (N_2890,N_2557,N_2627);
nand U2891 (N_2891,N_2552,N_2618);
and U2892 (N_2892,N_2583,N_2531);
nand U2893 (N_2893,N_2651,N_2703);
nand U2894 (N_2894,N_2735,N_2694);
nand U2895 (N_2895,N_2592,N_2711);
and U2896 (N_2896,N_2694,N_2618);
or U2897 (N_2897,N_2741,N_2606);
nor U2898 (N_2898,N_2584,N_2654);
nor U2899 (N_2899,N_2650,N_2744);
nand U2900 (N_2900,N_2637,N_2740);
or U2901 (N_2901,N_2712,N_2561);
nor U2902 (N_2902,N_2540,N_2656);
xnor U2903 (N_2903,N_2670,N_2565);
xnor U2904 (N_2904,N_2528,N_2515);
xor U2905 (N_2905,N_2745,N_2602);
nor U2906 (N_2906,N_2543,N_2542);
xor U2907 (N_2907,N_2622,N_2527);
or U2908 (N_2908,N_2722,N_2605);
xnor U2909 (N_2909,N_2654,N_2691);
or U2910 (N_2910,N_2685,N_2591);
or U2911 (N_2911,N_2699,N_2592);
and U2912 (N_2912,N_2713,N_2517);
nand U2913 (N_2913,N_2600,N_2690);
and U2914 (N_2914,N_2740,N_2502);
and U2915 (N_2915,N_2526,N_2502);
nor U2916 (N_2916,N_2668,N_2709);
nand U2917 (N_2917,N_2643,N_2556);
or U2918 (N_2918,N_2574,N_2562);
nor U2919 (N_2919,N_2561,N_2709);
and U2920 (N_2920,N_2672,N_2652);
xnor U2921 (N_2921,N_2738,N_2640);
nand U2922 (N_2922,N_2534,N_2659);
xor U2923 (N_2923,N_2536,N_2601);
xnor U2924 (N_2924,N_2560,N_2607);
or U2925 (N_2925,N_2563,N_2718);
nand U2926 (N_2926,N_2680,N_2541);
or U2927 (N_2927,N_2610,N_2644);
xor U2928 (N_2928,N_2748,N_2506);
nor U2929 (N_2929,N_2641,N_2729);
or U2930 (N_2930,N_2665,N_2663);
xnor U2931 (N_2931,N_2686,N_2733);
nor U2932 (N_2932,N_2681,N_2722);
nand U2933 (N_2933,N_2573,N_2697);
xnor U2934 (N_2934,N_2621,N_2646);
nor U2935 (N_2935,N_2522,N_2737);
or U2936 (N_2936,N_2531,N_2726);
and U2937 (N_2937,N_2655,N_2717);
or U2938 (N_2938,N_2704,N_2695);
nand U2939 (N_2939,N_2654,N_2747);
xnor U2940 (N_2940,N_2654,N_2534);
and U2941 (N_2941,N_2608,N_2538);
xor U2942 (N_2942,N_2648,N_2538);
xor U2943 (N_2943,N_2736,N_2558);
nor U2944 (N_2944,N_2651,N_2713);
and U2945 (N_2945,N_2636,N_2735);
and U2946 (N_2946,N_2718,N_2542);
nor U2947 (N_2947,N_2666,N_2519);
or U2948 (N_2948,N_2686,N_2650);
nand U2949 (N_2949,N_2572,N_2501);
nand U2950 (N_2950,N_2593,N_2694);
and U2951 (N_2951,N_2555,N_2529);
and U2952 (N_2952,N_2669,N_2574);
and U2953 (N_2953,N_2647,N_2664);
and U2954 (N_2954,N_2668,N_2722);
xnor U2955 (N_2955,N_2597,N_2557);
nand U2956 (N_2956,N_2640,N_2513);
nand U2957 (N_2957,N_2695,N_2614);
and U2958 (N_2958,N_2604,N_2720);
and U2959 (N_2959,N_2613,N_2726);
nor U2960 (N_2960,N_2538,N_2683);
nor U2961 (N_2961,N_2632,N_2652);
and U2962 (N_2962,N_2554,N_2655);
xnor U2963 (N_2963,N_2632,N_2612);
nand U2964 (N_2964,N_2728,N_2670);
nor U2965 (N_2965,N_2623,N_2654);
and U2966 (N_2966,N_2503,N_2522);
nand U2967 (N_2967,N_2629,N_2736);
nand U2968 (N_2968,N_2668,N_2527);
xor U2969 (N_2969,N_2572,N_2641);
nand U2970 (N_2970,N_2513,N_2623);
or U2971 (N_2971,N_2523,N_2670);
nand U2972 (N_2972,N_2611,N_2721);
or U2973 (N_2973,N_2511,N_2677);
nor U2974 (N_2974,N_2600,N_2581);
nor U2975 (N_2975,N_2728,N_2574);
or U2976 (N_2976,N_2635,N_2708);
nand U2977 (N_2977,N_2749,N_2519);
xnor U2978 (N_2978,N_2506,N_2633);
nor U2979 (N_2979,N_2594,N_2626);
nand U2980 (N_2980,N_2531,N_2634);
xor U2981 (N_2981,N_2653,N_2508);
nand U2982 (N_2982,N_2521,N_2718);
xnor U2983 (N_2983,N_2623,N_2607);
nor U2984 (N_2984,N_2636,N_2646);
nor U2985 (N_2985,N_2559,N_2585);
xor U2986 (N_2986,N_2571,N_2556);
or U2987 (N_2987,N_2559,N_2631);
nand U2988 (N_2988,N_2640,N_2605);
or U2989 (N_2989,N_2693,N_2648);
nor U2990 (N_2990,N_2730,N_2686);
nand U2991 (N_2991,N_2635,N_2650);
nand U2992 (N_2992,N_2670,N_2597);
nor U2993 (N_2993,N_2530,N_2654);
nand U2994 (N_2994,N_2632,N_2715);
nand U2995 (N_2995,N_2616,N_2565);
nor U2996 (N_2996,N_2714,N_2504);
or U2997 (N_2997,N_2701,N_2644);
and U2998 (N_2998,N_2534,N_2527);
nand U2999 (N_2999,N_2621,N_2559);
and U3000 (N_3000,N_2752,N_2825);
and U3001 (N_3001,N_2780,N_2760);
nor U3002 (N_3002,N_2824,N_2893);
nand U3003 (N_3003,N_2977,N_2890);
xnor U3004 (N_3004,N_2902,N_2971);
and U3005 (N_3005,N_2910,N_2874);
xnor U3006 (N_3006,N_2914,N_2815);
nor U3007 (N_3007,N_2771,N_2882);
nor U3008 (N_3008,N_2932,N_2940);
xnor U3009 (N_3009,N_2952,N_2949);
nand U3010 (N_3010,N_2983,N_2966);
nand U3011 (N_3011,N_2984,N_2770);
nor U3012 (N_3012,N_2931,N_2895);
or U3013 (N_3013,N_2772,N_2998);
xnor U3014 (N_3014,N_2894,N_2967);
nand U3015 (N_3015,N_2816,N_2935);
or U3016 (N_3016,N_2963,N_2887);
or U3017 (N_3017,N_2997,N_2828);
or U3018 (N_3018,N_2797,N_2805);
xor U3019 (N_3019,N_2776,N_2833);
nand U3020 (N_3020,N_2988,N_2858);
nand U3021 (N_3021,N_2899,N_2958);
nand U3022 (N_3022,N_2991,N_2925);
nor U3023 (N_3023,N_2996,N_2981);
or U3024 (N_3024,N_2853,N_2994);
xnor U3025 (N_3025,N_2809,N_2827);
nor U3026 (N_3026,N_2927,N_2830);
nor U3027 (N_3027,N_2870,N_2869);
xor U3028 (N_3028,N_2905,N_2802);
nand U3029 (N_3029,N_2938,N_2908);
and U3030 (N_3030,N_2856,N_2775);
or U3031 (N_3031,N_2982,N_2987);
nor U3032 (N_3032,N_2970,N_2754);
nor U3033 (N_3033,N_2992,N_2916);
nand U3034 (N_3034,N_2785,N_2876);
nor U3035 (N_3035,N_2959,N_2912);
and U3036 (N_3036,N_2803,N_2884);
nand U3037 (N_3037,N_2814,N_2821);
xnor U3038 (N_3038,N_2961,N_2791);
or U3039 (N_3039,N_2753,N_2964);
nand U3040 (N_3040,N_2751,N_2843);
nor U3041 (N_3041,N_2778,N_2855);
or U3042 (N_3042,N_2857,N_2948);
or U3043 (N_3043,N_2784,N_2980);
xor U3044 (N_3044,N_2946,N_2906);
or U3045 (N_3045,N_2919,N_2817);
xnor U3046 (N_3046,N_2877,N_2755);
nor U3047 (N_3047,N_2936,N_2937);
nor U3048 (N_3048,N_2807,N_2800);
and U3049 (N_3049,N_2781,N_2873);
nand U3050 (N_3050,N_2818,N_2774);
nor U3051 (N_3051,N_2831,N_2757);
nand U3052 (N_3052,N_2768,N_2832);
xor U3053 (N_3053,N_2993,N_2954);
nand U3054 (N_3054,N_2889,N_2974);
and U3055 (N_3055,N_2806,N_2872);
nor U3056 (N_3056,N_2786,N_2903);
or U3057 (N_3057,N_2866,N_2897);
and U3058 (N_3058,N_2922,N_2849);
and U3059 (N_3059,N_2837,N_2978);
and U3060 (N_3060,N_2947,N_2841);
and U3061 (N_3061,N_2883,N_2792);
or U3062 (N_3062,N_2799,N_2808);
nor U3063 (N_3063,N_2955,N_2864);
nand U3064 (N_3064,N_2926,N_2813);
and U3065 (N_3065,N_2852,N_2846);
nand U3066 (N_3066,N_2999,N_2933);
xnor U3067 (N_3067,N_2823,N_2979);
nand U3068 (N_3068,N_2787,N_2962);
nor U3069 (N_3069,N_2811,N_2801);
nor U3070 (N_3070,N_2860,N_2795);
nor U3071 (N_3071,N_2756,N_2779);
and U3072 (N_3072,N_2995,N_2915);
or U3073 (N_3073,N_2838,N_2920);
nor U3074 (N_3074,N_2879,N_2759);
and U3075 (N_3075,N_2796,N_2763);
nor U3076 (N_3076,N_2851,N_2924);
and U3077 (N_3077,N_2904,N_2812);
xnor U3078 (N_3078,N_2941,N_2945);
nor U3079 (N_3079,N_2875,N_2975);
and U3080 (N_3080,N_2794,N_2867);
nand U3081 (N_3081,N_2842,N_2826);
xnor U3082 (N_3082,N_2868,N_2848);
and U3083 (N_3083,N_2976,N_2892);
and U3084 (N_3084,N_2764,N_2942);
and U3085 (N_3085,N_2845,N_2769);
nor U3086 (N_3086,N_2834,N_2790);
and U3087 (N_3087,N_2973,N_2844);
nand U3088 (N_3088,N_2944,N_2835);
nand U3089 (N_3089,N_2953,N_2782);
and U3090 (N_3090,N_2863,N_2839);
xor U3091 (N_3091,N_2957,N_2777);
nand U3092 (N_3092,N_2819,N_2901);
and U3093 (N_3093,N_2750,N_2871);
nor U3094 (N_3094,N_2886,N_2985);
nand U3095 (N_3095,N_2859,N_2972);
or U3096 (N_3096,N_2990,N_2934);
nor U3097 (N_3097,N_2798,N_2921);
and U3098 (N_3098,N_2822,N_2951);
nor U3099 (N_3099,N_2930,N_2854);
xnor U3100 (N_3100,N_2939,N_2758);
nor U3101 (N_3101,N_2783,N_2888);
or U3102 (N_3102,N_2896,N_2766);
nand U3103 (N_3103,N_2960,N_2850);
and U3104 (N_3104,N_2881,N_2898);
xor U3105 (N_3105,N_2986,N_2928);
nor U3106 (N_3106,N_2761,N_2810);
nand U3107 (N_3107,N_2773,N_2917);
and U3108 (N_3108,N_2865,N_2918);
xor U3109 (N_3109,N_2965,N_2891);
nand U3110 (N_3110,N_2885,N_2968);
nand U3111 (N_3111,N_2911,N_2956);
xor U3112 (N_3112,N_2880,N_2788);
and U3113 (N_3113,N_2861,N_2793);
xnor U3114 (N_3114,N_2943,N_2929);
nor U3115 (N_3115,N_2907,N_2847);
nand U3116 (N_3116,N_2862,N_2820);
or U3117 (N_3117,N_2989,N_2923);
or U3118 (N_3118,N_2913,N_2950);
xnor U3119 (N_3119,N_2900,N_2909);
and U3120 (N_3120,N_2836,N_2765);
and U3121 (N_3121,N_2789,N_2762);
nand U3122 (N_3122,N_2829,N_2767);
xor U3123 (N_3123,N_2840,N_2878);
xnor U3124 (N_3124,N_2804,N_2969);
nand U3125 (N_3125,N_2985,N_2986);
and U3126 (N_3126,N_2879,N_2975);
or U3127 (N_3127,N_2981,N_2844);
nand U3128 (N_3128,N_2899,N_2842);
nand U3129 (N_3129,N_2948,N_2932);
or U3130 (N_3130,N_2924,N_2910);
nand U3131 (N_3131,N_2841,N_2962);
or U3132 (N_3132,N_2750,N_2766);
nor U3133 (N_3133,N_2783,N_2777);
and U3134 (N_3134,N_2788,N_2769);
and U3135 (N_3135,N_2975,N_2768);
and U3136 (N_3136,N_2884,N_2785);
and U3137 (N_3137,N_2899,N_2996);
or U3138 (N_3138,N_2965,N_2756);
xnor U3139 (N_3139,N_2989,N_2992);
xnor U3140 (N_3140,N_2947,N_2866);
or U3141 (N_3141,N_2980,N_2796);
nand U3142 (N_3142,N_2806,N_2915);
nor U3143 (N_3143,N_2878,N_2993);
nand U3144 (N_3144,N_2899,N_2888);
nand U3145 (N_3145,N_2986,N_2954);
or U3146 (N_3146,N_2814,N_2802);
nand U3147 (N_3147,N_2884,N_2831);
xor U3148 (N_3148,N_2920,N_2965);
nor U3149 (N_3149,N_2866,N_2854);
nand U3150 (N_3150,N_2850,N_2796);
and U3151 (N_3151,N_2994,N_2803);
nor U3152 (N_3152,N_2808,N_2952);
xor U3153 (N_3153,N_2774,N_2806);
or U3154 (N_3154,N_2996,N_2907);
or U3155 (N_3155,N_2926,N_2958);
xnor U3156 (N_3156,N_2923,N_2787);
xor U3157 (N_3157,N_2903,N_2750);
nand U3158 (N_3158,N_2864,N_2913);
or U3159 (N_3159,N_2982,N_2988);
nand U3160 (N_3160,N_2868,N_2875);
nand U3161 (N_3161,N_2897,N_2756);
and U3162 (N_3162,N_2981,N_2914);
xor U3163 (N_3163,N_2944,N_2868);
and U3164 (N_3164,N_2989,N_2945);
nor U3165 (N_3165,N_2981,N_2937);
or U3166 (N_3166,N_2911,N_2851);
nor U3167 (N_3167,N_2876,N_2840);
xor U3168 (N_3168,N_2761,N_2993);
or U3169 (N_3169,N_2789,N_2937);
and U3170 (N_3170,N_2800,N_2956);
or U3171 (N_3171,N_2999,N_2802);
and U3172 (N_3172,N_2768,N_2949);
nor U3173 (N_3173,N_2891,N_2893);
and U3174 (N_3174,N_2939,N_2907);
and U3175 (N_3175,N_2912,N_2968);
and U3176 (N_3176,N_2777,N_2932);
xor U3177 (N_3177,N_2874,N_2816);
or U3178 (N_3178,N_2976,N_2917);
nand U3179 (N_3179,N_2809,N_2873);
or U3180 (N_3180,N_2827,N_2905);
nor U3181 (N_3181,N_2778,N_2764);
nand U3182 (N_3182,N_2874,N_2814);
or U3183 (N_3183,N_2788,N_2957);
or U3184 (N_3184,N_2833,N_2899);
or U3185 (N_3185,N_2821,N_2910);
nor U3186 (N_3186,N_2953,N_2819);
xor U3187 (N_3187,N_2843,N_2847);
nand U3188 (N_3188,N_2872,N_2941);
and U3189 (N_3189,N_2980,N_2825);
and U3190 (N_3190,N_2944,N_2893);
nor U3191 (N_3191,N_2831,N_2917);
nand U3192 (N_3192,N_2753,N_2798);
or U3193 (N_3193,N_2826,N_2763);
nand U3194 (N_3194,N_2838,N_2935);
xor U3195 (N_3195,N_2951,N_2767);
nand U3196 (N_3196,N_2846,N_2779);
or U3197 (N_3197,N_2995,N_2863);
and U3198 (N_3198,N_2834,N_2828);
xor U3199 (N_3199,N_2809,N_2994);
nand U3200 (N_3200,N_2815,N_2986);
and U3201 (N_3201,N_2886,N_2791);
or U3202 (N_3202,N_2977,N_2898);
or U3203 (N_3203,N_2954,N_2990);
or U3204 (N_3204,N_2802,N_2765);
and U3205 (N_3205,N_2835,N_2958);
nor U3206 (N_3206,N_2799,N_2833);
nand U3207 (N_3207,N_2826,N_2986);
nor U3208 (N_3208,N_2827,N_2929);
or U3209 (N_3209,N_2786,N_2897);
and U3210 (N_3210,N_2828,N_2774);
nand U3211 (N_3211,N_2871,N_2909);
and U3212 (N_3212,N_2770,N_2970);
or U3213 (N_3213,N_2973,N_2865);
and U3214 (N_3214,N_2964,N_2954);
xor U3215 (N_3215,N_2829,N_2793);
nand U3216 (N_3216,N_2999,N_2845);
xor U3217 (N_3217,N_2905,N_2855);
or U3218 (N_3218,N_2972,N_2871);
xnor U3219 (N_3219,N_2948,N_2813);
and U3220 (N_3220,N_2773,N_2781);
nor U3221 (N_3221,N_2897,N_2999);
nor U3222 (N_3222,N_2943,N_2893);
and U3223 (N_3223,N_2802,N_2858);
or U3224 (N_3224,N_2814,N_2893);
and U3225 (N_3225,N_2951,N_2807);
nor U3226 (N_3226,N_2991,N_2820);
or U3227 (N_3227,N_2903,N_2860);
nand U3228 (N_3228,N_2797,N_2766);
or U3229 (N_3229,N_2824,N_2970);
nand U3230 (N_3230,N_2981,N_2986);
nand U3231 (N_3231,N_2793,N_2878);
nor U3232 (N_3232,N_2754,N_2778);
xnor U3233 (N_3233,N_2771,N_2926);
xor U3234 (N_3234,N_2834,N_2966);
or U3235 (N_3235,N_2872,N_2967);
nor U3236 (N_3236,N_2945,N_2908);
and U3237 (N_3237,N_2845,N_2855);
or U3238 (N_3238,N_2921,N_2759);
xnor U3239 (N_3239,N_2845,N_2939);
and U3240 (N_3240,N_2948,N_2830);
nor U3241 (N_3241,N_2881,N_2985);
nand U3242 (N_3242,N_2993,N_2977);
and U3243 (N_3243,N_2759,N_2899);
nor U3244 (N_3244,N_2795,N_2867);
nor U3245 (N_3245,N_2753,N_2845);
nor U3246 (N_3246,N_2798,N_2879);
and U3247 (N_3247,N_2836,N_2886);
nand U3248 (N_3248,N_2839,N_2945);
nor U3249 (N_3249,N_2754,N_2957);
or U3250 (N_3250,N_3058,N_3238);
or U3251 (N_3251,N_3249,N_3118);
or U3252 (N_3252,N_3237,N_3092);
xor U3253 (N_3253,N_3038,N_3245);
xnor U3254 (N_3254,N_3147,N_3207);
nand U3255 (N_3255,N_3088,N_3208);
nand U3256 (N_3256,N_3137,N_3043);
nand U3257 (N_3257,N_3091,N_3124);
and U3258 (N_3258,N_3136,N_3093);
and U3259 (N_3259,N_3046,N_3212);
xnor U3260 (N_3260,N_3177,N_3206);
or U3261 (N_3261,N_3050,N_3047);
nand U3262 (N_3262,N_3142,N_3102);
xnor U3263 (N_3263,N_3191,N_3174);
xor U3264 (N_3264,N_3014,N_3133);
xnor U3265 (N_3265,N_3157,N_3134);
or U3266 (N_3266,N_3203,N_3227);
nor U3267 (N_3267,N_3200,N_3016);
nand U3268 (N_3268,N_3117,N_3051);
and U3269 (N_3269,N_3247,N_3153);
and U3270 (N_3270,N_3108,N_3195);
nor U3271 (N_3271,N_3151,N_3004);
nor U3272 (N_3272,N_3018,N_3034);
nor U3273 (N_3273,N_3010,N_3183);
and U3274 (N_3274,N_3175,N_3022);
and U3275 (N_3275,N_3193,N_3064);
or U3276 (N_3276,N_3055,N_3216);
and U3277 (N_3277,N_3218,N_3094);
nor U3278 (N_3278,N_3170,N_3128);
xor U3279 (N_3279,N_3192,N_3156);
and U3280 (N_3280,N_3244,N_3221);
nand U3281 (N_3281,N_3052,N_3048);
or U3282 (N_3282,N_3150,N_3072);
nand U3283 (N_3283,N_3057,N_3190);
nand U3284 (N_3284,N_3225,N_3205);
or U3285 (N_3285,N_3148,N_3180);
and U3286 (N_3286,N_3029,N_3103);
or U3287 (N_3287,N_3146,N_3032);
nor U3288 (N_3288,N_3025,N_3239);
xor U3289 (N_3289,N_3197,N_3228);
or U3290 (N_3290,N_3235,N_3054);
or U3291 (N_3291,N_3063,N_3067);
xnor U3292 (N_3292,N_3161,N_3021);
or U3293 (N_3293,N_3158,N_3083);
xor U3294 (N_3294,N_3223,N_3005);
or U3295 (N_3295,N_3155,N_3104);
or U3296 (N_3296,N_3166,N_3074);
or U3297 (N_3297,N_3111,N_3220);
xor U3298 (N_3298,N_3209,N_3028);
and U3299 (N_3299,N_3009,N_3100);
and U3300 (N_3300,N_3179,N_3248);
and U3301 (N_3301,N_3226,N_3084);
or U3302 (N_3302,N_3178,N_3199);
nor U3303 (N_3303,N_3187,N_3070);
or U3304 (N_3304,N_3098,N_3138);
or U3305 (N_3305,N_3086,N_3246);
and U3306 (N_3306,N_3123,N_3078);
nor U3307 (N_3307,N_3107,N_3017);
nor U3308 (N_3308,N_3131,N_3075);
nand U3309 (N_3309,N_3140,N_3096);
xnor U3310 (N_3310,N_3236,N_3020);
or U3311 (N_3311,N_3154,N_3068);
or U3312 (N_3312,N_3113,N_3119);
xnor U3313 (N_3313,N_3186,N_3061);
xor U3314 (N_3314,N_3152,N_3090);
and U3315 (N_3315,N_3087,N_3030);
or U3316 (N_3316,N_3015,N_3184);
xnor U3317 (N_3317,N_3230,N_3233);
xnor U3318 (N_3318,N_3143,N_3172);
nor U3319 (N_3319,N_3234,N_3196);
or U3320 (N_3320,N_3066,N_3112);
or U3321 (N_3321,N_3132,N_3085);
and U3322 (N_3322,N_3006,N_3039);
nor U3323 (N_3323,N_3003,N_3173);
or U3324 (N_3324,N_3026,N_3149);
nand U3325 (N_3325,N_3243,N_3144);
or U3326 (N_3326,N_3232,N_3115);
nor U3327 (N_3327,N_3027,N_3000);
nor U3328 (N_3328,N_3012,N_3210);
nand U3329 (N_3329,N_3031,N_3194);
and U3330 (N_3330,N_3163,N_3019);
xor U3331 (N_3331,N_3201,N_3049);
or U3332 (N_3332,N_3229,N_3167);
or U3333 (N_3333,N_3007,N_3073);
or U3334 (N_3334,N_3164,N_3171);
nand U3335 (N_3335,N_3219,N_3041);
nor U3336 (N_3336,N_3109,N_3224);
xor U3337 (N_3337,N_3116,N_3242);
or U3338 (N_3338,N_3069,N_3106);
or U3339 (N_3339,N_3129,N_3077);
xor U3340 (N_3340,N_3071,N_3145);
nand U3341 (N_3341,N_3169,N_3122);
and U3342 (N_3342,N_3099,N_3079);
nor U3343 (N_3343,N_3080,N_3002);
nor U3344 (N_3344,N_3044,N_3198);
xnor U3345 (N_3345,N_3125,N_3105);
nand U3346 (N_3346,N_3182,N_3231);
xnor U3347 (N_3347,N_3040,N_3141);
nor U3348 (N_3348,N_3062,N_3222);
or U3349 (N_3349,N_3160,N_3176);
nor U3350 (N_3350,N_3065,N_3037);
or U3351 (N_3351,N_3053,N_3013);
nor U3352 (N_3352,N_3240,N_3188);
or U3353 (N_3353,N_3082,N_3011);
nor U3354 (N_3354,N_3023,N_3127);
xnor U3355 (N_3355,N_3130,N_3135);
nand U3356 (N_3356,N_3101,N_3089);
and U3357 (N_3357,N_3204,N_3211);
nand U3358 (N_3358,N_3213,N_3202);
and U3359 (N_3359,N_3081,N_3185);
nand U3360 (N_3360,N_3114,N_3042);
nor U3361 (N_3361,N_3036,N_3060);
nor U3362 (N_3362,N_3008,N_3189);
and U3363 (N_3363,N_3159,N_3024);
or U3364 (N_3364,N_3165,N_3120);
nor U3365 (N_3365,N_3139,N_3033);
and U3366 (N_3366,N_3214,N_3045);
nand U3367 (N_3367,N_3001,N_3215);
and U3368 (N_3368,N_3056,N_3095);
and U3369 (N_3369,N_3217,N_3035);
nor U3370 (N_3370,N_3241,N_3181);
and U3371 (N_3371,N_3097,N_3076);
and U3372 (N_3372,N_3059,N_3162);
or U3373 (N_3373,N_3168,N_3126);
or U3374 (N_3374,N_3121,N_3110);
and U3375 (N_3375,N_3024,N_3223);
or U3376 (N_3376,N_3103,N_3119);
nor U3377 (N_3377,N_3013,N_3169);
xor U3378 (N_3378,N_3129,N_3161);
xor U3379 (N_3379,N_3032,N_3068);
or U3380 (N_3380,N_3017,N_3074);
and U3381 (N_3381,N_3057,N_3024);
xnor U3382 (N_3382,N_3056,N_3237);
and U3383 (N_3383,N_3124,N_3127);
or U3384 (N_3384,N_3075,N_3129);
nor U3385 (N_3385,N_3080,N_3066);
nor U3386 (N_3386,N_3209,N_3104);
or U3387 (N_3387,N_3030,N_3047);
nand U3388 (N_3388,N_3066,N_3070);
nand U3389 (N_3389,N_3120,N_3158);
xor U3390 (N_3390,N_3189,N_3103);
nand U3391 (N_3391,N_3171,N_3096);
and U3392 (N_3392,N_3216,N_3205);
nor U3393 (N_3393,N_3106,N_3012);
xor U3394 (N_3394,N_3157,N_3066);
and U3395 (N_3395,N_3205,N_3041);
and U3396 (N_3396,N_3073,N_3122);
and U3397 (N_3397,N_3231,N_3175);
xor U3398 (N_3398,N_3029,N_3134);
and U3399 (N_3399,N_3072,N_3046);
or U3400 (N_3400,N_3223,N_3241);
xnor U3401 (N_3401,N_3143,N_3179);
nor U3402 (N_3402,N_3057,N_3112);
or U3403 (N_3403,N_3138,N_3226);
nor U3404 (N_3404,N_3187,N_3013);
or U3405 (N_3405,N_3174,N_3222);
nand U3406 (N_3406,N_3176,N_3114);
xor U3407 (N_3407,N_3112,N_3073);
xor U3408 (N_3408,N_3138,N_3147);
nand U3409 (N_3409,N_3144,N_3109);
nand U3410 (N_3410,N_3229,N_3151);
and U3411 (N_3411,N_3042,N_3245);
nor U3412 (N_3412,N_3039,N_3199);
nand U3413 (N_3413,N_3144,N_3068);
nand U3414 (N_3414,N_3242,N_3020);
or U3415 (N_3415,N_3047,N_3151);
and U3416 (N_3416,N_3223,N_3128);
nand U3417 (N_3417,N_3062,N_3012);
nor U3418 (N_3418,N_3155,N_3122);
nor U3419 (N_3419,N_3196,N_3217);
or U3420 (N_3420,N_3173,N_3054);
xor U3421 (N_3421,N_3188,N_3016);
nand U3422 (N_3422,N_3023,N_3154);
xnor U3423 (N_3423,N_3212,N_3159);
or U3424 (N_3424,N_3232,N_3099);
xor U3425 (N_3425,N_3066,N_3049);
xnor U3426 (N_3426,N_3026,N_3140);
and U3427 (N_3427,N_3103,N_3213);
nor U3428 (N_3428,N_3240,N_3236);
xnor U3429 (N_3429,N_3023,N_3039);
and U3430 (N_3430,N_3087,N_3155);
xnor U3431 (N_3431,N_3219,N_3168);
or U3432 (N_3432,N_3037,N_3145);
and U3433 (N_3433,N_3032,N_3013);
and U3434 (N_3434,N_3169,N_3139);
nor U3435 (N_3435,N_3135,N_3062);
xor U3436 (N_3436,N_3057,N_3041);
nor U3437 (N_3437,N_3167,N_3071);
and U3438 (N_3438,N_3116,N_3034);
and U3439 (N_3439,N_3217,N_3018);
nor U3440 (N_3440,N_3249,N_3180);
nand U3441 (N_3441,N_3226,N_3197);
or U3442 (N_3442,N_3051,N_3104);
nand U3443 (N_3443,N_3183,N_3084);
or U3444 (N_3444,N_3225,N_3101);
and U3445 (N_3445,N_3015,N_3181);
nand U3446 (N_3446,N_3222,N_3003);
nand U3447 (N_3447,N_3138,N_3075);
and U3448 (N_3448,N_3226,N_3165);
nor U3449 (N_3449,N_3201,N_3057);
nor U3450 (N_3450,N_3244,N_3095);
and U3451 (N_3451,N_3137,N_3045);
and U3452 (N_3452,N_3149,N_3184);
or U3453 (N_3453,N_3071,N_3060);
xor U3454 (N_3454,N_3057,N_3177);
or U3455 (N_3455,N_3158,N_3041);
xor U3456 (N_3456,N_3148,N_3193);
or U3457 (N_3457,N_3092,N_3113);
or U3458 (N_3458,N_3028,N_3227);
xor U3459 (N_3459,N_3217,N_3156);
or U3460 (N_3460,N_3044,N_3020);
nor U3461 (N_3461,N_3136,N_3249);
or U3462 (N_3462,N_3004,N_3024);
xor U3463 (N_3463,N_3063,N_3001);
and U3464 (N_3464,N_3242,N_3016);
nor U3465 (N_3465,N_3027,N_3022);
nand U3466 (N_3466,N_3133,N_3028);
and U3467 (N_3467,N_3064,N_3091);
and U3468 (N_3468,N_3098,N_3008);
nor U3469 (N_3469,N_3042,N_3054);
nand U3470 (N_3470,N_3156,N_3115);
xnor U3471 (N_3471,N_3192,N_3114);
or U3472 (N_3472,N_3042,N_3169);
nor U3473 (N_3473,N_3045,N_3082);
nand U3474 (N_3474,N_3215,N_3134);
or U3475 (N_3475,N_3032,N_3207);
and U3476 (N_3476,N_3049,N_3060);
or U3477 (N_3477,N_3149,N_3181);
and U3478 (N_3478,N_3196,N_3141);
nor U3479 (N_3479,N_3031,N_3131);
nand U3480 (N_3480,N_3042,N_3241);
or U3481 (N_3481,N_3090,N_3036);
or U3482 (N_3482,N_3074,N_3111);
nor U3483 (N_3483,N_3085,N_3168);
nand U3484 (N_3484,N_3249,N_3041);
nand U3485 (N_3485,N_3019,N_3079);
nor U3486 (N_3486,N_3094,N_3165);
nand U3487 (N_3487,N_3219,N_3024);
nand U3488 (N_3488,N_3067,N_3192);
nand U3489 (N_3489,N_3117,N_3037);
and U3490 (N_3490,N_3172,N_3151);
xnor U3491 (N_3491,N_3040,N_3041);
and U3492 (N_3492,N_3026,N_3233);
or U3493 (N_3493,N_3182,N_3022);
nand U3494 (N_3494,N_3009,N_3068);
xnor U3495 (N_3495,N_3039,N_3084);
or U3496 (N_3496,N_3193,N_3026);
nand U3497 (N_3497,N_3119,N_3179);
xor U3498 (N_3498,N_3082,N_3001);
xor U3499 (N_3499,N_3065,N_3032);
nor U3500 (N_3500,N_3425,N_3495);
or U3501 (N_3501,N_3436,N_3309);
and U3502 (N_3502,N_3492,N_3255);
nand U3503 (N_3503,N_3479,N_3493);
nand U3504 (N_3504,N_3481,N_3362);
and U3505 (N_3505,N_3339,N_3369);
and U3506 (N_3506,N_3423,N_3424);
nor U3507 (N_3507,N_3464,N_3389);
xnor U3508 (N_3508,N_3406,N_3461);
or U3509 (N_3509,N_3494,N_3471);
nor U3510 (N_3510,N_3390,N_3416);
and U3511 (N_3511,N_3364,N_3407);
nor U3512 (N_3512,N_3330,N_3378);
or U3513 (N_3513,N_3395,N_3371);
nor U3514 (N_3514,N_3392,N_3289);
or U3515 (N_3515,N_3281,N_3463);
nor U3516 (N_3516,N_3284,N_3473);
or U3517 (N_3517,N_3365,N_3264);
nand U3518 (N_3518,N_3460,N_3270);
nand U3519 (N_3519,N_3363,N_3344);
nor U3520 (N_3520,N_3429,N_3311);
nand U3521 (N_3521,N_3455,N_3312);
nor U3522 (N_3522,N_3431,N_3253);
xnor U3523 (N_3523,N_3262,N_3469);
nand U3524 (N_3524,N_3306,N_3250);
nand U3525 (N_3525,N_3408,N_3279);
and U3526 (N_3526,N_3437,N_3432);
nand U3527 (N_3527,N_3329,N_3334);
xor U3528 (N_3528,N_3440,N_3490);
xor U3529 (N_3529,N_3428,N_3417);
and U3530 (N_3530,N_3295,N_3486);
or U3531 (N_3531,N_3263,N_3442);
or U3532 (N_3532,N_3265,N_3487);
nor U3533 (N_3533,N_3458,N_3393);
xor U3534 (N_3534,N_3256,N_3433);
nor U3535 (N_3535,N_3405,N_3475);
or U3536 (N_3536,N_3370,N_3385);
and U3537 (N_3537,N_3454,N_3497);
or U3538 (N_3538,N_3271,N_3323);
xnor U3539 (N_3539,N_3478,N_3391);
nand U3540 (N_3540,N_3489,N_3419);
or U3541 (N_3541,N_3287,N_3468);
xor U3542 (N_3542,N_3350,N_3354);
or U3543 (N_3543,N_3411,N_3360);
and U3544 (N_3544,N_3269,N_3285);
and U3545 (N_3545,N_3310,N_3485);
nor U3546 (N_3546,N_3348,N_3333);
nand U3547 (N_3547,N_3278,N_3274);
xor U3548 (N_3548,N_3465,N_3276);
nor U3549 (N_3549,N_3418,N_3317);
or U3550 (N_3550,N_3366,N_3252);
or U3551 (N_3551,N_3273,N_3450);
and U3552 (N_3552,N_3327,N_3325);
nand U3553 (N_3553,N_3452,N_3387);
nor U3554 (N_3554,N_3413,N_3380);
and U3555 (N_3555,N_3466,N_3328);
nand U3556 (N_3556,N_3474,N_3304);
or U3557 (N_3557,N_3298,N_3291);
nor U3558 (N_3558,N_3335,N_3351);
nor U3559 (N_3559,N_3403,N_3379);
xor U3560 (N_3560,N_3373,N_3449);
nor U3561 (N_3561,N_3410,N_3318);
xnor U3562 (N_3562,N_3401,N_3314);
nor U3563 (N_3563,N_3361,N_3320);
xnor U3564 (N_3564,N_3305,N_3297);
xor U3565 (N_3565,N_3377,N_3342);
nor U3566 (N_3566,N_3260,N_3375);
xor U3567 (N_3567,N_3331,N_3315);
xor U3568 (N_3568,N_3445,N_3496);
or U3569 (N_3569,N_3277,N_3352);
nor U3570 (N_3570,N_3254,N_3347);
nor U3571 (N_3571,N_3321,N_3421);
nand U3572 (N_3572,N_3343,N_3316);
nor U3573 (N_3573,N_3346,N_3482);
nor U3574 (N_3574,N_3345,N_3415);
nand U3575 (N_3575,N_3286,N_3448);
or U3576 (N_3576,N_3462,N_3319);
nor U3577 (N_3577,N_3374,N_3399);
and U3578 (N_3578,N_3400,N_3447);
xnor U3579 (N_3579,N_3355,N_3409);
or U3580 (N_3580,N_3384,N_3300);
nand U3581 (N_3581,N_3275,N_3337);
and U3582 (N_3582,N_3292,N_3357);
xnor U3583 (N_3583,N_3290,N_3484);
and U3584 (N_3584,N_3324,N_3258);
or U3585 (N_3585,N_3336,N_3457);
nor U3586 (N_3586,N_3368,N_3280);
or U3587 (N_3587,N_3422,N_3376);
nand U3588 (N_3588,N_3446,N_3439);
and U3589 (N_3589,N_3259,N_3326);
xor U3590 (N_3590,N_3426,N_3268);
nor U3591 (N_3591,N_3451,N_3476);
nand U3592 (N_3592,N_3480,N_3459);
and U3593 (N_3593,N_3435,N_3356);
and U3594 (N_3594,N_3443,N_3301);
or U3595 (N_3595,N_3308,N_3434);
and U3596 (N_3596,N_3251,N_3467);
and U3597 (N_3597,N_3358,N_3322);
xnor U3598 (N_3598,N_3444,N_3420);
nand U3599 (N_3599,N_3472,N_3272);
nand U3600 (N_3600,N_3470,N_3341);
or U3601 (N_3601,N_3288,N_3396);
xnor U3602 (N_3602,N_3372,N_3453);
or U3603 (N_3603,N_3313,N_3266);
nor U3604 (N_3604,N_3499,N_3386);
nand U3605 (N_3605,N_3488,N_3402);
nand U3606 (N_3606,N_3491,N_3353);
xnor U3607 (N_3607,N_3302,N_3261);
nor U3608 (N_3608,N_3257,N_3349);
xnor U3609 (N_3609,N_3307,N_3441);
and U3610 (N_3610,N_3412,N_3430);
nand U3611 (N_3611,N_3299,N_3294);
xor U3612 (N_3612,N_3359,N_3338);
and U3613 (N_3613,N_3398,N_3394);
nand U3614 (N_3614,N_3303,N_3498);
nand U3615 (N_3615,N_3381,N_3483);
xor U3616 (N_3616,N_3296,N_3388);
xnor U3617 (N_3617,N_3382,N_3267);
and U3618 (N_3618,N_3383,N_3456);
nor U3619 (N_3619,N_3477,N_3367);
nand U3620 (N_3620,N_3397,N_3293);
nor U3621 (N_3621,N_3414,N_3282);
and U3622 (N_3622,N_3427,N_3283);
or U3623 (N_3623,N_3340,N_3438);
nand U3624 (N_3624,N_3404,N_3332);
xor U3625 (N_3625,N_3306,N_3365);
or U3626 (N_3626,N_3254,N_3314);
xnor U3627 (N_3627,N_3343,N_3378);
xor U3628 (N_3628,N_3320,N_3316);
xor U3629 (N_3629,N_3433,N_3389);
nor U3630 (N_3630,N_3333,N_3432);
nor U3631 (N_3631,N_3490,N_3461);
nor U3632 (N_3632,N_3498,N_3306);
nor U3633 (N_3633,N_3497,N_3455);
or U3634 (N_3634,N_3432,N_3385);
nand U3635 (N_3635,N_3456,N_3253);
nand U3636 (N_3636,N_3410,N_3251);
nand U3637 (N_3637,N_3311,N_3385);
xor U3638 (N_3638,N_3465,N_3349);
nand U3639 (N_3639,N_3294,N_3327);
nor U3640 (N_3640,N_3397,N_3473);
xnor U3641 (N_3641,N_3469,N_3352);
or U3642 (N_3642,N_3432,N_3470);
xor U3643 (N_3643,N_3272,N_3266);
or U3644 (N_3644,N_3486,N_3417);
nand U3645 (N_3645,N_3386,N_3266);
or U3646 (N_3646,N_3443,N_3277);
or U3647 (N_3647,N_3339,N_3319);
and U3648 (N_3648,N_3292,N_3417);
or U3649 (N_3649,N_3353,N_3497);
nor U3650 (N_3650,N_3468,N_3285);
nor U3651 (N_3651,N_3324,N_3459);
or U3652 (N_3652,N_3389,N_3388);
nand U3653 (N_3653,N_3274,N_3378);
xor U3654 (N_3654,N_3372,N_3275);
nand U3655 (N_3655,N_3392,N_3437);
xor U3656 (N_3656,N_3269,N_3381);
or U3657 (N_3657,N_3434,N_3351);
or U3658 (N_3658,N_3338,N_3377);
and U3659 (N_3659,N_3392,N_3468);
nand U3660 (N_3660,N_3391,N_3367);
nand U3661 (N_3661,N_3448,N_3433);
nor U3662 (N_3662,N_3401,N_3380);
nand U3663 (N_3663,N_3250,N_3373);
and U3664 (N_3664,N_3434,N_3282);
nor U3665 (N_3665,N_3361,N_3497);
xor U3666 (N_3666,N_3473,N_3487);
nor U3667 (N_3667,N_3412,N_3402);
and U3668 (N_3668,N_3389,N_3497);
nor U3669 (N_3669,N_3472,N_3366);
xnor U3670 (N_3670,N_3381,N_3395);
or U3671 (N_3671,N_3341,N_3465);
nor U3672 (N_3672,N_3495,N_3275);
xor U3673 (N_3673,N_3343,N_3465);
and U3674 (N_3674,N_3307,N_3331);
or U3675 (N_3675,N_3292,N_3351);
nand U3676 (N_3676,N_3278,N_3454);
nor U3677 (N_3677,N_3405,N_3483);
or U3678 (N_3678,N_3347,N_3291);
nand U3679 (N_3679,N_3462,N_3441);
nor U3680 (N_3680,N_3299,N_3414);
nand U3681 (N_3681,N_3481,N_3448);
xor U3682 (N_3682,N_3361,N_3440);
and U3683 (N_3683,N_3373,N_3254);
xor U3684 (N_3684,N_3491,N_3329);
or U3685 (N_3685,N_3280,N_3485);
nand U3686 (N_3686,N_3319,N_3431);
nor U3687 (N_3687,N_3431,N_3474);
nand U3688 (N_3688,N_3404,N_3261);
xnor U3689 (N_3689,N_3331,N_3281);
xnor U3690 (N_3690,N_3272,N_3327);
xor U3691 (N_3691,N_3362,N_3368);
nor U3692 (N_3692,N_3373,N_3295);
or U3693 (N_3693,N_3297,N_3352);
nor U3694 (N_3694,N_3498,N_3305);
and U3695 (N_3695,N_3383,N_3277);
nor U3696 (N_3696,N_3293,N_3374);
and U3697 (N_3697,N_3436,N_3394);
or U3698 (N_3698,N_3483,N_3439);
nor U3699 (N_3699,N_3384,N_3445);
xnor U3700 (N_3700,N_3375,N_3364);
nand U3701 (N_3701,N_3485,N_3480);
or U3702 (N_3702,N_3387,N_3430);
nand U3703 (N_3703,N_3487,N_3469);
nand U3704 (N_3704,N_3444,N_3279);
or U3705 (N_3705,N_3378,N_3319);
nor U3706 (N_3706,N_3495,N_3482);
xnor U3707 (N_3707,N_3397,N_3443);
or U3708 (N_3708,N_3280,N_3430);
xnor U3709 (N_3709,N_3360,N_3483);
or U3710 (N_3710,N_3394,N_3282);
xor U3711 (N_3711,N_3332,N_3383);
nand U3712 (N_3712,N_3481,N_3327);
and U3713 (N_3713,N_3491,N_3380);
or U3714 (N_3714,N_3374,N_3466);
and U3715 (N_3715,N_3312,N_3368);
nor U3716 (N_3716,N_3284,N_3297);
nor U3717 (N_3717,N_3407,N_3424);
xnor U3718 (N_3718,N_3483,N_3377);
or U3719 (N_3719,N_3410,N_3488);
xnor U3720 (N_3720,N_3328,N_3306);
or U3721 (N_3721,N_3479,N_3454);
and U3722 (N_3722,N_3354,N_3492);
nand U3723 (N_3723,N_3329,N_3459);
nor U3724 (N_3724,N_3299,N_3269);
xnor U3725 (N_3725,N_3347,N_3355);
nand U3726 (N_3726,N_3297,N_3369);
xnor U3727 (N_3727,N_3397,N_3457);
xnor U3728 (N_3728,N_3259,N_3379);
xnor U3729 (N_3729,N_3350,N_3484);
nand U3730 (N_3730,N_3283,N_3409);
nand U3731 (N_3731,N_3405,N_3396);
nor U3732 (N_3732,N_3468,N_3319);
nor U3733 (N_3733,N_3396,N_3295);
or U3734 (N_3734,N_3261,N_3281);
or U3735 (N_3735,N_3365,N_3332);
nor U3736 (N_3736,N_3385,N_3436);
nand U3737 (N_3737,N_3467,N_3316);
nor U3738 (N_3738,N_3490,N_3274);
nand U3739 (N_3739,N_3457,N_3435);
xor U3740 (N_3740,N_3425,N_3317);
and U3741 (N_3741,N_3466,N_3417);
or U3742 (N_3742,N_3256,N_3463);
xor U3743 (N_3743,N_3428,N_3402);
and U3744 (N_3744,N_3285,N_3350);
and U3745 (N_3745,N_3474,N_3458);
or U3746 (N_3746,N_3283,N_3464);
nand U3747 (N_3747,N_3273,N_3416);
nor U3748 (N_3748,N_3458,N_3407);
nand U3749 (N_3749,N_3331,N_3272);
and U3750 (N_3750,N_3704,N_3683);
nand U3751 (N_3751,N_3669,N_3581);
or U3752 (N_3752,N_3722,N_3736);
or U3753 (N_3753,N_3530,N_3610);
nor U3754 (N_3754,N_3630,N_3588);
nand U3755 (N_3755,N_3573,N_3502);
and U3756 (N_3756,N_3519,N_3522);
and U3757 (N_3757,N_3737,N_3615);
and U3758 (N_3758,N_3526,N_3641);
nand U3759 (N_3759,N_3727,N_3734);
xor U3760 (N_3760,N_3532,N_3744);
or U3761 (N_3761,N_3720,N_3512);
xnor U3762 (N_3762,N_3620,N_3693);
and U3763 (N_3763,N_3567,N_3743);
nand U3764 (N_3764,N_3673,N_3516);
and U3765 (N_3765,N_3724,N_3679);
nor U3766 (N_3766,N_3728,N_3591);
nand U3767 (N_3767,N_3699,N_3680);
xor U3768 (N_3768,N_3583,N_3510);
and U3769 (N_3769,N_3675,N_3738);
and U3770 (N_3770,N_3569,N_3652);
nor U3771 (N_3771,N_3730,N_3623);
and U3772 (N_3772,N_3600,N_3681);
nor U3773 (N_3773,N_3646,N_3568);
and U3774 (N_3774,N_3625,N_3501);
nor U3775 (N_3775,N_3678,N_3655);
xnor U3776 (N_3776,N_3705,N_3657);
or U3777 (N_3777,N_3564,N_3701);
nand U3778 (N_3778,N_3672,N_3715);
nor U3779 (N_3779,N_3554,N_3609);
or U3780 (N_3780,N_3645,N_3595);
nor U3781 (N_3781,N_3710,N_3662);
nand U3782 (N_3782,N_3556,N_3732);
xor U3783 (N_3783,N_3674,N_3647);
or U3784 (N_3784,N_3521,N_3713);
and U3785 (N_3785,N_3515,N_3575);
xnor U3786 (N_3786,N_3636,N_3634);
nand U3787 (N_3787,N_3565,N_3700);
and U3788 (N_3788,N_3541,N_3540);
and U3789 (N_3789,N_3659,N_3542);
xnor U3790 (N_3790,N_3518,N_3686);
or U3791 (N_3791,N_3572,N_3505);
nor U3792 (N_3792,N_3702,N_3629);
or U3793 (N_3793,N_3597,N_3548);
xnor U3794 (N_3794,N_3719,N_3690);
or U3795 (N_3795,N_3513,N_3546);
xor U3796 (N_3796,N_3577,N_3692);
nor U3797 (N_3797,N_3626,N_3632);
xor U3798 (N_3798,N_3711,N_3579);
nand U3799 (N_3799,N_3716,N_3698);
xor U3800 (N_3800,N_3741,N_3534);
or U3801 (N_3801,N_3621,N_3691);
xor U3802 (N_3802,N_3566,N_3533);
nand U3803 (N_3803,N_3555,N_3687);
or U3804 (N_3804,N_3592,N_3633);
nor U3805 (N_3805,N_3605,N_3648);
xnor U3806 (N_3806,N_3653,N_3547);
or U3807 (N_3807,N_3538,N_3587);
nand U3808 (N_3808,N_3685,N_3520);
nor U3809 (N_3809,N_3525,N_3539);
nor U3810 (N_3810,N_3644,N_3658);
or U3811 (N_3811,N_3714,N_3689);
nand U3812 (N_3812,N_3557,N_3740);
nor U3813 (N_3813,N_3561,N_3523);
nand U3814 (N_3814,N_3553,N_3649);
xnor U3815 (N_3815,N_3551,N_3514);
and U3816 (N_3816,N_3617,N_3654);
nand U3817 (N_3817,N_3742,N_3593);
nand U3818 (N_3818,N_3650,N_3584);
or U3819 (N_3819,N_3739,N_3661);
or U3820 (N_3820,N_3580,N_3717);
and U3821 (N_3821,N_3718,N_3706);
or U3822 (N_3822,N_3535,N_3589);
xor U3823 (N_3823,N_3624,N_3576);
or U3824 (N_3824,N_3747,N_3614);
and U3825 (N_3825,N_3545,N_3552);
or U3826 (N_3826,N_3560,N_3723);
xnor U3827 (N_3827,N_3616,N_3570);
and U3828 (N_3828,N_3503,N_3746);
xnor U3829 (N_3829,N_3642,N_3651);
xnor U3830 (N_3830,N_3694,N_3638);
and U3831 (N_3831,N_3663,N_3612);
xor U3832 (N_3832,N_3712,N_3725);
nand U3833 (N_3833,N_3735,N_3660);
and U3834 (N_3834,N_3676,N_3618);
xnor U3835 (N_3835,N_3586,N_3606);
nor U3836 (N_3836,N_3549,N_3506);
or U3837 (N_3837,N_3598,N_3622);
xor U3838 (N_3838,N_3524,N_3517);
xor U3839 (N_3839,N_3745,N_3696);
xnor U3840 (N_3840,N_3504,N_3508);
and U3841 (N_3841,N_3709,N_3582);
nand U3842 (N_3842,N_3627,N_3639);
nor U3843 (N_3843,N_3550,N_3559);
nor U3844 (N_3844,N_3668,N_3544);
and U3845 (N_3845,N_3602,N_3599);
xnor U3846 (N_3846,N_3608,N_3585);
and U3847 (N_3847,N_3604,N_3628);
or U3848 (N_3848,N_3733,N_3731);
nor U3849 (N_3849,N_3596,N_3601);
and U3850 (N_3850,N_3677,N_3637);
xor U3851 (N_3851,N_3666,N_3603);
nor U3852 (N_3852,N_3571,N_3590);
nand U3853 (N_3853,N_3721,N_3619);
or U3854 (N_3854,N_3500,N_3665);
nor U3855 (N_3855,N_3529,N_3682);
nor U3856 (N_3856,N_3670,N_3509);
or U3857 (N_3857,N_3726,N_3631);
xor U3858 (N_3858,N_3749,N_3563);
nand U3859 (N_3859,N_3729,N_3578);
nor U3860 (N_3860,N_3536,N_3656);
nand U3861 (N_3861,N_3688,N_3664);
nor U3862 (N_3862,N_3528,N_3543);
nand U3863 (N_3863,N_3611,N_3607);
nor U3864 (N_3864,N_3594,N_3695);
nor U3865 (N_3865,N_3531,N_3562);
xnor U3866 (N_3866,N_3527,N_3558);
nand U3867 (N_3867,N_3697,N_3635);
and U3868 (N_3868,N_3507,N_3643);
and U3869 (N_3869,N_3640,N_3684);
nand U3870 (N_3870,N_3511,N_3537);
or U3871 (N_3871,N_3708,N_3671);
or U3872 (N_3872,N_3707,N_3574);
xnor U3873 (N_3873,N_3748,N_3667);
and U3874 (N_3874,N_3703,N_3613);
nand U3875 (N_3875,N_3502,N_3614);
nand U3876 (N_3876,N_3644,N_3525);
or U3877 (N_3877,N_3623,N_3737);
nor U3878 (N_3878,N_3552,N_3650);
nand U3879 (N_3879,N_3737,N_3503);
or U3880 (N_3880,N_3507,N_3631);
nand U3881 (N_3881,N_3665,N_3707);
nand U3882 (N_3882,N_3699,N_3558);
nor U3883 (N_3883,N_3509,N_3674);
nor U3884 (N_3884,N_3514,N_3722);
or U3885 (N_3885,N_3730,N_3701);
or U3886 (N_3886,N_3501,N_3512);
xnor U3887 (N_3887,N_3599,N_3676);
nor U3888 (N_3888,N_3719,N_3603);
xor U3889 (N_3889,N_3735,N_3612);
nor U3890 (N_3890,N_3574,N_3544);
xnor U3891 (N_3891,N_3523,N_3686);
and U3892 (N_3892,N_3611,N_3576);
xnor U3893 (N_3893,N_3683,N_3603);
xor U3894 (N_3894,N_3573,N_3655);
and U3895 (N_3895,N_3572,N_3603);
or U3896 (N_3896,N_3747,N_3604);
and U3897 (N_3897,N_3552,N_3738);
and U3898 (N_3898,N_3648,N_3701);
xor U3899 (N_3899,N_3617,N_3601);
nor U3900 (N_3900,N_3617,N_3641);
and U3901 (N_3901,N_3704,N_3572);
or U3902 (N_3902,N_3645,N_3562);
and U3903 (N_3903,N_3699,N_3674);
nor U3904 (N_3904,N_3534,N_3505);
and U3905 (N_3905,N_3659,N_3610);
xnor U3906 (N_3906,N_3577,N_3619);
nand U3907 (N_3907,N_3617,N_3570);
nand U3908 (N_3908,N_3633,N_3540);
nor U3909 (N_3909,N_3563,N_3507);
xnor U3910 (N_3910,N_3568,N_3585);
and U3911 (N_3911,N_3591,N_3688);
xor U3912 (N_3912,N_3662,N_3690);
nor U3913 (N_3913,N_3749,N_3744);
nand U3914 (N_3914,N_3551,N_3602);
nand U3915 (N_3915,N_3556,N_3603);
nor U3916 (N_3916,N_3685,N_3674);
xor U3917 (N_3917,N_3652,N_3702);
nor U3918 (N_3918,N_3599,N_3613);
or U3919 (N_3919,N_3674,N_3712);
nor U3920 (N_3920,N_3640,N_3669);
and U3921 (N_3921,N_3500,N_3527);
and U3922 (N_3922,N_3561,N_3521);
or U3923 (N_3923,N_3625,N_3640);
or U3924 (N_3924,N_3695,N_3678);
xnor U3925 (N_3925,N_3673,N_3595);
nand U3926 (N_3926,N_3598,N_3530);
or U3927 (N_3927,N_3735,N_3575);
or U3928 (N_3928,N_3723,N_3531);
nor U3929 (N_3929,N_3529,N_3535);
nand U3930 (N_3930,N_3606,N_3749);
nand U3931 (N_3931,N_3503,N_3537);
nor U3932 (N_3932,N_3529,N_3635);
nand U3933 (N_3933,N_3675,N_3553);
or U3934 (N_3934,N_3653,N_3658);
or U3935 (N_3935,N_3609,N_3600);
or U3936 (N_3936,N_3668,N_3704);
nand U3937 (N_3937,N_3663,N_3700);
and U3938 (N_3938,N_3674,N_3672);
nor U3939 (N_3939,N_3701,N_3748);
xnor U3940 (N_3940,N_3638,N_3630);
or U3941 (N_3941,N_3681,N_3606);
nor U3942 (N_3942,N_3541,N_3502);
nor U3943 (N_3943,N_3675,N_3708);
nand U3944 (N_3944,N_3737,N_3579);
and U3945 (N_3945,N_3515,N_3672);
xor U3946 (N_3946,N_3734,N_3690);
nor U3947 (N_3947,N_3675,N_3732);
nor U3948 (N_3948,N_3555,N_3619);
nand U3949 (N_3949,N_3679,N_3528);
nor U3950 (N_3950,N_3593,N_3530);
xnor U3951 (N_3951,N_3520,N_3641);
nor U3952 (N_3952,N_3597,N_3560);
or U3953 (N_3953,N_3666,N_3598);
nor U3954 (N_3954,N_3539,N_3572);
nor U3955 (N_3955,N_3527,N_3694);
or U3956 (N_3956,N_3543,N_3585);
or U3957 (N_3957,N_3736,N_3522);
and U3958 (N_3958,N_3631,N_3573);
nor U3959 (N_3959,N_3723,N_3565);
and U3960 (N_3960,N_3548,N_3660);
nand U3961 (N_3961,N_3670,N_3598);
nor U3962 (N_3962,N_3586,N_3659);
or U3963 (N_3963,N_3746,N_3506);
or U3964 (N_3964,N_3513,N_3621);
nor U3965 (N_3965,N_3646,N_3686);
xor U3966 (N_3966,N_3522,N_3647);
and U3967 (N_3967,N_3568,N_3668);
xnor U3968 (N_3968,N_3549,N_3511);
xnor U3969 (N_3969,N_3720,N_3697);
xor U3970 (N_3970,N_3719,N_3643);
nand U3971 (N_3971,N_3611,N_3698);
and U3972 (N_3972,N_3673,N_3505);
nor U3973 (N_3973,N_3654,N_3504);
or U3974 (N_3974,N_3657,N_3648);
and U3975 (N_3975,N_3724,N_3638);
xnor U3976 (N_3976,N_3746,N_3729);
xnor U3977 (N_3977,N_3621,N_3641);
nand U3978 (N_3978,N_3633,N_3614);
and U3979 (N_3979,N_3554,N_3680);
and U3980 (N_3980,N_3707,N_3533);
nor U3981 (N_3981,N_3658,N_3680);
or U3982 (N_3982,N_3589,N_3696);
and U3983 (N_3983,N_3674,N_3630);
nand U3984 (N_3984,N_3636,N_3640);
or U3985 (N_3985,N_3653,N_3608);
nand U3986 (N_3986,N_3727,N_3562);
nand U3987 (N_3987,N_3691,N_3650);
nand U3988 (N_3988,N_3544,N_3692);
nor U3989 (N_3989,N_3688,N_3588);
and U3990 (N_3990,N_3741,N_3602);
and U3991 (N_3991,N_3506,N_3680);
nor U3992 (N_3992,N_3653,N_3711);
and U3993 (N_3993,N_3569,N_3725);
nand U3994 (N_3994,N_3656,N_3582);
or U3995 (N_3995,N_3543,N_3510);
xnor U3996 (N_3996,N_3664,N_3581);
and U3997 (N_3997,N_3568,N_3698);
xor U3998 (N_3998,N_3663,N_3701);
xnor U3999 (N_3999,N_3622,N_3649);
and U4000 (N_4000,N_3957,N_3757);
nor U4001 (N_4001,N_3769,N_3787);
or U4002 (N_4002,N_3981,N_3986);
xnor U4003 (N_4003,N_3804,N_3930);
xor U4004 (N_4004,N_3946,N_3810);
nor U4005 (N_4005,N_3928,N_3977);
or U4006 (N_4006,N_3851,N_3833);
and U4007 (N_4007,N_3888,N_3889);
or U4008 (N_4008,N_3947,N_3868);
or U4009 (N_4009,N_3931,N_3917);
nor U4010 (N_4010,N_3963,N_3879);
and U4011 (N_4011,N_3901,N_3873);
nor U4012 (N_4012,N_3759,N_3909);
nor U4013 (N_4013,N_3980,N_3786);
nor U4014 (N_4014,N_3993,N_3751);
xnor U4015 (N_4015,N_3781,N_3794);
nor U4016 (N_4016,N_3895,N_3960);
nand U4017 (N_4017,N_3784,N_3775);
xor U4018 (N_4018,N_3972,N_3850);
and U4019 (N_4019,N_3863,N_3893);
and U4020 (N_4020,N_3860,N_3970);
xnor U4021 (N_4021,N_3773,N_3820);
nand U4022 (N_4022,N_3882,N_3830);
xnor U4023 (N_4023,N_3813,N_3958);
nor U4024 (N_4024,N_3806,N_3840);
xor U4025 (N_4025,N_3811,N_3959);
xor U4026 (N_4026,N_3932,N_3886);
and U4027 (N_4027,N_3838,N_3832);
or U4028 (N_4028,N_3831,N_3877);
nor U4029 (N_4029,N_3808,N_3941);
xor U4030 (N_4030,N_3890,N_3964);
nor U4031 (N_4031,N_3899,N_3995);
nand U4032 (N_4032,N_3793,N_3921);
or U4033 (N_4033,N_3923,N_3907);
nor U4034 (N_4034,N_3968,N_3765);
xnor U4035 (N_4035,N_3861,N_3929);
nor U4036 (N_4036,N_3989,N_3918);
and U4037 (N_4037,N_3951,N_3783);
nor U4038 (N_4038,N_3798,N_3848);
or U4039 (N_4039,N_3991,N_3797);
nor U4040 (N_4040,N_3755,N_3939);
nor U4041 (N_4041,N_3903,N_3876);
nand U4042 (N_4042,N_3953,N_3900);
and U4043 (N_4043,N_3978,N_3912);
nand U4044 (N_4044,N_3764,N_3869);
nand U4045 (N_4045,N_3845,N_3884);
xor U4046 (N_4046,N_3814,N_3817);
and U4047 (N_4047,N_3846,N_3756);
xnor U4048 (N_4048,N_3770,N_3822);
nor U4049 (N_4049,N_3824,N_3996);
xor U4050 (N_4050,N_3844,N_3763);
and U4051 (N_4051,N_3880,N_3872);
or U4052 (N_4052,N_3774,N_3815);
and U4053 (N_4053,N_3896,N_3871);
xor U4054 (N_4054,N_3916,N_3983);
nand U4055 (N_4055,N_3842,N_3782);
nand U4056 (N_4056,N_3865,N_3809);
xnor U4057 (N_4057,N_3800,N_3979);
nor U4058 (N_4058,N_3937,N_3788);
nor U4059 (N_4059,N_3906,N_3789);
nand U4060 (N_4060,N_3936,N_3927);
nor U4061 (N_4061,N_3768,N_3988);
nor U4062 (N_4062,N_3950,N_3870);
and U4063 (N_4063,N_3952,N_3761);
and U4064 (N_4064,N_3966,N_3818);
and U4065 (N_4065,N_3892,N_3922);
and U4066 (N_4066,N_3949,N_3973);
and U4067 (N_4067,N_3802,N_3945);
and U4068 (N_4068,N_3881,N_3791);
nor U4069 (N_4069,N_3902,N_3827);
nand U4070 (N_4070,N_3938,N_3841);
nor U4071 (N_4071,N_3924,N_3854);
xor U4072 (N_4072,N_3867,N_3942);
xor U4073 (N_4073,N_3976,N_3792);
nor U4074 (N_4074,N_3992,N_3962);
nor U4075 (N_4075,N_3857,N_3935);
nand U4076 (N_4076,N_3771,N_3766);
xnor U4077 (N_4077,N_3969,N_3891);
nand U4078 (N_4078,N_3777,N_3785);
nand U4079 (N_4079,N_3898,N_3762);
xor U4080 (N_4080,N_3897,N_3853);
nand U4081 (N_4081,N_3883,N_3948);
xnor U4082 (N_4082,N_3894,N_3905);
nor U4083 (N_4083,N_3955,N_3999);
nand U4084 (N_4084,N_3984,N_3750);
nand U4085 (N_4085,N_3971,N_3826);
and U4086 (N_4086,N_3911,N_3925);
xor U4087 (N_4087,N_3779,N_3855);
and U4088 (N_4088,N_3837,N_3985);
xnor U4089 (N_4089,N_3862,N_3758);
nor U4090 (N_4090,N_3760,N_3908);
nand U4091 (N_4091,N_3974,N_3944);
nor U4092 (N_4092,N_3859,N_3965);
and U4093 (N_4093,N_3778,N_3796);
nor U4094 (N_4094,N_3864,N_3803);
and U4095 (N_4095,N_3856,N_3772);
nor U4096 (N_4096,N_3975,N_3816);
and U4097 (N_4097,N_3956,N_3812);
nor U4098 (N_4098,N_3829,N_3752);
and U4099 (N_4099,N_3767,N_3998);
nor U4100 (N_4100,N_3874,N_3780);
or U4101 (N_4101,N_3843,N_3753);
nand U4102 (N_4102,N_3994,N_3828);
or U4103 (N_4103,N_3836,N_3990);
and U4104 (N_4104,N_3934,N_3904);
or U4105 (N_4105,N_3943,N_3847);
nor U4106 (N_4106,N_3807,N_3913);
xnor U4107 (N_4107,N_3790,N_3858);
xor U4108 (N_4108,N_3885,N_3819);
nor U4109 (N_4109,N_3821,N_3801);
xor U4110 (N_4110,N_3776,N_3866);
nand U4111 (N_4111,N_3835,N_3887);
nor U4112 (N_4112,N_3967,N_3805);
nor U4113 (N_4113,N_3875,N_3940);
nor U4114 (N_4114,N_3825,N_3852);
nor U4115 (N_4115,N_3823,N_3839);
and U4116 (N_4116,N_3799,N_3961);
or U4117 (N_4117,N_3754,N_3920);
or U4118 (N_4118,N_3982,N_3954);
nand U4119 (N_4119,N_3878,N_3795);
and U4120 (N_4120,N_3926,N_3834);
or U4121 (N_4121,N_3915,N_3997);
xnor U4122 (N_4122,N_3914,N_3910);
or U4123 (N_4123,N_3919,N_3987);
nor U4124 (N_4124,N_3849,N_3933);
nor U4125 (N_4125,N_3772,N_3957);
xnor U4126 (N_4126,N_3784,N_3821);
nand U4127 (N_4127,N_3938,N_3928);
nand U4128 (N_4128,N_3908,N_3926);
nor U4129 (N_4129,N_3864,N_3773);
and U4130 (N_4130,N_3759,N_3957);
xnor U4131 (N_4131,N_3852,N_3917);
nor U4132 (N_4132,N_3926,N_3835);
and U4133 (N_4133,N_3805,N_3831);
nand U4134 (N_4134,N_3936,N_3997);
and U4135 (N_4135,N_3936,N_3865);
and U4136 (N_4136,N_3930,N_3825);
nor U4137 (N_4137,N_3988,N_3888);
or U4138 (N_4138,N_3933,N_3915);
nand U4139 (N_4139,N_3973,N_3958);
and U4140 (N_4140,N_3806,N_3974);
nor U4141 (N_4141,N_3893,N_3816);
or U4142 (N_4142,N_3857,N_3778);
nand U4143 (N_4143,N_3804,N_3995);
and U4144 (N_4144,N_3884,N_3813);
xnor U4145 (N_4145,N_3767,N_3895);
and U4146 (N_4146,N_3874,N_3841);
and U4147 (N_4147,N_3927,N_3793);
or U4148 (N_4148,N_3900,N_3861);
or U4149 (N_4149,N_3978,N_3913);
nor U4150 (N_4150,N_3883,N_3834);
nand U4151 (N_4151,N_3769,N_3973);
and U4152 (N_4152,N_3899,N_3808);
xnor U4153 (N_4153,N_3980,N_3940);
or U4154 (N_4154,N_3959,N_3894);
nand U4155 (N_4155,N_3948,N_3802);
nor U4156 (N_4156,N_3964,N_3773);
and U4157 (N_4157,N_3861,N_3846);
and U4158 (N_4158,N_3882,N_3973);
or U4159 (N_4159,N_3951,N_3792);
nand U4160 (N_4160,N_3816,N_3948);
or U4161 (N_4161,N_3858,N_3992);
and U4162 (N_4162,N_3862,N_3941);
nand U4163 (N_4163,N_3960,N_3774);
xor U4164 (N_4164,N_3863,N_3834);
nand U4165 (N_4165,N_3988,N_3921);
or U4166 (N_4166,N_3814,N_3957);
nor U4167 (N_4167,N_3805,N_3791);
xor U4168 (N_4168,N_3892,N_3751);
or U4169 (N_4169,N_3861,N_3901);
xor U4170 (N_4170,N_3879,N_3851);
and U4171 (N_4171,N_3953,N_3787);
nand U4172 (N_4172,N_3881,N_3812);
and U4173 (N_4173,N_3903,N_3918);
xor U4174 (N_4174,N_3750,N_3779);
xnor U4175 (N_4175,N_3965,N_3869);
nor U4176 (N_4176,N_3833,N_3976);
or U4177 (N_4177,N_3913,N_3817);
nand U4178 (N_4178,N_3787,N_3928);
nor U4179 (N_4179,N_3801,N_3788);
or U4180 (N_4180,N_3898,N_3971);
nand U4181 (N_4181,N_3760,N_3886);
nor U4182 (N_4182,N_3772,N_3835);
and U4183 (N_4183,N_3934,N_3885);
xnor U4184 (N_4184,N_3970,N_3980);
and U4185 (N_4185,N_3964,N_3872);
and U4186 (N_4186,N_3962,N_3832);
or U4187 (N_4187,N_3827,N_3773);
and U4188 (N_4188,N_3924,N_3795);
nor U4189 (N_4189,N_3865,N_3792);
or U4190 (N_4190,N_3810,N_3960);
xor U4191 (N_4191,N_3974,N_3978);
nor U4192 (N_4192,N_3917,N_3806);
xnor U4193 (N_4193,N_3764,N_3783);
nor U4194 (N_4194,N_3888,N_3782);
or U4195 (N_4195,N_3784,N_3891);
nand U4196 (N_4196,N_3891,N_3834);
nand U4197 (N_4197,N_3899,N_3770);
nor U4198 (N_4198,N_3994,N_3924);
nand U4199 (N_4199,N_3984,N_3962);
nand U4200 (N_4200,N_3820,N_3880);
or U4201 (N_4201,N_3829,N_3955);
or U4202 (N_4202,N_3774,N_3916);
nand U4203 (N_4203,N_3780,N_3838);
nor U4204 (N_4204,N_3872,N_3902);
xor U4205 (N_4205,N_3996,N_3867);
nor U4206 (N_4206,N_3976,N_3810);
nor U4207 (N_4207,N_3935,N_3825);
xnor U4208 (N_4208,N_3754,N_3793);
and U4209 (N_4209,N_3834,N_3762);
xor U4210 (N_4210,N_3981,N_3827);
nand U4211 (N_4211,N_3790,N_3962);
and U4212 (N_4212,N_3972,N_3802);
or U4213 (N_4213,N_3836,N_3872);
or U4214 (N_4214,N_3882,N_3776);
or U4215 (N_4215,N_3871,N_3764);
and U4216 (N_4216,N_3799,N_3996);
nor U4217 (N_4217,N_3808,N_3913);
nor U4218 (N_4218,N_3907,N_3967);
and U4219 (N_4219,N_3798,N_3777);
xnor U4220 (N_4220,N_3921,N_3819);
nand U4221 (N_4221,N_3942,N_3948);
or U4222 (N_4222,N_3990,N_3796);
nor U4223 (N_4223,N_3926,N_3848);
xor U4224 (N_4224,N_3913,N_3977);
and U4225 (N_4225,N_3902,N_3879);
xnor U4226 (N_4226,N_3979,N_3941);
or U4227 (N_4227,N_3886,N_3864);
or U4228 (N_4228,N_3836,N_3770);
and U4229 (N_4229,N_3870,N_3993);
nor U4230 (N_4230,N_3901,N_3756);
nor U4231 (N_4231,N_3773,N_3927);
or U4232 (N_4232,N_3941,N_3830);
xnor U4233 (N_4233,N_3767,N_3823);
xor U4234 (N_4234,N_3835,N_3924);
xnor U4235 (N_4235,N_3966,N_3762);
or U4236 (N_4236,N_3888,N_3908);
or U4237 (N_4237,N_3816,N_3843);
xnor U4238 (N_4238,N_3947,N_3831);
and U4239 (N_4239,N_3870,N_3896);
and U4240 (N_4240,N_3866,N_3841);
xor U4241 (N_4241,N_3959,N_3904);
or U4242 (N_4242,N_3934,N_3754);
and U4243 (N_4243,N_3806,N_3932);
xor U4244 (N_4244,N_3789,N_3956);
nand U4245 (N_4245,N_3754,N_3799);
or U4246 (N_4246,N_3970,N_3833);
nand U4247 (N_4247,N_3858,N_3933);
nand U4248 (N_4248,N_3954,N_3906);
or U4249 (N_4249,N_3973,N_3867);
and U4250 (N_4250,N_4029,N_4171);
and U4251 (N_4251,N_4182,N_4013);
nand U4252 (N_4252,N_4205,N_4112);
nand U4253 (N_4253,N_4093,N_4069);
nor U4254 (N_4254,N_4183,N_4044);
xor U4255 (N_4255,N_4051,N_4030);
nand U4256 (N_4256,N_4097,N_4215);
nand U4257 (N_4257,N_4165,N_4164);
and U4258 (N_4258,N_4054,N_4047);
or U4259 (N_4259,N_4218,N_4065);
xnor U4260 (N_4260,N_4192,N_4039);
xor U4261 (N_4261,N_4149,N_4007);
nor U4262 (N_4262,N_4163,N_4041);
nor U4263 (N_4263,N_4141,N_4177);
nor U4264 (N_4264,N_4080,N_4036);
xor U4265 (N_4265,N_4076,N_4175);
and U4266 (N_4266,N_4060,N_4020);
nor U4267 (N_4267,N_4114,N_4142);
and U4268 (N_4268,N_4168,N_4106);
xor U4269 (N_4269,N_4246,N_4074);
and U4270 (N_4270,N_4101,N_4116);
nand U4271 (N_4271,N_4123,N_4179);
nor U4272 (N_4272,N_4066,N_4063);
xnor U4273 (N_4273,N_4187,N_4092);
nand U4274 (N_4274,N_4237,N_4212);
or U4275 (N_4275,N_4008,N_4033);
nor U4276 (N_4276,N_4048,N_4005);
or U4277 (N_4277,N_4002,N_4023);
and U4278 (N_4278,N_4085,N_4242);
or U4279 (N_4279,N_4202,N_4089);
nand U4280 (N_4280,N_4040,N_4216);
or U4281 (N_4281,N_4102,N_4227);
nor U4282 (N_4282,N_4104,N_4245);
xnor U4283 (N_4283,N_4011,N_4127);
nand U4284 (N_4284,N_4121,N_4238);
xnor U4285 (N_4285,N_4028,N_4228);
nor U4286 (N_4286,N_4072,N_4208);
nand U4287 (N_4287,N_4026,N_4160);
nand U4288 (N_4288,N_4045,N_4061);
nor U4289 (N_4289,N_4022,N_4151);
xnor U4290 (N_4290,N_4220,N_4012);
and U4291 (N_4291,N_4197,N_4191);
or U4292 (N_4292,N_4094,N_4010);
xor U4293 (N_4293,N_4108,N_4064);
nor U4294 (N_4294,N_4118,N_4230);
nand U4295 (N_4295,N_4198,N_4009);
and U4296 (N_4296,N_4157,N_4052);
nor U4297 (N_4297,N_4243,N_4152);
nand U4298 (N_4298,N_4035,N_4158);
and U4299 (N_4299,N_4196,N_4099);
xnor U4300 (N_4300,N_4082,N_4224);
xnor U4301 (N_4301,N_4204,N_4049);
and U4302 (N_4302,N_4236,N_4043);
nor U4303 (N_4303,N_4225,N_4136);
xnor U4304 (N_4304,N_4219,N_4146);
xor U4305 (N_4305,N_4037,N_4103);
and U4306 (N_4306,N_4098,N_4100);
or U4307 (N_4307,N_4122,N_4113);
nand U4308 (N_4308,N_4095,N_4172);
nor U4309 (N_4309,N_4249,N_4042);
and U4310 (N_4310,N_4184,N_4129);
nor U4311 (N_4311,N_4148,N_4021);
nand U4312 (N_4312,N_4024,N_4159);
and U4313 (N_4313,N_4025,N_4071);
and U4314 (N_4314,N_4223,N_4248);
and U4315 (N_4315,N_4234,N_4133);
or U4316 (N_4316,N_4046,N_4214);
xnor U4317 (N_4317,N_4203,N_4147);
and U4318 (N_4318,N_4073,N_4130);
and U4319 (N_4319,N_4155,N_4156);
and U4320 (N_4320,N_4200,N_4153);
xnor U4321 (N_4321,N_4201,N_4078);
and U4322 (N_4322,N_4233,N_4015);
nor U4323 (N_4323,N_4195,N_4077);
nand U4324 (N_4324,N_4109,N_4124);
xor U4325 (N_4325,N_4018,N_4140);
xor U4326 (N_4326,N_4014,N_4126);
nand U4327 (N_4327,N_4134,N_4154);
xor U4328 (N_4328,N_4091,N_4190);
nor U4329 (N_4329,N_4161,N_4067);
nand U4330 (N_4330,N_4027,N_4016);
nor U4331 (N_4331,N_4240,N_4199);
nand U4332 (N_4332,N_4128,N_4235);
nand U4333 (N_4333,N_4070,N_4226);
or U4334 (N_4334,N_4173,N_4017);
or U4335 (N_4335,N_4081,N_4139);
and U4336 (N_4336,N_4001,N_4117);
nand U4337 (N_4337,N_4062,N_4229);
and U4338 (N_4338,N_4084,N_4111);
and U4339 (N_4339,N_4181,N_4170);
and U4340 (N_4340,N_4217,N_4207);
and U4341 (N_4341,N_4194,N_4150);
nand U4342 (N_4342,N_4239,N_4188);
nand U4343 (N_4343,N_4038,N_4176);
and U4344 (N_4344,N_4119,N_4055);
or U4345 (N_4345,N_4137,N_4232);
nand U4346 (N_4346,N_4120,N_4135);
nand U4347 (N_4347,N_4090,N_4169);
xor U4348 (N_4348,N_4034,N_4096);
or U4349 (N_4349,N_4222,N_4138);
or U4350 (N_4350,N_4000,N_4075);
and U4351 (N_4351,N_4213,N_4209);
nand U4352 (N_4352,N_4162,N_4211);
or U4353 (N_4353,N_4244,N_4004);
nand U4354 (N_4354,N_4210,N_4167);
nand U4355 (N_4355,N_4068,N_4087);
xor U4356 (N_4356,N_4180,N_4186);
xnor U4357 (N_4357,N_4125,N_4110);
nand U4358 (N_4358,N_4132,N_4144);
xnor U4359 (N_4359,N_4185,N_4019);
nand U4360 (N_4360,N_4032,N_4143);
nor U4361 (N_4361,N_4107,N_4059);
nor U4362 (N_4362,N_4057,N_4231);
nor U4363 (N_4363,N_4174,N_4003);
xnor U4364 (N_4364,N_4166,N_4241);
xnor U4365 (N_4365,N_4105,N_4115);
and U4366 (N_4366,N_4056,N_4053);
nand U4367 (N_4367,N_4079,N_4221);
nor U4368 (N_4368,N_4058,N_4050);
or U4369 (N_4369,N_4145,N_4088);
and U4370 (N_4370,N_4131,N_4086);
and U4371 (N_4371,N_4206,N_4083);
nand U4372 (N_4372,N_4006,N_4031);
and U4373 (N_4373,N_4189,N_4178);
and U4374 (N_4374,N_4193,N_4247);
nor U4375 (N_4375,N_4172,N_4064);
nand U4376 (N_4376,N_4196,N_4172);
or U4377 (N_4377,N_4156,N_4174);
nand U4378 (N_4378,N_4235,N_4073);
xnor U4379 (N_4379,N_4184,N_4036);
xor U4380 (N_4380,N_4222,N_4001);
nand U4381 (N_4381,N_4001,N_4150);
nor U4382 (N_4382,N_4128,N_4012);
and U4383 (N_4383,N_4032,N_4204);
xor U4384 (N_4384,N_4210,N_4196);
or U4385 (N_4385,N_4149,N_4117);
nor U4386 (N_4386,N_4190,N_4089);
nand U4387 (N_4387,N_4037,N_4102);
nand U4388 (N_4388,N_4001,N_4032);
nand U4389 (N_4389,N_4136,N_4189);
nor U4390 (N_4390,N_4036,N_4106);
xor U4391 (N_4391,N_4225,N_4082);
xor U4392 (N_4392,N_4220,N_4112);
xor U4393 (N_4393,N_4243,N_4015);
and U4394 (N_4394,N_4209,N_4050);
nand U4395 (N_4395,N_4194,N_4042);
nand U4396 (N_4396,N_4141,N_4111);
nand U4397 (N_4397,N_4125,N_4034);
or U4398 (N_4398,N_4030,N_4017);
xor U4399 (N_4399,N_4239,N_4052);
nor U4400 (N_4400,N_4077,N_4011);
nor U4401 (N_4401,N_4117,N_4182);
xnor U4402 (N_4402,N_4227,N_4057);
xor U4403 (N_4403,N_4189,N_4155);
nor U4404 (N_4404,N_4015,N_4161);
or U4405 (N_4405,N_4032,N_4172);
xnor U4406 (N_4406,N_4029,N_4160);
nor U4407 (N_4407,N_4007,N_4152);
nand U4408 (N_4408,N_4142,N_4178);
xnor U4409 (N_4409,N_4062,N_4171);
xnor U4410 (N_4410,N_4104,N_4078);
or U4411 (N_4411,N_4153,N_4168);
or U4412 (N_4412,N_4173,N_4057);
xor U4413 (N_4413,N_4166,N_4190);
or U4414 (N_4414,N_4007,N_4071);
nand U4415 (N_4415,N_4021,N_4079);
nand U4416 (N_4416,N_4173,N_4113);
or U4417 (N_4417,N_4041,N_4074);
xnor U4418 (N_4418,N_4211,N_4116);
xnor U4419 (N_4419,N_4107,N_4113);
or U4420 (N_4420,N_4042,N_4040);
and U4421 (N_4421,N_4105,N_4031);
xor U4422 (N_4422,N_4211,N_4017);
and U4423 (N_4423,N_4188,N_4216);
nor U4424 (N_4424,N_4041,N_4026);
or U4425 (N_4425,N_4129,N_4108);
and U4426 (N_4426,N_4098,N_4215);
nand U4427 (N_4427,N_4125,N_4016);
xnor U4428 (N_4428,N_4029,N_4138);
nor U4429 (N_4429,N_4078,N_4028);
and U4430 (N_4430,N_4003,N_4033);
nand U4431 (N_4431,N_4174,N_4005);
or U4432 (N_4432,N_4201,N_4138);
nor U4433 (N_4433,N_4016,N_4232);
or U4434 (N_4434,N_4249,N_4079);
nand U4435 (N_4435,N_4031,N_4088);
nor U4436 (N_4436,N_4204,N_4109);
nand U4437 (N_4437,N_4136,N_4173);
or U4438 (N_4438,N_4122,N_4173);
nand U4439 (N_4439,N_4009,N_4238);
and U4440 (N_4440,N_4097,N_4180);
and U4441 (N_4441,N_4049,N_4081);
and U4442 (N_4442,N_4226,N_4035);
nand U4443 (N_4443,N_4015,N_4206);
and U4444 (N_4444,N_4247,N_4121);
xnor U4445 (N_4445,N_4218,N_4007);
nor U4446 (N_4446,N_4164,N_4073);
nor U4447 (N_4447,N_4159,N_4027);
nand U4448 (N_4448,N_4145,N_4244);
and U4449 (N_4449,N_4052,N_4023);
nor U4450 (N_4450,N_4202,N_4172);
and U4451 (N_4451,N_4203,N_4180);
nor U4452 (N_4452,N_4084,N_4144);
xor U4453 (N_4453,N_4201,N_4008);
nand U4454 (N_4454,N_4059,N_4062);
xor U4455 (N_4455,N_4017,N_4235);
nand U4456 (N_4456,N_4033,N_4020);
or U4457 (N_4457,N_4102,N_4229);
nor U4458 (N_4458,N_4237,N_4127);
nor U4459 (N_4459,N_4059,N_4200);
nor U4460 (N_4460,N_4023,N_4009);
nor U4461 (N_4461,N_4151,N_4190);
or U4462 (N_4462,N_4228,N_4227);
and U4463 (N_4463,N_4019,N_4027);
or U4464 (N_4464,N_4220,N_4046);
or U4465 (N_4465,N_4054,N_4246);
nand U4466 (N_4466,N_4093,N_4013);
or U4467 (N_4467,N_4093,N_4230);
or U4468 (N_4468,N_4131,N_4016);
or U4469 (N_4469,N_4055,N_4050);
nor U4470 (N_4470,N_4177,N_4237);
nor U4471 (N_4471,N_4190,N_4239);
and U4472 (N_4472,N_4125,N_4073);
nand U4473 (N_4473,N_4020,N_4051);
xor U4474 (N_4474,N_4152,N_4113);
or U4475 (N_4475,N_4031,N_4171);
or U4476 (N_4476,N_4153,N_4148);
xor U4477 (N_4477,N_4127,N_4166);
nand U4478 (N_4478,N_4192,N_4146);
or U4479 (N_4479,N_4059,N_4070);
and U4480 (N_4480,N_4102,N_4015);
nor U4481 (N_4481,N_4127,N_4202);
nor U4482 (N_4482,N_4035,N_4131);
and U4483 (N_4483,N_4100,N_4188);
xor U4484 (N_4484,N_4055,N_4195);
nor U4485 (N_4485,N_4095,N_4222);
nor U4486 (N_4486,N_4127,N_4080);
nand U4487 (N_4487,N_4154,N_4048);
xnor U4488 (N_4488,N_4147,N_4172);
and U4489 (N_4489,N_4155,N_4136);
or U4490 (N_4490,N_4186,N_4230);
nor U4491 (N_4491,N_4245,N_4108);
xnor U4492 (N_4492,N_4098,N_4009);
and U4493 (N_4493,N_4053,N_4062);
and U4494 (N_4494,N_4207,N_4146);
or U4495 (N_4495,N_4162,N_4181);
nor U4496 (N_4496,N_4083,N_4224);
nand U4497 (N_4497,N_4038,N_4234);
and U4498 (N_4498,N_4029,N_4187);
nand U4499 (N_4499,N_4020,N_4086);
nor U4500 (N_4500,N_4266,N_4436);
or U4501 (N_4501,N_4471,N_4472);
or U4502 (N_4502,N_4394,N_4467);
nor U4503 (N_4503,N_4435,N_4364);
nand U4504 (N_4504,N_4265,N_4418);
nand U4505 (N_4505,N_4430,N_4365);
or U4506 (N_4506,N_4348,N_4315);
or U4507 (N_4507,N_4333,N_4360);
nor U4508 (N_4508,N_4465,N_4367);
and U4509 (N_4509,N_4393,N_4357);
nand U4510 (N_4510,N_4494,N_4496);
and U4511 (N_4511,N_4489,N_4449);
xor U4512 (N_4512,N_4480,N_4354);
nand U4513 (N_4513,N_4381,N_4481);
nand U4514 (N_4514,N_4391,N_4451);
nand U4515 (N_4515,N_4409,N_4476);
xor U4516 (N_4516,N_4323,N_4390);
nand U4517 (N_4517,N_4344,N_4400);
and U4518 (N_4518,N_4456,N_4340);
and U4519 (N_4519,N_4466,N_4299);
and U4520 (N_4520,N_4379,N_4253);
and U4521 (N_4521,N_4416,N_4268);
nor U4522 (N_4522,N_4450,N_4258);
nand U4523 (N_4523,N_4421,N_4305);
xnor U4524 (N_4524,N_4358,N_4377);
nor U4525 (N_4525,N_4342,N_4298);
nand U4526 (N_4526,N_4478,N_4479);
or U4527 (N_4527,N_4290,N_4458);
or U4528 (N_4528,N_4314,N_4433);
or U4529 (N_4529,N_4386,N_4495);
and U4530 (N_4530,N_4325,N_4288);
nor U4531 (N_4531,N_4291,N_4294);
xnor U4532 (N_4532,N_4426,N_4468);
nand U4533 (N_4533,N_4341,N_4279);
nand U4534 (N_4534,N_4427,N_4351);
and U4535 (N_4535,N_4371,N_4275);
or U4536 (N_4536,N_4499,N_4252);
nand U4537 (N_4537,N_4398,N_4303);
nor U4538 (N_4538,N_4281,N_4260);
nand U4539 (N_4539,N_4399,N_4493);
xnor U4540 (N_4540,N_4318,N_4332);
and U4541 (N_4541,N_4470,N_4292);
xnor U4542 (N_4542,N_4378,N_4259);
nor U4543 (N_4543,N_4272,N_4267);
and U4544 (N_4544,N_4492,N_4317);
xnor U4545 (N_4545,N_4335,N_4473);
nor U4546 (N_4546,N_4361,N_4431);
and U4547 (N_4547,N_4251,N_4331);
or U4548 (N_4548,N_4289,N_4432);
or U4549 (N_4549,N_4347,N_4469);
nand U4550 (N_4550,N_4271,N_4355);
xor U4551 (N_4551,N_4283,N_4475);
nand U4552 (N_4552,N_4376,N_4284);
and U4553 (N_4553,N_4413,N_4406);
xnor U4554 (N_4554,N_4363,N_4353);
and U4555 (N_4555,N_4422,N_4420);
nor U4556 (N_4556,N_4385,N_4359);
nor U4557 (N_4557,N_4308,N_4444);
nor U4558 (N_4558,N_4311,N_4424);
and U4559 (N_4559,N_4488,N_4405);
or U4560 (N_4560,N_4263,N_4309);
xor U4561 (N_4561,N_4368,N_4300);
xnor U4562 (N_4562,N_4445,N_4321);
and U4563 (N_4563,N_4434,N_4293);
nor U4564 (N_4564,N_4329,N_4285);
nor U4565 (N_4565,N_4350,N_4396);
and U4566 (N_4566,N_4278,N_4428);
nor U4567 (N_4567,N_4383,N_4440);
and U4568 (N_4568,N_4395,N_4255);
nand U4569 (N_4569,N_4446,N_4425);
or U4570 (N_4570,N_4498,N_4256);
nor U4571 (N_4571,N_4486,N_4336);
and U4572 (N_4572,N_4261,N_4487);
xnor U4573 (N_4573,N_4339,N_4372);
or U4574 (N_4574,N_4274,N_4410);
nor U4575 (N_4575,N_4464,N_4397);
or U4576 (N_4576,N_4273,N_4483);
nor U4577 (N_4577,N_4438,N_4334);
nand U4578 (N_4578,N_4454,N_4264);
nand U4579 (N_4579,N_4280,N_4384);
nor U4580 (N_4580,N_4388,N_4356);
or U4581 (N_4581,N_4419,N_4286);
xnor U4582 (N_4582,N_4338,N_4287);
nand U4583 (N_4583,N_4370,N_4277);
nor U4584 (N_4584,N_4262,N_4459);
nor U4585 (N_4585,N_4455,N_4448);
or U4586 (N_4586,N_4306,N_4382);
nor U4587 (N_4587,N_4457,N_4257);
nand U4588 (N_4588,N_4327,N_4282);
nor U4589 (N_4589,N_4328,N_4407);
and U4590 (N_4590,N_4460,N_4412);
nand U4591 (N_4591,N_4316,N_4414);
nor U4592 (N_4592,N_4392,N_4441);
or U4593 (N_4593,N_4408,N_4429);
nand U4594 (N_4594,N_4304,N_4463);
xnor U4595 (N_4595,N_4346,N_4415);
or U4596 (N_4596,N_4490,N_4362);
and U4597 (N_4597,N_4373,N_4319);
nor U4598 (N_4598,N_4337,N_4343);
nor U4599 (N_4599,N_4442,N_4374);
xor U4600 (N_4600,N_4387,N_4403);
nand U4601 (N_4601,N_4302,N_4254);
nor U4602 (N_4602,N_4404,N_4402);
nor U4603 (N_4603,N_4296,N_4295);
nor U4604 (N_4604,N_4276,N_4375);
or U4605 (N_4605,N_4447,N_4411);
nor U4606 (N_4606,N_4330,N_4369);
nand U4607 (N_4607,N_4452,N_4380);
nand U4608 (N_4608,N_4491,N_4482);
or U4609 (N_4609,N_4497,N_4443);
nand U4610 (N_4610,N_4474,N_4401);
nor U4611 (N_4611,N_4345,N_4439);
and U4612 (N_4612,N_4324,N_4461);
and U4613 (N_4613,N_4301,N_4437);
and U4614 (N_4614,N_4366,N_4423);
nor U4615 (N_4615,N_4349,N_4297);
nor U4616 (N_4616,N_4485,N_4312);
nand U4617 (N_4617,N_4352,N_4310);
or U4618 (N_4618,N_4389,N_4477);
nand U4619 (N_4619,N_4270,N_4307);
nor U4620 (N_4620,N_4484,N_4320);
and U4621 (N_4621,N_4326,N_4453);
nor U4622 (N_4622,N_4462,N_4250);
xnor U4623 (N_4623,N_4313,N_4417);
nand U4624 (N_4624,N_4322,N_4269);
nand U4625 (N_4625,N_4368,N_4259);
xor U4626 (N_4626,N_4336,N_4497);
nor U4627 (N_4627,N_4385,N_4419);
xor U4628 (N_4628,N_4363,N_4343);
or U4629 (N_4629,N_4318,N_4461);
and U4630 (N_4630,N_4390,N_4421);
or U4631 (N_4631,N_4324,N_4287);
and U4632 (N_4632,N_4255,N_4450);
xnor U4633 (N_4633,N_4263,N_4350);
nand U4634 (N_4634,N_4445,N_4298);
xor U4635 (N_4635,N_4411,N_4423);
nand U4636 (N_4636,N_4399,N_4416);
nor U4637 (N_4637,N_4255,N_4455);
nor U4638 (N_4638,N_4368,N_4377);
nor U4639 (N_4639,N_4294,N_4267);
nor U4640 (N_4640,N_4449,N_4461);
nor U4641 (N_4641,N_4280,N_4432);
or U4642 (N_4642,N_4393,N_4333);
or U4643 (N_4643,N_4490,N_4341);
nand U4644 (N_4644,N_4250,N_4422);
nand U4645 (N_4645,N_4441,N_4389);
nand U4646 (N_4646,N_4310,N_4382);
xnor U4647 (N_4647,N_4431,N_4476);
or U4648 (N_4648,N_4351,N_4480);
xor U4649 (N_4649,N_4437,N_4477);
and U4650 (N_4650,N_4495,N_4396);
and U4651 (N_4651,N_4314,N_4327);
nor U4652 (N_4652,N_4368,N_4402);
xor U4653 (N_4653,N_4454,N_4322);
nor U4654 (N_4654,N_4250,N_4257);
nor U4655 (N_4655,N_4496,N_4351);
nor U4656 (N_4656,N_4302,N_4384);
or U4657 (N_4657,N_4312,N_4319);
xnor U4658 (N_4658,N_4483,N_4385);
xor U4659 (N_4659,N_4276,N_4395);
nand U4660 (N_4660,N_4463,N_4474);
or U4661 (N_4661,N_4379,N_4394);
nor U4662 (N_4662,N_4432,N_4255);
or U4663 (N_4663,N_4357,N_4460);
xor U4664 (N_4664,N_4367,N_4461);
nor U4665 (N_4665,N_4487,N_4401);
or U4666 (N_4666,N_4369,N_4355);
nand U4667 (N_4667,N_4320,N_4497);
xor U4668 (N_4668,N_4432,N_4332);
xor U4669 (N_4669,N_4297,N_4324);
nand U4670 (N_4670,N_4328,N_4263);
xnor U4671 (N_4671,N_4431,N_4274);
xnor U4672 (N_4672,N_4498,N_4481);
xor U4673 (N_4673,N_4418,N_4398);
and U4674 (N_4674,N_4372,N_4380);
xnor U4675 (N_4675,N_4299,N_4353);
and U4676 (N_4676,N_4262,N_4250);
nor U4677 (N_4677,N_4341,N_4329);
or U4678 (N_4678,N_4456,N_4401);
nand U4679 (N_4679,N_4456,N_4270);
nor U4680 (N_4680,N_4350,N_4335);
nor U4681 (N_4681,N_4300,N_4464);
and U4682 (N_4682,N_4475,N_4420);
xor U4683 (N_4683,N_4303,N_4479);
xnor U4684 (N_4684,N_4372,N_4325);
or U4685 (N_4685,N_4477,N_4270);
or U4686 (N_4686,N_4291,N_4273);
or U4687 (N_4687,N_4404,N_4414);
nor U4688 (N_4688,N_4487,N_4288);
nor U4689 (N_4689,N_4263,N_4452);
or U4690 (N_4690,N_4423,N_4461);
nor U4691 (N_4691,N_4444,N_4477);
nor U4692 (N_4692,N_4486,N_4329);
nand U4693 (N_4693,N_4345,N_4384);
or U4694 (N_4694,N_4369,N_4442);
xor U4695 (N_4695,N_4421,N_4324);
nand U4696 (N_4696,N_4329,N_4357);
nand U4697 (N_4697,N_4489,N_4428);
or U4698 (N_4698,N_4409,N_4267);
or U4699 (N_4699,N_4328,N_4271);
and U4700 (N_4700,N_4286,N_4342);
or U4701 (N_4701,N_4255,N_4302);
nand U4702 (N_4702,N_4369,N_4441);
or U4703 (N_4703,N_4450,N_4366);
nand U4704 (N_4704,N_4301,N_4270);
and U4705 (N_4705,N_4453,N_4304);
xor U4706 (N_4706,N_4259,N_4467);
nor U4707 (N_4707,N_4424,N_4388);
nor U4708 (N_4708,N_4405,N_4384);
nor U4709 (N_4709,N_4459,N_4406);
nor U4710 (N_4710,N_4484,N_4352);
nor U4711 (N_4711,N_4274,N_4293);
nand U4712 (N_4712,N_4261,N_4338);
or U4713 (N_4713,N_4278,N_4291);
or U4714 (N_4714,N_4264,N_4493);
xor U4715 (N_4715,N_4381,N_4259);
and U4716 (N_4716,N_4351,N_4295);
and U4717 (N_4717,N_4344,N_4353);
nor U4718 (N_4718,N_4349,N_4370);
nand U4719 (N_4719,N_4255,N_4277);
nand U4720 (N_4720,N_4440,N_4290);
and U4721 (N_4721,N_4436,N_4437);
xnor U4722 (N_4722,N_4419,N_4401);
xor U4723 (N_4723,N_4379,N_4356);
nor U4724 (N_4724,N_4395,N_4250);
or U4725 (N_4725,N_4445,N_4489);
nor U4726 (N_4726,N_4296,N_4254);
nor U4727 (N_4727,N_4489,N_4396);
xnor U4728 (N_4728,N_4316,N_4346);
or U4729 (N_4729,N_4333,N_4370);
and U4730 (N_4730,N_4429,N_4385);
nand U4731 (N_4731,N_4264,N_4351);
nand U4732 (N_4732,N_4368,N_4253);
and U4733 (N_4733,N_4404,N_4334);
xnor U4734 (N_4734,N_4282,N_4361);
xnor U4735 (N_4735,N_4365,N_4341);
or U4736 (N_4736,N_4456,N_4495);
and U4737 (N_4737,N_4259,N_4476);
nand U4738 (N_4738,N_4309,N_4463);
xnor U4739 (N_4739,N_4300,N_4374);
nor U4740 (N_4740,N_4392,N_4474);
nand U4741 (N_4741,N_4337,N_4493);
or U4742 (N_4742,N_4332,N_4427);
or U4743 (N_4743,N_4436,N_4410);
or U4744 (N_4744,N_4340,N_4294);
nand U4745 (N_4745,N_4375,N_4433);
nor U4746 (N_4746,N_4292,N_4457);
nand U4747 (N_4747,N_4339,N_4411);
and U4748 (N_4748,N_4408,N_4377);
xor U4749 (N_4749,N_4367,N_4455);
or U4750 (N_4750,N_4621,N_4716);
or U4751 (N_4751,N_4518,N_4539);
and U4752 (N_4752,N_4597,N_4623);
nand U4753 (N_4753,N_4710,N_4672);
xor U4754 (N_4754,N_4543,N_4662);
and U4755 (N_4755,N_4692,N_4719);
nor U4756 (N_4756,N_4501,N_4584);
nand U4757 (N_4757,N_4661,N_4536);
xor U4758 (N_4758,N_4631,N_4547);
nor U4759 (N_4759,N_4728,N_4559);
xnor U4760 (N_4760,N_4553,N_4691);
or U4761 (N_4761,N_4571,N_4657);
nand U4762 (N_4762,N_4668,N_4713);
nand U4763 (N_4763,N_4565,N_4743);
or U4764 (N_4764,N_4731,N_4554);
or U4765 (N_4765,N_4715,N_4614);
and U4766 (N_4766,N_4737,N_4694);
and U4767 (N_4767,N_4511,N_4525);
xnor U4768 (N_4768,N_4749,N_4526);
nor U4769 (N_4769,N_4522,N_4706);
xor U4770 (N_4770,N_4517,N_4537);
nand U4771 (N_4771,N_4609,N_4549);
xor U4772 (N_4772,N_4697,N_4587);
xor U4773 (N_4773,N_4722,N_4588);
or U4774 (N_4774,N_4541,N_4574);
xor U4775 (N_4775,N_4508,N_4738);
nor U4776 (N_4776,N_4652,N_4600);
nand U4777 (N_4777,N_4717,N_4580);
nand U4778 (N_4778,N_4665,N_4681);
xnor U4779 (N_4779,N_4618,N_4573);
xnor U4780 (N_4780,N_4538,N_4700);
or U4781 (N_4781,N_4509,N_4646);
nor U4782 (N_4782,N_4653,N_4626);
nand U4783 (N_4783,N_4564,N_4688);
xor U4784 (N_4784,N_4568,N_4695);
nand U4785 (N_4785,N_4569,N_4707);
and U4786 (N_4786,N_4744,N_4578);
nand U4787 (N_4787,N_4582,N_4682);
xor U4788 (N_4788,N_4595,N_4612);
nand U4789 (N_4789,N_4581,N_4643);
nand U4790 (N_4790,N_4718,N_4669);
or U4791 (N_4791,N_4545,N_4555);
nor U4792 (N_4792,N_4640,N_4671);
nor U4793 (N_4793,N_4660,N_4528);
nor U4794 (N_4794,N_4693,N_4673);
nand U4795 (N_4795,N_4616,N_4577);
and U4796 (N_4796,N_4736,N_4685);
or U4797 (N_4797,N_4664,N_4603);
or U4798 (N_4798,N_4520,N_4666);
nand U4799 (N_4799,N_4644,N_4632);
nor U4800 (N_4800,N_4519,N_4594);
nor U4801 (N_4801,N_4670,N_4516);
nand U4802 (N_4802,N_4534,N_4727);
nor U4803 (N_4803,N_4610,N_4607);
nor U4804 (N_4804,N_4579,N_4570);
and U4805 (N_4805,N_4699,N_4724);
or U4806 (N_4806,N_4689,N_4637);
nor U4807 (N_4807,N_4676,N_4596);
nand U4808 (N_4808,N_4510,N_4655);
or U4809 (N_4809,N_4524,N_4502);
and U4810 (N_4810,N_4723,N_4659);
nand U4811 (N_4811,N_4720,N_4566);
nand U4812 (N_4812,N_4512,N_4567);
or U4813 (N_4813,N_4633,N_4507);
nand U4814 (N_4814,N_4506,N_4561);
nor U4815 (N_4815,N_4608,N_4550);
nand U4816 (N_4816,N_4540,N_4739);
nand U4817 (N_4817,N_4615,N_4601);
nand U4818 (N_4818,N_4557,N_4617);
nand U4819 (N_4819,N_4648,N_4514);
nand U4820 (N_4820,N_4642,N_4711);
and U4821 (N_4821,N_4551,N_4624);
and U4822 (N_4822,N_4732,N_4714);
or U4823 (N_4823,N_4687,N_4535);
or U4824 (N_4824,N_4638,N_4674);
xor U4825 (N_4825,N_4730,N_4544);
and U4826 (N_4826,N_4622,N_4599);
nand U4827 (N_4827,N_4639,N_4542);
nor U4828 (N_4828,N_4500,N_4531);
xor U4829 (N_4829,N_4556,N_4740);
nor U4830 (N_4830,N_4705,N_4513);
nor U4831 (N_4831,N_4735,N_4663);
nor U4832 (N_4832,N_4680,N_4654);
xnor U4833 (N_4833,N_4503,N_4683);
xnor U4834 (N_4834,N_4703,N_4729);
nor U4835 (N_4835,N_4641,N_4649);
nand U4836 (N_4836,N_4630,N_4529);
nand U4837 (N_4837,N_4678,N_4560);
nor U4838 (N_4838,N_4726,N_4656);
xnor U4839 (N_4839,N_4575,N_4734);
xnor U4840 (N_4840,N_4747,N_4667);
xor U4841 (N_4841,N_4576,N_4712);
nand U4842 (N_4842,N_4651,N_4530);
nor U4843 (N_4843,N_4690,N_4704);
nand U4844 (N_4844,N_4527,N_4546);
nand U4845 (N_4845,N_4558,N_4611);
nor U4846 (N_4846,N_4548,N_4505);
xnor U4847 (N_4847,N_4698,N_4515);
or U4848 (N_4848,N_4620,N_4625);
or U4849 (N_4849,N_4708,N_4628);
and U4850 (N_4850,N_4591,N_4590);
xor U4851 (N_4851,N_4701,N_4619);
nor U4852 (N_4852,N_4725,N_4650);
nand U4853 (N_4853,N_4746,N_4658);
xor U4854 (N_4854,N_4742,N_4585);
xnor U4855 (N_4855,N_4605,N_4586);
nor U4856 (N_4856,N_4702,N_4589);
nand U4857 (N_4857,N_4709,N_4613);
and U4858 (N_4858,N_4748,N_4686);
and U4859 (N_4859,N_4721,N_4733);
nand U4860 (N_4860,N_4745,N_4606);
nor U4861 (N_4861,N_4629,N_4593);
nand U4862 (N_4862,N_4675,N_4552);
nor U4863 (N_4863,N_4602,N_4521);
xnor U4864 (N_4864,N_4572,N_4679);
or U4865 (N_4865,N_4627,N_4533);
and U4866 (N_4866,N_4523,N_4598);
nor U4867 (N_4867,N_4583,N_4504);
nor U4868 (N_4868,N_4677,N_4604);
and U4869 (N_4869,N_4647,N_4634);
or U4870 (N_4870,N_4741,N_4532);
nor U4871 (N_4871,N_4684,N_4592);
nor U4872 (N_4872,N_4563,N_4645);
and U4873 (N_4873,N_4696,N_4636);
and U4874 (N_4874,N_4562,N_4635);
and U4875 (N_4875,N_4509,N_4614);
nor U4876 (N_4876,N_4710,N_4594);
nand U4877 (N_4877,N_4537,N_4570);
nor U4878 (N_4878,N_4714,N_4592);
and U4879 (N_4879,N_4595,N_4637);
or U4880 (N_4880,N_4628,N_4706);
and U4881 (N_4881,N_4506,N_4673);
and U4882 (N_4882,N_4530,N_4596);
nand U4883 (N_4883,N_4646,N_4638);
and U4884 (N_4884,N_4605,N_4525);
nor U4885 (N_4885,N_4738,N_4727);
xor U4886 (N_4886,N_4598,N_4710);
nor U4887 (N_4887,N_4643,N_4603);
or U4888 (N_4888,N_4686,N_4500);
nor U4889 (N_4889,N_4686,N_4664);
nor U4890 (N_4890,N_4615,N_4716);
nand U4891 (N_4891,N_4540,N_4621);
and U4892 (N_4892,N_4520,N_4544);
nor U4893 (N_4893,N_4657,N_4749);
nand U4894 (N_4894,N_4519,N_4622);
and U4895 (N_4895,N_4691,N_4665);
nor U4896 (N_4896,N_4560,N_4654);
or U4897 (N_4897,N_4721,N_4623);
nor U4898 (N_4898,N_4527,N_4519);
and U4899 (N_4899,N_4738,N_4643);
or U4900 (N_4900,N_4675,N_4561);
xnor U4901 (N_4901,N_4702,N_4646);
nor U4902 (N_4902,N_4712,N_4597);
and U4903 (N_4903,N_4594,N_4679);
or U4904 (N_4904,N_4640,N_4538);
xor U4905 (N_4905,N_4522,N_4634);
xor U4906 (N_4906,N_4546,N_4597);
or U4907 (N_4907,N_4629,N_4542);
nor U4908 (N_4908,N_4648,N_4737);
nor U4909 (N_4909,N_4643,N_4503);
nand U4910 (N_4910,N_4715,N_4733);
nand U4911 (N_4911,N_4641,N_4639);
or U4912 (N_4912,N_4562,N_4646);
xor U4913 (N_4913,N_4524,N_4676);
nand U4914 (N_4914,N_4549,N_4630);
xor U4915 (N_4915,N_4565,N_4598);
xnor U4916 (N_4916,N_4566,N_4685);
nor U4917 (N_4917,N_4745,N_4727);
or U4918 (N_4918,N_4600,N_4575);
or U4919 (N_4919,N_4610,N_4733);
nand U4920 (N_4920,N_4547,N_4676);
or U4921 (N_4921,N_4575,N_4504);
nand U4922 (N_4922,N_4565,N_4719);
and U4923 (N_4923,N_4719,N_4674);
and U4924 (N_4924,N_4576,N_4514);
or U4925 (N_4925,N_4728,N_4688);
or U4926 (N_4926,N_4647,N_4617);
nand U4927 (N_4927,N_4518,N_4610);
or U4928 (N_4928,N_4623,N_4595);
nor U4929 (N_4929,N_4642,N_4602);
nand U4930 (N_4930,N_4525,N_4696);
nand U4931 (N_4931,N_4586,N_4652);
xnor U4932 (N_4932,N_4673,N_4503);
xnor U4933 (N_4933,N_4607,N_4517);
xor U4934 (N_4934,N_4571,N_4559);
or U4935 (N_4935,N_4740,N_4637);
or U4936 (N_4936,N_4590,N_4674);
nor U4937 (N_4937,N_4625,N_4631);
or U4938 (N_4938,N_4561,N_4706);
nand U4939 (N_4939,N_4700,N_4520);
nand U4940 (N_4940,N_4639,N_4521);
and U4941 (N_4941,N_4671,N_4663);
or U4942 (N_4942,N_4558,N_4527);
or U4943 (N_4943,N_4718,N_4598);
xor U4944 (N_4944,N_4552,N_4614);
nand U4945 (N_4945,N_4709,N_4638);
or U4946 (N_4946,N_4514,N_4723);
and U4947 (N_4947,N_4652,N_4741);
nand U4948 (N_4948,N_4620,N_4636);
or U4949 (N_4949,N_4513,N_4700);
nor U4950 (N_4950,N_4660,N_4530);
nand U4951 (N_4951,N_4685,N_4608);
xnor U4952 (N_4952,N_4675,N_4725);
and U4953 (N_4953,N_4577,N_4622);
nand U4954 (N_4954,N_4739,N_4678);
nand U4955 (N_4955,N_4725,N_4646);
xnor U4956 (N_4956,N_4500,N_4549);
and U4957 (N_4957,N_4533,N_4587);
nor U4958 (N_4958,N_4554,N_4738);
and U4959 (N_4959,N_4687,N_4506);
nand U4960 (N_4960,N_4557,N_4748);
nor U4961 (N_4961,N_4530,N_4732);
or U4962 (N_4962,N_4649,N_4711);
nor U4963 (N_4963,N_4550,N_4619);
nand U4964 (N_4964,N_4676,N_4543);
xnor U4965 (N_4965,N_4697,N_4624);
xor U4966 (N_4966,N_4626,N_4608);
and U4967 (N_4967,N_4599,N_4527);
nor U4968 (N_4968,N_4586,N_4518);
and U4969 (N_4969,N_4509,N_4713);
nand U4970 (N_4970,N_4677,N_4695);
nand U4971 (N_4971,N_4610,N_4550);
nand U4972 (N_4972,N_4588,N_4743);
or U4973 (N_4973,N_4580,N_4649);
nand U4974 (N_4974,N_4552,N_4632);
nor U4975 (N_4975,N_4660,N_4657);
nor U4976 (N_4976,N_4579,N_4608);
nand U4977 (N_4977,N_4556,N_4735);
xnor U4978 (N_4978,N_4558,N_4637);
nand U4979 (N_4979,N_4552,N_4661);
xnor U4980 (N_4980,N_4621,N_4650);
or U4981 (N_4981,N_4565,N_4583);
or U4982 (N_4982,N_4628,N_4570);
xor U4983 (N_4983,N_4742,N_4677);
and U4984 (N_4984,N_4699,N_4578);
nand U4985 (N_4985,N_4579,N_4741);
and U4986 (N_4986,N_4646,N_4533);
nor U4987 (N_4987,N_4581,N_4547);
nor U4988 (N_4988,N_4666,N_4716);
xor U4989 (N_4989,N_4536,N_4642);
nand U4990 (N_4990,N_4636,N_4741);
xnor U4991 (N_4991,N_4682,N_4510);
nor U4992 (N_4992,N_4605,N_4738);
nor U4993 (N_4993,N_4543,N_4726);
and U4994 (N_4994,N_4731,N_4676);
or U4995 (N_4995,N_4672,N_4525);
xor U4996 (N_4996,N_4593,N_4702);
or U4997 (N_4997,N_4717,N_4729);
xor U4998 (N_4998,N_4738,N_4525);
and U4999 (N_4999,N_4536,N_4526);
and U5000 (N_5000,N_4817,N_4880);
xnor U5001 (N_5001,N_4751,N_4933);
xor U5002 (N_5002,N_4779,N_4780);
or U5003 (N_5003,N_4801,N_4839);
xor U5004 (N_5004,N_4938,N_4912);
nand U5005 (N_5005,N_4988,N_4800);
nor U5006 (N_5006,N_4840,N_4853);
and U5007 (N_5007,N_4883,N_4825);
nand U5008 (N_5008,N_4943,N_4927);
xor U5009 (N_5009,N_4815,N_4872);
xnor U5010 (N_5010,N_4925,N_4902);
nand U5011 (N_5011,N_4919,N_4841);
or U5012 (N_5012,N_4967,N_4945);
nor U5013 (N_5013,N_4984,N_4935);
xor U5014 (N_5014,N_4858,N_4990);
or U5015 (N_5015,N_4862,N_4784);
xnor U5016 (N_5016,N_4949,N_4766);
nand U5017 (N_5017,N_4964,N_4906);
nand U5018 (N_5018,N_4859,N_4824);
or U5019 (N_5019,N_4907,N_4834);
and U5020 (N_5020,N_4983,N_4956);
nor U5021 (N_5021,N_4994,N_4857);
nand U5022 (N_5022,N_4823,N_4837);
nand U5023 (N_5023,N_4977,N_4928);
or U5024 (N_5024,N_4820,N_4891);
or U5025 (N_5025,N_4856,N_4794);
and U5026 (N_5026,N_4830,N_4863);
and U5027 (N_5027,N_4917,N_4997);
or U5028 (N_5028,N_4923,N_4962);
or U5029 (N_5029,N_4878,N_4781);
or U5030 (N_5030,N_4852,N_4886);
nand U5031 (N_5031,N_4952,N_4851);
xnor U5032 (N_5032,N_4898,N_4969);
nor U5033 (N_5033,N_4768,N_4798);
nor U5034 (N_5034,N_4896,N_4941);
and U5035 (N_5035,N_4770,N_4805);
nand U5036 (N_5036,N_4826,N_4996);
nand U5037 (N_5037,N_4885,N_4774);
xnor U5038 (N_5038,N_4844,N_4995);
and U5039 (N_5039,N_4796,N_4909);
xnor U5040 (N_5040,N_4987,N_4921);
nor U5041 (N_5041,N_4910,N_4913);
nand U5042 (N_5042,N_4847,N_4953);
nand U5043 (N_5043,N_4842,N_4756);
or U5044 (N_5044,N_4973,N_4978);
nor U5045 (N_5045,N_4937,N_4991);
and U5046 (N_5046,N_4802,N_4992);
xor U5047 (N_5047,N_4777,N_4764);
xnor U5048 (N_5048,N_4870,N_4760);
xor U5049 (N_5049,N_4963,N_4835);
nor U5050 (N_5050,N_4793,N_4980);
xnor U5051 (N_5051,N_4915,N_4845);
nand U5052 (N_5052,N_4772,N_4931);
nand U5053 (N_5053,N_4888,N_4934);
nor U5054 (N_5054,N_4785,N_4783);
or U5055 (N_5055,N_4797,N_4976);
nor U5056 (N_5056,N_4877,N_4959);
or U5057 (N_5057,N_4754,N_4954);
nand U5058 (N_5058,N_4812,N_4979);
nor U5059 (N_5059,N_4951,N_4790);
or U5060 (N_5060,N_4871,N_4866);
nand U5061 (N_5061,N_4924,N_4892);
nand U5062 (N_5062,N_4828,N_4982);
nand U5063 (N_5063,N_4899,N_4811);
nor U5064 (N_5064,N_4832,N_4993);
xor U5065 (N_5065,N_4998,N_4763);
nand U5066 (N_5066,N_4788,N_4874);
nor U5067 (N_5067,N_4769,N_4855);
and U5068 (N_5068,N_4860,N_4838);
and U5069 (N_5069,N_4897,N_4961);
or U5070 (N_5070,N_4890,N_4960);
xor U5071 (N_5071,N_4776,N_4771);
nor U5072 (N_5072,N_4922,N_4803);
xnor U5073 (N_5073,N_4827,N_4867);
and U5074 (N_5074,N_4821,N_4848);
or U5075 (N_5075,N_4761,N_4882);
and U5076 (N_5076,N_4836,N_4986);
xnor U5077 (N_5077,N_4948,N_4787);
nand U5078 (N_5078,N_4799,N_4914);
and U5079 (N_5079,N_4905,N_4822);
nor U5080 (N_5080,N_4753,N_4829);
or U5081 (N_5081,N_4804,N_4939);
xor U5082 (N_5082,N_4791,N_4894);
or U5083 (N_5083,N_4846,N_4813);
or U5084 (N_5084,N_4895,N_4810);
xor U5085 (N_5085,N_4789,N_4775);
nand U5086 (N_5086,N_4833,N_4957);
nor U5087 (N_5087,N_4974,N_4970);
nand U5088 (N_5088,N_4981,N_4808);
and U5089 (N_5089,N_4965,N_4767);
and U5090 (N_5090,N_4792,N_4850);
or U5091 (N_5091,N_4989,N_4999);
xnor U5092 (N_5092,N_4819,N_4782);
nor U5093 (N_5093,N_4929,N_4889);
nand U5094 (N_5094,N_4750,N_4807);
nor U5095 (N_5095,N_4875,N_4975);
and U5096 (N_5096,N_4757,N_4849);
or U5097 (N_5097,N_4918,N_4814);
nor U5098 (N_5098,N_4958,N_4936);
or U5099 (N_5099,N_4985,N_4947);
nor U5100 (N_5100,N_4876,N_4904);
and U5101 (N_5101,N_4765,N_4762);
and U5102 (N_5102,N_4868,N_4786);
xnor U5103 (N_5103,N_4809,N_4893);
nor U5104 (N_5104,N_4887,N_4930);
and U5105 (N_5105,N_4944,N_4901);
or U5106 (N_5106,N_4865,N_4758);
nor U5107 (N_5107,N_4759,N_4903);
or U5108 (N_5108,N_4911,N_4778);
nand U5109 (N_5109,N_4752,N_4873);
xnor U5110 (N_5110,N_4773,N_4843);
and U5111 (N_5111,N_4955,N_4920);
nand U5112 (N_5112,N_4879,N_4816);
nor U5113 (N_5113,N_4806,N_4950);
xnor U5114 (N_5114,N_4966,N_4932);
xnor U5115 (N_5115,N_4946,N_4968);
xnor U5116 (N_5116,N_4972,N_4916);
nor U5117 (N_5117,N_4818,N_4831);
or U5118 (N_5118,N_4940,N_4861);
nor U5119 (N_5119,N_4854,N_4942);
and U5120 (N_5120,N_4908,N_4926);
nor U5121 (N_5121,N_4971,N_4869);
or U5122 (N_5122,N_4864,N_4900);
or U5123 (N_5123,N_4795,N_4755);
xnor U5124 (N_5124,N_4884,N_4881);
xor U5125 (N_5125,N_4854,N_4916);
and U5126 (N_5126,N_4825,N_4964);
nor U5127 (N_5127,N_4878,N_4826);
nor U5128 (N_5128,N_4764,N_4980);
nor U5129 (N_5129,N_4800,N_4920);
xor U5130 (N_5130,N_4752,N_4780);
and U5131 (N_5131,N_4833,N_4907);
nand U5132 (N_5132,N_4989,N_4796);
xor U5133 (N_5133,N_4876,N_4757);
xor U5134 (N_5134,N_4910,N_4911);
nand U5135 (N_5135,N_4895,N_4930);
or U5136 (N_5136,N_4883,N_4966);
nand U5137 (N_5137,N_4775,N_4955);
nand U5138 (N_5138,N_4832,N_4772);
xor U5139 (N_5139,N_4797,N_4917);
nand U5140 (N_5140,N_4994,N_4961);
or U5141 (N_5141,N_4936,N_4821);
and U5142 (N_5142,N_4878,N_4852);
xor U5143 (N_5143,N_4994,N_4850);
xor U5144 (N_5144,N_4870,N_4942);
or U5145 (N_5145,N_4918,N_4853);
or U5146 (N_5146,N_4821,N_4996);
or U5147 (N_5147,N_4990,N_4926);
or U5148 (N_5148,N_4841,N_4812);
xnor U5149 (N_5149,N_4948,N_4771);
nand U5150 (N_5150,N_4916,N_4981);
nor U5151 (N_5151,N_4852,N_4754);
nand U5152 (N_5152,N_4951,N_4800);
nor U5153 (N_5153,N_4789,N_4834);
or U5154 (N_5154,N_4920,N_4944);
xnor U5155 (N_5155,N_4957,N_4964);
nand U5156 (N_5156,N_4871,N_4863);
xor U5157 (N_5157,N_4881,N_4754);
nor U5158 (N_5158,N_4842,N_4826);
or U5159 (N_5159,N_4919,N_4907);
and U5160 (N_5160,N_4935,N_4847);
xor U5161 (N_5161,N_4931,N_4884);
nand U5162 (N_5162,N_4939,N_4922);
or U5163 (N_5163,N_4971,N_4871);
nand U5164 (N_5164,N_4822,N_4873);
xnor U5165 (N_5165,N_4760,N_4803);
nand U5166 (N_5166,N_4758,N_4798);
nand U5167 (N_5167,N_4796,N_4864);
xor U5168 (N_5168,N_4864,N_4848);
nor U5169 (N_5169,N_4819,N_4915);
and U5170 (N_5170,N_4888,N_4961);
nor U5171 (N_5171,N_4860,N_4873);
nand U5172 (N_5172,N_4824,N_4796);
nand U5173 (N_5173,N_4877,N_4776);
and U5174 (N_5174,N_4800,N_4971);
and U5175 (N_5175,N_4849,N_4884);
nor U5176 (N_5176,N_4879,N_4848);
or U5177 (N_5177,N_4794,N_4796);
nor U5178 (N_5178,N_4766,N_4898);
or U5179 (N_5179,N_4973,N_4967);
nor U5180 (N_5180,N_4861,N_4963);
and U5181 (N_5181,N_4807,N_4983);
xor U5182 (N_5182,N_4807,N_4814);
nor U5183 (N_5183,N_4917,N_4835);
nor U5184 (N_5184,N_4808,N_4937);
or U5185 (N_5185,N_4954,N_4854);
xnor U5186 (N_5186,N_4978,N_4844);
or U5187 (N_5187,N_4810,N_4848);
nor U5188 (N_5188,N_4945,N_4920);
nand U5189 (N_5189,N_4772,N_4816);
nor U5190 (N_5190,N_4959,N_4798);
and U5191 (N_5191,N_4863,N_4836);
or U5192 (N_5192,N_4772,N_4944);
nand U5193 (N_5193,N_4778,N_4866);
nand U5194 (N_5194,N_4891,N_4943);
xor U5195 (N_5195,N_4881,N_4785);
and U5196 (N_5196,N_4966,N_4886);
and U5197 (N_5197,N_4807,N_4808);
xnor U5198 (N_5198,N_4961,N_4989);
or U5199 (N_5199,N_4755,N_4826);
nand U5200 (N_5200,N_4993,N_4799);
xnor U5201 (N_5201,N_4763,N_4918);
nand U5202 (N_5202,N_4996,N_4981);
nor U5203 (N_5203,N_4861,N_4968);
or U5204 (N_5204,N_4998,N_4753);
nand U5205 (N_5205,N_4944,N_4941);
xor U5206 (N_5206,N_4755,N_4792);
or U5207 (N_5207,N_4919,N_4863);
nor U5208 (N_5208,N_4879,N_4819);
nand U5209 (N_5209,N_4944,N_4811);
nand U5210 (N_5210,N_4952,N_4860);
nor U5211 (N_5211,N_4773,N_4803);
nand U5212 (N_5212,N_4899,N_4794);
and U5213 (N_5213,N_4967,N_4832);
nand U5214 (N_5214,N_4961,N_4900);
or U5215 (N_5215,N_4933,N_4919);
xor U5216 (N_5216,N_4973,N_4936);
nor U5217 (N_5217,N_4759,N_4786);
nor U5218 (N_5218,N_4979,N_4784);
xnor U5219 (N_5219,N_4752,N_4916);
nor U5220 (N_5220,N_4972,N_4817);
nand U5221 (N_5221,N_4890,N_4848);
nand U5222 (N_5222,N_4800,N_4914);
nor U5223 (N_5223,N_4926,N_4913);
nor U5224 (N_5224,N_4824,N_4790);
nand U5225 (N_5225,N_4914,N_4868);
nand U5226 (N_5226,N_4857,N_4909);
nor U5227 (N_5227,N_4805,N_4919);
nor U5228 (N_5228,N_4918,N_4842);
nor U5229 (N_5229,N_4774,N_4824);
or U5230 (N_5230,N_4831,N_4893);
and U5231 (N_5231,N_4899,N_4824);
or U5232 (N_5232,N_4805,N_4759);
nand U5233 (N_5233,N_4913,N_4887);
or U5234 (N_5234,N_4823,N_4768);
or U5235 (N_5235,N_4896,N_4863);
nor U5236 (N_5236,N_4801,N_4905);
xnor U5237 (N_5237,N_4935,N_4998);
nor U5238 (N_5238,N_4753,N_4796);
xnor U5239 (N_5239,N_4938,N_4911);
nand U5240 (N_5240,N_4864,N_4869);
nand U5241 (N_5241,N_4756,N_4925);
or U5242 (N_5242,N_4779,N_4869);
xnor U5243 (N_5243,N_4884,N_4839);
or U5244 (N_5244,N_4829,N_4923);
or U5245 (N_5245,N_4893,N_4782);
nor U5246 (N_5246,N_4858,N_4914);
xnor U5247 (N_5247,N_4955,N_4841);
nand U5248 (N_5248,N_4842,N_4854);
xnor U5249 (N_5249,N_4885,N_4783);
nor U5250 (N_5250,N_5032,N_5216);
nor U5251 (N_5251,N_5057,N_5199);
or U5252 (N_5252,N_5123,N_5136);
nand U5253 (N_5253,N_5115,N_5087);
nand U5254 (N_5254,N_5065,N_5086);
nor U5255 (N_5255,N_5248,N_5177);
or U5256 (N_5256,N_5092,N_5074);
nand U5257 (N_5257,N_5040,N_5242);
and U5258 (N_5258,N_5240,N_5021);
or U5259 (N_5259,N_5193,N_5037);
nor U5260 (N_5260,N_5214,N_5091);
nor U5261 (N_5261,N_5130,N_5201);
or U5262 (N_5262,N_5102,N_5034);
and U5263 (N_5263,N_5150,N_5135);
xor U5264 (N_5264,N_5243,N_5129);
xor U5265 (N_5265,N_5134,N_5198);
nor U5266 (N_5266,N_5247,N_5112);
or U5267 (N_5267,N_5205,N_5159);
xor U5268 (N_5268,N_5111,N_5038);
nor U5269 (N_5269,N_5093,N_5015);
nand U5270 (N_5270,N_5067,N_5045);
nor U5271 (N_5271,N_5178,N_5025);
nor U5272 (N_5272,N_5225,N_5106);
nor U5273 (N_5273,N_5138,N_5189);
xnor U5274 (N_5274,N_5051,N_5039);
xnor U5275 (N_5275,N_5209,N_5171);
nor U5276 (N_5276,N_5071,N_5098);
or U5277 (N_5277,N_5140,N_5008);
or U5278 (N_5278,N_5104,N_5126);
xor U5279 (N_5279,N_5089,N_5174);
and U5280 (N_5280,N_5183,N_5195);
or U5281 (N_5281,N_5192,N_5233);
xor U5282 (N_5282,N_5128,N_5097);
nor U5283 (N_5283,N_5033,N_5110);
xor U5284 (N_5284,N_5223,N_5185);
or U5285 (N_5285,N_5167,N_5131);
and U5286 (N_5286,N_5113,N_5127);
nor U5287 (N_5287,N_5217,N_5068);
and U5288 (N_5288,N_5179,N_5244);
or U5289 (N_5289,N_5002,N_5011);
and U5290 (N_5290,N_5017,N_5026);
xnor U5291 (N_5291,N_5157,N_5154);
xnor U5292 (N_5292,N_5031,N_5180);
nor U5293 (N_5293,N_5018,N_5082);
nand U5294 (N_5294,N_5058,N_5095);
xor U5295 (N_5295,N_5121,N_5103);
and U5296 (N_5296,N_5149,N_5050);
nand U5297 (N_5297,N_5156,N_5190);
nor U5298 (N_5298,N_5213,N_5004);
or U5299 (N_5299,N_5063,N_5191);
and U5300 (N_5300,N_5084,N_5020);
or U5301 (N_5301,N_5224,N_5054);
nor U5302 (N_5302,N_5206,N_5030);
nor U5303 (N_5303,N_5062,N_5083);
xor U5304 (N_5304,N_5114,N_5194);
nand U5305 (N_5305,N_5125,N_5022);
nand U5306 (N_5306,N_5215,N_5064);
nor U5307 (N_5307,N_5028,N_5075);
nand U5308 (N_5308,N_5047,N_5066);
nand U5309 (N_5309,N_5186,N_5155);
nor U5310 (N_5310,N_5007,N_5220);
nor U5311 (N_5311,N_5073,N_5006);
nand U5312 (N_5312,N_5041,N_5145);
and U5313 (N_5313,N_5212,N_5019);
nor U5314 (N_5314,N_5117,N_5148);
nand U5315 (N_5315,N_5096,N_5188);
nand U5316 (N_5316,N_5056,N_5230);
or U5317 (N_5317,N_5184,N_5196);
nand U5318 (N_5318,N_5202,N_5099);
nor U5319 (N_5319,N_5000,N_5181);
nand U5320 (N_5320,N_5200,N_5035);
nor U5321 (N_5321,N_5236,N_5070);
and U5322 (N_5322,N_5118,N_5053);
nand U5323 (N_5323,N_5228,N_5119);
nor U5324 (N_5324,N_5080,N_5059);
and U5325 (N_5325,N_5218,N_5010);
or U5326 (N_5326,N_5078,N_5061);
or U5327 (N_5327,N_5014,N_5237);
xnor U5328 (N_5328,N_5208,N_5085);
nor U5329 (N_5329,N_5101,N_5153);
or U5330 (N_5330,N_5162,N_5163);
and U5331 (N_5331,N_5133,N_5023);
nand U5332 (N_5332,N_5197,N_5175);
xor U5333 (N_5333,N_5235,N_5120);
nor U5334 (N_5334,N_5219,N_5108);
nand U5335 (N_5335,N_5234,N_5029);
xor U5336 (N_5336,N_5227,N_5144);
nor U5337 (N_5337,N_5147,N_5081);
xnor U5338 (N_5338,N_5168,N_5001);
and U5339 (N_5339,N_5207,N_5165);
xnor U5340 (N_5340,N_5158,N_5222);
nor U5341 (N_5341,N_5048,N_5241);
xnor U5342 (N_5342,N_5152,N_5012);
or U5343 (N_5343,N_5164,N_5076);
nor U5344 (N_5344,N_5079,N_5170);
nand U5345 (N_5345,N_5210,N_5043);
and U5346 (N_5346,N_5146,N_5166);
xor U5347 (N_5347,N_5060,N_5042);
xnor U5348 (N_5348,N_5109,N_5049);
and U5349 (N_5349,N_5116,N_5169);
and U5350 (N_5350,N_5239,N_5069);
xor U5351 (N_5351,N_5203,N_5231);
and U5352 (N_5352,N_5088,N_5238);
xnor U5353 (N_5353,N_5094,N_5182);
and U5354 (N_5354,N_5142,N_5055);
and U5355 (N_5355,N_5211,N_5132);
or U5356 (N_5356,N_5124,N_5221);
and U5357 (N_5357,N_5016,N_5141);
or U5358 (N_5358,N_5077,N_5122);
or U5359 (N_5359,N_5100,N_5249);
and U5360 (N_5360,N_5090,N_5027);
or U5361 (N_5361,N_5105,N_5151);
nor U5362 (N_5362,N_5107,N_5046);
xor U5363 (N_5363,N_5160,N_5173);
nand U5364 (N_5364,N_5176,N_5226);
and U5365 (N_5365,N_5003,N_5187);
xnor U5366 (N_5366,N_5204,N_5137);
and U5367 (N_5367,N_5246,N_5005);
xor U5368 (N_5368,N_5161,N_5013);
xor U5369 (N_5369,N_5009,N_5072);
xnor U5370 (N_5370,N_5232,N_5044);
xnor U5371 (N_5371,N_5139,N_5245);
nand U5372 (N_5372,N_5172,N_5052);
nor U5373 (N_5373,N_5024,N_5229);
xnor U5374 (N_5374,N_5143,N_5036);
xnor U5375 (N_5375,N_5059,N_5139);
xor U5376 (N_5376,N_5136,N_5188);
xor U5377 (N_5377,N_5140,N_5247);
nor U5378 (N_5378,N_5053,N_5054);
xnor U5379 (N_5379,N_5016,N_5130);
and U5380 (N_5380,N_5104,N_5177);
xnor U5381 (N_5381,N_5135,N_5051);
nand U5382 (N_5382,N_5214,N_5028);
nand U5383 (N_5383,N_5208,N_5048);
and U5384 (N_5384,N_5182,N_5148);
nor U5385 (N_5385,N_5207,N_5105);
nand U5386 (N_5386,N_5184,N_5032);
or U5387 (N_5387,N_5055,N_5149);
or U5388 (N_5388,N_5177,N_5240);
nor U5389 (N_5389,N_5067,N_5033);
and U5390 (N_5390,N_5086,N_5061);
and U5391 (N_5391,N_5050,N_5206);
or U5392 (N_5392,N_5079,N_5222);
nor U5393 (N_5393,N_5202,N_5025);
nand U5394 (N_5394,N_5012,N_5107);
nand U5395 (N_5395,N_5039,N_5144);
nand U5396 (N_5396,N_5007,N_5040);
nand U5397 (N_5397,N_5247,N_5216);
or U5398 (N_5398,N_5215,N_5002);
nor U5399 (N_5399,N_5173,N_5062);
xor U5400 (N_5400,N_5108,N_5064);
and U5401 (N_5401,N_5044,N_5109);
and U5402 (N_5402,N_5097,N_5104);
nand U5403 (N_5403,N_5153,N_5063);
nor U5404 (N_5404,N_5155,N_5177);
and U5405 (N_5405,N_5045,N_5192);
nand U5406 (N_5406,N_5160,N_5242);
or U5407 (N_5407,N_5169,N_5032);
or U5408 (N_5408,N_5147,N_5012);
or U5409 (N_5409,N_5237,N_5104);
or U5410 (N_5410,N_5048,N_5069);
and U5411 (N_5411,N_5110,N_5248);
nor U5412 (N_5412,N_5029,N_5022);
nor U5413 (N_5413,N_5066,N_5232);
nor U5414 (N_5414,N_5067,N_5145);
nor U5415 (N_5415,N_5147,N_5204);
xnor U5416 (N_5416,N_5039,N_5228);
and U5417 (N_5417,N_5235,N_5068);
nand U5418 (N_5418,N_5075,N_5209);
or U5419 (N_5419,N_5120,N_5193);
xnor U5420 (N_5420,N_5168,N_5242);
or U5421 (N_5421,N_5018,N_5172);
and U5422 (N_5422,N_5107,N_5064);
or U5423 (N_5423,N_5202,N_5237);
xnor U5424 (N_5424,N_5222,N_5047);
or U5425 (N_5425,N_5027,N_5111);
or U5426 (N_5426,N_5242,N_5028);
nor U5427 (N_5427,N_5187,N_5097);
and U5428 (N_5428,N_5032,N_5179);
or U5429 (N_5429,N_5243,N_5132);
xor U5430 (N_5430,N_5233,N_5051);
xnor U5431 (N_5431,N_5099,N_5174);
and U5432 (N_5432,N_5240,N_5184);
xnor U5433 (N_5433,N_5176,N_5177);
nand U5434 (N_5434,N_5232,N_5040);
or U5435 (N_5435,N_5040,N_5082);
nand U5436 (N_5436,N_5003,N_5063);
nand U5437 (N_5437,N_5222,N_5057);
nor U5438 (N_5438,N_5077,N_5189);
nor U5439 (N_5439,N_5051,N_5035);
nor U5440 (N_5440,N_5064,N_5126);
xnor U5441 (N_5441,N_5155,N_5139);
and U5442 (N_5442,N_5148,N_5210);
and U5443 (N_5443,N_5162,N_5085);
xnor U5444 (N_5444,N_5014,N_5195);
and U5445 (N_5445,N_5017,N_5223);
nand U5446 (N_5446,N_5072,N_5217);
nor U5447 (N_5447,N_5204,N_5085);
nand U5448 (N_5448,N_5098,N_5117);
nor U5449 (N_5449,N_5066,N_5243);
nand U5450 (N_5450,N_5137,N_5032);
xnor U5451 (N_5451,N_5106,N_5144);
and U5452 (N_5452,N_5063,N_5083);
and U5453 (N_5453,N_5087,N_5226);
xnor U5454 (N_5454,N_5229,N_5187);
and U5455 (N_5455,N_5231,N_5017);
xnor U5456 (N_5456,N_5025,N_5194);
nor U5457 (N_5457,N_5023,N_5049);
nand U5458 (N_5458,N_5128,N_5069);
and U5459 (N_5459,N_5203,N_5035);
and U5460 (N_5460,N_5199,N_5073);
xnor U5461 (N_5461,N_5107,N_5034);
xor U5462 (N_5462,N_5058,N_5198);
or U5463 (N_5463,N_5203,N_5173);
or U5464 (N_5464,N_5123,N_5024);
nor U5465 (N_5465,N_5132,N_5227);
or U5466 (N_5466,N_5174,N_5110);
nor U5467 (N_5467,N_5056,N_5117);
or U5468 (N_5468,N_5120,N_5080);
nor U5469 (N_5469,N_5005,N_5125);
nor U5470 (N_5470,N_5175,N_5001);
xor U5471 (N_5471,N_5038,N_5087);
or U5472 (N_5472,N_5062,N_5244);
nor U5473 (N_5473,N_5039,N_5225);
or U5474 (N_5474,N_5127,N_5155);
nor U5475 (N_5475,N_5082,N_5189);
nor U5476 (N_5476,N_5184,N_5232);
xor U5477 (N_5477,N_5227,N_5220);
and U5478 (N_5478,N_5077,N_5162);
nand U5479 (N_5479,N_5042,N_5208);
xnor U5480 (N_5480,N_5148,N_5198);
and U5481 (N_5481,N_5123,N_5082);
nand U5482 (N_5482,N_5210,N_5208);
nand U5483 (N_5483,N_5179,N_5071);
and U5484 (N_5484,N_5206,N_5122);
nand U5485 (N_5485,N_5194,N_5238);
xnor U5486 (N_5486,N_5216,N_5014);
xor U5487 (N_5487,N_5150,N_5183);
or U5488 (N_5488,N_5134,N_5217);
xor U5489 (N_5489,N_5000,N_5108);
or U5490 (N_5490,N_5189,N_5159);
or U5491 (N_5491,N_5061,N_5179);
or U5492 (N_5492,N_5106,N_5205);
or U5493 (N_5493,N_5113,N_5063);
xor U5494 (N_5494,N_5102,N_5099);
and U5495 (N_5495,N_5093,N_5086);
nand U5496 (N_5496,N_5196,N_5171);
xnor U5497 (N_5497,N_5245,N_5035);
or U5498 (N_5498,N_5209,N_5193);
xnor U5499 (N_5499,N_5144,N_5069);
and U5500 (N_5500,N_5345,N_5419);
xnor U5501 (N_5501,N_5466,N_5301);
xnor U5502 (N_5502,N_5258,N_5333);
and U5503 (N_5503,N_5274,N_5424);
and U5504 (N_5504,N_5308,N_5457);
and U5505 (N_5505,N_5487,N_5423);
nand U5506 (N_5506,N_5484,N_5366);
and U5507 (N_5507,N_5417,N_5414);
nand U5508 (N_5508,N_5488,N_5287);
nor U5509 (N_5509,N_5281,N_5320);
nand U5510 (N_5510,N_5363,N_5260);
or U5511 (N_5511,N_5275,N_5293);
xor U5512 (N_5512,N_5328,N_5398);
or U5513 (N_5513,N_5490,N_5339);
nand U5514 (N_5514,N_5409,N_5393);
xor U5515 (N_5515,N_5462,N_5364);
and U5516 (N_5516,N_5429,N_5412);
nand U5517 (N_5517,N_5324,N_5459);
or U5518 (N_5518,N_5430,N_5476);
xor U5519 (N_5519,N_5439,N_5420);
nand U5520 (N_5520,N_5288,N_5388);
xor U5521 (N_5521,N_5331,N_5317);
nand U5522 (N_5522,N_5332,N_5486);
and U5523 (N_5523,N_5370,N_5468);
or U5524 (N_5524,N_5456,N_5277);
and U5525 (N_5525,N_5355,N_5329);
nand U5526 (N_5526,N_5407,N_5471);
nor U5527 (N_5527,N_5338,N_5432);
xor U5528 (N_5528,N_5428,N_5455);
or U5529 (N_5529,N_5498,N_5313);
and U5530 (N_5530,N_5465,N_5481);
and U5531 (N_5531,N_5304,N_5305);
nand U5532 (N_5532,N_5375,N_5403);
nor U5533 (N_5533,N_5354,N_5292);
and U5534 (N_5534,N_5434,N_5336);
xnor U5535 (N_5535,N_5376,N_5306);
nor U5536 (N_5536,N_5289,N_5342);
xor U5537 (N_5537,N_5351,N_5368);
or U5538 (N_5538,N_5461,N_5349);
xor U5539 (N_5539,N_5440,N_5426);
and U5540 (N_5540,N_5493,N_5496);
or U5541 (N_5541,N_5437,N_5259);
nand U5542 (N_5542,N_5396,N_5372);
nand U5543 (N_5543,N_5371,N_5452);
nor U5544 (N_5544,N_5431,N_5299);
xnor U5545 (N_5545,N_5296,N_5385);
nand U5546 (N_5546,N_5489,N_5261);
and U5547 (N_5547,N_5491,N_5360);
or U5548 (N_5548,N_5279,N_5374);
and U5549 (N_5549,N_5446,N_5303);
nand U5550 (N_5550,N_5365,N_5254);
xnor U5551 (N_5551,N_5290,N_5425);
nor U5552 (N_5552,N_5369,N_5482);
and U5553 (N_5553,N_5350,N_5269);
and U5554 (N_5554,N_5282,N_5264);
xor U5555 (N_5555,N_5309,N_5356);
or U5556 (N_5556,N_5415,N_5447);
xnor U5557 (N_5557,N_5251,N_5340);
or U5558 (N_5558,N_5458,N_5294);
xor U5559 (N_5559,N_5470,N_5344);
and U5560 (N_5560,N_5319,N_5367);
nand U5561 (N_5561,N_5406,N_5266);
or U5562 (N_5562,N_5353,N_5358);
nor U5563 (N_5563,N_5322,N_5394);
and U5564 (N_5564,N_5255,N_5302);
nor U5565 (N_5565,N_5312,N_5474);
and U5566 (N_5566,N_5263,N_5454);
and U5567 (N_5567,N_5435,N_5257);
xor U5568 (N_5568,N_5479,N_5335);
xnor U5569 (N_5569,N_5381,N_5323);
nor U5570 (N_5570,N_5295,N_5390);
nor U5571 (N_5571,N_5438,N_5377);
and U5572 (N_5572,N_5444,N_5327);
nand U5573 (N_5573,N_5405,N_5485);
nand U5574 (N_5574,N_5271,N_5348);
nand U5575 (N_5575,N_5283,N_5291);
or U5576 (N_5576,N_5300,N_5421);
or U5577 (N_5577,N_5399,N_5341);
or U5578 (N_5578,N_5347,N_5418);
or U5579 (N_5579,N_5285,N_5453);
xnor U5580 (N_5580,N_5361,N_5298);
xor U5581 (N_5581,N_5495,N_5443);
nor U5582 (N_5582,N_5463,N_5416);
nor U5583 (N_5583,N_5422,N_5404);
nand U5584 (N_5584,N_5270,N_5460);
nand U5585 (N_5585,N_5478,N_5326);
or U5586 (N_5586,N_5383,N_5497);
or U5587 (N_5587,N_5473,N_5330);
or U5588 (N_5588,N_5448,N_5411);
xnor U5589 (N_5589,N_5307,N_5252);
nor U5590 (N_5590,N_5362,N_5262);
nand U5591 (N_5591,N_5256,N_5286);
and U5592 (N_5592,N_5268,N_5494);
nor U5593 (N_5593,N_5265,N_5278);
nand U5594 (N_5594,N_5310,N_5314);
xnor U5595 (N_5595,N_5397,N_5472);
nand U5596 (N_5596,N_5284,N_5402);
nand U5597 (N_5597,N_5389,N_5311);
nor U5598 (N_5598,N_5445,N_5373);
and U5599 (N_5599,N_5475,N_5343);
nand U5600 (N_5600,N_5469,N_5410);
or U5601 (N_5601,N_5273,N_5467);
nor U5602 (N_5602,N_5321,N_5413);
xor U5603 (N_5603,N_5386,N_5387);
nand U5604 (N_5604,N_5315,N_5280);
nand U5605 (N_5605,N_5441,N_5400);
or U5606 (N_5606,N_5427,N_5297);
and U5607 (N_5607,N_5357,N_5449);
xnor U5608 (N_5608,N_5253,N_5442);
or U5609 (N_5609,N_5352,N_5382);
nor U5610 (N_5610,N_5408,N_5276);
nand U5611 (N_5611,N_5325,N_5378);
xor U5612 (N_5612,N_5483,N_5334);
nand U5613 (N_5613,N_5337,N_5499);
or U5614 (N_5614,N_5379,N_5267);
nor U5615 (N_5615,N_5451,N_5359);
xnor U5616 (N_5616,N_5480,N_5250);
nor U5617 (N_5617,N_5346,N_5392);
or U5618 (N_5618,N_5316,N_5391);
or U5619 (N_5619,N_5384,N_5436);
or U5620 (N_5620,N_5492,N_5401);
or U5621 (N_5621,N_5395,N_5318);
nand U5622 (N_5622,N_5272,N_5380);
nand U5623 (N_5623,N_5464,N_5450);
and U5624 (N_5624,N_5433,N_5477);
nand U5625 (N_5625,N_5447,N_5483);
nor U5626 (N_5626,N_5289,N_5381);
xor U5627 (N_5627,N_5393,N_5384);
and U5628 (N_5628,N_5403,N_5320);
nand U5629 (N_5629,N_5387,N_5300);
nor U5630 (N_5630,N_5254,N_5389);
and U5631 (N_5631,N_5261,N_5370);
nand U5632 (N_5632,N_5320,N_5283);
nand U5633 (N_5633,N_5454,N_5488);
or U5634 (N_5634,N_5307,N_5415);
or U5635 (N_5635,N_5380,N_5491);
or U5636 (N_5636,N_5273,N_5404);
nor U5637 (N_5637,N_5254,N_5470);
xnor U5638 (N_5638,N_5405,N_5429);
nand U5639 (N_5639,N_5323,N_5339);
nand U5640 (N_5640,N_5387,N_5480);
and U5641 (N_5641,N_5269,N_5361);
xor U5642 (N_5642,N_5335,N_5373);
xor U5643 (N_5643,N_5317,N_5453);
nand U5644 (N_5644,N_5357,N_5364);
nand U5645 (N_5645,N_5285,N_5377);
or U5646 (N_5646,N_5489,N_5279);
xnor U5647 (N_5647,N_5364,N_5288);
and U5648 (N_5648,N_5450,N_5472);
and U5649 (N_5649,N_5365,N_5267);
nand U5650 (N_5650,N_5445,N_5398);
or U5651 (N_5651,N_5288,N_5335);
nand U5652 (N_5652,N_5347,N_5273);
xor U5653 (N_5653,N_5289,N_5306);
nand U5654 (N_5654,N_5264,N_5357);
xor U5655 (N_5655,N_5448,N_5384);
or U5656 (N_5656,N_5337,N_5270);
nand U5657 (N_5657,N_5262,N_5496);
nor U5658 (N_5658,N_5464,N_5447);
xnor U5659 (N_5659,N_5305,N_5384);
xnor U5660 (N_5660,N_5256,N_5311);
and U5661 (N_5661,N_5490,N_5323);
and U5662 (N_5662,N_5295,N_5482);
nor U5663 (N_5663,N_5408,N_5346);
and U5664 (N_5664,N_5420,N_5292);
and U5665 (N_5665,N_5419,N_5349);
nor U5666 (N_5666,N_5267,N_5479);
nor U5667 (N_5667,N_5324,N_5330);
or U5668 (N_5668,N_5331,N_5428);
nor U5669 (N_5669,N_5434,N_5403);
or U5670 (N_5670,N_5301,N_5359);
nor U5671 (N_5671,N_5314,N_5415);
nor U5672 (N_5672,N_5341,N_5423);
and U5673 (N_5673,N_5423,N_5493);
or U5674 (N_5674,N_5469,N_5271);
nor U5675 (N_5675,N_5334,N_5265);
xnor U5676 (N_5676,N_5376,N_5413);
nand U5677 (N_5677,N_5275,N_5470);
nor U5678 (N_5678,N_5319,N_5254);
and U5679 (N_5679,N_5331,N_5464);
nor U5680 (N_5680,N_5257,N_5275);
xnor U5681 (N_5681,N_5478,N_5464);
xnor U5682 (N_5682,N_5351,N_5404);
and U5683 (N_5683,N_5468,N_5397);
nor U5684 (N_5684,N_5285,N_5444);
nand U5685 (N_5685,N_5391,N_5393);
nor U5686 (N_5686,N_5465,N_5469);
xnor U5687 (N_5687,N_5355,N_5310);
and U5688 (N_5688,N_5282,N_5287);
nor U5689 (N_5689,N_5454,N_5419);
and U5690 (N_5690,N_5387,N_5430);
xor U5691 (N_5691,N_5454,N_5407);
nand U5692 (N_5692,N_5270,N_5349);
and U5693 (N_5693,N_5266,N_5448);
nand U5694 (N_5694,N_5314,N_5281);
and U5695 (N_5695,N_5313,N_5334);
and U5696 (N_5696,N_5490,N_5292);
nand U5697 (N_5697,N_5282,N_5260);
nor U5698 (N_5698,N_5459,N_5322);
nor U5699 (N_5699,N_5264,N_5365);
nor U5700 (N_5700,N_5306,N_5283);
nor U5701 (N_5701,N_5261,N_5280);
and U5702 (N_5702,N_5334,N_5452);
nor U5703 (N_5703,N_5252,N_5386);
or U5704 (N_5704,N_5423,N_5305);
or U5705 (N_5705,N_5359,N_5387);
and U5706 (N_5706,N_5288,N_5400);
and U5707 (N_5707,N_5328,N_5385);
or U5708 (N_5708,N_5351,N_5296);
nor U5709 (N_5709,N_5349,N_5494);
and U5710 (N_5710,N_5420,N_5402);
nor U5711 (N_5711,N_5371,N_5341);
xnor U5712 (N_5712,N_5386,N_5428);
and U5713 (N_5713,N_5462,N_5293);
nand U5714 (N_5714,N_5254,N_5458);
or U5715 (N_5715,N_5335,N_5372);
or U5716 (N_5716,N_5494,N_5403);
or U5717 (N_5717,N_5318,N_5476);
nor U5718 (N_5718,N_5494,N_5450);
nor U5719 (N_5719,N_5363,N_5303);
nor U5720 (N_5720,N_5420,N_5344);
or U5721 (N_5721,N_5355,N_5412);
nor U5722 (N_5722,N_5309,N_5471);
or U5723 (N_5723,N_5306,N_5349);
and U5724 (N_5724,N_5481,N_5380);
xor U5725 (N_5725,N_5392,N_5282);
nor U5726 (N_5726,N_5373,N_5285);
or U5727 (N_5727,N_5366,N_5452);
or U5728 (N_5728,N_5343,N_5401);
nor U5729 (N_5729,N_5427,N_5260);
nor U5730 (N_5730,N_5411,N_5369);
xor U5731 (N_5731,N_5409,N_5499);
xor U5732 (N_5732,N_5496,N_5382);
nor U5733 (N_5733,N_5376,N_5276);
and U5734 (N_5734,N_5395,N_5421);
nor U5735 (N_5735,N_5328,N_5387);
nand U5736 (N_5736,N_5488,N_5427);
xor U5737 (N_5737,N_5431,N_5324);
nor U5738 (N_5738,N_5256,N_5272);
xor U5739 (N_5739,N_5336,N_5421);
or U5740 (N_5740,N_5282,N_5294);
nand U5741 (N_5741,N_5497,N_5378);
nand U5742 (N_5742,N_5412,N_5286);
nand U5743 (N_5743,N_5276,N_5304);
nor U5744 (N_5744,N_5445,N_5409);
nand U5745 (N_5745,N_5370,N_5421);
nand U5746 (N_5746,N_5446,N_5316);
xnor U5747 (N_5747,N_5265,N_5446);
or U5748 (N_5748,N_5473,N_5357);
nand U5749 (N_5749,N_5472,N_5344);
or U5750 (N_5750,N_5650,N_5523);
nand U5751 (N_5751,N_5694,N_5656);
or U5752 (N_5752,N_5545,N_5647);
and U5753 (N_5753,N_5689,N_5516);
or U5754 (N_5754,N_5531,N_5681);
xnor U5755 (N_5755,N_5646,N_5543);
xnor U5756 (N_5756,N_5594,N_5620);
xor U5757 (N_5757,N_5500,N_5574);
and U5758 (N_5758,N_5718,N_5624);
nand U5759 (N_5759,N_5520,N_5706);
xor U5760 (N_5760,N_5579,N_5611);
nor U5761 (N_5761,N_5577,N_5599);
and U5762 (N_5762,N_5726,N_5617);
xnor U5763 (N_5763,N_5512,N_5600);
nand U5764 (N_5764,N_5648,N_5583);
nand U5765 (N_5765,N_5566,N_5502);
or U5766 (N_5766,N_5697,N_5544);
and U5767 (N_5767,N_5526,N_5529);
xor U5768 (N_5768,N_5559,N_5554);
nand U5769 (N_5769,N_5614,N_5735);
or U5770 (N_5770,N_5572,N_5567);
xor U5771 (N_5771,N_5597,N_5503);
nand U5772 (N_5772,N_5524,N_5743);
and U5773 (N_5773,N_5513,N_5675);
nor U5774 (N_5774,N_5685,N_5549);
xor U5775 (N_5775,N_5686,N_5608);
xor U5776 (N_5776,N_5716,N_5717);
nor U5777 (N_5777,N_5683,N_5514);
and U5778 (N_5778,N_5555,N_5507);
xor U5779 (N_5779,N_5619,N_5715);
and U5780 (N_5780,N_5562,N_5542);
nand U5781 (N_5781,N_5655,N_5505);
nand U5782 (N_5782,N_5688,N_5664);
nand U5783 (N_5783,N_5584,N_5733);
nor U5784 (N_5784,N_5713,N_5571);
xnor U5785 (N_5785,N_5747,N_5746);
and U5786 (N_5786,N_5725,N_5556);
nor U5787 (N_5787,N_5720,N_5532);
xnor U5788 (N_5788,N_5744,N_5628);
nand U5789 (N_5789,N_5588,N_5550);
or U5790 (N_5790,N_5652,N_5727);
nand U5791 (N_5791,N_5721,N_5527);
or U5792 (N_5792,N_5602,N_5616);
nor U5793 (N_5793,N_5712,N_5690);
or U5794 (N_5794,N_5667,N_5615);
or U5795 (N_5795,N_5639,N_5724);
xnor U5796 (N_5796,N_5504,N_5642);
nand U5797 (N_5797,N_5591,N_5636);
or U5798 (N_5798,N_5530,N_5623);
xor U5799 (N_5799,N_5578,N_5627);
nand U5800 (N_5800,N_5569,N_5573);
and U5801 (N_5801,N_5719,N_5576);
or U5802 (N_5802,N_5547,N_5551);
nand U5803 (N_5803,N_5593,N_5691);
nor U5804 (N_5804,N_5737,N_5640);
xor U5805 (N_5805,N_5643,N_5748);
nor U5806 (N_5806,N_5663,N_5708);
xnor U5807 (N_5807,N_5680,N_5638);
nor U5808 (N_5808,N_5651,N_5521);
and U5809 (N_5809,N_5560,N_5687);
nand U5810 (N_5810,N_5590,N_5739);
nor U5811 (N_5811,N_5672,N_5604);
xnor U5812 (N_5812,N_5509,N_5536);
nand U5813 (N_5813,N_5632,N_5580);
xor U5814 (N_5814,N_5618,N_5700);
xor U5815 (N_5815,N_5671,N_5666);
nand U5816 (N_5816,N_5695,N_5653);
nor U5817 (N_5817,N_5629,N_5511);
xor U5818 (N_5818,N_5607,N_5541);
or U5819 (N_5819,N_5561,N_5501);
and U5820 (N_5820,N_5654,N_5519);
and U5821 (N_5821,N_5563,N_5709);
xnor U5822 (N_5822,N_5538,N_5670);
or U5823 (N_5823,N_5621,N_5644);
nand U5824 (N_5824,N_5601,N_5575);
nand U5825 (N_5825,N_5701,N_5609);
nor U5826 (N_5826,N_5525,N_5634);
and U5827 (N_5827,N_5605,N_5741);
and U5828 (N_5828,N_5635,N_5728);
nand U5829 (N_5829,N_5669,N_5696);
nand U5830 (N_5830,N_5722,N_5613);
and U5831 (N_5831,N_5676,N_5630);
or U5832 (N_5832,N_5537,N_5692);
nor U5833 (N_5833,N_5649,N_5587);
or U5834 (N_5834,N_5714,N_5658);
or U5835 (N_5835,N_5533,N_5535);
xnor U5836 (N_5836,N_5645,N_5506);
nor U5837 (N_5837,N_5704,N_5564);
nor U5838 (N_5838,N_5592,N_5665);
and U5839 (N_5839,N_5582,N_5702);
nor U5840 (N_5840,N_5633,N_5699);
nor U5841 (N_5841,N_5570,N_5707);
nor U5842 (N_5842,N_5585,N_5657);
nor U5843 (N_5843,N_5610,N_5534);
and U5844 (N_5844,N_5711,N_5673);
and U5845 (N_5845,N_5738,N_5581);
nand U5846 (N_5846,N_5606,N_5703);
nand U5847 (N_5847,N_5732,N_5661);
or U5848 (N_5848,N_5729,N_5742);
xor U5849 (N_5849,N_5622,N_5625);
nor U5850 (N_5850,N_5595,N_5518);
or U5851 (N_5851,N_5659,N_5730);
nand U5852 (N_5852,N_5603,N_5734);
nor U5853 (N_5853,N_5693,N_5705);
nor U5854 (N_5854,N_5517,N_5598);
xor U5855 (N_5855,N_5508,N_5522);
xor U5856 (N_5856,N_5510,N_5745);
and U5857 (N_5857,N_5612,N_5710);
or U5858 (N_5858,N_5552,N_5684);
or U5859 (N_5859,N_5631,N_5637);
or U5860 (N_5860,N_5540,N_5586);
or U5861 (N_5861,N_5723,N_5641);
xnor U5862 (N_5862,N_5553,N_5679);
xnor U5863 (N_5863,N_5558,N_5660);
xnor U5864 (N_5864,N_5749,N_5589);
and U5865 (N_5865,N_5668,N_5736);
nand U5866 (N_5866,N_5565,N_5626);
and U5867 (N_5867,N_5568,N_5596);
and U5868 (N_5868,N_5678,N_5548);
and U5869 (N_5869,N_5515,N_5662);
xnor U5870 (N_5870,N_5698,N_5740);
and U5871 (N_5871,N_5677,N_5731);
nor U5872 (N_5872,N_5528,N_5557);
nor U5873 (N_5873,N_5682,N_5539);
nand U5874 (N_5874,N_5674,N_5546);
and U5875 (N_5875,N_5727,N_5717);
and U5876 (N_5876,N_5562,N_5513);
or U5877 (N_5877,N_5505,N_5657);
or U5878 (N_5878,N_5569,N_5636);
or U5879 (N_5879,N_5698,N_5607);
and U5880 (N_5880,N_5628,N_5524);
and U5881 (N_5881,N_5707,N_5552);
nor U5882 (N_5882,N_5744,N_5625);
and U5883 (N_5883,N_5617,N_5660);
and U5884 (N_5884,N_5714,N_5724);
nand U5885 (N_5885,N_5523,N_5695);
xor U5886 (N_5886,N_5549,N_5619);
nor U5887 (N_5887,N_5514,N_5631);
or U5888 (N_5888,N_5688,N_5553);
xnor U5889 (N_5889,N_5524,N_5701);
nor U5890 (N_5890,N_5513,N_5554);
xnor U5891 (N_5891,N_5716,N_5654);
nor U5892 (N_5892,N_5558,N_5506);
nor U5893 (N_5893,N_5625,N_5726);
nor U5894 (N_5894,N_5585,N_5543);
and U5895 (N_5895,N_5588,N_5634);
nand U5896 (N_5896,N_5526,N_5670);
xor U5897 (N_5897,N_5615,N_5581);
nor U5898 (N_5898,N_5550,N_5608);
nor U5899 (N_5899,N_5700,N_5623);
nand U5900 (N_5900,N_5674,N_5729);
xnor U5901 (N_5901,N_5730,N_5561);
or U5902 (N_5902,N_5715,N_5601);
or U5903 (N_5903,N_5614,N_5641);
and U5904 (N_5904,N_5720,N_5728);
nand U5905 (N_5905,N_5506,N_5540);
or U5906 (N_5906,N_5511,N_5634);
or U5907 (N_5907,N_5518,N_5611);
nor U5908 (N_5908,N_5673,N_5610);
xnor U5909 (N_5909,N_5520,N_5730);
nand U5910 (N_5910,N_5533,N_5604);
nand U5911 (N_5911,N_5674,N_5747);
xnor U5912 (N_5912,N_5515,N_5645);
nand U5913 (N_5913,N_5706,N_5749);
or U5914 (N_5914,N_5526,N_5664);
nand U5915 (N_5915,N_5517,N_5571);
or U5916 (N_5916,N_5609,N_5594);
or U5917 (N_5917,N_5654,N_5721);
nand U5918 (N_5918,N_5593,N_5592);
and U5919 (N_5919,N_5686,N_5551);
nor U5920 (N_5920,N_5583,N_5532);
and U5921 (N_5921,N_5526,N_5594);
nor U5922 (N_5922,N_5742,N_5555);
xnor U5923 (N_5923,N_5626,N_5517);
nand U5924 (N_5924,N_5571,N_5742);
and U5925 (N_5925,N_5652,N_5621);
nand U5926 (N_5926,N_5681,N_5506);
and U5927 (N_5927,N_5531,N_5710);
nand U5928 (N_5928,N_5519,N_5686);
or U5929 (N_5929,N_5573,N_5732);
or U5930 (N_5930,N_5542,N_5663);
nand U5931 (N_5931,N_5715,N_5646);
xnor U5932 (N_5932,N_5559,N_5603);
and U5933 (N_5933,N_5690,N_5521);
or U5934 (N_5934,N_5716,N_5718);
and U5935 (N_5935,N_5636,N_5713);
or U5936 (N_5936,N_5668,N_5572);
or U5937 (N_5937,N_5583,N_5683);
or U5938 (N_5938,N_5502,N_5583);
nand U5939 (N_5939,N_5644,N_5503);
nand U5940 (N_5940,N_5749,N_5600);
nor U5941 (N_5941,N_5595,N_5668);
and U5942 (N_5942,N_5523,N_5661);
xor U5943 (N_5943,N_5500,N_5593);
and U5944 (N_5944,N_5569,N_5703);
nand U5945 (N_5945,N_5680,N_5731);
xnor U5946 (N_5946,N_5560,N_5602);
or U5947 (N_5947,N_5520,N_5743);
nand U5948 (N_5948,N_5613,N_5738);
or U5949 (N_5949,N_5586,N_5535);
xnor U5950 (N_5950,N_5690,N_5500);
xnor U5951 (N_5951,N_5550,N_5648);
or U5952 (N_5952,N_5672,N_5733);
xor U5953 (N_5953,N_5616,N_5605);
nand U5954 (N_5954,N_5591,N_5516);
nand U5955 (N_5955,N_5742,N_5720);
xor U5956 (N_5956,N_5525,N_5588);
and U5957 (N_5957,N_5512,N_5505);
nor U5958 (N_5958,N_5534,N_5740);
xor U5959 (N_5959,N_5643,N_5647);
or U5960 (N_5960,N_5542,N_5642);
xnor U5961 (N_5961,N_5568,N_5585);
and U5962 (N_5962,N_5567,N_5659);
nor U5963 (N_5963,N_5709,N_5602);
or U5964 (N_5964,N_5511,N_5674);
and U5965 (N_5965,N_5730,N_5698);
xnor U5966 (N_5966,N_5714,N_5512);
and U5967 (N_5967,N_5725,N_5715);
nor U5968 (N_5968,N_5740,N_5744);
xor U5969 (N_5969,N_5554,N_5664);
nand U5970 (N_5970,N_5587,N_5701);
nand U5971 (N_5971,N_5611,N_5506);
xnor U5972 (N_5972,N_5698,N_5732);
nor U5973 (N_5973,N_5683,N_5585);
or U5974 (N_5974,N_5510,N_5657);
nor U5975 (N_5975,N_5524,N_5693);
nand U5976 (N_5976,N_5598,N_5688);
xor U5977 (N_5977,N_5686,N_5727);
xor U5978 (N_5978,N_5748,N_5588);
nor U5979 (N_5979,N_5557,N_5627);
and U5980 (N_5980,N_5512,N_5510);
xor U5981 (N_5981,N_5513,N_5528);
or U5982 (N_5982,N_5742,N_5740);
nand U5983 (N_5983,N_5708,N_5727);
nand U5984 (N_5984,N_5592,N_5594);
xnor U5985 (N_5985,N_5596,N_5648);
and U5986 (N_5986,N_5545,N_5565);
xnor U5987 (N_5987,N_5714,N_5509);
nor U5988 (N_5988,N_5615,N_5571);
nand U5989 (N_5989,N_5736,N_5656);
xnor U5990 (N_5990,N_5666,N_5715);
and U5991 (N_5991,N_5645,N_5712);
and U5992 (N_5992,N_5676,N_5527);
and U5993 (N_5993,N_5530,N_5732);
or U5994 (N_5994,N_5557,N_5529);
nor U5995 (N_5995,N_5609,N_5639);
or U5996 (N_5996,N_5678,N_5547);
nand U5997 (N_5997,N_5720,N_5633);
nor U5998 (N_5998,N_5748,N_5572);
or U5999 (N_5999,N_5644,N_5529);
nor U6000 (N_6000,N_5789,N_5775);
and U6001 (N_6001,N_5885,N_5995);
and U6002 (N_6002,N_5809,N_5982);
nand U6003 (N_6003,N_5968,N_5977);
nand U6004 (N_6004,N_5957,N_5847);
nand U6005 (N_6005,N_5931,N_5910);
nor U6006 (N_6006,N_5822,N_5973);
nand U6007 (N_6007,N_5853,N_5862);
nor U6008 (N_6008,N_5932,N_5793);
xor U6009 (N_6009,N_5859,N_5891);
or U6010 (N_6010,N_5949,N_5807);
or U6011 (N_6011,N_5941,N_5839);
nor U6012 (N_6012,N_5904,N_5796);
nor U6013 (N_6013,N_5780,N_5980);
xor U6014 (N_6014,N_5756,N_5886);
or U6015 (N_6015,N_5971,N_5769);
and U6016 (N_6016,N_5844,N_5909);
and U6017 (N_6017,N_5905,N_5959);
and U6018 (N_6018,N_5781,N_5843);
nor U6019 (N_6019,N_5820,N_5928);
xnor U6020 (N_6020,N_5837,N_5962);
or U6021 (N_6021,N_5933,N_5774);
xnor U6022 (N_6022,N_5879,N_5895);
nor U6023 (N_6023,N_5875,N_5892);
nor U6024 (N_6024,N_5950,N_5898);
nor U6025 (N_6025,N_5752,N_5947);
nand U6026 (N_6026,N_5848,N_5794);
nor U6027 (N_6027,N_5979,N_5758);
nand U6028 (N_6028,N_5825,N_5812);
xnor U6029 (N_6029,N_5930,N_5817);
xor U6030 (N_6030,N_5976,N_5896);
nor U6031 (N_6031,N_5911,N_5795);
or U6032 (N_6032,N_5906,N_5922);
nand U6033 (N_6033,N_5916,N_5923);
or U6034 (N_6034,N_5969,N_5926);
nand U6035 (N_6035,N_5924,N_5888);
nor U6036 (N_6036,N_5835,N_5763);
xnor U6037 (N_6037,N_5764,N_5889);
and U6038 (N_6038,N_5802,N_5967);
or U6039 (N_6039,N_5899,N_5983);
and U6040 (N_6040,N_5913,N_5773);
or U6041 (N_6041,N_5777,N_5818);
xor U6042 (N_6042,N_5944,N_5893);
nor U6043 (N_6043,N_5830,N_5877);
and U6044 (N_6044,N_5869,N_5804);
xor U6045 (N_6045,N_5964,N_5993);
nand U6046 (N_6046,N_5961,N_5801);
nor U6047 (N_6047,N_5841,N_5754);
or U6048 (N_6048,N_5782,N_5870);
xnor U6049 (N_6049,N_5988,N_5954);
nor U6050 (N_6050,N_5786,N_5824);
or U6051 (N_6051,N_5806,N_5936);
nor U6052 (N_6052,N_5890,N_5831);
or U6053 (N_6053,N_5978,N_5797);
and U6054 (N_6054,N_5943,N_5826);
xor U6055 (N_6055,N_5791,N_5760);
xnor U6056 (N_6056,N_5766,N_5884);
and U6057 (N_6057,N_5881,N_5914);
xnor U6058 (N_6058,N_5778,N_5813);
and U6059 (N_6059,N_5863,N_5985);
or U6060 (N_6060,N_5938,N_5960);
or U6061 (N_6061,N_5998,N_5838);
nor U6062 (N_6062,N_5920,N_5787);
or U6063 (N_6063,N_5942,N_5770);
and U6064 (N_6064,N_5987,N_5940);
nand U6065 (N_6065,N_5999,N_5846);
xnor U6066 (N_6066,N_5970,N_5965);
nor U6067 (N_6067,N_5955,N_5912);
nand U6068 (N_6068,N_5894,N_5832);
and U6069 (N_6069,N_5878,N_5819);
xor U6070 (N_6070,N_5811,N_5776);
nor U6071 (N_6071,N_5860,N_5919);
nor U6072 (N_6072,N_5972,N_5945);
nand U6073 (N_6073,N_5934,N_5966);
nand U6074 (N_6074,N_5784,N_5915);
nor U6075 (N_6075,N_5867,N_5779);
and U6076 (N_6076,N_5986,N_5814);
xor U6077 (N_6077,N_5921,N_5850);
and U6078 (N_6078,N_5883,N_5866);
or U6079 (N_6079,N_5753,N_5948);
or U6080 (N_6080,N_5935,N_5855);
and U6081 (N_6081,N_5992,N_5790);
xor U6082 (N_6082,N_5788,N_5974);
nand U6083 (N_6083,N_5808,N_5816);
or U6084 (N_6084,N_5887,N_5876);
xor U6085 (N_6085,N_5827,N_5792);
nand U6086 (N_6086,N_5865,N_5861);
nor U6087 (N_6087,N_5989,N_5842);
nand U6088 (N_6088,N_5901,N_5975);
nand U6089 (N_6089,N_5958,N_5907);
nand U6090 (N_6090,N_5925,N_5997);
and U6091 (N_6091,N_5840,N_5854);
nand U6092 (N_6092,N_5851,N_5810);
and U6093 (N_6093,N_5897,N_5902);
nor U6094 (N_6094,N_5852,N_5937);
xor U6095 (N_6095,N_5990,N_5917);
or U6096 (N_6096,N_5956,N_5761);
and U6097 (N_6097,N_5951,N_5903);
xnor U6098 (N_6098,N_5857,N_5805);
nor U6099 (N_6099,N_5864,N_5953);
and U6100 (N_6100,N_5880,N_5755);
nand U6101 (N_6101,N_5751,N_5759);
nor U6102 (N_6102,N_5849,N_5828);
and U6103 (N_6103,N_5994,N_5856);
nand U6104 (N_6104,N_5952,N_5946);
xor U6105 (N_6105,N_5836,N_5772);
xor U6106 (N_6106,N_5874,N_5783);
and U6107 (N_6107,N_5927,N_5963);
nand U6108 (N_6108,N_5929,N_5868);
or U6109 (N_6109,N_5871,N_5918);
or U6110 (N_6110,N_5762,N_5803);
and U6111 (N_6111,N_5981,N_5872);
xor U6112 (N_6112,N_5996,N_5984);
xor U6113 (N_6113,N_5882,N_5991);
and U6114 (N_6114,N_5757,N_5765);
nor U6115 (N_6115,N_5799,N_5873);
nand U6116 (N_6116,N_5829,N_5939);
or U6117 (N_6117,N_5908,N_5768);
xnor U6118 (N_6118,N_5823,N_5750);
or U6119 (N_6119,N_5785,N_5845);
or U6120 (N_6120,N_5834,N_5798);
xnor U6121 (N_6121,N_5767,N_5858);
nand U6122 (N_6122,N_5900,N_5815);
xnor U6123 (N_6123,N_5833,N_5800);
xnor U6124 (N_6124,N_5821,N_5771);
or U6125 (N_6125,N_5997,N_5923);
nand U6126 (N_6126,N_5954,N_5908);
nor U6127 (N_6127,N_5809,N_5930);
xnor U6128 (N_6128,N_5996,N_5874);
xor U6129 (N_6129,N_5786,N_5769);
xor U6130 (N_6130,N_5827,N_5785);
or U6131 (N_6131,N_5923,N_5880);
or U6132 (N_6132,N_5850,N_5904);
nor U6133 (N_6133,N_5851,N_5823);
or U6134 (N_6134,N_5945,N_5770);
nand U6135 (N_6135,N_5802,N_5951);
nand U6136 (N_6136,N_5915,N_5881);
nand U6137 (N_6137,N_5831,N_5901);
and U6138 (N_6138,N_5909,N_5846);
xnor U6139 (N_6139,N_5901,N_5962);
or U6140 (N_6140,N_5914,N_5851);
nor U6141 (N_6141,N_5783,N_5937);
nor U6142 (N_6142,N_5855,N_5797);
nor U6143 (N_6143,N_5983,N_5917);
or U6144 (N_6144,N_5833,N_5926);
xor U6145 (N_6145,N_5952,N_5759);
nand U6146 (N_6146,N_5955,N_5956);
nor U6147 (N_6147,N_5795,N_5943);
and U6148 (N_6148,N_5867,N_5968);
or U6149 (N_6149,N_5940,N_5773);
nand U6150 (N_6150,N_5871,N_5866);
nand U6151 (N_6151,N_5874,N_5943);
and U6152 (N_6152,N_5820,N_5817);
and U6153 (N_6153,N_5827,N_5778);
nand U6154 (N_6154,N_5962,N_5996);
or U6155 (N_6155,N_5757,N_5857);
nor U6156 (N_6156,N_5796,N_5845);
nand U6157 (N_6157,N_5968,N_5913);
and U6158 (N_6158,N_5866,N_5910);
and U6159 (N_6159,N_5764,N_5848);
and U6160 (N_6160,N_5878,N_5756);
and U6161 (N_6161,N_5960,N_5875);
xnor U6162 (N_6162,N_5978,N_5954);
and U6163 (N_6163,N_5751,N_5952);
or U6164 (N_6164,N_5954,N_5914);
or U6165 (N_6165,N_5795,N_5915);
nand U6166 (N_6166,N_5833,N_5902);
or U6167 (N_6167,N_5911,N_5945);
or U6168 (N_6168,N_5915,N_5964);
xnor U6169 (N_6169,N_5858,N_5892);
or U6170 (N_6170,N_5850,N_5874);
and U6171 (N_6171,N_5797,N_5839);
nor U6172 (N_6172,N_5950,N_5920);
nand U6173 (N_6173,N_5831,N_5961);
or U6174 (N_6174,N_5946,N_5882);
nand U6175 (N_6175,N_5922,N_5761);
xor U6176 (N_6176,N_5854,N_5871);
xnor U6177 (N_6177,N_5863,N_5819);
and U6178 (N_6178,N_5988,N_5870);
and U6179 (N_6179,N_5892,N_5759);
nand U6180 (N_6180,N_5858,N_5862);
or U6181 (N_6181,N_5978,N_5951);
nand U6182 (N_6182,N_5935,N_5863);
or U6183 (N_6183,N_5808,N_5798);
xnor U6184 (N_6184,N_5840,N_5842);
nand U6185 (N_6185,N_5890,N_5760);
xor U6186 (N_6186,N_5904,N_5815);
and U6187 (N_6187,N_5805,N_5864);
and U6188 (N_6188,N_5956,N_5865);
and U6189 (N_6189,N_5964,N_5793);
nand U6190 (N_6190,N_5854,N_5932);
or U6191 (N_6191,N_5769,N_5803);
xnor U6192 (N_6192,N_5853,N_5999);
nand U6193 (N_6193,N_5876,N_5909);
xor U6194 (N_6194,N_5929,N_5941);
nand U6195 (N_6195,N_5820,N_5784);
or U6196 (N_6196,N_5891,N_5977);
nand U6197 (N_6197,N_5944,N_5979);
nor U6198 (N_6198,N_5798,N_5976);
and U6199 (N_6199,N_5870,N_5871);
nor U6200 (N_6200,N_5875,N_5917);
and U6201 (N_6201,N_5856,N_5808);
and U6202 (N_6202,N_5826,N_5866);
and U6203 (N_6203,N_5979,N_5825);
and U6204 (N_6204,N_5987,N_5802);
nand U6205 (N_6205,N_5940,N_5844);
xnor U6206 (N_6206,N_5902,N_5845);
nand U6207 (N_6207,N_5904,N_5861);
and U6208 (N_6208,N_5804,N_5966);
xnor U6209 (N_6209,N_5927,N_5907);
and U6210 (N_6210,N_5886,N_5897);
or U6211 (N_6211,N_5815,N_5992);
nor U6212 (N_6212,N_5924,N_5918);
or U6213 (N_6213,N_5869,N_5846);
nor U6214 (N_6214,N_5985,N_5955);
xnor U6215 (N_6215,N_5845,N_5940);
or U6216 (N_6216,N_5874,N_5858);
nor U6217 (N_6217,N_5871,N_5892);
xnor U6218 (N_6218,N_5772,N_5800);
nor U6219 (N_6219,N_5849,N_5806);
and U6220 (N_6220,N_5765,N_5756);
nor U6221 (N_6221,N_5859,N_5980);
xor U6222 (N_6222,N_5876,N_5948);
or U6223 (N_6223,N_5987,N_5812);
or U6224 (N_6224,N_5822,N_5946);
xor U6225 (N_6225,N_5778,N_5759);
xor U6226 (N_6226,N_5893,N_5833);
xnor U6227 (N_6227,N_5862,N_5938);
nand U6228 (N_6228,N_5793,N_5947);
nor U6229 (N_6229,N_5818,N_5892);
or U6230 (N_6230,N_5782,N_5895);
nor U6231 (N_6231,N_5997,N_5828);
xor U6232 (N_6232,N_5878,N_5963);
or U6233 (N_6233,N_5926,N_5944);
xnor U6234 (N_6234,N_5776,N_5883);
nand U6235 (N_6235,N_5782,N_5754);
xnor U6236 (N_6236,N_5922,N_5769);
or U6237 (N_6237,N_5854,N_5993);
or U6238 (N_6238,N_5842,N_5950);
nor U6239 (N_6239,N_5976,N_5855);
nand U6240 (N_6240,N_5876,N_5873);
nand U6241 (N_6241,N_5903,N_5864);
or U6242 (N_6242,N_5945,N_5989);
xnor U6243 (N_6243,N_5755,N_5763);
nand U6244 (N_6244,N_5765,N_5973);
xor U6245 (N_6245,N_5938,N_5962);
nand U6246 (N_6246,N_5913,N_5791);
nor U6247 (N_6247,N_5917,N_5873);
xor U6248 (N_6248,N_5793,N_5769);
and U6249 (N_6249,N_5836,N_5873);
xor U6250 (N_6250,N_6158,N_6093);
and U6251 (N_6251,N_6052,N_6155);
and U6252 (N_6252,N_6121,N_6075);
nand U6253 (N_6253,N_6243,N_6110);
nor U6254 (N_6254,N_6101,N_6117);
and U6255 (N_6255,N_6216,N_6127);
xnor U6256 (N_6256,N_6061,N_6106);
or U6257 (N_6257,N_6193,N_6038);
nor U6258 (N_6258,N_6034,N_6004);
or U6259 (N_6259,N_6192,N_6051);
and U6260 (N_6260,N_6217,N_6103);
nand U6261 (N_6261,N_6073,N_6013);
or U6262 (N_6262,N_6238,N_6000);
nand U6263 (N_6263,N_6007,N_6149);
nand U6264 (N_6264,N_6125,N_6231);
nor U6265 (N_6265,N_6076,N_6249);
and U6266 (N_6266,N_6172,N_6197);
xnor U6267 (N_6267,N_6042,N_6150);
nor U6268 (N_6268,N_6186,N_6068);
nor U6269 (N_6269,N_6138,N_6078);
xnor U6270 (N_6270,N_6210,N_6119);
and U6271 (N_6271,N_6173,N_6129);
xnor U6272 (N_6272,N_6050,N_6234);
nor U6273 (N_6273,N_6136,N_6124);
or U6274 (N_6274,N_6229,N_6104);
nor U6275 (N_6275,N_6028,N_6220);
nor U6276 (N_6276,N_6091,N_6097);
and U6277 (N_6277,N_6037,N_6226);
xor U6278 (N_6278,N_6182,N_6139);
nand U6279 (N_6279,N_6159,N_6146);
xor U6280 (N_6280,N_6072,N_6089);
nand U6281 (N_6281,N_6026,N_6245);
nand U6282 (N_6282,N_6029,N_6137);
or U6283 (N_6283,N_6203,N_6005);
and U6284 (N_6284,N_6118,N_6165);
and U6285 (N_6285,N_6166,N_6200);
xnor U6286 (N_6286,N_6170,N_6211);
and U6287 (N_6287,N_6019,N_6001);
and U6288 (N_6288,N_6017,N_6080);
nand U6289 (N_6289,N_6223,N_6039);
nand U6290 (N_6290,N_6112,N_6087);
xnor U6291 (N_6291,N_6134,N_6218);
xor U6292 (N_6292,N_6088,N_6175);
nor U6293 (N_6293,N_6180,N_6070);
nand U6294 (N_6294,N_6053,N_6048);
or U6295 (N_6295,N_6135,N_6247);
nor U6296 (N_6296,N_6160,N_6188);
and U6297 (N_6297,N_6195,N_6108);
and U6298 (N_6298,N_6041,N_6140);
nor U6299 (N_6299,N_6151,N_6094);
nor U6300 (N_6300,N_6077,N_6233);
or U6301 (N_6301,N_6115,N_6027);
nor U6302 (N_6302,N_6126,N_6058);
and U6303 (N_6303,N_6095,N_6168);
nor U6304 (N_6304,N_6063,N_6036);
and U6305 (N_6305,N_6123,N_6147);
or U6306 (N_6306,N_6099,N_6107);
xor U6307 (N_6307,N_6128,N_6092);
nand U6308 (N_6308,N_6062,N_6246);
xnor U6309 (N_6309,N_6179,N_6020);
nor U6310 (N_6310,N_6012,N_6096);
or U6311 (N_6311,N_6171,N_6049);
nand U6312 (N_6312,N_6214,N_6174);
xor U6313 (N_6313,N_6157,N_6154);
xor U6314 (N_6314,N_6069,N_6225);
xor U6315 (N_6315,N_6145,N_6130);
or U6316 (N_6316,N_6178,N_6060);
or U6317 (N_6317,N_6116,N_6064);
and U6318 (N_6318,N_6105,N_6065);
nor U6319 (N_6319,N_6232,N_6066);
nand U6320 (N_6320,N_6240,N_6023);
nor U6321 (N_6321,N_6043,N_6224);
nand U6322 (N_6322,N_6142,N_6181);
nand U6323 (N_6323,N_6074,N_6006);
or U6324 (N_6324,N_6055,N_6040);
nand U6325 (N_6325,N_6212,N_6024);
and U6326 (N_6326,N_6194,N_6009);
and U6327 (N_6327,N_6114,N_6184);
xor U6328 (N_6328,N_6016,N_6098);
or U6329 (N_6329,N_6189,N_6241);
nand U6330 (N_6330,N_6067,N_6057);
nand U6331 (N_6331,N_6102,N_6011);
xnor U6332 (N_6332,N_6228,N_6236);
or U6333 (N_6333,N_6100,N_6230);
or U6334 (N_6334,N_6003,N_6071);
or U6335 (N_6335,N_6083,N_6046);
or U6336 (N_6336,N_6018,N_6082);
xnor U6337 (N_6337,N_6132,N_6190);
nand U6338 (N_6338,N_6152,N_6176);
xnor U6339 (N_6339,N_6219,N_6148);
and U6340 (N_6340,N_6208,N_6153);
nor U6341 (N_6341,N_6047,N_6109);
xor U6342 (N_6342,N_6035,N_6185);
xor U6343 (N_6343,N_6045,N_6222);
xor U6344 (N_6344,N_6221,N_6010);
xor U6345 (N_6345,N_6227,N_6086);
or U6346 (N_6346,N_6131,N_6025);
xor U6347 (N_6347,N_6161,N_6202);
or U6348 (N_6348,N_6059,N_6164);
or U6349 (N_6349,N_6133,N_6033);
nand U6350 (N_6350,N_6242,N_6177);
nand U6351 (N_6351,N_6213,N_6090);
xor U6352 (N_6352,N_6031,N_6022);
or U6353 (N_6353,N_6205,N_6002);
nor U6354 (N_6354,N_6162,N_6248);
or U6355 (N_6355,N_6244,N_6081);
xor U6356 (N_6356,N_6237,N_6191);
nor U6357 (N_6357,N_6206,N_6207);
nand U6358 (N_6358,N_6044,N_6156);
and U6359 (N_6359,N_6167,N_6032);
and U6360 (N_6360,N_6201,N_6183);
nand U6361 (N_6361,N_6143,N_6120);
xor U6362 (N_6362,N_6144,N_6209);
and U6363 (N_6363,N_6187,N_6014);
nand U6364 (N_6364,N_6198,N_6204);
or U6365 (N_6365,N_6239,N_6056);
nand U6366 (N_6366,N_6196,N_6111);
nand U6367 (N_6367,N_6079,N_6084);
xor U6368 (N_6368,N_6113,N_6054);
nor U6369 (N_6369,N_6021,N_6030);
or U6370 (N_6370,N_6163,N_6015);
nor U6371 (N_6371,N_6122,N_6169);
or U6372 (N_6372,N_6235,N_6215);
nand U6373 (N_6373,N_6085,N_6008);
nor U6374 (N_6374,N_6199,N_6141);
nand U6375 (N_6375,N_6057,N_6103);
xor U6376 (N_6376,N_6173,N_6171);
or U6377 (N_6377,N_6072,N_6226);
or U6378 (N_6378,N_6157,N_6054);
nor U6379 (N_6379,N_6150,N_6077);
nor U6380 (N_6380,N_6062,N_6032);
and U6381 (N_6381,N_6097,N_6036);
xnor U6382 (N_6382,N_6048,N_6069);
xor U6383 (N_6383,N_6172,N_6190);
nand U6384 (N_6384,N_6153,N_6110);
nor U6385 (N_6385,N_6095,N_6247);
and U6386 (N_6386,N_6227,N_6223);
nor U6387 (N_6387,N_6027,N_6220);
or U6388 (N_6388,N_6037,N_6094);
or U6389 (N_6389,N_6241,N_6091);
or U6390 (N_6390,N_6035,N_6081);
or U6391 (N_6391,N_6195,N_6213);
and U6392 (N_6392,N_6063,N_6119);
or U6393 (N_6393,N_6128,N_6140);
and U6394 (N_6394,N_6100,N_6143);
nand U6395 (N_6395,N_6230,N_6187);
nand U6396 (N_6396,N_6131,N_6106);
nand U6397 (N_6397,N_6132,N_6000);
or U6398 (N_6398,N_6222,N_6152);
or U6399 (N_6399,N_6146,N_6233);
and U6400 (N_6400,N_6226,N_6158);
nand U6401 (N_6401,N_6030,N_6234);
xor U6402 (N_6402,N_6207,N_6066);
or U6403 (N_6403,N_6020,N_6191);
or U6404 (N_6404,N_6094,N_6247);
and U6405 (N_6405,N_6112,N_6212);
and U6406 (N_6406,N_6065,N_6164);
xor U6407 (N_6407,N_6056,N_6123);
xnor U6408 (N_6408,N_6125,N_6068);
nor U6409 (N_6409,N_6004,N_6193);
xor U6410 (N_6410,N_6246,N_6108);
nand U6411 (N_6411,N_6206,N_6095);
nand U6412 (N_6412,N_6247,N_6077);
or U6413 (N_6413,N_6150,N_6182);
or U6414 (N_6414,N_6101,N_6162);
and U6415 (N_6415,N_6097,N_6154);
nand U6416 (N_6416,N_6232,N_6247);
nand U6417 (N_6417,N_6215,N_6163);
or U6418 (N_6418,N_6000,N_6026);
xnor U6419 (N_6419,N_6171,N_6133);
xnor U6420 (N_6420,N_6037,N_6085);
nand U6421 (N_6421,N_6031,N_6014);
or U6422 (N_6422,N_6099,N_6203);
or U6423 (N_6423,N_6216,N_6071);
and U6424 (N_6424,N_6158,N_6086);
xnor U6425 (N_6425,N_6039,N_6207);
nand U6426 (N_6426,N_6012,N_6124);
and U6427 (N_6427,N_6158,N_6214);
nand U6428 (N_6428,N_6201,N_6083);
and U6429 (N_6429,N_6016,N_6226);
xor U6430 (N_6430,N_6006,N_6093);
nor U6431 (N_6431,N_6065,N_6013);
and U6432 (N_6432,N_6149,N_6124);
and U6433 (N_6433,N_6202,N_6200);
nor U6434 (N_6434,N_6182,N_6092);
nor U6435 (N_6435,N_6155,N_6208);
nor U6436 (N_6436,N_6119,N_6019);
or U6437 (N_6437,N_6112,N_6033);
or U6438 (N_6438,N_6068,N_6175);
and U6439 (N_6439,N_6082,N_6065);
nor U6440 (N_6440,N_6072,N_6224);
or U6441 (N_6441,N_6232,N_6108);
nand U6442 (N_6442,N_6045,N_6243);
nand U6443 (N_6443,N_6081,N_6200);
and U6444 (N_6444,N_6249,N_6150);
xor U6445 (N_6445,N_6051,N_6246);
and U6446 (N_6446,N_6201,N_6101);
nor U6447 (N_6447,N_6223,N_6031);
nand U6448 (N_6448,N_6217,N_6133);
and U6449 (N_6449,N_6015,N_6012);
and U6450 (N_6450,N_6084,N_6222);
xor U6451 (N_6451,N_6242,N_6011);
and U6452 (N_6452,N_6215,N_6144);
and U6453 (N_6453,N_6145,N_6011);
nand U6454 (N_6454,N_6013,N_6086);
nand U6455 (N_6455,N_6153,N_6159);
xnor U6456 (N_6456,N_6063,N_6223);
nand U6457 (N_6457,N_6051,N_6081);
xnor U6458 (N_6458,N_6084,N_6135);
nand U6459 (N_6459,N_6175,N_6162);
xor U6460 (N_6460,N_6216,N_6052);
xnor U6461 (N_6461,N_6045,N_6065);
or U6462 (N_6462,N_6202,N_6192);
and U6463 (N_6463,N_6165,N_6100);
nand U6464 (N_6464,N_6080,N_6035);
nand U6465 (N_6465,N_6095,N_6087);
nand U6466 (N_6466,N_6237,N_6215);
and U6467 (N_6467,N_6107,N_6071);
nor U6468 (N_6468,N_6093,N_6108);
or U6469 (N_6469,N_6106,N_6229);
nor U6470 (N_6470,N_6072,N_6167);
nor U6471 (N_6471,N_6243,N_6203);
or U6472 (N_6472,N_6112,N_6049);
nor U6473 (N_6473,N_6106,N_6024);
xnor U6474 (N_6474,N_6134,N_6101);
nor U6475 (N_6475,N_6120,N_6049);
nand U6476 (N_6476,N_6228,N_6118);
and U6477 (N_6477,N_6127,N_6006);
nor U6478 (N_6478,N_6022,N_6020);
and U6479 (N_6479,N_6005,N_6201);
nor U6480 (N_6480,N_6148,N_6150);
nand U6481 (N_6481,N_6091,N_6123);
nor U6482 (N_6482,N_6103,N_6031);
nand U6483 (N_6483,N_6015,N_6232);
nor U6484 (N_6484,N_6180,N_6035);
or U6485 (N_6485,N_6005,N_6186);
nand U6486 (N_6486,N_6095,N_6246);
and U6487 (N_6487,N_6145,N_6080);
and U6488 (N_6488,N_6033,N_6169);
or U6489 (N_6489,N_6113,N_6046);
and U6490 (N_6490,N_6072,N_6018);
and U6491 (N_6491,N_6227,N_6040);
or U6492 (N_6492,N_6142,N_6220);
and U6493 (N_6493,N_6240,N_6184);
or U6494 (N_6494,N_6219,N_6194);
and U6495 (N_6495,N_6086,N_6029);
nand U6496 (N_6496,N_6034,N_6145);
xor U6497 (N_6497,N_6064,N_6092);
or U6498 (N_6498,N_6010,N_6156);
nand U6499 (N_6499,N_6076,N_6097);
nor U6500 (N_6500,N_6348,N_6364);
xor U6501 (N_6501,N_6442,N_6366);
nor U6502 (N_6502,N_6395,N_6378);
nor U6503 (N_6503,N_6339,N_6313);
nand U6504 (N_6504,N_6267,N_6338);
xor U6505 (N_6505,N_6477,N_6495);
and U6506 (N_6506,N_6493,N_6250);
or U6507 (N_6507,N_6490,N_6298);
nor U6508 (N_6508,N_6353,N_6406);
xnor U6509 (N_6509,N_6259,N_6371);
xnor U6510 (N_6510,N_6454,N_6380);
nand U6511 (N_6511,N_6296,N_6479);
xor U6512 (N_6512,N_6377,N_6285);
and U6513 (N_6513,N_6488,N_6476);
xnor U6514 (N_6514,N_6290,N_6438);
nor U6515 (N_6515,N_6398,N_6478);
xor U6516 (N_6516,N_6449,N_6459);
or U6517 (N_6517,N_6452,N_6425);
nand U6518 (N_6518,N_6391,N_6421);
nand U6519 (N_6519,N_6480,N_6357);
nor U6520 (N_6520,N_6458,N_6324);
or U6521 (N_6521,N_6263,N_6274);
nor U6522 (N_6522,N_6319,N_6356);
nand U6523 (N_6523,N_6289,N_6355);
nand U6524 (N_6524,N_6426,N_6292);
or U6525 (N_6525,N_6261,N_6389);
xor U6526 (N_6526,N_6360,N_6253);
nor U6527 (N_6527,N_6252,N_6288);
xor U6528 (N_6528,N_6270,N_6394);
or U6529 (N_6529,N_6419,N_6322);
or U6530 (N_6530,N_6434,N_6424);
xor U6531 (N_6531,N_6379,N_6260);
nand U6532 (N_6532,N_6472,N_6475);
nor U6533 (N_6533,N_6486,N_6436);
xnor U6534 (N_6534,N_6372,N_6496);
nor U6535 (N_6535,N_6325,N_6423);
nor U6536 (N_6536,N_6291,N_6315);
and U6537 (N_6537,N_6365,N_6310);
xor U6538 (N_6538,N_6441,N_6411);
nor U6539 (N_6539,N_6401,N_6376);
nor U6540 (N_6540,N_6402,N_6497);
nand U6541 (N_6541,N_6435,N_6382);
xnor U6542 (N_6542,N_6381,N_6418);
xnor U6543 (N_6543,N_6409,N_6273);
nand U6544 (N_6544,N_6400,N_6330);
and U6545 (N_6545,N_6404,N_6264);
and U6546 (N_6546,N_6331,N_6323);
and U6547 (N_6547,N_6427,N_6275);
nor U6548 (N_6548,N_6337,N_6386);
nor U6549 (N_6549,N_6284,N_6367);
nand U6550 (N_6550,N_6384,N_6336);
or U6551 (N_6551,N_6305,N_6368);
or U6552 (N_6552,N_6489,N_6299);
and U6553 (N_6553,N_6363,N_6326);
nor U6554 (N_6554,N_6347,N_6375);
xnor U6555 (N_6555,N_6450,N_6494);
nand U6556 (N_6556,N_6433,N_6370);
and U6557 (N_6557,N_6302,N_6446);
or U6558 (N_6558,N_6272,N_6388);
or U6559 (N_6559,N_6465,N_6440);
xnor U6560 (N_6560,N_6271,N_6354);
xor U6561 (N_6561,N_6445,N_6414);
xnor U6562 (N_6562,N_6278,N_6255);
nor U6563 (N_6563,N_6309,N_6460);
and U6564 (N_6564,N_6254,N_6349);
nand U6565 (N_6565,N_6361,N_6358);
nand U6566 (N_6566,N_6407,N_6374);
and U6567 (N_6567,N_6471,N_6469);
and U6568 (N_6568,N_6341,N_6399);
or U6569 (N_6569,N_6405,N_6464);
xor U6570 (N_6570,N_6327,N_6332);
nor U6571 (N_6571,N_6462,N_6487);
xnor U6572 (N_6572,N_6328,N_6457);
and U6573 (N_6573,N_6334,N_6373);
nor U6574 (N_6574,N_6258,N_6257);
and U6575 (N_6575,N_6320,N_6293);
xor U6576 (N_6576,N_6316,N_6413);
nor U6577 (N_6577,N_6467,N_6483);
nor U6578 (N_6578,N_6312,N_6306);
or U6579 (N_6579,N_6279,N_6453);
nor U6580 (N_6580,N_6422,N_6444);
and U6581 (N_6581,N_6256,N_6390);
and U6582 (N_6582,N_6432,N_6335);
or U6583 (N_6583,N_6437,N_6304);
or U6584 (N_6584,N_6383,N_6329);
and U6585 (N_6585,N_6342,N_6420);
nor U6586 (N_6586,N_6481,N_6351);
xnor U6587 (N_6587,N_6485,N_6403);
nor U6588 (N_6588,N_6340,N_6396);
xnor U6589 (N_6589,N_6268,N_6369);
nand U6590 (N_6590,N_6499,N_6468);
nor U6591 (N_6591,N_6287,N_6317);
nor U6592 (N_6592,N_6412,N_6393);
and U6593 (N_6593,N_6276,N_6294);
and U6594 (N_6594,N_6286,N_6301);
nor U6595 (N_6595,N_6482,N_6352);
nand U6596 (N_6596,N_6346,N_6429);
xor U6597 (N_6597,N_6303,N_6463);
or U6598 (N_6598,N_6308,N_6265);
nand U6599 (N_6599,N_6392,N_6456);
xor U6600 (N_6600,N_6461,N_6451);
nor U6601 (N_6601,N_6318,N_6344);
or U6602 (N_6602,N_6428,N_6295);
nor U6603 (N_6603,N_6417,N_6281);
and U6604 (N_6604,N_6498,N_6470);
or U6605 (N_6605,N_6416,N_6321);
xnor U6606 (N_6606,N_6359,N_6314);
or U6607 (N_6607,N_6455,N_6415);
and U6608 (N_6608,N_6473,N_6280);
nand U6609 (N_6609,N_6277,N_6474);
nor U6610 (N_6610,N_6283,N_6297);
xnor U6611 (N_6611,N_6266,N_6447);
xor U6612 (N_6612,N_6430,N_6387);
nand U6613 (N_6613,N_6343,N_6333);
nor U6614 (N_6614,N_6466,N_6443);
and U6615 (N_6615,N_6408,N_6350);
xnor U6616 (N_6616,N_6307,N_6345);
and U6617 (N_6617,N_6269,N_6397);
xor U6618 (N_6618,N_6262,N_6484);
and U6619 (N_6619,N_6439,N_6410);
and U6620 (N_6620,N_6311,N_6251);
nand U6621 (N_6621,N_6362,N_6448);
nand U6622 (N_6622,N_6431,N_6492);
nor U6623 (N_6623,N_6300,N_6282);
or U6624 (N_6624,N_6385,N_6491);
nand U6625 (N_6625,N_6297,N_6279);
and U6626 (N_6626,N_6377,N_6269);
xor U6627 (N_6627,N_6297,N_6364);
xor U6628 (N_6628,N_6344,N_6376);
nor U6629 (N_6629,N_6403,N_6346);
or U6630 (N_6630,N_6385,N_6416);
xnor U6631 (N_6631,N_6444,N_6483);
xnor U6632 (N_6632,N_6363,N_6485);
nor U6633 (N_6633,N_6492,N_6343);
and U6634 (N_6634,N_6266,N_6451);
and U6635 (N_6635,N_6496,N_6475);
xor U6636 (N_6636,N_6332,N_6375);
or U6637 (N_6637,N_6280,N_6467);
xnor U6638 (N_6638,N_6360,N_6343);
or U6639 (N_6639,N_6284,N_6253);
xnor U6640 (N_6640,N_6360,N_6317);
nand U6641 (N_6641,N_6334,N_6451);
nor U6642 (N_6642,N_6273,N_6326);
nand U6643 (N_6643,N_6480,N_6259);
or U6644 (N_6644,N_6466,N_6411);
and U6645 (N_6645,N_6364,N_6391);
or U6646 (N_6646,N_6256,N_6481);
nand U6647 (N_6647,N_6400,N_6283);
nand U6648 (N_6648,N_6441,N_6252);
nand U6649 (N_6649,N_6317,N_6368);
nor U6650 (N_6650,N_6487,N_6409);
or U6651 (N_6651,N_6266,N_6417);
xor U6652 (N_6652,N_6273,N_6368);
and U6653 (N_6653,N_6386,N_6484);
nor U6654 (N_6654,N_6482,N_6328);
nor U6655 (N_6655,N_6418,N_6285);
and U6656 (N_6656,N_6278,N_6262);
nand U6657 (N_6657,N_6339,N_6285);
xor U6658 (N_6658,N_6458,N_6276);
nand U6659 (N_6659,N_6334,N_6423);
and U6660 (N_6660,N_6420,N_6387);
or U6661 (N_6661,N_6494,N_6499);
xor U6662 (N_6662,N_6311,N_6385);
nor U6663 (N_6663,N_6475,N_6354);
nor U6664 (N_6664,N_6301,N_6336);
nand U6665 (N_6665,N_6418,N_6407);
and U6666 (N_6666,N_6403,N_6434);
and U6667 (N_6667,N_6417,N_6412);
xor U6668 (N_6668,N_6353,N_6308);
xor U6669 (N_6669,N_6429,N_6322);
nand U6670 (N_6670,N_6261,N_6485);
and U6671 (N_6671,N_6344,N_6343);
nor U6672 (N_6672,N_6302,N_6358);
or U6673 (N_6673,N_6367,N_6260);
and U6674 (N_6674,N_6488,N_6415);
and U6675 (N_6675,N_6342,N_6456);
or U6676 (N_6676,N_6252,N_6460);
and U6677 (N_6677,N_6451,N_6297);
and U6678 (N_6678,N_6469,N_6484);
or U6679 (N_6679,N_6251,N_6430);
nor U6680 (N_6680,N_6340,N_6409);
nor U6681 (N_6681,N_6277,N_6343);
nor U6682 (N_6682,N_6405,N_6305);
and U6683 (N_6683,N_6311,N_6475);
nor U6684 (N_6684,N_6350,N_6382);
xor U6685 (N_6685,N_6472,N_6364);
nor U6686 (N_6686,N_6496,N_6263);
nand U6687 (N_6687,N_6344,N_6499);
nand U6688 (N_6688,N_6325,N_6453);
nor U6689 (N_6689,N_6330,N_6452);
or U6690 (N_6690,N_6321,N_6314);
nor U6691 (N_6691,N_6273,N_6317);
xor U6692 (N_6692,N_6313,N_6255);
nor U6693 (N_6693,N_6280,N_6432);
nand U6694 (N_6694,N_6379,N_6382);
and U6695 (N_6695,N_6455,N_6459);
nand U6696 (N_6696,N_6353,N_6306);
nand U6697 (N_6697,N_6402,N_6477);
and U6698 (N_6698,N_6256,N_6363);
nand U6699 (N_6699,N_6326,N_6497);
or U6700 (N_6700,N_6415,N_6330);
nor U6701 (N_6701,N_6272,N_6413);
nor U6702 (N_6702,N_6254,N_6257);
or U6703 (N_6703,N_6293,N_6257);
xnor U6704 (N_6704,N_6384,N_6429);
nor U6705 (N_6705,N_6473,N_6322);
nor U6706 (N_6706,N_6381,N_6366);
nand U6707 (N_6707,N_6408,N_6487);
or U6708 (N_6708,N_6450,N_6389);
nor U6709 (N_6709,N_6256,N_6338);
xor U6710 (N_6710,N_6373,N_6386);
xnor U6711 (N_6711,N_6345,N_6314);
nor U6712 (N_6712,N_6272,N_6409);
nor U6713 (N_6713,N_6305,N_6460);
and U6714 (N_6714,N_6453,N_6379);
and U6715 (N_6715,N_6358,N_6258);
and U6716 (N_6716,N_6334,N_6458);
or U6717 (N_6717,N_6284,N_6414);
nand U6718 (N_6718,N_6337,N_6261);
or U6719 (N_6719,N_6289,N_6379);
nand U6720 (N_6720,N_6307,N_6499);
nand U6721 (N_6721,N_6400,N_6341);
and U6722 (N_6722,N_6466,N_6367);
and U6723 (N_6723,N_6465,N_6368);
nor U6724 (N_6724,N_6404,N_6484);
and U6725 (N_6725,N_6391,N_6429);
nand U6726 (N_6726,N_6251,N_6491);
nor U6727 (N_6727,N_6480,N_6428);
xor U6728 (N_6728,N_6251,N_6382);
nor U6729 (N_6729,N_6400,N_6358);
and U6730 (N_6730,N_6365,N_6434);
nor U6731 (N_6731,N_6476,N_6498);
nand U6732 (N_6732,N_6466,N_6253);
xnor U6733 (N_6733,N_6424,N_6291);
nand U6734 (N_6734,N_6487,N_6329);
or U6735 (N_6735,N_6382,N_6418);
and U6736 (N_6736,N_6268,N_6431);
or U6737 (N_6737,N_6331,N_6438);
or U6738 (N_6738,N_6333,N_6279);
xnor U6739 (N_6739,N_6301,N_6363);
and U6740 (N_6740,N_6393,N_6278);
nand U6741 (N_6741,N_6357,N_6290);
xnor U6742 (N_6742,N_6440,N_6470);
and U6743 (N_6743,N_6411,N_6392);
nor U6744 (N_6744,N_6336,N_6339);
nand U6745 (N_6745,N_6472,N_6340);
and U6746 (N_6746,N_6433,N_6389);
xnor U6747 (N_6747,N_6303,N_6453);
nor U6748 (N_6748,N_6454,N_6477);
nand U6749 (N_6749,N_6480,N_6443);
nor U6750 (N_6750,N_6732,N_6722);
and U6751 (N_6751,N_6544,N_6510);
and U6752 (N_6752,N_6681,N_6626);
and U6753 (N_6753,N_6589,N_6630);
nor U6754 (N_6754,N_6647,N_6598);
or U6755 (N_6755,N_6559,N_6620);
nor U6756 (N_6756,N_6508,N_6699);
xnor U6757 (N_6757,N_6608,N_6622);
nor U6758 (N_6758,N_6580,N_6616);
xnor U6759 (N_6759,N_6652,N_6542);
nor U6760 (N_6760,N_6605,N_6674);
nand U6761 (N_6761,N_6726,N_6554);
nor U6762 (N_6762,N_6507,N_6697);
or U6763 (N_6763,N_6635,N_6724);
or U6764 (N_6764,N_6685,N_6680);
or U6765 (N_6765,N_6617,N_6569);
nand U6766 (N_6766,N_6594,N_6541);
and U6767 (N_6767,N_6537,N_6684);
or U6768 (N_6768,N_6606,N_6659);
nor U6769 (N_6769,N_6624,N_6553);
or U6770 (N_6770,N_6528,N_6536);
or U6771 (N_6771,N_6702,N_6664);
or U6772 (N_6772,N_6566,N_6596);
and U6773 (N_6773,N_6698,N_6708);
xor U6774 (N_6774,N_6540,N_6695);
and U6775 (N_6775,N_6551,N_6637);
or U6776 (N_6776,N_6517,N_6648);
or U6777 (N_6777,N_6650,N_6646);
xor U6778 (N_6778,N_6714,N_6644);
or U6779 (N_6779,N_6511,N_6704);
nor U6780 (N_6780,N_6675,N_6607);
xnor U6781 (N_6781,N_6745,N_6671);
and U6782 (N_6782,N_6661,N_6656);
nand U6783 (N_6783,N_6666,N_6523);
xor U6784 (N_6784,N_6619,N_6518);
or U6785 (N_6785,N_6677,N_6582);
xor U6786 (N_6786,N_6513,N_6557);
nor U6787 (N_6787,N_6565,N_6627);
xor U6788 (N_6788,N_6590,N_6723);
nand U6789 (N_6789,N_6515,N_6602);
and U6790 (N_6790,N_6632,N_6678);
nor U6791 (N_6791,N_6641,N_6735);
and U6792 (N_6792,N_6501,N_6567);
or U6793 (N_6793,N_6509,N_6693);
and U6794 (N_6794,N_6526,N_6595);
or U6795 (N_6795,N_6625,N_6662);
xnor U6796 (N_6796,N_6690,N_6586);
or U6797 (N_6797,N_6728,N_6749);
nor U6798 (N_6798,N_6581,N_6663);
nor U6799 (N_6799,N_6547,N_6642);
xnor U6800 (N_6800,N_6700,N_6623);
xnor U6801 (N_6801,N_6657,N_6601);
nand U6802 (N_6802,N_6563,N_6731);
xor U6803 (N_6803,N_6585,N_6709);
xor U6804 (N_6804,N_6730,N_6592);
xnor U6805 (N_6805,N_6578,N_6711);
xnor U6806 (N_6806,N_6686,N_6670);
and U6807 (N_6807,N_6688,N_6621);
and U6808 (N_6808,N_6719,N_6548);
nor U6809 (N_6809,N_6747,N_6696);
nor U6810 (N_6810,N_6529,N_6733);
nand U6811 (N_6811,N_6527,N_6679);
nand U6812 (N_6812,N_6564,N_6505);
nor U6813 (N_6813,N_6612,N_6676);
nand U6814 (N_6814,N_6593,N_6654);
or U6815 (N_6815,N_6742,N_6524);
or U6816 (N_6816,N_6744,N_6737);
xor U6817 (N_6817,N_6614,N_6721);
nand U6818 (N_6818,N_6633,N_6504);
nand U6819 (N_6819,N_6734,N_6550);
or U6820 (N_6820,N_6568,N_6574);
nand U6821 (N_6821,N_6741,N_6532);
and U6822 (N_6822,N_6636,N_6748);
or U6823 (N_6823,N_6599,N_6613);
nor U6824 (N_6824,N_6672,N_6706);
or U6825 (N_6825,N_6716,N_6687);
xor U6826 (N_6826,N_6611,N_6555);
and U6827 (N_6827,N_6500,N_6655);
or U6828 (N_6828,N_6736,N_6502);
and U6829 (N_6829,N_6519,N_6600);
nor U6830 (N_6830,N_6558,N_6660);
nand U6831 (N_6831,N_6653,N_6571);
and U6832 (N_6832,N_6521,N_6673);
nor U6833 (N_6833,N_6514,N_6520);
or U6834 (N_6834,N_6552,N_6573);
xnor U6835 (N_6835,N_6597,N_6682);
xor U6836 (N_6836,N_6668,N_6603);
and U6837 (N_6837,N_6665,N_6651);
nand U6838 (N_6838,N_6538,N_6591);
nor U6839 (N_6839,N_6535,N_6579);
and U6840 (N_6840,N_6629,N_6530);
nand U6841 (N_6841,N_6584,N_6743);
or U6842 (N_6842,N_6587,N_6639);
nor U6843 (N_6843,N_6543,N_6705);
xnor U6844 (N_6844,N_6531,N_6707);
or U6845 (N_6845,N_6549,N_6583);
nand U6846 (N_6846,N_6522,N_6572);
nand U6847 (N_6847,N_6720,N_6746);
nor U6848 (N_6848,N_6539,N_6525);
xor U6849 (N_6849,N_6645,N_6576);
nand U6850 (N_6850,N_6588,N_6643);
xor U6851 (N_6851,N_6512,N_6718);
nor U6852 (N_6852,N_6667,N_6506);
nor U6853 (N_6853,N_6577,N_6715);
or U6854 (N_6854,N_6701,N_6609);
or U6855 (N_6855,N_6713,N_6727);
nor U6856 (N_6856,N_6546,N_6560);
nand U6857 (N_6857,N_6691,N_6649);
xor U6858 (N_6858,N_6631,N_6610);
or U6859 (N_6859,N_6615,N_6534);
and U6860 (N_6860,N_6692,N_6694);
xnor U6861 (N_6861,N_6561,N_6689);
or U6862 (N_6862,N_6729,N_6503);
and U6863 (N_6863,N_6628,N_6738);
xnor U6864 (N_6864,N_6710,N_6562);
nor U6865 (N_6865,N_6604,N_6740);
nand U6866 (N_6866,N_6516,N_6717);
and U6867 (N_6867,N_6739,N_6683);
xnor U6868 (N_6868,N_6638,N_6703);
nor U6869 (N_6869,N_6658,N_6533);
xor U6870 (N_6870,N_6556,N_6669);
xor U6871 (N_6871,N_6640,N_6634);
and U6872 (N_6872,N_6570,N_6618);
xor U6873 (N_6873,N_6725,N_6712);
nor U6874 (N_6874,N_6575,N_6545);
xor U6875 (N_6875,N_6534,N_6688);
nor U6876 (N_6876,N_6561,N_6600);
and U6877 (N_6877,N_6715,N_6619);
and U6878 (N_6878,N_6529,N_6504);
xnor U6879 (N_6879,N_6543,N_6724);
and U6880 (N_6880,N_6630,N_6550);
nor U6881 (N_6881,N_6560,N_6555);
nor U6882 (N_6882,N_6672,N_6680);
xnor U6883 (N_6883,N_6549,N_6569);
xnor U6884 (N_6884,N_6522,N_6710);
nand U6885 (N_6885,N_6743,N_6745);
or U6886 (N_6886,N_6724,N_6609);
nand U6887 (N_6887,N_6733,N_6547);
and U6888 (N_6888,N_6504,N_6551);
nand U6889 (N_6889,N_6562,N_6574);
nor U6890 (N_6890,N_6510,N_6528);
nor U6891 (N_6891,N_6529,N_6584);
or U6892 (N_6892,N_6656,N_6548);
xor U6893 (N_6893,N_6748,N_6613);
xor U6894 (N_6894,N_6593,N_6597);
xor U6895 (N_6895,N_6685,N_6569);
xnor U6896 (N_6896,N_6748,N_6701);
and U6897 (N_6897,N_6553,N_6586);
nor U6898 (N_6898,N_6714,N_6658);
or U6899 (N_6899,N_6534,N_6679);
or U6900 (N_6900,N_6703,N_6719);
nand U6901 (N_6901,N_6511,N_6738);
and U6902 (N_6902,N_6596,N_6578);
and U6903 (N_6903,N_6623,N_6648);
nand U6904 (N_6904,N_6676,N_6589);
and U6905 (N_6905,N_6593,N_6570);
and U6906 (N_6906,N_6540,N_6663);
and U6907 (N_6907,N_6621,N_6682);
nand U6908 (N_6908,N_6547,N_6624);
nand U6909 (N_6909,N_6707,N_6506);
xnor U6910 (N_6910,N_6588,N_6580);
or U6911 (N_6911,N_6566,N_6616);
nand U6912 (N_6912,N_6571,N_6563);
xor U6913 (N_6913,N_6519,N_6554);
nor U6914 (N_6914,N_6522,N_6698);
nor U6915 (N_6915,N_6595,N_6515);
xor U6916 (N_6916,N_6743,N_6738);
xnor U6917 (N_6917,N_6726,N_6562);
and U6918 (N_6918,N_6599,N_6747);
nand U6919 (N_6919,N_6563,N_6685);
nand U6920 (N_6920,N_6669,N_6672);
or U6921 (N_6921,N_6566,N_6559);
or U6922 (N_6922,N_6712,N_6666);
nand U6923 (N_6923,N_6720,N_6646);
nor U6924 (N_6924,N_6661,N_6555);
xor U6925 (N_6925,N_6546,N_6744);
xor U6926 (N_6926,N_6550,N_6593);
xor U6927 (N_6927,N_6653,N_6617);
nor U6928 (N_6928,N_6557,N_6673);
nor U6929 (N_6929,N_6665,N_6743);
xnor U6930 (N_6930,N_6720,N_6614);
nand U6931 (N_6931,N_6695,N_6675);
and U6932 (N_6932,N_6744,N_6696);
xnor U6933 (N_6933,N_6639,N_6633);
and U6934 (N_6934,N_6604,N_6670);
or U6935 (N_6935,N_6624,N_6702);
nand U6936 (N_6936,N_6746,N_6562);
and U6937 (N_6937,N_6736,N_6726);
and U6938 (N_6938,N_6579,N_6586);
and U6939 (N_6939,N_6690,N_6689);
nor U6940 (N_6940,N_6567,N_6653);
nor U6941 (N_6941,N_6533,N_6589);
nor U6942 (N_6942,N_6648,N_6516);
or U6943 (N_6943,N_6607,N_6541);
or U6944 (N_6944,N_6652,N_6650);
nand U6945 (N_6945,N_6736,N_6506);
and U6946 (N_6946,N_6564,N_6619);
and U6947 (N_6947,N_6702,N_6673);
nand U6948 (N_6948,N_6611,N_6700);
nand U6949 (N_6949,N_6583,N_6604);
xor U6950 (N_6950,N_6678,N_6578);
or U6951 (N_6951,N_6534,N_6620);
xnor U6952 (N_6952,N_6602,N_6725);
nor U6953 (N_6953,N_6633,N_6699);
nor U6954 (N_6954,N_6738,N_6647);
nand U6955 (N_6955,N_6609,N_6700);
nor U6956 (N_6956,N_6539,N_6597);
or U6957 (N_6957,N_6583,N_6703);
nand U6958 (N_6958,N_6511,N_6608);
xor U6959 (N_6959,N_6722,N_6671);
or U6960 (N_6960,N_6594,N_6534);
or U6961 (N_6961,N_6698,N_6524);
nor U6962 (N_6962,N_6520,N_6676);
and U6963 (N_6963,N_6695,N_6567);
xnor U6964 (N_6964,N_6631,N_6655);
xor U6965 (N_6965,N_6655,N_6718);
nor U6966 (N_6966,N_6651,N_6552);
nor U6967 (N_6967,N_6558,N_6645);
nand U6968 (N_6968,N_6610,N_6681);
or U6969 (N_6969,N_6705,N_6599);
xnor U6970 (N_6970,N_6523,N_6705);
or U6971 (N_6971,N_6517,N_6689);
or U6972 (N_6972,N_6524,N_6613);
xnor U6973 (N_6973,N_6744,N_6618);
nor U6974 (N_6974,N_6617,N_6674);
nor U6975 (N_6975,N_6659,N_6572);
xnor U6976 (N_6976,N_6572,N_6529);
nor U6977 (N_6977,N_6529,N_6592);
or U6978 (N_6978,N_6678,N_6728);
nand U6979 (N_6979,N_6554,N_6561);
nor U6980 (N_6980,N_6749,N_6621);
nand U6981 (N_6981,N_6709,N_6600);
nor U6982 (N_6982,N_6633,N_6561);
and U6983 (N_6983,N_6509,N_6680);
nand U6984 (N_6984,N_6677,N_6684);
nor U6985 (N_6985,N_6553,N_6743);
or U6986 (N_6986,N_6691,N_6695);
or U6987 (N_6987,N_6588,N_6675);
or U6988 (N_6988,N_6613,N_6672);
nor U6989 (N_6989,N_6568,N_6566);
nor U6990 (N_6990,N_6502,N_6507);
xor U6991 (N_6991,N_6548,N_6566);
nor U6992 (N_6992,N_6620,N_6557);
xnor U6993 (N_6993,N_6686,N_6749);
nand U6994 (N_6994,N_6560,N_6541);
nor U6995 (N_6995,N_6508,N_6622);
nor U6996 (N_6996,N_6656,N_6743);
and U6997 (N_6997,N_6640,N_6543);
or U6998 (N_6998,N_6517,N_6737);
xor U6999 (N_6999,N_6738,N_6599);
and U7000 (N_7000,N_6902,N_6912);
or U7001 (N_7001,N_6849,N_6751);
or U7002 (N_7002,N_6790,N_6783);
or U7003 (N_7003,N_6752,N_6908);
and U7004 (N_7004,N_6796,N_6981);
xor U7005 (N_7005,N_6788,N_6773);
xor U7006 (N_7006,N_6910,N_6924);
or U7007 (N_7007,N_6854,N_6915);
or U7008 (N_7008,N_6850,N_6944);
nor U7009 (N_7009,N_6866,N_6777);
and U7010 (N_7010,N_6918,N_6835);
nor U7011 (N_7011,N_6989,N_6757);
nand U7012 (N_7012,N_6846,N_6890);
xor U7013 (N_7013,N_6815,N_6807);
xnor U7014 (N_7014,N_6838,N_6802);
and U7015 (N_7015,N_6913,N_6909);
and U7016 (N_7016,N_6922,N_6960);
xor U7017 (N_7017,N_6855,N_6775);
nand U7018 (N_7018,N_6999,N_6889);
or U7019 (N_7019,N_6774,N_6950);
or U7020 (N_7020,N_6834,N_6929);
xor U7021 (N_7021,N_6977,N_6818);
or U7022 (N_7022,N_6776,N_6871);
xnor U7023 (N_7023,N_6853,N_6831);
and U7024 (N_7024,N_6847,N_6780);
or U7025 (N_7025,N_6794,N_6969);
and U7026 (N_7026,N_6819,N_6760);
or U7027 (N_7027,N_6856,N_6882);
xnor U7028 (N_7028,N_6933,N_6920);
nand U7029 (N_7029,N_6869,N_6958);
nand U7030 (N_7030,N_6753,N_6931);
nor U7031 (N_7031,N_6903,N_6984);
or U7032 (N_7032,N_6972,N_6945);
nor U7033 (N_7033,N_6892,N_6857);
xor U7034 (N_7034,N_6824,N_6928);
and U7035 (N_7035,N_6956,N_6822);
nor U7036 (N_7036,N_6916,N_6754);
or U7037 (N_7037,N_6859,N_6870);
or U7038 (N_7038,N_6820,N_6996);
nor U7039 (N_7039,N_6848,N_6957);
and U7040 (N_7040,N_6768,N_6755);
xor U7041 (N_7041,N_6888,N_6809);
nand U7042 (N_7042,N_6800,N_6940);
nor U7043 (N_7043,N_6875,N_6844);
and U7044 (N_7044,N_6836,N_6879);
xor U7045 (N_7045,N_6832,N_6821);
nand U7046 (N_7046,N_6979,N_6837);
and U7047 (N_7047,N_6826,N_6771);
nand U7048 (N_7048,N_6795,N_6936);
nand U7049 (N_7049,N_6954,N_6782);
xor U7050 (N_7050,N_6813,N_6978);
and U7051 (N_7051,N_6970,N_6860);
or U7052 (N_7052,N_6816,N_6986);
nor U7053 (N_7053,N_6914,N_6965);
xnor U7054 (N_7054,N_6982,N_6801);
xor U7055 (N_7055,N_6759,N_6939);
and U7056 (N_7056,N_6937,N_6943);
nor U7057 (N_7057,N_6948,N_6842);
nor U7058 (N_7058,N_6881,N_6803);
xor U7059 (N_7059,N_6865,N_6786);
nand U7060 (N_7060,N_6798,N_6907);
or U7061 (N_7061,N_6799,N_6787);
nor U7062 (N_7062,N_6906,N_6845);
nand U7063 (N_7063,N_6756,N_6806);
xor U7064 (N_7064,N_6961,N_6825);
nor U7065 (N_7065,N_6867,N_6941);
nor U7066 (N_7066,N_6827,N_6991);
and U7067 (N_7067,N_6963,N_6814);
nor U7068 (N_7068,N_6765,N_6952);
and U7069 (N_7069,N_6877,N_6810);
or U7070 (N_7070,N_6811,N_6898);
or U7071 (N_7071,N_6988,N_6926);
nand U7072 (N_7072,N_6885,N_6804);
and U7073 (N_7073,N_6829,N_6947);
nand U7074 (N_7074,N_6962,N_6993);
xnor U7075 (N_7075,N_6817,N_6925);
nor U7076 (N_7076,N_6942,N_6887);
nor U7077 (N_7077,N_6992,N_6919);
xor U7078 (N_7078,N_6935,N_6808);
xor U7079 (N_7079,N_6967,N_6784);
xor U7080 (N_7080,N_6873,N_6767);
or U7081 (N_7081,N_6964,N_6772);
and U7082 (N_7082,N_6861,N_6872);
nand U7083 (N_7083,N_6874,N_6823);
or U7084 (N_7084,N_6997,N_6949);
and U7085 (N_7085,N_6864,N_6959);
or U7086 (N_7086,N_6990,N_6900);
nor U7087 (N_7087,N_6770,N_6761);
or U7088 (N_7088,N_6901,N_6934);
or U7089 (N_7089,N_6778,N_6971);
and U7090 (N_7090,N_6841,N_6897);
nor U7091 (N_7091,N_6781,N_6797);
nor U7092 (N_7092,N_6975,N_6995);
and U7093 (N_7093,N_6880,N_6974);
or U7094 (N_7094,N_6828,N_6793);
or U7095 (N_7095,N_6805,N_6884);
xor U7096 (N_7096,N_6985,N_6868);
xor U7097 (N_7097,N_6750,N_6966);
nor U7098 (N_7098,N_6994,N_6953);
xnor U7099 (N_7099,N_6863,N_6764);
and U7100 (N_7100,N_6899,N_6973);
and U7101 (N_7101,N_6830,N_6792);
nor U7102 (N_7102,N_6785,N_6833);
nand U7103 (N_7103,N_6946,N_6758);
or U7104 (N_7104,N_6852,N_6923);
nand U7105 (N_7105,N_6904,N_6769);
or U7106 (N_7106,N_6894,N_6789);
nand U7107 (N_7107,N_6905,N_6862);
and U7108 (N_7108,N_6927,N_6911);
nand U7109 (N_7109,N_6951,N_6878);
xnor U7110 (N_7110,N_6976,N_6932);
xnor U7111 (N_7111,N_6762,N_6843);
or U7112 (N_7112,N_6779,N_6840);
or U7113 (N_7113,N_6886,N_6763);
and U7114 (N_7114,N_6791,N_6930);
or U7115 (N_7115,N_6766,N_6895);
xnor U7116 (N_7116,N_6955,N_6896);
nand U7117 (N_7117,N_6876,N_6839);
and U7118 (N_7118,N_6851,N_6917);
nor U7119 (N_7119,N_6858,N_6893);
or U7120 (N_7120,N_6938,N_6998);
nor U7121 (N_7121,N_6968,N_6980);
or U7122 (N_7122,N_6983,N_6921);
nand U7123 (N_7123,N_6891,N_6812);
nand U7124 (N_7124,N_6883,N_6987);
nor U7125 (N_7125,N_6904,N_6828);
and U7126 (N_7126,N_6944,N_6820);
nor U7127 (N_7127,N_6866,N_6765);
nand U7128 (N_7128,N_6903,N_6803);
xnor U7129 (N_7129,N_6821,N_6868);
xor U7130 (N_7130,N_6954,N_6842);
nand U7131 (N_7131,N_6904,N_6952);
nand U7132 (N_7132,N_6780,N_6752);
or U7133 (N_7133,N_6936,N_6875);
nand U7134 (N_7134,N_6994,N_6860);
nand U7135 (N_7135,N_6997,N_6829);
nor U7136 (N_7136,N_6861,N_6763);
nor U7137 (N_7137,N_6843,N_6947);
or U7138 (N_7138,N_6957,N_6934);
or U7139 (N_7139,N_6860,N_6756);
and U7140 (N_7140,N_6806,N_6940);
and U7141 (N_7141,N_6984,N_6785);
nor U7142 (N_7142,N_6947,N_6802);
xor U7143 (N_7143,N_6985,N_6993);
nor U7144 (N_7144,N_6883,N_6896);
nand U7145 (N_7145,N_6752,N_6787);
nor U7146 (N_7146,N_6984,N_6962);
or U7147 (N_7147,N_6916,N_6842);
nand U7148 (N_7148,N_6963,N_6887);
xnor U7149 (N_7149,N_6963,N_6940);
nand U7150 (N_7150,N_6901,N_6988);
and U7151 (N_7151,N_6900,N_6940);
nand U7152 (N_7152,N_6817,N_6770);
nor U7153 (N_7153,N_6843,N_6838);
nor U7154 (N_7154,N_6773,N_6820);
xor U7155 (N_7155,N_6872,N_6903);
xnor U7156 (N_7156,N_6779,N_6896);
and U7157 (N_7157,N_6918,N_6763);
and U7158 (N_7158,N_6848,N_6781);
and U7159 (N_7159,N_6872,N_6801);
and U7160 (N_7160,N_6940,N_6943);
and U7161 (N_7161,N_6877,N_6799);
nand U7162 (N_7162,N_6781,N_6989);
and U7163 (N_7163,N_6983,N_6886);
xnor U7164 (N_7164,N_6925,N_6845);
and U7165 (N_7165,N_6896,N_6771);
nand U7166 (N_7166,N_6824,N_6813);
and U7167 (N_7167,N_6994,N_6934);
and U7168 (N_7168,N_6899,N_6959);
or U7169 (N_7169,N_6990,N_6979);
nand U7170 (N_7170,N_6779,N_6764);
nor U7171 (N_7171,N_6860,N_6805);
xnor U7172 (N_7172,N_6894,N_6877);
nor U7173 (N_7173,N_6937,N_6851);
or U7174 (N_7174,N_6868,N_6755);
xnor U7175 (N_7175,N_6851,N_6862);
xnor U7176 (N_7176,N_6894,N_6820);
nor U7177 (N_7177,N_6807,N_6818);
nand U7178 (N_7178,N_6946,N_6996);
nor U7179 (N_7179,N_6947,N_6760);
nor U7180 (N_7180,N_6845,N_6867);
nor U7181 (N_7181,N_6786,N_6946);
nand U7182 (N_7182,N_6934,N_6834);
xnor U7183 (N_7183,N_6905,N_6783);
nor U7184 (N_7184,N_6908,N_6961);
nor U7185 (N_7185,N_6876,N_6913);
or U7186 (N_7186,N_6881,N_6795);
and U7187 (N_7187,N_6788,N_6764);
or U7188 (N_7188,N_6983,N_6766);
or U7189 (N_7189,N_6858,N_6913);
xor U7190 (N_7190,N_6852,N_6795);
xor U7191 (N_7191,N_6909,N_6862);
and U7192 (N_7192,N_6798,N_6868);
and U7193 (N_7193,N_6891,N_6956);
nand U7194 (N_7194,N_6910,N_6918);
xnor U7195 (N_7195,N_6996,N_6926);
or U7196 (N_7196,N_6800,N_6997);
xnor U7197 (N_7197,N_6862,N_6987);
or U7198 (N_7198,N_6780,N_6985);
xnor U7199 (N_7199,N_6964,N_6953);
or U7200 (N_7200,N_6958,N_6909);
nand U7201 (N_7201,N_6956,N_6996);
nor U7202 (N_7202,N_6901,N_6850);
xor U7203 (N_7203,N_6898,N_6940);
or U7204 (N_7204,N_6843,N_6892);
nand U7205 (N_7205,N_6939,N_6958);
xor U7206 (N_7206,N_6843,N_6801);
or U7207 (N_7207,N_6925,N_6751);
nand U7208 (N_7208,N_6848,N_6754);
nor U7209 (N_7209,N_6963,N_6900);
nor U7210 (N_7210,N_6990,N_6961);
or U7211 (N_7211,N_6810,N_6853);
or U7212 (N_7212,N_6906,N_6773);
nand U7213 (N_7213,N_6866,N_6954);
nor U7214 (N_7214,N_6938,N_6919);
or U7215 (N_7215,N_6914,N_6897);
xor U7216 (N_7216,N_6962,N_6841);
xor U7217 (N_7217,N_6815,N_6818);
nand U7218 (N_7218,N_6833,N_6858);
xnor U7219 (N_7219,N_6896,N_6953);
nand U7220 (N_7220,N_6791,N_6851);
nand U7221 (N_7221,N_6752,N_6792);
nor U7222 (N_7222,N_6862,N_6753);
nor U7223 (N_7223,N_6877,N_6833);
or U7224 (N_7224,N_6844,N_6837);
or U7225 (N_7225,N_6970,N_6823);
and U7226 (N_7226,N_6825,N_6821);
xnor U7227 (N_7227,N_6998,N_6804);
nand U7228 (N_7228,N_6845,N_6992);
xor U7229 (N_7229,N_6916,N_6750);
or U7230 (N_7230,N_6754,N_6898);
nand U7231 (N_7231,N_6949,N_6763);
xor U7232 (N_7232,N_6997,N_6802);
nor U7233 (N_7233,N_6914,N_6794);
and U7234 (N_7234,N_6822,N_6765);
or U7235 (N_7235,N_6836,N_6874);
nor U7236 (N_7236,N_6811,N_6928);
or U7237 (N_7237,N_6986,N_6851);
xor U7238 (N_7238,N_6872,N_6955);
xnor U7239 (N_7239,N_6808,N_6982);
xnor U7240 (N_7240,N_6954,N_6913);
nand U7241 (N_7241,N_6864,N_6851);
xor U7242 (N_7242,N_6819,N_6972);
nor U7243 (N_7243,N_6994,N_6851);
and U7244 (N_7244,N_6885,N_6914);
nor U7245 (N_7245,N_6881,N_6854);
xnor U7246 (N_7246,N_6858,N_6973);
xnor U7247 (N_7247,N_6979,N_6750);
nor U7248 (N_7248,N_6810,N_6826);
nor U7249 (N_7249,N_6938,N_6825);
or U7250 (N_7250,N_7149,N_7022);
or U7251 (N_7251,N_7024,N_7220);
nor U7252 (N_7252,N_7103,N_7215);
nand U7253 (N_7253,N_7240,N_7241);
xnor U7254 (N_7254,N_7042,N_7162);
xnor U7255 (N_7255,N_7067,N_7147);
nand U7256 (N_7256,N_7048,N_7237);
xnor U7257 (N_7257,N_7111,N_7191);
xor U7258 (N_7258,N_7221,N_7195);
and U7259 (N_7259,N_7193,N_7213);
or U7260 (N_7260,N_7112,N_7035);
and U7261 (N_7261,N_7157,N_7011);
xnor U7262 (N_7262,N_7141,N_7206);
nand U7263 (N_7263,N_7094,N_7093);
nor U7264 (N_7264,N_7085,N_7100);
nand U7265 (N_7265,N_7080,N_7090);
or U7266 (N_7266,N_7197,N_7102);
xnor U7267 (N_7267,N_7163,N_7124);
xor U7268 (N_7268,N_7155,N_7075);
or U7269 (N_7269,N_7010,N_7176);
or U7270 (N_7270,N_7228,N_7107);
or U7271 (N_7271,N_7079,N_7095);
or U7272 (N_7272,N_7236,N_7173);
nand U7273 (N_7273,N_7091,N_7232);
nor U7274 (N_7274,N_7072,N_7201);
xnor U7275 (N_7275,N_7226,N_7225);
and U7276 (N_7276,N_7105,N_7086);
and U7277 (N_7277,N_7019,N_7012);
and U7278 (N_7278,N_7152,N_7247);
and U7279 (N_7279,N_7199,N_7202);
nand U7280 (N_7280,N_7055,N_7205);
xnor U7281 (N_7281,N_7164,N_7222);
xor U7282 (N_7282,N_7229,N_7003);
and U7283 (N_7283,N_7006,N_7127);
nand U7284 (N_7284,N_7002,N_7170);
and U7285 (N_7285,N_7099,N_7243);
nand U7286 (N_7286,N_7101,N_7181);
and U7287 (N_7287,N_7119,N_7244);
and U7288 (N_7288,N_7078,N_7219);
and U7289 (N_7289,N_7023,N_7016);
or U7290 (N_7290,N_7144,N_7059);
nor U7291 (N_7291,N_7027,N_7177);
nor U7292 (N_7292,N_7097,N_7092);
xor U7293 (N_7293,N_7041,N_7005);
xor U7294 (N_7294,N_7039,N_7077);
nor U7295 (N_7295,N_7029,N_7212);
nand U7296 (N_7296,N_7131,N_7031);
and U7297 (N_7297,N_7040,N_7081);
and U7298 (N_7298,N_7200,N_7053);
and U7299 (N_7299,N_7187,N_7064);
nor U7300 (N_7300,N_7044,N_7110);
or U7301 (N_7301,N_7139,N_7113);
nor U7302 (N_7302,N_7218,N_7142);
nand U7303 (N_7303,N_7207,N_7179);
or U7304 (N_7304,N_7118,N_7037);
xor U7305 (N_7305,N_7242,N_7117);
xnor U7306 (N_7306,N_7061,N_7208);
xor U7307 (N_7307,N_7058,N_7125);
nand U7308 (N_7308,N_7194,N_7146);
xnor U7309 (N_7309,N_7216,N_7183);
or U7310 (N_7310,N_7180,N_7057);
xor U7311 (N_7311,N_7063,N_7030);
nand U7312 (N_7312,N_7234,N_7106);
nor U7313 (N_7313,N_7043,N_7128);
or U7314 (N_7314,N_7083,N_7231);
or U7315 (N_7315,N_7089,N_7135);
nor U7316 (N_7316,N_7096,N_7088);
and U7317 (N_7317,N_7188,N_7238);
nand U7318 (N_7318,N_7123,N_7013);
or U7319 (N_7319,N_7008,N_7084);
nor U7320 (N_7320,N_7069,N_7122);
nand U7321 (N_7321,N_7196,N_7174);
nand U7322 (N_7322,N_7115,N_7098);
nor U7323 (N_7323,N_7018,N_7223);
xor U7324 (N_7324,N_7120,N_7217);
and U7325 (N_7325,N_7049,N_7192);
or U7326 (N_7326,N_7026,N_7082);
and U7327 (N_7327,N_7121,N_7235);
nor U7328 (N_7328,N_7065,N_7038);
or U7329 (N_7329,N_7108,N_7066);
nand U7330 (N_7330,N_7143,N_7071);
and U7331 (N_7331,N_7116,N_7172);
and U7332 (N_7332,N_7000,N_7233);
nand U7333 (N_7333,N_7015,N_7004);
and U7334 (N_7334,N_7211,N_7129);
nand U7335 (N_7335,N_7045,N_7017);
and U7336 (N_7336,N_7070,N_7076);
xnor U7337 (N_7337,N_7150,N_7165);
nand U7338 (N_7338,N_7246,N_7214);
nand U7339 (N_7339,N_7209,N_7034);
nor U7340 (N_7340,N_7132,N_7136);
nor U7341 (N_7341,N_7148,N_7114);
nor U7342 (N_7342,N_7014,N_7198);
and U7343 (N_7343,N_7186,N_7073);
nand U7344 (N_7344,N_7052,N_7140);
or U7345 (N_7345,N_7060,N_7074);
and U7346 (N_7346,N_7166,N_7230);
xnor U7347 (N_7347,N_7046,N_7032);
and U7348 (N_7348,N_7134,N_7167);
or U7349 (N_7349,N_7068,N_7001);
and U7350 (N_7350,N_7227,N_7054);
or U7351 (N_7351,N_7007,N_7204);
nor U7352 (N_7352,N_7028,N_7009);
and U7353 (N_7353,N_7050,N_7190);
nand U7354 (N_7354,N_7145,N_7137);
and U7355 (N_7355,N_7189,N_7154);
xor U7356 (N_7356,N_7020,N_7160);
or U7357 (N_7357,N_7249,N_7175);
nor U7358 (N_7358,N_7104,N_7248);
xor U7359 (N_7359,N_7153,N_7130);
and U7360 (N_7360,N_7158,N_7178);
and U7361 (N_7361,N_7056,N_7087);
xnor U7362 (N_7362,N_7169,N_7036);
and U7363 (N_7363,N_7025,N_7185);
and U7364 (N_7364,N_7210,N_7156);
nor U7365 (N_7365,N_7161,N_7159);
nor U7366 (N_7366,N_7133,N_7182);
or U7367 (N_7367,N_7033,N_7171);
nand U7368 (N_7368,N_7126,N_7203);
nor U7369 (N_7369,N_7062,N_7047);
nor U7370 (N_7370,N_7109,N_7224);
nand U7371 (N_7371,N_7051,N_7239);
or U7372 (N_7372,N_7151,N_7138);
or U7373 (N_7373,N_7245,N_7184);
xor U7374 (N_7374,N_7168,N_7021);
nand U7375 (N_7375,N_7147,N_7219);
nand U7376 (N_7376,N_7111,N_7062);
xnor U7377 (N_7377,N_7153,N_7116);
nor U7378 (N_7378,N_7083,N_7149);
and U7379 (N_7379,N_7107,N_7012);
and U7380 (N_7380,N_7099,N_7030);
and U7381 (N_7381,N_7118,N_7196);
xor U7382 (N_7382,N_7051,N_7064);
or U7383 (N_7383,N_7174,N_7212);
xnor U7384 (N_7384,N_7208,N_7074);
nor U7385 (N_7385,N_7184,N_7169);
nor U7386 (N_7386,N_7051,N_7056);
nand U7387 (N_7387,N_7237,N_7197);
xor U7388 (N_7388,N_7075,N_7097);
and U7389 (N_7389,N_7032,N_7088);
and U7390 (N_7390,N_7237,N_7227);
xor U7391 (N_7391,N_7235,N_7100);
nor U7392 (N_7392,N_7151,N_7191);
xnor U7393 (N_7393,N_7245,N_7208);
xor U7394 (N_7394,N_7011,N_7112);
nand U7395 (N_7395,N_7015,N_7089);
nor U7396 (N_7396,N_7047,N_7136);
xnor U7397 (N_7397,N_7157,N_7230);
nor U7398 (N_7398,N_7216,N_7133);
or U7399 (N_7399,N_7079,N_7142);
nor U7400 (N_7400,N_7195,N_7048);
xor U7401 (N_7401,N_7028,N_7114);
or U7402 (N_7402,N_7029,N_7075);
or U7403 (N_7403,N_7099,N_7024);
and U7404 (N_7404,N_7178,N_7084);
or U7405 (N_7405,N_7093,N_7128);
nor U7406 (N_7406,N_7145,N_7080);
xnor U7407 (N_7407,N_7153,N_7018);
and U7408 (N_7408,N_7199,N_7121);
nor U7409 (N_7409,N_7169,N_7083);
nor U7410 (N_7410,N_7146,N_7161);
and U7411 (N_7411,N_7175,N_7164);
nand U7412 (N_7412,N_7140,N_7208);
xnor U7413 (N_7413,N_7091,N_7210);
nor U7414 (N_7414,N_7082,N_7137);
or U7415 (N_7415,N_7057,N_7225);
nand U7416 (N_7416,N_7179,N_7059);
nor U7417 (N_7417,N_7115,N_7035);
xnor U7418 (N_7418,N_7104,N_7212);
or U7419 (N_7419,N_7140,N_7023);
xnor U7420 (N_7420,N_7061,N_7205);
nand U7421 (N_7421,N_7109,N_7129);
xor U7422 (N_7422,N_7225,N_7163);
xor U7423 (N_7423,N_7003,N_7043);
nand U7424 (N_7424,N_7236,N_7131);
and U7425 (N_7425,N_7151,N_7157);
or U7426 (N_7426,N_7141,N_7169);
or U7427 (N_7427,N_7227,N_7182);
or U7428 (N_7428,N_7063,N_7014);
and U7429 (N_7429,N_7060,N_7048);
xor U7430 (N_7430,N_7017,N_7192);
xor U7431 (N_7431,N_7073,N_7196);
or U7432 (N_7432,N_7060,N_7176);
or U7433 (N_7433,N_7164,N_7242);
nand U7434 (N_7434,N_7248,N_7163);
nand U7435 (N_7435,N_7169,N_7010);
xor U7436 (N_7436,N_7181,N_7091);
nand U7437 (N_7437,N_7196,N_7012);
and U7438 (N_7438,N_7133,N_7206);
and U7439 (N_7439,N_7102,N_7029);
or U7440 (N_7440,N_7248,N_7136);
xnor U7441 (N_7441,N_7023,N_7193);
and U7442 (N_7442,N_7131,N_7055);
and U7443 (N_7443,N_7069,N_7011);
nor U7444 (N_7444,N_7192,N_7119);
nand U7445 (N_7445,N_7131,N_7147);
and U7446 (N_7446,N_7141,N_7190);
nand U7447 (N_7447,N_7144,N_7241);
and U7448 (N_7448,N_7073,N_7131);
or U7449 (N_7449,N_7051,N_7029);
nor U7450 (N_7450,N_7234,N_7049);
and U7451 (N_7451,N_7145,N_7239);
xor U7452 (N_7452,N_7229,N_7034);
or U7453 (N_7453,N_7057,N_7137);
nor U7454 (N_7454,N_7037,N_7066);
nand U7455 (N_7455,N_7062,N_7174);
xnor U7456 (N_7456,N_7212,N_7222);
xnor U7457 (N_7457,N_7087,N_7034);
xor U7458 (N_7458,N_7149,N_7142);
nor U7459 (N_7459,N_7098,N_7090);
or U7460 (N_7460,N_7002,N_7246);
or U7461 (N_7461,N_7194,N_7181);
xor U7462 (N_7462,N_7015,N_7157);
or U7463 (N_7463,N_7105,N_7043);
or U7464 (N_7464,N_7127,N_7176);
and U7465 (N_7465,N_7054,N_7214);
xnor U7466 (N_7466,N_7190,N_7133);
nor U7467 (N_7467,N_7081,N_7236);
xnor U7468 (N_7468,N_7020,N_7071);
or U7469 (N_7469,N_7138,N_7105);
nand U7470 (N_7470,N_7123,N_7161);
nand U7471 (N_7471,N_7102,N_7200);
nor U7472 (N_7472,N_7225,N_7010);
and U7473 (N_7473,N_7217,N_7181);
nand U7474 (N_7474,N_7211,N_7232);
or U7475 (N_7475,N_7095,N_7085);
xor U7476 (N_7476,N_7060,N_7146);
nand U7477 (N_7477,N_7220,N_7053);
and U7478 (N_7478,N_7244,N_7013);
or U7479 (N_7479,N_7192,N_7166);
xor U7480 (N_7480,N_7181,N_7207);
nand U7481 (N_7481,N_7008,N_7136);
and U7482 (N_7482,N_7063,N_7074);
and U7483 (N_7483,N_7034,N_7227);
nor U7484 (N_7484,N_7128,N_7097);
and U7485 (N_7485,N_7211,N_7072);
nor U7486 (N_7486,N_7131,N_7194);
and U7487 (N_7487,N_7177,N_7248);
or U7488 (N_7488,N_7055,N_7061);
nand U7489 (N_7489,N_7208,N_7233);
or U7490 (N_7490,N_7078,N_7186);
or U7491 (N_7491,N_7115,N_7028);
xor U7492 (N_7492,N_7139,N_7126);
or U7493 (N_7493,N_7054,N_7226);
or U7494 (N_7494,N_7043,N_7149);
nand U7495 (N_7495,N_7188,N_7185);
xor U7496 (N_7496,N_7162,N_7138);
xnor U7497 (N_7497,N_7009,N_7221);
xor U7498 (N_7498,N_7088,N_7202);
nand U7499 (N_7499,N_7147,N_7114);
xor U7500 (N_7500,N_7487,N_7350);
or U7501 (N_7501,N_7343,N_7328);
and U7502 (N_7502,N_7275,N_7490);
xor U7503 (N_7503,N_7498,N_7437);
or U7504 (N_7504,N_7379,N_7286);
and U7505 (N_7505,N_7363,N_7268);
xnor U7506 (N_7506,N_7340,N_7297);
nand U7507 (N_7507,N_7464,N_7494);
xor U7508 (N_7508,N_7351,N_7289);
nand U7509 (N_7509,N_7395,N_7489);
xor U7510 (N_7510,N_7336,N_7321);
xnor U7511 (N_7511,N_7406,N_7266);
or U7512 (N_7512,N_7305,N_7491);
or U7513 (N_7513,N_7307,N_7377);
nand U7514 (N_7514,N_7484,N_7454);
nand U7515 (N_7515,N_7356,N_7427);
and U7516 (N_7516,N_7346,N_7418);
nand U7517 (N_7517,N_7287,N_7369);
or U7518 (N_7518,N_7374,N_7326);
xnor U7519 (N_7519,N_7358,N_7252);
and U7520 (N_7520,N_7412,N_7482);
nand U7521 (N_7521,N_7315,N_7253);
xnor U7522 (N_7522,N_7388,N_7259);
nor U7523 (N_7523,N_7302,N_7338);
and U7524 (N_7524,N_7462,N_7345);
nand U7525 (N_7525,N_7308,N_7444);
and U7526 (N_7526,N_7257,N_7354);
nor U7527 (N_7527,N_7455,N_7389);
and U7528 (N_7528,N_7411,N_7323);
xnor U7529 (N_7529,N_7283,N_7399);
nor U7530 (N_7530,N_7263,N_7341);
nand U7531 (N_7531,N_7457,N_7443);
nor U7532 (N_7532,N_7276,N_7274);
xnor U7533 (N_7533,N_7471,N_7461);
or U7534 (N_7534,N_7265,N_7278);
nor U7535 (N_7535,N_7314,N_7474);
and U7536 (N_7536,N_7386,N_7292);
or U7537 (N_7537,N_7282,N_7367);
xnor U7538 (N_7538,N_7296,N_7415);
or U7539 (N_7539,N_7273,N_7331);
nand U7540 (N_7540,N_7322,N_7258);
xor U7541 (N_7541,N_7360,N_7256);
and U7542 (N_7542,N_7285,N_7353);
or U7543 (N_7543,N_7335,N_7352);
and U7544 (N_7544,N_7311,N_7410);
or U7545 (N_7545,N_7463,N_7365);
nor U7546 (N_7546,N_7277,N_7419);
and U7547 (N_7547,N_7378,N_7394);
and U7548 (N_7548,N_7324,N_7445);
xnor U7549 (N_7549,N_7486,N_7434);
or U7550 (N_7550,N_7425,N_7451);
xor U7551 (N_7551,N_7261,N_7327);
nor U7552 (N_7552,N_7312,N_7495);
xor U7553 (N_7553,N_7468,N_7480);
nor U7554 (N_7554,N_7404,N_7436);
nor U7555 (N_7555,N_7342,N_7272);
nand U7556 (N_7556,N_7349,N_7301);
nand U7557 (N_7557,N_7413,N_7403);
nand U7558 (N_7558,N_7250,N_7485);
and U7559 (N_7559,N_7381,N_7368);
nor U7560 (N_7560,N_7255,N_7458);
or U7561 (N_7561,N_7375,N_7251);
and U7562 (N_7562,N_7380,N_7447);
xor U7563 (N_7563,N_7361,N_7325);
nor U7564 (N_7564,N_7304,N_7370);
nor U7565 (N_7565,N_7392,N_7372);
or U7566 (N_7566,N_7478,N_7319);
nor U7567 (N_7567,N_7488,N_7313);
xnor U7568 (N_7568,N_7473,N_7357);
and U7569 (N_7569,N_7284,N_7267);
xor U7570 (N_7570,N_7429,N_7470);
xnor U7571 (N_7571,N_7280,N_7409);
nor U7572 (N_7572,N_7477,N_7481);
nor U7573 (N_7573,N_7387,N_7371);
nand U7574 (N_7574,N_7396,N_7294);
xnor U7575 (N_7575,N_7400,N_7414);
or U7576 (N_7576,N_7420,N_7408);
nand U7577 (N_7577,N_7422,N_7366);
nor U7578 (N_7578,N_7450,N_7448);
nand U7579 (N_7579,N_7337,N_7456);
xor U7580 (N_7580,N_7332,N_7339);
and U7581 (N_7581,N_7417,N_7497);
or U7582 (N_7582,N_7334,N_7475);
xnor U7583 (N_7583,N_7433,N_7303);
nor U7584 (N_7584,N_7320,N_7393);
xor U7585 (N_7585,N_7460,N_7431);
or U7586 (N_7586,N_7318,N_7279);
xnor U7587 (N_7587,N_7383,N_7452);
nor U7588 (N_7588,N_7359,N_7401);
and U7589 (N_7589,N_7439,N_7391);
and U7590 (N_7590,N_7344,N_7459);
nand U7591 (N_7591,N_7329,N_7330);
nand U7592 (N_7592,N_7428,N_7281);
nand U7593 (N_7593,N_7288,N_7309);
xor U7594 (N_7594,N_7446,N_7333);
nand U7595 (N_7595,N_7316,N_7469);
nand U7596 (N_7596,N_7269,N_7348);
nor U7597 (N_7597,N_7385,N_7493);
nand U7598 (N_7598,N_7432,N_7298);
nor U7599 (N_7599,N_7260,N_7483);
nor U7600 (N_7600,N_7466,N_7310);
or U7601 (N_7601,N_7438,N_7397);
and U7602 (N_7602,N_7496,N_7254);
nand U7603 (N_7603,N_7300,N_7421);
nor U7604 (N_7604,N_7476,N_7376);
and U7605 (N_7605,N_7364,N_7424);
nor U7606 (N_7606,N_7440,N_7373);
nor U7607 (N_7607,N_7416,N_7384);
xnor U7608 (N_7608,N_7355,N_7398);
and U7609 (N_7609,N_7347,N_7264);
nor U7610 (N_7610,N_7293,N_7435);
or U7611 (N_7611,N_7306,N_7492);
and U7612 (N_7612,N_7499,N_7270);
or U7613 (N_7613,N_7423,N_7295);
xnor U7614 (N_7614,N_7317,N_7362);
nor U7615 (N_7615,N_7390,N_7467);
or U7616 (N_7616,N_7402,N_7271);
nor U7617 (N_7617,N_7291,N_7407);
nand U7618 (N_7618,N_7479,N_7430);
xor U7619 (N_7619,N_7262,N_7299);
nor U7620 (N_7620,N_7290,N_7426);
and U7621 (N_7621,N_7453,N_7405);
nand U7622 (N_7622,N_7472,N_7465);
xor U7623 (N_7623,N_7441,N_7382);
and U7624 (N_7624,N_7449,N_7442);
xnor U7625 (N_7625,N_7421,N_7472);
and U7626 (N_7626,N_7433,N_7313);
nor U7627 (N_7627,N_7335,N_7299);
or U7628 (N_7628,N_7413,N_7416);
or U7629 (N_7629,N_7363,N_7353);
xor U7630 (N_7630,N_7426,N_7440);
or U7631 (N_7631,N_7432,N_7376);
xor U7632 (N_7632,N_7488,N_7465);
xor U7633 (N_7633,N_7351,N_7296);
or U7634 (N_7634,N_7271,N_7254);
or U7635 (N_7635,N_7340,N_7367);
xor U7636 (N_7636,N_7288,N_7395);
nor U7637 (N_7637,N_7398,N_7290);
and U7638 (N_7638,N_7437,N_7289);
nor U7639 (N_7639,N_7443,N_7392);
or U7640 (N_7640,N_7276,N_7370);
nor U7641 (N_7641,N_7414,N_7322);
nor U7642 (N_7642,N_7314,N_7453);
nor U7643 (N_7643,N_7443,N_7303);
nor U7644 (N_7644,N_7458,N_7424);
and U7645 (N_7645,N_7451,N_7320);
or U7646 (N_7646,N_7476,N_7429);
xnor U7647 (N_7647,N_7270,N_7343);
xor U7648 (N_7648,N_7330,N_7465);
nor U7649 (N_7649,N_7443,N_7480);
nand U7650 (N_7650,N_7462,N_7430);
nand U7651 (N_7651,N_7402,N_7299);
xor U7652 (N_7652,N_7333,N_7488);
nand U7653 (N_7653,N_7298,N_7338);
nand U7654 (N_7654,N_7480,N_7446);
xnor U7655 (N_7655,N_7419,N_7431);
nand U7656 (N_7656,N_7473,N_7372);
nor U7657 (N_7657,N_7326,N_7267);
and U7658 (N_7658,N_7380,N_7345);
and U7659 (N_7659,N_7449,N_7459);
nor U7660 (N_7660,N_7405,N_7346);
or U7661 (N_7661,N_7362,N_7346);
and U7662 (N_7662,N_7299,N_7462);
and U7663 (N_7663,N_7273,N_7485);
nand U7664 (N_7664,N_7440,N_7368);
nand U7665 (N_7665,N_7473,N_7286);
nor U7666 (N_7666,N_7321,N_7368);
or U7667 (N_7667,N_7288,N_7477);
nand U7668 (N_7668,N_7291,N_7449);
or U7669 (N_7669,N_7381,N_7471);
and U7670 (N_7670,N_7315,N_7272);
nand U7671 (N_7671,N_7313,N_7461);
nand U7672 (N_7672,N_7422,N_7335);
nor U7673 (N_7673,N_7359,N_7279);
xor U7674 (N_7674,N_7397,N_7421);
and U7675 (N_7675,N_7411,N_7327);
nand U7676 (N_7676,N_7315,N_7345);
and U7677 (N_7677,N_7488,N_7266);
nand U7678 (N_7678,N_7489,N_7429);
nor U7679 (N_7679,N_7376,N_7429);
xnor U7680 (N_7680,N_7257,N_7375);
nand U7681 (N_7681,N_7487,N_7439);
nand U7682 (N_7682,N_7359,N_7463);
nand U7683 (N_7683,N_7313,N_7274);
nand U7684 (N_7684,N_7378,N_7310);
nor U7685 (N_7685,N_7303,N_7305);
nand U7686 (N_7686,N_7434,N_7420);
nand U7687 (N_7687,N_7452,N_7345);
nor U7688 (N_7688,N_7270,N_7406);
or U7689 (N_7689,N_7345,N_7414);
nand U7690 (N_7690,N_7459,N_7418);
and U7691 (N_7691,N_7330,N_7397);
nand U7692 (N_7692,N_7469,N_7261);
or U7693 (N_7693,N_7261,N_7455);
or U7694 (N_7694,N_7253,N_7462);
or U7695 (N_7695,N_7300,N_7275);
or U7696 (N_7696,N_7491,N_7395);
or U7697 (N_7697,N_7348,N_7485);
or U7698 (N_7698,N_7378,N_7422);
nand U7699 (N_7699,N_7273,N_7251);
nand U7700 (N_7700,N_7313,N_7441);
nand U7701 (N_7701,N_7433,N_7251);
nand U7702 (N_7702,N_7370,N_7485);
nand U7703 (N_7703,N_7377,N_7445);
xor U7704 (N_7704,N_7368,N_7295);
nor U7705 (N_7705,N_7379,N_7351);
nor U7706 (N_7706,N_7273,N_7420);
nand U7707 (N_7707,N_7497,N_7439);
or U7708 (N_7708,N_7250,N_7404);
nor U7709 (N_7709,N_7486,N_7413);
nor U7710 (N_7710,N_7287,N_7390);
nor U7711 (N_7711,N_7310,N_7463);
or U7712 (N_7712,N_7484,N_7495);
nor U7713 (N_7713,N_7303,N_7415);
xor U7714 (N_7714,N_7459,N_7305);
nand U7715 (N_7715,N_7300,N_7496);
or U7716 (N_7716,N_7470,N_7393);
nor U7717 (N_7717,N_7456,N_7378);
nor U7718 (N_7718,N_7480,N_7334);
xnor U7719 (N_7719,N_7358,N_7486);
nor U7720 (N_7720,N_7380,N_7358);
xor U7721 (N_7721,N_7317,N_7455);
nand U7722 (N_7722,N_7390,N_7405);
nand U7723 (N_7723,N_7304,N_7433);
xor U7724 (N_7724,N_7344,N_7381);
nand U7725 (N_7725,N_7316,N_7367);
xnor U7726 (N_7726,N_7496,N_7311);
nand U7727 (N_7727,N_7381,N_7412);
nand U7728 (N_7728,N_7415,N_7384);
or U7729 (N_7729,N_7369,N_7278);
or U7730 (N_7730,N_7334,N_7327);
nand U7731 (N_7731,N_7344,N_7270);
nor U7732 (N_7732,N_7268,N_7318);
or U7733 (N_7733,N_7336,N_7365);
nor U7734 (N_7734,N_7344,N_7499);
xor U7735 (N_7735,N_7366,N_7445);
and U7736 (N_7736,N_7465,N_7387);
nor U7737 (N_7737,N_7488,N_7303);
and U7738 (N_7738,N_7465,N_7474);
and U7739 (N_7739,N_7419,N_7433);
nand U7740 (N_7740,N_7299,N_7482);
xor U7741 (N_7741,N_7401,N_7309);
and U7742 (N_7742,N_7365,N_7391);
xor U7743 (N_7743,N_7378,N_7353);
xnor U7744 (N_7744,N_7404,N_7398);
and U7745 (N_7745,N_7481,N_7438);
xor U7746 (N_7746,N_7256,N_7442);
xnor U7747 (N_7747,N_7445,N_7255);
nand U7748 (N_7748,N_7324,N_7406);
nor U7749 (N_7749,N_7428,N_7482);
xor U7750 (N_7750,N_7739,N_7733);
nor U7751 (N_7751,N_7563,N_7720);
or U7752 (N_7752,N_7725,N_7533);
nand U7753 (N_7753,N_7669,N_7741);
xnor U7754 (N_7754,N_7664,N_7527);
nor U7755 (N_7755,N_7514,N_7536);
and U7756 (N_7756,N_7510,N_7593);
or U7757 (N_7757,N_7690,N_7652);
nor U7758 (N_7758,N_7695,N_7608);
nand U7759 (N_7759,N_7526,N_7622);
and U7760 (N_7760,N_7645,N_7516);
nor U7761 (N_7761,N_7700,N_7687);
nand U7762 (N_7762,N_7512,N_7522);
or U7763 (N_7763,N_7542,N_7599);
or U7764 (N_7764,N_7618,N_7709);
and U7765 (N_7765,N_7619,N_7661);
and U7766 (N_7766,N_7578,N_7559);
or U7767 (N_7767,N_7565,N_7665);
nor U7768 (N_7768,N_7683,N_7705);
nand U7769 (N_7769,N_7631,N_7585);
and U7770 (N_7770,N_7576,N_7572);
xor U7771 (N_7771,N_7553,N_7701);
and U7772 (N_7772,N_7660,N_7505);
nand U7773 (N_7773,N_7630,N_7719);
nor U7774 (N_7774,N_7677,N_7688);
xnor U7775 (N_7775,N_7525,N_7580);
nand U7776 (N_7776,N_7551,N_7693);
and U7777 (N_7777,N_7646,N_7625);
and U7778 (N_7778,N_7515,N_7543);
and U7779 (N_7779,N_7714,N_7595);
nand U7780 (N_7780,N_7600,N_7513);
nand U7781 (N_7781,N_7518,N_7666);
or U7782 (N_7782,N_7567,N_7612);
or U7783 (N_7783,N_7623,N_7712);
or U7784 (N_7784,N_7636,N_7644);
nor U7785 (N_7785,N_7579,N_7744);
or U7786 (N_7786,N_7703,N_7570);
nor U7787 (N_7787,N_7606,N_7642);
nor U7788 (N_7788,N_7696,N_7633);
nand U7789 (N_7789,N_7562,N_7707);
xor U7790 (N_7790,N_7643,N_7564);
nor U7791 (N_7791,N_7745,N_7655);
nor U7792 (N_7792,N_7710,N_7603);
nor U7793 (N_7793,N_7508,N_7601);
nand U7794 (N_7794,N_7742,N_7651);
nand U7795 (N_7795,N_7632,N_7748);
and U7796 (N_7796,N_7596,N_7722);
nor U7797 (N_7797,N_7502,N_7503);
nand U7798 (N_7798,N_7523,N_7738);
nand U7799 (N_7799,N_7674,N_7587);
nand U7800 (N_7800,N_7684,N_7528);
or U7801 (N_7801,N_7620,N_7604);
or U7802 (N_7802,N_7629,N_7552);
and U7803 (N_7803,N_7500,N_7656);
nand U7804 (N_7804,N_7659,N_7548);
xor U7805 (N_7805,N_7511,N_7726);
nand U7806 (N_7806,N_7749,N_7718);
or U7807 (N_7807,N_7501,N_7546);
or U7808 (N_7808,N_7521,N_7544);
nand U7809 (N_7809,N_7734,N_7680);
xnor U7810 (N_7810,N_7694,N_7556);
nand U7811 (N_7811,N_7654,N_7713);
xor U7812 (N_7812,N_7716,N_7557);
nor U7813 (N_7813,N_7727,N_7624);
nor U7814 (N_7814,N_7535,N_7699);
nor U7815 (N_7815,N_7678,N_7628);
nand U7816 (N_7816,N_7594,N_7743);
xnor U7817 (N_7817,N_7532,N_7602);
and U7818 (N_7818,N_7747,N_7607);
xnor U7819 (N_7819,N_7673,N_7653);
nand U7820 (N_7820,N_7698,N_7592);
xnor U7821 (N_7821,N_7735,N_7702);
nor U7822 (N_7822,N_7638,N_7583);
or U7823 (N_7823,N_7547,N_7626);
nand U7824 (N_7824,N_7686,N_7611);
xnor U7825 (N_7825,N_7708,N_7724);
or U7826 (N_7826,N_7520,N_7537);
xor U7827 (N_7827,N_7697,N_7517);
nand U7828 (N_7828,N_7584,N_7641);
nor U7829 (N_7829,N_7617,N_7550);
nor U7830 (N_7830,N_7574,N_7715);
xor U7831 (N_7831,N_7635,N_7582);
xnor U7832 (N_7832,N_7706,N_7568);
xor U7833 (N_7833,N_7679,N_7692);
or U7834 (N_7834,N_7569,N_7627);
nor U7835 (N_7835,N_7598,N_7740);
nor U7836 (N_7836,N_7558,N_7621);
or U7837 (N_7837,N_7730,N_7682);
or U7838 (N_7838,N_7541,N_7614);
xnor U7839 (N_7839,N_7589,N_7723);
nor U7840 (N_7840,N_7507,N_7610);
xnor U7841 (N_7841,N_7615,N_7681);
or U7842 (N_7842,N_7650,N_7555);
nor U7843 (N_7843,N_7634,N_7605);
xor U7844 (N_7844,N_7721,N_7717);
or U7845 (N_7845,N_7529,N_7577);
xor U7846 (N_7846,N_7561,N_7581);
xnor U7847 (N_7847,N_7658,N_7524);
and U7848 (N_7848,N_7554,N_7663);
and U7849 (N_7849,N_7675,N_7647);
and U7850 (N_7850,N_7530,N_7609);
nand U7851 (N_7851,N_7731,N_7540);
nor U7852 (N_7852,N_7746,N_7616);
nor U7853 (N_7853,N_7685,N_7639);
xor U7854 (N_7854,N_7509,N_7591);
xnor U7855 (N_7855,N_7670,N_7597);
nor U7856 (N_7856,N_7649,N_7668);
nand U7857 (N_7857,N_7573,N_7560);
or U7858 (N_7858,N_7566,N_7691);
nor U7859 (N_7859,N_7671,N_7711);
or U7860 (N_7860,N_7539,N_7640);
nor U7861 (N_7861,N_7545,N_7504);
nor U7862 (N_7862,N_7531,N_7538);
nor U7863 (N_7863,N_7737,N_7672);
xnor U7864 (N_7864,N_7729,N_7590);
xor U7865 (N_7865,N_7736,N_7586);
nand U7866 (N_7866,N_7676,N_7662);
and U7867 (N_7867,N_7648,N_7657);
xor U7868 (N_7868,N_7728,N_7704);
nor U7869 (N_7869,N_7637,N_7732);
xnor U7870 (N_7870,N_7519,N_7689);
nand U7871 (N_7871,N_7571,N_7575);
xor U7872 (N_7872,N_7667,N_7506);
xor U7873 (N_7873,N_7588,N_7613);
nand U7874 (N_7874,N_7549,N_7534);
nand U7875 (N_7875,N_7564,N_7728);
xnor U7876 (N_7876,N_7654,N_7674);
or U7877 (N_7877,N_7644,N_7624);
xnor U7878 (N_7878,N_7664,N_7687);
xor U7879 (N_7879,N_7693,N_7549);
nand U7880 (N_7880,N_7523,N_7585);
nor U7881 (N_7881,N_7594,N_7551);
and U7882 (N_7882,N_7654,N_7672);
and U7883 (N_7883,N_7645,N_7600);
nand U7884 (N_7884,N_7671,N_7582);
and U7885 (N_7885,N_7731,N_7739);
or U7886 (N_7886,N_7685,N_7728);
nor U7887 (N_7887,N_7604,N_7586);
or U7888 (N_7888,N_7591,N_7557);
xor U7889 (N_7889,N_7744,N_7745);
and U7890 (N_7890,N_7540,N_7553);
nor U7891 (N_7891,N_7681,N_7561);
xor U7892 (N_7892,N_7526,N_7539);
and U7893 (N_7893,N_7579,N_7585);
xnor U7894 (N_7894,N_7501,N_7653);
or U7895 (N_7895,N_7712,N_7579);
or U7896 (N_7896,N_7595,N_7702);
xor U7897 (N_7897,N_7526,N_7746);
xor U7898 (N_7898,N_7553,N_7748);
and U7899 (N_7899,N_7612,N_7702);
nand U7900 (N_7900,N_7605,N_7508);
and U7901 (N_7901,N_7637,N_7600);
nand U7902 (N_7902,N_7590,N_7516);
or U7903 (N_7903,N_7604,N_7592);
xnor U7904 (N_7904,N_7610,N_7705);
and U7905 (N_7905,N_7731,N_7718);
nand U7906 (N_7906,N_7564,N_7657);
xnor U7907 (N_7907,N_7733,N_7591);
and U7908 (N_7908,N_7686,N_7709);
nor U7909 (N_7909,N_7692,N_7570);
and U7910 (N_7910,N_7719,N_7540);
and U7911 (N_7911,N_7591,N_7654);
xnor U7912 (N_7912,N_7693,N_7700);
nor U7913 (N_7913,N_7572,N_7548);
and U7914 (N_7914,N_7661,N_7679);
nand U7915 (N_7915,N_7566,N_7673);
or U7916 (N_7916,N_7607,N_7506);
and U7917 (N_7917,N_7697,N_7618);
nand U7918 (N_7918,N_7590,N_7647);
nor U7919 (N_7919,N_7711,N_7704);
nor U7920 (N_7920,N_7699,N_7722);
nand U7921 (N_7921,N_7714,N_7633);
nand U7922 (N_7922,N_7580,N_7513);
or U7923 (N_7923,N_7687,N_7564);
nor U7924 (N_7924,N_7560,N_7556);
xnor U7925 (N_7925,N_7504,N_7619);
nand U7926 (N_7926,N_7690,N_7657);
nand U7927 (N_7927,N_7696,N_7613);
or U7928 (N_7928,N_7583,N_7712);
or U7929 (N_7929,N_7709,N_7534);
and U7930 (N_7930,N_7672,N_7670);
nor U7931 (N_7931,N_7712,N_7555);
or U7932 (N_7932,N_7734,N_7673);
xnor U7933 (N_7933,N_7598,N_7664);
xor U7934 (N_7934,N_7522,N_7507);
nand U7935 (N_7935,N_7600,N_7687);
xnor U7936 (N_7936,N_7713,N_7516);
nand U7937 (N_7937,N_7606,N_7696);
nand U7938 (N_7938,N_7560,N_7727);
xor U7939 (N_7939,N_7635,N_7597);
nor U7940 (N_7940,N_7626,N_7553);
nor U7941 (N_7941,N_7533,N_7698);
nand U7942 (N_7942,N_7708,N_7550);
nand U7943 (N_7943,N_7729,N_7646);
and U7944 (N_7944,N_7558,N_7653);
or U7945 (N_7945,N_7518,N_7571);
and U7946 (N_7946,N_7675,N_7602);
xor U7947 (N_7947,N_7701,N_7544);
nand U7948 (N_7948,N_7567,N_7723);
nand U7949 (N_7949,N_7527,N_7608);
nor U7950 (N_7950,N_7614,N_7637);
and U7951 (N_7951,N_7691,N_7734);
and U7952 (N_7952,N_7558,N_7572);
nand U7953 (N_7953,N_7553,N_7529);
and U7954 (N_7954,N_7670,N_7605);
and U7955 (N_7955,N_7525,N_7557);
or U7956 (N_7956,N_7686,N_7541);
nor U7957 (N_7957,N_7537,N_7522);
nand U7958 (N_7958,N_7601,N_7609);
xor U7959 (N_7959,N_7678,N_7734);
xnor U7960 (N_7960,N_7695,N_7563);
xnor U7961 (N_7961,N_7651,N_7597);
or U7962 (N_7962,N_7521,N_7631);
nor U7963 (N_7963,N_7657,N_7655);
xor U7964 (N_7964,N_7689,N_7580);
nor U7965 (N_7965,N_7679,N_7723);
nand U7966 (N_7966,N_7570,N_7706);
nor U7967 (N_7967,N_7607,N_7662);
nand U7968 (N_7968,N_7643,N_7607);
or U7969 (N_7969,N_7658,N_7595);
xor U7970 (N_7970,N_7673,N_7725);
and U7971 (N_7971,N_7700,N_7510);
xnor U7972 (N_7972,N_7528,N_7614);
or U7973 (N_7973,N_7623,N_7664);
nand U7974 (N_7974,N_7651,N_7734);
or U7975 (N_7975,N_7615,N_7534);
nor U7976 (N_7976,N_7604,N_7723);
nor U7977 (N_7977,N_7567,N_7571);
and U7978 (N_7978,N_7715,N_7539);
or U7979 (N_7979,N_7707,N_7656);
or U7980 (N_7980,N_7655,N_7634);
nor U7981 (N_7981,N_7686,N_7694);
nor U7982 (N_7982,N_7722,N_7614);
xor U7983 (N_7983,N_7508,N_7562);
xnor U7984 (N_7984,N_7688,N_7570);
nand U7985 (N_7985,N_7661,N_7682);
and U7986 (N_7986,N_7635,N_7515);
nand U7987 (N_7987,N_7564,N_7641);
nand U7988 (N_7988,N_7650,N_7668);
nand U7989 (N_7989,N_7722,N_7540);
or U7990 (N_7990,N_7615,N_7501);
nor U7991 (N_7991,N_7628,N_7737);
nor U7992 (N_7992,N_7657,N_7516);
and U7993 (N_7993,N_7734,N_7517);
and U7994 (N_7994,N_7637,N_7585);
and U7995 (N_7995,N_7548,N_7730);
or U7996 (N_7996,N_7677,N_7518);
and U7997 (N_7997,N_7591,N_7517);
xnor U7998 (N_7998,N_7642,N_7714);
xor U7999 (N_7999,N_7652,N_7747);
or U8000 (N_8000,N_7857,N_7800);
xnor U8001 (N_8001,N_7779,N_7867);
nor U8002 (N_8002,N_7765,N_7823);
xnor U8003 (N_8003,N_7991,N_7829);
nand U8004 (N_8004,N_7752,N_7842);
and U8005 (N_8005,N_7882,N_7750);
and U8006 (N_8006,N_7903,N_7878);
or U8007 (N_8007,N_7845,N_7997);
xor U8008 (N_8008,N_7865,N_7944);
or U8009 (N_8009,N_7910,N_7898);
and U8010 (N_8010,N_7843,N_7858);
or U8011 (N_8011,N_7951,N_7978);
nand U8012 (N_8012,N_7848,N_7818);
or U8013 (N_8013,N_7837,N_7982);
or U8014 (N_8014,N_7941,N_7953);
xor U8015 (N_8015,N_7753,N_7912);
nor U8016 (N_8016,N_7851,N_7946);
and U8017 (N_8017,N_7854,N_7956);
nand U8018 (N_8018,N_7799,N_7899);
or U8019 (N_8019,N_7762,N_7985);
nor U8020 (N_8020,N_7841,N_7918);
nor U8021 (N_8021,N_7963,N_7862);
xnor U8022 (N_8022,N_7873,N_7785);
and U8023 (N_8023,N_7839,N_7846);
and U8024 (N_8024,N_7889,N_7988);
and U8025 (N_8025,N_7947,N_7817);
or U8026 (N_8026,N_7945,N_7916);
nor U8027 (N_8027,N_7776,N_7897);
nor U8028 (N_8028,N_7763,N_7900);
nand U8029 (N_8029,N_7879,N_7911);
or U8030 (N_8030,N_7754,N_7925);
nand U8031 (N_8031,N_7852,N_7774);
nand U8032 (N_8032,N_7801,N_7767);
nand U8033 (N_8033,N_7780,N_7964);
xor U8034 (N_8034,N_7870,N_7908);
and U8035 (N_8035,N_7836,N_7980);
nor U8036 (N_8036,N_7977,N_7827);
nand U8037 (N_8037,N_7772,N_7797);
nand U8038 (N_8038,N_7975,N_7995);
or U8039 (N_8039,N_7814,N_7933);
nand U8040 (N_8040,N_7810,N_7824);
nand U8041 (N_8041,N_7812,N_7955);
xor U8042 (N_8042,N_7914,N_7840);
nor U8043 (N_8043,N_7961,N_7808);
or U8044 (N_8044,N_7755,N_7969);
nor U8045 (N_8045,N_7877,N_7864);
and U8046 (N_8046,N_7771,N_7863);
xnor U8047 (N_8047,N_7819,N_7787);
nand U8048 (N_8048,N_7777,N_7850);
xnor U8049 (N_8049,N_7904,N_7815);
nand U8050 (N_8050,N_7883,N_7983);
nor U8051 (N_8051,N_7761,N_7935);
and U8052 (N_8052,N_7884,N_7805);
and U8053 (N_8053,N_7893,N_7793);
nor U8054 (N_8054,N_7902,N_7775);
and U8055 (N_8055,N_7838,N_7967);
or U8056 (N_8056,N_7920,N_7960);
and U8057 (N_8057,N_7913,N_7782);
xnor U8058 (N_8058,N_7751,N_7990);
nor U8059 (N_8059,N_7807,N_7943);
xnor U8060 (N_8060,N_7970,N_7923);
nand U8061 (N_8061,N_7968,N_7936);
xnor U8062 (N_8062,N_7756,N_7871);
nand U8063 (N_8063,N_7948,N_7804);
nor U8064 (N_8064,N_7950,N_7784);
nor U8065 (N_8065,N_7932,N_7887);
nor U8066 (N_8066,N_7981,N_7798);
nor U8067 (N_8067,N_7781,N_7766);
xor U8068 (N_8068,N_7994,N_7929);
nor U8069 (N_8069,N_7796,N_7821);
xor U8070 (N_8070,N_7986,N_7820);
or U8071 (N_8071,N_7949,N_7758);
nand U8072 (N_8072,N_7917,N_7965);
xor U8073 (N_8073,N_7874,N_7802);
nand U8074 (N_8074,N_7778,N_7919);
xnor U8075 (N_8075,N_7938,N_7895);
nand U8076 (N_8076,N_7973,N_7888);
nand U8077 (N_8077,N_7927,N_7795);
and U8078 (N_8078,N_7924,N_7987);
xnor U8079 (N_8079,N_7966,N_7816);
and U8080 (N_8080,N_7825,N_7789);
nand U8081 (N_8081,N_7834,N_7830);
nor U8082 (N_8082,N_7926,N_7764);
or U8083 (N_8083,N_7790,N_7849);
and U8084 (N_8084,N_7915,N_7826);
and U8085 (N_8085,N_7921,N_7868);
nor U8086 (N_8086,N_7783,N_7760);
or U8087 (N_8087,N_7835,N_7930);
nor U8088 (N_8088,N_7999,N_7939);
or U8089 (N_8089,N_7769,N_7832);
xnor U8090 (N_8090,N_7962,N_7768);
and U8091 (N_8091,N_7928,N_7869);
or U8092 (N_8092,N_7876,N_7892);
nor U8093 (N_8093,N_7940,N_7861);
and U8094 (N_8094,N_7979,N_7792);
and U8095 (N_8095,N_7909,N_7885);
or U8096 (N_8096,N_7880,N_7809);
xnor U8097 (N_8097,N_7993,N_7937);
nor U8098 (N_8098,N_7757,N_7803);
and U8099 (N_8099,N_7791,N_7976);
xnor U8100 (N_8100,N_7958,N_7859);
nor U8101 (N_8101,N_7992,N_7907);
and U8102 (N_8102,N_7984,N_7860);
nand U8103 (N_8103,N_7855,N_7847);
nand U8104 (N_8104,N_7794,N_7957);
xor U8105 (N_8105,N_7989,N_7813);
nand U8106 (N_8106,N_7856,N_7853);
and U8107 (N_8107,N_7931,N_7866);
nand U8108 (N_8108,N_7896,N_7786);
xnor U8109 (N_8109,N_7922,N_7806);
or U8110 (N_8110,N_7905,N_7954);
xnor U8111 (N_8111,N_7881,N_7788);
or U8112 (N_8112,N_7942,N_7759);
nor U8113 (N_8113,N_7872,N_7833);
nand U8114 (N_8114,N_7971,N_7770);
xnor U8115 (N_8115,N_7998,N_7901);
and U8116 (N_8116,N_7906,N_7822);
nor U8117 (N_8117,N_7773,N_7996);
and U8118 (N_8118,N_7831,N_7875);
or U8119 (N_8119,N_7974,N_7886);
nor U8120 (N_8120,N_7959,N_7952);
or U8121 (N_8121,N_7890,N_7828);
xor U8122 (N_8122,N_7972,N_7934);
xnor U8123 (N_8123,N_7811,N_7894);
nand U8124 (N_8124,N_7891,N_7844);
nor U8125 (N_8125,N_7915,N_7813);
or U8126 (N_8126,N_7879,N_7781);
or U8127 (N_8127,N_7890,N_7750);
or U8128 (N_8128,N_7997,N_7881);
xor U8129 (N_8129,N_7991,N_7877);
or U8130 (N_8130,N_7812,N_7782);
or U8131 (N_8131,N_7806,N_7863);
or U8132 (N_8132,N_7848,N_7962);
nor U8133 (N_8133,N_7931,N_7972);
xor U8134 (N_8134,N_7911,N_7853);
nand U8135 (N_8135,N_7872,N_7811);
xnor U8136 (N_8136,N_7816,N_7827);
xor U8137 (N_8137,N_7932,N_7985);
nor U8138 (N_8138,N_7938,N_7961);
and U8139 (N_8139,N_7977,N_7836);
nand U8140 (N_8140,N_7772,N_7970);
nand U8141 (N_8141,N_7999,N_7977);
or U8142 (N_8142,N_7937,N_7759);
and U8143 (N_8143,N_7765,N_7795);
nand U8144 (N_8144,N_7763,N_7859);
nor U8145 (N_8145,N_7963,N_7988);
or U8146 (N_8146,N_7962,N_7778);
nand U8147 (N_8147,N_7817,N_7792);
nor U8148 (N_8148,N_7784,N_7882);
nor U8149 (N_8149,N_7954,N_7846);
nand U8150 (N_8150,N_7794,N_7809);
nand U8151 (N_8151,N_7753,N_7836);
or U8152 (N_8152,N_7877,N_7968);
and U8153 (N_8153,N_7925,N_7903);
nor U8154 (N_8154,N_7914,N_7879);
nor U8155 (N_8155,N_7755,N_7835);
xor U8156 (N_8156,N_7994,N_7762);
nor U8157 (N_8157,N_7827,N_7998);
or U8158 (N_8158,N_7780,N_7992);
nand U8159 (N_8159,N_7771,N_7767);
xor U8160 (N_8160,N_7911,N_7842);
or U8161 (N_8161,N_7763,N_7916);
xnor U8162 (N_8162,N_7909,N_7981);
or U8163 (N_8163,N_7896,N_7937);
or U8164 (N_8164,N_7950,N_7808);
or U8165 (N_8165,N_7791,N_7948);
nor U8166 (N_8166,N_7861,N_7994);
nor U8167 (N_8167,N_7793,N_7979);
nand U8168 (N_8168,N_7947,N_7924);
and U8169 (N_8169,N_7823,N_7830);
nand U8170 (N_8170,N_7893,N_7810);
and U8171 (N_8171,N_7944,N_7959);
or U8172 (N_8172,N_7983,N_7991);
xor U8173 (N_8173,N_7800,N_7988);
xor U8174 (N_8174,N_7898,N_7801);
or U8175 (N_8175,N_7770,N_7782);
or U8176 (N_8176,N_7811,N_7984);
or U8177 (N_8177,N_7782,N_7850);
or U8178 (N_8178,N_7858,N_7810);
nor U8179 (N_8179,N_7870,N_7817);
nor U8180 (N_8180,N_7968,N_7853);
xor U8181 (N_8181,N_7999,N_7880);
nand U8182 (N_8182,N_7777,N_7797);
nand U8183 (N_8183,N_7971,N_7938);
xnor U8184 (N_8184,N_7996,N_7847);
nand U8185 (N_8185,N_7869,N_7972);
nand U8186 (N_8186,N_7860,N_7909);
or U8187 (N_8187,N_7944,N_7814);
or U8188 (N_8188,N_7862,N_7824);
xor U8189 (N_8189,N_7930,N_7811);
and U8190 (N_8190,N_7765,N_7961);
and U8191 (N_8191,N_7764,N_7959);
nor U8192 (N_8192,N_7874,N_7880);
nor U8193 (N_8193,N_7837,N_7890);
or U8194 (N_8194,N_7954,N_7889);
nor U8195 (N_8195,N_7851,N_7833);
xnor U8196 (N_8196,N_7888,N_7812);
and U8197 (N_8197,N_7866,N_7781);
and U8198 (N_8198,N_7990,N_7899);
and U8199 (N_8199,N_7889,N_7880);
or U8200 (N_8200,N_7803,N_7852);
and U8201 (N_8201,N_7973,N_7928);
nor U8202 (N_8202,N_7798,N_7763);
or U8203 (N_8203,N_7987,N_7896);
xor U8204 (N_8204,N_7859,N_7876);
and U8205 (N_8205,N_7987,N_7851);
nand U8206 (N_8206,N_7789,N_7890);
xor U8207 (N_8207,N_7758,N_7877);
nand U8208 (N_8208,N_7997,N_7964);
nand U8209 (N_8209,N_7997,N_7768);
nor U8210 (N_8210,N_7993,N_7887);
or U8211 (N_8211,N_7864,N_7807);
nor U8212 (N_8212,N_7953,N_7831);
nor U8213 (N_8213,N_7832,N_7787);
or U8214 (N_8214,N_7996,N_7981);
or U8215 (N_8215,N_7962,N_7797);
and U8216 (N_8216,N_7951,N_7874);
nor U8217 (N_8217,N_7837,N_7791);
nor U8218 (N_8218,N_7919,N_7989);
xor U8219 (N_8219,N_7761,N_7985);
or U8220 (N_8220,N_7986,N_7783);
nand U8221 (N_8221,N_7989,N_7811);
xor U8222 (N_8222,N_7955,N_7766);
or U8223 (N_8223,N_7909,N_7903);
xor U8224 (N_8224,N_7807,N_7849);
nor U8225 (N_8225,N_7834,N_7992);
nor U8226 (N_8226,N_7828,N_7761);
xnor U8227 (N_8227,N_7812,N_7956);
and U8228 (N_8228,N_7859,N_7990);
or U8229 (N_8229,N_7830,N_7923);
or U8230 (N_8230,N_7827,N_7987);
or U8231 (N_8231,N_7893,N_7766);
or U8232 (N_8232,N_7880,N_7771);
and U8233 (N_8233,N_7784,N_7873);
and U8234 (N_8234,N_7781,N_7817);
xnor U8235 (N_8235,N_7958,N_7903);
xor U8236 (N_8236,N_7944,N_7758);
or U8237 (N_8237,N_7969,N_7976);
and U8238 (N_8238,N_7942,N_7801);
and U8239 (N_8239,N_7954,N_7817);
and U8240 (N_8240,N_7876,N_7935);
nand U8241 (N_8241,N_7867,N_7994);
xnor U8242 (N_8242,N_7942,N_7795);
nand U8243 (N_8243,N_7867,N_7914);
nand U8244 (N_8244,N_7946,N_7824);
nor U8245 (N_8245,N_7820,N_7950);
xor U8246 (N_8246,N_7906,N_7840);
xor U8247 (N_8247,N_7874,N_7962);
xor U8248 (N_8248,N_7883,N_7834);
nor U8249 (N_8249,N_7758,N_7811);
nor U8250 (N_8250,N_8031,N_8076);
xnor U8251 (N_8251,N_8219,N_8059);
nand U8252 (N_8252,N_8021,N_8224);
nand U8253 (N_8253,N_8129,N_8081);
and U8254 (N_8254,N_8140,N_8045);
xor U8255 (N_8255,N_8092,N_8112);
nor U8256 (N_8256,N_8187,N_8157);
xor U8257 (N_8257,N_8223,N_8018);
nand U8258 (N_8258,N_8009,N_8134);
and U8259 (N_8259,N_8012,N_8124);
xor U8260 (N_8260,N_8028,N_8069);
or U8261 (N_8261,N_8054,N_8132);
nand U8262 (N_8262,N_8185,N_8207);
nor U8263 (N_8263,N_8068,N_8143);
nand U8264 (N_8264,N_8073,N_8195);
xnor U8265 (N_8265,N_8179,N_8024);
and U8266 (N_8266,N_8089,N_8145);
nand U8267 (N_8267,N_8019,N_8041);
xnor U8268 (N_8268,N_8171,N_8199);
and U8269 (N_8269,N_8096,N_8088);
nand U8270 (N_8270,N_8040,N_8232);
or U8271 (N_8271,N_8161,N_8177);
xnor U8272 (N_8272,N_8244,N_8015);
xor U8273 (N_8273,N_8033,N_8097);
nor U8274 (N_8274,N_8027,N_8101);
nand U8275 (N_8275,N_8078,N_8048);
xor U8276 (N_8276,N_8236,N_8052);
or U8277 (N_8277,N_8198,N_8065);
nand U8278 (N_8278,N_8020,N_8104);
xnor U8279 (N_8279,N_8102,N_8047);
and U8280 (N_8280,N_8062,N_8095);
and U8281 (N_8281,N_8010,N_8220);
or U8282 (N_8282,N_8231,N_8113);
and U8283 (N_8283,N_8154,N_8038);
xnor U8284 (N_8284,N_8135,N_8043);
nand U8285 (N_8285,N_8230,N_8148);
or U8286 (N_8286,N_8166,N_8123);
and U8287 (N_8287,N_8227,N_8082);
nor U8288 (N_8288,N_8007,N_8190);
xor U8289 (N_8289,N_8201,N_8079);
nand U8290 (N_8290,N_8246,N_8245);
nor U8291 (N_8291,N_8149,N_8165);
nand U8292 (N_8292,N_8050,N_8167);
or U8293 (N_8293,N_8049,N_8111);
and U8294 (N_8294,N_8013,N_8058);
nand U8295 (N_8295,N_8093,N_8211);
nand U8296 (N_8296,N_8042,N_8006);
nor U8297 (N_8297,N_8128,N_8011);
nor U8298 (N_8298,N_8130,N_8080);
nor U8299 (N_8299,N_8233,N_8127);
and U8300 (N_8300,N_8239,N_8215);
and U8301 (N_8301,N_8109,N_8032);
nor U8302 (N_8302,N_8114,N_8138);
or U8303 (N_8303,N_8036,N_8071);
and U8304 (N_8304,N_8151,N_8105);
nand U8305 (N_8305,N_8242,N_8213);
nand U8306 (N_8306,N_8182,N_8051);
and U8307 (N_8307,N_8221,N_8090);
and U8308 (N_8308,N_8086,N_8170);
and U8309 (N_8309,N_8248,N_8240);
nor U8310 (N_8310,N_8016,N_8172);
or U8311 (N_8311,N_8098,N_8204);
nor U8312 (N_8312,N_8053,N_8125);
and U8313 (N_8313,N_8162,N_8247);
nand U8314 (N_8314,N_8234,N_8175);
or U8315 (N_8315,N_8188,N_8064);
and U8316 (N_8316,N_8226,N_8160);
nand U8317 (N_8317,N_8137,N_8212);
nor U8318 (N_8318,N_8122,N_8196);
and U8319 (N_8319,N_8063,N_8243);
nor U8320 (N_8320,N_8200,N_8181);
or U8321 (N_8321,N_8099,N_8218);
xor U8322 (N_8322,N_8017,N_8115);
and U8323 (N_8323,N_8235,N_8110);
xor U8324 (N_8324,N_8003,N_8152);
nor U8325 (N_8325,N_8014,N_8202);
and U8326 (N_8326,N_8150,N_8156);
or U8327 (N_8327,N_8203,N_8084);
or U8328 (N_8328,N_8029,N_8026);
xnor U8329 (N_8329,N_8205,N_8142);
nor U8330 (N_8330,N_8023,N_8158);
xnor U8331 (N_8331,N_8008,N_8066);
and U8332 (N_8332,N_8168,N_8214);
or U8333 (N_8333,N_8210,N_8094);
nor U8334 (N_8334,N_8237,N_8163);
and U8335 (N_8335,N_8193,N_8209);
nor U8336 (N_8336,N_8136,N_8216);
xnor U8337 (N_8337,N_8189,N_8091);
xnor U8338 (N_8338,N_8060,N_8118);
and U8339 (N_8339,N_8222,N_8249);
nand U8340 (N_8340,N_8119,N_8035);
xnor U8341 (N_8341,N_8001,N_8169);
or U8342 (N_8342,N_8085,N_8192);
nor U8343 (N_8343,N_8139,N_8002);
nand U8344 (N_8344,N_8238,N_8141);
and U8345 (N_8345,N_8037,N_8004);
and U8346 (N_8346,N_8044,N_8184);
xor U8347 (N_8347,N_8133,N_8030);
or U8348 (N_8348,N_8106,N_8208);
nor U8349 (N_8349,N_8108,N_8159);
nand U8350 (N_8350,N_8180,N_8022);
or U8351 (N_8351,N_8146,N_8000);
and U8352 (N_8352,N_8072,N_8228);
nand U8353 (N_8353,N_8155,N_8075);
xor U8354 (N_8354,N_8057,N_8206);
nor U8355 (N_8355,N_8039,N_8178);
or U8356 (N_8356,N_8117,N_8191);
nand U8357 (N_8357,N_8087,N_8241);
nand U8358 (N_8358,N_8131,N_8194);
or U8359 (N_8359,N_8121,N_8153);
nand U8360 (N_8360,N_8103,N_8083);
nor U8361 (N_8361,N_8183,N_8025);
nand U8362 (N_8362,N_8077,N_8120);
and U8363 (N_8363,N_8217,N_8107);
nor U8364 (N_8364,N_8225,N_8174);
nand U8365 (N_8365,N_8074,N_8055);
xnor U8366 (N_8366,N_8067,N_8164);
xor U8367 (N_8367,N_8046,N_8056);
or U8368 (N_8368,N_8034,N_8173);
xnor U8369 (N_8369,N_8144,N_8061);
nor U8370 (N_8370,N_8229,N_8070);
nand U8371 (N_8371,N_8126,N_8186);
nand U8372 (N_8372,N_8100,N_8197);
xnor U8373 (N_8373,N_8147,N_8176);
nor U8374 (N_8374,N_8116,N_8005);
and U8375 (N_8375,N_8168,N_8037);
nor U8376 (N_8376,N_8002,N_8156);
or U8377 (N_8377,N_8182,N_8106);
nand U8378 (N_8378,N_8154,N_8111);
nor U8379 (N_8379,N_8013,N_8232);
xor U8380 (N_8380,N_8090,N_8117);
nor U8381 (N_8381,N_8086,N_8146);
xor U8382 (N_8382,N_8143,N_8037);
or U8383 (N_8383,N_8146,N_8149);
and U8384 (N_8384,N_8031,N_8025);
or U8385 (N_8385,N_8128,N_8126);
xnor U8386 (N_8386,N_8141,N_8199);
nor U8387 (N_8387,N_8231,N_8147);
and U8388 (N_8388,N_8154,N_8127);
nor U8389 (N_8389,N_8097,N_8125);
or U8390 (N_8390,N_8028,N_8203);
nand U8391 (N_8391,N_8152,N_8234);
and U8392 (N_8392,N_8014,N_8174);
and U8393 (N_8393,N_8124,N_8185);
nor U8394 (N_8394,N_8234,N_8181);
and U8395 (N_8395,N_8001,N_8003);
nor U8396 (N_8396,N_8007,N_8118);
and U8397 (N_8397,N_8227,N_8221);
nand U8398 (N_8398,N_8203,N_8026);
and U8399 (N_8399,N_8031,N_8085);
nor U8400 (N_8400,N_8245,N_8122);
xor U8401 (N_8401,N_8025,N_8234);
xnor U8402 (N_8402,N_8086,N_8178);
and U8403 (N_8403,N_8083,N_8130);
nor U8404 (N_8404,N_8097,N_8022);
xnor U8405 (N_8405,N_8007,N_8032);
or U8406 (N_8406,N_8116,N_8240);
and U8407 (N_8407,N_8243,N_8184);
xor U8408 (N_8408,N_8171,N_8172);
or U8409 (N_8409,N_8231,N_8134);
xnor U8410 (N_8410,N_8190,N_8131);
nor U8411 (N_8411,N_8230,N_8181);
nor U8412 (N_8412,N_8038,N_8045);
or U8413 (N_8413,N_8208,N_8076);
and U8414 (N_8414,N_8052,N_8102);
nor U8415 (N_8415,N_8147,N_8017);
and U8416 (N_8416,N_8138,N_8070);
xor U8417 (N_8417,N_8185,N_8248);
and U8418 (N_8418,N_8196,N_8223);
nand U8419 (N_8419,N_8021,N_8169);
or U8420 (N_8420,N_8110,N_8085);
or U8421 (N_8421,N_8061,N_8224);
xnor U8422 (N_8422,N_8166,N_8074);
nor U8423 (N_8423,N_8241,N_8091);
xor U8424 (N_8424,N_8173,N_8121);
xnor U8425 (N_8425,N_8246,N_8034);
nor U8426 (N_8426,N_8210,N_8056);
nand U8427 (N_8427,N_8059,N_8121);
or U8428 (N_8428,N_8004,N_8060);
nand U8429 (N_8429,N_8237,N_8206);
or U8430 (N_8430,N_8037,N_8241);
nor U8431 (N_8431,N_8039,N_8003);
and U8432 (N_8432,N_8013,N_8241);
and U8433 (N_8433,N_8107,N_8037);
and U8434 (N_8434,N_8010,N_8143);
and U8435 (N_8435,N_8222,N_8066);
or U8436 (N_8436,N_8216,N_8129);
xnor U8437 (N_8437,N_8101,N_8070);
and U8438 (N_8438,N_8196,N_8212);
or U8439 (N_8439,N_8112,N_8123);
nor U8440 (N_8440,N_8106,N_8094);
xnor U8441 (N_8441,N_8232,N_8011);
nor U8442 (N_8442,N_8106,N_8131);
or U8443 (N_8443,N_8141,N_8139);
nor U8444 (N_8444,N_8160,N_8089);
nand U8445 (N_8445,N_8021,N_8210);
nor U8446 (N_8446,N_8136,N_8075);
nand U8447 (N_8447,N_8177,N_8112);
nand U8448 (N_8448,N_8159,N_8187);
xnor U8449 (N_8449,N_8106,N_8069);
or U8450 (N_8450,N_8228,N_8076);
and U8451 (N_8451,N_8004,N_8239);
or U8452 (N_8452,N_8041,N_8122);
nor U8453 (N_8453,N_8109,N_8020);
nand U8454 (N_8454,N_8135,N_8067);
and U8455 (N_8455,N_8244,N_8086);
nor U8456 (N_8456,N_8180,N_8228);
or U8457 (N_8457,N_8142,N_8211);
and U8458 (N_8458,N_8088,N_8191);
xnor U8459 (N_8459,N_8210,N_8036);
nor U8460 (N_8460,N_8179,N_8204);
xor U8461 (N_8461,N_8078,N_8047);
xor U8462 (N_8462,N_8185,N_8194);
or U8463 (N_8463,N_8022,N_8161);
and U8464 (N_8464,N_8155,N_8077);
and U8465 (N_8465,N_8084,N_8202);
xor U8466 (N_8466,N_8216,N_8083);
or U8467 (N_8467,N_8030,N_8249);
nor U8468 (N_8468,N_8164,N_8036);
xor U8469 (N_8469,N_8057,N_8150);
xor U8470 (N_8470,N_8039,N_8172);
and U8471 (N_8471,N_8080,N_8067);
and U8472 (N_8472,N_8164,N_8119);
nor U8473 (N_8473,N_8139,N_8178);
and U8474 (N_8474,N_8167,N_8168);
or U8475 (N_8475,N_8082,N_8067);
or U8476 (N_8476,N_8219,N_8146);
nand U8477 (N_8477,N_8106,N_8217);
or U8478 (N_8478,N_8103,N_8021);
nor U8479 (N_8479,N_8007,N_8101);
and U8480 (N_8480,N_8217,N_8183);
xor U8481 (N_8481,N_8092,N_8234);
nand U8482 (N_8482,N_8199,N_8105);
xor U8483 (N_8483,N_8183,N_8242);
nand U8484 (N_8484,N_8081,N_8082);
or U8485 (N_8485,N_8169,N_8220);
and U8486 (N_8486,N_8166,N_8020);
xor U8487 (N_8487,N_8213,N_8186);
xor U8488 (N_8488,N_8211,N_8241);
or U8489 (N_8489,N_8079,N_8129);
and U8490 (N_8490,N_8000,N_8159);
nor U8491 (N_8491,N_8133,N_8022);
nand U8492 (N_8492,N_8001,N_8081);
and U8493 (N_8493,N_8142,N_8063);
and U8494 (N_8494,N_8142,N_8165);
or U8495 (N_8495,N_8153,N_8235);
or U8496 (N_8496,N_8103,N_8178);
and U8497 (N_8497,N_8185,N_8011);
nand U8498 (N_8498,N_8152,N_8157);
xnor U8499 (N_8499,N_8005,N_8053);
xor U8500 (N_8500,N_8302,N_8464);
nor U8501 (N_8501,N_8262,N_8462);
xor U8502 (N_8502,N_8398,N_8466);
nor U8503 (N_8503,N_8424,N_8475);
and U8504 (N_8504,N_8470,N_8385);
or U8505 (N_8505,N_8368,N_8279);
or U8506 (N_8506,N_8371,N_8311);
nand U8507 (N_8507,N_8375,N_8281);
or U8508 (N_8508,N_8253,N_8408);
nand U8509 (N_8509,N_8312,N_8482);
nor U8510 (N_8510,N_8391,N_8294);
nand U8511 (N_8511,N_8357,N_8359);
nand U8512 (N_8512,N_8303,N_8372);
xnor U8513 (N_8513,N_8492,N_8423);
and U8514 (N_8514,N_8386,N_8373);
nand U8515 (N_8515,N_8333,N_8257);
nor U8516 (N_8516,N_8336,N_8293);
xor U8517 (N_8517,N_8439,N_8277);
nand U8518 (N_8518,N_8289,N_8345);
and U8519 (N_8519,N_8347,N_8494);
or U8520 (N_8520,N_8282,N_8477);
xnor U8521 (N_8521,N_8271,N_8425);
nand U8522 (N_8522,N_8348,N_8411);
nor U8523 (N_8523,N_8396,N_8432);
and U8524 (N_8524,N_8451,N_8445);
xnor U8525 (N_8525,N_8453,N_8319);
or U8526 (N_8526,N_8321,N_8349);
or U8527 (N_8527,N_8484,N_8363);
nand U8528 (N_8528,N_8285,N_8463);
xnor U8529 (N_8529,N_8374,N_8370);
nor U8530 (N_8530,N_8471,N_8428);
xor U8531 (N_8531,N_8338,N_8387);
and U8532 (N_8532,N_8360,N_8328);
or U8533 (N_8533,N_8269,N_8365);
xnor U8534 (N_8534,N_8409,N_8326);
xor U8535 (N_8535,N_8358,N_8459);
or U8536 (N_8536,N_8317,N_8329);
or U8537 (N_8537,N_8497,N_8255);
and U8538 (N_8538,N_8342,N_8467);
xnor U8539 (N_8539,N_8498,N_8456);
xnor U8540 (N_8540,N_8272,N_8320);
or U8541 (N_8541,N_8399,N_8256);
nor U8542 (N_8542,N_8378,N_8380);
nor U8543 (N_8543,N_8313,N_8297);
nor U8544 (N_8544,N_8413,N_8406);
and U8545 (N_8545,N_8325,N_8286);
xnor U8546 (N_8546,N_8496,N_8487);
nor U8547 (N_8547,N_8438,N_8404);
nand U8548 (N_8548,N_8437,N_8377);
nand U8549 (N_8549,N_8383,N_8280);
or U8550 (N_8550,N_8296,N_8324);
nand U8551 (N_8551,N_8292,N_8481);
nand U8552 (N_8552,N_8364,N_8488);
nand U8553 (N_8553,N_8354,N_8352);
nand U8554 (N_8554,N_8491,N_8429);
nor U8555 (N_8555,N_8486,N_8400);
or U8556 (N_8556,N_8460,N_8299);
nor U8557 (N_8557,N_8483,N_8332);
xor U8558 (N_8558,N_8476,N_8300);
xnor U8559 (N_8559,N_8489,N_8351);
nor U8560 (N_8560,N_8421,N_8304);
and U8561 (N_8561,N_8306,N_8275);
xor U8562 (N_8562,N_8434,N_8427);
nand U8563 (N_8563,N_8310,N_8447);
and U8564 (N_8564,N_8376,N_8499);
nand U8565 (N_8565,N_8307,N_8393);
xnor U8566 (N_8566,N_8441,N_8252);
or U8567 (N_8567,N_8250,N_8394);
and U8568 (N_8568,N_8474,N_8254);
xnor U8569 (N_8569,N_8258,N_8444);
nand U8570 (N_8570,N_8287,N_8323);
nand U8571 (N_8571,N_8457,N_8267);
or U8572 (N_8572,N_8443,N_8327);
xnor U8573 (N_8573,N_8436,N_8414);
or U8574 (N_8574,N_8490,N_8263);
or U8575 (N_8575,N_8454,N_8335);
or U8576 (N_8576,N_8426,N_8330);
xor U8577 (N_8577,N_8495,N_8417);
nor U8578 (N_8578,N_8343,N_8397);
xor U8579 (N_8579,N_8346,N_8401);
xor U8580 (N_8580,N_8339,N_8341);
nand U8581 (N_8581,N_8308,N_8407);
xnor U8582 (N_8582,N_8265,N_8270);
nand U8583 (N_8583,N_8448,N_8353);
nor U8584 (N_8584,N_8435,N_8468);
or U8585 (N_8585,N_8440,N_8422);
nand U8586 (N_8586,N_8259,N_8480);
or U8587 (N_8587,N_8465,N_8251);
and U8588 (N_8588,N_8412,N_8384);
or U8589 (N_8589,N_8260,N_8381);
nor U8590 (N_8590,N_8379,N_8301);
nor U8591 (N_8591,N_8337,N_8366);
and U8592 (N_8592,N_8388,N_8315);
xor U8593 (N_8593,N_8361,N_8278);
or U8594 (N_8594,N_8461,N_8340);
or U8595 (N_8595,N_8367,N_8309);
xnor U8596 (N_8596,N_8485,N_8314);
nand U8597 (N_8597,N_8449,N_8318);
xnor U8598 (N_8598,N_8276,N_8355);
nand U8599 (N_8599,N_8369,N_8418);
nor U8600 (N_8600,N_8455,N_8433);
and U8601 (N_8601,N_8392,N_8273);
xnor U8602 (N_8602,N_8350,N_8322);
nand U8603 (N_8603,N_8402,N_8450);
xor U8604 (N_8604,N_8291,N_8452);
or U8605 (N_8605,N_8283,N_8442);
and U8606 (N_8606,N_8472,N_8389);
and U8607 (N_8607,N_8419,N_8420);
xnor U8608 (N_8608,N_8316,N_8469);
or U8609 (N_8609,N_8446,N_8431);
and U8610 (N_8610,N_8290,N_8382);
nor U8611 (N_8611,N_8298,N_8268);
xnor U8612 (N_8612,N_8390,N_8331);
nand U8613 (N_8613,N_8416,N_8305);
nand U8614 (N_8614,N_8334,N_8479);
nand U8615 (N_8615,N_8458,N_8430);
and U8616 (N_8616,N_8295,N_8284);
xor U8617 (N_8617,N_8403,N_8478);
or U8618 (N_8618,N_8274,N_8264);
nor U8619 (N_8619,N_8344,N_8405);
nor U8620 (N_8620,N_8493,N_8356);
nand U8621 (N_8621,N_8261,N_8288);
nor U8622 (N_8622,N_8415,N_8410);
nor U8623 (N_8623,N_8362,N_8266);
xor U8624 (N_8624,N_8473,N_8395);
and U8625 (N_8625,N_8497,N_8287);
and U8626 (N_8626,N_8352,N_8444);
nand U8627 (N_8627,N_8328,N_8486);
or U8628 (N_8628,N_8266,N_8343);
xor U8629 (N_8629,N_8453,N_8385);
or U8630 (N_8630,N_8461,N_8429);
nor U8631 (N_8631,N_8297,N_8334);
and U8632 (N_8632,N_8345,N_8383);
and U8633 (N_8633,N_8448,N_8465);
or U8634 (N_8634,N_8349,N_8327);
nand U8635 (N_8635,N_8345,N_8394);
nand U8636 (N_8636,N_8344,N_8431);
nor U8637 (N_8637,N_8434,N_8498);
or U8638 (N_8638,N_8285,N_8411);
and U8639 (N_8639,N_8359,N_8422);
xnor U8640 (N_8640,N_8254,N_8345);
or U8641 (N_8641,N_8330,N_8498);
nor U8642 (N_8642,N_8287,N_8458);
nand U8643 (N_8643,N_8380,N_8394);
nor U8644 (N_8644,N_8494,N_8479);
xnor U8645 (N_8645,N_8302,N_8487);
nand U8646 (N_8646,N_8419,N_8388);
or U8647 (N_8647,N_8433,N_8363);
xor U8648 (N_8648,N_8453,N_8306);
nand U8649 (N_8649,N_8396,N_8475);
and U8650 (N_8650,N_8421,N_8491);
or U8651 (N_8651,N_8378,N_8314);
and U8652 (N_8652,N_8364,N_8349);
nand U8653 (N_8653,N_8264,N_8424);
xor U8654 (N_8654,N_8283,N_8308);
xor U8655 (N_8655,N_8492,N_8477);
or U8656 (N_8656,N_8280,N_8456);
xor U8657 (N_8657,N_8266,N_8387);
or U8658 (N_8658,N_8433,N_8286);
nand U8659 (N_8659,N_8432,N_8393);
nor U8660 (N_8660,N_8386,N_8337);
and U8661 (N_8661,N_8488,N_8348);
or U8662 (N_8662,N_8257,N_8340);
xor U8663 (N_8663,N_8456,N_8462);
nor U8664 (N_8664,N_8439,N_8350);
or U8665 (N_8665,N_8252,N_8335);
or U8666 (N_8666,N_8302,N_8275);
nor U8667 (N_8667,N_8495,N_8401);
or U8668 (N_8668,N_8369,N_8353);
nor U8669 (N_8669,N_8433,N_8292);
xnor U8670 (N_8670,N_8330,N_8406);
and U8671 (N_8671,N_8361,N_8297);
xor U8672 (N_8672,N_8355,N_8258);
or U8673 (N_8673,N_8298,N_8460);
xor U8674 (N_8674,N_8408,N_8420);
xnor U8675 (N_8675,N_8300,N_8274);
xor U8676 (N_8676,N_8323,N_8277);
or U8677 (N_8677,N_8252,N_8430);
xor U8678 (N_8678,N_8374,N_8292);
xnor U8679 (N_8679,N_8365,N_8257);
xnor U8680 (N_8680,N_8254,N_8250);
nor U8681 (N_8681,N_8304,N_8434);
or U8682 (N_8682,N_8410,N_8358);
nor U8683 (N_8683,N_8360,N_8494);
or U8684 (N_8684,N_8301,N_8298);
nor U8685 (N_8685,N_8386,N_8481);
xnor U8686 (N_8686,N_8473,N_8486);
nor U8687 (N_8687,N_8390,N_8453);
nor U8688 (N_8688,N_8430,N_8385);
and U8689 (N_8689,N_8329,N_8498);
xor U8690 (N_8690,N_8473,N_8276);
or U8691 (N_8691,N_8479,N_8332);
nand U8692 (N_8692,N_8350,N_8485);
nand U8693 (N_8693,N_8270,N_8395);
nor U8694 (N_8694,N_8303,N_8386);
or U8695 (N_8695,N_8483,N_8328);
and U8696 (N_8696,N_8372,N_8331);
nand U8697 (N_8697,N_8333,N_8416);
and U8698 (N_8698,N_8480,N_8309);
nor U8699 (N_8699,N_8257,N_8286);
nor U8700 (N_8700,N_8282,N_8255);
or U8701 (N_8701,N_8338,N_8287);
and U8702 (N_8702,N_8495,N_8268);
xnor U8703 (N_8703,N_8399,N_8371);
nand U8704 (N_8704,N_8278,N_8271);
or U8705 (N_8705,N_8322,N_8421);
xor U8706 (N_8706,N_8415,N_8349);
nand U8707 (N_8707,N_8492,N_8259);
nand U8708 (N_8708,N_8404,N_8433);
xnor U8709 (N_8709,N_8306,N_8350);
or U8710 (N_8710,N_8447,N_8415);
and U8711 (N_8711,N_8422,N_8279);
nand U8712 (N_8712,N_8369,N_8318);
and U8713 (N_8713,N_8338,N_8307);
nand U8714 (N_8714,N_8250,N_8298);
nor U8715 (N_8715,N_8342,N_8320);
nand U8716 (N_8716,N_8452,N_8402);
nor U8717 (N_8717,N_8478,N_8287);
and U8718 (N_8718,N_8432,N_8254);
nand U8719 (N_8719,N_8430,N_8256);
nand U8720 (N_8720,N_8413,N_8390);
xor U8721 (N_8721,N_8261,N_8428);
nor U8722 (N_8722,N_8367,N_8426);
nor U8723 (N_8723,N_8352,N_8450);
or U8724 (N_8724,N_8298,N_8340);
nor U8725 (N_8725,N_8273,N_8420);
and U8726 (N_8726,N_8250,N_8459);
nor U8727 (N_8727,N_8396,N_8300);
nand U8728 (N_8728,N_8476,N_8387);
or U8729 (N_8729,N_8280,N_8407);
and U8730 (N_8730,N_8495,N_8322);
nand U8731 (N_8731,N_8414,N_8325);
nand U8732 (N_8732,N_8412,N_8432);
nor U8733 (N_8733,N_8487,N_8260);
or U8734 (N_8734,N_8329,N_8344);
nand U8735 (N_8735,N_8321,N_8426);
xnor U8736 (N_8736,N_8276,N_8378);
xnor U8737 (N_8737,N_8424,N_8489);
nand U8738 (N_8738,N_8351,N_8449);
nor U8739 (N_8739,N_8275,N_8270);
xor U8740 (N_8740,N_8287,N_8452);
or U8741 (N_8741,N_8482,N_8480);
nand U8742 (N_8742,N_8315,N_8441);
xor U8743 (N_8743,N_8273,N_8259);
or U8744 (N_8744,N_8277,N_8395);
and U8745 (N_8745,N_8329,N_8450);
nand U8746 (N_8746,N_8392,N_8402);
nand U8747 (N_8747,N_8324,N_8254);
and U8748 (N_8748,N_8461,N_8498);
nand U8749 (N_8749,N_8422,N_8477);
and U8750 (N_8750,N_8623,N_8555);
or U8751 (N_8751,N_8545,N_8645);
xor U8752 (N_8752,N_8706,N_8606);
or U8753 (N_8753,N_8710,N_8632);
and U8754 (N_8754,N_8601,N_8746);
and U8755 (N_8755,N_8633,N_8748);
nor U8756 (N_8756,N_8622,N_8513);
nand U8757 (N_8757,N_8727,N_8556);
nand U8758 (N_8758,N_8559,N_8547);
and U8759 (N_8759,N_8616,N_8560);
nor U8760 (N_8760,N_8707,N_8569);
nor U8761 (N_8761,N_8735,N_8517);
and U8762 (N_8762,N_8600,N_8716);
or U8763 (N_8763,N_8612,N_8535);
or U8764 (N_8764,N_8652,N_8644);
and U8765 (N_8765,N_8672,N_8566);
and U8766 (N_8766,N_8639,N_8507);
and U8767 (N_8767,N_8641,N_8646);
or U8768 (N_8768,N_8531,N_8609);
or U8769 (N_8769,N_8694,N_8574);
xor U8770 (N_8770,N_8651,N_8564);
and U8771 (N_8771,N_8551,N_8658);
xor U8772 (N_8772,N_8691,N_8553);
xnor U8773 (N_8773,N_8557,N_8515);
nand U8774 (N_8774,N_8740,N_8525);
or U8775 (N_8775,N_8687,N_8656);
xor U8776 (N_8776,N_8544,N_8508);
and U8777 (N_8777,N_8734,N_8621);
and U8778 (N_8778,N_8540,N_8543);
xor U8779 (N_8779,N_8567,N_8587);
nor U8780 (N_8780,N_8561,N_8520);
nor U8781 (N_8781,N_8703,N_8638);
or U8782 (N_8782,N_8733,N_8728);
xor U8783 (N_8783,N_8677,N_8550);
nand U8784 (N_8784,N_8693,N_8722);
xnor U8785 (N_8785,N_8620,N_8577);
xor U8786 (N_8786,N_8685,N_8744);
xnor U8787 (N_8787,N_8699,N_8604);
xnor U8788 (N_8788,N_8676,N_8701);
xnor U8789 (N_8789,N_8618,N_8709);
nor U8790 (N_8790,N_8665,N_8666);
or U8791 (N_8791,N_8558,N_8675);
or U8792 (N_8792,N_8714,N_8503);
and U8793 (N_8793,N_8669,N_8527);
nand U8794 (N_8794,N_8501,N_8681);
or U8795 (N_8795,N_8537,N_8625);
nor U8796 (N_8796,N_8530,N_8529);
nand U8797 (N_8797,N_8749,N_8590);
nand U8798 (N_8798,N_8667,N_8648);
or U8799 (N_8799,N_8584,N_8607);
or U8800 (N_8800,N_8702,N_8598);
nand U8801 (N_8801,N_8522,N_8689);
nand U8802 (N_8802,N_8659,N_8662);
or U8803 (N_8803,N_8649,N_8673);
nor U8804 (N_8804,N_8581,N_8713);
xor U8805 (N_8805,N_8512,N_8663);
or U8806 (N_8806,N_8614,N_8653);
nand U8807 (N_8807,N_8700,N_8745);
xor U8808 (N_8808,N_8660,N_8736);
or U8809 (N_8809,N_8636,N_8511);
nor U8810 (N_8810,N_8549,N_8536);
nand U8811 (N_8811,N_8631,N_8548);
xnor U8812 (N_8812,N_8500,N_8690);
nor U8813 (N_8813,N_8519,N_8715);
nand U8814 (N_8814,N_8592,N_8747);
or U8815 (N_8815,N_8708,N_8720);
xor U8816 (N_8816,N_8610,N_8628);
or U8817 (N_8817,N_8533,N_8657);
xnor U8818 (N_8818,N_8647,N_8719);
xor U8819 (N_8819,N_8554,N_8724);
nand U8820 (N_8820,N_8552,N_8627);
nor U8821 (N_8821,N_8718,N_8576);
xnor U8822 (N_8822,N_8717,N_8615);
nand U8823 (N_8823,N_8741,N_8640);
or U8824 (N_8824,N_8596,N_8509);
and U8825 (N_8825,N_8626,N_8534);
xnor U8826 (N_8826,N_8729,N_8504);
xor U8827 (N_8827,N_8588,N_8580);
or U8828 (N_8828,N_8603,N_8505);
nand U8829 (N_8829,N_8679,N_8650);
xor U8830 (N_8830,N_8664,N_8506);
or U8831 (N_8831,N_8518,N_8562);
and U8832 (N_8832,N_8629,N_8682);
and U8833 (N_8833,N_8661,N_8686);
and U8834 (N_8834,N_8680,N_8613);
nand U8835 (N_8835,N_8605,N_8670);
xnor U8836 (N_8836,N_8565,N_8726);
or U8837 (N_8837,N_8583,N_8698);
and U8838 (N_8838,N_8688,N_8668);
nand U8839 (N_8839,N_8510,N_8643);
nand U8840 (N_8840,N_8573,N_8723);
nor U8841 (N_8841,N_8619,N_8739);
nor U8842 (N_8842,N_8538,N_8542);
and U8843 (N_8843,N_8696,N_8575);
and U8844 (N_8844,N_8711,N_8526);
or U8845 (N_8845,N_8705,N_8630);
and U8846 (N_8846,N_8524,N_8602);
nand U8847 (N_8847,N_8743,N_8563);
nand U8848 (N_8848,N_8582,N_8683);
nor U8849 (N_8849,N_8608,N_8528);
nand U8850 (N_8850,N_8697,N_8617);
and U8851 (N_8851,N_8571,N_8655);
nand U8852 (N_8852,N_8731,N_8585);
and U8853 (N_8853,N_8704,N_8572);
or U8854 (N_8854,N_8586,N_8635);
and U8855 (N_8855,N_8502,N_8732);
or U8856 (N_8856,N_8611,N_8599);
nand U8857 (N_8857,N_8712,N_8725);
nand U8858 (N_8858,N_8695,N_8597);
or U8859 (N_8859,N_8521,N_8595);
nor U8860 (N_8860,N_8546,N_8654);
nand U8861 (N_8861,N_8568,N_8541);
nor U8862 (N_8862,N_8579,N_8578);
nand U8863 (N_8863,N_8684,N_8637);
xnor U8864 (N_8864,N_8523,N_8570);
nor U8865 (N_8865,N_8532,N_8642);
xnor U8866 (N_8866,N_8594,N_8514);
nand U8867 (N_8867,N_8671,N_8593);
nand U8868 (N_8868,N_8721,N_8737);
nor U8869 (N_8869,N_8634,N_8539);
nor U8870 (N_8870,N_8591,N_8624);
nand U8871 (N_8871,N_8692,N_8674);
xor U8872 (N_8872,N_8678,N_8516);
nor U8873 (N_8873,N_8730,N_8589);
or U8874 (N_8874,N_8742,N_8738);
nand U8875 (N_8875,N_8694,N_8675);
nor U8876 (N_8876,N_8661,N_8722);
and U8877 (N_8877,N_8687,N_8691);
and U8878 (N_8878,N_8737,N_8688);
nand U8879 (N_8879,N_8749,N_8673);
and U8880 (N_8880,N_8633,N_8597);
or U8881 (N_8881,N_8582,N_8539);
or U8882 (N_8882,N_8694,N_8578);
xor U8883 (N_8883,N_8670,N_8612);
nand U8884 (N_8884,N_8612,N_8724);
xor U8885 (N_8885,N_8538,N_8651);
nor U8886 (N_8886,N_8606,N_8687);
or U8887 (N_8887,N_8525,N_8674);
and U8888 (N_8888,N_8631,N_8697);
nor U8889 (N_8889,N_8526,N_8665);
and U8890 (N_8890,N_8655,N_8600);
xnor U8891 (N_8891,N_8674,N_8658);
nand U8892 (N_8892,N_8712,N_8722);
xor U8893 (N_8893,N_8733,N_8720);
xnor U8894 (N_8894,N_8503,N_8647);
and U8895 (N_8895,N_8716,N_8695);
and U8896 (N_8896,N_8619,N_8648);
nor U8897 (N_8897,N_8667,N_8558);
xor U8898 (N_8898,N_8644,N_8699);
nor U8899 (N_8899,N_8645,N_8623);
or U8900 (N_8900,N_8729,N_8624);
nor U8901 (N_8901,N_8720,N_8651);
nor U8902 (N_8902,N_8685,N_8619);
nand U8903 (N_8903,N_8746,N_8618);
and U8904 (N_8904,N_8558,N_8549);
nor U8905 (N_8905,N_8503,N_8610);
and U8906 (N_8906,N_8614,N_8746);
xor U8907 (N_8907,N_8740,N_8710);
nand U8908 (N_8908,N_8522,N_8510);
xor U8909 (N_8909,N_8652,N_8612);
xor U8910 (N_8910,N_8507,N_8546);
and U8911 (N_8911,N_8532,N_8637);
nand U8912 (N_8912,N_8542,N_8724);
nor U8913 (N_8913,N_8606,N_8554);
xnor U8914 (N_8914,N_8647,N_8603);
nor U8915 (N_8915,N_8576,N_8583);
xnor U8916 (N_8916,N_8572,N_8500);
and U8917 (N_8917,N_8678,N_8612);
nand U8918 (N_8918,N_8524,N_8743);
and U8919 (N_8919,N_8746,N_8668);
or U8920 (N_8920,N_8617,N_8554);
xnor U8921 (N_8921,N_8719,N_8708);
nor U8922 (N_8922,N_8612,N_8738);
nor U8923 (N_8923,N_8740,N_8504);
xnor U8924 (N_8924,N_8669,N_8509);
nor U8925 (N_8925,N_8538,N_8582);
nand U8926 (N_8926,N_8740,N_8623);
nand U8927 (N_8927,N_8556,N_8706);
or U8928 (N_8928,N_8651,N_8565);
nor U8929 (N_8929,N_8531,N_8625);
xnor U8930 (N_8930,N_8615,N_8672);
and U8931 (N_8931,N_8584,N_8658);
or U8932 (N_8932,N_8659,N_8736);
nor U8933 (N_8933,N_8626,N_8688);
nor U8934 (N_8934,N_8707,N_8566);
and U8935 (N_8935,N_8614,N_8726);
or U8936 (N_8936,N_8548,N_8553);
and U8937 (N_8937,N_8635,N_8674);
nor U8938 (N_8938,N_8605,N_8596);
or U8939 (N_8939,N_8557,N_8520);
xor U8940 (N_8940,N_8706,N_8680);
nand U8941 (N_8941,N_8582,N_8552);
or U8942 (N_8942,N_8673,N_8657);
xnor U8943 (N_8943,N_8690,N_8633);
xnor U8944 (N_8944,N_8628,N_8728);
or U8945 (N_8945,N_8692,N_8673);
nand U8946 (N_8946,N_8661,N_8625);
or U8947 (N_8947,N_8735,N_8615);
nor U8948 (N_8948,N_8612,N_8579);
or U8949 (N_8949,N_8747,N_8705);
or U8950 (N_8950,N_8684,N_8643);
nor U8951 (N_8951,N_8559,N_8589);
or U8952 (N_8952,N_8740,N_8575);
and U8953 (N_8953,N_8597,N_8637);
or U8954 (N_8954,N_8597,N_8500);
or U8955 (N_8955,N_8601,N_8588);
or U8956 (N_8956,N_8531,N_8630);
xnor U8957 (N_8957,N_8638,N_8739);
xor U8958 (N_8958,N_8635,N_8676);
nor U8959 (N_8959,N_8637,N_8638);
or U8960 (N_8960,N_8632,N_8566);
nand U8961 (N_8961,N_8607,N_8616);
nand U8962 (N_8962,N_8639,N_8627);
nand U8963 (N_8963,N_8579,N_8521);
or U8964 (N_8964,N_8656,N_8623);
or U8965 (N_8965,N_8606,N_8708);
or U8966 (N_8966,N_8713,N_8605);
and U8967 (N_8967,N_8711,N_8692);
nand U8968 (N_8968,N_8577,N_8665);
and U8969 (N_8969,N_8562,N_8513);
nor U8970 (N_8970,N_8537,N_8573);
xor U8971 (N_8971,N_8574,N_8663);
or U8972 (N_8972,N_8743,N_8693);
nor U8973 (N_8973,N_8653,N_8644);
xor U8974 (N_8974,N_8509,N_8555);
and U8975 (N_8975,N_8551,N_8659);
or U8976 (N_8976,N_8634,N_8534);
nand U8977 (N_8977,N_8607,N_8707);
nand U8978 (N_8978,N_8556,N_8692);
and U8979 (N_8979,N_8609,N_8707);
nor U8980 (N_8980,N_8690,N_8558);
nor U8981 (N_8981,N_8578,N_8587);
xnor U8982 (N_8982,N_8644,N_8505);
nand U8983 (N_8983,N_8561,N_8704);
or U8984 (N_8984,N_8672,N_8520);
or U8985 (N_8985,N_8745,N_8727);
and U8986 (N_8986,N_8605,N_8686);
and U8987 (N_8987,N_8718,N_8719);
and U8988 (N_8988,N_8712,N_8657);
nand U8989 (N_8989,N_8718,N_8667);
nand U8990 (N_8990,N_8596,N_8602);
nand U8991 (N_8991,N_8505,N_8723);
nand U8992 (N_8992,N_8646,N_8725);
or U8993 (N_8993,N_8658,N_8502);
and U8994 (N_8994,N_8719,N_8649);
xnor U8995 (N_8995,N_8550,N_8586);
and U8996 (N_8996,N_8595,N_8585);
xnor U8997 (N_8997,N_8575,N_8703);
nand U8998 (N_8998,N_8668,N_8528);
or U8999 (N_8999,N_8695,N_8589);
or U9000 (N_9000,N_8902,N_8926);
and U9001 (N_9001,N_8766,N_8942);
xnor U9002 (N_9002,N_8952,N_8818);
or U9003 (N_9003,N_8806,N_8887);
nand U9004 (N_9004,N_8807,N_8870);
nor U9005 (N_9005,N_8830,N_8827);
nand U9006 (N_9006,N_8900,N_8854);
xnor U9007 (N_9007,N_8963,N_8773);
or U9008 (N_9008,N_8915,N_8856);
nor U9009 (N_9009,N_8792,N_8759);
or U9010 (N_9010,N_8767,N_8780);
or U9011 (N_9011,N_8757,N_8891);
xor U9012 (N_9012,N_8785,N_8927);
nand U9013 (N_9013,N_8871,N_8947);
and U9014 (N_9014,N_8760,N_8881);
xor U9015 (N_9015,N_8844,N_8933);
and U9016 (N_9016,N_8974,N_8916);
and U9017 (N_9017,N_8843,N_8869);
or U9018 (N_9018,N_8992,N_8850);
xor U9019 (N_9019,N_8803,N_8975);
xor U9020 (N_9020,N_8978,N_8839);
nand U9021 (N_9021,N_8977,N_8875);
nor U9022 (N_9022,N_8953,N_8834);
xnor U9023 (N_9023,N_8795,N_8802);
nand U9024 (N_9024,N_8804,N_8849);
xor U9025 (N_9025,N_8790,N_8815);
xor U9026 (N_9026,N_8980,N_8903);
or U9027 (N_9027,N_8973,N_8880);
xnor U9028 (N_9028,N_8946,N_8838);
nor U9029 (N_9029,N_8884,N_8750);
nor U9030 (N_9030,N_8886,N_8833);
or U9031 (N_9031,N_8805,N_8841);
and U9032 (N_9032,N_8829,N_8883);
nand U9033 (N_9033,N_8812,N_8832);
nand U9034 (N_9034,N_8852,N_8799);
nor U9035 (N_9035,N_8752,N_8996);
and U9036 (N_9036,N_8896,N_8999);
nand U9037 (N_9037,N_8961,N_8855);
xnor U9038 (N_9038,N_8986,N_8965);
or U9039 (N_9039,N_8761,N_8816);
nor U9040 (N_9040,N_8800,N_8779);
nor U9041 (N_9041,N_8835,N_8956);
nor U9042 (N_9042,N_8894,N_8840);
or U9043 (N_9043,N_8948,N_8879);
or U9044 (N_9044,N_8905,N_8967);
xor U9045 (N_9045,N_8866,N_8922);
and U9046 (N_9046,N_8808,N_8983);
xor U9047 (N_9047,N_8958,N_8971);
or U9048 (N_9048,N_8831,N_8837);
and U9049 (N_9049,N_8984,N_8814);
nand U9050 (N_9050,N_8899,N_8794);
xnor U9051 (N_9051,N_8964,N_8796);
xnor U9052 (N_9052,N_8774,N_8867);
or U9053 (N_9053,N_8888,N_8991);
nand U9054 (N_9054,N_8758,N_8817);
and U9055 (N_9055,N_8826,N_8824);
and U9056 (N_9056,N_8931,N_8770);
and U9057 (N_9057,N_8929,N_8819);
and U9058 (N_9058,N_8797,N_8951);
xor U9059 (N_9059,N_8823,N_8810);
xor U9060 (N_9060,N_8784,N_8865);
and U9061 (N_9061,N_8943,N_8876);
nand U9062 (N_9062,N_8783,N_8775);
or U9063 (N_9063,N_8782,N_8919);
nand U9064 (N_9064,N_8845,N_8861);
nand U9065 (N_9065,N_8987,N_8889);
nor U9066 (N_9066,N_8908,N_8938);
and U9067 (N_9067,N_8921,N_8769);
or U9068 (N_9068,N_8914,N_8968);
and U9069 (N_9069,N_8918,N_8836);
nor U9070 (N_9070,N_8930,N_8842);
nor U9071 (N_9071,N_8828,N_8937);
nand U9072 (N_9072,N_8753,N_8853);
nor U9073 (N_9073,N_8771,N_8972);
nand U9074 (N_9074,N_8940,N_8923);
xnor U9075 (N_9075,N_8872,N_8962);
nor U9076 (N_9076,N_8847,N_8990);
nor U9077 (N_9077,N_8960,N_8939);
or U9078 (N_9078,N_8778,N_8901);
or U9079 (N_9079,N_8787,N_8859);
or U9080 (N_9080,N_8910,N_8995);
or U9081 (N_9081,N_8955,N_8981);
nor U9082 (N_9082,N_8925,N_8890);
and U9083 (N_9083,N_8954,N_8820);
xor U9084 (N_9084,N_8957,N_8885);
nand U9085 (N_9085,N_8873,N_8928);
or U9086 (N_9086,N_8920,N_8906);
and U9087 (N_9087,N_8979,N_8959);
nor U9088 (N_9088,N_8825,N_8976);
nor U9089 (N_9089,N_8950,N_8811);
xnor U9090 (N_9090,N_8858,N_8907);
or U9091 (N_9091,N_8864,N_8913);
nand U9092 (N_9092,N_8988,N_8949);
or U9093 (N_9093,N_8801,N_8966);
nand U9094 (N_9094,N_8944,N_8993);
xor U9095 (N_9095,N_8932,N_8763);
nor U9096 (N_9096,N_8776,N_8821);
nand U9097 (N_9097,N_8848,N_8851);
nand U9098 (N_9098,N_8789,N_8989);
or U9099 (N_9099,N_8809,N_8893);
nand U9100 (N_9100,N_8764,N_8762);
xnor U9101 (N_9101,N_8904,N_8924);
nor U9102 (N_9102,N_8998,N_8982);
nand U9103 (N_9103,N_8897,N_8765);
nand U9104 (N_9104,N_8970,N_8863);
nor U9105 (N_9105,N_8781,N_8935);
xnor U9106 (N_9106,N_8868,N_8917);
nor U9107 (N_9107,N_8911,N_8882);
and U9108 (N_9108,N_8934,N_8877);
nand U9109 (N_9109,N_8754,N_8822);
nor U9110 (N_9110,N_8912,N_8941);
xnor U9111 (N_9111,N_8846,N_8793);
or U9112 (N_9112,N_8878,N_8788);
nor U9113 (N_9113,N_8985,N_8751);
nor U9114 (N_9114,N_8874,N_8756);
nand U9115 (N_9115,N_8777,N_8945);
nand U9116 (N_9116,N_8791,N_8857);
nand U9117 (N_9117,N_8772,N_8994);
or U9118 (N_9118,N_8860,N_8755);
nor U9119 (N_9119,N_8909,N_8768);
xnor U9120 (N_9120,N_8895,N_8892);
xor U9121 (N_9121,N_8997,N_8969);
nor U9122 (N_9122,N_8936,N_8813);
xnor U9123 (N_9123,N_8786,N_8798);
nand U9124 (N_9124,N_8898,N_8862);
xor U9125 (N_9125,N_8819,N_8956);
and U9126 (N_9126,N_8912,N_8787);
nor U9127 (N_9127,N_8778,N_8804);
or U9128 (N_9128,N_8993,N_8968);
and U9129 (N_9129,N_8818,N_8910);
nand U9130 (N_9130,N_8949,N_8971);
xor U9131 (N_9131,N_8920,N_8867);
nand U9132 (N_9132,N_8891,N_8879);
nand U9133 (N_9133,N_8918,N_8961);
nand U9134 (N_9134,N_8963,N_8800);
and U9135 (N_9135,N_8793,N_8925);
nor U9136 (N_9136,N_8788,N_8985);
and U9137 (N_9137,N_8903,N_8970);
xor U9138 (N_9138,N_8851,N_8818);
nor U9139 (N_9139,N_8770,N_8867);
nand U9140 (N_9140,N_8812,N_8889);
nand U9141 (N_9141,N_8872,N_8964);
nand U9142 (N_9142,N_8847,N_8757);
or U9143 (N_9143,N_8771,N_8897);
and U9144 (N_9144,N_8771,N_8882);
or U9145 (N_9145,N_8793,N_8921);
xor U9146 (N_9146,N_8953,N_8944);
and U9147 (N_9147,N_8903,N_8993);
xor U9148 (N_9148,N_8951,N_8914);
and U9149 (N_9149,N_8793,N_8895);
xor U9150 (N_9150,N_8819,N_8855);
nand U9151 (N_9151,N_8964,N_8816);
xor U9152 (N_9152,N_8782,N_8762);
or U9153 (N_9153,N_8821,N_8799);
or U9154 (N_9154,N_8816,N_8820);
or U9155 (N_9155,N_8870,N_8788);
and U9156 (N_9156,N_8946,N_8777);
nand U9157 (N_9157,N_8772,N_8919);
nand U9158 (N_9158,N_8764,N_8943);
nand U9159 (N_9159,N_8779,N_8926);
or U9160 (N_9160,N_8926,N_8764);
nand U9161 (N_9161,N_8785,N_8900);
or U9162 (N_9162,N_8892,N_8853);
nand U9163 (N_9163,N_8812,N_8928);
nand U9164 (N_9164,N_8850,N_8918);
or U9165 (N_9165,N_8800,N_8851);
xor U9166 (N_9166,N_8821,N_8793);
xnor U9167 (N_9167,N_8908,N_8755);
nand U9168 (N_9168,N_8835,N_8826);
nand U9169 (N_9169,N_8781,N_8762);
or U9170 (N_9170,N_8798,N_8933);
nor U9171 (N_9171,N_8942,N_8974);
and U9172 (N_9172,N_8764,N_8990);
nor U9173 (N_9173,N_8866,N_8970);
nand U9174 (N_9174,N_8889,N_8794);
nor U9175 (N_9175,N_8941,N_8993);
xnor U9176 (N_9176,N_8974,N_8767);
or U9177 (N_9177,N_8821,N_8964);
nand U9178 (N_9178,N_8916,N_8889);
xnor U9179 (N_9179,N_8913,N_8954);
xnor U9180 (N_9180,N_8821,N_8862);
and U9181 (N_9181,N_8815,N_8831);
or U9182 (N_9182,N_8905,N_8861);
or U9183 (N_9183,N_8991,N_8955);
xor U9184 (N_9184,N_8919,N_8945);
or U9185 (N_9185,N_8930,N_8925);
xor U9186 (N_9186,N_8793,N_8773);
xor U9187 (N_9187,N_8783,N_8862);
xnor U9188 (N_9188,N_8959,N_8931);
nand U9189 (N_9189,N_8917,N_8855);
nand U9190 (N_9190,N_8897,N_8940);
xnor U9191 (N_9191,N_8755,N_8854);
nand U9192 (N_9192,N_8785,N_8805);
xor U9193 (N_9193,N_8959,N_8858);
nand U9194 (N_9194,N_8945,N_8974);
or U9195 (N_9195,N_8859,N_8981);
nor U9196 (N_9196,N_8918,N_8765);
and U9197 (N_9197,N_8789,N_8952);
nor U9198 (N_9198,N_8928,N_8891);
xnor U9199 (N_9199,N_8915,N_8783);
nor U9200 (N_9200,N_8786,N_8869);
nor U9201 (N_9201,N_8939,N_8918);
nand U9202 (N_9202,N_8825,N_8967);
and U9203 (N_9203,N_8879,N_8881);
nor U9204 (N_9204,N_8788,N_8955);
nand U9205 (N_9205,N_8825,N_8923);
xor U9206 (N_9206,N_8991,N_8788);
xor U9207 (N_9207,N_8992,N_8907);
and U9208 (N_9208,N_8969,N_8868);
or U9209 (N_9209,N_8775,N_8903);
nor U9210 (N_9210,N_8958,N_8999);
nor U9211 (N_9211,N_8836,N_8945);
nor U9212 (N_9212,N_8913,N_8852);
xor U9213 (N_9213,N_8911,N_8762);
and U9214 (N_9214,N_8814,N_8972);
and U9215 (N_9215,N_8859,N_8941);
xnor U9216 (N_9216,N_8762,N_8786);
and U9217 (N_9217,N_8983,N_8831);
xnor U9218 (N_9218,N_8893,N_8899);
nand U9219 (N_9219,N_8987,N_8890);
or U9220 (N_9220,N_8842,N_8803);
and U9221 (N_9221,N_8919,N_8849);
nor U9222 (N_9222,N_8968,N_8970);
and U9223 (N_9223,N_8833,N_8962);
nor U9224 (N_9224,N_8930,N_8979);
xnor U9225 (N_9225,N_8878,N_8848);
and U9226 (N_9226,N_8845,N_8943);
xnor U9227 (N_9227,N_8929,N_8974);
nor U9228 (N_9228,N_8795,N_8970);
and U9229 (N_9229,N_8990,N_8961);
and U9230 (N_9230,N_8822,N_8835);
nor U9231 (N_9231,N_8871,N_8780);
or U9232 (N_9232,N_8812,N_8929);
and U9233 (N_9233,N_8981,N_8809);
and U9234 (N_9234,N_8973,N_8882);
xor U9235 (N_9235,N_8991,N_8927);
or U9236 (N_9236,N_8796,N_8920);
nor U9237 (N_9237,N_8984,N_8777);
or U9238 (N_9238,N_8795,N_8879);
nand U9239 (N_9239,N_8913,N_8956);
nor U9240 (N_9240,N_8788,N_8905);
or U9241 (N_9241,N_8769,N_8898);
nor U9242 (N_9242,N_8838,N_8985);
nand U9243 (N_9243,N_8792,N_8844);
and U9244 (N_9244,N_8868,N_8973);
xnor U9245 (N_9245,N_8972,N_8839);
or U9246 (N_9246,N_8806,N_8904);
nor U9247 (N_9247,N_8968,N_8861);
nand U9248 (N_9248,N_8813,N_8784);
nor U9249 (N_9249,N_8802,N_8787);
nand U9250 (N_9250,N_9066,N_9138);
or U9251 (N_9251,N_9087,N_9054);
or U9252 (N_9252,N_9188,N_9210);
nand U9253 (N_9253,N_9043,N_9103);
xor U9254 (N_9254,N_9102,N_9203);
nor U9255 (N_9255,N_9244,N_9115);
nand U9256 (N_9256,N_9129,N_9093);
or U9257 (N_9257,N_9196,N_9169);
xnor U9258 (N_9258,N_9029,N_9187);
nand U9259 (N_9259,N_9100,N_9040);
and U9260 (N_9260,N_9032,N_9194);
nor U9261 (N_9261,N_9070,N_9174);
and U9262 (N_9262,N_9038,N_9033);
or U9263 (N_9263,N_9160,N_9171);
nor U9264 (N_9264,N_9105,N_9081);
or U9265 (N_9265,N_9155,N_9168);
nor U9266 (N_9266,N_9104,N_9112);
xor U9267 (N_9267,N_9120,N_9075);
nand U9268 (N_9268,N_9123,N_9204);
or U9269 (N_9269,N_9201,N_9215);
nor U9270 (N_9270,N_9128,N_9202);
and U9271 (N_9271,N_9064,N_9190);
nand U9272 (N_9272,N_9072,N_9118);
nand U9273 (N_9273,N_9246,N_9036);
nor U9274 (N_9274,N_9000,N_9111);
or U9275 (N_9275,N_9022,N_9079);
nor U9276 (N_9276,N_9021,N_9230);
or U9277 (N_9277,N_9228,N_9052);
xor U9278 (N_9278,N_9065,N_9183);
or U9279 (N_9279,N_9011,N_9216);
and U9280 (N_9280,N_9165,N_9058);
nor U9281 (N_9281,N_9213,N_9071);
nand U9282 (N_9282,N_9047,N_9229);
and U9283 (N_9283,N_9019,N_9224);
nand U9284 (N_9284,N_9220,N_9141);
xnor U9285 (N_9285,N_9232,N_9122);
and U9286 (N_9286,N_9031,N_9221);
nor U9287 (N_9287,N_9090,N_9113);
nand U9288 (N_9288,N_9146,N_9226);
or U9289 (N_9289,N_9025,N_9170);
nand U9290 (N_9290,N_9243,N_9086);
or U9291 (N_9291,N_9208,N_9062);
nand U9292 (N_9292,N_9092,N_9042);
xnor U9293 (N_9293,N_9055,N_9008);
nor U9294 (N_9294,N_9248,N_9069);
xnor U9295 (N_9295,N_9152,N_9217);
and U9296 (N_9296,N_9006,N_9009);
and U9297 (N_9297,N_9164,N_9094);
xor U9298 (N_9298,N_9001,N_9097);
or U9299 (N_9299,N_9067,N_9214);
and U9300 (N_9300,N_9109,N_9057);
and U9301 (N_9301,N_9088,N_9017);
nand U9302 (N_9302,N_9119,N_9083);
xnor U9303 (N_9303,N_9212,N_9101);
nand U9304 (N_9304,N_9245,N_9020);
xor U9305 (N_9305,N_9219,N_9063);
or U9306 (N_9306,N_9049,N_9110);
nand U9307 (N_9307,N_9108,N_9180);
nor U9308 (N_9308,N_9028,N_9015);
or U9309 (N_9309,N_9048,N_9184);
xor U9310 (N_9310,N_9172,N_9162);
and U9311 (N_9311,N_9073,N_9237);
nand U9312 (N_9312,N_9197,N_9178);
nand U9313 (N_9313,N_9089,N_9241);
xnor U9314 (N_9314,N_9041,N_9023);
or U9315 (N_9315,N_9124,N_9167);
or U9316 (N_9316,N_9233,N_9247);
and U9317 (N_9317,N_9140,N_9091);
nand U9318 (N_9318,N_9193,N_9211);
nor U9319 (N_9319,N_9234,N_9099);
and U9320 (N_9320,N_9147,N_9084);
xor U9321 (N_9321,N_9225,N_9161);
nand U9322 (N_9322,N_9240,N_9045);
xnor U9323 (N_9323,N_9127,N_9151);
and U9324 (N_9324,N_9061,N_9175);
and U9325 (N_9325,N_9034,N_9231);
nand U9326 (N_9326,N_9207,N_9205);
nor U9327 (N_9327,N_9150,N_9035);
nand U9328 (N_9328,N_9238,N_9195);
or U9329 (N_9329,N_9242,N_9218);
and U9330 (N_9330,N_9181,N_9116);
nor U9331 (N_9331,N_9153,N_9051);
nor U9332 (N_9332,N_9010,N_9030);
and U9333 (N_9333,N_9098,N_9177);
and U9334 (N_9334,N_9080,N_9074);
and U9335 (N_9335,N_9027,N_9134);
xor U9336 (N_9336,N_9209,N_9173);
nor U9337 (N_9337,N_9199,N_9085);
and U9338 (N_9338,N_9222,N_9012);
xor U9339 (N_9339,N_9026,N_9133);
or U9340 (N_9340,N_9235,N_9056);
nor U9341 (N_9341,N_9013,N_9107);
nor U9342 (N_9342,N_9163,N_9179);
or U9343 (N_9343,N_9157,N_9077);
and U9344 (N_9344,N_9018,N_9082);
xor U9345 (N_9345,N_9148,N_9206);
nor U9346 (N_9346,N_9142,N_9044);
or U9347 (N_9347,N_9249,N_9046);
nand U9348 (N_9348,N_9039,N_9198);
or U9349 (N_9349,N_9076,N_9132);
nand U9350 (N_9350,N_9139,N_9126);
xor U9351 (N_9351,N_9159,N_9078);
nand U9352 (N_9352,N_9223,N_9053);
nand U9353 (N_9353,N_9166,N_9125);
nand U9354 (N_9354,N_9037,N_9137);
nand U9355 (N_9355,N_9186,N_9185);
and U9356 (N_9356,N_9182,N_9144);
or U9357 (N_9357,N_9121,N_9024);
nor U9358 (N_9358,N_9158,N_9014);
nand U9359 (N_9359,N_9200,N_9149);
xnor U9360 (N_9360,N_9143,N_9156);
nor U9361 (N_9361,N_9130,N_9145);
nand U9362 (N_9362,N_9007,N_9154);
or U9363 (N_9363,N_9176,N_9239);
nor U9364 (N_9364,N_9096,N_9016);
xor U9365 (N_9365,N_9068,N_9191);
and U9366 (N_9366,N_9003,N_9227);
or U9367 (N_9367,N_9135,N_9060);
nor U9368 (N_9368,N_9005,N_9004);
xnor U9369 (N_9369,N_9136,N_9050);
nor U9370 (N_9370,N_9189,N_9106);
nand U9371 (N_9371,N_9236,N_9117);
or U9372 (N_9372,N_9002,N_9059);
nand U9373 (N_9373,N_9192,N_9095);
nor U9374 (N_9374,N_9114,N_9131);
nor U9375 (N_9375,N_9236,N_9084);
nor U9376 (N_9376,N_9041,N_9224);
xor U9377 (N_9377,N_9018,N_9194);
xnor U9378 (N_9378,N_9183,N_9086);
or U9379 (N_9379,N_9189,N_9170);
nand U9380 (N_9380,N_9112,N_9010);
and U9381 (N_9381,N_9217,N_9190);
or U9382 (N_9382,N_9132,N_9195);
nor U9383 (N_9383,N_9075,N_9220);
and U9384 (N_9384,N_9209,N_9176);
nor U9385 (N_9385,N_9248,N_9096);
or U9386 (N_9386,N_9175,N_9139);
nand U9387 (N_9387,N_9117,N_9220);
or U9388 (N_9388,N_9195,N_9114);
nand U9389 (N_9389,N_9008,N_9014);
nor U9390 (N_9390,N_9246,N_9067);
nor U9391 (N_9391,N_9179,N_9100);
or U9392 (N_9392,N_9036,N_9154);
or U9393 (N_9393,N_9173,N_9160);
nand U9394 (N_9394,N_9176,N_9106);
nand U9395 (N_9395,N_9138,N_9181);
nand U9396 (N_9396,N_9216,N_9185);
xor U9397 (N_9397,N_9217,N_9067);
or U9398 (N_9398,N_9081,N_9095);
and U9399 (N_9399,N_9162,N_9040);
and U9400 (N_9400,N_9181,N_9106);
and U9401 (N_9401,N_9076,N_9242);
or U9402 (N_9402,N_9229,N_9091);
and U9403 (N_9403,N_9035,N_9208);
or U9404 (N_9404,N_9104,N_9091);
xnor U9405 (N_9405,N_9155,N_9096);
or U9406 (N_9406,N_9205,N_9224);
nor U9407 (N_9407,N_9180,N_9010);
and U9408 (N_9408,N_9182,N_9006);
or U9409 (N_9409,N_9160,N_9215);
and U9410 (N_9410,N_9162,N_9072);
or U9411 (N_9411,N_9166,N_9021);
and U9412 (N_9412,N_9213,N_9155);
nor U9413 (N_9413,N_9102,N_9210);
nor U9414 (N_9414,N_9135,N_9236);
nand U9415 (N_9415,N_9176,N_9105);
xnor U9416 (N_9416,N_9187,N_9237);
or U9417 (N_9417,N_9049,N_9007);
or U9418 (N_9418,N_9133,N_9046);
nand U9419 (N_9419,N_9158,N_9119);
nor U9420 (N_9420,N_9091,N_9224);
xor U9421 (N_9421,N_9201,N_9240);
nand U9422 (N_9422,N_9205,N_9059);
nand U9423 (N_9423,N_9024,N_9155);
nand U9424 (N_9424,N_9014,N_9212);
and U9425 (N_9425,N_9100,N_9045);
nand U9426 (N_9426,N_9144,N_9020);
nor U9427 (N_9427,N_9228,N_9029);
nand U9428 (N_9428,N_9242,N_9130);
xor U9429 (N_9429,N_9082,N_9078);
nand U9430 (N_9430,N_9119,N_9029);
nor U9431 (N_9431,N_9108,N_9094);
or U9432 (N_9432,N_9234,N_9176);
xnor U9433 (N_9433,N_9090,N_9162);
or U9434 (N_9434,N_9093,N_9014);
nor U9435 (N_9435,N_9058,N_9039);
nand U9436 (N_9436,N_9038,N_9186);
or U9437 (N_9437,N_9221,N_9092);
nand U9438 (N_9438,N_9126,N_9108);
xnor U9439 (N_9439,N_9011,N_9031);
or U9440 (N_9440,N_9152,N_9087);
or U9441 (N_9441,N_9133,N_9234);
nand U9442 (N_9442,N_9136,N_9074);
xor U9443 (N_9443,N_9228,N_9089);
nand U9444 (N_9444,N_9117,N_9141);
nor U9445 (N_9445,N_9170,N_9218);
xor U9446 (N_9446,N_9099,N_9201);
or U9447 (N_9447,N_9059,N_9167);
or U9448 (N_9448,N_9221,N_9107);
or U9449 (N_9449,N_9032,N_9097);
or U9450 (N_9450,N_9023,N_9192);
or U9451 (N_9451,N_9162,N_9077);
xnor U9452 (N_9452,N_9128,N_9149);
xnor U9453 (N_9453,N_9242,N_9111);
nor U9454 (N_9454,N_9033,N_9196);
and U9455 (N_9455,N_9222,N_9216);
or U9456 (N_9456,N_9068,N_9188);
and U9457 (N_9457,N_9053,N_9173);
or U9458 (N_9458,N_9005,N_9128);
and U9459 (N_9459,N_9228,N_9056);
xnor U9460 (N_9460,N_9136,N_9057);
or U9461 (N_9461,N_9248,N_9177);
and U9462 (N_9462,N_9132,N_9218);
or U9463 (N_9463,N_9097,N_9103);
nor U9464 (N_9464,N_9096,N_9231);
and U9465 (N_9465,N_9111,N_9236);
or U9466 (N_9466,N_9210,N_9145);
and U9467 (N_9467,N_9096,N_9199);
xor U9468 (N_9468,N_9145,N_9229);
nor U9469 (N_9469,N_9090,N_9233);
nand U9470 (N_9470,N_9166,N_9042);
nand U9471 (N_9471,N_9218,N_9068);
and U9472 (N_9472,N_9011,N_9206);
xor U9473 (N_9473,N_9158,N_9223);
xor U9474 (N_9474,N_9156,N_9023);
xnor U9475 (N_9475,N_9232,N_9084);
or U9476 (N_9476,N_9164,N_9055);
xor U9477 (N_9477,N_9112,N_9075);
or U9478 (N_9478,N_9138,N_9061);
xor U9479 (N_9479,N_9149,N_9219);
xor U9480 (N_9480,N_9055,N_9176);
and U9481 (N_9481,N_9197,N_9189);
nand U9482 (N_9482,N_9049,N_9022);
nor U9483 (N_9483,N_9222,N_9090);
xnor U9484 (N_9484,N_9018,N_9037);
or U9485 (N_9485,N_9087,N_9190);
or U9486 (N_9486,N_9020,N_9130);
xnor U9487 (N_9487,N_9000,N_9053);
or U9488 (N_9488,N_9005,N_9000);
nand U9489 (N_9489,N_9169,N_9014);
nor U9490 (N_9490,N_9058,N_9183);
nand U9491 (N_9491,N_9080,N_9121);
and U9492 (N_9492,N_9098,N_9076);
xor U9493 (N_9493,N_9135,N_9196);
nor U9494 (N_9494,N_9137,N_9157);
or U9495 (N_9495,N_9083,N_9216);
or U9496 (N_9496,N_9042,N_9156);
nand U9497 (N_9497,N_9180,N_9042);
nor U9498 (N_9498,N_9138,N_9174);
nand U9499 (N_9499,N_9044,N_9119);
or U9500 (N_9500,N_9309,N_9422);
nand U9501 (N_9501,N_9417,N_9280);
nand U9502 (N_9502,N_9390,N_9394);
xnor U9503 (N_9503,N_9263,N_9445);
xor U9504 (N_9504,N_9452,N_9456);
nor U9505 (N_9505,N_9400,N_9382);
and U9506 (N_9506,N_9478,N_9260);
and U9507 (N_9507,N_9454,N_9251);
and U9508 (N_9508,N_9277,N_9285);
nand U9509 (N_9509,N_9250,N_9471);
nand U9510 (N_9510,N_9377,N_9376);
xor U9511 (N_9511,N_9428,N_9396);
nor U9512 (N_9512,N_9437,N_9499);
xnor U9513 (N_9513,N_9397,N_9365);
xnor U9514 (N_9514,N_9259,N_9385);
nor U9515 (N_9515,N_9279,N_9322);
and U9516 (N_9516,N_9481,N_9436);
and U9517 (N_9517,N_9367,N_9342);
and U9518 (N_9518,N_9393,N_9283);
and U9519 (N_9519,N_9266,N_9363);
or U9520 (N_9520,N_9380,N_9496);
nor U9521 (N_9521,N_9387,N_9371);
nand U9522 (N_9522,N_9491,N_9401);
nand U9523 (N_9523,N_9489,N_9355);
and U9524 (N_9524,N_9483,N_9281);
and U9525 (N_9525,N_9440,N_9340);
nor U9526 (N_9526,N_9423,N_9354);
and U9527 (N_9527,N_9271,N_9378);
and U9528 (N_9528,N_9439,N_9357);
xnor U9529 (N_9529,N_9392,N_9487);
or U9530 (N_9530,N_9461,N_9414);
or U9531 (N_9531,N_9264,N_9288);
and U9532 (N_9532,N_9362,N_9446);
nand U9533 (N_9533,N_9448,N_9465);
and U9534 (N_9534,N_9399,N_9389);
or U9535 (N_9535,N_9284,N_9408);
nor U9536 (N_9536,N_9334,N_9457);
and U9537 (N_9537,N_9438,N_9493);
or U9538 (N_9538,N_9300,N_9484);
nand U9539 (N_9539,N_9391,N_9314);
xnor U9540 (N_9540,N_9412,N_9292);
nor U9541 (N_9541,N_9435,N_9459);
and U9542 (N_9542,N_9287,N_9337);
xor U9543 (N_9543,N_9336,N_9282);
nor U9544 (N_9544,N_9286,N_9321);
or U9545 (N_9545,N_9326,N_9482);
nor U9546 (N_9546,N_9498,N_9419);
nor U9547 (N_9547,N_9324,N_9333);
nor U9548 (N_9548,N_9290,N_9274);
xor U9549 (N_9549,N_9494,N_9407);
or U9550 (N_9550,N_9318,N_9313);
or U9551 (N_9551,N_9303,N_9375);
or U9552 (N_9552,N_9455,N_9479);
or U9553 (N_9553,N_9298,N_9254);
xnor U9554 (N_9554,N_9386,N_9291);
or U9555 (N_9555,N_9403,N_9449);
xnor U9556 (N_9556,N_9344,N_9372);
and U9557 (N_9557,N_9364,N_9405);
or U9558 (N_9558,N_9335,N_9262);
nor U9559 (N_9559,N_9307,N_9270);
nand U9560 (N_9560,N_9466,N_9480);
nor U9561 (N_9561,N_9325,N_9346);
and U9562 (N_9562,N_9299,N_9488);
nand U9563 (N_9563,N_9497,N_9312);
nand U9564 (N_9564,N_9383,N_9369);
xnor U9565 (N_9565,N_9268,N_9311);
and U9566 (N_9566,N_9370,N_9431);
xnor U9567 (N_9567,N_9304,N_9373);
or U9568 (N_9568,N_9442,N_9273);
and U9569 (N_9569,N_9305,N_9252);
or U9570 (N_9570,N_9433,N_9469);
xnor U9571 (N_9571,N_9495,N_9427);
or U9572 (N_9572,N_9257,N_9330);
and U9573 (N_9573,N_9265,N_9424);
nor U9574 (N_9574,N_9486,N_9297);
and U9575 (N_9575,N_9474,N_9310);
nor U9576 (N_9576,N_9490,N_9293);
nor U9577 (N_9577,N_9475,N_9315);
nor U9578 (N_9578,N_9352,N_9319);
nand U9579 (N_9579,N_9272,N_9295);
xnor U9580 (N_9580,N_9416,N_9413);
nor U9581 (N_9581,N_9443,N_9430);
xnor U9582 (N_9582,N_9356,N_9415);
nand U9583 (N_9583,N_9464,N_9381);
or U9584 (N_9584,N_9256,N_9294);
or U9585 (N_9585,N_9351,N_9366);
nand U9586 (N_9586,N_9429,N_9338);
and U9587 (N_9587,N_9349,N_9358);
xnor U9588 (N_9588,N_9331,N_9368);
nand U9589 (N_9589,N_9388,N_9398);
nand U9590 (N_9590,N_9451,N_9477);
nand U9591 (N_9591,N_9395,N_9341);
nor U9592 (N_9592,N_9406,N_9470);
xor U9593 (N_9593,N_9347,N_9306);
xor U9594 (N_9594,N_9261,N_9379);
nand U9595 (N_9595,N_9275,N_9434);
nand U9596 (N_9596,N_9345,N_9432);
nand U9597 (N_9597,N_9447,N_9276);
nor U9598 (N_9598,N_9289,N_9492);
and U9599 (N_9599,N_9402,N_9343);
or U9600 (N_9600,N_9374,N_9296);
nor U9601 (N_9601,N_9317,N_9426);
xor U9602 (N_9602,N_9332,N_9485);
nor U9603 (N_9603,N_9359,N_9278);
or U9604 (N_9604,N_9421,N_9302);
nand U9605 (N_9605,N_9460,N_9441);
or U9606 (N_9606,N_9410,N_9404);
xor U9607 (N_9607,N_9353,N_9350);
nand U9608 (N_9608,N_9255,N_9418);
nand U9609 (N_9609,N_9323,N_9467);
nor U9610 (N_9610,N_9339,N_9444);
xor U9611 (N_9611,N_9329,N_9462);
and U9612 (N_9612,N_9409,N_9269);
nor U9613 (N_9613,N_9328,N_9453);
nor U9614 (N_9614,N_9360,N_9472);
nand U9615 (N_9615,N_9308,N_9361);
nand U9616 (N_9616,N_9327,N_9316);
or U9617 (N_9617,N_9420,N_9253);
and U9618 (N_9618,N_9258,N_9267);
and U9619 (N_9619,N_9463,N_9450);
nand U9620 (N_9620,N_9468,N_9473);
or U9621 (N_9621,N_9301,N_9384);
and U9622 (N_9622,N_9348,N_9476);
nor U9623 (N_9623,N_9320,N_9411);
xor U9624 (N_9624,N_9458,N_9425);
nand U9625 (N_9625,N_9261,N_9481);
or U9626 (N_9626,N_9422,N_9429);
nand U9627 (N_9627,N_9465,N_9417);
and U9628 (N_9628,N_9498,N_9472);
xnor U9629 (N_9629,N_9413,N_9490);
nand U9630 (N_9630,N_9269,N_9403);
or U9631 (N_9631,N_9272,N_9488);
xor U9632 (N_9632,N_9446,N_9272);
and U9633 (N_9633,N_9321,N_9329);
xor U9634 (N_9634,N_9293,N_9287);
xnor U9635 (N_9635,N_9468,N_9426);
nand U9636 (N_9636,N_9326,N_9299);
and U9637 (N_9637,N_9278,N_9458);
nor U9638 (N_9638,N_9377,N_9483);
nand U9639 (N_9639,N_9426,N_9409);
nand U9640 (N_9640,N_9319,N_9347);
and U9641 (N_9641,N_9295,N_9492);
nand U9642 (N_9642,N_9422,N_9432);
and U9643 (N_9643,N_9302,N_9346);
nand U9644 (N_9644,N_9497,N_9315);
or U9645 (N_9645,N_9358,N_9448);
xnor U9646 (N_9646,N_9254,N_9289);
and U9647 (N_9647,N_9290,N_9442);
and U9648 (N_9648,N_9488,N_9254);
nor U9649 (N_9649,N_9357,N_9372);
or U9650 (N_9650,N_9491,N_9273);
nor U9651 (N_9651,N_9340,N_9376);
and U9652 (N_9652,N_9253,N_9440);
or U9653 (N_9653,N_9462,N_9336);
nand U9654 (N_9654,N_9380,N_9473);
xnor U9655 (N_9655,N_9401,N_9325);
and U9656 (N_9656,N_9483,N_9299);
nand U9657 (N_9657,N_9428,N_9285);
nand U9658 (N_9658,N_9311,N_9497);
nand U9659 (N_9659,N_9378,N_9284);
nand U9660 (N_9660,N_9280,N_9362);
nor U9661 (N_9661,N_9378,N_9343);
nand U9662 (N_9662,N_9346,N_9435);
or U9663 (N_9663,N_9435,N_9381);
nor U9664 (N_9664,N_9479,N_9368);
nand U9665 (N_9665,N_9292,N_9418);
xnor U9666 (N_9666,N_9270,N_9282);
and U9667 (N_9667,N_9461,N_9465);
nor U9668 (N_9668,N_9334,N_9336);
and U9669 (N_9669,N_9359,N_9306);
xor U9670 (N_9670,N_9410,N_9417);
nand U9671 (N_9671,N_9339,N_9430);
and U9672 (N_9672,N_9251,N_9481);
xnor U9673 (N_9673,N_9396,N_9487);
nor U9674 (N_9674,N_9442,N_9438);
or U9675 (N_9675,N_9313,N_9374);
nor U9676 (N_9676,N_9478,N_9335);
nand U9677 (N_9677,N_9461,N_9334);
or U9678 (N_9678,N_9299,N_9285);
and U9679 (N_9679,N_9259,N_9492);
and U9680 (N_9680,N_9444,N_9416);
nand U9681 (N_9681,N_9349,N_9497);
and U9682 (N_9682,N_9328,N_9349);
nand U9683 (N_9683,N_9454,N_9440);
nor U9684 (N_9684,N_9355,N_9378);
and U9685 (N_9685,N_9499,N_9307);
and U9686 (N_9686,N_9276,N_9412);
xor U9687 (N_9687,N_9257,N_9485);
xnor U9688 (N_9688,N_9403,N_9357);
and U9689 (N_9689,N_9282,N_9335);
or U9690 (N_9690,N_9340,N_9455);
and U9691 (N_9691,N_9301,N_9329);
nand U9692 (N_9692,N_9432,N_9258);
and U9693 (N_9693,N_9451,N_9289);
nor U9694 (N_9694,N_9463,N_9437);
xor U9695 (N_9695,N_9463,N_9434);
xnor U9696 (N_9696,N_9302,N_9365);
nand U9697 (N_9697,N_9353,N_9304);
nand U9698 (N_9698,N_9412,N_9452);
or U9699 (N_9699,N_9311,N_9341);
nor U9700 (N_9700,N_9316,N_9489);
nand U9701 (N_9701,N_9473,N_9366);
and U9702 (N_9702,N_9253,N_9409);
xnor U9703 (N_9703,N_9348,N_9336);
or U9704 (N_9704,N_9459,N_9291);
or U9705 (N_9705,N_9322,N_9420);
nor U9706 (N_9706,N_9329,N_9331);
or U9707 (N_9707,N_9434,N_9340);
and U9708 (N_9708,N_9295,N_9395);
or U9709 (N_9709,N_9480,N_9331);
nor U9710 (N_9710,N_9309,N_9360);
xor U9711 (N_9711,N_9398,N_9309);
nand U9712 (N_9712,N_9371,N_9276);
xnor U9713 (N_9713,N_9296,N_9475);
and U9714 (N_9714,N_9491,N_9315);
or U9715 (N_9715,N_9409,N_9259);
nor U9716 (N_9716,N_9461,N_9342);
or U9717 (N_9717,N_9481,N_9282);
or U9718 (N_9718,N_9428,N_9278);
nand U9719 (N_9719,N_9412,N_9330);
nor U9720 (N_9720,N_9468,N_9454);
xnor U9721 (N_9721,N_9417,N_9256);
xnor U9722 (N_9722,N_9484,N_9435);
nand U9723 (N_9723,N_9434,N_9265);
or U9724 (N_9724,N_9460,N_9443);
and U9725 (N_9725,N_9268,N_9468);
and U9726 (N_9726,N_9281,N_9319);
nand U9727 (N_9727,N_9427,N_9287);
nor U9728 (N_9728,N_9328,N_9323);
xor U9729 (N_9729,N_9317,N_9432);
or U9730 (N_9730,N_9346,N_9270);
xor U9731 (N_9731,N_9288,N_9422);
nand U9732 (N_9732,N_9270,N_9493);
and U9733 (N_9733,N_9441,N_9480);
nor U9734 (N_9734,N_9330,N_9316);
nand U9735 (N_9735,N_9366,N_9464);
and U9736 (N_9736,N_9285,N_9499);
nor U9737 (N_9737,N_9404,N_9377);
and U9738 (N_9738,N_9297,N_9391);
nand U9739 (N_9739,N_9276,N_9327);
or U9740 (N_9740,N_9474,N_9368);
nor U9741 (N_9741,N_9383,N_9476);
xnor U9742 (N_9742,N_9251,N_9366);
and U9743 (N_9743,N_9357,N_9446);
and U9744 (N_9744,N_9392,N_9385);
xnor U9745 (N_9745,N_9273,N_9270);
or U9746 (N_9746,N_9437,N_9257);
nand U9747 (N_9747,N_9334,N_9354);
and U9748 (N_9748,N_9281,N_9271);
nand U9749 (N_9749,N_9323,N_9498);
nor U9750 (N_9750,N_9711,N_9520);
or U9751 (N_9751,N_9543,N_9553);
nor U9752 (N_9752,N_9531,N_9588);
or U9753 (N_9753,N_9594,N_9592);
nor U9754 (N_9754,N_9534,N_9618);
nand U9755 (N_9755,N_9569,N_9736);
nor U9756 (N_9756,N_9686,N_9576);
and U9757 (N_9757,N_9586,N_9741);
and U9758 (N_9758,N_9591,N_9521);
nor U9759 (N_9759,N_9662,N_9734);
and U9760 (N_9760,N_9743,N_9615);
and U9761 (N_9761,N_9633,N_9682);
and U9762 (N_9762,N_9562,N_9705);
xor U9763 (N_9763,N_9696,N_9581);
nand U9764 (N_9764,N_9621,N_9637);
xnor U9765 (N_9765,N_9503,N_9720);
and U9766 (N_9766,N_9539,N_9599);
xnor U9767 (N_9767,N_9574,N_9676);
nand U9768 (N_9768,N_9693,N_9533);
nand U9769 (N_9769,N_9622,N_9642);
xnor U9770 (N_9770,N_9724,N_9738);
and U9771 (N_9771,N_9613,N_9578);
nand U9772 (N_9772,N_9607,N_9546);
or U9773 (N_9773,N_9611,N_9663);
or U9774 (N_9774,N_9744,N_9597);
or U9775 (N_9775,N_9629,N_9668);
nand U9776 (N_9776,N_9645,N_9502);
or U9777 (N_9777,N_9683,N_9679);
nor U9778 (N_9778,N_9602,N_9656);
or U9779 (N_9779,N_9589,N_9707);
nor U9780 (N_9780,N_9582,N_9598);
nor U9781 (N_9781,N_9567,N_9687);
xor U9782 (N_9782,N_9708,N_9623);
or U9783 (N_9783,N_9701,N_9745);
and U9784 (N_9784,N_9641,N_9530);
xor U9785 (N_9785,N_9665,N_9580);
nand U9786 (N_9786,N_9620,N_9700);
xnor U9787 (N_9787,N_9608,N_9517);
xnor U9788 (N_9788,N_9635,N_9625);
xnor U9789 (N_9789,N_9654,N_9575);
or U9790 (N_9790,N_9748,N_9699);
or U9791 (N_9791,N_9508,N_9630);
nor U9792 (N_9792,N_9747,N_9587);
xor U9793 (N_9793,N_9570,N_9674);
or U9794 (N_9794,N_9740,N_9609);
nor U9795 (N_9795,N_9703,N_9634);
xnor U9796 (N_9796,N_9566,N_9695);
nor U9797 (N_9797,N_9522,N_9524);
or U9798 (N_9798,N_9554,N_9712);
and U9799 (N_9799,N_9737,N_9704);
or U9800 (N_9800,N_9667,N_9512);
nor U9801 (N_9801,N_9706,N_9550);
xor U9802 (N_9802,N_9600,N_9643);
and U9803 (N_9803,N_9614,N_9639);
nor U9804 (N_9804,N_9518,N_9572);
nand U9805 (N_9805,N_9514,N_9713);
or U9806 (N_9806,N_9739,N_9593);
or U9807 (N_9807,N_9515,N_9505);
xor U9808 (N_9808,N_9544,N_9604);
or U9809 (N_9809,N_9525,N_9732);
nand U9810 (N_9810,N_9536,N_9547);
nor U9811 (N_9811,N_9722,N_9605);
xor U9812 (N_9812,N_9650,N_9673);
nor U9813 (N_9813,N_9549,N_9644);
xnor U9814 (N_9814,N_9649,N_9727);
or U9815 (N_9815,N_9681,N_9595);
nor U9816 (N_9816,N_9715,N_9532);
or U9817 (N_9817,N_9504,N_9661);
or U9818 (N_9818,N_9556,N_9551);
xnor U9819 (N_9819,N_9677,N_9612);
or U9820 (N_9820,N_9564,N_9717);
nor U9821 (N_9821,N_9716,N_9709);
nand U9822 (N_9822,N_9729,N_9728);
xnor U9823 (N_9823,N_9627,N_9718);
nor U9824 (N_9824,N_9610,N_9573);
and U9825 (N_9825,N_9684,N_9670);
and U9826 (N_9826,N_9601,N_9535);
nand U9827 (N_9827,N_9628,N_9733);
xnor U9828 (N_9828,N_9672,N_9555);
nand U9829 (N_9829,N_9640,N_9527);
and U9830 (N_9830,N_9606,N_9617);
nand U9831 (N_9831,N_9537,N_9568);
and U9832 (N_9832,N_9719,N_9690);
and U9833 (N_9833,N_9552,N_9660);
nor U9834 (N_9834,N_9730,N_9746);
and U9835 (N_9835,N_9710,N_9500);
nand U9836 (N_9836,N_9749,N_9565);
and U9837 (N_9837,N_9506,N_9528);
and U9838 (N_9838,N_9655,N_9584);
nand U9839 (N_9839,N_9742,N_9509);
and U9840 (N_9840,N_9511,N_9579);
xnor U9841 (N_9841,N_9638,N_9513);
nand U9842 (N_9842,N_9501,N_9726);
or U9843 (N_9843,N_9559,N_9735);
and U9844 (N_9844,N_9725,N_9590);
or U9845 (N_9845,N_9702,N_9697);
nand U9846 (N_9846,N_9563,N_9685);
and U9847 (N_9847,N_9510,N_9624);
and U9848 (N_9848,N_9653,N_9652);
xnor U9849 (N_9849,N_9666,N_9558);
nand U9850 (N_9850,N_9557,N_9659);
nand U9851 (N_9851,N_9688,N_9619);
nand U9852 (N_9852,N_9636,N_9664);
and U9853 (N_9853,N_9631,N_9669);
or U9854 (N_9854,N_9548,N_9577);
and U9855 (N_9855,N_9603,N_9538);
and U9856 (N_9856,N_9692,N_9585);
nand U9857 (N_9857,N_9675,N_9523);
or U9858 (N_9858,N_9671,N_9632);
or U9859 (N_9859,N_9583,N_9721);
nand U9860 (N_9860,N_9526,N_9596);
xnor U9861 (N_9861,N_9694,N_9646);
xor U9862 (N_9862,N_9651,N_9658);
and U9863 (N_9863,N_9519,N_9542);
nand U9864 (N_9864,N_9657,N_9529);
or U9865 (N_9865,N_9689,N_9507);
nand U9866 (N_9866,N_9561,N_9648);
xnor U9867 (N_9867,N_9647,N_9560);
nand U9868 (N_9868,N_9616,N_9678);
and U9869 (N_9869,N_9731,N_9723);
nand U9870 (N_9870,N_9626,N_9540);
or U9871 (N_9871,N_9571,N_9714);
nand U9872 (N_9872,N_9698,N_9541);
nor U9873 (N_9873,N_9545,N_9691);
xor U9874 (N_9874,N_9516,N_9680);
nand U9875 (N_9875,N_9724,N_9735);
nand U9876 (N_9876,N_9552,N_9548);
xor U9877 (N_9877,N_9566,N_9544);
nor U9878 (N_9878,N_9685,N_9696);
and U9879 (N_9879,N_9730,N_9502);
xor U9880 (N_9880,N_9722,N_9638);
nor U9881 (N_9881,N_9622,N_9723);
xnor U9882 (N_9882,N_9547,N_9559);
or U9883 (N_9883,N_9720,N_9592);
nand U9884 (N_9884,N_9608,N_9510);
nand U9885 (N_9885,N_9650,N_9550);
or U9886 (N_9886,N_9536,N_9533);
or U9887 (N_9887,N_9661,N_9643);
nand U9888 (N_9888,N_9733,N_9578);
and U9889 (N_9889,N_9573,N_9689);
and U9890 (N_9890,N_9659,N_9516);
and U9891 (N_9891,N_9711,N_9564);
nor U9892 (N_9892,N_9620,N_9689);
and U9893 (N_9893,N_9734,N_9680);
nand U9894 (N_9894,N_9655,N_9610);
or U9895 (N_9895,N_9714,N_9635);
nand U9896 (N_9896,N_9641,N_9537);
and U9897 (N_9897,N_9733,N_9722);
or U9898 (N_9898,N_9549,N_9573);
or U9899 (N_9899,N_9554,N_9577);
nor U9900 (N_9900,N_9719,N_9567);
and U9901 (N_9901,N_9658,N_9728);
or U9902 (N_9902,N_9523,N_9620);
xor U9903 (N_9903,N_9652,N_9627);
nand U9904 (N_9904,N_9631,N_9596);
xnor U9905 (N_9905,N_9635,N_9515);
or U9906 (N_9906,N_9501,N_9596);
nand U9907 (N_9907,N_9599,N_9526);
xor U9908 (N_9908,N_9612,N_9582);
or U9909 (N_9909,N_9640,N_9631);
nand U9910 (N_9910,N_9634,N_9632);
or U9911 (N_9911,N_9623,N_9539);
nand U9912 (N_9912,N_9641,N_9647);
nor U9913 (N_9913,N_9535,N_9502);
xor U9914 (N_9914,N_9612,N_9515);
and U9915 (N_9915,N_9543,N_9700);
and U9916 (N_9916,N_9509,N_9571);
nor U9917 (N_9917,N_9677,N_9515);
xor U9918 (N_9918,N_9615,N_9509);
nor U9919 (N_9919,N_9547,N_9530);
xnor U9920 (N_9920,N_9651,N_9673);
nor U9921 (N_9921,N_9647,N_9738);
xor U9922 (N_9922,N_9720,N_9717);
nor U9923 (N_9923,N_9658,N_9650);
nand U9924 (N_9924,N_9693,N_9634);
nand U9925 (N_9925,N_9672,N_9614);
xnor U9926 (N_9926,N_9559,N_9672);
or U9927 (N_9927,N_9652,N_9573);
or U9928 (N_9928,N_9587,N_9731);
xnor U9929 (N_9929,N_9510,N_9543);
xnor U9930 (N_9930,N_9713,N_9731);
nor U9931 (N_9931,N_9525,N_9589);
xor U9932 (N_9932,N_9660,N_9527);
xnor U9933 (N_9933,N_9590,N_9569);
nor U9934 (N_9934,N_9703,N_9626);
or U9935 (N_9935,N_9597,N_9643);
nand U9936 (N_9936,N_9569,N_9579);
xor U9937 (N_9937,N_9692,N_9731);
nor U9938 (N_9938,N_9543,N_9545);
and U9939 (N_9939,N_9625,N_9628);
xnor U9940 (N_9940,N_9617,N_9722);
nor U9941 (N_9941,N_9730,N_9694);
xnor U9942 (N_9942,N_9671,N_9733);
nor U9943 (N_9943,N_9503,N_9654);
nand U9944 (N_9944,N_9524,N_9630);
xnor U9945 (N_9945,N_9581,N_9558);
or U9946 (N_9946,N_9710,N_9729);
or U9947 (N_9947,N_9615,N_9740);
nand U9948 (N_9948,N_9673,N_9547);
or U9949 (N_9949,N_9536,N_9594);
and U9950 (N_9950,N_9719,N_9515);
or U9951 (N_9951,N_9694,N_9510);
nor U9952 (N_9952,N_9690,N_9650);
nand U9953 (N_9953,N_9625,N_9734);
nand U9954 (N_9954,N_9608,N_9601);
xor U9955 (N_9955,N_9611,N_9503);
and U9956 (N_9956,N_9689,N_9731);
and U9957 (N_9957,N_9691,N_9681);
xnor U9958 (N_9958,N_9556,N_9654);
nand U9959 (N_9959,N_9599,N_9689);
nor U9960 (N_9960,N_9704,N_9547);
and U9961 (N_9961,N_9638,N_9746);
nand U9962 (N_9962,N_9688,N_9618);
or U9963 (N_9963,N_9676,N_9630);
nor U9964 (N_9964,N_9591,N_9510);
nor U9965 (N_9965,N_9688,N_9653);
or U9966 (N_9966,N_9693,N_9737);
nor U9967 (N_9967,N_9632,N_9546);
nor U9968 (N_9968,N_9546,N_9553);
xor U9969 (N_9969,N_9548,N_9571);
nor U9970 (N_9970,N_9502,N_9550);
or U9971 (N_9971,N_9597,N_9505);
or U9972 (N_9972,N_9653,N_9647);
nor U9973 (N_9973,N_9665,N_9556);
nor U9974 (N_9974,N_9580,N_9544);
and U9975 (N_9975,N_9557,N_9649);
xor U9976 (N_9976,N_9697,N_9592);
and U9977 (N_9977,N_9514,N_9524);
nand U9978 (N_9978,N_9558,N_9570);
and U9979 (N_9979,N_9539,N_9584);
nand U9980 (N_9980,N_9555,N_9505);
nand U9981 (N_9981,N_9731,N_9520);
and U9982 (N_9982,N_9543,N_9544);
xnor U9983 (N_9983,N_9505,N_9728);
xor U9984 (N_9984,N_9555,N_9576);
nor U9985 (N_9985,N_9663,N_9744);
xor U9986 (N_9986,N_9564,N_9682);
or U9987 (N_9987,N_9593,N_9566);
xnor U9988 (N_9988,N_9568,N_9640);
nand U9989 (N_9989,N_9691,N_9524);
nand U9990 (N_9990,N_9691,N_9680);
nor U9991 (N_9991,N_9557,N_9601);
xor U9992 (N_9992,N_9732,N_9644);
or U9993 (N_9993,N_9574,N_9630);
xnor U9994 (N_9994,N_9652,N_9527);
nor U9995 (N_9995,N_9529,N_9614);
nand U9996 (N_9996,N_9588,N_9740);
and U9997 (N_9997,N_9554,N_9656);
nor U9998 (N_9998,N_9526,N_9610);
or U9999 (N_9999,N_9624,N_9542);
or U10000 (N_10000,N_9800,N_9868);
xnor U10001 (N_10001,N_9825,N_9924);
nand U10002 (N_10002,N_9981,N_9834);
nor U10003 (N_10003,N_9956,N_9859);
or U10004 (N_10004,N_9842,N_9758);
and U10005 (N_10005,N_9880,N_9887);
and U10006 (N_10006,N_9870,N_9847);
or U10007 (N_10007,N_9909,N_9864);
nor U10008 (N_10008,N_9942,N_9939);
nand U10009 (N_10009,N_9986,N_9934);
nor U10010 (N_10010,N_9879,N_9994);
nand U10011 (N_10011,N_9849,N_9788);
xor U10012 (N_10012,N_9972,N_9973);
nor U10013 (N_10013,N_9894,N_9941);
xor U10014 (N_10014,N_9971,N_9872);
and U10015 (N_10015,N_9853,N_9767);
nor U10016 (N_10016,N_9888,N_9764);
nand U10017 (N_10017,N_9759,N_9836);
or U10018 (N_10018,N_9866,N_9858);
xnor U10019 (N_10019,N_9773,N_9821);
and U10020 (N_10020,N_9856,N_9768);
or U10021 (N_10021,N_9938,N_9948);
nand U10022 (N_10022,N_9962,N_9835);
and U10023 (N_10023,N_9782,N_9996);
and U10024 (N_10024,N_9969,N_9937);
xor U10025 (N_10025,N_9976,N_9995);
xor U10026 (N_10026,N_9807,N_9947);
nor U10027 (N_10027,N_9778,N_9829);
and U10028 (N_10028,N_9885,N_9926);
xnor U10029 (N_10029,N_9774,N_9997);
xor U10030 (N_10030,N_9755,N_9979);
nor U10031 (N_10031,N_9891,N_9884);
or U10032 (N_10032,N_9918,N_9946);
xnor U10033 (N_10033,N_9812,N_9935);
or U10034 (N_10034,N_9786,N_9832);
xnor U10035 (N_10035,N_9913,N_9878);
nand U10036 (N_10036,N_9865,N_9968);
nor U10037 (N_10037,N_9923,N_9988);
and U10038 (N_10038,N_9949,N_9895);
nand U10039 (N_10039,N_9809,N_9910);
nor U10040 (N_10040,N_9876,N_9945);
or U10041 (N_10041,N_9780,N_9857);
nor U10042 (N_10042,N_9925,N_9933);
and U10043 (N_10043,N_9796,N_9890);
and U10044 (N_10044,N_9801,N_9823);
nand U10045 (N_10045,N_9882,N_9843);
or U10046 (N_10046,N_9792,N_9966);
nand U10047 (N_10047,N_9898,N_9958);
or U10048 (N_10048,N_9911,N_9928);
nand U10049 (N_10049,N_9874,N_9803);
or U10050 (N_10050,N_9756,N_9959);
and U10051 (N_10051,N_9932,N_9920);
xnor U10052 (N_10052,N_9751,N_9804);
nand U10053 (N_10053,N_9886,N_9815);
and U10054 (N_10054,N_9875,N_9952);
or U10055 (N_10055,N_9833,N_9819);
nor U10056 (N_10056,N_9760,N_9987);
xnor U10057 (N_10057,N_9787,N_9921);
nand U10058 (N_10058,N_9953,N_9850);
and U10059 (N_10059,N_9810,N_9827);
nor U10060 (N_10060,N_9783,N_9776);
or U10061 (N_10061,N_9957,N_9960);
xnor U10062 (N_10062,N_9944,N_9862);
and U10063 (N_10063,N_9839,N_9917);
nor U10064 (N_10064,N_9816,N_9845);
or U10065 (N_10065,N_9838,N_9769);
nor U10066 (N_10066,N_9931,N_9813);
or U10067 (N_10067,N_9817,N_9900);
or U10068 (N_10068,N_9989,N_9936);
or U10069 (N_10069,N_9795,N_9855);
xnor U10070 (N_10070,N_9848,N_9974);
nand U10071 (N_10071,N_9781,N_9943);
nor U10072 (N_10072,N_9808,N_9922);
xor U10073 (N_10073,N_9970,N_9984);
nor U10074 (N_10074,N_9919,N_9790);
nor U10075 (N_10075,N_9975,N_9791);
nand U10076 (N_10076,N_9770,N_9861);
nor U10077 (N_10077,N_9914,N_9761);
nand U10078 (N_10078,N_9784,N_9798);
xor U10079 (N_10079,N_9982,N_9951);
nor U10080 (N_10080,N_9963,N_9901);
and U10081 (N_10081,N_9852,N_9955);
and U10082 (N_10082,N_9851,N_9822);
nand U10083 (N_10083,N_9814,N_9867);
nor U10084 (N_10084,N_9820,N_9753);
nand U10085 (N_10085,N_9828,N_9954);
and U10086 (N_10086,N_9883,N_9991);
nand U10087 (N_10087,N_9837,N_9830);
xor U10088 (N_10088,N_9779,N_9775);
nor U10089 (N_10089,N_9765,N_9992);
or U10090 (N_10090,N_9762,N_9860);
or U10091 (N_10091,N_9785,N_9802);
and U10092 (N_10092,N_9896,N_9877);
or U10093 (N_10093,N_9998,N_9927);
or U10094 (N_10094,N_9916,N_9754);
xor U10095 (N_10095,N_9950,N_9840);
xor U10096 (N_10096,N_9965,N_9863);
and U10097 (N_10097,N_9772,N_9805);
and U10098 (N_10098,N_9899,N_9818);
nor U10099 (N_10099,N_9797,N_9752);
xnor U10100 (N_10100,N_9854,N_9881);
and U10101 (N_10101,N_9831,N_9967);
nand U10102 (N_10102,N_9766,N_9869);
and U10103 (N_10103,N_9844,N_9824);
nor U10104 (N_10104,N_9897,N_9893);
and U10105 (N_10105,N_9799,N_9908);
nor U10106 (N_10106,N_9912,N_9841);
or U10107 (N_10107,N_9794,N_9929);
nand U10108 (N_10108,N_9806,N_9905);
xnor U10109 (N_10109,N_9889,N_9930);
nor U10110 (N_10110,N_9811,N_9980);
or U10111 (N_10111,N_9993,N_9892);
nand U10112 (N_10112,N_9940,N_9871);
nor U10113 (N_10113,N_9990,N_9902);
xor U10114 (N_10114,N_9903,N_9907);
and U10115 (N_10115,N_9964,N_9983);
or U10116 (N_10116,N_9977,N_9873);
or U10117 (N_10117,N_9826,N_9750);
or U10118 (N_10118,N_9763,N_9777);
nand U10119 (N_10119,N_9793,N_9904);
and U10120 (N_10120,N_9906,N_9985);
and U10121 (N_10121,N_9757,N_9789);
nand U10122 (N_10122,N_9978,N_9999);
nor U10123 (N_10123,N_9961,N_9846);
nand U10124 (N_10124,N_9771,N_9915);
nand U10125 (N_10125,N_9890,N_9828);
nor U10126 (N_10126,N_9783,N_9932);
nor U10127 (N_10127,N_9826,N_9941);
and U10128 (N_10128,N_9812,N_9979);
nor U10129 (N_10129,N_9810,N_9941);
nor U10130 (N_10130,N_9764,N_9984);
nand U10131 (N_10131,N_9765,N_9943);
xor U10132 (N_10132,N_9836,N_9863);
xnor U10133 (N_10133,N_9786,N_9951);
or U10134 (N_10134,N_9868,N_9930);
and U10135 (N_10135,N_9991,N_9803);
nor U10136 (N_10136,N_9833,N_9761);
xor U10137 (N_10137,N_9923,N_9877);
and U10138 (N_10138,N_9947,N_9787);
or U10139 (N_10139,N_9915,N_9953);
nor U10140 (N_10140,N_9969,N_9977);
nor U10141 (N_10141,N_9831,N_9990);
or U10142 (N_10142,N_9841,N_9839);
nand U10143 (N_10143,N_9824,N_9884);
nand U10144 (N_10144,N_9794,N_9936);
or U10145 (N_10145,N_9837,N_9969);
or U10146 (N_10146,N_9785,N_9921);
nand U10147 (N_10147,N_9819,N_9878);
nand U10148 (N_10148,N_9965,N_9838);
or U10149 (N_10149,N_9798,N_9813);
nor U10150 (N_10150,N_9894,N_9793);
nand U10151 (N_10151,N_9778,N_9751);
nor U10152 (N_10152,N_9896,N_9902);
and U10153 (N_10153,N_9919,N_9970);
nand U10154 (N_10154,N_9997,N_9859);
or U10155 (N_10155,N_9770,N_9834);
and U10156 (N_10156,N_9771,N_9785);
nor U10157 (N_10157,N_9873,N_9788);
nor U10158 (N_10158,N_9993,N_9871);
or U10159 (N_10159,N_9783,N_9960);
nand U10160 (N_10160,N_9978,N_9974);
and U10161 (N_10161,N_9796,N_9874);
xnor U10162 (N_10162,N_9901,N_9825);
nor U10163 (N_10163,N_9916,N_9877);
and U10164 (N_10164,N_9924,N_9922);
xnor U10165 (N_10165,N_9784,N_9976);
xor U10166 (N_10166,N_9807,N_9825);
nor U10167 (N_10167,N_9764,N_9946);
xnor U10168 (N_10168,N_9981,N_9788);
nand U10169 (N_10169,N_9961,N_9980);
xor U10170 (N_10170,N_9753,N_9754);
nor U10171 (N_10171,N_9986,N_9989);
or U10172 (N_10172,N_9972,N_9781);
nand U10173 (N_10173,N_9895,N_9967);
xor U10174 (N_10174,N_9954,N_9792);
or U10175 (N_10175,N_9993,N_9970);
or U10176 (N_10176,N_9862,N_9941);
nand U10177 (N_10177,N_9804,N_9875);
and U10178 (N_10178,N_9750,N_9896);
nor U10179 (N_10179,N_9920,N_9819);
and U10180 (N_10180,N_9860,N_9922);
nor U10181 (N_10181,N_9954,N_9853);
nand U10182 (N_10182,N_9775,N_9926);
and U10183 (N_10183,N_9975,N_9771);
nand U10184 (N_10184,N_9942,N_9833);
or U10185 (N_10185,N_9773,N_9786);
nor U10186 (N_10186,N_9900,N_9781);
xnor U10187 (N_10187,N_9750,N_9779);
or U10188 (N_10188,N_9964,N_9789);
and U10189 (N_10189,N_9978,N_9964);
or U10190 (N_10190,N_9826,N_9883);
and U10191 (N_10191,N_9930,N_9756);
nor U10192 (N_10192,N_9920,N_9949);
nand U10193 (N_10193,N_9860,N_9803);
or U10194 (N_10194,N_9812,N_9894);
or U10195 (N_10195,N_9828,N_9794);
and U10196 (N_10196,N_9924,N_9884);
nor U10197 (N_10197,N_9899,N_9852);
or U10198 (N_10198,N_9894,N_9977);
or U10199 (N_10199,N_9800,N_9899);
and U10200 (N_10200,N_9967,N_9891);
or U10201 (N_10201,N_9931,N_9780);
nor U10202 (N_10202,N_9880,N_9920);
and U10203 (N_10203,N_9815,N_9868);
and U10204 (N_10204,N_9867,N_9872);
nand U10205 (N_10205,N_9800,N_9795);
nand U10206 (N_10206,N_9968,N_9893);
and U10207 (N_10207,N_9773,N_9754);
and U10208 (N_10208,N_9872,N_9966);
nand U10209 (N_10209,N_9865,N_9891);
xor U10210 (N_10210,N_9774,N_9888);
nor U10211 (N_10211,N_9904,N_9963);
nand U10212 (N_10212,N_9960,N_9886);
nor U10213 (N_10213,N_9816,N_9833);
nand U10214 (N_10214,N_9853,N_9888);
and U10215 (N_10215,N_9753,N_9768);
nor U10216 (N_10216,N_9867,N_9925);
and U10217 (N_10217,N_9758,N_9754);
and U10218 (N_10218,N_9984,N_9954);
or U10219 (N_10219,N_9945,N_9798);
or U10220 (N_10220,N_9921,N_9810);
nor U10221 (N_10221,N_9758,N_9858);
nand U10222 (N_10222,N_9907,N_9981);
or U10223 (N_10223,N_9779,N_9755);
nand U10224 (N_10224,N_9929,N_9810);
nand U10225 (N_10225,N_9793,N_9914);
nor U10226 (N_10226,N_9876,N_9824);
xor U10227 (N_10227,N_9870,N_9787);
nand U10228 (N_10228,N_9863,N_9786);
or U10229 (N_10229,N_9958,N_9914);
and U10230 (N_10230,N_9773,N_9994);
nor U10231 (N_10231,N_9956,N_9772);
xnor U10232 (N_10232,N_9968,N_9950);
xnor U10233 (N_10233,N_9810,N_9886);
nand U10234 (N_10234,N_9893,N_9915);
nor U10235 (N_10235,N_9984,N_9995);
and U10236 (N_10236,N_9801,N_9891);
or U10237 (N_10237,N_9859,N_9899);
xnor U10238 (N_10238,N_9855,N_9821);
nor U10239 (N_10239,N_9792,N_9920);
nor U10240 (N_10240,N_9935,N_9957);
nor U10241 (N_10241,N_9799,N_9842);
nor U10242 (N_10242,N_9751,N_9892);
xor U10243 (N_10243,N_9814,N_9907);
or U10244 (N_10244,N_9816,N_9805);
and U10245 (N_10245,N_9778,N_9816);
and U10246 (N_10246,N_9815,N_9811);
and U10247 (N_10247,N_9763,N_9950);
nand U10248 (N_10248,N_9830,N_9944);
and U10249 (N_10249,N_9810,N_9845);
or U10250 (N_10250,N_10181,N_10084);
nor U10251 (N_10251,N_10225,N_10151);
or U10252 (N_10252,N_10071,N_10247);
nand U10253 (N_10253,N_10104,N_10092);
xor U10254 (N_10254,N_10055,N_10143);
nand U10255 (N_10255,N_10230,N_10050);
and U10256 (N_10256,N_10034,N_10097);
xor U10257 (N_10257,N_10188,N_10073);
xnor U10258 (N_10258,N_10138,N_10124);
or U10259 (N_10259,N_10173,N_10194);
nand U10260 (N_10260,N_10160,N_10117);
nor U10261 (N_10261,N_10053,N_10171);
nand U10262 (N_10262,N_10113,N_10003);
nand U10263 (N_10263,N_10129,N_10144);
nand U10264 (N_10264,N_10083,N_10208);
nor U10265 (N_10265,N_10169,N_10079);
xnor U10266 (N_10266,N_10018,N_10014);
nor U10267 (N_10267,N_10044,N_10091);
and U10268 (N_10268,N_10161,N_10217);
nor U10269 (N_10269,N_10037,N_10075);
nor U10270 (N_10270,N_10038,N_10226);
nor U10271 (N_10271,N_10004,N_10158);
nand U10272 (N_10272,N_10146,N_10140);
nor U10273 (N_10273,N_10135,N_10043);
or U10274 (N_10274,N_10166,N_10235);
nor U10275 (N_10275,N_10072,N_10116);
xor U10276 (N_10276,N_10076,N_10110);
xnor U10277 (N_10277,N_10216,N_10179);
or U10278 (N_10278,N_10148,N_10047);
and U10279 (N_10279,N_10224,N_10157);
nand U10280 (N_10280,N_10105,N_10036);
nand U10281 (N_10281,N_10085,N_10021);
nor U10282 (N_10282,N_10184,N_10039);
nor U10283 (N_10283,N_10081,N_10142);
or U10284 (N_10284,N_10139,N_10199);
xor U10285 (N_10285,N_10098,N_10243);
xor U10286 (N_10286,N_10242,N_10249);
nand U10287 (N_10287,N_10177,N_10219);
nand U10288 (N_10288,N_10193,N_10220);
nor U10289 (N_10289,N_10115,N_10172);
or U10290 (N_10290,N_10095,N_10229);
or U10291 (N_10291,N_10223,N_10245);
nand U10292 (N_10292,N_10012,N_10168);
or U10293 (N_10293,N_10145,N_10125);
and U10294 (N_10294,N_10241,N_10227);
and U10295 (N_10295,N_10048,N_10207);
nand U10296 (N_10296,N_10137,N_10213);
nor U10297 (N_10297,N_10045,N_10127);
xor U10298 (N_10298,N_10074,N_10154);
and U10299 (N_10299,N_10210,N_10130);
nor U10300 (N_10300,N_10093,N_10244);
and U10301 (N_10301,N_10035,N_10164);
nor U10302 (N_10302,N_10159,N_10052);
and U10303 (N_10303,N_10100,N_10101);
nand U10304 (N_10304,N_10096,N_10061);
and U10305 (N_10305,N_10011,N_10180);
xor U10306 (N_10306,N_10109,N_10186);
or U10307 (N_10307,N_10212,N_10010);
nor U10308 (N_10308,N_10002,N_10240);
nor U10309 (N_10309,N_10106,N_10060);
nand U10310 (N_10310,N_10024,N_10078);
xnor U10311 (N_10311,N_10183,N_10228);
nand U10312 (N_10312,N_10178,N_10232);
xor U10313 (N_10313,N_10058,N_10202);
or U10314 (N_10314,N_10205,N_10068);
or U10315 (N_10315,N_10119,N_10167);
nor U10316 (N_10316,N_10248,N_10017);
and U10317 (N_10317,N_10170,N_10112);
or U10318 (N_10318,N_10136,N_10046);
nor U10319 (N_10319,N_10118,N_10218);
nand U10320 (N_10320,N_10040,N_10132);
xnor U10321 (N_10321,N_10201,N_10111);
nor U10322 (N_10322,N_10114,N_10153);
nand U10323 (N_10323,N_10051,N_10057);
nand U10324 (N_10324,N_10175,N_10238);
or U10325 (N_10325,N_10203,N_10088);
xor U10326 (N_10326,N_10214,N_10233);
and U10327 (N_10327,N_10102,N_10000);
nand U10328 (N_10328,N_10077,N_10067);
xor U10329 (N_10329,N_10182,N_10231);
nand U10330 (N_10330,N_10086,N_10094);
nor U10331 (N_10331,N_10070,N_10246);
or U10332 (N_10332,N_10222,N_10192);
nand U10333 (N_10333,N_10056,N_10023);
or U10334 (N_10334,N_10197,N_10033);
or U10335 (N_10335,N_10195,N_10019);
or U10336 (N_10336,N_10082,N_10156);
nor U10337 (N_10337,N_10090,N_10028);
nor U10338 (N_10338,N_10099,N_10121);
nand U10339 (N_10339,N_10089,N_10031);
xnor U10340 (N_10340,N_10041,N_10131);
or U10341 (N_10341,N_10234,N_10027);
nand U10342 (N_10342,N_10025,N_10087);
or U10343 (N_10343,N_10063,N_10128);
or U10344 (N_10344,N_10126,N_10065);
or U10345 (N_10345,N_10133,N_10064);
or U10346 (N_10346,N_10069,N_10141);
nand U10347 (N_10347,N_10054,N_10009);
or U10348 (N_10348,N_10108,N_10221);
nand U10349 (N_10349,N_10174,N_10215);
and U10350 (N_10350,N_10236,N_10007);
nand U10351 (N_10351,N_10029,N_10107);
xnor U10352 (N_10352,N_10200,N_10165);
or U10353 (N_10353,N_10015,N_10062);
xor U10354 (N_10354,N_10122,N_10198);
and U10355 (N_10355,N_10080,N_10211);
nor U10356 (N_10356,N_10020,N_10134);
or U10357 (N_10357,N_10032,N_10155);
nor U10358 (N_10358,N_10013,N_10190);
and U10359 (N_10359,N_10189,N_10026);
nand U10360 (N_10360,N_10059,N_10006);
nor U10361 (N_10361,N_10206,N_10196);
nand U10362 (N_10362,N_10049,N_10150);
xnor U10363 (N_10363,N_10209,N_10239);
or U10364 (N_10364,N_10185,N_10005);
nor U10365 (N_10365,N_10163,N_10123);
and U10366 (N_10366,N_10030,N_10022);
nand U10367 (N_10367,N_10001,N_10149);
or U10368 (N_10368,N_10204,N_10103);
nor U10369 (N_10369,N_10066,N_10016);
nor U10370 (N_10370,N_10147,N_10237);
nor U10371 (N_10371,N_10176,N_10162);
nand U10372 (N_10372,N_10187,N_10191);
or U10373 (N_10373,N_10120,N_10152);
xnor U10374 (N_10374,N_10008,N_10042);
and U10375 (N_10375,N_10082,N_10094);
xnor U10376 (N_10376,N_10059,N_10037);
nand U10377 (N_10377,N_10062,N_10221);
nand U10378 (N_10378,N_10184,N_10038);
nand U10379 (N_10379,N_10212,N_10060);
and U10380 (N_10380,N_10209,N_10041);
and U10381 (N_10381,N_10068,N_10211);
xnor U10382 (N_10382,N_10057,N_10147);
and U10383 (N_10383,N_10088,N_10048);
nor U10384 (N_10384,N_10156,N_10136);
nor U10385 (N_10385,N_10185,N_10234);
or U10386 (N_10386,N_10017,N_10072);
nand U10387 (N_10387,N_10065,N_10150);
or U10388 (N_10388,N_10146,N_10025);
and U10389 (N_10389,N_10195,N_10208);
xnor U10390 (N_10390,N_10027,N_10187);
or U10391 (N_10391,N_10034,N_10194);
nand U10392 (N_10392,N_10189,N_10029);
xnor U10393 (N_10393,N_10156,N_10238);
or U10394 (N_10394,N_10031,N_10135);
nor U10395 (N_10395,N_10153,N_10230);
xnor U10396 (N_10396,N_10054,N_10177);
xnor U10397 (N_10397,N_10231,N_10139);
xnor U10398 (N_10398,N_10016,N_10086);
nand U10399 (N_10399,N_10059,N_10007);
and U10400 (N_10400,N_10235,N_10048);
or U10401 (N_10401,N_10103,N_10009);
nor U10402 (N_10402,N_10023,N_10212);
and U10403 (N_10403,N_10238,N_10150);
nand U10404 (N_10404,N_10133,N_10080);
nand U10405 (N_10405,N_10113,N_10151);
nor U10406 (N_10406,N_10169,N_10199);
nor U10407 (N_10407,N_10015,N_10170);
and U10408 (N_10408,N_10165,N_10186);
nor U10409 (N_10409,N_10122,N_10196);
and U10410 (N_10410,N_10107,N_10017);
nand U10411 (N_10411,N_10210,N_10133);
nand U10412 (N_10412,N_10024,N_10036);
xor U10413 (N_10413,N_10175,N_10042);
nand U10414 (N_10414,N_10105,N_10093);
nor U10415 (N_10415,N_10092,N_10148);
nor U10416 (N_10416,N_10081,N_10223);
or U10417 (N_10417,N_10152,N_10131);
xnor U10418 (N_10418,N_10233,N_10176);
or U10419 (N_10419,N_10211,N_10034);
and U10420 (N_10420,N_10079,N_10202);
xor U10421 (N_10421,N_10174,N_10236);
and U10422 (N_10422,N_10108,N_10096);
and U10423 (N_10423,N_10067,N_10116);
nand U10424 (N_10424,N_10234,N_10106);
and U10425 (N_10425,N_10214,N_10040);
nand U10426 (N_10426,N_10181,N_10064);
nand U10427 (N_10427,N_10119,N_10040);
nor U10428 (N_10428,N_10058,N_10159);
nand U10429 (N_10429,N_10229,N_10208);
or U10430 (N_10430,N_10032,N_10065);
nand U10431 (N_10431,N_10070,N_10170);
or U10432 (N_10432,N_10091,N_10042);
xor U10433 (N_10433,N_10009,N_10180);
nor U10434 (N_10434,N_10130,N_10200);
and U10435 (N_10435,N_10224,N_10162);
nor U10436 (N_10436,N_10150,N_10166);
nand U10437 (N_10437,N_10081,N_10076);
or U10438 (N_10438,N_10197,N_10133);
nand U10439 (N_10439,N_10222,N_10241);
nand U10440 (N_10440,N_10235,N_10004);
xnor U10441 (N_10441,N_10235,N_10173);
xnor U10442 (N_10442,N_10071,N_10138);
or U10443 (N_10443,N_10136,N_10203);
xnor U10444 (N_10444,N_10207,N_10032);
xor U10445 (N_10445,N_10081,N_10003);
xnor U10446 (N_10446,N_10097,N_10175);
and U10447 (N_10447,N_10068,N_10105);
xor U10448 (N_10448,N_10066,N_10202);
nand U10449 (N_10449,N_10058,N_10151);
and U10450 (N_10450,N_10221,N_10090);
nand U10451 (N_10451,N_10117,N_10080);
or U10452 (N_10452,N_10235,N_10247);
nor U10453 (N_10453,N_10054,N_10026);
xor U10454 (N_10454,N_10057,N_10228);
nor U10455 (N_10455,N_10113,N_10203);
nor U10456 (N_10456,N_10081,N_10227);
and U10457 (N_10457,N_10153,N_10203);
or U10458 (N_10458,N_10119,N_10220);
and U10459 (N_10459,N_10182,N_10101);
and U10460 (N_10460,N_10012,N_10174);
or U10461 (N_10461,N_10163,N_10195);
or U10462 (N_10462,N_10119,N_10128);
xnor U10463 (N_10463,N_10180,N_10195);
and U10464 (N_10464,N_10107,N_10060);
nand U10465 (N_10465,N_10043,N_10021);
nor U10466 (N_10466,N_10046,N_10096);
or U10467 (N_10467,N_10124,N_10207);
nor U10468 (N_10468,N_10137,N_10099);
nand U10469 (N_10469,N_10171,N_10228);
xnor U10470 (N_10470,N_10086,N_10004);
or U10471 (N_10471,N_10141,N_10159);
xnor U10472 (N_10472,N_10020,N_10153);
nand U10473 (N_10473,N_10202,N_10113);
nand U10474 (N_10474,N_10010,N_10038);
nand U10475 (N_10475,N_10137,N_10032);
and U10476 (N_10476,N_10024,N_10053);
or U10477 (N_10477,N_10112,N_10036);
nor U10478 (N_10478,N_10212,N_10012);
and U10479 (N_10479,N_10184,N_10054);
or U10480 (N_10480,N_10026,N_10005);
or U10481 (N_10481,N_10064,N_10146);
and U10482 (N_10482,N_10139,N_10085);
nand U10483 (N_10483,N_10025,N_10110);
nand U10484 (N_10484,N_10086,N_10160);
or U10485 (N_10485,N_10201,N_10187);
nor U10486 (N_10486,N_10143,N_10209);
or U10487 (N_10487,N_10179,N_10214);
xnor U10488 (N_10488,N_10148,N_10228);
and U10489 (N_10489,N_10090,N_10068);
xor U10490 (N_10490,N_10066,N_10022);
xor U10491 (N_10491,N_10242,N_10196);
or U10492 (N_10492,N_10097,N_10062);
and U10493 (N_10493,N_10098,N_10162);
xnor U10494 (N_10494,N_10178,N_10017);
nand U10495 (N_10495,N_10056,N_10114);
and U10496 (N_10496,N_10159,N_10148);
xor U10497 (N_10497,N_10121,N_10215);
xnor U10498 (N_10498,N_10042,N_10040);
or U10499 (N_10499,N_10162,N_10017);
nand U10500 (N_10500,N_10365,N_10415);
nand U10501 (N_10501,N_10437,N_10447);
or U10502 (N_10502,N_10299,N_10474);
xnor U10503 (N_10503,N_10412,N_10488);
xor U10504 (N_10504,N_10453,N_10306);
xor U10505 (N_10505,N_10411,N_10404);
nor U10506 (N_10506,N_10267,N_10392);
xor U10507 (N_10507,N_10426,N_10377);
xor U10508 (N_10508,N_10280,N_10398);
nor U10509 (N_10509,N_10304,N_10316);
xnor U10510 (N_10510,N_10328,N_10250);
nor U10511 (N_10511,N_10309,N_10346);
or U10512 (N_10512,N_10472,N_10445);
and U10513 (N_10513,N_10349,N_10450);
xnor U10514 (N_10514,N_10266,N_10329);
or U10515 (N_10515,N_10489,N_10448);
nor U10516 (N_10516,N_10492,N_10458);
nor U10517 (N_10517,N_10495,N_10423);
or U10518 (N_10518,N_10491,N_10345);
nor U10519 (N_10519,N_10255,N_10397);
or U10520 (N_10520,N_10473,N_10406);
nor U10521 (N_10521,N_10361,N_10278);
and U10522 (N_10522,N_10360,N_10371);
nand U10523 (N_10523,N_10457,N_10442);
nand U10524 (N_10524,N_10425,N_10486);
nand U10525 (N_10525,N_10376,N_10369);
and U10526 (N_10526,N_10494,N_10296);
and U10527 (N_10527,N_10362,N_10387);
and U10528 (N_10528,N_10318,N_10413);
or U10529 (N_10529,N_10339,N_10419);
xnor U10530 (N_10530,N_10301,N_10321);
or U10531 (N_10531,N_10275,N_10300);
xnor U10532 (N_10532,N_10394,N_10270);
and U10533 (N_10533,N_10452,N_10320);
nand U10534 (N_10534,N_10253,N_10390);
xnor U10535 (N_10535,N_10348,N_10324);
nand U10536 (N_10536,N_10310,N_10281);
or U10537 (N_10537,N_10483,N_10338);
and U10538 (N_10538,N_10443,N_10436);
xor U10539 (N_10539,N_10433,N_10340);
xnor U10540 (N_10540,N_10432,N_10468);
and U10541 (N_10541,N_10277,N_10272);
nand U10542 (N_10542,N_10289,N_10359);
nand U10543 (N_10543,N_10375,N_10493);
nor U10544 (N_10544,N_10414,N_10265);
xor U10545 (N_10545,N_10370,N_10481);
and U10546 (N_10546,N_10342,N_10274);
or U10547 (N_10547,N_10259,N_10416);
or U10548 (N_10548,N_10459,N_10322);
nand U10549 (N_10549,N_10422,N_10288);
nor U10550 (N_10550,N_10262,N_10254);
xor U10551 (N_10551,N_10395,N_10367);
xnor U10552 (N_10552,N_10388,N_10302);
or U10553 (N_10553,N_10334,N_10393);
nor U10554 (N_10554,N_10373,N_10283);
and U10555 (N_10555,N_10383,N_10444);
and U10556 (N_10556,N_10421,N_10261);
xor U10557 (N_10557,N_10396,N_10356);
and U10558 (N_10558,N_10344,N_10276);
nand U10559 (N_10559,N_10385,N_10333);
nand U10560 (N_10560,N_10456,N_10308);
or U10561 (N_10561,N_10279,N_10497);
xnor U10562 (N_10562,N_10311,N_10382);
nor U10563 (N_10563,N_10460,N_10363);
nor U10564 (N_10564,N_10366,N_10330);
xnor U10565 (N_10565,N_10462,N_10409);
xor U10566 (N_10566,N_10418,N_10268);
nand U10567 (N_10567,N_10455,N_10490);
xnor U10568 (N_10568,N_10285,N_10297);
xor U10569 (N_10569,N_10314,N_10401);
nand U10570 (N_10570,N_10343,N_10487);
and U10571 (N_10571,N_10358,N_10368);
xor U10572 (N_10572,N_10496,N_10251);
nor U10573 (N_10573,N_10391,N_10446);
and U10574 (N_10574,N_10260,N_10323);
nor U10575 (N_10575,N_10464,N_10400);
xor U10576 (N_10576,N_10417,N_10264);
or U10577 (N_10577,N_10410,N_10440);
or U10578 (N_10578,N_10466,N_10303);
nand U10579 (N_10579,N_10485,N_10336);
and U10580 (N_10580,N_10461,N_10357);
xor U10581 (N_10581,N_10313,N_10307);
or U10582 (N_10582,N_10364,N_10386);
nor U10583 (N_10583,N_10498,N_10479);
and U10584 (N_10584,N_10287,N_10438);
nor U10585 (N_10585,N_10429,N_10298);
nand U10586 (N_10586,N_10273,N_10290);
and U10587 (N_10587,N_10355,N_10374);
nand U10588 (N_10588,N_10331,N_10469);
nor U10589 (N_10589,N_10332,N_10312);
and U10590 (N_10590,N_10381,N_10431);
nand U10591 (N_10591,N_10449,N_10263);
nor U10592 (N_10592,N_10292,N_10325);
xor U10593 (N_10593,N_10352,N_10317);
and U10594 (N_10594,N_10405,N_10258);
and U10595 (N_10595,N_10293,N_10454);
and U10596 (N_10596,N_10480,N_10294);
or U10597 (N_10597,N_10257,N_10428);
nor U10598 (N_10598,N_10402,N_10271);
or U10599 (N_10599,N_10284,N_10335);
xor U10600 (N_10600,N_10439,N_10477);
or U10601 (N_10601,N_10291,N_10403);
xnor U10602 (N_10602,N_10399,N_10476);
xor U10603 (N_10603,N_10389,N_10471);
nand U10604 (N_10604,N_10347,N_10380);
nand U10605 (N_10605,N_10475,N_10315);
xnor U10606 (N_10606,N_10484,N_10408);
nor U10607 (N_10607,N_10282,N_10435);
xor U10608 (N_10608,N_10420,N_10465);
xor U10609 (N_10609,N_10482,N_10354);
xnor U10610 (N_10610,N_10326,N_10378);
nor U10611 (N_10611,N_10463,N_10319);
and U10612 (N_10612,N_10286,N_10427);
and U10613 (N_10613,N_10499,N_10379);
and U10614 (N_10614,N_10256,N_10353);
nor U10615 (N_10615,N_10451,N_10351);
nand U10616 (N_10616,N_10372,N_10350);
or U10617 (N_10617,N_10407,N_10341);
or U10618 (N_10618,N_10478,N_10252);
xor U10619 (N_10619,N_10295,N_10434);
nand U10620 (N_10620,N_10467,N_10305);
or U10621 (N_10621,N_10430,N_10441);
nand U10622 (N_10622,N_10327,N_10470);
or U10623 (N_10623,N_10269,N_10424);
and U10624 (N_10624,N_10384,N_10337);
nand U10625 (N_10625,N_10434,N_10484);
nand U10626 (N_10626,N_10336,N_10493);
nand U10627 (N_10627,N_10274,N_10476);
nor U10628 (N_10628,N_10432,N_10270);
nand U10629 (N_10629,N_10287,N_10327);
or U10630 (N_10630,N_10415,N_10466);
xor U10631 (N_10631,N_10312,N_10339);
nor U10632 (N_10632,N_10364,N_10340);
xnor U10633 (N_10633,N_10377,N_10423);
nor U10634 (N_10634,N_10357,N_10293);
or U10635 (N_10635,N_10423,N_10372);
xnor U10636 (N_10636,N_10404,N_10456);
and U10637 (N_10637,N_10402,N_10426);
and U10638 (N_10638,N_10348,N_10476);
and U10639 (N_10639,N_10427,N_10360);
nand U10640 (N_10640,N_10482,N_10387);
xnor U10641 (N_10641,N_10386,N_10255);
or U10642 (N_10642,N_10414,N_10447);
nand U10643 (N_10643,N_10412,N_10447);
xor U10644 (N_10644,N_10452,N_10281);
xor U10645 (N_10645,N_10476,N_10434);
and U10646 (N_10646,N_10380,N_10255);
xor U10647 (N_10647,N_10257,N_10370);
nand U10648 (N_10648,N_10467,N_10375);
nor U10649 (N_10649,N_10262,N_10343);
xor U10650 (N_10650,N_10328,N_10474);
xor U10651 (N_10651,N_10325,N_10290);
nand U10652 (N_10652,N_10305,N_10309);
xor U10653 (N_10653,N_10499,N_10334);
and U10654 (N_10654,N_10314,N_10265);
nor U10655 (N_10655,N_10466,N_10423);
xor U10656 (N_10656,N_10328,N_10371);
nand U10657 (N_10657,N_10344,N_10285);
xor U10658 (N_10658,N_10279,N_10357);
nand U10659 (N_10659,N_10422,N_10375);
xnor U10660 (N_10660,N_10470,N_10264);
or U10661 (N_10661,N_10344,N_10458);
nor U10662 (N_10662,N_10352,N_10276);
xor U10663 (N_10663,N_10420,N_10336);
or U10664 (N_10664,N_10427,N_10317);
nor U10665 (N_10665,N_10409,N_10393);
and U10666 (N_10666,N_10296,N_10331);
nor U10667 (N_10667,N_10278,N_10453);
nand U10668 (N_10668,N_10388,N_10456);
nand U10669 (N_10669,N_10278,N_10443);
and U10670 (N_10670,N_10428,N_10430);
or U10671 (N_10671,N_10483,N_10355);
nand U10672 (N_10672,N_10358,N_10445);
xnor U10673 (N_10673,N_10348,N_10384);
nand U10674 (N_10674,N_10416,N_10497);
nand U10675 (N_10675,N_10270,N_10287);
or U10676 (N_10676,N_10289,N_10346);
and U10677 (N_10677,N_10282,N_10341);
nor U10678 (N_10678,N_10483,N_10417);
nand U10679 (N_10679,N_10252,N_10400);
xnor U10680 (N_10680,N_10416,N_10362);
nor U10681 (N_10681,N_10278,N_10486);
nor U10682 (N_10682,N_10445,N_10422);
nand U10683 (N_10683,N_10266,N_10372);
and U10684 (N_10684,N_10415,N_10445);
nand U10685 (N_10685,N_10484,N_10299);
nand U10686 (N_10686,N_10342,N_10281);
and U10687 (N_10687,N_10367,N_10254);
xnor U10688 (N_10688,N_10381,N_10463);
xnor U10689 (N_10689,N_10268,N_10338);
nor U10690 (N_10690,N_10459,N_10440);
and U10691 (N_10691,N_10311,N_10357);
xnor U10692 (N_10692,N_10327,N_10473);
nand U10693 (N_10693,N_10487,N_10311);
or U10694 (N_10694,N_10454,N_10419);
and U10695 (N_10695,N_10459,N_10347);
xnor U10696 (N_10696,N_10465,N_10409);
xor U10697 (N_10697,N_10283,N_10277);
xnor U10698 (N_10698,N_10421,N_10349);
nor U10699 (N_10699,N_10379,N_10469);
xor U10700 (N_10700,N_10397,N_10388);
or U10701 (N_10701,N_10377,N_10325);
and U10702 (N_10702,N_10485,N_10453);
and U10703 (N_10703,N_10342,N_10464);
nor U10704 (N_10704,N_10401,N_10385);
nand U10705 (N_10705,N_10340,N_10253);
or U10706 (N_10706,N_10474,N_10379);
xor U10707 (N_10707,N_10439,N_10290);
nand U10708 (N_10708,N_10275,N_10260);
nand U10709 (N_10709,N_10322,N_10390);
or U10710 (N_10710,N_10476,N_10346);
nand U10711 (N_10711,N_10466,N_10460);
or U10712 (N_10712,N_10413,N_10390);
and U10713 (N_10713,N_10289,N_10433);
and U10714 (N_10714,N_10261,N_10266);
nand U10715 (N_10715,N_10465,N_10391);
nor U10716 (N_10716,N_10325,N_10415);
xnor U10717 (N_10717,N_10331,N_10309);
nor U10718 (N_10718,N_10276,N_10462);
and U10719 (N_10719,N_10309,N_10449);
and U10720 (N_10720,N_10294,N_10253);
nand U10721 (N_10721,N_10300,N_10357);
xnor U10722 (N_10722,N_10455,N_10454);
nand U10723 (N_10723,N_10392,N_10335);
or U10724 (N_10724,N_10488,N_10438);
nor U10725 (N_10725,N_10446,N_10330);
nor U10726 (N_10726,N_10299,N_10349);
or U10727 (N_10727,N_10294,N_10448);
nand U10728 (N_10728,N_10427,N_10302);
xnor U10729 (N_10729,N_10482,N_10270);
and U10730 (N_10730,N_10312,N_10495);
nand U10731 (N_10731,N_10393,N_10437);
nor U10732 (N_10732,N_10457,N_10467);
xnor U10733 (N_10733,N_10357,N_10342);
or U10734 (N_10734,N_10395,N_10284);
nand U10735 (N_10735,N_10485,N_10302);
and U10736 (N_10736,N_10422,N_10347);
xor U10737 (N_10737,N_10497,N_10415);
and U10738 (N_10738,N_10479,N_10252);
or U10739 (N_10739,N_10336,N_10334);
and U10740 (N_10740,N_10374,N_10283);
nand U10741 (N_10741,N_10378,N_10412);
nand U10742 (N_10742,N_10391,N_10382);
and U10743 (N_10743,N_10414,N_10475);
nand U10744 (N_10744,N_10279,N_10371);
nor U10745 (N_10745,N_10418,N_10459);
and U10746 (N_10746,N_10467,N_10324);
xor U10747 (N_10747,N_10304,N_10411);
or U10748 (N_10748,N_10279,N_10338);
or U10749 (N_10749,N_10385,N_10463);
or U10750 (N_10750,N_10584,N_10577);
xnor U10751 (N_10751,N_10725,N_10718);
or U10752 (N_10752,N_10695,N_10533);
and U10753 (N_10753,N_10563,N_10682);
and U10754 (N_10754,N_10711,N_10660);
nand U10755 (N_10755,N_10747,N_10652);
nand U10756 (N_10756,N_10578,N_10740);
and U10757 (N_10757,N_10648,N_10672);
nand U10758 (N_10758,N_10524,N_10614);
and U10759 (N_10759,N_10576,N_10624);
and U10760 (N_10760,N_10516,N_10690);
or U10761 (N_10761,N_10523,N_10553);
and U10762 (N_10762,N_10592,N_10691);
or U10763 (N_10763,N_10650,N_10673);
nand U10764 (N_10764,N_10509,N_10728);
xnor U10765 (N_10765,N_10591,N_10529);
nor U10766 (N_10766,N_10595,N_10670);
nand U10767 (N_10767,N_10735,N_10649);
nor U10768 (N_10768,N_10579,N_10598);
xor U10769 (N_10769,N_10603,N_10580);
nand U10770 (N_10770,N_10638,N_10558);
nand U10771 (N_10771,N_10730,N_10743);
and U10772 (N_10772,N_10572,N_10643);
nor U10773 (N_10773,N_10560,N_10583);
xnor U10774 (N_10774,N_10688,N_10681);
nor U10775 (N_10775,N_10678,N_10706);
or U10776 (N_10776,N_10604,N_10539);
nor U10777 (N_10777,N_10525,N_10664);
xor U10778 (N_10778,N_10582,N_10731);
or U10779 (N_10779,N_10641,N_10712);
nor U10780 (N_10780,N_10587,N_10645);
xor U10781 (N_10781,N_10503,N_10552);
nor U10782 (N_10782,N_10676,N_10601);
nand U10783 (N_10783,N_10703,N_10658);
xnor U10784 (N_10784,N_10659,N_10713);
or U10785 (N_10785,N_10547,N_10651);
nor U10786 (N_10786,N_10510,N_10683);
xor U10787 (N_10787,N_10543,N_10520);
nor U10788 (N_10788,N_10722,N_10668);
or U10789 (N_10789,N_10692,N_10541);
nand U10790 (N_10790,N_10554,N_10551);
nor U10791 (N_10791,N_10530,N_10654);
and U10792 (N_10792,N_10644,N_10517);
nor U10793 (N_10793,N_10732,N_10693);
nor U10794 (N_10794,N_10656,N_10586);
xnor U10795 (N_10795,N_10617,N_10736);
xor U10796 (N_10796,N_10506,N_10663);
and U10797 (N_10797,N_10636,N_10540);
or U10798 (N_10798,N_10669,N_10561);
nand U10799 (N_10799,N_10719,N_10502);
or U10800 (N_10800,N_10628,N_10640);
nor U10801 (N_10801,N_10720,N_10627);
and U10802 (N_10802,N_10737,N_10613);
and U10803 (N_10803,N_10568,N_10610);
or U10804 (N_10804,N_10618,N_10570);
and U10805 (N_10805,N_10635,N_10723);
and U10806 (N_10806,N_10704,N_10705);
nand U10807 (N_10807,N_10620,N_10549);
xnor U10808 (N_10808,N_10702,N_10744);
or U10809 (N_10809,N_10653,N_10504);
and U10810 (N_10810,N_10545,N_10684);
or U10811 (N_10811,N_10528,N_10581);
nand U10812 (N_10812,N_10689,N_10544);
xor U10813 (N_10813,N_10536,N_10514);
and U10814 (N_10814,N_10697,N_10671);
nor U10815 (N_10815,N_10675,N_10694);
or U10816 (N_10816,N_10745,N_10527);
nor U10817 (N_10817,N_10749,N_10526);
and U10818 (N_10818,N_10622,N_10519);
nand U10819 (N_10819,N_10642,N_10521);
nor U10820 (N_10820,N_10593,N_10607);
nor U10821 (N_10821,N_10639,N_10542);
xor U10822 (N_10822,N_10512,N_10585);
or U10823 (N_10823,N_10726,N_10507);
xnor U10824 (N_10824,N_10707,N_10500);
xor U10825 (N_10825,N_10559,N_10655);
and U10826 (N_10826,N_10714,N_10634);
and U10827 (N_10827,N_10715,N_10606);
nor U10828 (N_10828,N_10727,N_10569);
or U10829 (N_10829,N_10602,N_10698);
and U10830 (N_10830,N_10710,N_10615);
or U10831 (N_10831,N_10612,N_10665);
nor U10832 (N_10832,N_10637,N_10616);
xor U10833 (N_10833,N_10729,N_10531);
or U10834 (N_10834,N_10511,N_10501);
nand U10835 (N_10835,N_10629,N_10708);
xnor U10836 (N_10836,N_10573,N_10619);
nor U10837 (N_10837,N_10522,N_10608);
nand U10838 (N_10838,N_10657,N_10538);
xnor U10839 (N_10839,N_10716,N_10696);
xnor U10840 (N_10840,N_10646,N_10661);
nand U10841 (N_10841,N_10574,N_10590);
or U10842 (N_10842,N_10537,N_10700);
xnor U10843 (N_10843,N_10515,N_10550);
nand U10844 (N_10844,N_10633,N_10662);
nor U10845 (N_10845,N_10566,N_10605);
xnor U10846 (N_10846,N_10596,N_10738);
nor U10847 (N_10847,N_10709,N_10599);
xnor U10848 (N_10848,N_10600,N_10609);
xor U10849 (N_10849,N_10724,N_10647);
and U10850 (N_10850,N_10734,N_10679);
nor U10851 (N_10851,N_10748,N_10631);
nor U10852 (N_10852,N_10623,N_10666);
nor U10853 (N_10853,N_10733,N_10701);
nand U10854 (N_10854,N_10546,N_10741);
nor U10855 (N_10855,N_10532,N_10611);
or U10856 (N_10856,N_10567,N_10564);
nor U10857 (N_10857,N_10575,N_10508);
and U10858 (N_10858,N_10626,N_10680);
or U10859 (N_10859,N_10687,N_10667);
xor U10860 (N_10860,N_10571,N_10621);
and U10861 (N_10861,N_10505,N_10746);
nor U10862 (N_10862,N_10548,N_10555);
or U10863 (N_10863,N_10742,N_10589);
nor U10864 (N_10864,N_10534,N_10565);
xnor U10865 (N_10865,N_10674,N_10677);
and U10866 (N_10866,N_10739,N_10562);
xor U10867 (N_10867,N_10625,N_10588);
nor U10868 (N_10868,N_10518,N_10513);
nor U10869 (N_10869,N_10557,N_10597);
nand U10870 (N_10870,N_10630,N_10594);
nor U10871 (N_10871,N_10556,N_10717);
and U10872 (N_10872,N_10535,N_10699);
nand U10873 (N_10873,N_10721,N_10685);
nor U10874 (N_10874,N_10686,N_10632);
xor U10875 (N_10875,N_10745,N_10744);
nand U10876 (N_10876,N_10575,N_10522);
and U10877 (N_10877,N_10696,N_10557);
xnor U10878 (N_10878,N_10694,N_10742);
xor U10879 (N_10879,N_10560,N_10676);
and U10880 (N_10880,N_10539,N_10524);
xnor U10881 (N_10881,N_10514,N_10653);
nand U10882 (N_10882,N_10594,N_10615);
xnor U10883 (N_10883,N_10694,N_10673);
or U10884 (N_10884,N_10722,N_10667);
and U10885 (N_10885,N_10664,N_10679);
nor U10886 (N_10886,N_10662,N_10690);
xor U10887 (N_10887,N_10653,N_10626);
and U10888 (N_10888,N_10642,N_10512);
or U10889 (N_10889,N_10550,N_10686);
or U10890 (N_10890,N_10565,N_10561);
nand U10891 (N_10891,N_10630,N_10607);
and U10892 (N_10892,N_10744,N_10579);
nand U10893 (N_10893,N_10738,N_10619);
nor U10894 (N_10894,N_10601,N_10693);
nor U10895 (N_10895,N_10687,N_10502);
and U10896 (N_10896,N_10694,N_10617);
and U10897 (N_10897,N_10741,N_10540);
nor U10898 (N_10898,N_10521,N_10694);
nor U10899 (N_10899,N_10727,N_10665);
and U10900 (N_10900,N_10565,N_10720);
and U10901 (N_10901,N_10701,N_10512);
xnor U10902 (N_10902,N_10726,N_10567);
or U10903 (N_10903,N_10596,N_10549);
nor U10904 (N_10904,N_10635,N_10537);
or U10905 (N_10905,N_10669,N_10677);
or U10906 (N_10906,N_10699,N_10646);
and U10907 (N_10907,N_10665,N_10569);
nor U10908 (N_10908,N_10712,N_10643);
xor U10909 (N_10909,N_10698,N_10504);
nor U10910 (N_10910,N_10567,N_10536);
nor U10911 (N_10911,N_10744,N_10633);
xnor U10912 (N_10912,N_10733,N_10707);
and U10913 (N_10913,N_10712,N_10576);
and U10914 (N_10914,N_10571,N_10601);
or U10915 (N_10915,N_10630,N_10591);
xnor U10916 (N_10916,N_10637,N_10609);
nor U10917 (N_10917,N_10602,N_10574);
nand U10918 (N_10918,N_10549,N_10588);
or U10919 (N_10919,N_10655,N_10735);
nor U10920 (N_10920,N_10705,N_10691);
nor U10921 (N_10921,N_10736,N_10603);
xor U10922 (N_10922,N_10542,N_10728);
and U10923 (N_10923,N_10636,N_10677);
or U10924 (N_10924,N_10631,N_10671);
and U10925 (N_10925,N_10524,N_10535);
nand U10926 (N_10926,N_10626,N_10643);
nor U10927 (N_10927,N_10612,N_10502);
nor U10928 (N_10928,N_10718,N_10533);
nand U10929 (N_10929,N_10656,N_10608);
or U10930 (N_10930,N_10534,N_10749);
or U10931 (N_10931,N_10594,N_10721);
or U10932 (N_10932,N_10507,N_10737);
and U10933 (N_10933,N_10541,N_10584);
and U10934 (N_10934,N_10631,N_10507);
nand U10935 (N_10935,N_10584,N_10546);
nand U10936 (N_10936,N_10506,N_10548);
or U10937 (N_10937,N_10637,N_10578);
nand U10938 (N_10938,N_10542,N_10657);
nor U10939 (N_10939,N_10698,N_10722);
nor U10940 (N_10940,N_10661,N_10525);
nand U10941 (N_10941,N_10579,N_10505);
xor U10942 (N_10942,N_10536,N_10663);
nor U10943 (N_10943,N_10733,N_10621);
or U10944 (N_10944,N_10620,N_10734);
and U10945 (N_10945,N_10590,N_10652);
nand U10946 (N_10946,N_10536,N_10676);
nor U10947 (N_10947,N_10698,N_10692);
nand U10948 (N_10948,N_10535,N_10715);
nor U10949 (N_10949,N_10661,N_10609);
xnor U10950 (N_10950,N_10605,N_10542);
nand U10951 (N_10951,N_10644,N_10728);
nand U10952 (N_10952,N_10707,N_10699);
nand U10953 (N_10953,N_10535,N_10542);
and U10954 (N_10954,N_10549,N_10574);
and U10955 (N_10955,N_10635,N_10726);
nand U10956 (N_10956,N_10744,N_10515);
xor U10957 (N_10957,N_10647,N_10690);
and U10958 (N_10958,N_10563,N_10704);
nor U10959 (N_10959,N_10519,N_10643);
or U10960 (N_10960,N_10579,N_10643);
or U10961 (N_10961,N_10658,N_10585);
and U10962 (N_10962,N_10685,N_10693);
nor U10963 (N_10963,N_10546,N_10705);
and U10964 (N_10964,N_10577,N_10711);
and U10965 (N_10965,N_10734,N_10538);
nor U10966 (N_10966,N_10689,N_10633);
xnor U10967 (N_10967,N_10672,N_10697);
xor U10968 (N_10968,N_10560,N_10651);
nand U10969 (N_10969,N_10730,N_10562);
xnor U10970 (N_10970,N_10686,N_10609);
nand U10971 (N_10971,N_10653,N_10516);
and U10972 (N_10972,N_10521,N_10503);
or U10973 (N_10973,N_10639,N_10708);
and U10974 (N_10974,N_10745,N_10703);
or U10975 (N_10975,N_10587,N_10506);
nand U10976 (N_10976,N_10645,N_10546);
nor U10977 (N_10977,N_10732,N_10694);
or U10978 (N_10978,N_10718,N_10667);
nor U10979 (N_10979,N_10591,N_10654);
nand U10980 (N_10980,N_10525,N_10615);
or U10981 (N_10981,N_10674,N_10690);
xnor U10982 (N_10982,N_10528,N_10613);
and U10983 (N_10983,N_10579,N_10708);
and U10984 (N_10984,N_10615,N_10630);
xnor U10985 (N_10985,N_10565,N_10613);
nand U10986 (N_10986,N_10690,N_10644);
nor U10987 (N_10987,N_10645,N_10726);
xor U10988 (N_10988,N_10601,N_10606);
nor U10989 (N_10989,N_10669,N_10666);
and U10990 (N_10990,N_10573,N_10533);
xor U10991 (N_10991,N_10516,N_10584);
xor U10992 (N_10992,N_10714,N_10517);
or U10993 (N_10993,N_10545,N_10530);
and U10994 (N_10994,N_10701,N_10599);
and U10995 (N_10995,N_10665,N_10552);
nor U10996 (N_10996,N_10515,N_10597);
and U10997 (N_10997,N_10681,N_10555);
xnor U10998 (N_10998,N_10524,N_10627);
nand U10999 (N_10999,N_10521,N_10522);
nor U11000 (N_11000,N_10996,N_10992);
or U11001 (N_11001,N_10813,N_10897);
and U11002 (N_11002,N_10987,N_10852);
nand U11003 (N_11003,N_10957,N_10836);
or U11004 (N_11004,N_10910,N_10796);
and U11005 (N_11005,N_10809,N_10899);
and U11006 (N_11006,N_10798,N_10985);
nor U11007 (N_11007,N_10898,N_10845);
or U11008 (N_11008,N_10860,N_10922);
nor U11009 (N_11009,N_10909,N_10811);
xor U11010 (N_11010,N_10810,N_10993);
nor U11011 (N_11011,N_10953,N_10853);
or U11012 (N_11012,N_10858,N_10850);
or U11013 (N_11013,N_10812,N_10808);
nand U11014 (N_11014,N_10893,N_10924);
and U11015 (N_11015,N_10989,N_10762);
or U11016 (N_11016,N_10849,N_10753);
and U11017 (N_11017,N_10838,N_10966);
or U11018 (N_11018,N_10948,N_10946);
and U11019 (N_11019,N_10821,N_10815);
and U11020 (N_11020,N_10831,N_10759);
and U11021 (N_11021,N_10889,N_10965);
or U11022 (N_11022,N_10926,N_10894);
or U11023 (N_11023,N_10886,N_10940);
and U11024 (N_11024,N_10766,N_10859);
or U11025 (N_11025,N_10915,N_10997);
or U11026 (N_11026,N_10869,N_10863);
or U11027 (N_11027,N_10846,N_10844);
and U11028 (N_11028,N_10829,N_10760);
nand U11029 (N_11029,N_10991,N_10871);
and U11030 (N_11030,N_10961,N_10925);
nor U11031 (N_11031,N_10941,N_10960);
nor U11032 (N_11032,N_10947,N_10873);
and U11033 (N_11033,N_10778,N_10783);
xnor U11034 (N_11034,N_10972,N_10772);
nor U11035 (N_11035,N_10819,N_10883);
and U11036 (N_11036,N_10968,N_10930);
xor U11037 (N_11037,N_10804,N_10781);
nor U11038 (N_11038,N_10773,N_10980);
nand U11039 (N_11039,N_10801,N_10867);
nor U11040 (N_11040,N_10785,N_10769);
nor U11041 (N_11041,N_10887,N_10822);
or U11042 (N_11042,N_10955,N_10788);
nor U11043 (N_11043,N_10876,N_10929);
xnor U11044 (N_11044,N_10761,N_10837);
xnor U11045 (N_11045,N_10994,N_10782);
and U11046 (N_11046,N_10750,N_10891);
and U11047 (N_11047,N_10807,N_10881);
and U11048 (N_11048,N_10979,N_10864);
xor U11049 (N_11049,N_10904,N_10885);
xor U11050 (N_11050,N_10905,N_10959);
nor U11051 (N_11051,N_10865,N_10903);
nand U11052 (N_11052,N_10916,N_10868);
or U11053 (N_11053,N_10779,N_10956);
xnor U11054 (N_11054,N_10981,N_10938);
nor U11055 (N_11055,N_10751,N_10847);
nor U11056 (N_11056,N_10877,N_10839);
nand U11057 (N_11057,N_10900,N_10862);
xor U11058 (N_11058,N_10793,N_10990);
xnor U11059 (N_11059,N_10918,N_10984);
or U11060 (N_11060,N_10952,N_10848);
xnor U11061 (N_11061,N_10817,N_10902);
nand U11062 (N_11062,N_10917,N_10874);
nand U11063 (N_11063,N_10920,N_10911);
xnor U11064 (N_11064,N_10791,N_10857);
nand U11065 (N_11065,N_10835,N_10976);
nand U11066 (N_11066,N_10971,N_10816);
and U11067 (N_11067,N_10906,N_10878);
xor U11068 (N_11068,N_10828,N_10776);
xnor U11069 (N_11069,N_10927,N_10777);
nand U11070 (N_11070,N_10832,N_10943);
nand U11071 (N_11071,N_10919,N_10901);
nand U11072 (N_11072,N_10977,N_10907);
nand U11073 (N_11073,N_10870,N_10752);
xor U11074 (N_11074,N_10842,N_10784);
nor U11075 (N_11075,N_10833,N_10823);
nor U11076 (N_11076,N_10888,N_10824);
xnor U11077 (N_11077,N_10950,N_10855);
or U11078 (N_11078,N_10795,N_10937);
nand U11079 (N_11079,N_10935,N_10914);
and U11080 (N_11080,N_10970,N_10789);
nand U11081 (N_11081,N_10806,N_10774);
nand U11082 (N_11082,N_10814,N_10963);
xnor U11083 (N_11083,N_10913,N_10792);
xnor U11084 (N_11084,N_10770,N_10999);
nand U11085 (N_11085,N_10825,N_10764);
nand U11086 (N_11086,N_10756,N_10767);
or U11087 (N_11087,N_10800,N_10958);
and U11088 (N_11088,N_10843,N_10939);
nor U11089 (N_11089,N_10763,N_10866);
xor U11090 (N_11090,N_10962,N_10802);
or U11091 (N_11091,N_10896,N_10780);
nand U11092 (N_11092,N_10969,N_10890);
nor U11093 (N_11093,N_10771,N_10973);
xor U11094 (N_11094,N_10933,N_10797);
and U11095 (N_11095,N_10978,N_10923);
xor U11096 (N_11096,N_10754,N_10936);
and U11097 (N_11097,N_10787,N_10967);
xnor U11098 (N_11098,N_10840,N_10954);
and U11099 (N_11099,N_10945,N_10934);
xor U11100 (N_11100,N_10892,N_10758);
or U11101 (N_11101,N_10820,N_10988);
nor U11102 (N_11102,N_10872,N_10786);
or U11103 (N_11103,N_10912,N_10799);
nor U11104 (N_11104,N_10964,N_10951);
xor U11105 (N_11105,N_10851,N_10982);
xor U11106 (N_11106,N_10768,N_10775);
or U11107 (N_11107,N_10931,N_10765);
or U11108 (N_11108,N_10928,N_10884);
nand U11109 (N_11109,N_10998,N_10880);
or U11110 (N_11110,N_10921,N_10879);
nand U11111 (N_11111,N_10932,N_10830);
xnor U11112 (N_11112,N_10983,N_10875);
nand U11113 (N_11113,N_10944,N_10790);
or U11114 (N_11114,N_10827,N_10854);
and U11115 (N_11115,N_10882,N_10908);
or U11116 (N_11116,N_10757,N_10986);
or U11117 (N_11117,N_10755,N_10861);
xnor U11118 (N_11118,N_10895,N_10818);
nor U11119 (N_11119,N_10834,N_10805);
nand U11120 (N_11120,N_10803,N_10975);
nor U11121 (N_11121,N_10856,N_10794);
nand U11122 (N_11122,N_10949,N_10995);
or U11123 (N_11123,N_10826,N_10841);
nor U11124 (N_11124,N_10974,N_10942);
nand U11125 (N_11125,N_10899,N_10990);
and U11126 (N_11126,N_10936,N_10918);
xor U11127 (N_11127,N_10969,N_10945);
or U11128 (N_11128,N_10786,N_10796);
nand U11129 (N_11129,N_10961,N_10972);
and U11130 (N_11130,N_10902,N_10947);
nand U11131 (N_11131,N_10785,N_10996);
or U11132 (N_11132,N_10863,N_10940);
and U11133 (N_11133,N_10876,N_10956);
and U11134 (N_11134,N_10926,N_10844);
nand U11135 (N_11135,N_10753,N_10839);
xnor U11136 (N_11136,N_10886,N_10986);
nand U11137 (N_11137,N_10840,N_10845);
and U11138 (N_11138,N_10948,N_10840);
nor U11139 (N_11139,N_10756,N_10813);
and U11140 (N_11140,N_10884,N_10864);
and U11141 (N_11141,N_10838,N_10808);
nor U11142 (N_11142,N_10753,N_10898);
xor U11143 (N_11143,N_10754,N_10839);
xor U11144 (N_11144,N_10758,N_10901);
nand U11145 (N_11145,N_10962,N_10828);
xor U11146 (N_11146,N_10941,N_10869);
nor U11147 (N_11147,N_10910,N_10986);
nand U11148 (N_11148,N_10915,N_10771);
or U11149 (N_11149,N_10910,N_10920);
and U11150 (N_11150,N_10836,N_10926);
nor U11151 (N_11151,N_10897,N_10875);
xnor U11152 (N_11152,N_10788,N_10871);
nand U11153 (N_11153,N_10962,N_10904);
and U11154 (N_11154,N_10772,N_10824);
or U11155 (N_11155,N_10861,N_10979);
xnor U11156 (N_11156,N_10919,N_10949);
nor U11157 (N_11157,N_10856,N_10845);
or U11158 (N_11158,N_10914,N_10962);
nand U11159 (N_11159,N_10968,N_10891);
nor U11160 (N_11160,N_10884,N_10926);
and U11161 (N_11161,N_10757,N_10959);
nor U11162 (N_11162,N_10769,N_10786);
and U11163 (N_11163,N_10972,N_10982);
or U11164 (N_11164,N_10853,N_10971);
or U11165 (N_11165,N_10973,N_10791);
xnor U11166 (N_11166,N_10755,N_10941);
nor U11167 (N_11167,N_10853,N_10919);
xor U11168 (N_11168,N_10901,N_10783);
nor U11169 (N_11169,N_10900,N_10769);
nand U11170 (N_11170,N_10770,N_10898);
nand U11171 (N_11171,N_10908,N_10902);
or U11172 (N_11172,N_10827,N_10998);
or U11173 (N_11173,N_10980,N_10892);
or U11174 (N_11174,N_10777,N_10955);
and U11175 (N_11175,N_10793,N_10863);
xnor U11176 (N_11176,N_10829,N_10871);
nand U11177 (N_11177,N_10814,N_10956);
or U11178 (N_11178,N_10924,N_10880);
or U11179 (N_11179,N_10843,N_10871);
nand U11180 (N_11180,N_10836,N_10788);
or U11181 (N_11181,N_10773,N_10924);
or U11182 (N_11182,N_10896,N_10794);
nor U11183 (N_11183,N_10897,N_10784);
xor U11184 (N_11184,N_10939,N_10753);
nor U11185 (N_11185,N_10778,N_10932);
and U11186 (N_11186,N_10800,N_10993);
nand U11187 (N_11187,N_10860,N_10923);
and U11188 (N_11188,N_10942,N_10766);
xor U11189 (N_11189,N_10853,N_10865);
nor U11190 (N_11190,N_10859,N_10783);
and U11191 (N_11191,N_10896,N_10754);
and U11192 (N_11192,N_10833,N_10896);
and U11193 (N_11193,N_10806,N_10879);
nor U11194 (N_11194,N_10976,N_10954);
xnor U11195 (N_11195,N_10834,N_10771);
xor U11196 (N_11196,N_10836,N_10874);
nand U11197 (N_11197,N_10804,N_10816);
nor U11198 (N_11198,N_10873,N_10936);
nand U11199 (N_11199,N_10813,N_10987);
and U11200 (N_11200,N_10972,N_10958);
and U11201 (N_11201,N_10857,N_10807);
xnor U11202 (N_11202,N_10880,N_10944);
xor U11203 (N_11203,N_10758,N_10806);
nor U11204 (N_11204,N_10858,N_10995);
or U11205 (N_11205,N_10751,N_10865);
and U11206 (N_11206,N_10798,N_10768);
or U11207 (N_11207,N_10917,N_10845);
or U11208 (N_11208,N_10818,N_10845);
nor U11209 (N_11209,N_10810,N_10950);
or U11210 (N_11210,N_10842,N_10773);
or U11211 (N_11211,N_10948,N_10870);
nor U11212 (N_11212,N_10769,N_10990);
xnor U11213 (N_11213,N_10919,N_10787);
nand U11214 (N_11214,N_10880,N_10815);
nand U11215 (N_11215,N_10892,N_10755);
xnor U11216 (N_11216,N_10908,N_10841);
or U11217 (N_11217,N_10969,N_10757);
xor U11218 (N_11218,N_10940,N_10829);
or U11219 (N_11219,N_10764,N_10959);
xor U11220 (N_11220,N_10860,N_10825);
xor U11221 (N_11221,N_10997,N_10900);
nor U11222 (N_11222,N_10859,N_10907);
or U11223 (N_11223,N_10759,N_10877);
nand U11224 (N_11224,N_10968,N_10755);
xnor U11225 (N_11225,N_10753,N_10822);
nor U11226 (N_11226,N_10750,N_10895);
nand U11227 (N_11227,N_10930,N_10878);
and U11228 (N_11228,N_10938,N_10976);
nor U11229 (N_11229,N_10862,N_10937);
and U11230 (N_11230,N_10916,N_10943);
or U11231 (N_11231,N_10915,N_10936);
nor U11232 (N_11232,N_10759,N_10942);
nand U11233 (N_11233,N_10804,N_10888);
nor U11234 (N_11234,N_10847,N_10776);
nor U11235 (N_11235,N_10995,N_10783);
or U11236 (N_11236,N_10994,N_10862);
xor U11237 (N_11237,N_10775,N_10840);
or U11238 (N_11238,N_10885,N_10918);
xnor U11239 (N_11239,N_10966,N_10897);
or U11240 (N_11240,N_10954,N_10831);
or U11241 (N_11241,N_10824,N_10805);
xor U11242 (N_11242,N_10977,N_10879);
nand U11243 (N_11243,N_10840,N_10838);
and U11244 (N_11244,N_10898,N_10936);
xnor U11245 (N_11245,N_10985,N_10772);
nor U11246 (N_11246,N_10917,N_10772);
or U11247 (N_11247,N_10881,N_10898);
and U11248 (N_11248,N_10852,N_10903);
nand U11249 (N_11249,N_10979,N_10969);
or U11250 (N_11250,N_11001,N_11125);
nor U11251 (N_11251,N_11110,N_11219);
or U11252 (N_11252,N_11004,N_11170);
nor U11253 (N_11253,N_11053,N_11213);
or U11254 (N_11254,N_11018,N_11077);
or U11255 (N_11255,N_11039,N_11247);
or U11256 (N_11256,N_11058,N_11090);
or U11257 (N_11257,N_11105,N_11181);
xnor U11258 (N_11258,N_11082,N_11231);
nor U11259 (N_11259,N_11071,N_11028);
nand U11260 (N_11260,N_11176,N_11148);
xor U11261 (N_11261,N_11098,N_11000);
or U11262 (N_11262,N_11218,N_11024);
nand U11263 (N_11263,N_11042,N_11134);
and U11264 (N_11264,N_11162,N_11052);
nor U11265 (N_11265,N_11107,N_11164);
or U11266 (N_11266,N_11179,N_11221);
or U11267 (N_11267,N_11238,N_11241);
nand U11268 (N_11268,N_11232,N_11021);
nand U11269 (N_11269,N_11009,N_11067);
and U11270 (N_11270,N_11233,N_11166);
or U11271 (N_11271,N_11045,N_11036);
and U11272 (N_11272,N_11037,N_11212);
nand U11273 (N_11273,N_11124,N_11126);
xnor U11274 (N_11274,N_11050,N_11153);
or U11275 (N_11275,N_11074,N_11234);
nor U11276 (N_11276,N_11189,N_11088);
xnor U11277 (N_11277,N_11132,N_11177);
xor U11278 (N_11278,N_11183,N_11133);
nand U11279 (N_11279,N_11111,N_11222);
and U11280 (N_11280,N_11121,N_11094);
nand U11281 (N_11281,N_11034,N_11008);
and U11282 (N_11282,N_11243,N_11122);
xor U11283 (N_11283,N_11048,N_11165);
nand U11284 (N_11284,N_11227,N_11249);
and U11285 (N_11285,N_11112,N_11178);
xnor U11286 (N_11286,N_11207,N_11242);
nor U11287 (N_11287,N_11204,N_11041);
and U11288 (N_11288,N_11031,N_11097);
nor U11289 (N_11289,N_11210,N_11230);
and U11290 (N_11290,N_11143,N_11220);
nand U11291 (N_11291,N_11186,N_11025);
and U11292 (N_11292,N_11159,N_11091);
nor U11293 (N_11293,N_11038,N_11119);
and U11294 (N_11294,N_11020,N_11196);
and U11295 (N_11295,N_11044,N_11182);
nor U11296 (N_11296,N_11073,N_11062);
nor U11297 (N_11297,N_11145,N_11078);
nor U11298 (N_11298,N_11099,N_11194);
or U11299 (N_11299,N_11137,N_11104);
or U11300 (N_11300,N_11026,N_11236);
nor U11301 (N_11301,N_11011,N_11016);
or U11302 (N_11302,N_11205,N_11055);
and U11303 (N_11303,N_11065,N_11014);
and U11304 (N_11304,N_11158,N_11072);
and U11305 (N_11305,N_11128,N_11237);
nand U11306 (N_11306,N_11129,N_11101);
or U11307 (N_11307,N_11087,N_11149);
or U11308 (N_11308,N_11108,N_11120);
and U11309 (N_11309,N_11086,N_11171);
or U11310 (N_11310,N_11115,N_11069);
nand U11311 (N_11311,N_11136,N_11084);
or U11312 (N_11312,N_11118,N_11172);
nor U11313 (N_11313,N_11224,N_11163);
nor U11314 (N_11314,N_11027,N_11175);
or U11315 (N_11315,N_11075,N_11187);
nor U11316 (N_11316,N_11089,N_11017);
xnor U11317 (N_11317,N_11198,N_11225);
xor U11318 (N_11318,N_11216,N_11195);
and U11319 (N_11319,N_11199,N_11223);
xor U11320 (N_11320,N_11206,N_11197);
xor U11321 (N_11321,N_11208,N_11096);
nand U11322 (N_11322,N_11015,N_11190);
or U11323 (N_11323,N_11217,N_11192);
and U11324 (N_11324,N_11063,N_11092);
nor U11325 (N_11325,N_11157,N_11054);
or U11326 (N_11326,N_11146,N_11180);
nor U11327 (N_11327,N_11123,N_11010);
or U11328 (N_11328,N_11167,N_11142);
and U11329 (N_11329,N_11013,N_11135);
nor U11330 (N_11330,N_11049,N_11211);
nor U11331 (N_11331,N_11066,N_11076);
nor U11332 (N_11332,N_11007,N_11023);
xor U11333 (N_11333,N_11174,N_11202);
and U11334 (N_11334,N_11151,N_11169);
nand U11335 (N_11335,N_11200,N_11060);
nand U11336 (N_11336,N_11047,N_11184);
xor U11337 (N_11337,N_11035,N_11154);
nand U11338 (N_11338,N_11117,N_11070);
xnor U11339 (N_11339,N_11019,N_11229);
or U11340 (N_11340,N_11131,N_11002);
nand U11341 (N_11341,N_11141,N_11239);
nor U11342 (N_11342,N_11064,N_11160);
and U11343 (N_11343,N_11147,N_11155);
nand U11344 (N_11344,N_11095,N_11046);
and U11345 (N_11345,N_11106,N_11057);
or U11346 (N_11346,N_11127,N_11056);
or U11347 (N_11347,N_11006,N_11085);
nand U11348 (N_11348,N_11188,N_11240);
and U11349 (N_11349,N_11244,N_11103);
or U11350 (N_11350,N_11168,N_11140);
nand U11351 (N_11351,N_11003,N_11051);
nand U11352 (N_11352,N_11139,N_11138);
or U11353 (N_11353,N_11012,N_11203);
xnor U11354 (N_11354,N_11191,N_11248);
nand U11355 (N_11355,N_11030,N_11114);
or U11356 (N_11356,N_11079,N_11152);
nor U11357 (N_11357,N_11246,N_11113);
nor U11358 (N_11358,N_11235,N_11005);
and U11359 (N_11359,N_11193,N_11059);
nor U11360 (N_11360,N_11032,N_11093);
and U11361 (N_11361,N_11116,N_11080);
nand U11362 (N_11362,N_11109,N_11185);
xor U11363 (N_11363,N_11061,N_11201);
nor U11364 (N_11364,N_11156,N_11102);
nand U11365 (N_11365,N_11215,N_11173);
or U11366 (N_11366,N_11161,N_11209);
nand U11367 (N_11367,N_11214,N_11130);
nand U11368 (N_11368,N_11040,N_11083);
nand U11369 (N_11369,N_11043,N_11029);
nand U11370 (N_11370,N_11144,N_11150);
nand U11371 (N_11371,N_11068,N_11100);
xnor U11372 (N_11372,N_11228,N_11033);
nor U11373 (N_11373,N_11245,N_11226);
and U11374 (N_11374,N_11081,N_11022);
or U11375 (N_11375,N_11047,N_11239);
and U11376 (N_11376,N_11158,N_11227);
nor U11377 (N_11377,N_11192,N_11066);
xor U11378 (N_11378,N_11003,N_11149);
and U11379 (N_11379,N_11139,N_11039);
xor U11380 (N_11380,N_11146,N_11218);
or U11381 (N_11381,N_11202,N_11186);
and U11382 (N_11382,N_11203,N_11215);
xnor U11383 (N_11383,N_11036,N_11091);
nor U11384 (N_11384,N_11044,N_11208);
nor U11385 (N_11385,N_11221,N_11110);
nand U11386 (N_11386,N_11085,N_11165);
nor U11387 (N_11387,N_11103,N_11137);
xor U11388 (N_11388,N_11067,N_11086);
nor U11389 (N_11389,N_11182,N_11047);
nor U11390 (N_11390,N_11200,N_11000);
nand U11391 (N_11391,N_11196,N_11126);
or U11392 (N_11392,N_11152,N_11073);
or U11393 (N_11393,N_11194,N_11083);
nand U11394 (N_11394,N_11203,N_11116);
nor U11395 (N_11395,N_11052,N_11227);
and U11396 (N_11396,N_11216,N_11006);
or U11397 (N_11397,N_11156,N_11231);
and U11398 (N_11398,N_11017,N_11139);
nor U11399 (N_11399,N_11158,N_11105);
nor U11400 (N_11400,N_11102,N_11135);
nor U11401 (N_11401,N_11133,N_11154);
xor U11402 (N_11402,N_11160,N_11237);
or U11403 (N_11403,N_11131,N_11150);
and U11404 (N_11404,N_11203,N_11083);
nor U11405 (N_11405,N_11100,N_11080);
xor U11406 (N_11406,N_11179,N_11126);
and U11407 (N_11407,N_11078,N_11093);
xnor U11408 (N_11408,N_11214,N_11176);
nand U11409 (N_11409,N_11239,N_11199);
xnor U11410 (N_11410,N_11189,N_11086);
nor U11411 (N_11411,N_11126,N_11021);
nand U11412 (N_11412,N_11229,N_11237);
nand U11413 (N_11413,N_11155,N_11064);
xnor U11414 (N_11414,N_11137,N_11162);
nor U11415 (N_11415,N_11198,N_11084);
and U11416 (N_11416,N_11183,N_11025);
and U11417 (N_11417,N_11167,N_11161);
xnor U11418 (N_11418,N_11219,N_11025);
nand U11419 (N_11419,N_11063,N_11238);
and U11420 (N_11420,N_11068,N_11145);
nand U11421 (N_11421,N_11231,N_11209);
nand U11422 (N_11422,N_11223,N_11085);
nand U11423 (N_11423,N_11103,N_11167);
xor U11424 (N_11424,N_11150,N_11015);
xor U11425 (N_11425,N_11065,N_11042);
nor U11426 (N_11426,N_11059,N_11204);
nand U11427 (N_11427,N_11013,N_11209);
xnor U11428 (N_11428,N_11221,N_11019);
and U11429 (N_11429,N_11010,N_11151);
xor U11430 (N_11430,N_11033,N_11051);
nor U11431 (N_11431,N_11244,N_11223);
nor U11432 (N_11432,N_11073,N_11048);
nand U11433 (N_11433,N_11116,N_11019);
nor U11434 (N_11434,N_11233,N_11154);
nand U11435 (N_11435,N_11186,N_11084);
or U11436 (N_11436,N_11147,N_11215);
and U11437 (N_11437,N_11092,N_11133);
nor U11438 (N_11438,N_11047,N_11114);
nand U11439 (N_11439,N_11021,N_11245);
or U11440 (N_11440,N_11084,N_11164);
xor U11441 (N_11441,N_11041,N_11045);
nand U11442 (N_11442,N_11178,N_11184);
xor U11443 (N_11443,N_11058,N_11070);
nand U11444 (N_11444,N_11013,N_11206);
nor U11445 (N_11445,N_11236,N_11178);
or U11446 (N_11446,N_11011,N_11170);
and U11447 (N_11447,N_11092,N_11065);
and U11448 (N_11448,N_11042,N_11120);
and U11449 (N_11449,N_11080,N_11117);
nor U11450 (N_11450,N_11232,N_11002);
or U11451 (N_11451,N_11206,N_11231);
nand U11452 (N_11452,N_11216,N_11106);
nor U11453 (N_11453,N_11176,N_11029);
nand U11454 (N_11454,N_11039,N_11119);
xnor U11455 (N_11455,N_11181,N_11231);
nand U11456 (N_11456,N_11089,N_11014);
xor U11457 (N_11457,N_11241,N_11138);
or U11458 (N_11458,N_11027,N_11185);
and U11459 (N_11459,N_11022,N_11139);
nor U11460 (N_11460,N_11040,N_11224);
nand U11461 (N_11461,N_11165,N_11089);
nor U11462 (N_11462,N_11189,N_11099);
or U11463 (N_11463,N_11159,N_11137);
and U11464 (N_11464,N_11234,N_11063);
xor U11465 (N_11465,N_11082,N_11200);
and U11466 (N_11466,N_11024,N_11066);
xnor U11467 (N_11467,N_11029,N_11207);
nor U11468 (N_11468,N_11082,N_11023);
xnor U11469 (N_11469,N_11151,N_11038);
nor U11470 (N_11470,N_11087,N_11092);
nand U11471 (N_11471,N_11173,N_11150);
and U11472 (N_11472,N_11022,N_11075);
nor U11473 (N_11473,N_11190,N_11187);
nand U11474 (N_11474,N_11116,N_11074);
nand U11475 (N_11475,N_11181,N_11180);
xnor U11476 (N_11476,N_11249,N_11048);
and U11477 (N_11477,N_11238,N_11204);
and U11478 (N_11478,N_11018,N_11199);
nor U11479 (N_11479,N_11042,N_11076);
nand U11480 (N_11480,N_11226,N_11153);
and U11481 (N_11481,N_11168,N_11132);
or U11482 (N_11482,N_11021,N_11040);
xor U11483 (N_11483,N_11150,N_11179);
xnor U11484 (N_11484,N_11131,N_11091);
nor U11485 (N_11485,N_11132,N_11032);
or U11486 (N_11486,N_11208,N_11161);
and U11487 (N_11487,N_11229,N_11184);
or U11488 (N_11488,N_11068,N_11207);
or U11489 (N_11489,N_11008,N_11234);
nand U11490 (N_11490,N_11244,N_11128);
nor U11491 (N_11491,N_11062,N_11059);
or U11492 (N_11492,N_11116,N_11010);
and U11493 (N_11493,N_11147,N_11028);
nand U11494 (N_11494,N_11106,N_11021);
xnor U11495 (N_11495,N_11068,N_11228);
nand U11496 (N_11496,N_11148,N_11089);
or U11497 (N_11497,N_11155,N_11128);
xnor U11498 (N_11498,N_11228,N_11133);
nand U11499 (N_11499,N_11183,N_11173);
nor U11500 (N_11500,N_11499,N_11314);
and U11501 (N_11501,N_11487,N_11444);
nand U11502 (N_11502,N_11372,N_11349);
xnor U11503 (N_11503,N_11262,N_11451);
xor U11504 (N_11504,N_11343,N_11332);
nor U11505 (N_11505,N_11449,N_11356);
and U11506 (N_11506,N_11261,N_11410);
nand U11507 (N_11507,N_11497,N_11468);
or U11508 (N_11508,N_11279,N_11369);
and U11509 (N_11509,N_11429,N_11266);
xor U11510 (N_11510,N_11294,N_11267);
and U11511 (N_11511,N_11309,N_11387);
xor U11512 (N_11512,N_11443,N_11341);
or U11513 (N_11513,N_11482,N_11424);
nor U11514 (N_11514,N_11463,N_11345);
and U11515 (N_11515,N_11300,N_11358);
or U11516 (N_11516,N_11475,N_11278);
and U11517 (N_11517,N_11337,N_11286);
xnor U11518 (N_11518,N_11269,N_11447);
or U11519 (N_11519,N_11400,N_11318);
or U11520 (N_11520,N_11473,N_11275);
and U11521 (N_11521,N_11273,N_11256);
nand U11522 (N_11522,N_11394,N_11464);
nor U11523 (N_11523,N_11265,N_11259);
and U11524 (N_11524,N_11385,N_11493);
xnor U11525 (N_11525,N_11362,N_11373);
and U11526 (N_11526,N_11289,N_11287);
xor U11527 (N_11527,N_11455,N_11371);
and U11528 (N_11528,N_11317,N_11325);
nand U11529 (N_11529,N_11353,N_11474);
nor U11530 (N_11530,N_11333,N_11411);
xor U11531 (N_11531,N_11305,N_11321);
xor U11532 (N_11532,N_11389,N_11361);
and U11533 (N_11533,N_11340,N_11360);
or U11534 (N_11534,N_11351,N_11396);
and U11535 (N_11535,N_11498,N_11397);
or U11536 (N_11536,N_11303,N_11272);
nor U11537 (N_11537,N_11288,N_11291);
or U11538 (N_11538,N_11476,N_11307);
nor U11539 (N_11539,N_11326,N_11485);
and U11540 (N_11540,N_11384,N_11460);
or U11541 (N_11541,N_11430,N_11324);
and U11542 (N_11542,N_11442,N_11469);
nand U11543 (N_11543,N_11403,N_11328);
or U11544 (N_11544,N_11470,N_11479);
or U11545 (N_11545,N_11408,N_11329);
nor U11546 (N_11546,N_11282,N_11330);
or U11547 (N_11547,N_11494,N_11402);
nand U11548 (N_11548,N_11458,N_11301);
nor U11549 (N_11549,N_11364,N_11375);
and U11550 (N_11550,N_11370,N_11454);
nand U11551 (N_11551,N_11365,N_11441);
nand U11552 (N_11552,N_11334,N_11290);
or U11553 (N_11553,N_11302,N_11298);
and U11554 (N_11554,N_11417,N_11274);
or U11555 (N_11555,N_11270,N_11407);
xor U11556 (N_11556,N_11338,N_11415);
or U11557 (N_11557,N_11486,N_11393);
and U11558 (N_11558,N_11462,N_11435);
nand U11559 (N_11559,N_11461,N_11355);
and U11560 (N_11560,N_11392,N_11336);
nand U11561 (N_11561,N_11354,N_11357);
and U11562 (N_11562,N_11453,N_11496);
or U11563 (N_11563,N_11297,N_11299);
and U11564 (N_11564,N_11280,N_11439);
xnor U11565 (N_11565,N_11374,N_11271);
or U11566 (N_11566,N_11450,N_11490);
or U11567 (N_11567,N_11346,N_11315);
xor U11568 (N_11568,N_11320,N_11283);
nand U11569 (N_11569,N_11304,N_11477);
nand U11570 (N_11570,N_11412,N_11457);
and U11571 (N_11571,N_11401,N_11339);
nand U11572 (N_11572,N_11446,N_11255);
nor U11573 (N_11573,N_11292,N_11434);
xor U11574 (N_11574,N_11311,N_11491);
or U11575 (N_11575,N_11319,N_11478);
xnor U11576 (N_11576,N_11293,N_11347);
or U11577 (N_11577,N_11484,N_11495);
nand U11578 (N_11578,N_11363,N_11483);
nand U11579 (N_11579,N_11335,N_11310);
or U11580 (N_11580,N_11465,N_11359);
and U11581 (N_11581,N_11331,N_11448);
and U11582 (N_11582,N_11428,N_11382);
nand U11583 (N_11583,N_11268,N_11257);
and U11584 (N_11584,N_11492,N_11284);
or U11585 (N_11585,N_11308,N_11432);
nor U11586 (N_11586,N_11431,N_11426);
and U11587 (N_11587,N_11251,N_11250);
and U11588 (N_11588,N_11421,N_11344);
and U11589 (N_11589,N_11306,N_11253);
or U11590 (N_11590,N_11381,N_11433);
nor U11591 (N_11591,N_11348,N_11488);
nor U11592 (N_11592,N_11416,N_11377);
nand U11593 (N_11593,N_11263,N_11342);
nor U11594 (N_11594,N_11419,N_11350);
or U11595 (N_11595,N_11456,N_11471);
xor U11596 (N_11596,N_11391,N_11366);
xnor U11597 (N_11597,N_11489,N_11383);
nand U11598 (N_11598,N_11260,N_11388);
xnor U11599 (N_11599,N_11399,N_11409);
nand U11600 (N_11600,N_11425,N_11467);
nor U11601 (N_11601,N_11380,N_11277);
and U11602 (N_11602,N_11445,N_11480);
and U11603 (N_11603,N_11312,N_11395);
and U11604 (N_11604,N_11285,N_11313);
and U11605 (N_11605,N_11390,N_11472);
nand U11606 (N_11606,N_11405,N_11258);
nand U11607 (N_11607,N_11323,N_11376);
xor U11608 (N_11608,N_11368,N_11427);
xor U11609 (N_11609,N_11252,N_11367);
and U11610 (N_11610,N_11436,N_11440);
xor U11611 (N_11611,N_11438,N_11459);
nor U11612 (N_11612,N_11418,N_11404);
nor U11613 (N_11613,N_11420,N_11406);
xnor U11614 (N_11614,N_11281,N_11386);
nand U11615 (N_11615,N_11413,N_11423);
or U11616 (N_11616,N_11254,N_11452);
or U11617 (N_11617,N_11379,N_11481);
nor U11618 (N_11618,N_11276,N_11352);
nor U11619 (N_11619,N_11264,N_11378);
nand U11620 (N_11620,N_11296,N_11398);
xnor U11621 (N_11621,N_11414,N_11322);
and U11622 (N_11622,N_11437,N_11466);
and U11623 (N_11623,N_11316,N_11422);
and U11624 (N_11624,N_11295,N_11327);
and U11625 (N_11625,N_11485,N_11494);
and U11626 (N_11626,N_11308,N_11283);
nor U11627 (N_11627,N_11318,N_11293);
and U11628 (N_11628,N_11364,N_11494);
nand U11629 (N_11629,N_11449,N_11472);
nand U11630 (N_11630,N_11250,N_11446);
and U11631 (N_11631,N_11478,N_11494);
xor U11632 (N_11632,N_11458,N_11394);
nand U11633 (N_11633,N_11346,N_11447);
and U11634 (N_11634,N_11284,N_11377);
and U11635 (N_11635,N_11331,N_11451);
xnor U11636 (N_11636,N_11313,N_11482);
or U11637 (N_11637,N_11463,N_11431);
and U11638 (N_11638,N_11415,N_11394);
nand U11639 (N_11639,N_11376,N_11260);
nand U11640 (N_11640,N_11292,N_11483);
nor U11641 (N_11641,N_11367,N_11464);
xor U11642 (N_11642,N_11299,N_11322);
nand U11643 (N_11643,N_11299,N_11433);
or U11644 (N_11644,N_11307,N_11427);
or U11645 (N_11645,N_11412,N_11323);
nor U11646 (N_11646,N_11394,N_11427);
nand U11647 (N_11647,N_11359,N_11260);
xor U11648 (N_11648,N_11357,N_11407);
or U11649 (N_11649,N_11276,N_11307);
nor U11650 (N_11650,N_11251,N_11385);
xor U11651 (N_11651,N_11299,N_11367);
xnor U11652 (N_11652,N_11256,N_11408);
nor U11653 (N_11653,N_11258,N_11331);
or U11654 (N_11654,N_11280,N_11434);
nor U11655 (N_11655,N_11349,N_11466);
and U11656 (N_11656,N_11398,N_11353);
nand U11657 (N_11657,N_11253,N_11438);
nor U11658 (N_11658,N_11327,N_11334);
nand U11659 (N_11659,N_11406,N_11482);
nand U11660 (N_11660,N_11447,N_11451);
and U11661 (N_11661,N_11275,N_11470);
nor U11662 (N_11662,N_11420,N_11363);
nand U11663 (N_11663,N_11408,N_11259);
or U11664 (N_11664,N_11266,N_11370);
and U11665 (N_11665,N_11251,N_11325);
nor U11666 (N_11666,N_11367,N_11406);
or U11667 (N_11667,N_11353,N_11473);
nor U11668 (N_11668,N_11316,N_11457);
and U11669 (N_11669,N_11326,N_11281);
nand U11670 (N_11670,N_11255,N_11295);
xor U11671 (N_11671,N_11477,N_11349);
or U11672 (N_11672,N_11280,N_11461);
nand U11673 (N_11673,N_11284,N_11391);
and U11674 (N_11674,N_11474,N_11425);
and U11675 (N_11675,N_11355,N_11306);
xnor U11676 (N_11676,N_11455,N_11258);
or U11677 (N_11677,N_11330,N_11369);
nand U11678 (N_11678,N_11498,N_11420);
or U11679 (N_11679,N_11277,N_11322);
or U11680 (N_11680,N_11428,N_11419);
nor U11681 (N_11681,N_11375,N_11317);
nor U11682 (N_11682,N_11466,N_11385);
nor U11683 (N_11683,N_11336,N_11393);
nor U11684 (N_11684,N_11443,N_11368);
nand U11685 (N_11685,N_11337,N_11401);
and U11686 (N_11686,N_11490,N_11276);
nand U11687 (N_11687,N_11433,N_11275);
nand U11688 (N_11688,N_11494,N_11396);
nand U11689 (N_11689,N_11329,N_11266);
or U11690 (N_11690,N_11325,N_11341);
xor U11691 (N_11691,N_11316,N_11429);
or U11692 (N_11692,N_11356,N_11495);
or U11693 (N_11693,N_11319,N_11276);
and U11694 (N_11694,N_11286,N_11428);
xor U11695 (N_11695,N_11431,N_11464);
nor U11696 (N_11696,N_11273,N_11305);
or U11697 (N_11697,N_11312,N_11256);
nand U11698 (N_11698,N_11272,N_11277);
and U11699 (N_11699,N_11329,N_11269);
nor U11700 (N_11700,N_11319,N_11492);
xnor U11701 (N_11701,N_11487,N_11308);
nand U11702 (N_11702,N_11444,N_11442);
nand U11703 (N_11703,N_11305,N_11488);
or U11704 (N_11704,N_11373,N_11403);
xnor U11705 (N_11705,N_11342,N_11412);
and U11706 (N_11706,N_11257,N_11477);
xor U11707 (N_11707,N_11378,N_11421);
or U11708 (N_11708,N_11297,N_11374);
nor U11709 (N_11709,N_11391,N_11263);
xnor U11710 (N_11710,N_11388,N_11376);
and U11711 (N_11711,N_11286,N_11394);
or U11712 (N_11712,N_11469,N_11272);
nor U11713 (N_11713,N_11439,N_11339);
and U11714 (N_11714,N_11395,N_11321);
xor U11715 (N_11715,N_11342,N_11376);
and U11716 (N_11716,N_11334,N_11428);
and U11717 (N_11717,N_11407,N_11319);
nand U11718 (N_11718,N_11471,N_11391);
nand U11719 (N_11719,N_11272,N_11316);
and U11720 (N_11720,N_11316,N_11383);
and U11721 (N_11721,N_11490,N_11480);
nor U11722 (N_11722,N_11489,N_11313);
and U11723 (N_11723,N_11439,N_11392);
or U11724 (N_11724,N_11333,N_11493);
nand U11725 (N_11725,N_11403,N_11353);
nand U11726 (N_11726,N_11358,N_11282);
or U11727 (N_11727,N_11279,N_11388);
nand U11728 (N_11728,N_11466,N_11389);
and U11729 (N_11729,N_11466,N_11327);
xor U11730 (N_11730,N_11252,N_11279);
or U11731 (N_11731,N_11321,N_11311);
nand U11732 (N_11732,N_11463,N_11464);
and U11733 (N_11733,N_11413,N_11254);
nor U11734 (N_11734,N_11327,N_11376);
nor U11735 (N_11735,N_11313,N_11376);
nor U11736 (N_11736,N_11284,N_11365);
nand U11737 (N_11737,N_11443,N_11412);
nand U11738 (N_11738,N_11377,N_11407);
xor U11739 (N_11739,N_11465,N_11398);
nor U11740 (N_11740,N_11382,N_11339);
and U11741 (N_11741,N_11400,N_11294);
and U11742 (N_11742,N_11270,N_11347);
and U11743 (N_11743,N_11482,N_11465);
nor U11744 (N_11744,N_11459,N_11416);
nor U11745 (N_11745,N_11280,N_11447);
and U11746 (N_11746,N_11343,N_11435);
xor U11747 (N_11747,N_11413,N_11449);
and U11748 (N_11748,N_11256,N_11270);
nand U11749 (N_11749,N_11284,N_11476);
and U11750 (N_11750,N_11557,N_11594);
xnor U11751 (N_11751,N_11539,N_11609);
nand U11752 (N_11752,N_11650,N_11549);
nand U11753 (N_11753,N_11604,N_11649);
or U11754 (N_11754,N_11666,N_11714);
xor U11755 (N_11755,N_11631,N_11728);
nand U11756 (N_11756,N_11700,N_11507);
xnor U11757 (N_11757,N_11702,N_11677);
and U11758 (N_11758,N_11580,N_11566);
or U11759 (N_11759,N_11589,N_11737);
and U11760 (N_11760,N_11554,N_11526);
nand U11761 (N_11761,N_11538,N_11708);
xnor U11762 (N_11762,N_11721,N_11643);
nand U11763 (N_11763,N_11591,N_11640);
and U11764 (N_11764,N_11691,N_11656);
nand U11765 (N_11765,N_11681,N_11593);
xnor U11766 (N_11766,N_11583,N_11573);
or U11767 (N_11767,N_11610,N_11525);
xnor U11768 (N_11768,N_11732,N_11546);
xor U11769 (N_11769,N_11560,N_11688);
nor U11770 (N_11770,N_11603,N_11724);
xnor U11771 (N_11771,N_11717,N_11742);
nand U11772 (N_11772,N_11596,N_11586);
xnor U11773 (N_11773,N_11530,N_11633);
and U11774 (N_11774,N_11627,N_11613);
or U11775 (N_11775,N_11680,N_11703);
xnor U11776 (N_11776,N_11652,N_11731);
xnor U11777 (N_11777,N_11644,N_11520);
or U11778 (N_11778,N_11564,N_11535);
nor U11779 (N_11779,N_11692,N_11616);
nor U11780 (N_11780,N_11571,N_11660);
nand U11781 (N_11781,N_11563,N_11706);
nand U11782 (N_11782,N_11622,N_11661);
or U11783 (N_11783,N_11712,N_11541);
xor U11784 (N_11784,N_11522,N_11715);
nor U11785 (N_11785,N_11506,N_11602);
nand U11786 (N_11786,N_11518,N_11587);
xnor U11787 (N_11787,N_11555,N_11730);
nand U11788 (N_11788,N_11673,N_11572);
xor U11789 (N_11789,N_11588,N_11690);
or U11790 (N_11790,N_11705,N_11646);
and U11791 (N_11791,N_11701,N_11685);
and U11792 (N_11792,N_11598,N_11623);
nand U11793 (N_11793,N_11581,N_11567);
nor U11794 (N_11794,N_11519,N_11727);
nand U11795 (N_11795,N_11533,N_11606);
and U11796 (N_11796,N_11537,N_11720);
nand U11797 (N_11797,N_11707,N_11508);
or U11798 (N_11798,N_11693,N_11647);
nand U11799 (N_11799,N_11529,N_11632);
nor U11800 (N_11800,N_11618,N_11582);
or U11801 (N_11801,N_11628,N_11741);
or U11802 (N_11802,N_11653,N_11625);
nor U11803 (N_11803,N_11561,N_11745);
xnor U11804 (N_11804,N_11679,N_11663);
or U11805 (N_11805,N_11515,N_11542);
nand U11806 (N_11806,N_11501,N_11575);
nand U11807 (N_11807,N_11577,N_11574);
and U11808 (N_11808,N_11615,N_11619);
or U11809 (N_11809,N_11669,N_11699);
nor U11810 (N_11810,N_11734,N_11709);
or U11811 (N_11811,N_11686,N_11634);
xor U11812 (N_11812,N_11713,N_11551);
and U11813 (N_11813,N_11527,N_11639);
nand U11814 (N_11814,N_11553,N_11536);
or U11815 (N_11815,N_11614,N_11570);
and U11816 (N_11816,N_11547,N_11675);
nand U11817 (N_11817,N_11540,N_11735);
nand U11818 (N_11818,N_11523,N_11558);
nand U11819 (N_11819,N_11534,N_11543);
nand U11820 (N_11820,N_11642,N_11565);
and U11821 (N_11821,N_11621,N_11626);
nand U11822 (N_11822,N_11667,N_11722);
nor U11823 (N_11823,N_11504,N_11568);
and U11824 (N_11824,N_11704,N_11674);
and U11825 (N_11825,N_11683,N_11531);
nand U11826 (N_11826,N_11695,N_11739);
and U11827 (N_11827,N_11637,N_11636);
nand U11828 (N_11828,N_11716,N_11524);
nand U11829 (N_11829,N_11676,N_11658);
nor U11830 (N_11830,N_11548,N_11746);
or U11831 (N_11831,N_11694,N_11687);
nand U11832 (N_11832,N_11726,N_11592);
xnor U11833 (N_11833,N_11597,N_11559);
nor U11834 (N_11834,N_11678,N_11641);
xnor U11835 (N_11835,N_11725,N_11585);
nor U11836 (N_11836,N_11502,N_11648);
nor U11837 (N_11837,N_11729,N_11738);
nand U11838 (N_11838,N_11595,N_11612);
nor U11839 (N_11839,N_11620,N_11511);
xnor U11840 (N_11840,N_11599,N_11749);
and U11841 (N_11841,N_11509,N_11605);
nor U11842 (N_11842,N_11600,N_11576);
or U11843 (N_11843,N_11670,N_11513);
nand U11844 (N_11844,N_11645,N_11651);
xnor U11845 (N_11845,N_11552,N_11578);
nor U11846 (N_11846,N_11654,N_11635);
xnor U11847 (N_11847,N_11516,N_11723);
or U11848 (N_11848,N_11659,N_11744);
xor U11849 (N_11849,N_11521,N_11517);
nor U11850 (N_11850,N_11655,N_11664);
nand U11851 (N_11851,N_11733,N_11569);
or U11852 (N_11852,N_11689,N_11638);
xor U11853 (N_11853,N_11710,N_11611);
nand U11854 (N_11854,N_11514,N_11698);
xor U11855 (N_11855,N_11662,N_11697);
and U11856 (N_11856,N_11711,N_11607);
xor U11857 (N_11857,N_11624,N_11743);
nor U11858 (N_11858,N_11510,N_11528);
xnor U11859 (N_11859,N_11505,N_11748);
nor U11860 (N_11860,N_11696,N_11682);
xnor U11861 (N_11861,N_11562,N_11740);
or U11862 (N_11862,N_11630,N_11503);
xor U11863 (N_11863,N_11747,N_11665);
and U11864 (N_11864,N_11719,N_11590);
nor U11865 (N_11865,N_11584,N_11512);
nor U11866 (N_11866,N_11718,N_11608);
xor U11867 (N_11867,N_11671,N_11545);
nand U11868 (N_11868,N_11629,N_11672);
nor U11869 (N_11869,N_11579,N_11736);
nor U11870 (N_11870,N_11601,N_11617);
and U11871 (N_11871,N_11532,N_11500);
nor U11872 (N_11872,N_11556,N_11550);
nand U11873 (N_11873,N_11544,N_11657);
xor U11874 (N_11874,N_11684,N_11668);
nand U11875 (N_11875,N_11501,N_11510);
and U11876 (N_11876,N_11505,N_11736);
xor U11877 (N_11877,N_11700,N_11697);
nand U11878 (N_11878,N_11677,N_11636);
xor U11879 (N_11879,N_11668,N_11649);
or U11880 (N_11880,N_11727,N_11680);
or U11881 (N_11881,N_11718,N_11560);
nor U11882 (N_11882,N_11605,N_11679);
or U11883 (N_11883,N_11579,N_11544);
xnor U11884 (N_11884,N_11601,N_11724);
xor U11885 (N_11885,N_11508,N_11672);
nor U11886 (N_11886,N_11546,N_11666);
or U11887 (N_11887,N_11720,N_11556);
and U11888 (N_11888,N_11746,N_11632);
or U11889 (N_11889,N_11581,N_11545);
and U11890 (N_11890,N_11604,N_11684);
nor U11891 (N_11891,N_11728,N_11547);
and U11892 (N_11892,N_11587,N_11530);
and U11893 (N_11893,N_11675,N_11712);
nand U11894 (N_11894,N_11668,N_11555);
xnor U11895 (N_11895,N_11725,N_11688);
nor U11896 (N_11896,N_11545,N_11557);
or U11897 (N_11897,N_11576,N_11632);
nor U11898 (N_11898,N_11636,N_11727);
nand U11899 (N_11899,N_11597,N_11676);
and U11900 (N_11900,N_11558,N_11635);
or U11901 (N_11901,N_11569,N_11725);
or U11902 (N_11902,N_11524,N_11726);
or U11903 (N_11903,N_11511,N_11567);
nor U11904 (N_11904,N_11718,N_11666);
or U11905 (N_11905,N_11704,N_11546);
or U11906 (N_11906,N_11552,N_11646);
nor U11907 (N_11907,N_11726,N_11593);
and U11908 (N_11908,N_11563,N_11719);
and U11909 (N_11909,N_11688,N_11705);
xnor U11910 (N_11910,N_11518,N_11617);
nand U11911 (N_11911,N_11520,N_11609);
nor U11912 (N_11912,N_11656,N_11528);
xor U11913 (N_11913,N_11555,N_11559);
nor U11914 (N_11914,N_11581,N_11748);
or U11915 (N_11915,N_11686,N_11521);
nor U11916 (N_11916,N_11747,N_11680);
xnor U11917 (N_11917,N_11693,N_11590);
nand U11918 (N_11918,N_11572,N_11575);
or U11919 (N_11919,N_11610,N_11644);
nand U11920 (N_11920,N_11704,N_11569);
xor U11921 (N_11921,N_11520,N_11705);
xor U11922 (N_11922,N_11569,N_11711);
nand U11923 (N_11923,N_11564,N_11584);
xor U11924 (N_11924,N_11502,N_11604);
and U11925 (N_11925,N_11604,N_11691);
xnor U11926 (N_11926,N_11707,N_11668);
nand U11927 (N_11927,N_11640,N_11729);
xnor U11928 (N_11928,N_11699,N_11702);
xor U11929 (N_11929,N_11578,N_11517);
nand U11930 (N_11930,N_11700,N_11559);
nor U11931 (N_11931,N_11526,N_11591);
nor U11932 (N_11932,N_11542,N_11708);
xnor U11933 (N_11933,N_11655,N_11724);
xnor U11934 (N_11934,N_11621,N_11741);
or U11935 (N_11935,N_11619,N_11637);
nor U11936 (N_11936,N_11702,N_11548);
xor U11937 (N_11937,N_11579,N_11551);
and U11938 (N_11938,N_11621,N_11718);
nor U11939 (N_11939,N_11604,N_11723);
or U11940 (N_11940,N_11518,N_11664);
nand U11941 (N_11941,N_11653,N_11703);
or U11942 (N_11942,N_11589,N_11540);
xnor U11943 (N_11943,N_11548,N_11599);
nand U11944 (N_11944,N_11535,N_11563);
xor U11945 (N_11945,N_11662,N_11522);
or U11946 (N_11946,N_11685,N_11552);
xnor U11947 (N_11947,N_11724,N_11581);
nor U11948 (N_11948,N_11563,N_11596);
nand U11949 (N_11949,N_11546,N_11663);
or U11950 (N_11950,N_11668,N_11611);
xnor U11951 (N_11951,N_11505,N_11519);
nand U11952 (N_11952,N_11654,N_11538);
nor U11953 (N_11953,N_11694,N_11572);
nand U11954 (N_11954,N_11548,N_11624);
or U11955 (N_11955,N_11655,N_11721);
or U11956 (N_11956,N_11627,N_11702);
nor U11957 (N_11957,N_11657,N_11567);
xnor U11958 (N_11958,N_11733,N_11707);
nor U11959 (N_11959,N_11676,N_11732);
nand U11960 (N_11960,N_11734,N_11596);
or U11961 (N_11961,N_11622,N_11517);
xor U11962 (N_11962,N_11707,N_11711);
and U11963 (N_11963,N_11697,N_11539);
nand U11964 (N_11964,N_11547,N_11542);
nor U11965 (N_11965,N_11528,N_11628);
xnor U11966 (N_11966,N_11736,N_11519);
and U11967 (N_11967,N_11586,N_11537);
and U11968 (N_11968,N_11658,N_11737);
xnor U11969 (N_11969,N_11666,N_11698);
xor U11970 (N_11970,N_11723,N_11596);
xnor U11971 (N_11971,N_11733,N_11739);
or U11972 (N_11972,N_11703,N_11626);
or U11973 (N_11973,N_11585,N_11537);
nor U11974 (N_11974,N_11543,N_11646);
nand U11975 (N_11975,N_11525,N_11697);
nand U11976 (N_11976,N_11643,N_11733);
nor U11977 (N_11977,N_11696,N_11742);
nand U11978 (N_11978,N_11582,N_11655);
nand U11979 (N_11979,N_11735,N_11693);
xnor U11980 (N_11980,N_11529,N_11644);
and U11981 (N_11981,N_11545,N_11715);
and U11982 (N_11982,N_11651,N_11575);
and U11983 (N_11983,N_11516,N_11565);
and U11984 (N_11984,N_11651,N_11557);
nand U11985 (N_11985,N_11724,N_11696);
or U11986 (N_11986,N_11682,N_11674);
or U11987 (N_11987,N_11658,N_11537);
nand U11988 (N_11988,N_11584,N_11514);
or U11989 (N_11989,N_11695,N_11558);
nor U11990 (N_11990,N_11501,N_11547);
and U11991 (N_11991,N_11638,N_11595);
xnor U11992 (N_11992,N_11532,N_11695);
nor U11993 (N_11993,N_11718,N_11705);
nor U11994 (N_11994,N_11524,N_11549);
xor U11995 (N_11995,N_11607,N_11744);
xnor U11996 (N_11996,N_11659,N_11746);
and U11997 (N_11997,N_11540,N_11695);
nor U11998 (N_11998,N_11546,N_11545);
nor U11999 (N_11999,N_11630,N_11717);
nand U12000 (N_12000,N_11751,N_11953);
nand U12001 (N_12001,N_11904,N_11846);
nand U12002 (N_12002,N_11948,N_11930);
or U12003 (N_12003,N_11901,N_11884);
xor U12004 (N_12004,N_11760,N_11862);
xnor U12005 (N_12005,N_11844,N_11783);
nand U12006 (N_12006,N_11972,N_11796);
nor U12007 (N_12007,N_11855,N_11755);
nand U12008 (N_12008,N_11975,N_11898);
nor U12009 (N_12009,N_11807,N_11778);
or U12010 (N_12010,N_11922,N_11759);
or U12011 (N_12011,N_11874,N_11978);
xnor U12012 (N_12012,N_11985,N_11771);
or U12013 (N_12013,N_11879,N_11983);
xor U12014 (N_12014,N_11761,N_11940);
nor U12015 (N_12015,N_11750,N_11960);
and U12016 (N_12016,N_11765,N_11961);
or U12017 (N_12017,N_11753,N_11838);
or U12018 (N_12018,N_11909,N_11872);
nand U12019 (N_12019,N_11908,N_11896);
xnor U12020 (N_12020,N_11925,N_11852);
or U12021 (N_12021,N_11918,N_11957);
or U12022 (N_12022,N_11973,N_11780);
or U12023 (N_12023,N_11934,N_11938);
nor U12024 (N_12024,N_11882,N_11890);
nand U12025 (N_12025,N_11829,N_11928);
and U12026 (N_12026,N_11979,N_11955);
or U12027 (N_12027,N_11980,N_11757);
and U12028 (N_12028,N_11790,N_11939);
nor U12029 (N_12029,N_11993,N_11963);
nand U12030 (N_12030,N_11770,N_11839);
or U12031 (N_12031,N_11802,N_11769);
xor U12032 (N_12032,N_11830,N_11988);
nor U12033 (N_12033,N_11989,N_11917);
nand U12034 (N_12034,N_11817,N_11804);
xnor U12035 (N_12035,N_11854,N_11950);
nand U12036 (N_12036,N_11946,N_11792);
and U12037 (N_12037,N_11986,N_11810);
or U12038 (N_12038,N_11789,N_11767);
nor U12039 (N_12039,N_11840,N_11895);
or U12040 (N_12040,N_11870,N_11886);
or U12041 (N_12041,N_11808,N_11977);
nand U12042 (N_12042,N_11956,N_11856);
or U12043 (N_12043,N_11861,N_11818);
xor U12044 (N_12044,N_11784,N_11915);
or U12045 (N_12045,N_11837,N_11831);
xor U12046 (N_12046,N_11984,N_11793);
xnor U12047 (N_12047,N_11995,N_11777);
nor U12048 (N_12048,N_11774,N_11903);
nand U12049 (N_12049,N_11875,N_11819);
xor U12050 (N_12050,N_11869,N_11809);
nand U12051 (N_12051,N_11906,N_11987);
nor U12052 (N_12052,N_11924,N_11814);
xor U12053 (N_12053,N_11944,N_11942);
and U12054 (N_12054,N_11880,N_11954);
and U12055 (N_12055,N_11833,N_11974);
and U12056 (N_12056,N_11969,N_11785);
nand U12057 (N_12057,N_11899,N_11902);
and U12058 (N_12058,N_11763,N_11990);
and U12059 (N_12059,N_11991,N_11826);
nor U12060 (N_12060,N_11820,N_11965);
or U12061 (N_12061,N_11968,N_11834);
nor U12062 (N_12062,N_11877,N_11916);
xnor U12063 (N_12063,N_11821,N_11794);
nand U12064 (N_12064,N_11788,N_11900);
nand U12065 (N_12065,N_11923,N_11764);
xor U12066 (N_12066,N_11897,N_11883);
nor U12067 (N_12067,N_11920,N_11822);
nor U12068 (N_12068,N_11756,N_11997);
xnor U12069 (N_12069,N_11964,N_11813);
or U12070 (N_12070,N_11867,N_11781);
and U12071 (N_12071,N_11935,N_11982);
xor U12072 (N_12072,N_11888,N_11945);
nor U12073 (N_12073,N_11959,N_11931);
and U12074 (N_12074,N_11921,N_11805);
nand U12075 (N_12075,N_11871,N_11791);
nand U12076 (N_12076,N_11932,N_11943);
nor U12077 (N_12077,N_11803,N_11762);
nor U12078 (N_12078,N_11966,N_11999);
nand U12079 (N_12079,N_11912,N_11801);
nand U12080 (N_12080,N_11949,N_11787);
or U12081 (N_12081,N_11828,N_11779);
nand U12082 (N_12082,N_11845,N_11927);
or U12083 (N_12083,N_11892,N_11775);
or U12084 (N_12084,N_11911,N_11841);
nand U12085 (N_12085,N_11926,N_11768);
or U12086 (N_12086,N_11752,N_11849);
or U12087 (N_12087,N_11811,N_11981);
and U12088 (N_12088,N_11782,N_11952);
xnor U12089 (N_12089,N_11859,N_11848);
nor U12090 (N_12090,N_11976,N_11958);
and U12091 (N_12091,N_11891,N_11816);
nor U12092 (N_12092,N_11827,N_11815);
and U12093 (N_12093,N_11967,N_11893);
and U12094 (N_12094,N_11850,N_11951);
nand U12095 (N_12095,N_11864,N_11842);
and U12096 (N_12096,N_11876,N_11786);
nor U12097 (N_12097,N_11936,N_11878);
and U12098 (N_12098,N_11825,N_11835);
nor U12099 (N_12099,N_11772,N_11843);
and U12100 (N_12100,N_11933,N_11868);
and U12101 (N_12101,N_11797,N_11919);
xnor U12102 (N_12102,N_11863,N_11776);
and U12103 (N_12103,N_11941,N_11866);
nor U12104 (N_12104,N_11907,N_11798);
nor U12105 (N_12105,N_11851,N_11795);
nand U12106 (N_12106,N_11887,N_11836);
xor U12107 (N_12107,N_11799,N_11894);
or U12108 (N_12108,N_11847,N_11992);
and U12109 (N_12109,N_11937,N_11914);
and U12110 (N_12110,N_11800,N_11910);
nand U12111 (N_12111,N_11885,N_11929);
and U12112 (N_12112,N_11754,N_11970);
or U12113 (N_12113,N_11832,N_11998);
or U12114 (N_12114,N_11971,N_11857);
nor U12115 (N_12115,N_11913,N_11766);
and U12116 (N_12116,N_11873,N_11889);
xor U12117 (N_12117,N_11905,N_11758);
and U12118 (N_12118,N_11881,N_11994);
nand U12119 (N_12119,N_11996,N_11806);
nand U12120 (N_12120,N_11824,N_11773);
or U12121 (N_12121,N_11823,N_11962);
or U12122 (N_12122,N_11865,N_11860);
or U12123 (N_12123,N_11812,N_11858);
xnor U12124 (N_12124,N_11947,N_11853);
xor U12125 (N_12125,N_11838,N_11921);
or U12126 (N_12126,N_11824,N_11923);
nand U12127 (N_12127,N_11977,N_11893);
or U12128 (N_12128,N_11812,N_11940);
and U12129 (N_12129,N_11752,N_11993);
nand U12130 (N_12130,N_11767,N_11934);
nand U12131 (N_12131,N_11908,N_11933);
nand U12132 (N_12132,N_11878,N_11992);
or U12133 (N_12133,N_11817,N_11819);
nor U12134 (N_12134,N_11999,N_11823);
nand U12135 (N_12135,N_11927,N_11964);
nand U12136 (N_12136,N_11912,N_11785);
xnor U12137 (N_12137,N_11921,N_11893);
and U12138 (N_12138,N_11828,N_11849);
and U12139 (N_12139,N_11925,N_11838);
and U12140 (N_12140,N_11997,N_11937);
and U12141 (N_12141,N_11788,N_11851);
and U12142 (N_12142,N_11823,N_11856);
nor U12143 (N_12143,N_11775,N_11969);
nor U12144 (N_12144,N_11835,N_11913);
xor U12145 (N_12145,N_11759,N_11995);
nand U12146 (N_12146,N_11882,N_11880);
and U12147 (N_12147,N_11828,N_11813);
nor U12148 (N_12148,N_11825,N_11947);
nor U12149 (N_12149,N_11953,N_11991);
and U12150 (N_12150,N_11809,N_11922);
nor U12151 (N_12151,N_11813,N_11901);
and U12152 (N_12152,N_11910,N_11808);
xnor U12153 (N_12153,N_11935,N_11995);
and U12154 (N_12154,N_11751,N_11764);
nand U12155 (N_12155,N_11906,N_11944);
xnor U12156 (N_12156,N_11814,N_11838);
or U12157 (N_12157,N_11957,N_11991);
xor U12158 (N_12158,N_11894,N_11804);
nand U12159 (N_12159,N_11987,N_11812);
xnor U12160 (N_12160,N_11854,N_11968);
nand U12161 (N_12161,N_11971,N_11896);
and U12162 (N_12162,N_11803,N_11826);
nand U12163 (N_12163,N_11788,N_11933);
or U12164 (N_12164,N_11764,N_11890);
nor U12165 (N_12165,N_11779,N_11814);
xor U12166 (N_12166,N_11760,N_11876);
xnor U12167 (N_12167,N_11789,N_11885);
nand U12168 (N_12168,N_11934,N_11784);
or U12169 (N_12169,N_11869,N_11950);
and U12170 (N_12170,N_11934,N_11975);
and U12171 (N_12171,N_11872,N_11979);
nand U12172 (N_12172,N_11950,N_11876);
nor U12173 (N_12173,N_11940,N_11856);
nand U12174 (N_12174,N_11872,N_11898);
nand U12175 (N_12175,N_11797,N_11912);
nor U12176 (N_12176,N_11927,N_11848);
nor U12177 (N_12177,N_11851,N_11823);
or U12178 (N_12178,N_11808,N_11872);
nand U12179 (N_12179,N_11981,N_11909);
or U12180 (N_12180,N_11829,N_11764);
xnor U12181 (N_12181,N_11841,N_11993);
or U12182 (N_12182,N_11815,N_11790);
nor U12183 (N_12183,N_11853,N_11960);
and U12184 (N_12184,N_11971,N_11922);
and U12185 (N_12185,N_11896,N_11927);
nor U12186 (N_12186,N_11905,N_11943);
and U12187 (N_12187,N_11916,N_11893);
nor U12188 (N_12188,N_11809,N_11941);
nand U12189 (N_12189,N_11863,N_11819);
and U12190 (N_12190,N_11993,N_11839);
nor U12191 (N_12191,N_11827,N_11995);
nor U12192 (N_12192,N_11959,N_11761);
and U12193 (N_12193,N_11855,N_11851);
or U12194 (N_12194,N_11798,N_11914);
or U12195 (N_12195,N_11863,N_11853);
and U12196 (N_12196,N_11906,N_11941);
xnor U12197 (N_12197,N_11823,N_11943);
nor U12198 (N_12198,N_11797,N_11973);
and U12199 (N_12199,N_11865,N_11897);
or U12200 (N_12200,N_11918,N_11810);
and U12201 (N_12201,N_11900,N_11818);
or U12202 (N_12202,N_11813,N_11903);
xor U12203 (N_12203,N_11974,N_11961);
nand U12204 (N_12204,N_11911,N_11918);
nor U12205 (N_12205,N_11925,N_11943);
nand U12206 (N_12206,N_11839,N_11850);
and U12207 (N_12207,N_11875,N_11988);
or U12208 (N_12208,N_11930,N_11866);
or U12209 (N_12209,N_11984,N_11898);
and U12210 (N_12210,N_11773,N_11850);
xnor U12211 (N_12211,N_11853,N_11782);
or U12212 (N_12212,N_11999,N_11974);
nor U12213 (N_12213,N_11793,N_11921);
and U12214 (N_12214,N_11926,N_11932);
xnor U12215 (N_12215,N_11840,N_11916);
and U12216 (N_12216,N_11790,N_11874);
nand U12217 (N_12217,N_11814,N_11986);
and U12218 (N_12218,N_11936,N_11990);
nand U12219 (N_12219,N_11752,N_11827);
xnor U12220 (N_12220,N_11767,N_11855);
xor U12221 (N_12221,N_11979,N_11769);
and U12222 (N_12222,N_11846,N_11852);
xor U12223 (N_12223,N_11754,N_11967);
nor U12224 (N_12224,N_11885,N_11888);
nor U12225 (N_12225,N_11925,N_11788);
or U12226 (N_12226,N_11971,N_11994);
nor U12227 (N_12227,N_11909,N_11926);
nand U12228 (N_12228,N_11863,N_11879);
nor U12229 (N_12229,N_11991,N_11785);
nand U12230 (N_12230,N_11776,N_11919);
xnor U12231 (N_12231,N_11901,N_11764);
or U12232 (N_12232,N_11790,N_11996);
xnor U12233 (N_12233,N_11802,N_11973);
nand U12234 (N_12234,N_11876,N_11886);
or U12235 (N_12235,N_11861,N_11885);
nand U12236 (N_12236,N_11787,N_11993);
and U12237 (N_12237,N_11970,N_11774);
and U12238 (N_12238,N_11950,N_11810);
and U12239 (N_12239,N_11823,N_11889);
nand U12240 (N_12240,N_11782,N_11808);
or U12241 (N_12241,N_11902,N_11851);
xnor U12242 (N_12242,N_11856,N_11829);
or U12243 (N_12243,N_11789,N_11985);
or U12244 (N_12244,N_11760,N_11964);
nor U12245 (N_12245,N_11960,N_11879);
nand U12246 (N_12246,N_11875,N_11901);
or U12247 (N_12247,N_11974,N_11939);
xor U12248 (N_12248,N_11888,N_11764);
nand U12249 (N_12249,N_11881,N_11800);
or U12250 (N_12250,N_12093,N_12173);
xnor U12251 (N_12251,N_12113,N_12199);
nand U12252 (N_12252,N_12114,N_12068);
nor U12253 (N_12253,N_12181,N_12030);
or U12254 (N_12254,N_12134,N_12174);
or U12255 (N_12255,N_12154,N_12130);
xor U12256 (N_12256,N_12020,N_12131);
or U12257 (N_12257,N_12119,N_12015);
or U12258 (N_12258,N_12230,N_12115);
nor U12259 (N_12259,N_12249,N_12246);
xnor U12260 (N_12260,N_12140,N_12200);
nand U12261 (N_12261,N_12097,N_12108);
xnor U12262 (N_12262,N_12229,N_12214);
or U12263 (N_12263,N_12195,N_12079);
and U12264 (N_12264,N_12002,N_12009);
nor U12265 (N_12265,N_12024,N_12233);
or U12266 (N_12266,N_12117,N_12208);
xor U12267 (N_12267,N_12186,N_12071);
or U12268 (N_12268,N_12092,N_12087);
nand U12269 (N_12269,N_12135,N_12044);
nand U12270 (N_12270,N_12143,N_12047);
and U12271 (N_12271,N_12228,N_12045);
or U12272 (N_12272,N_12061,N_12172);
nand U12273 (N_12273,N_12083,N_12243);
xor U12274 (N_12274,N_12039,N_12125);
nand U12275 (N_12275,N_12217,N_12060);
nand U12276 (N_12276,N_12112,N_12150);
xnor U12277 (N_12277,N_12120,N_12185);
nand U12278 (N_12278,N_12162,N_12157);
nand U12279 (N_12279,N_12056,N_12042);
and U12280 (N_12280,N_12003,N_12189);
nor U12281 (N_12281,N_12239,N_12095);
xor U12282 (N_12282,N_12167,N_12212);
xor U12283 (N_12283,N_12025,N_12164);
nand U12284 (N_12284,N_12171,N_12098);
nor U12285 (N_12285,N_12161,N_12057);
nor U12286 (N_12286,N_12219,N_12192);
nand U12287 (N_12287,N_12197,N_12031);
and U12288 (N_12288,N_12000,N_12138);
or U12289 (N_12289,N_12067,N_12180);
xor U12290 (N_12290,N_12139,N_12218);
nor U12291 (N_12291,N_12160,N_12220);
nor U12292 (N_12292,N_12158,N_12211);
and U12293 (N_12293,N_12129,N_12017);
xnor U12294 (N_12294,N_12149,N_12038);
nand U12295 (N_12295,N_12175,N_12101);
xor U12296 (N_12296,N_12123,N_12032);
nor U12297 (N_12297,N_12078,N_12063);
and U12298 (N_12298,N_12238,N_12204);
or U12299 (N_12299,N_12145,N_12155);
or U12300 (N_12300,N_12035,N_12216);
nand U12301 (N_12301,N_12245,N_12178);
or U12302 (N_12302,N_12176,N_12247);
xnor U12303 (N_12303,N_12053,N_12111);
nand U12304 (N_12304,N_12116,N_12001);
or U12305 (N_12305,N_12077,N_12223);
xnor U12306 (N_12306,N_12187,N_12102);
xnor U12307 (N_12307,N_12037,N_12016);
xnor U12308 (N_12308,N_12148,N_12052);
and U12309 (N_12309,N_12069,N_12225);
or U12310 (N_12310,N_12036,N_12088);
nor U12311 (N_12311,N_12232,N_12051);
xor U12312 (N_12312,N_12075,N_12054);
xnor U12313 (N_12313,N_12007,N_12137);
nor U12314 (N_12314,N_12029,N_12151);
or U12315 (N_12315,N_12146,N_12182);
nand U12316 (N_12316,N_12207,N_12248);
nand U12317 (N_12317,N_12072,N_12221);
and U12318 (N_12318,N_12109,N_12065);
nand U12319 (N_12319,N_12118,N_12122);
and U12320 (N_12320,N_12226,N_12004);
nand U12321 (N_12321,N_12023,N_12234);
and U12322 (N_12322,N_12144,N_12177);
or U12323 (N_12323,N_12011,N_12086);
or U12324 (N_12324,N_12124,N_12188);
or U12325 (N_12325,N_12240,N_12099);
nand U12326 (N_12326,N_12074,N_12126);
or U12327 (N_12327,N_12106,N_12210);
nand U12328 (N_12328,N_12152,N_12190);
or U12329 (N_12329,N_12170,N_12222);
nor U12330 (N_12330,N_12046,N_12227);
and U12331 (N_12331,N_12048,N_12013);
or U12332 (N_12332,N_12209,N_12235);
or U12333 (N_12333,N_12085,N_12132);
and U12334 (N_12334,N_12136,N_12034);
or U12335 (N_12335,N_12159,N_12033);
or U12336 (N_12336,N_12121,N_12049);
nor U12337 (N_12337,N_12213,N_12165);
nand U12338 (N_12338,N_12191,N_12215);
or U12339 (N_12339,N_12066,N_12094);
and U12340 (N_12340,N_12163,N_12014);
nand U12341 (N_12341,N_12019,N_12147);
and U12342 (N_12342,N_12076,N_12169);
nor U12343 (N_12343,N_12059,N_12018);
nand U12344 (N_12344,N_12153,N_12107);
and U12345 (N_12345,N_12103,N_12242);
xnor U12346 (N_12346,N_12205,N_12105);
nor U12347 (N_12347,N_12082,N_12231);
and U12348 (N_12348,N_12201,N_12091);
xor U12349 (N_12349,N_12142,N_12168);
nor U12350 (N_12350,N_12008,N_12133);
nand U12351 (N_12351,N_12183,N_12110);
xor U12352 (N_12352,N_12028,N_12080);
nor U12353 (N_12353,N_12237,N_12202);
or U12354 (N_12354,N_12128,N_12179);
xnor U12355 (N_12355,N_12203,N_12058);
and U12356 (N_12356,N_12027,N_12198);
and U12357 (N_12357,N_12193,N_12194);
and U12358 (N_12358,N_12096,N_12062);
xnor U12359 (N_12359,N_12070,N_12184);
and U12360 (N_12360,N_12084,N_12026);
or U12361 (N_12361,N_12100,N_12021);
xor U12362 (N_12362,N_12156,N_12166);
or U12363 (N_12363,N_12236,N_12104);
xnor U12364 (N_12364,N_12141,N_12050);
or U12365 (N_12365,N_12081,N_12012);
nand U12366 (N_12366,N_12073,N_12244);
nand U12367 (N_12367,N_12005,N_12043);
nand U12368 (N_12368,N_12010,N_12064);
or U12369 (N_12369,N_12196,N_12089);
or U12370 (N_12370,N_12041,N_12224);
xor U12371 (N_12371,N_12206,N_12241);
and U12372 (N_12372,N_12090,N_12055);
or U12373 (N_12373,N_12127,N_12006);
xor U12374 (N_12374,N_12040,N_12022);
or U12375 (N_12375,N_12226,N_12181);
and U12376 (N_12376,N_12105,N_12033);
or U12377 (N_12377,N_12020,N_12000);
and U12378 (N_12378,N_12169,N_12034);
nand U12379 (N_12379,N_12125,N_12216);
nor U12380 (N_12380,N_12033,N_12023);
nor U12381 (N_12381,N_12152,N_12240);
xor U12382 (N_12382,N_12229,N_12233);
or U12383 (N_12383,N_12088,N_12181);
nor U12384 (N_12384,N_12245,N_12028);
and U12385 (N_12385,N_12061,N_12065);
or U12386 (N_12386,N_12204,N_12225);
xnor U12387 (N_12387,N_12088,N_12105);
nand U12388 (N_12388,N_12099,N_12155);
xnor U12389 (N_12389,N_12115,N_12240);
nor U12390 (N_12390,N_12144,N_12203);
xor U12391 (N_12391,N_12157,N_12165);
nor U12392 (N_12392,N_12236,N_12157);
nand U12393 (N_12393,N_12128,N_12172);
nand U12394 (N_12394,N_12031,N_12236);
nand U12395 (N_12395,N_12220,N_12123);
nor U12396 (N_12396,N_12019,N_12021);
nand U12397 (N_12397,N_12132,N_12241);
nand U12398 (N_12398,N_12000,N_12091);
nand U12399 (N_12399,N_12038,N_12237);
xor U12400 (N_12400,N_12139,N_12155);
xnor U12401 (N_12401,N_12113,N_12147);
xnor U12402 (N_12402,N_12029,N_12006);
nor U12403 (N_12403,N_12173,N_12025);
and U12404 (N_12404,N_12159,N_12093);
xor U12405 (N_12405,N_12210,N_12163);
xor U12406 (N_12406,N_12210,N_12223);
or U12407 (N_12407,N_12135,N_12107);
or U12408 (N_12408,N_12060,N_12079);
and U12409 (N_12409,N_12005,N_12152);
nor U12410 (N_12410,N_12052,N_12149);
nor U12411 (N_12411,N_12136,N_12009);
nor U12412 (N_12412,N_12221,N_12118);
nand U12413 (N_12413,N_12015,N_12110);
and U12414 (N_12414,N_12145,N_12175);
and U12415 (N_12415,N_12133,N_12205);
nor U12416 (N_12416,N_12051,N_12082);
or U12417 (N_12417,N_12173,N_12008);
and U12418 (N_12418,N_12040,N_12109);
or U12419 (N_12419,N_12089,N_12074);
nor U12420 (N_12420,N_12240,N_12237);
and U12421 (N_12421,N_12060,N_12017);
xor U12422 (N_12422,N_12158,N_12139);
nor U12423 (N_12423,N_12015,N_12002);
and U12424 (N_12424,N_12017,N_12055);
nand U12425 (N_12425,N_12237,N_12239);
or U12426 (N_12426,N_12093,N_12240);
or U12427 (N_12427,N_12126,N_12231);
nand U12428 (N_12428,N_12003,N_12068);
and U12429 (N_12429,N_12178,N_12065);
nor U12430 (N_12430,N_12138,N_12123);
nand U12431 (N_12431,N_12010,N_12114);
and U12432 (N_12432,N_12002,N_12133);
or U12433 (N_12433,N_12042,N_12039);
and U12434 (N_12434,N_12008,N_12040);
xnor U12435 (N_12435,N_12167,N_12126);
or U12436 (N_12436,N_12137,N_12198);
or U12437 (N_12437,N_12149,N_12136);
and U12438 (N_12438,N_12193,N_12062);
and U12439 (N_12439,N_12020,N_12127);
nand U12440 (N_12440,N_12176,N_12067);
or U12441 (N_12441,N_12228,N_12056);
and U12442 (N_12442,N_12137,N_12128);
nand U12443 (N_12443,N_12038,N_12210);
and U12444 (N_12444,N_12000,N_12093);
nor U12445 (N_12445,N_12234,N_12197);
nand U12446 (N_12446,N_12238,N_12128);
nor U12447 (N_12447,N_12215,N_12085);
nor U12448 (N_12448,N_12065,N_12062);
nand U12449 (N_12449,N_12011,N_12041);
xor U12450 (N_12450,N_12153,N_12066);
and U12451 (N_12451,N_12176,N_12119);
and U12452 (N_12452,N_12005,N_12237);
and U12453 (N_12453,N_12053,N_12240);
and U12454 (N_12454,N_12140,N_12057);
nor U12455 (N_12455,N_12031,N_12140);
xor U12456 (N_12456,N_12088,N_12167);
or U12457 (N_12457,N_12063,N_12180);
xnor U12458 (N_12458,N_12215,N_12233);
or U12459 (N_12459,N_12152,N_12228);
and U12460 (N_12460,N_12219,N_12098);
xnor U12461 (N_12461,N_12178,N_12024);
or U12462 (N_12462,N_12026,N_12136);
xor U12463 (N_12463,N_12133,N_12024);
or U12464 (N_12464,N_12122,N_12199);
and U12465 (N_12465,N_12162,N_12116);
nand U12466 (N_12466,N_12136,N_12100);
xnor U12467 (N_12467,N_12022,N_12186);
xnor U12468 (N_12468,N_12021,N_12015);
nand U12469 (N_12469,N_12245,N_12190);
and U12470 (N_12470,N_12118,N_12134);
and U12471 (N_12471,N_12100,N_12104);
xnor U12472 (N_12472,N_12232,N_12208);
nand U12473 (N_12473,N_12129,N_12043);
and U12474 (N_12474,N_12056,N_12153);
nand U12475 (N_12475,N_12021,N_12193);
nand U12476 (N_12476,N_12193,N_12165);
nand U12477 (N_12477,N_12195,N_12072);
and U12478 (N_12478,N_12174,N_12106);
xor U12479 (N_12479,N_12142,N_12162);
or U12480 (N_12480,N_12096,N_12237);
xor U12481 (N_12481,N_12042,N_12052);
nand U12482 (N_12482,N_12136,N_12107);
xnor U12483 (N_12483,N_12004,N_12003);
xnor U12484 (N_12484,N_12155,N_12112);
nor U12485 (N_12485,N_12072,N_12140);
or U12486 (N_12486,N_12160,N_12130);
or U12487 (N_12487,N_12025,N_12030);
xnor U12488 (N_12488,N_12035,N_12045);
xor U12489 (N_12489,N_12247,N_12119);
or U12490 (N_12490,N_12164,N_12179);
nor U12491 (N_12491,N_12078,N_12005);
or U12492 (N_12492,N_12084,N_12037);
or U12493 (N_12493,N_12125,N_12074);
xnor U12494 (N_12494,N_12080,N_12124);
or U12495 (N_12495,N_12228,N_12168);
nand U12496 (N_12496,N_12216,N_12205);
nand U12497 (N_12497,N_12242,N_12247);
or U12498 (N_12498,N_12040,N_12186);
nand U12499 (N_12499,N_12226,N_12192);
nor U12500 (N_12500,N_12364,N_12462);
xnor U12501 (N_12501,N_12468,N_12386);
nand U12502 (N_12502,N_12343,N_12328);
xor U12503 (N_12503,N_12342,N_12282);
xor U12504 (N_12504,N_12313,N_12287);
and U12505 (N_12505,N_12330,N_12493);
nor U12506 (N_12506,N_12374,N_12351);
nor U12507 (N_12507,N_12469,N_12266);
xor U12508 (N_12508,N_12329,N_12379);
nand U12509 (N_12509,N_12354,N_12339);
and U12510 (N_12510,N_12292,N_12293);
xnor U12511 (N_12511,N_12346,N_12263);
and U12512 (N_12512,N_12479,N_12410);
nand U12513 (N_12513,N_12481,N_12378);
nand U12514 (N_12514,N_12483,N_12412);
and U12515 (N_12515,N_12480,N_12419);
nor U12516 (N_12516,N_12411,N_12471);
and U12517 (N_12517,N_12448,N_12392);
and U12518 (N_12518,N_12432,N_12338);
xor U12519 (N_12519,N_12417,N_12256);
or U12520 (N_12520,N_12421,N_12439);
or U12521 (N_12521,N_12390,N_12358);
xnor U12522 (N_12522,N_12350,N_12490);
nand U12523 (N_12523,N_12436,N_12425);
nor U12524 (N_12524,N_12395,N_12359);
xor U12525 (N_12525,N_12445,N_12290);
and U12526 (N_12526,N_12265,N_12472);
nor U12527 (N_12527,N_12305,N_12482);
nor U12528 (N_12528,N_12435,N_12262);
or U12529 (N_12529,N_12406,N_12443);
and U12530 (N_12530,N_12405,N_12444);
nor U12531 (N_12531,N_12408,N_12487);
nand U12532 (N_12532,N_12294,N_12366);
or U12533 (N_12533,N_12474,N_12463);
nand U12534 (N_12534,N_12333,N_12401);
nor U12535 (N_12535,N_12324,N_12409);
xnor U12536 (N_12536,N_12486,N_12433);
and U12537 (N_12537,N_12459,N_12475);
or U12538 (N_12538,N_12377,N_12465);
nand U12539 (N_12539,N_12437,N_12428);
xor U12540 (N_12540,N_12326,N_12438);
nand U12541 (N_12541,N_12488,N_12347);
nor U12542 (N_12542,N_12309,N_12385);
and U12543 (N_12543,N_12283,N_12277);
xnor U12544 (N_12544,N_12356,N_12344);
and U12545 (N_12545,N_12306,N_12296);
and U12546 (N_12546,N_12272,N_12260);
or U12547 (N_12547,N_12253,N_12279);
nand U12548 (N_12548,N_12301,N_12431);
and U12549 (N_12549,N_12278,N_12460);
and U12550 (N_12550,N_12457,N_12461);
or U12551 (N_12551,N_12255,N_12372);
nor U12552 (N_12552,N_12335,N_12491);
nor U12553 (N_12553,N_12496,N_12414);
nor U12554 (N_12554,N_12456,N_12319);
nor U12555 (N_12555,N_12284,N_12434);
or U12556 (N_12556,N_12275,N_12316);
xnor U12557 (N_12557,N_12302,N_12273);
or U12558 (N_12558,N_12363,N_12494);
nand U12559 (N_12559,N_12349,N_12447);
nand U12560 (N_12560,N_12391,N_12477);
nor U12561 (N_12561,N_12375,N_12394);
and U12562 (N_12562,N_12258,N_12402);
and U12563 (N_12563,N_12357,N_12365);
nor U12564 (N_12564,N_12449,N_12452);
nand U12565 (N_12565,N_12424,N_12369);
xor U12566 (N_12566,N_12300,N_12389);
nand U12567 (N_12567,N_12362,N_12478);
nor U12568 (N_12568,N_12484,N_12336);
or U12569 (N_12569,N_12257,N_12345);
nor U12570 (N_12570,N_12413,N_12250);
xnor U12571 (N_12571,N_12495,N_12485);
or U12572 (N_12572,N_12321,N_12426);
xor U12573 (N_12573,N_12361,N_12367);
and U12574 (N_12574,N_12322,N_12458);
and U12575 (N_12575,N_12397,N_12427);
and U12576 (N_12576,N_12418,N_12286);
nor U12577 (N_12577,N_12360,N_12476);
nand U12578 (N_12578,N_12341,N_12276);
nand U12579 (N_12579,N_12274,N_12308);
and U12580 (N_12580,N_12314,N_12289);
nor U12581 (N_12581,N_12251,N_12499);
and U12582 (N_12582,N_12353,N_12489);
xor U12583 (N_12583,N_12252,N_12285);
nand U12584 (N_12584,N_12270,N_12403);
nor U12585 (N_12585,N_12298,N_12430);
xnor U12586 (N_12586,N_12454,N_12268);
and U12587 (N_12587,N_12381,N_12291);
xor U12588 (N_12588,N_12370,N_12295);
nand U12589 (N_12589,N_12384,N_12254);
or U12590 (N_12590,N_12323,N_12376);
nand U12591 (N_12591,N_12399,N_12267);
nand U12592 (N_12592,N_12422,N_12334);
nand U12593 (N_12593,N_12441,N_12396);
and U12594 (N_12594,N_12470,N_12497);
xor U12595 (N_12595,N_12440,N_12311);
nor U12596 (N_12596,N_12492,N_12280);
xnor U12597 (N_12597,N_12467,N_12315);
and U12598 (N_12598,N_12498,N_12371);
nand U12599 (N_12599,N_12400,N_12320);
nand U12600 (N_12600,N_12310,N_12261);
nor U12601 (N_12601,N_12331,N_12352);
and U12602 (N_12602,N_12317,N_12325);
or U12603 (N_12603,N_12416,N_12393);
nor U12604 (N_12604,N_12380,N_12259);
xnor U12605 (N_12605,N_12451,N_12312);
and U12606 (N_12606,N_12383,N_12327);
nand U12607 (N_12607,N_12404,N_12382);
nand U12608 (N_12608,N_12423,N_12398);
or U12609 (N_12609,N_12332,N_12373);
nand U12610 (N_12610,N_12318,N_12368);
or U12611 (N_12611,N_12303,N_12281);
xor U12612 (N_12612,N_12307,N_12455);
nand U12613 (N_12613,N_12407,N_12453);
or U12614 (N_12614,N_12288,N_12387);
nor U12615 (N_12615,N_12297,N_12420);
xnor U12616 (N_12616,N_12429,N_12415);
xnor U12617 (N_12617,N_12299,N_12340);
or U12618 (N_12618,N_12388,N_12348);
xor U12619 (N_12619,N_12450,N_12355);
nor U12620 (N_12620,N_12466,N_12264);
nor U12621 (N_12621,N_12446,N_12442);
nor U12622 (N_12622,N_12337,N_12464);
xor U12623 (N_12623,N_12269,N_12271);
nor U12624 (N_12624,N_12304,N_12473);
nand U12625 (N_12625,N_12404,N_12332);
xnor U12626 (N_12626,N_12496,N_12417);
or U12627 (N_12627,N_12484,N_12333);
or U12628 (N_12628,N_12479,N_12450);
xor U12629 (N_12629,N_12480,N_12492);
and U12630 (N_12630,N_12392,N_12489);
nor U12631 (N_12631,N_12268,N_12399);
nor U12632 (N_12632,N_12472,N_12266);
nor U12633 (N_12633,N_12262,N_12338);
and U12634 (N_12634,N_12341,N_12383);
xnor U12635 (N_12635,N_12319,N_12391);
nor U12636 (N_12636,N_12479,N_12253);
or U12637 (N_12637,N_12478,N_12305);
xnor U12638 (N_12638,N_12414,N_12451);
or U12639 (N_12639,N_12311,N_12485);
xnor U12640 (N_12640,N_12480,N_12494);
and U12641 (N_12641,N_12368,N_12383);
nand U12642 (N_12642,N_12289,N_12306);
or U12643 (N_12643,N_12284,N_12312);
xnor U12644 (N_12644,N_12478,N_12396);
nor U12645 (N_12645,N_12281,N_12333);
and U12646 (N_12646,N_12266,N_12384);
nand U12647 (N_12647,N_12273,N_12380);
or U12648 (N_12648,N_12382,N_12492);
xor U12649 (N_12649,N_12455,N_12352);
nor U12650 (N_12650,N_12376,N_12329);
and U12651 (N_12651,N_12423,N_12330);
xnor U12652 (N_12652,N_12440,N_12338);
and U12653 (N_12653,N_12447,N_12262);
or U12654 (N_12654,N_12397,N_12374);
and U12655 (N_12655,N_12483,N_12277);
nand U12656 (N_12656,N_12467,N_12430);
or U12657 (N_12657,N_12340,N_12418);
or U12658 (N_12658,N_12375,N_12288);
nand U12659 (N_12659,N_12483,N_12259);
xor U12660 (N_12660,N_12475,N_12361);
and U12661 (N_12661,N_12255,N_12281);
nand U12662 (N_12662,N_12403,N_12354);
and U12663 (N_12663,N_12382,N_12357);
nor U12664 (N_12664,N_12310,N_12426);
nand U12665 (N_12665,N_12328,N_12319);
xnor U12666 (N_12666,N_12313,N_12345);
and U12667 (N_12667,N_12343,N_12427);
nand U12668 (N_12668,N_12271,N_12356);
or U12669 (N_12669,N_12289,N_12278);
xnor U12670 (N_12670,N_12464,N_12471);
xor U12671 (N_12671,N_12484,N_12278);
nor U12672 (N_12672,N_12351,N_12360);
nand U12673 (N_12673,N_12477,N_12312);
nand U12674 (N_12674,N_12358,N_12439);
and U12675 (N_12675,N_12302,N_12323);
xor U12676 (N_12676,N_12460,N_12302);
and U12677 (N_12677,N_12498,N_12397);
nor U12678 (N_12678,N_12473,N_12263);
nor U12679 (N_12679,N_12301,N_12295);
xor U12680 (N_12680,N_12482,N_12294);
and U12681 (N_12681,N_12409,N_12314);
and U12682 (N_12682,N_12468,N_12493);
or U12683 (N_12683,N_12472,N_12313);
xnor U12684 (N_12684,N_12326,N_12388);
xnor U12685 (N_12685,N_12318,N_12467);
and U12686 (N_12686,N_12400,N_12346);
nand U12687 (N_12687,N_12311,N_12496);
and U12688 (N_12688,N_12483,N_12421);
nand U12689 (N_12689,N_12378,N_12398);
nor U12690 (N_12690,N_12470,N_12329);
nand U12691 (N_12691,N_12322,N_12329);
and U12692 (N_12692,N_12286,N_12297);
or U12693 (N_12693,N_12494,N_12392);
nor U12694 (N_12694,N_12460,N_12344);
or U12695 (N_12695,N_12329,N_12381);
or U12696 (N_12696,N_12421,N_12327);
nor U12697 (N_12697,N_12317,N_12366);
or U12698 (N_12698,N_12364,N_12283);
nor U12699 (N_12699,N_12469,N_12390);
and U12700 (N_12700,N_12254,N_12479);
and U12701 (N_12701,N_12250,N_12376);
or U12702 (N_12702,N_12458,N_12404);
nor U12703 (N_12703,N_12451,N_12429);
xor U12704 (N_12704,N_12384,N_12332);
or U12705 (N_12705,N_12379,N_12303);
xnor U12706 (N_12706,N_12462,N_12273);
or U12707 (N_12707,N_12332,N_12371);
xnor U12708 (N_12708,N_12260,N_12261);
or U12709 (N_12709,N_12481,N_12456);
nor U12710 (N_12710,N_12482,N_12284);
and U12711 (N_12711,N_12302,N_12305);
xnor U12712 (N_12712,N_12299,N_12415);
xnor U12713 (N_12713,N_12370,N_12371);
or U12714 (N_12714,N_12308,N_12498);
nor U12715 (N_12715,N_12321,N_12293);
and U12716 (N_12716,N_12273,N_12456);
nor U12717 (N_12717,N_12424,N_12477);
xor U12718 (N_12718,N_12325,N_12272);
nor U12719 (N_12719,N_12369,N_12291);
or U12720 (N_12720,N_12454,N_12453);
nor U12721 (N_12721,N_12259,N_12480);
xor U12722 (N_12722,N_12337,N_12315);
xnor U12723 (N_12723,N_12361,N_12264);
nand U12724 (N_12724,N_12379,N_12431);
or U12725 (N_12725,N_12373,N_12289);
nor U12726 (N_12726,N_12289,N_12405);
nor U12727 (N_12727,N_12447,N_12269);
nand U12728 (N_12728,N_12452,N_12297);
xnor U12729 (N_12729,N_12456,N_12330);
and U12730 (N_12730,N_12471,N_12491);
nor U12731 (N_12731,N_12277,N_12350);
nor U12732 (N_12732,N_12259,N_12287);
xor U12733 (N_12733,N_12377,N_12480);
xor U12734 (N_12734,N_12251,N_12297);
nor U12735 (N_12735,N_12254,N_12441);
xnor U12736 (N_12736,N_12300,N_12324);
nand U12737 (N_12737,N_12387,N_12337);
or U12738 (N_12738,N_12352,N_12328);
nor U12739 (N_12739,N_12433,N_12301);
or U12740 (N_12740,N_12358,N_12308);
nand U12741 (N_12741,N_12465,N_12453);
nand U12742 (N_12742,N_12261,N_12441);
and U12743 (N_12743,N_12461,N_12278);
xnor U12744 (N_12744,N_12449,N_12380);
nand U12745 (N_12745,N_12407,N_12310);
nand U12746 (N_12746,N_12294,N_12443);
xor U12747 (N_12747,N_12291,N_12427);
nand U12748 (N_12748,N_12345,N_12376);
xor U12749 (N_12749,N_12387,N_12457);
and U12750 (N_12750,N_12662,N_12588);
nor U12751 (N_12751,N_12676,N_12720);
nor U12752 (N_12752,N_12749,N_12734);
nor U12753 (N_12753,N_12630,N_12637);
nand U12754 (N_12754,N_12555,N_12642);
and U12755 (N_12755,N_12505,N_12686);
and U12756 (N_12756,N_12681,N_12595);
and U12757 (N_12757,N_12671,N_12638);
nor U12758 (N_12758,N_12509,N_12668);
and U12759 (N_12759,N_12692,N_12738);
nand U12760 (N_12760,N_12551,N_12612);
xor U12761 (N_12761,N_12565,N_12733);
nor U12762 (N_12762,N_12573,N_12598);
and U12763 (N_12763,N_12504,N_12521);
or U12764 (N_12764,N_12552,N_12541);
and U12765 (N_12765,N_12589,N_12661);
or U12766 (N_12766,N_12506,N_12633);
and U12767 (N_12767,N_12643,N_12714);
and U12768 (N_12768,N_12512,N_12649);
nand U12769 (N_12769,N_12557,N_12539);
or U12770 (N_12770,N_12648,N_12583);
nor U12771 (N_12771,N_12655,N_12650);
or U12772 (N_12772,N_12625,N_12561);
nand U12773 (N_12773,N_12729,N_12663);
or U12774 (N_12774,N_12707,N_12695);
nor U12775 (N_12775,N_12568,N_12558);
and U12776 (N_12776,N_12702,N_12622);
nand U12777 (N_12777,N_12659,N_12629);
nand U12778 (N_12778,N_12654,N_12691);
and U12779 (N_12779,N_12617,N_12596);
nor U12780 (N_12780,N_12586,N_12678);
and U12781 (N_12781,N_12582,N_12605);
and U12782 (N_12782,N_12694,N_12682);
xnor U12783 (N_12783,N_12604,N_12571);
nor U12784 (N_12784,N_12653,N_12722);
or U12785 (N_12785,N_12546,N_12584);
and U12786 (N_12786,N_12687,N_12531);
xor U12787 (N_12787,N_12545,N_12549);
xor U12788 (N_12788,N_12743,N_12550);
nand U12789 (N_12789,N_12685,N_12665);
nand U12790 (N_12790,N_12741,N_12697);
nand U12791 (N_12791,N_12726,N_12658);
and U12792 (N_12792,N_12600,N_12574);
nand U12793 (N_12793,N_12587,N_12526);
xnor U12794 (N_12794,N_12689,N_12656);
xnor U12795 (N_12795,N_12579,N_12613);
xor U12796 (N_12796,N_12516,N_12543);
nor U12797 (N_12797,N_12511,N_12544);
nor U12798 (N_12798,N_12675,N_12652);
and U12799 (N_12799,N_12501,N_12632);
nand U12800 (N_12800,N_12581,N_12556);
nand U12801 (N_12801,N_12560,N_12519);
xor U12802 (N_12802,N_12507,N_12532);
nand U12803 (N_12803,N_12510,N_12537);
xnor U12804 (N_12804,N_12721,N_12747);
nand U12805 (N_12805,N_12708,N_12610);
nand U12806 (N_12806,N_12534,N_12576);
or U12807 (N_12807,N_12578,N_12683);
and U12808 (N_12808,N_12580,N_12730);
xor U12809 (N_12809,N_12706,N_12620);
nor U12810 (N_12810,N_12572,N_12614);
or U12811 (N_12811,N_12503,N_12684);
and U12812 (N_12812,N_12547,N_12674);
nor U12813 (N_12813,N_12530,N_12611);
xnor U12814 (N_12814,N_12575,N_12536);
nand U12815 (N_12815,N_12715,N_12524);
xor U12816 (N_12816,N_12615,N_12623);
nor U12817 (N_12817,N_12716,N_12677);
and U12818 (N_12818,N_12713,N_12562);
and U12819 (N_12819,N_12641,N_12701);
nor U12820 (N_12820,N_12732,N_12711);
xor U12821 (N_12821,N_12538,N_12728);
nand U12822 (N_12822,N_12592,N_12693);
nand U12823 (N_12823,N_12688,N_12626);
or U12824 (N_12824,N_12727,N_12705);
and U12825 (N_12825,N_12523,N_12528);
nor U12826 (N_12826,N_12670,N_12567);
xor U12827 (N_12827,N_12748,N_12508);
nand U12828 (N_12828,N_12651,N_12672);
and U12829 (N_12829,N_12680,N_12570);
nor U12830 (N_12830,N_12717,N_12522);
and U12831 (N_12831,N_12597,N_12513);
nor U12832 (N_12832,N_12569,N_12725);
or U12833 (N_12833,N_12599,N_12679);
or U12834 (N_12834,N_12603,N_12640);
nand U12835 (N_12835,N_12664,N_12529);
nor U12836 (N_12836,N_12628,N_12515);
or U12837 (N_12837,N_12517,N_12644);
xnor U12838 (N_12838,N_12608,N_12593);
xor U12839 (N_12839,N_12639,N_12673);
xor U12840 (N_12840,N_12616,N_12709);
nand U12841 (N_12841,N_12619,N_12627);
and U12842 (N_12842,N_12742,N_12563);
nand U12843 (N_12843,N_12636,N_12621);
and U12844 (N_12844,N_12718,N_12548);
or U12845 (N_12845,N_12591,N_12553);
or U12846 (N_12846,N_12525,N_12590);
or U12847 (N_12847,N_12699,N_12667);
xnor U12848 (N_12848,N_12696,N_12585);
xnor U12849 (N_12849,N_12533,N_12602);
nor U12850 (N_12850,N_12698,N_12564);
nand U12851 (N_12851,N_12527,N_12657);
and U12852 (N_12852,N_12739,N_12735);
nand U12853 (N_12853,N_12634,N_12624);
nor U12854 (N_12854,N_12645,N_12669);
nand U12855 (N_12855,N_12744,N_12594);
or U12856 (N_12856,N_12609,N_12737);
nand U12857 (N_12857,N_12745,N_12666);
xor U12858 (N_12858,N_12635,N_12746);
xor U12859 (N_12859,N_12631,N_12740);
and U12860 (N_12860,N_12618,N_12647);
nand U12861 (N_12861,N_12559,N_12700);
nand U12862 (N_12862,N_12646,N_12554);
or U12863 (N_12863,N_12731,N_12712);
or U12864 (N_12864,N_12719,N_12520);
and U12865 (N_12865,N_12502,N_12514);
xor U12866 (N_12866,N_12736,N_12566);
nand U12867 (N_12867,N_12607,N_12660);
xor U12868 (N_12868,N_12540,N_12724);
xor U12869 (N_12869,N_12690,N_12710);
and U12870 (N_12870,N_12518,N_12542);
nand U12871 (N_12871,N_12723,N_12535);
nor U12872 (N_12872,N_12601,N_12577);
nor U12873 (N_12873,N_12704,N_12703);
nand U12874 (N_12874,N_12500,N_12606);
nor U12875 (N_12875,N_12535,N_12635);
nand U12876 (N_12876,N_12593,N_12626);
and U12877 (N_12877,N_12613,N_12580);
nand U12878 (N_12878,N_12577,N_12731);
and U12879 (N_12879,N_12737,N_12693);
nand U12880 (N_12880,N_12525,N_12683);
or U12881 (N_12881,N_12740,N_12609);
xnor U12882 (N_12882,N_12657,N_12678);
xnor U12883 (N_12883,N_12538,N_12586);
and U12884 (N_12884,N_12732,N_12595);
nor U12885 (N_12885,N_12554,N_12538);
xor U12886 (N_12886,N_12710,N_12742);
and U12887 (N_12887,N_12551,N_12647);
and U12888 (N_12888,N_12607,N_12684);
and U12889 (N_12889,N_12578,N_12563);
xor U12890 (N_12890,N_12592,N_12686);
nor U12891 (N_12891,N_12541,N_12569);
xor U12892 (N_12892,N_12630,N_12617);
and U12893 (N_12893,N_12511,N_12683);
nand U12894 (N_12894,N_12724,N_12670);
nand U12895 (N_12895,N_12659,N_12603);
and U12896 (N_12896,N_12680,N_12633);
nor U12897 (N_12897,N_12671,N_12513);
xnor U12898 (N_12898,N_12544,N_12731);
xor U12899 (N_12899,N_12665,N_12641);
xnor U12900 (N_12900,N_12690,N_12584);
nor U12901 (N_12901,N_12602,N_12649);
and U12902 (N_12902,N_12622,N_12749);
xor U12903 (N_12903,N_12518,N_12688);
and U12904 (N_12904,N_12613,N_12619);
and U12905 (N_12905,N_12541,N_12673);
nand U12906 (N_12906,N_12595,N_12677);
or U12907 (N_12907,N_12693,N_12559);
nor U12908 (N_12908,N_12719,N_12575);
nor U12909 (N_12909,N_12749,N_12539);
and U12910 (N_12910,N_12591,N_12506);
nand U12911 (N_12911,N_12726,N_12506);
nand U12912 (N_12912,N_12675,N_12641);
or U12913 (N_12913,N_12630,N_12725);
and U12914 (N_12914,N_12723,N_12608);
and U12915 (N_12915,N_12592,N_12671);
nor U12916 (N_12916,N_12727,N_12669);
nor U12917 (N_12917,N_12679,N_12702);
nand U12918 (N_12918,N_12603,N_12651);
xnor U12919 (N_12919,N_12728,N_12590);
and U12920 (N_12920,N_12572,N_12512);
xnor U12921 (N_12921,N_12650,N_12641);
xnor U12922 (N_12922,N_12583,N_12532);
nor U12923 (N_12923,N_12734,N_12521);
xnor U12924 (N_12924,N_12543,N_12539);
or U12925 (N_12925,N_12695,N_12514);
nor U12926 (N_12926,N_12744,N_12598);
or U12927 (N_12927,N_12629,N_12552);
nand U12928 (N_12928,N_12572,N_12504);
xor U12929 (N_12929,N_12609,N_12699);
nand U12930 (N_12930,N_12562,N_12657);
or U12931 (N_12931,N_12611,N_12666);
or U12932 (N_12932,N_12501,N_12627);
nor U12933 (N_12933,N_12583,N_12557);
nand U12934 (N_12934,N_12665,N_12600);
and U12935 (N_12935,N_12663,N_12542);
or U12936 (N_12936,N_12624,N_12745);
or U12937 (N_12937,N_12643,N_12631);
and U12938 (N_12938,N_12733,N_12699);
nor U12939 (N_12939,N_12695,N_12725);
nand U12940 (N_12940,N_12635,N_12680);
and U12941 (N_12941,N_12680,N_12578);
nand U12942 (N_12942,N_12677,N_12679);
and U12943 (N_12943,N_12661,N_12645);
xnor U12944 (N_12944,N_12512,N_12622);
and U12945 (N_12945,N_12684,N_12675);
or U12946 (N_12946,N_12659,N_12563);
and U12947 (N_12947,N_12501,N_12713);
or U12948 (N_12948,N_12712,N_12598);
or U12949 (N_12949,N_12673,N_12737);
nand U12950 (N_12950,N_12579,N_12623);
nand U12951 (N_12951,N_12605,N_12679);
xor U12952 (N_12952,N_12628,N_12660);
and U12953 (N_12953,N_12517,N_12558);
xnor U12954 (N_12954,N_12671,N_12575);
nor U12955 (N_12955,N_12577,N_12663);
and U12956 (N_12956,N_12543,N_12550);
xor U12957 (N_12957,N_12587,N_12640);
nand U12958 (N_12958,N_12514,N_12708);
and U12959 (N_12959,N_12747,N_12577);
nand U12960 (N_12960,N_12721,N_12690);
or U12961 (N_12961,N_12539,N_12565);
xor U12962 (N_12962,N_12693,N_12744);
nand U12963 (N_12963,N_12724,N_12517);
or U12964 (N_12964,N_12625,N_12513);
xor U12965 (N_12965,N_12597,N_12503);
and U12966 (N_12966,N_12530,N_12679);
and U12967 (N_12967,N_12657,N_12504);
nand U12968 (N_12968,N_12697,N_12657);
nor U12969 (N_12969,N_12608,N_12552);
nor U12970 (N_12970,N_12728,N_12690);
nor U12971 (N_12971,N_12575,N_12741);
and U12972 (N_12972,N_12715,N_12608);
or U12973 (N_12973,N_12517,N_12685);
nor U12974 (N_12974,N_12581,N_12619);
nand U12975 (N_12975,N_12602,N_12641);
and U12976 (N_12976,N_12708,N_12599);
nor U12977 (N_12977,N_12731,N_12521);
or U12978 (N_12978,N_12690,N_12550);
nor U12979 (N_12979,N_12640,N_12581);
and U12980 (N_12980,N_12595,N_12650);
nand U12981 (N_12981,N_12738,N_12502);
xnor U12982 (N_12982,N_12610,N_12617);
nor U12983 (N_12983,N_12691,N_12723);
xnor U12984 (N_12984,N_12734,N_12690);
and U12985 (N_12985,N_12714,N_12621);
nand U12986 (N_12986,N_12639,N_12558);
or U12987 (N_12987,N_12520,N_12721);
nand U12988 (N_12988,N_12696,N_12641);
or U12989 (N_12989,N_12722,N_12614);
or U12990 (N_12990,N_12661,N_12698);
xnor U12991 (N_12991,N_12529,N_12731);
nand U12992 (N_12992,N_12648,N_12544);
xor U12993 (N_12993,N_12738,N_12593);
nand U12994 (N_12994,N_12727,N_12554);
or U12995 (N_12995,N_12584,N_12686);
nor U12996 (N_12996,N_12718,N_12712);
or U12997 (N_12997,N_12688,N_12618);
nor U12998 (N_12998,N_12666,N_12569);
and U12999 (N_12999,N_12728,N_12631);
nand U13000 (N_13000,N_12922,N_12827);
nand U13001 (N_13001,N_12866,N_12873);
nand U13002 (N_13002,N_12856,N_12841);
xnor U13003 (N_13003,N_12989,N_12778);
nand U13004 (N_13004,N_12983,N_12941);
and U13005 (N_13005,N_12790,N_12880);
xnor U13006 (N_13006,N_12946,N_12795);
and U13007 (N_13007,N_12882,N_12846);
or U13008 (N_13008,N_12998,N_12826);
nand U13009 (N_13009,N_12943,N_12945);
nand U13010 (N_13010,N_12937,N_12988);
nor U13011 (N_13011,N_12987,N_12949);
xor U13012 (N_13012,N_12973,N_12766);
nor U13013 (N_13013,N_12888,N_12854);
or U13014 (N_13014,N_12979,N_12847);
nor U13015 (N_13015,N_12972,N_12978);
xor U13016 (N_13016,N_12966,N_12984);
or U13017 (N_13017,N_12874,N_12883);
nand U13018 (N_13018,N_12954,N_12785);
and U13019 (N_13019,N_12812,N_12770);
or U13020 (N_13020,N_12982,N_12992);
nor U13021 (N_13021,N_12892,N_12980);
nand U13022 (N_13022,N_12898,N_12835);
nor U13023 (N_13023,N_12840,N_12993);
nor U13024 (N_13024,N_12833,N_12773);
or U13025 (N_13025,N_12764,N_12936);
xnor U13026 (N_13026,N_12905,N_12761);
nand U13027 (N_13027,N_12916,N_12800);
xor U13028 (N_13028,N_12959,N_12902);
and U13029 (N_13029,N_12801,N_12893);
nand U13030 (N_13030,N_12863,N_12806);
and U13031 (N_13031,N_12853,N_12895);
nand U13032 (N_13032,N_12926,N_12923);
nor U13033 (N_13033,N_12821,N_12828);
or U13034 (N_13034,N_12932,N_12901);
and U13035 (N_13035,N_12855,N_12877);
nor U13036 (N_13036,N_12900,N_12974);
or U13037 (N_13037,N_12842,N_12804);
and U13038 (N_13038,N_12951,N_12756);
or U13039 (N_13039,N_12997,N_12931);
and U13040 (N_13040,N_12849,N_12963);
and U13041 (N_13041,N_12875,N_12985);
xor U13042 (N_13042,N_12769,N_12844);
or U13043 (N_13043,N_12782,N_12861);
or U13044 (N_13044,N_12825,N_12890);
or U13045 (N_13045,N_12768,N_12869);
nand U13046 (N_13046,N_12798,N_12851);
nor U13047 (N_13047,N_12816,N_12948);
nand U13048 (N_13048,N_12817,N_12793);
and U13049 (N_13049,N_12969,N_12934);
and U13050 (N_13050,N_12789,N_12908);
xnor U13051 (N_13051,N_12794,N_12876);
and U13052 (N_13052,N_12956,N_12791);
xor U13053 (N_13053,N_12957,N_12837);
nor U13054 (N_13054,N_12942,N_12824);
nor U13055 (N_13055,N_12965,N_12788);
xnor U13056 (N_13056,N_12899,N_12811);
xor U13057 (N_13057,N_12935,N_12753);
nor U13058 (N_13058,N_12970,N_12832);
xor U13059 (N_13059,N_12810,N_12962);
nand U13060 (N_13060,N_12912,N_12792);
or U13061 (N_13061,N_12994,N_12903);
or U13062 (N_13062,N_12750,N_12759);
nand U13063 (N_13063,N_12975,N_12894);
xnor U13064 (N_13064,N_12848,N_12961);
nand U13065 (N_13065,N_12771,N_12868);
nand U13066 (N_13066,N_12781,N_12830);
nand U13067 (N_13067,N_12762,N_12885);
or U13068 (N_13068,N_12838,N_12917);
and U13069 (N_13069,N_12990,N_12952);
nor U13070 (N_13070,N_12843,N_12991);
nor U13071 (N_13071,N_12796,N_12818);
and U13072 (N_13072,N_12807,N_12813);
and U13073 (N_13073,N_12967,N_12907);
and U13074 (N_13074,N_12999,N_12822);
nor U13075 (N_13075,N_12995,N_12802);
nor U13076 (N_13076,N_12919,N_12865);
and U13077 (N_13077,N_12754,N_12808);
nand U13078 (N_13078,N_12797,N_12784);
xnor U13079 (N_13079,N_12918,N_12776);
and U13080 (N_13080,N_12889,N_12925);
nor U13081 (N_13081,N_12783,N_12938);
xor U13082 (N_13082,N_12976,N_12968);
or U13083 (N_13083,N_12953,N_12763);
or U13084 (N_13084,N_12870,N_12779);
xor U13085 (N_13085,N_12915,N_12755);
or U13086 (N_13086,N_12820,N_12777);
and U13087 (N_13087,N_12928,N_12864);
and U13088 (N_13088,N_12920,N_12887);
or U13089 (N_13089,N_12921,N_12947);
nand U13090 (N_13090,N_12891,N_12977);
or U13091 (N_13091,N_12872,N_12904);
or U13092 (N_13092,N_12960,N_12758);
or U13093 (N_13093,N_12772,N_12829);
nand U13094 (N_13094,N_12787,N_12867);
or U13095 (N_13095,N_12906,N_12859);
xor U13096 (N_13096,N_12751,N_12886);
xor U13097 (N_13097,N_12857,N_12819);
and U13098 (N_13098,N_12845,N_12958);
nand U13099 (N_13099,N_12775,N_12871);
nor U13100 (N_13100,N_12955,N_12757);
and U13101 (N_13101,N_12839,N_12814);
xor U13102 (N_13102,N_12913,N_12786);
and U13103 (N_13103,N_12809,N_12940);
nand U13104 (N_13104,N_12950,N_12860);
or U13105 (N_13105,N_12939,N_12927);
nor U13106 (N_13106,N_12858,N_12914);
nand U13107 (N_13107,N_12752,N_12981);
nand U13108 (N_13108,N_12836,N_12964);
nor U13109 (N_13109,N_12971,N_12852);
and U13110 (N_13110,N_12850,N_12911);
or U13111 (N_13111,N_12897,N_12996);
nand U13112 (N_13112,N_12933,N_12910);
nor U13113 (N_13113,N_12896,N_12815);
nand U13114 (N_13114,N_12803,N_12831);
nor U13115 (N_13115,N_12780,N_12834);
xnor U13116 (N_13116,N_12767,N_12929);
nor U13117 (N_13117,N_12884,N_12909);
and U13118 (N_13118,N_12799,N_12924);
or U13119 (N_13119,N_12805,N_12823);
nand U13120 (N_13120,N_12878,N_12944);
or U13121 (N_13121,N_12881,N_12774);
and U13122 (N_13122,N_12986,N_12765);
or U13123 (N_13123,N_12760,N_12879);
xor U13124 (N_13124,N_12930,N_12862);
nand U13125 (N_13125,N_12941,N_12970);
nor U13126 (N_13126,N_12978,N_12769);
nor U13127 (N_13127,N_12799,N_12832);
or U13128 (N_13128,N_12946,N_12840);
and U13129 (N_13129,N_12961,N_12875);
and U13130 (N_13130,N_12937,N_12916);
xnor U13131 (N_13131,N_12889,N_12954);
nand U13132 (N_13132,N_12883,N_12985);
nand U13133 (N_13133,N_12902,N_12933);
xor U13134 (N_13134,N_12941,N_12854);
xor U13135 (N_13135,N_12941,N_12872);
xor U13136 (N_13136,N_12977,N_12832);
and U13137 (N_13137,N_12924,N_12969);
nor U13138 (N_13138,N_12767,N_12751);
nor U13139 (N_13139,N_12909,N_12772);
or U13140 (N_13140,N_12854,N_12918);
nor U13141 (N_13141,N_12886,N_12935);
nand U13142 (N_13142,N_12983,N_12916);
or U13143 (N_13143,N_12798,N_12997);
xnor U13144 (N_13144,N_12986,N_12914);
nor U13145 (N_13145,N_12990,N_12805);
nor U13146 (N_13146,N_12804,N_12996);
nor U13147 (N_13147,N_12985,N_12876);
nand U13148 (N_13148,N_12847,N_12948);
or U13149 (N_13149,N_12991,N_12995);
nor U13150 (N_13150,N_12902,N_12883);
and U13151 (N_13151,N_12956,N_12921);
or U13152 (N_13152,N_12824,N_12948);
or U13153 (N_13153,N_12987,N_12776);
xor U13154 (N_13154,N_12989,N_12759);
and U13155 (N_13155,N_12941,N_12871);
xor U13156 (N_13156,N_12798,N_12806);
and U13157 (N_13157,N_12867,N_12838);
or U13158 (N_13158,N_12861,N_12938);
nand U13159 (N_13159,N_12953,N_12766);
or U13160 (N_13160,N_12919,N_12999);
or U13161 (N_13161,N_12796,N_12768);
and U13162 (N_13162,N_12813,N_12872);
nand U13163 (N_13163,N_12845,N_12849);
xnor U13164 (N_13164,N_12809,N_12797);
nand U13165 (N_13165,N_12952,N_12859);
and U13166 (N_13166,N_12862,N_12908);
xnor U13167 (N_13167,N_12819,N_12850);
nand U13168 (N_13168,N_12930,N_12863);
or U13169 (N_13169,N_12824,N_12878);
xor U13170 (N_13170,N_12888,N_12960);
nor U13171 (N_13171,N_12754,N_12799);
and U13172 (N_13172,N_12830,N_12751);
nand U13173 (N_13173,N_12913,N_12978);
and U13174 (N_13174,N_12884,N_12930);
or U13175 (N_13175,N_12823,N_12803);
nand U13176 (N_13176,N_12966,N_12969);
xnor U13177 (N_13177,N_12912,N_12814);
nor U13178 (N_13178,N_12756,N_12861);
or U13179 (N_13179,N_12936,N_12914);
or U13180 (N_13180,N_12980,N_12904);
nor U13181 (N_13181,N_12986,N_12955);
or U13182 (N_13182,N_12879,N_12801);
nand U13183 (N_13183,N_12757,N_12804);
nand U13184 (N_13184,N_12781,N_12779);
nor U13185 (N_13185,N_12963,N_12870);
and U13186 (N_13186,N_12766,N_12967);
xor U13187 (N_13187,N_12923,N_12928);
nor U13188 (N_13188,N_12857,N_12887);
nand U13189 (N_13189,N_12992,N_12865);
nor U13190 (N_13190,N_12956,N_12927);
xnor U13191 (N_13191,N_12759,N_12922);
and U13192 (N_13192,N_12838,N_12784);
nor U13193 (N_13193,N_12913,N_12969);
nor U13194 (N_13194,N_12950,N_12883);
and U13195 (N_13195,N_12968,N_12914);
nand U13196 (N_13196,N_12755,N_12916);
nand U13197 (N_13197,N_12895,N_12804);
nand U13198 (N_13198,N_12808,N_12993);
nand U13199 (N_13199,N_12785,N_12794);
xnor U13200 (N_13200,N_12787,N_12760);
and U13201 (N_13201,N_12900,N_12895);
and U13202 (N_13202,N_12811,N_12923);
nand U13203 (N_13203,N_12752,N_12784);
nor U13204 (N_13204,N_12940,N_12926);
xor U13205 (N_13205,N_12852,N_12961);
xnor U13206 (N_13206,N_12959,N_12944);
nand U13207 (N_13207,N_12923,N_12785);
or U13208 (N_13208,N_12975,N_12820);
and U13209 (N_13209,N_12943,N_12985);
xnor U13210 (N_13210,N_12877,N_12819);
and U13211 (N_13211,N_12996,N_12751);
nor U13212 (N_13212,N_12970,N_12753);
xnor U13213 (N_13213,N_12927,N_12806);
or U13214 (N_13214,N_12940,N_12942);
or U13215 (N_13215,N_12795,N_12813);
and U13216 (N_13216,N_12758,N_12987);
xnor U13217 (N_13217,N_12997,N_12769);
or U13218 (N_13218,N_12881,N_12901);
and U13219 (N_13219,N_12923,N_12924);
and U13220 (N_13220,N_12958,N_12831);
and U13221 (N_13221,N_12838,N_12989);
nor U13222 (N_13222,N_12975,N_12953);
nand U13223 (N_13223,N_12858,N_12962);
and U13224 (N_13224,N_12802,N_12800);
nor U13225 (N_13225,N_12820,N_12899);
and U13226 (N_13226,N_12932,N_12800);
nand U13227 (N_13227,N_12957,N_12768);
or U13228 (N_13228,N_12905,N_12843);
and U13229 (N_13229,N_12925,N_12766);
or U13230 (N_13230,N_12968,N_12787);
or U13231 (N_13231,N_12964,N_12775);
nor U13232 (N_13232,N_12877,N_12964);
nor U13233 (N_13233,N_12822,N_12804);
and U13234 (N_13234,N_12832,N_12997);
and U13235 (N_13235,N_12934,N_12819);
and U13236 (N_13236,N_12791,N_12887);
nor U13237 (N_13237,N_12799,N_12865);
and U13238 (N_13238,N_12870,N_12766);
and U13239 (N_13239,N_12795,N_12954);
nand U13240 (N_13240,N_12942,N_12933);
and U13241 (N_13241,N_12929,N_12848);
or U13242 (N_13242,N_12758,N_12861);
or U13243 (N_13243,N_12810,N_12882);
nor U13244 (N_13244,N_12888,N_12991);
xor U13245 (N_13245,N_12870,N_12842);
nor U13246 (N_13246,N_12937,N_12993);
xnor U13247 (N_13247,N_12947,N_12967);
nand U13248 (N_13248,N_12878,N_12772);
or U13249 (N_13249,N_12790,N_12872);
nor U13250 (N_13250,N_13146,N_13213);
nand U13251 (N_13251,N_13081,N_13182);
nand U13252 (N_13252,N_13050,N_13041);
nor U13253 (N_13253,N_13190,N_13038);
nand U13254 (N_13254,N_13226,N_13045);
and U13255 (N_13255,N_13234,N_13046);
or U13256 (N_13256,N_13012,N_13183);
and U13257 (N_13257,N_13002,N_13119);
or U13258 (N_13258,N_13205,N_13063);
and U13259 (N_13259,N_13096,N_13082);
and U13260 (N_13260,N_13169,N_13080);
or U13261 (N_13261,N_13061,N_13189);
xor U13262 (N_13262,N_13031,N_13125);
nand U13263 (N_13263,N_13152,N_13070);
or U13264 (N_13264,N_13037,N_13200);
nor U13265 (N_13265,N_13199,N_13043);
or U13266 (N_13266,N_13153,N_13073);
xor U13267 (N_13267,N_13239,N_13197);
and U13268 (N_13268,N_13042,N_13051);
and U13269 (N_13269,N_13033,N_13140);
nand U13270 (N_13270,N_13206,N_13222);
or U13271 (N_13271,N_13230,N_13207);
or U13272 (N_13272,N_13001,N_13009);
xor U13273 (N_13273,N_13139,N_13204);
nor U13274 (N_13274,N_13167,N_13118);
nand U13275 (N_13275,N_13157,N_13210);
and U13276 (N_13276,N_13220,N_13129);
nor U13277 (N_13277,N_13021,N_13191);
nand U13278 (N_13278,N_13128,N_13163);
and U13279 (N_13279,N_13006,N_13180);
nand U13280 (N_13280,N_13241,N_13121);
xnor U13281 (N_13281,N_13086,N_13236);
xor U13282 (N_13282,N_13104,N_13074);
xnor U13283 (N_13283,N_13211,N_13114);
nor U13284 (N_13284,N_13170,N_13148);
or U13285 (N_13285,N_13087,N_13245);
xnor U13286 (N_13286,N_13202,N_13177);
nand U13287 (N_13287,N_13229,N_13039);
and U13288 (N_13288,N_13161,N_13011);
nand U13289 (N_13289,N_13158,N_13126);
nor U13290 (N_13290,N_13243,N_13181);
and U13291 (N_13291,N_13151,N_13173);
nor U13292 (N_13292,N_13123,N_13249);
nand U13293 (N_13293,N_13069,N_13093);
xnor U13294 (N_13294,N_13075,N_13171);
or U13295 (N_13295,N_13088,N_13165);
or U13296 (N_13296,N_13116,N_13164);
nor U13297 (N_13297,N_13224,N_13195);
xor U13298 (N_13298,N_13036,N_13134);
and U13299 (N_13299,N_13055,N_13174);
nand U13300 (N_13300,N_13247,N_13184);
and U13301 (N_13301,N_13018,N_13168);
xor U13302 (N_13302,N_13099,N_13023);
nor U13303 (N_13303,N_13137,N_13192);
xnor U13304 (N_13304,N_13242,N_13185);
and U13305 (N_13305,N_13106,N_13112);
nor U13306 (N_13306,N_13113,N_13136);
nand U13307 (N_13307,N_13246,N_13024);
or U13308 (N_13308,N_13048,N_13107);
nand U13309 (N_13309,N_13067,N_13054);
or U13310 (N_13310,N_13193,N_13216);
nor U13311 (N_13311,N_13115,N_13143);
nor U13312 (N_13312,N_13060,N_13016);
or U13313 (N_13313,N_13231,N_13217);
and U13314 (N_13314,N_13237,N_13155);
nor U13315 (N_13315,N_13208,N_13223);
or U13316 (N_13316,N_13218,N_13227);
and U13317 (N_13317,N_13248,N_13221);
and U13318 (N_13318,N_13166,N_13003);
or U13319 (N_13319,N_13000,N_13147);
nor U13320 (N_13320,N_13117,N_13131);
and U13321 (N_13321,N_13138,N_13215);
nor U13322 (N_13322,N_13133,N_13065);
nor U13323 (N_13323,N_13201,N_13032);
nor U13324 (N_13324,N_13066,N_13029);
xnor U13325 (N_13325,N_13007,N_13035);
xnor U13326 (N_13326,N_13090,N_13240);
and U13327 (N_13327,N_13145,N_13219);
xnor U13328 (N_13328,N_13044,N_13110);
xnor U13329 (N_13329,N_13056,N_13127);
and U13330 (N_13330,N_13142,N_13076);
or U13331 (N_13331,N_13238,N_13130);
or U13332 (N_13332,N_13162,N_13228);
and U13333 (N_13333,N_13053,N_13034);
nand U13334 (N_13334,N_13052,N_13124);
and U13335 (N_13335,N_13178,N_13072);
nor U13336 (N_13336,N_13109,N_13233);
xor U13337 (N_13337,N_13194,N_13062);
or U13338 (N_13338,N_13186,N_13159);
or U13339 (N_13339,N_13111,N_13026);
nor U13340 (N_13340,N_13100,N_13103);
nand U13341 (N_13341,N_13049,N_13198);
xor U13342 (N_13342,N_13014,N_13244);
nor U13343 (N_13343,N_13179,N_13008);
nor U13344 (N_13344,N_13028,N_13025);
xnor U13345 (N_13345,N_13078,N_13089);
nor U13346 (N_13346,N_13122,N_13225);
nor U13347 (N_13347,N_13149,N_13156);
xor U13348 (N_13348,N_13172,N_13105);
or U13349 (N_13349,N_13141,N_13077);
xor U13350 (N_13350,N_13150,N_13098);
nor U13351 (N_13351,N_13132,N_13209);
or U13352 (N_13352,N_13059,N_13004);
or U13353 (N_13353,N_13203,N_13083);
and U13354 (N_13354,N_13010,N_13188);
nand U13355 (N_13355,N_13101,N_13092);
xnor U13356 (N_13356,N_13064,N_13097);
or U13357 (N_13357,N_13154,N_13068);
nand U13358 (N_13358,N_13108,N_13091);
or U13359 (N_13359,N_13017,N_13212);
or U13360 (N_13360,N_13022,N_13235);
or U13361 (N_13361,N_13160,N_13102);
xnor U13362 (N_13362,N_13071,N_13058);
and U13363 (N_13363,N_13196,N_13020);
xor U13364 (N_13364,N_13214,N_13094);
nor U13365 (N_13365,N_13013,N_13095);
xnor U13366 (N_13366,N_13144,N_13019);
or U13367 (N_13367,N_13176,N_13047);
or U13368 (N_13368,N_13187,N_13057);
nor U13369 (N_13369,N_13135,N_13120);
and U13370 (N_13370,N_13232,N_13079);
xor U13371 (N_13371,N_13085,N_13015);
nand U13372 (N_13372,N_13040,N_13005);
or U13373 (N_13373,N_13030,N_13027);
nand U13374 (N_13374,N_13084,N_13175);
or U13375 (N_13375,N_13129,N_13187);
or U13376 (N_13376,N_13198,N_13135);
and U13377 (N_13377,N_13177,N_13210);
nand U13378 (N_13378,N_13235,N_13246);
nand U13379 (N_13379,N_13029,N_13065);
xor U13380 (N_13380,N_13093,N_13081);
nor U13381 (N_13381,N_13068,N_13096);
and U13382 (N_13382,N_13176,N_13048);
nand U13383 (N_13383,N_13110,N_13028);
or U13384 (N_13384,N_13211,N_13207);
nor U13385 (N_13385,N_13166,N_13125);
nor U13386 (N_13386,N_13045,N_13128);
xnor U13387 (N_13387,N_13068,N_13210);
or U13388 (N_13388,N_13196,N_13199);
nor U13389 (N_13389,N_13132,N_13078);
nor U13390 (N_13390,N_13104,N_13070);
and U13391 (N_13391,N_13218,N_13153);
xnor U13392 (N_13392,N_13132,N_13030);
or U13393 (N_13393,N_13022,N_13225);
or U13394 (N_13394,N_13192,N_13111);
nor U13395 (N_13395,N_13078,N_13033);
or U13396 (N_13396,N_13167,N_13093);
nor U13397 (N_13397,N_13114,N_13144);
nand U13398 (N_13398,N_13160,N_13211);
xnor U13399 (N_13399,N_13100,N_13241);
nand U13400 (N_13400,N_13170,N_13039);
or U13401 (N_13401,N_13165,N_13180);
or U13402 (N_13402,N_13219,N_13125);
or U13403 (N_13403,N_13091,N_13077);
xor U13404 (N_13404,N_13096,N_13122);
xor U13405 (N_13405,N_13130,N_13096);
nor U13406 (N_13406,N_13059,N_13079);
nor U13407 (N_13407,N_13082,N_13026);
or U13408 (N_13408,N_13045,N_13059);
nand U13409 (N_13409,N_13001,N_13135);
nor U13410 (N_13410,N_13013,N_13023);
xor U13411 (N_13411,N_13031,N_13073);
xnor U13412 (N_13412,N_13034,N_13159);
nor U13413 (N_13413,N_13162,N_13085);
nor U13414 (N_13414,N_13229,N_13006);
nor U13415 (N_13415,N_13153,N_13063);
or U13416 (N_13416,N_13104,N_13041);
and U13417 (N_13417,N_13128,N_13086);
and U13418 (N_13418,N_13114,N_13089);
or U13419 (N_13419,N_13117,N_13144);
or U13420 (N_13420,N_13122,N_13094);
nand U13421 (N_13421,N_13108,N_13147);
nand U13422 (N_13422,N_13097,N_13225);
nand U13423 (N_13423,N_13023,N_13198);
or U13424 (N_13424,N_13103,N_13038);
and U13425 (N_13425,N_13140,N_13079);
or U13426 (N_13426,N_13075,N_13219);
and U13427 (N_13427,N_13015,N_13148);
xor U13428 (N_13428,N_13005,N_13180);
nand U13429 (N_13429,N_13128,N_13191);
nand U13430 (N_13430,N_13115,N_13153);
and U13431 (N_13431,N_13173,N_13220);
or U13432 (N_13432,N_13114,N_13035);
xnor U13433 (N_13433,N_13061,N_13154);
nand U13434 (N_13434,N_13195,N_13058);
xor U13435 (N_13435,N_13246,N_13040);
nor U13436 (N_13436,N_13023,N_13174);
xnor U13437 (N_13437,N_13184,N_13085);
and U13438 (N_13438,N_13181,N_13136);
xor U13439 (N_13439,N_13227,N_13074);
nor U13440 (N_13440,N_13139,N_13229);
nand U13441 (N_13441,N_13223,N_13000);
or U13442 (N_13442,N_13030,N_13249);
nand U13443 (N_13443,N_13133,N_13231);
and U13444 (N_13444,N_13231,N_13042);
or U13445 (N_13445,N_13228,N_13035);
xor U13446 (N_13446,N_13015,N_13230);
or U13447 (N_13447,N_13046,N_13196);
and U13448 (N_13448,N_13132,N_13105);
xnor U13449 (N_13449,N_13200,N_13022);
nand U13450 (N_13450,N_13167,N_13135);
nand U13451 (N_13451,N_13011,N_13127);
nand U13452 (N_13452,N_13108,N_13100);
or U13453 (N_13453,N_13005,N_13016);
and U13454 (N_13454,N_13036,N_13133);
or U13455 (N_13455,N_13206,N_13009);
nand U13456 (N_13456,N_13109,N_13074);
or U13457 (N_13457,N_13134,N_13076);
nor U13458 (N_13458,N_13123,N_13095);
and U13459 (N_13459,N_13209,N_13086);
nor U13460 (N_13460,N_13106,N_13030);
nand U13461 (N_13461,N_13097,N_13029);
and U13462 (N_13462,N_13086,N_13233);
and U13463 (N_13463,N_13142,N_13056);
nor U13464 (N_13464,N_13017,N_13244);
xnor U13465 (N_13465,N_13219,N_13198);
and U13466 (N_13466,N_13086,N_13178);
nand U13467 (N_13467,N_13220,N_13026);
nand U13468 (N_13468,N_13115,N_13038);
nor U13469 (N_13469,N_13222,N_13239);
nand U13470 (N_13470,N_13195,N_13149);
and U13471 (N_13471,N_13024,N_13110);
nor U13472 (N_13472,N_13106,N_13241);
or U13473 (N_13473,N_13103,N_13097);
or U13474 (N_13474,N_13192,N_13023);
nor U13475 (N_13475,N_13248,N_13049);
xor U13476 (N_13476,N_13113,N_13079);
nor U13477 (N_13477,N_13125,N_13041);
and U13478 (N_13478,N_13166,N_13169);
xor U13479 (N_13479,N_13072,N_13165);
or U13480 (N_13480,N_13145,N_13018);
nand U13481 (N_13481,N_13245,N_13214);
nand U13482 (N_13482,N_13163,N_13079);
or U13483 (N_13483,N_13058,N_13130);
and U13484 (N_13484,N_13082,N_13190);
or U13485 (N_13485,N_13084,N_13235);
xor U13486 (N_13486,N_13092,N_13127);
and U13487 (N_13487,N_13030,N_13148);
or U13488 (N_13488,N_13165,N_13136);
nor U13489 (N_13489,N_13143,N_13019);
or U13490 (N_13490,N_13074,N_13170);
nor U13491 (N_13491,N_13113,N_13184);
nand U13492 (N_13492,N_13083,N_13208);
or U13493 (N_13493,N_13087,N_13144);
xnor U13494 (N_13494,N_13199,N_13011);
nand U13495 (N_13495,N_13023,N_13026);
nand U13496 (N_13496,N_13171,N_13175);
nor U13497 (N_13497,N_13182,N_13188);
xor U13498 (N_13498,N_13154,N_13006);
nand U13499 (N_13499,N_13176,N_13014);
or U13500 (N_13500,N_13260,N_13469);
and U13501 (N_13501,N_13493,N_13452);
xor U13502 (N_13502,N_13278,N_13333);
nand U13503 (N_13503,N_13398,N_13303);
or U13504 (N_13504,N_13270,N_13450);
nand U13505 (N_13505,N_13297,N_13269);
nor U13506 (N_13506,N_13461,N_13313);
xnor U13507 (N_13507,N_13264,N_13390);
and U13508 (N_13508,N_13408,N_13361);
or U13509 (N_13509,N_13349,N_13419);
and U13510 (N_13510,N_13432,N_13251);
or U13511 (N_13511,N_13319,N_13271);
nor U13512 (N_13512,N_13388,N_13379);
nand U13513 (N_13513,N_13306,N_13327);
nor U13514 (N_13514,N_13287,N_13475);
and U13515 (N_13515,N_13410,N_13401);
and U13516 (N_13516,N_13321,N_13425);
nor U13517 (N_13517,N_13268,N_13371);
nor U13518 (N_13518,N_13355,N_13320);
nor U13519 (N_13519,N_13433,N_13441);
nand U13520 (N_13520,N_13274,N_13257);
xnor U13521 (N_13521,N_13487,N_13359);
and U13522 (N_13522,N_13498,N_13276);
nand U13523 (N_13523,N_13266,N_13395);
and U13524 (N_13524,N_13326,N_13434);
and U13525 (N_13525,N_13404,N_13442);
and U13526 (N_13526,N_13362,N_13440);
or U13527 (N_13527,N_13405,N_13284);
xnor U13528 (N_13528,N_13311,N_13288);
or U13529 (N_13529,N_13314,N_13343);
nand U13530 (N_13530,N_13275,N_13399);
and U13531 (N_13531,N_13444,N_13252);
or U13532 (N_13532,N_13344,N_13310);
nand U13533 (N_13533,N_13402,N_13483);
xor U13534 (N_13534,N_13439,N_13463);
nand U13535 (N_13535,N_13457,N_13340);
nand U13536 (N_13536,N_13367,N_13486);
or U13537 (N_13537,N_13446,N_13323);
or U13538 (N_13538,N_13467,N_13280);
or U13539 (N_13539,N_13345,N_13403);
or U13540 (N_13540,N_13392,N_13298);
and U13541 (N_13541,N_13305,N_13341);
or U13542 (N_13542,N_13347,N_13447);
or U13543 (N_13543,N_13406,N_13482);
or U13544 (N_13544,N_13292,N_13337);
and U13545 (N_13545,N_13254,N_13473);
or U13546 (N_13546,N_13331,N_13332);
and U13547 (N_13547,N_13316,N_13397);
nor U13548 (N_13548,N_13256,N_13329);
and U13549 (N_13549,N_13293,N_13272);
or U13550 (N_13550,N_13296,N_13476);
nor U13551 (N_13551,N_13428,N_13365);
and U13552 (N_13552,N_13477,N_13346);
or U13553 (N_13553,N_13424,N_13449);
and U13554 (N_13554,N_13464,N_13330);
or U13555 (N_13555,N_13466,N_13499);
and U13556 (N_13556,N_13422,N_13282);
nor U13557 (N_13557,N_13334,N_13437);
nand U13558 (N_13558,N_13281,N_13290);
or U13559 (N_13559,N_13438,N_13380);
nor U13560 (N_13560,N_13435,N_13259);
nor U13561 (N_13561,N_13263,N_13415);
nand U13562 (N_13562,N_13471,N_13423);
or U13563 (N_13563,N_13363,N_13400);
and U13564 (N_13564,N_13356,N_13462);
or U13565 (N_13565,N_13352,N_13373);
or U13566 (N_13566,N_13478,N_13265);
nor U13567 (N_13567,N_13324,N_13407);
nand U13568 (N_13568,N_13368,N_13308);
nand U13569 (N_13569,N_13325,N_13456);
nand U13570 (N_13570,N_13258,N_13317);
nor U13571 (N_13571,N_13351,N_13430);
and U13572 (N_13572,N_13304,N_13250);
nand U13573 (N_13573,N_13262,N_13366);
nor U13574 (N_13574,N_13391,N_13335);
and U13575 (N_13575,N_13490,N_13378);
and U13576 (N_13576,N_13374,N_13387);
or U13577 (N_13577,N_13448,N_13307);
or U13578 (N_13578,N_13429,N_13385);
xnor U13579 (N_13579,N_13382,N_13375);
xor U13580 (N_13580,N_13465,N_13383);
nor U13581 (N_13581,N_13372,N_13459);
xor U13582 (N_13582,N_13291,N_13411);
xnor U13583 (N_13583,N_13494,N_13255);
or U13584 (N_13584,N_13328,N_13492);
nand U13585 (N_13585,N_13458,N_13445);
nand U13586 (N_13586,N_13451,N_13470);
nand U13587 (N_13587,N_13417,N_13315);
nand U13588 (N_13588,N_13360,N_13289);
nor U13589 (N_13589,N_13302,N_13354);
xnor U13590 (N_13590,N_13443,N_13485);
xor U13591 (N_13591,N_13427,N_13342);
nor U13592 (N_13592,N_13468,N_13436);
or U13593 (N_13593,N_13357,N_13489);
nor U13594 (N_13594,N_13299,N_13312);
nand U13595 (N_13595,N_13460,N_13283);
xnor U13596 (N_13596,N_13393,N_13396);
or U13597 (N_13597,N_13267,N_13394);
nand U13598 (N_13598,N_13426,N_13496);
and U13599 (N_13599,N_13453,N_13484);
xnor U13600 (N_13600,N_13294,N_13350);
nand U13601 (N_13601,N_13386,N_13420);
xnor U13602 (N_13602,N_13273,N_13421);
nor U13603 (N_13603,N_13455,N_13377);
xnor U13604 (N_13604,N_13338,N_13412);
or U13605 (N_13605,N_13339,N_13300);
or U13606 (N_13606,N_13409,N_13253);
or U13607 (N_13607,N_13416,N_13318);
nor U13608 (N_13608,N_13480,N_13413);
xor U13609 (N_13609,N_13348,N_13389);
xor U13610 (N_13610,N_13454,N_13322);
nor U13611 (N_13611,N_13497,N_13495);
xor U13612 (N_13612,N_13261,N_13370);
and U13613 (N_13613,N_13414,N_13336);
nand U13614 (N_13614,N_13286,N_13358);
nor U13615 (N_13615,N_13488,N_13376);
xor U13616 (N_13616,N_13295,N_13491);
nand U13617 (N_13617,N_13353,N_13418);
nand U13618 (N_13618,N_13479,N_13369);
xnor U13619 (N_13619,N_13381,N_13431);
nor U13620 (N_13620,N_13309,N_13285);
and U13621 (N_13621,N_13301,N_13481);
or U13622 (N_13622,N_13472,N_13364);
nor U13623 (N_13623,N_13277,N_13474);
nand U13624 (N_13624,N_13384,N_13279);
xor U13625 (N_13625,N_13307,N_13375);
xor U13626 (N_13626,N_13396,N_13272);
xor U13627 (N_13627,N_13308,N_13409);
or U13628 (N_13628,N_13475,N_13398);
nor U13629 (N_13629,N_13471,N_13459);
and U13630 (N_13630,N_13322,N_13363);
nand U13631 (N_13631,N_13323,N_13388);
and U13632 (N_13632,N_13277,N_13302);
and U13633 (N_13633,N_13459,N_13437);
xnor U13634 (N_13634,N_13256,N_13343);
or U13635 (N_13635,N_13352,N_13403);
nand U13636 (N_13636,N_13387,N_13351);
xor U13637 (N_13637,N_13465,N_13380);
or U13638 (N_13638,N_13411,N_13268);
and U13639 (N_13639,N_13289,N_13373);
xnor U13640 (N_13640,N_13285,N_13259);
or U13641 (N_13641,N_13460,N_13338);
nand U13642 (N_13642,N_13315,N_13346);
and U13643 (N_13643,N_13297,N_13415);
or U13644 (N_13644,N_13436,N_13308);
or U13645 (N_13645,N_13261,N_13310);
xor U13646 (N_13646,N_13410,N_13324);
xor U13647 (N_13647,N_13313,N_13331);
nand U13648 (N_13648,N_13284,N_13299);
nand U13649 (N_13649,N_13253,N_13455);
and U13650 (N_13650,N_13345,N_13307);
nand U13651 (N_13651,N_13281,N_13253);
or U13652 (N_13652,N_13250,N_13349);
nor U13653 (N_13653,N_13403,N_13336);
nand U13654 (N_13654,N_13383,N_13269);
or U13655 (N_13655,N_13279,N_13250);
xnor U13656 (N_13656,N_13296,N_13256);
nor U13657 (N_13657,N_13304,N_13410);
nand U13658 (N_13658,N_13303,N_13429);
xor U13659 (N_13659,N_13464,N_13385);
and U13660 (N_13660,N_13362,N_13377);
nand U13661 (N_13661,N_13282,N_13319);
or U13662 (N_13662,N_13330,N_13436);
or U13663 (N_13663,N_13419,N_13270);
or U13664 (N_13664,N_13438,N_13487);
xnor U13665 (N_13665,N_13313,N_13452);
xor U13666 (N_13666,N_13395,N_13333);
and U13667 (N_13667,N_13485,N_13392);
xor U13668 (N_13668,N_13487,N_13485);
nor U13669 (N_13669,N_13434,N_13415);
xor U13670 (N_13670,N_13434,N_13443);
nand U13671 (N_13671,N_13263,N_13446);
xnor U13672 (N_13672,N_13423,N_13452);
nor U13673 (N_13673,N_13436,N_13367);
and U13674 (N_13674,N_13367,N_13393);
nand U13675 (N_13675,N_13387,N_13280);
or U13676 (N_13676,N_13261,N_13356);
and U13677 (N_13677,N_13458,N_13455);
and U13678 (N_13678,N_13383,N_13313);
nand U13679 (N_13679,N_13461,N_13462);
or U13680 (N_13680,N_13353,N_13346);
nor U13681 (N_13681,N_13285,N_13436);
and U13682 (N_13682,N_13471,N_13453);
or U13683 (N_13683,N_13370,N_13278);
or U13684 (N_13684,N_13391,N_13484);
xnor U13685 (N_13685,N_13282,N_13393);
and U13686 (N_13686,N_13414,N_13388);
nor U13687 (N_13687,N_13325,N_13321);
and U13688 (N_13688,N_13279,N_13493);
nor U13689 (N_13689,N_13261,N_13305);
or U13690 (N_13690,N_13403,N_13317);
nor U13691 (N_13691,N_13494,N_13282);
and U13692 (N_13692,N_13324,N_13276);
nor U13693 (N_13693,N_13288,N_13420);
and U13694 (N_13694,N_13388,N_13333);
xor U13695 (N_13695,N_13464,N_13303);
xor U13696 (N_13696,N_13294,N_13470);
xnor U13697 (N_13697,N_13298,N_13297);
nor U13698 (N_13698,N_13316,N_13314);
nand U13699 (N_13699,N_13466,N_13457);
nand U13700 (N_13700,N_13360,N_13335);
nand U13701 (N_13701,N_13331,N_13464);
nor U13702 (N_13702,N_13466,N_13384);
xnor U13703 (N_13703,N_13492,N_13414);
nor U13704 (N_13704,N_13392,N_13448);
nand U13705 (N_13705,N_13274,N_13386);
nand U13706 (N_13706,N_13403,N_13385);
nor U13707 (N_13707,N_13386,N_13487);
and U13708 (N_13708,N_13498,N_13433);
or U13709 (N_13709,N_13383,N_13444);
or U13710 (N_13710,N_13331,N_13351);
nor U13711 (N_13711,N_13320,N_13309);
and U13712 (N_13712,N_13391,N_13425);
and U13713 (N_13713,N_13284,N_13270);
xnor U13714 (N_13714,N_13490,N_13359);
nor U13715 (N_13715,N_13399,N_13390);
nand U13716 (N_13716,N_13306,N_13456);
or U13717 (N_13717,N_13331,N_13446);
xor U13718 (N_13718,N_13498,N_13267);
nor U13719 (N_13719,N_13347,N_13316);
xor U13720 (N_13720,N_13304,N_13408);
nand U13721 (N_13721,N_13492,N_13375);
and U13722 (N_13722,N_13342,N_13328);
xor U13723 (N_13723,N_13462,N_13445);
xor U13724 (N_13724,N_13321,N_13267);
xor U13725 (N_13725,N_13313,N_13299);
nand U13726 (N_13726,N_13280,N_13407);
nand U13727 (N_13727,N_13304,N_13482);
nor U13728 (N_13728,N_13270,N_13471);
and U13729 (N_13729,N_13274,N_13401);
or U13730 (N_13730,N_13415,N_13404);
xor U13731 (N_13731,N_13307,N_13351);
xnor U13732 (N_13732,N_13260,N_13353);
xor U13733 (N_13733,N_13373,N_13366);
and U13734 (N_13734,N_13369,N_13474);
xnor U13735 (N_13735,N_13468,N_13256);
and U13736 (N_13736,N_13318,N_13412);
xor U13737 (N_13737,N_13376,N_13454);
nor U13738 (N_13738,N_13444,N_13427);
xor U13739 (N_13739,N_13300,N_13434);
nand U13740 (N_13740,N_13408,N_13257);
xnor U13741 (N_13741,N_13428,N_13482);
or U13742 (N_13742,N_13474,N_13366);
xnor U13743 (N_13743,N_13396,N_13410);
nand U13744 (N_13744,N_13263,N_13305);
and U13745 (N_13745,N_13400,N_13402);
and U13746 (N_13746,N_13361,N_13403);
xor U13747 (N_13747,N_13305,N_13478);
and U13748 (N_13748,N_13481,N_13308);
xnor U13749 (N_13749,N_13318,N_13252);
and U13750 (N_13750,N_13632,N_13601);
or U13751 (N_13751,N_13722,N_13688);
nand U13752 (N_13752,N_13524,N_13686);
nor U13753 (N_13753,N_13531,N_13642);
or U13754 (N_13754,N_13626,N_13634);
nand U13755 (N_13755,N_13578,N_13528);
nor U13756 (N_13756,N_13682,N_13542);
and U13757 (N_13757,N_13681,N_13523);
nor U13758 (N_13758,N_13639,N_13584);
nand U13759 (N_13759,N_13699,N_13662);
nor U13760 (N_13760,N_13705,N_13532);
and U13761 (N_13761,N_13510,N_13549);
and U13762 (N_13762,N_13514,N_13679);
nand U13763 (N_13763,N_13534,N_13719);
xnor U13764 (N_13764,N_13627,N_13697);
or U13765 (N_13765,N_13658,N_13690);
nand U13766 (N_13766,N_13741,N_13515);
xnor U13767 (N_13767,N_13502,N_13712);
or U13768 (N_13768,N_13565,N_13620);
nor U13769 (N_13769,N_13689,N_13605);
or U13770 (N_13770,N_13715,N_13596);
xor U13771 (N_13771,N_13587,N_13656);
or U13772 (N_13772,N_13527,N_13543);
or U13773 (N_13773,N_13691,N_13588);
or U13774 (N_13774,N_13695,N_13635);
nor U13775 (N_13775,N_13659,N_13551);
xnor U13776 (N_13776,N_13538,N_13641);
or U13777 (N_13777,N_13663,N_13591);
xor U13778 (N_13778,N_13667,N_13582);
xor U13779 (N_13779,N_13700,N_13537);
and U13780 (N_13780,N_13513,N_13579);
and U13781 (N_13781,N_13671,N_13678);
nand U13782 (N_13782,N_13604,N_13598);
nand U13783 (N_13783,N_13512,N_13501);
xor U13784 (N_13784,N_13736,N_13676);
and U13785 (N_13785,N_13693,N_13580);
or U13786 (N_13786,N_13516,N_13713);
or U13787 (N_13787,N_13680,N_13717);
or U13788 (N_13788,N_13692,N_13685);
xor U13789 (N_13789,N_13526,N_13603);
nor U13790 (N_13790,N_13555,N_13743);
or U13791 (N_13791,N_13657,N_13540);
nor U13792 (N_13792,N_13638,N_13651);
nor U13793 (N_13793,N_13599,N_13730);
or U13794 (N_13794,N_13535,N_13547);
and U13795 (N_13795,N_13594,N_13572);
xor U13796 (N_13796,N_13684,N_13511);
or U13797 (N_13797,N_13552,N_13640);
nand U13798 (N_13798,N_13560,N_13665);
and U13799 (N_13799,N_13623,N_13561);
or U13800 (N_13800,N_13602,N_13728);
nand U13801 (N_13801,N_13586,N_13739);
nand U13802 (N_13802,N_13747,N_13738);
or U13803 (N_13803,N_13742,N_13731);
and U13804 (N_13804,N_13711,N_13646);
nor U13805 (N_13805,N_13624,N_13725);
nand U13806 (N_13806,N_13718,N_13675);
nand U13807 (N_13807,N_13734,N_13593);
or U13808 (N_13808,N_13727,N_13687);
and U13809 (N_13809,N_13619,N_13517);
nor U13810 (N_13810,N_13648,N_13546);
or U13811 (N_13811,N_13660,N_13649);
nor U13812 (N_13812,N_13589,N_13563);
and U13813 (N_13813,N_13608,N_13597);
nor U13814 (N_13814,N_13655,N_13530);
and U13815 (N_13815,N_13557,N_13567);
or U13816 (N_13816,N_13669,N_13503);
nand U13817 (N_13817,N_13569,N_13744);
and U13818 (N_13818,N_13606,N_13653);
or U13819 (N_13819,N_13545,N_13698);
and U13820 (N_13820,N_13643,N_13518);
xor U13821 (N_13821,N_13745,N_13637);
nor U13822 (N_13822,N_13702,N_13574);
nor U13823 (N_13823,N_13664,N_13625);
or U13824 (N_13824,N_13612,N_13726);
or U13825 (N_13825,N_13670,N_13600);
nor U13826 (N_13826,N_13696,N_13735);
xnor U13827 (N_13827,N_13721,N_13716);
nand U13828 (N_13828,N_13708,N_13611);
nand U13829 (N_13829,N_13720,N_13674);
nor U13830 (N_13830,N_13581,N_13654);
nand U13831 (N_13831,N_13729,N_13577);
or U13832 (N_13832,N_13746,N_13616);
nor U13833 (N_13833,N_13585,N_13628);
nand U13834 (N_13834,N_13500,N_13749);
nor U13835 (N_13835,N_13519,N_13607);
or U13836 (N_13836,N_13701,N_13710);
xnor U13837 (N_13837,N_13590,N_13553);
nor U13838 (N_13838,N_13615,N_13522);
nand U13839 (N_13839,N_13703,N_13748);
xnor U13840 (N_13840,N_13570,N_13737);
xor U13841 (N_13841,N_13507,N_13521);
and U13842 (N_13842,N_13566,N_13568);
nand U13843 (N_13843,N_13592,N_13617);
nor U13844 (N_13844,N_13723,N_13505);
and U13845 (N_13845,N_13571,N_13652);
or U13846 (N_13846,N_13683,N_13694);
and U13847 (N_13847,N_13707,N_13595);
or U13848 (N_13848,N_13550,N_13520);
nand U13849 (N_13849,N_13621,N_13554);
nand U13850 (N_13850,N_13610,N_13508);
nand U13851 (N_13851,N_13645,N_13740);
and U13852 (N_13852,N_13525,N_13509);
nor U13853 (N_13853,N_13544,N_13614);
nand U13854 (N_13854,N_13636,N_13558);
or U13855 (N_13855,N_13541,N_13673);
or U13856 (N_13856,N_13644,N_13733);
and U13857 (N_13857,N_13564,N_13622);
or U13858 (N_13858,N_13633,N_13706);
nor U13859 (N_13859,N_13539,N_13573);
and U13860 (N_13860,N_13732,N_13672);
or U13861 (N_13861,N_13668,N_13576);
nor U13862 (N_13862,N_13548,N_13562);
or U13863 (N_13863,N_13629,N_13724);
or U13864 (N_13864,N_13609,N_13704);
nor U13865 (N_13865,N_13618,N_13661);
nand U13866 (N_13866,N_13666,N_13583);
and U13867 (N_13867,N_13556,N_13613);
xor U13868 (N_13868,N_13559,N_13647);
xnor U13869 (N_13869,N_13506,N_13536);
and U13870 (N_13870,N_13630,N_13575);
xnor U13871 (N_13871,N_13677,N_13529);
nor U13872 (N_13872,N_13533,N_13709);
nor U13873 (N_13873,N_13650,N_13504);
or U13874 (N_13874,N_13631,N_13714);
xor U13875 (N_13875,N_13699,N_13726);
xor U13876 (N_13876,N_13573,N_13630);
xor U13877 (N_13877,N_13664,N_13606);
nor U13878 (N_13878,N_13579,N_13619);
nand U13879 (N_13879,N_13598,N_13642);
xnor U13880 (N_13880,N_13533,N_13577);
nand U13881 (N_13881,N_13551,N_13518);
or U13882 (N_13882,N_13514,N_13593);
and U13883 (N_13883,N_13655,N_13701);
or U13884 (N_13884,N_13574,N_13620);
nor U13885 (N_13885,N_13613,N_13514);
xor U13886 (N_13886,N_13617,N_13519);
nor U13887 (N_13887,N_13719,N_13614);
or U13888 (N_13888,N_13556,N_13696);
nor U13889 (N_13889,N_13671,N_13598);
and U13890 (N_13890,N_13697,N_13502);
nand U13891 (N_13891,N_13573,N_13619);
nand U13892 (N_13892,N_13676,N_13738);
nor U13893 (N_13893,N_13503,N_13543);
nand U13894 (N_13894,N_13646,N_13552);
or U13895 (N_13895,N_13659,N_13685);
nor U13896 (N_13896,N_13541,N_13679);
and U13897 (N_13897,N_13598,N_13709);
or U13898 (N_13898,N_13568,N_13608);
nor U13899 (N_13899,N_13658,N_13637);
nand U13900 (N_13900,N_13536,N_13670);
nor U13901 (N_13901,N_13701,N_13554);
nand U13902 (N_13902,N_13748,N_13712);
or U13903 (N_13903,N_13500,N_13591);
and U13904 (N_13904,N_13707,N_13637);
nor U13905 (N_13905,N_13714,N_13609);
or U13906 (N_13906,N_13561,N_13648);
or U13907 (N_13907,N_13683,N_13543);
nor U13908 (N_13908,N_13606,N_13582);
nor U13909 (N_13909,N_13678,N_13701);
or U13910 (N_13910,N_13564,N_13662);
and U13911 (N_13911,N_13647,N_13573);
nor U13912 (N_13912,N_13555,N_13666);
and U13913 (N_13913,N_13598,N_13555);
xnor U13914 (N_13914,N_13735,N_13561);
or U13915 (N_13915,N_13742,N_13513);
or U13916 (N_13916,N_13503,N_13625);
and U13917 (N_13917,N_13614,N_13532);
and U13918 (N_13918,N_13632,N_13721);
xor U13919 (N_13919,N_13550,N_13724);
xnor U13920 (N_13920,N_13632,N_13635);
nand U13921 (N_13921,N_13524,N_13644);
xnor U13922 (N_13922,N_13545,N_13593);
xor U13923 (N_13923,N_13627,N_13626);
and U13924 (N_13924,N_13637,N_13569);
xor U13925 (N_13925,N_13702,N_13593);
nand U13926 (N_13926,N_13539,N_13611);
xor U13927 (N_13927,N_13546,N_13683);
and U13928 (N_13928,N_13553,N_13620);
nand U13929 (N_13929,N_13638,N_13527);
nor U13930 (N_13930,N_13504,N_13573);
nand U13931 (N_13931,N_13672,N_13521);
xor U13932 (N_13932,N_13537,N_13531);
nand U13933 (N_13933,N_13688,N_13501);
nand U13934 (N_13934,N_13528,N_13747);
or U13935 (N_13935,N_13563,N_13556);
and U13936 (N_13936,N_13661,N_13729);
nor U13937 (N_13937,N_13725,N_13545);
and U13938 (N_13938,N_13673,N_13566);
nor U13939 (N_13939,N_13604,N_13681);
and U13940 (N_13940,N_13595,N_13747);
or U13941 (N_13941,N_13551,N_13582);
xnor U13942 (N_13942,N_13560,N_13545);
nor U13943 (N_13943,N_13732,N_13668);
xnor U13944 (N_13944,N_13602,N_13650);
xnor U13945 (N_13945,N_13518,N_13620);
or U13946 (N_13946,N_13646,N_13632);
nor U13947 (N_13947,N_13593,N_13510);
or U13948 (N_13948,N_13640,N_13606);
nor U13949 (N_13949,N_13509,N_13516);
or U13950 (N_13950,N_13720,N_13721);
nor U13951 (N_13951,N_13605,N_13741);
nor U13952 (N_13952,N_13547,N_13653);
or U13953 (N_13953,N_13650,N_13557);
and U13954 (N_13954,N_13575,N_13733);
and U13955 (N_13955,N_13563,N_13718);
xnor U13956 (N_13956,N_13557,N_13520);
and U13957 (N_13957,N_13561,N_13674);
or U13958 (N_13958,N_13546,N_13684);
or U13959 (N_13959,N_13620,N_13506);
or U13960 (N_13960,N_13588,N_13634);
nor U13961 (N_13961,N_13543,N_13676);
and U13962 (N_13962,N_13552,N_13557);
xor U13963 (N_13963,N_13615,N_13711);
and U13964 (N_13964,N_13627,N_13568);
xnor U13965 (N_13965,N_13632,N_13675);
and U13966 (N_13966,N_13631,N_13691);
and U13967 (N_13967,N_13549,N_13602);
nor U13968 (N_13968,N_13668,N_13549);
nor U13969 (N_13969,N_13585,N_13575);
and U13970 (N_13970,N_13657,N_13573);
nand U13971 (N_13971,N_13685,N_13637);
xnor U13972 (N_13972,N_13747,N_13630);
nor U13973 (N_13973,N_13645,N_13643);
and U13974 (N_13974,N_13669,N_13592);
xor U13975 (N_13975,N_13564,N_13682);
or U13976 (N_13976,N_13709,N_13728);
nor U13977 (N_13977,N_13584,N_13548);
nor U13978 (N_13978,N_13642,N_13744);
or U13979 (N_13979,N_13573,N_13701);
and U13980 (N_13980,N_13718,N_13600);
nand U13981 (N_13981,N_13713,N_13711);
nand U13982 (N_13982,N_13554,N_13684);
nand U13983 (N_13983,N_13545,N_13723);
or U13984 (N_13984,N_13664,N_13547);
or U13985 (N_13985,N_13589,N_13705);
nand U13986 (N_13986,N_13710,N_13630);
and U13987 (N_13987,N_13586,N_13609);
xor U13988 (N_13988,N_13731,N_13608);
nand U13989 (N_13989,N_13590,N_13510);
or U13990 (N_13990,N_13608,N_13707);
and U13991 (N_13991,N_13601,N_13631);
nor U13992 (N_13992,N_13552,N_13689);
xor U13993 (N_13993,N_13561,N_13652);
nand U13994 (N_13994,N_13707,N_13516);
or U13995 (N_13995,N_13551,N_13605);
or U13996 (N_13996,N_13588,N_13663);
nor U13997 (N_13997,N_13717,N_13638);
nand U13998 (N_13998,N_13564,N_13687);
xor U13999 (N_13999,N_13649,N_13708);
or U14000 (N_14000,N_13770,N_13951);
and U14001 (N_14001,N_13983,N_13782);
or U14002 (N_14002,N_13979,N_13808);
xnor U14003 (N_14003,N_13755,N_13781);
nor U14004 (N_14004,N_13860,N_13812);
nor U14005 (N_14005,N_13879,N_13785);
xnor U14006 (N_14006,N_13955,N_13882);
nand U14007 (N_14007,N_13997,N_13884);
or U14008 (N_14008,N_13995,N_13837);
or U14009 (N_14009,N_13801,N_13934);
nand U14010 (N_14010,N_13780,N_13810);
nand U14011 (N_14011,N_13757,N_13965);
nor U14012 (N_14012,N_13855,N_13805);
nor U14013 (N_14013,N_13830,N_13952);
or U14014 (N_14014,N_13849,N_13896);
and U14015 (N_14015,N_13799,N_13767);
xor U14016 (N_14016,N_13838,N_13821);
and U14017 (N_14017,N_13897,N_13829);
or U14018 (N_14018,N_13888,N_13859);
and U14019 (N_14019,N_13998,N_13809);
and U14020 (N_14020,N_13779,N_13921);
and U14021 (N_14021,N_13793,N_13803);
xor U14022 (N_14022,N_13929,N_13914);
nor U14023 (N_14023,N_13777,N_13958);
xnor U14024 (N_14024,N_13906,N_13806);
nand U14025 (N_14025,N_13794,N_13786);
and U14026 (N_14026,N_13971,N_13970);
xor U14027 (N_14027,N_13993,N_13950);
and U14028 (N_14028,N_13870,N_13769);
or U14029 (N_14029,N_13807,N_13956);
nand U14030 (N_14030,N_13824,N_13845);
nor U14031 (N_14031,N_13788,N_13828);
or U14032 (N_14032,N_13834,N_13835);
xor U14033 (N_14033,N_13823,N_13947);
nand U14034 (N_14034,N_13865,N_13848);
nor U14035 (N_14035,N_13917,N_13899);
nor U14036 (N_14036,N_13844,N_13945);
nand U14037 (N_14037,N_13866,N_13831);
nor U14038 (N_14038,N_13832,N_13762);
and U14039 (N_14039,N_13774,N_13992);
nor U14040 (N_14040,N_13861,N_13802);
nand U14041 (N_14041,N_13811,N_13927);
nor U14042 (N_14042,N_13939,N_13797);
or U14043 (N_14043,N_13880,N_13900);
nor U14044 (N_14044,N_13854,N_13969);
nor U14045 (N_14045,N_13911,N_13820);
nand U14046 (N_14046,N_13907,N_13874);
xnor U14047 (N_14047,N_13846,N_13887);
nor U14048 (N_14048,N_13856,N_13964);
and U14049 (N_14049,N_13814,N_13852);
nor U14050 (N_14050,N_13875,N_13940);
nor U14051 (N_14051,N_13954,N_13763);
and U14052 (N_14052,N_13825,N_13949);
and U14053 (N_14053,N_13923,N_13822);
nor U14054 (N_14054,N_13817,N_13815);
and U14055 (N_14055,N_13905,N_13759);
or U14056 (N_14056,N_13885,N_13839);
and U14057 (N_14057,N_13862,N_13919);
and U14058 (N_14058,N_13932,N_13761);
xnor U14059 (N_14059,N_13873,N_13858);
or U14060 (N_14060,N_13959,N_13991);
nor U14061 (N_14061,N_13904,N_13864);
nor U14062 (N_14062,N_13922,N_13756);
nand U14063 (N_14063,N_13981,N_13894);
nand U14064 (N_14064,N_13840,N_13760);
nor U14065 (N_14065,N_13913,N_13843);
xnor U14066 (N_14066,N_13942,N_13912);
xnor U14067 (N_14067,N_13881,N_13868);
nor U14068 (N_14068,N_13957,N_13863);
nor U14069 (N_14069,N_13902,N_13903);
or U14070 (N_14070,N_13754,N_13961);
nor U14071 (N_14071,N_13893,N_13765);
nor U14072 (N_14072,N_13768,N_13982);
nor U14073 (N_14073,N_13851,N_13918);
xnor U14074 (N_14074,N_13924,N_13909);
or U14075 (N_14075,N_13999,N_13751);
xnor U14076 (N_14076,N_13818,N_13773);
nor U14077 (N_14077,N_13977,N_13928);
or U14078 (N_14078,N_13766,N_13816);
nand U14079 (N_14079,N_13842,N_13935);
nor U14080 (N_14080,N_13791,N_13867);
nor U14081 (N_14081,N_13938,N_13968);
or U14082 (N_14082,N_13790,N_13976);
xor U14083 (N_14083,N_13853,N_13784);
xnor U14084 (N_14084,N_13776,N_13895);
nor U14085 (N_14085,N_13871,N_13850);
or U14086 (N_14086,N_13892,N_13994);
nor U14087 (N_14087,N_13778,N_13944);
and U14088 (N_14088,N_13847,N_13869);
or U14089 (N_14089,N_13986,N_13985);
and U14090 (N_14090,N_13877,N_13883);
and U14091 (N_14091,N_13787,N_13987);
and U14092 (N_14092,N_13978,N_13876);
and U14093 (N_14093,N_13975,N_13931);
nor U14094 (N_14094,N_13750,N_13920);
xnor U14095 (N_14095,N_13990,N_13819);
or U14096 (N_14096,N_13795,N_13967);
xor U14097 (N_14097,N_13836,N_13775);
or U14098 (N_14098,N_13890,N_13953);
and U14099 (N_14099,N_13827,N_13963);
nor U14100 (N_14100,N_13941,N_13792);
nor U14101 (N_14101,N_13915,N_13783);
or U14102 (N_14102,N_13796,N_13984);
xor U14103 (N_14103,N_13800,N_13996);
or U14104 (N_14104,N_13798,N_13908);
nand U14105 (N_14105,N_13925,N_13753);
nor U14106 (N_14106,N_13764,N_13933);
nand U14107 (N_14107,N_13841,N_13813);
and U14108 (N_14108,N_13988,N_13960);
and U14109 (N_14109,N_13889,N_13930);
nor U14110 (N_14110,N_13962,N_13857);
xnor U14111 (N_14111,N_13946,N_13804);
and U14112 (N_14112,N_13826,N_13789);
xnor U14113 (N_14113,N_13872,N_13937);
or U14114 (N_14114,N_13771,N_13916);
or U14115 (N_14115,N_13926,N_13752);
xnor U14116 (N_14116,N_13878,N_13772);
nand U14117 (N_14117,N_13948,N_13980);
and U14118 (N_14118,N_13898,N_13891);
and U14119 (N_14119,N_13910,N_13972);
or U14120 (N_14120,N_13833,N_13901);
nand U14121 (N_14121,N_13966,N_13974);
xnor U14122 (N_14122,N_13943,N_13989);
and U14123 (N_14123,N_13758,N_13973);
xor U14124 (N_14124,N_13936,N_13886);
nand U14125 (N_14125,N_13986,N_13863);
and U14126 (N_14126,N_13827,N_13760);
or U14127 (N_14127,N_13959,N_13946);
nor U14128 (N_14128,N_13897,N_13997);
nand U14129 (N_14129,N_13932,N_13865);
or U14130 (N_14130,N_13909,N_13795);
nand U14131 (N_14131,N_13913,N_13902);
nor U14132 (N_14132,N_13873,N_13963);
nor U14133 (N_14133,N_13760,N_13868);
xnor U14134 (N_14134,N_13768,N_13945);
nand U14135 (N_14135,N_13841,N_13979);
xor U14136 (N_14136,N_13924,N_13969);
nand U14137 (N_14137,N_13909,N_13753);
and U14138 (N_14138,N_13936,N_13871);
or U14139 (N_14139,N_13972,N_13839);
xnor U14140 (N_14140,N_13932,N_13995);
nand U14141 (N_14141,N_13865,N_13958);
and U14142 (N_14142,N_13916,N_13828);
or U14143 (N_14143,N_13955,N_13847);
xor U14144 (N_14144,N_13806,N_13856);
and U14145 (N_14145,N_13948,N_13996);
or U14146 (N_14146,N_13791,N_13806);
xor U14147 (N_14147,N_13756,N_13785);
nand U14148 (N_14148,N_13800,N_13976);
nor U14149 (N_14149,N_13786,N_13765);
nand U14150 (N_14150,N_13828,N_13914);
and U14151 (N_14151,N_13925,N_13835);
nand U14152 (N_14152,N_13944,N_13919);
and U14153 (N_14153,N_13925,N_13983);
xor U14154 (N_14154,N_13891,N_13861);
and U14155 (N_14155,N_13846,N_13914);
nor U14156 (N_14156,N_13933,N_13984);
xnor U14157 (N_14157,N_13847,N_13827);
xnor U14158 (N_14158,N_13895,N_13889);
or U14159 (N_14159,N_13819,N_13971);
or U14160 (N_14160,N_13847,N_13794);
nand U14161 (N_14161,N_13983,N_13778);
xnor U14162 (N_14162,N_13888,N_13882);
nor U14163 (N_14163,N_13997,N_13906);
nand U14164 (N_14164,N_13870,N_13805);
xnor U14165 (N_14165,N_13790,N_13936);
and U14166 (N_14166,N_13972,N_13954);
xnor U14167 (N_14167,N_13815,N_13890);
nor U14168 (N_14168,N_13766,N_13819);
and U14169 (N_14169,N_13852,N_13998);
nor U14170 (N_14170,N_13817,N_13999);
or U14171 (N_14171,N_13829,N_13813);
or U14172 (N_14172,N_13886,N_13852);
xor U14173 (N_14173,N_13760,N_13932);
xnor U14174 (N_14174,N_13923,N_13836);
nor U14175 (N_14175,N_13779,N_13879);
or U14176 (N_14176,N_13763,N_13875);
or U14177 (N_14177,N_13758,N_13980);
nand U14178 (N_14178,N_13801,N_13992);
xor U14179 (N_14179,N_13893,N_13976);
nor U14180 (N_14180,N_13953,N_13788);
nand U14181 (N_14181,N_13858,N_13989);
or U14182 (N_14182,N_13795,N_13814);
nor U14183 (N_14183,N_13779,N_13791);
nand U14184 (N_14184,N_13908,N_13853);
and U14185 (N_14185,N_13792,N_13940);
or U14186 (N_14186,N_13958,N_13822);
xor U14187 (N_14187,N_13851,N_13869);
nor U14188 (N_14188,N_13842,N_13864);
or U14189 (N_14189,N_13961,N_13879);
xnor U14190 (N_14190,N_13913,N_13924);
nor U14191 (N_14191,N_13842,N_13809);
nor U14192 (N_14192,N_13810,N_13760);
xnor U14193 (N_14193,N_13930,N_13882);
and U14194 (N_14194,N_13969,N_13821);
nand U14195 (N_14195,N_13880,N_13838);
and U14196 (N_14196,N_13883,N_13929);
and U14197 (N_14197,N_13773,N_13894);
nor U14198 (N_14198,N_13903,N_13885);
nor U14199 (N_14199,N_13802,N_13958);
nor U14200 (N_14200,N_13803,N_13837);
nor U14201 (N_14201,N_13973,N_13870);
xor U14202 (N_14202,N_13809,N_13833);
xnor U14203 (N_14203,N_13888,N_13969);
nand U14204 (N_14204,N_13942,N_13859);
xnor U14205 (N_14205,N_13824,N_13976);
nor U14206 (N_14206,N_13900,N_13985);
or U14207 (N_14207,N_13804,N_13797);
nor U14208 (N_14208,N_13790,N_13964);
nor U14209 (N_14209,N_13761,N_13846);
xor U14210 (N_14210,N_13892,N_13914);
nor U14211 (N_14211,N_13990,N_13959);
and U14212 (N_14212,N_13859,N_13782);
nor U14213 (N_14213,N_13913,N_13922);
nand U14214 (N_14214,N_13786,N_13952);
nand U14215 (N_14215,N_13988,N_13790);
xnor U14216 (N_14216,N_13797,N_13887);
nand U14217 (N_14217,N_13838,N_13927);
xor U14218 (N_14218,N_13963,N_13814);
xnor U14219 (N_14219,N_13974,N_13859);
and U14220 (N_14220,N_13968,N_13866);
nor U14221 (N_14221,N_13937,N_13899);
or U14222 (N_14222,N_13914,N_13880);
nor U14223 (N_14223,N_13971,N_13790);
nand U14224 (N_14224,N_13882,N_13813);
nor U14225 (N_14225,N_13844,N_13793);
or U14226 (N_14226,N_13873,N_13985);
and U14227 (N_14227,N_13841,N_13784);
or U14228 (N_14228,N_13876,N_13753);
xnor U14229 (N_14229,N_13937,N_13866);
xor U14230 (N_14230,N_13888,N_13986);
nand U14231 (N_14231,N_13921,N_13808);
nor U14232 (N_14232,N_13777,N_13902);
xnor U14233 (N_14233,N_13772,N_13879);
or U14234 (N_14234,N_13806,N_13809);
nor U14235 (N_14235,N_13765,N_13857);
or U14236 (N_14236,N_13840,N_13893);
or U14237 (N_14237,N_13869,N_13854);
nand U14238 (N_14238,N_13843,N_13762);
nand U14239 (N_14239,N_13894,N_13966);
or U14240 (N_14240,N_13797,N_13832);
xor U14241 (N_14241,N_13971,N_13782);
nand U14242 (N_14242,N_13795,N_13847);
and U14243 (N_14243,N_13857,N_13850);
xnor U14244 (N_14244,N_13936,N_13777);
xor U14245 (N_14245,N_13918,N_13828);
nor U14246 (N_14246,N_13891,N_13801);
and U14247 (N_14247,N_13924,N_13949);
xnor U14248 (N_14248,N_13863,N_13859);
xor U14249 (N_14249,N_13958,N_13783);
and U14250 (N_14250,N_14198,N_14125);
xor U14251 (N_14251,N_14050,N_14011);
nor U14252 (N_14252,N_14237,N_14022);
xnor U14253 (N_14253,N_14194,N_14021);
nand U14254 (N_14254,N_14238,N_14215);
xnor U14255 (N_14255,N_14025,N_14212);
nor U14256 (N_14256,N_14034,N_14063);
nand U14257 (N_14257,N_14110,N_14195);
nand U14258 (N_14258,N_14071,N_14189);
or U14259 (N_14259,N_14039,N_14166);
nand U14260 (N_14260,N_14245,N_14133);
xnor U14261 (N_14261,N_14056,N_14054);
xor U14262 (N_14262,N_14154,N_14134);
and U14263 (N_14263,N_14089,N_14053);
nor U14264 (N_14264,N_14099,N_14144);
xor U14265 (N_14265,N_14219,N_14102);
xnor U14266 (N_14266,N_14159,N_14182);
xnor U14267 (N_14267,N_14140,N_14074);
and U14268 (N_14268,N_14038,N_14059);
or U14269 (N_14269,N_14120,N_14127);
or U14270 (N_14270,N_14139,N_14216);
or U14271 (N_14271,N_14170,N_14206);
or U14272 (N_14272,N_14168,N_14242);
nand U14273 (N_14273,N_14131,N_14181);
and U14274 (N_14274,N_14044,N_14136);
or U14275 (N_14275,N_14001,N_14118);
and U14276 (N_14276,N_14014,N_14183);
or U14277 (N_14277,N_14057,N_14147);
or U14278 (N_14278,N_14041,N_14000);
nor U14279 (N_14279,N_14043,N_14178);
nor U14280 (N_14280,N_14106,N_14151);
and U14281 (N_14281,N_14224,N_14150);
xnor U14282 (N_14282,N_14076,N_14023);
nand U14283 (N_14283,N_14180,N_14213);
nand U14284 (N_14284,N_14163,N_14153);
xor U14285 (N_14285,N_14003,N_14072);
or U14286 (N_14286,N_14184,N_14040);
and U14287 (N_14287,N_14130,N_14008);
nor U14288 (N_14288,N_14239,N_14006);
nand U14289 (N_14289,N_14103,N_14177);
and U14290 (N_14290,N_14094,N_14046);
or U14291 (N_14291,N_14061,N_14217);
xnor U14292 (N_14292,N_14193,N_14160);
nand U14293 (N_14293,N_14049,N_14088);
and U14294 (N_14294,N_14135,N_14109);
nand U14295 (N_14295,N_14176,N_14188);
xnor U14296 (N_14296,N_14079,N_14143);
and U14297 (N_14297,N_14016,N_14027);
nand U14298 (N_14298,N_14197,N_14205);
or U14299 (N_14299,N_14165,N_14155);
nand U14300 (N_14300,N_14062,N_14124);
and U14301 (N_14301,N_14007,N_14248);
nor U14302 (N_14302,N_14161,N_14013);
and U14303 (N_14303,N_14231,N_14164);
xnor U14304 (N_14304,N_14087,N_14029);
nand U14305 (N_14305,N_14080,N_14210);
nor U14306 (N_14306,N_14077,N_14241);
xnor U14307 (N_14307,N_14012,N_14171);
xor U14308 (N_14308,N_14233,N_14209);
and U14309 (N_14309,N_14086,N_14247);
and U14310 (N_14310,N_14146,N_14107);
nand U14311 (N_14311,N_14128,N_14032);
and U14312 (N_14312,N_14031,N_14100);
or U14313 (N_14313,N_14232,N_14112);
xnor U14314 (N_14314,N_14081,N_14185);
and U14315 (N_14315,N_14018,N_14200);
or U14316 (N_14316,N_14226,N_14234);
and U14317 (N_14317,N_14202,N_14048);
nand U14318 (N_14318,N_14036,N_14104);
or U14319 (N_14319,N_14249,N_14052);
xnor U14320 (N_14320,N_14114,N_14098);
and U14321 (N_14321,N_14190,N_14045);
nor U14322 (N_14322,N_14228,N_14169);
nand U14323 (N_14323,N_14019,N_14122);
nor U14324 (N_14324,N_14230,N_14175);
nor U14325 (N_14325,N_14196,N_14204);
or U14326 (N_14326,N_14158,N_14083);
xnor U14327 (N_14327,N_14141,N_14167);
nor U14328 (N_14328,N_14220,N_14117);
xnor U14329 (N_14329,N_14152,N_14187);
xnor U14330 (N_14330,N_14075,N_14101);
or U14331 (N_14331,N_14156,N_14218);
nand U14332 (N_14332,N_14084,N_14119);
nand U14333 (N_14333,N_14108,N_14243);
and U14334 (N_14334,N_14028,N_14010);
or U14335 (N_14335,N_14097,N_14129);
nand U14336 (N_14336,N_14055,N_14223);
xnor U14337 (N_14337,N_14111,N_14191);
nand U14338 (N_14338,N_14020,N_14042);
xor U14339 (N_14339,N_14015,N_14090);
nor U14340 (N_14340,N_14174,N_14142);
nand U14341 (N_14341,N_14069,N_14067);
nor U14342 (N_14342,N_14179,N_14207);
nand U14343 (N_14343,N_14082,N_14236);
and U14344 (N_14344,N_14035,N_14095);
and U14345 (N_14345,N_14145,N_14192);
nor U14346 (N_14346,N_14004,N_14068);
nand U14347 (N_14347,N_14225,N_14246);
or U14348 (N_14348,N_14186,N_14033);
and U14349 (N_14349,N_14024,N_14047);
nand U14350 (N_14350,N_14173,N_14137);
xnor U14351 (N_14351,N_14214,N_14244);
nor U14352 (N_14352,N_14199,N_14064);
or U14353 (N_14353,N_14126,N_14211);
and U14354 (N_14354,N_14037,N_14005);
xnor U14355 (N_14355,N_14093,N_14009);
xor U14356 (N_14356,N_14051,N_14066);
xnor U14357 (N_14357,N_14123,N_14149);
and U14358 (N_14358,N_14065,N_14115);
or U14359 (N_14359,N_14092,N_14132);
or U14360 (N_14360,N_14105,N_14073);
nor U14361 (N_14361,N_14240,N_14070);
or U14362 (N_14362,N_14060,N_14201);
xor U14363 (N_14363,N_14091,N_14116);
nor U14364 (N_14364,N_14229,N_14058);
or U14365 (N_14365,N_14157,N_14030);
nand U14366 (N_14366,N_14121,N_14162);
nor U14367 (N_14367,N_14221,N_14002);
xnor U14368 (N_14368,N_14026,N_14227);
xor U14369 (N_14369,N_14208,N_14017);
xnor U14370 (N_14370,N_14148,N_14085);
nand U14371 (N_14371,N_14203,N_14172);
nor U14372 (N_14372,N_14113,N_14138);
and U14373 (N_14373,N_14235,N_14222);
nor U14374 (N_14374,N_14096,N_14078);
xnor U14375 (N_14375,N_14157,N_14059);
and U14376 (N_14376,N_14194,N_14128);
nor U14377 (N_14377,N_14056,N_14237);
xnor U14378 (N_14378,N_14168,N_14095);
xnor U14379 (N_14379,N_14239,N_14069);
xor U14380 (N_14380,N_14234,N_14211);
nand U14381 (N_14381,N_14083,N_14134);
and U14382 (N_14382,N_14213,N_14097);
and U14383 (N_14383,N_14039,N_14030);
and U14384 (N_14384,N_14167,N_14162);
or U14385 (N_14385,N_14200,N_14129);
nor U14386 (N_14386,N_14014,N_14093);
or U14387 (N_14387,N_14170,N_14005);
nand U14388 (N_14388,N_14192,N_14003);
nor U14389 (N_14389,N_14239,N_14093);
or U14390 (N_14390,N_14150,N_14235);
nand U14391 (N_14391,N_14098,N_14237);
nand U14392 (N_14392,N_14055,N_14102);
xnor U14393 (N_14393,N_14079,N_14043);
or U14394 (N_14394,N_14018,N_14092);
or U14395 (N_14395,N_14150,N_14061);
nor U14396 (N_14396,N_14004,N_14191);
xnor U14397 (N_14397,N_14181,N_14203);
nand U14398 (N_14398,N_14216,N_14026);
and U14399 (N_14399,N_14007,N_14002);
nand U14400 (N_14400,N_14157,N_14208);
or U14401 (N_14401,N_14220,N_14192);
nor U14402 (N_14402,N_14148,N_14034);
nor U14403 (N_14403,N_14176,N_14046);
xnor U14404 (N_14404,N_14080,N_14199);
nand U14405 (N_14405,N_14009,N_14030);
and U14406 (N_14406,N_14084,N_14118);
xor U14407 (N_14407,N_14117,N_14061);
or U14408 (N_14408,N_14027,N_14231);
or U14409 (N_14409,N_14063,N_14050);
xor U14410 (N_14410,N_14201,N_14117);
or U14411 (N_14411,N_14207,N_14177);
and U14412 (N_14412,N_14227,N_14085);
and U14413 (N_14413,N_14214,N_14109);
nand U14414 (N_14414,N_14229,N_14045);
nor U14415 (N_14415,N_14214,N_14015);
and U14416 (N_14416,N_14018,N_14025);
or U14417 (N_14417,N_14083,N_14229);
xnor U14418 (N_14418,N_14135,N_14150);
or U14419 (N_14419,N_14084,N_14191);
and U14420 (N_14420,N_14204,N_14215);
nand U14421 (N_14421,N_14017,N_14190);
or U14422 (N_14422,N_14035,N_14213);
nor U14423 (N_14423,N_14072,N_14148);
nand U14424 (N_14424,N_14245,N_14033);
nor U14425 (N_14425,N_14116,N_14190);
nand U14426 (N_14426,N_14003,N_14249);
nand U14427 (N_14427,N_14218,N_14200);
and U14428 (N_14428,N_14003,N_14220);
nand U14429 (N_14429,N_14249,N_14203);
and U14430 (N_14430,N_14011,N_14164);
nand U14431 (N_14431,N_14006,N_14124);
or U14432 (N_14432,N_14224,N_14125);
nor U14433 (N_14433,N_14119,N_14011);
xor U14434 (N_14434,N_14175,N_14169);
nor U14435 (N_14435,N_14242,N_14191);
nor U14436 (N_14436,N_14118,N_14169);
and U14437 (N_14437,N_14115,N_14076);
nor U14438 (N_14438,N_14023,N_14009);
nand U14439 (N_14439,N_14197,N_14009);
and U14440 (N_14440,N_14160,N_14205);
nor U14441 (N_14441,N_14178,N_14172);
xor U14442 (N_14442,N_14232,N_14193);
xor U14443 (N_14443,N_14232,N_14192);
nand U14444 (N_14444,N_14156,N_14225);
and U14445 (N_14445,N_14152,N_14110);
xor U14446 (N_14446,N_14182,N_14241);
nand U14447 (N_14447,N_14155,N_14068);
xnor U14448 (N_14448,N_14141,N_14200);
or U14449 (N_14449,N_14068,N_14050);
nand U14450 (N_14450,N_14159,N_14245);
nand U14451 (N_14451,N_14151,N_14007);
nor U14452 (N_14452,N_14243,N_14155);
nand U14453 (N_14453,N_14142,N_14062);
or U14454 (N_14454,N_14201,N_14161);
nand U14455 (N_14455,N_14003,N_14068);
nor U14456 (N_14456,N_14014,N_14236);
nand U14457 (N_14457,N_14089,N_14126);
and U14458 (N_14458,N_14137,N_14157);
nand U14459 (N_14459,N_14174,N_14001);
or U14460 (N_14460,N_14218,N_14033);
nor U14461 (N_14461,N_14236,N_14227);
xnor U14462 (N_14462,N_14094,N_14161);
nor U14463 (N_14463,N_14029,N_14138);
xnor U14464 (N_14464,N_14046,N_14000);
and U14465 (N_14465,N_14053,N_14073);
and U14466 (N_14466,N_14163,N_14074);
or U14467 (N_14467,N_14091,N_14215);
xor U14468 (N_14468,N_14197,N_14047);
nand U14469 (N_14469,N_14121,N_14001);
nor U14470 (N_14470,N_14019,N_14006);
nor U14471 (N_14471,N_14047,N_14233);
nor U14472 (N_14472,N_14169,N_14225);
or U14473 (N_14473,N_14167,N_14103);
and U14474 (N_14474,N_14036,N_14213);
nand U14475 (N_14475,N_14112,N_14061);
nor U14476 (N_14476,N_14173,N_14022);
nor U14477 (N_14477,N_14144,N_14077);
and U14478 (N_14478,N_14141,N_14034);
nand U14479 (N_14479,N_14075,N_14089);
nand U14480 (N_14480,N_14111,N_14011);
nand U14481 (N_14481,N_14131,N_14099);
or U14482 (N_14482,N_14063,N_14017);
nand U14483 (N_14483,N_14246,N_14126);
xor U14484 (N_14484,N_14171,N_14129);
nand U14485 (N_14485,N_14037,N_14043);
or U14486 (N_14486,N_14074,N_14236);
nor U14487 (N_14487,N_14236,N_14015);
nand U14488 (N_14488,N_14125,N_14200);
nand U14489 (N_14489,N_14218,N_14097);
xor U14490 (N_14490,N_14073,N_14087);
or U14491 (N_14491,N_14006,N_14051);
and U14492 (N_14492,N_14242,N_14037);
xnor U14493 (N_14493,N_14130,N_14215);
xnor U14494 (N_14494,N_14129,N_14233);
xor U14495 (N_14495,N_14097,N_14090);
xnor U14496 (N_14496,N_14216,N_14209);
nor U14497 (N_14497,N_14218,N_14194);
xnor U14498 (N_14498,N_14196,N_14049);
nand U14499 (N_14499,N_14125,N_14038);
or U14500 (N_14500,N_14482,N_14400);
or U14501 (N_14501,N_14479,N_14258);
and U14502 (N_14502,N_14309,N_14364);
nor U14503 (N_14503,N_14466,N_14279);
and U14504 (N_14504,N_14444,N_14282);
and U14505 (N_14505,N_14292,N_14326);
xor U14506 (N_14506,N_14461,N_14446);
nor U14507 (N_14507,N_14419,N_14273);
xnor U14508 (N_14508,N_14266,N_14306);
or U14509 (N_14509,N_14412,N_14286);
nand U14510 (N_14510,N_14311,N_14449);
nand U14511 (N_14511,N_14344,N_14434);
nor U14512 (N_14512,N_14381,N_14391);
or U14513 (N_14513,N_14353,N_14437);
nor U14514 (N_14514,N_14432,N_14475);
nand U14515 (N_14515,N_14267,N_14350);
nor U14516 (N_14516,N_14301,N_14483);
nand U14517 (N_14517,N_14293,N_14428);
nand U14518 (N_14518,N_14331,N_14342);
nand U14519 (N_14519,N_14290,N_14407);
nor U14520 (N_14520,N_14442,N_14313);
nand U14521 (N_14521,N_14341,N_14374);
xnor U14522 (N_14522,N_14263,N_14480);
or U14523 (N_14523,N_14300,N_14287);
and U14524 (N_14524,N_14430,N_14276);
xnor U14525 (N_14525,N_14455,N_14278);
nor U14526 (N_14526,N_14431,N_14392);
nor U14527 (N_14527,N_14406,N_14348);
or U14528 (N_14528,N_14369,N_14421);
and U14529 (N_14529,N_14302,N_14396);
xor U14530 (N_14530,N_14425,N_14285);
xor U14531 (N_14531,N_14349,N_14260);
or U14532 (N_14532,N_14498,N_14321);
nor U14533 (N_14533,N_14297,N_14308);
and U14534 (N_14534,N_14433,N_14254);
nand U14535 (N_14535,N_14320,N_14315);
or U14536 (N_14536,N_14394,N_14305);
xnor U14537 (N_14537,N_14274,N_14459);
and U14538 (N_14538,N_14457,N_14351);
nor U14539 (N_14539,N_14271,N_14436);
nor U14540 (N_14540,N_14485,N_14365);
or U14541 (N_14541,N_14423,N_14397);
or U14542 (N_14542,N_14403,N_14484);
nor U14543 (N_14543,N_14384,N_14473);
or U14544 (N_14544,N_14490,N_14337);
nand U14545 (N_14545,N_14332,N_14317);
nand U14546 (N_14546,N_14354,N_14357);
or U14547 (N_14547,N_14343,N_14265);
or U14548 (N_14548,N_14486,N_14335);
nor U14549 (N_14549,N_14383,N_14415);
or U14550 (N_14550,N_14465,N_14316);
nor U14551 (N_14551,N_14451,N_14499);
and U14552 (N_14552,N_14426,N_14359);
and U14553 (N_14553,N_14307,N_14438);
or U14554 (N_14554,N_14356,N_14323);
xor U14555 (N_14555,N_14445,N_14280);
and U14556 (N_14556,N_14358,N_14340);
and U14557 (N_14557,N_14454,N_14288);
or U14558 (N_14558,N_14439,N_14452);
nor U14559 (N_14559,N_14252,N_14324);
nor U14560 (N_14560,N_14330,N_14462);
nand U14561 (N_14561,N_14471,N_14319);
nor U14562 (N_14562,N_14450,N_14399);
and U14563 (N_14563,N_14377,N_14424);
and U14564 (N_14564,N_14289,N_14296);
nand U14565 (N_14565,N_14472,N_14314);
nand U14566 (N_14566,N_14420,N_14338);
nand U14567 (N_14567,N_14382,N_14310);
or U14568 (N_14568,N_14322,N_14492);
nor U14569 (N_14569,N_14496,N_14277);
nor U14570 (N_14570,N_14262,N_14256);
or U14571 (N_14571,N_14489,N_14275);
nand U14572 (N_14572,N_14257,N_14495);
and U14573 (N_14573,N_14367,N_14410);
and U14574 (N_14574,N_14468,N_14390);
and U14575 (N_14575,N_14417,N_14464);
nor U14576 (N_14576,N_14378,N_14270);
xnor U14577 (N_14577,N_14268,N_14360);
and U14578 (N_14578,N_14371,N_14339);
or U14579 (N_14579,N_14398,N_14447);
nand U14580 (N_14580,N_14476,N_14404);
xnor U14581 (N_14581,N_14352,N_14469);
xnor U14582 (N_14582,N_14272,N_14477);
and U14583 (N_14583,N_14251,N_14427);
nand U14584 (N_14584,N_14481,N_14304);
and U14585 (N_14585,N_14418,N_14422);
or U14586 (N_14586,N_14474,N_14453);
nor U14587 (N_14587,N_14488,N_14416);
nand U14588 (N_14588,N_14386,N_14405);
nor U14589 (N_14589,N_14387,N_14456);
or U14590 (N_14590,N_14328,N_14376);
nor U14591 (N_14591,N_14372,N_14366);
or U14592 (N_14592,N_14470,N_14478);
nor U14593 (N_14593,N_14284,N_14346);
nand U14594 (N_14594,N_14291,N_14259);
or U14595 (N_14595,N_14264,N_14361);
or U14596 (N_14596,N_14312,N_14443);
or U14597 (N_14597,N_14298,N_14409);
or U14598 (N_14598,N_14435,N_14333);
xor U14599 (N_14599,N_14295,N_14380);
and U14600 (N_14600,N_14299,N_14318);
xnor U14601 (N_14601,N_14334,N_14497);
and U14602 (N_14602,N_14375,N_14463);
nor U14603 (N_14603,N_14379,N_14325);
and U14604 (N_14604,N_14253,N_14283);
nor U14605 (N_14605,N_14336,N_14458);
xor U14606 (N_14606,N_14460,N_14355);
and U14607 (N_14607,N_14363,N_14368);
or U14608 (N_14608,N_14493,N_14281);
and U14609 (N_14609,N_14401,N_14429);
or U14610 (N_14610,N_14491,N_14441);
or U14611 (N_14611,N_14362,N_14345);
and U14612 (N_14612,N_14347,N_14303);
xor U14613 (N_14613,N_14494,N_14373);
and U14614 (N_14614,N_14294,N_14402);
or U14615 (N_14615,N_14255,N_14487);
or U14616 (N_14616,N_14250,N_14411);
xnor U14617 (N_14617,N_14389,N_14395);
nor U14618 (N_14618,N_14440,N_14385);
xnor U14619 (N_14619,N_14393,N_14467);
and U14620 (N_14620,N_14327,N_14261);
nand U14621 (N_14621,N_14448,N_14388);
or U14622 (N_14622,N_14329,N_14414);
or U14623 (N_14623,N_14413,N_14269);
nor U14624 (N_14624,N_14408,N_14370);
nand U14625 (N_14625,N_14350,N_14414);
nor U14626 (N_14626,N_14371,N_14351);
or U14627 (N_14627,N_14412,N_14468);
and U14628 (N_14628,N_14498,N_14452);
or U14629 (N_14629,N_14399,N_14445);
or U14630 (N_14630,N_14375,N_14250);
nand U14631 (N_14631,N_14327,N_14484);
and U14632 (N_14632,N_14361,N_14467);
and U14633 (N_14633,N_14274,N_14350);
nand U14634 (N_14634,N_14454,N_14464);
or U14635 (N_14635,N_14470,N_14450);
and U14636 (N_14636,N_14311,N_14411);
nand U14637 (N_14637,N_14337,N_14291);
and U14638 (N_14638,N_14289,N_14445);
nor U14639 (N_14639,N_14403,N_14329);
nand U14640 (N_14640,N_14478,N_14336);
nand U14641 (N_14641,N_14405,N_14268);
or U14642 (N_14642,N_14444,N_14347);
or U14643 (N_14643,N_14327,N_14368);
or U14644 (N_14644,N_14270,N_14377);
xnor U14645 (N_14645,N_14452,N_14491);
or U14646 (N_14646,N_14376,N_14436);
xnor U14647 (N_14647,N_14406,N_14378);
nand U14648 (N_14648,N_14425,N_14381);
or U14649 (N_14649,N_14275,N_14391);
or U14650 (N_14650,N_14461,N_14499);
and U14651 (N_14651,N_14311,N_14256);
or U14652 (N_14652,N_14250,N_14339);
nor U14653 (N_14653,N_14289,N_14491);
nor U14654 (N_14654,N_14402,N_14381);
or U14655 (N_14655,N_14301,N_14484);
or U14656 (N_14656,N_14270,N_14468);
nor U14657 (N_14657,N_14495,N_14482);
nand U14658 (N_14658,N_14259,N_14354);
or U14659 (N_14659,N_14353,N_14412);
nand U14660 (N_14660,N_14281,N_14342);
nand U14661 (N_14661,N_14401,N_14423);
xor U14662 (N_14662,N_14422,N_14401);
nor U14663 (N_14663,N_14444,N_14426);
and U14664 (N_14664,N_14448,N_14451);
or U14665 (N_14665,N_14422,N_14497);
nand U14666 (N_14666,N_14438,N_14284);
xor U14667 (N_14667,N_14448,N_14378);
nand U14668 (N_14668,N_14355,N_14325);
xor U14669 (N_14669,N_14410,N_14282);
nor U14670 (N_14670,N_14330,N_14387);
xnor U14671 (N_14671,N_14355,N_14391);
nor U14672 (N_14672,N_14281,N_14339);
and U14673 (N_14673,N_14472,N_14347);
xnor U14674 (N_14674,N_14342,N_14371);
and U14675 (N_14675,N_14250,N_14454);
nor U14676 (N_14676,N_14482,N_14450);
nand U14677 (N_14677,N_14498,N_14361);
nor U14678 (N_14678,N_14365,N_14337);
nor U14679 (N_14679,N_14297,N_14400);
or U14680 (N_14680,N_14277,N_14328);
xnor U14681 (N_14681,N_14252,N_14320);
and U14682 (N_14682,N_14440,N_14404);
or U14683 (N_14683,N_14373,N_14477);
or U14684 (N_14684,N_14482,N_14388);
or U14685 (N_14685,N_14442,N_14408);
nor U14686 (N_14686,N_14478,N_14319);
nand U14687 (N_14687,N_14395,N_14281);
and U14688 (N_14688,N_14467,N_14452);
and U14689 (N_14689,N_14435,N_14392);
and U14690 (N_14690,N_14381,N_14337);
nor U14691 (N_14691,N_14383,N_14253);
nor U14692 (N_14692,N_14345,N_14464);
or U14693 (N_14693,N_14455,N_14393);
and U14694 (N_14694,N_14479,N_14381);
or U14695 (N_14695,N_14466,N_14411);
nand U14696 (N_14696,N_14465,N_14276);
nand U14697 (N_14697,N_14294,N_14421);
and U14698 (N_14698,N_14377,N_14323);
or U14699 (N_14699,N_14257,N_14426);
xnor U14700 (N_14700,N_14321,N_14259);
and U14701 (N_14701,N_14296,N_14443);
nand U14702 (N_14702,N_14286,N_14464);
and U14703 (N_14703,N_14497,N_14474);
or U14704 (N_14704,N_14302,N_14397);
xor U14705 (N_14705,N_14470,N_14418);
nor U14706 (N_14706,N_14499,N_14372);
nor U14707 (N_14707,N_14359,N_14332);
nor U14708 (N_14708,N_14445,N_14389);
or U14709 (N_14709,N_14356,N_14449);
nand U14710 (N_14710,N_14470,N_14277);
and U14711 (N_14711,N_14455,N_14258);
or U14712 (N_14712,N_14251,N_14300);
xnor U14713 (N_14713,N_14316,N_14345);
nand U14714 (N_14714,N_14342,N_14486);
xor U14715 (N_14715,N_14422,N_14326);
xor U14716 (N_14716,N_14483,N_14365);
nor U14717 (N_14717,N_14362,N_14288);
xor U14718 (N_14718,N_14453,N_14343);
xnor U14719 (N_14719,N_14262,N_14495);
nand U14720 (N_14720,N_14250,N_14347);
and U14721 (N_14721,N_14411,N_14318);
nand U14722 (N_14722,N_14400,N_14475);
or U14723 (N_14723,N_14417,N_14337);
xnor U14724 (N_14724,N_14414,N_14305);
nor U14725 (N_14725,N_14489,N_14363);
nand U14726 (N_14726,N_14436,N_14374);
nand U14727 (N_14727,N_14477,N_14320);
and U14728 (N_14728,N_14431,N_14315);
or U14729 (N_14729,N_14368,N_14393);
nor U14730 (N_14730,N_14450,N_14483);
and U14731 (N_14731,N_14339,N_14374);
nor U14732 (N_14732,N_14416,N_14271);
or U14733 (N_14733,N_14256,N_14424);
nor U14734 (N_14734,N_14486,N_14365);
and U14735 (N_14735,N_14298,N_14472);
or U14736 (N_14736,N_14276,N_14323);
and U14737 (N_14737,N_14257,N_14412);
and U14738 (N_14738,N_14260,N_14305);
or U14739 (N_14739,N_14446,N_14386);
nor U14740 (N_14740,N_14490,N_14343);
xor U14741 (N_14741,N_14348,N_14448);
xor U14742 (N_14742,N_14405,N_14282);
xnor U14743 (N_14743,N_14476,N_14490);
and U14744 (N_14744,N_14451,N_14479);
nand U14745 (N_14745,N_14312,N_14407);
or U14746 (N_14746,N_14452,N_14372);
nor U14747 (N_14747,N_14405,N_14438);
or U14748 (N_14748,N_14267,N_14441);
xnor U14749 (N_14749,N_14359,N_14440);
and U14750 (N_14750,N_14610,N_14609);
nor U14751 (N_14751,N_14580,N_14732);
xor U14752 (N_14752,N_14548,N_14730);
nor U14753 (N_14753,N_14574,N_14526);
nor U14754 (N_14754,N_14571,N_14691);
nand U14755 (N_14755,N_14563,N_14601);
and U14756 (N_14756,N_14722,N_14659);
xnor U14757 (N_14757,N_14662,N_14668);
nor U14758 (N_14758,N_14648,N_14694);
or U14759 (N_14759,N_14674,N_14724);
xnor U14760 (N_14760,N_14746,N_14565);
or U14761 (N_14761,N_14581,N_14573);
and U14762 (N_14762,N_14529,N_14602);
or U14763 (N_14763,N_14592,N_14585);
nand U14764 (N_14764,N_14608,N_14567);
xor U14765 (N_14765,N_14530,N_14670);
or U14766 (N_14766,N_14699,N_14544);
nand U14767 (N_14767,N_14644,N_14560);
xor U14768 (N_14768,N_14647,N_14540);
nor U14769 (N_14769,N_14693,N_14531);
xor U14770 (N_14770,N_14742,N_14595);
or U14771 (N_14771,N_14539,N_14711);
nand U14772 (N_14772,N_14717,N_14702);
nand U14773 (N_14773,N_14664,N_14700);
and U14774 (N_14774,N_14527,N_14558);
and U14775 (N_14775,N_14577,N_14709);
or U14776 (N_14776,N_14721,N_14587);
nor U14777 (N_14777,N_14532,N_14626);
and U14778 (N_14778,N_14502,N_14666);
nand U14779 (N_14779,N_14656,N_14625);
nand U14780 (N_14780,N_14658,N_14553);
and U14781 (N_14781,N_14521,N_14590);
and U14782 (N_14782,N_14615,N_14569);
nand U14783 (N_14783,N_14679,N_14593);
and U14784 (N_14784,N_14661,N_14708);
or U14785 (N_14785,N_14634,N_14586);
nand U14786 (N_14786,N_14597,N_14507);
xnor U14787 (N_14787,N_14740,N_14589);
or U14788 (N_14788,N_14554,N_14506);
xor U14789 (N_14789,N_14641,N_14617);
xnor U14790 (N_14790,N_14747,N_14510);
nor U14791 (N_14791,N_14734,N_14672);
nand U14792 (N_14792,N_14542,N_14519);
or U14793 (N_14793,N_14728,N_14524);
and U14794 (N_14794,N_14528,N_14657);
and U14795 (N_14795,N_14618,N_14547);
or U14796 (N_14796,N_14516,N_14718);
and U14797 (N_14797,N_14624,N_14683);
xnor U14798 (N_14798,N_14652,N_14578);
nor U14799 (N_14799,N_14619,N_14605);
xnor U14800 (N_14800,N_14512,N_14714);
nor U14801 (N_14801,N_14745,N_14522);
and U14802 (N_14802,N_14534,N_14523);
xor U14803 (N_14803,N_14695,N_14703);
nor U14804 (N_14804,N_14564,N_14645);
nand U14805 (N_14805,N_14705,N_14704);
or U14806 (N_14806,N_14599,N_14729);
nand U14807 (N_14807,N_14551,N_14616);
xor U14808 (N_14808,N_14701,N_14737);
and U14809 (N_14809,N_14621,N_14690);
or U14810 (N_14810,N_14576,N_14628);
or U14811 (N_14811,N_14665,N_14552);
nand U14812 (N_14812,N_14513,N_14557);
or U14813 (N_14813,N_14603,N_14543);
nor U14814 (N_14814,N_14583,N_14686);
or U14815 (N_14815,N_14655,N_14632);
nor U14816 (N_14816,N_14749,N_14725);
xor U14817 (N_14817,N_14562,N_14606);
or U14818 (N_14818,N_14692,N_14505);
xnor U14819 (N_14819,N_14678,N_14735);
and U14820 (N_14820,N_14741,N_14653);
nand U14821 (N_14821,N_14640,N_14535);
or U14822 (N_14822,N_14623,N_14720);
xor U14823 (N_14823,N_14698,N_14520);
xor U14824 (N_14824,N_14533,N_14639);
nand U14825 (N_14825,N_14622,N_14651);
and U14826 (N_14826,N_14660,N_14739);
and U14827 (N_14827,N_14685,N_14509);
and U14828 (N_14828,N_14707,N_14712);
nor U14829 (N_14829,N_14575,N_14676);
xor U14830 (N_14830,N_14715,N_14604);
or U14831 (N_14831,N_14631,N_14566);
or U14832 (N_14832,N_14591,N_14546);
or U14833 (N_14833,N_14637,N_14663);
or U14834 (N_14834,N_14681,N_14550);
nor U14835 (N_14835,N_14517,N_14504);
nand U14836 (N_14836,N_14500,N_14738);
nor U14837 (N_14837,N_14514,N_14736);
nor U14838 (N_14838,N_14538,N_14620);
xor U14839 (N_14839,N_14518,N_14588);
xor U14840 (N_14840,N_14677,N_14646);
nor U14841 (N_14841,N_14508,N_14682);
xnor U14842 (N_14842,N_14525,N_14727);
xor U14843 (N_14843,N_14680,N_14555);
and U14844 (N_14844,N_14630,N_14688);
xnor U14845 (N_14845,N_14537,N_14697);
or U14846 (N_14846,N_14561,N_14598);
or U14847 (N_14847,N_14684,N_14613);
xor U14848 (N_14848,N_14614,N_14633);
or U14849 (N_14849,N_14570,N_14612);
nor U14850 (N_14850,N_14596,N_14654);
or U14851 (N_14851,N_14549,N_14669);
nand U14852 (N_14852,N_14638,N_14673);
nand U14853 (N_14853,N_14719,N_14600);
xnor U14854 (N_14854,N_14744,N_14748);
xnor U14855 (N_14855,N_14594,N_14642);
or U14856 (N_14856,N_14501,N_14667);
xnor U14857 (N_14857,N_14579,N_14733);
or U14858 (N_14858,N_14643,N_14545);
and U14859 (N_14859,N_14536,N_14696);
nor U14860 (N_14860,N_14515,N_14636);
nor U14861 (N_14861,N_14503,N_14706);
nor U14862 (N_14862,N_14627,N_14743);
nand U14863 (N_14863,N_14582,N_14726);
or U14864 (N_14864,N_14687,N_14559);
or U14865 (N_14865,N_14584,N_14629);
xnor U14866 (N_14866,N_14710,N_14556);
or U14867 (N_14867,N_14568,N_14611);
xor U14868 (N_14868,N_14723,N_14713);
xor U14869 (N_14869,N_14650,N_14675);
nand U14870 (N_14870,N_14635,N_14607);
or U14871 (N_14871,N_14572,N_14649);
or U14872 (N_14872,N_14541,N_14671);
and U14873 (N_14873,N_14689,N_14731);
nand U14874 (N_14874,N_14511,N_14716);
or U14875 (N_14875,N_14715,N_14539);
xor U14876 (N_14876,N_14705,N_14571);
nand U14877 (N_14877,N_14749,N_14503);
nand U14878 (N_14878,N_14629,N_14572);
xnor U14879 (N_14879,N_14526,N_14516);
nand U14880 (N_14880,N_14717,N_14516);
or U14881 (N_14881,N_14651,N_14733);
and U14882 (N_14882,N_14743,N_14565);
nor U14883 (N_14883,N_14744,N_14735);
xnor U14884 (N_14884,N_14621,N_14747);
nand U14885 (N_14885,N_14583,N_14567);
xor U14886 (N_14886,N_14709,N_14606);
xor U14887 (N_14887,N_14738,N_14634);
and U14888 (N_14888,N_14541,N_14505);
xor U14889 (N_14889,N_14531,N_14599);
nor U14890 (N_14890,N_14531,N_14696);
nor U14891 (N_14891,N_14553,N_14586);
nand U14892 (N_14892,N_14502,N_14548);
or U14893 (N_14893,N_14580,N_14560);
nor U14894 (N_14894,N_14552,N_14657);
and U14895 (N_14895,N_14559,N_14575);
xor U14896 (N_14896,N_14571,N_14657);
nor U14897 (N_14897,N_14691,N_14623);
nand U14898 (N_14898,N_14710,N_14534);
and U14899 (N_14899,N_14633,N_14598);
xor U14900 (N_14900,N_14732,N_14535);
or U14901 (N_14901,N_14616,N_14744);
or U14902 (N_14902,N_14525,N_14643);
nand U14903 (N_14903,N_14533,N_14530);
nor U14904 (N_14904,N_14600,N_14688);
xnor U14905 (N_14905,N_14689,N_14516);
xor U14906 (N_14906,N_14581,N_14680);
or U14907 (N_14907,N_14728,N_14644);
xor U14908 (N_14908,N_14705,N_14643);
xor U14909 (N_14909,N_14739,N_14604);
or U14910 (N_14910,N_14685,N_14562);
xnor U14911 (N_14911,N_14665,N_14728);
and U14912 (N_14912,N_14612,N_14704);
xnor U14913 (N_14913,N_14558,N_14695);
nor U14914 (N_14914,N_14696,N_14584);
nand U14915 (N_14915,N_14595,N_14574);
xnor U14916 (N_14916,N_14562,N_14531);
and U14917 (N_14917,N_14655,N_14664);
xor U14918 (N_14918,N_14501,N_14706);
or U14919 (N_14919,N_14743,N_14519);
nor U14920 (N_14920,N_14679,N_14672);
nor U14921 (N_14921,N_14554,N_14575);
xor U14922 (N_14922,N_14515,N_14669);
nand U14923 (N_14923,N_14727,N_14642);
xnor U14924 (N_14924,N_14708,N_14511);
or U14925 (N_14925,N_14589,N_14700);
nor U14926 (N_14926,N_14699,N_14654);
nand U14927 (N_14927,N_14685,N_14695);
xnor U14928 (N_14928,N_14601,N_14598);
xor U14929 (N_14929,N_14742,N_14569);
nand U14930 (N_14930,N_14748,N_14607);
xnor U14931 (N_14931,N_14662,N_14704);
nor U14932 (N_14932,N_14630,N_14611);
and U14933 (N_14933,N_14530,N_14623);
xnor U14934 (N_14934,N_14513,N_14729);
or U14935 (N_14935,N_14687,N_14682);
and U14936 (N_14936,N_14682,N_14740);
nand U14937 (N_14937,N_14710,N_14729);
nand U14938 (N_14938,N_14547,N_14651);
or U14939 (N_14939,N_14567,N_14519);
and U14940 (N_14940,N_14582,N_14515);
nor U14941 (N_14941,N_14664,N_14500);
nor U14942 (N_14942,N_14511,N_14705);
nand U14943 (N_14943,N_14658,N_14645);
and U14944 (N_14944,N_14508,N_14701);
xnor U14945 (N_14945,N_14577,N_14596);
or U14946 (N_14946,N_14506,N_14557);
nor U14947 (N_14947,N_14617,N_14505);
or U14948 (N_14948,N_14748,N_14511);
xor U14949 (N_14949,N_14659,N_14725);
nand U14950 (N_14950,N_14650,N_14602);
xor U14951 (N_14951,N_14502,N_14550);
xor U14952 (N_14952,N_14572,N_14637);
xor U14953 (N_14953,N_14555,N_14673);
or U14954 (N_14954,N_14571,N_14609);
and U14955 (N_14955,N_14646,N_14669);
nand U14956 (N_14956,N_14669,N_14729);
xor U14957 (N_14957,N_14500,N_14635);
nor U14958 (N_14958,N_14574,N_14693);
or U14959 (N_14959,N_14579,N_14604);
nor U14960 (N_14960,N_14638,N_14557);
nor U14961 (N_14961,N_14526,N_14529);
and U14962 (N_14962,N_14693,N_14736);
or U14963 (N_14963,N_14711,N_14741);
and U14964 (N_14964,N_14561,N_14570);
nor U14965 (N_14965,N_14646,N_14687);
and U14966 (N_14966,N_14601,N_14605);
nor U14967 (N_14967,N_14513,N_14666);
xor U14968 (N_14968,N_14683,N_14656);
or U14969 (N_14969,N_14652,N_14609);
xnor U14970 (N_14970,N_14618,N_14506);
nand U14971 (N_14971,N_14523,N_14505);
xor U14972 (N_14972,N_14684,N_14601);
nor U14973 (N_14973,N_14582,N_14674);
and U14974 (N_14974,N_14524,N_14583);
nand U14975 (N_14975,N_14522,N_14587);
and U14976 (N_14976,N_14544,N_14620);
nor U14977 (N_14977,N_14535,N_14525);
xnor U14978 (N_14978,N_14743,N_14513);
xor U14979 (N_14979,N_14744,N_14677);
and U14980 (N_14980,N_14652,N_14631);
nor U14981 (N_14981,N_14506,N_14502);
xnor U14982 (N_14982,N_14660,N_14686);
and U14983 (N_14983,N_14632,N_14626);
or U14984 (N_14984,N_14537,N_14741);
xor U14985 (N_14985,N_14733,N_14596);
or U14986 (N_14986,N_14710,N_14638);
nor U14987 (N_14987,N_14516,N_14661);
xor U14988 (N_14988,N_14742,N_14667);
or U14989 (N_14989,N_14583,N_14704);
or U14990 (N_14990,N_14622,N_14579);
nor U14991 (N_14991,N_14734,N_14612);
nand U14992 (N_14992,N_14663,N_14720);
nor U14993 (N_14993,N_14677,N_14708);
xor U14994 (N_14994,N_14505,N_14642);
and U14995 (N_14995,N_14575,N_14741);
nand U14996 (N_14996,N_14578,N_14624);
or U14997 (N_14997,N_14590,N_14527);
nor U14998 (N_14998,N_14699,N_14565);
nor U14999 (N_14999,N_14570,N_14536);
xnor U15000 (N_15000,N_14874,N_14995);
xnor U15001 (N_15001,N_14821,N_14921);
and U15002 (N_15002,N_14970,N_14992);
and U15003 (N_15003,N_14952,N_14752);
nand U15004 (N_15004,N_14839,N_14953);
nor U15005 (N_15005,N_14768,N_14879);
and U15006 (N_15006,N_14816,N_14846);
xnor U15007 (N_15007,N_14875,N_14803);
and U15008 (N_15008,N_14829,N_14907);
xnor U15009 (N_15009,N_14905,N_14864);
and U15010 (N_15010,N_14994,N_14997);
nor U15011 (N_15011,N_14884,N_14851);
nor U15012 (N_15012,N_14765,N_14840);
or U15013 (N_15013,N_14871,N_14947);
nor U15014 (N_15014,N_14893,N_14842);
nor U15015 (N_15015,N_14764,N_14941);
and U15016 (N_15016,N_14909,N_14770);
nand U15017 (N_15017,N_14781,N_14996);
or U15018 (N_15018,N_14800,N_14918);
or U15019 (N_15019,N_14930,N_14799);
nand U15020 (N_15020,N_14859,N_14956);
and U15021 (N_15021,N_14906,N_14903);
and U15022 (N_15022,N_14991,N_14807);
xnor U15023 (N_15023,N_14900,N_14759);
nand U15024 (N_15024,N_14897,N_14901);
xnor U15025 (N_15025,N_14817,N_14966);
nor U15026 (N_15026,N_14868,N_14757);
nor U15027 (N_15027,N_14820,N_14965);
xnor U15028 (N_15028,N_14876,N_14910);
nor U15029 (N_15029,N_14948,N_14769);
nand U15030 (N_15030,N_14946,N_14852);
nand U15031 (N_15031,N_14772,N_14908);
nand U15032 (N_15032,N_14976,N_14832);
nor U15033 (N_15033,N_14793,N_14955);
or U15034 (N_15034,N_14964,N_14819);
xnor U15035 (N_15035,N_14971,N_14945);
and U15036 (N_15036,N_14944,N_14830);
or U15037 (N_15037,N_14828,N_14860);
nor U15038 (N_15038,N_14914,N_14806);
and U15039 (N_15039,N_14891,N_14778);
nor U15040 (N_15040,N_14797,N_14935);
nor U15041 (N_15041,N_14812,N_14957);
xnor U15042 (N_15042,N_14815,N_14767);
nand U15043 (N_15043,N_14932,N_14887);
and U15044 (N_15044,N_14889,N_14805);
xnor U15045 (N_15045,N_14755,N_14967);
or U15046 (N_15046,N_14916,N_14831);
or U15047 (N_15047,N_14931,N_14870);
and U15048 (N_15048,N_14766,N_14802);
or U15049 (N_15049,N_14890,N_14938);
or U15050 (N_15050,N_14998,N_14885);
nand U15051 (N_15051,N_14969,N_14934);
xnor U15052 (N_15052,N_14989,N_14915);
xnor U15053 (N_15053,N_14977,N_14895);
nor U15054 (N_15054,N_14827,N_14987);
and U15055 (N_15055,N_14773,N_14788);
or U15056 (N_15056,N_14863,N_14758);
nand U15057 (N_15057,N_14818,N_14974);
nand U15058 (N_15058,N_14917,N_14779);
xor U15059 (N_15059,N_14942,N_14960);
xnor U15060 (N_15060,N_14980,N_14902);
and U15061 (N_15061,N_14867,N_14865);
or U15062 (N_15062,N_14933,N_14954);
nand U15063 (N_15063,N_14795,N_14899);
nand U15064 (N_15064,N_14973,N_14801);
xor U15065 (N_15065,N_14894,N_14858);
nand U15066 (N_15066,N_14835,N_14959);
nand U15067 (N_15067,N_14873,N_14883);
nor U15068 (N_15068,N_14898,N_14754);
nor U15069 (N_15069,N_14784,N_14882);
xnor U15070 (N_15070,N_14928,N_14990);
xor U15071 (N_15071,N_14834,N_14920);
or U15072 (N_15072,N_14927,N_14872);
or U15073 (N_15073,N_14854,N_14822);
xor U15074 (N_15074,N_14913,N_14923);
or U15075 (N_15075,N_14837,N_14789);
xnor U15076 (N_15076,N_14792,N_14919);
nor U15077 (N_15077,N_14826,N_14937);
xnor U15078 (N_15078,N_14975,N_14986);
and U15079 (N_15079,N_14787,N_14940);
nor U15080 (N_15080,N_14836,N_14968);
or U15081 (N_15081,N_14763,N_14813);
nor U15082 (N_15082,N_14929,N_14753);
nor U15083 (N_15083,N_14774,N_14847);
nand U15084 (N_15084,N_14783,N_14841);
nand U15085 (N_15085,N_14825,N_14756);
nand U15086 (N_15086,N_14886,N_14843);
or U15087 (N_15087,N_14888,N_14761);
nand U15088 (N_15088,N_14866,N_14896);
xnor U15089 (N_15089,N_14809,N_14869);
nor U15090 (N_15090,N_14877,N_14853);
xor U15091 (N_15091,N_14939,N_14861);
nand U15092 (N_15092,N_14911,N_14750);
nor U15093 (N_15093,N_14833,N_14862);
xnor U15094 (N_15094,N_14762,N_14985);
or U15095 (N_15095,N_14979,N_14777);
nand U15096 (N_15096,N_14844,N_14760);
xor U15097 (N_15097,N_14904,N_14785);
or U15098 (N_15098,N_14892,N_14978);
nor U15099 (N_15099,N_14961,N_14982);
or U15100 (N_15100,N_14924,N_14811);
nor U15101 (N_15101,N_14776,N_14845);
nor U15102 (N_15102,N_14775,N_14925);
xnor U15103 (N_15103,N_14880,N_14878);
xnor U15104 (N_15104,N_14856,N_14824);
or U15105 (N_15105,N_14855,N_14962);
nand U15106 (N_15106,N_14780,N_14798);
nand U15107 (N_15107,N_14796,N_14771);
xor U15108 (N_15108,N_14794,N_14786);
xnor U15109 (N_15109,N_14988,N_14814);
nand U15110 (N_15110,N_14823,N_14848);
or U15111 (N_15111,N_14912,N_14850);
nor U15112 (N_15112,N_14922,N_14782);
xnor U15113 (N_15113,N_14936,N_14972);
and U15114 (N_15114,N_14810,N_14808);
nor U15115 (N_15115,N_14838,N_14881);
xor U15116 (N_15116,N_14857,N_14981);
and U15117 (N_15117,N_14791,N_14849);
nor U15118 (N_15118,N_14984,N_14993);
nor U15119 (N_15119,N_14804,N_14983);
and U15120 (N_15120,N_14951,N_14943);
or U15121 (N_15121,N_14949,N_14790);
xor U15122 (N_15122,N_14963,N_14926);
xnor U15123 (N_15123,N_14958,N_14950);
or U15124 (N_15124,N_14751,N_14999);
nor U15125 (N_15125,N_14827,N_14883);
or U15126 (N_15126,N_14911,N_14801);
and U15127 (N_15127,N_14978,N_14816);
nor U15128 (N_15128,N_14864,N_14990);
nor U15129 (N_15129,N_14909,N_14824);
nor U15130 (N_15130,N_14997,N_14973);
or U15131 (N_15131,N_14984,N_14798);
xor U15132 (N_15132,N_14772,N_14881);
nor U15133 (N_15133,N_14887,N_14935);
xor U15134 (N_15134,N_14993,N_14856);
xnor U15135 (N_15135,N_14790,N_14774);
or U15136 (N_15136,N_14926,N_14817);
xor U15137 (N_15137,N_14825,N_14827);
and U15138 (N_15138,N_14818,N_14939);
xor U15139 (N_15139,N_14822,N_14751);
or U15140 (N_15140,N_14920,N_14840);
or U15141 (N_15141,N_14878,N_14943);
and U15142 (N_15142,N_14885,N_14831);
nor U15143 (N_15143,N_14900,N_14810);
nor U15144 (N_15144,N_14817,N_14792);
nand U15145 (N_15145,N_14942,N_14982);
or U15146 (N_15146,N_14960,N_14868);
nor U15147 (N_15147,N_14989,N_14978);
or U15148 (N_15148,N_14938,N_14972);
xnor U15149 (N_15149,N_14857,N_14975);
or U15150 (N_15150,N_14892,N_14998);
xnor U15151 (N_15151,N_14942,N_14941);
nor U15152 (N_15152,N_14773,N_14913);
and U15153 (N_15153,N_14821,N_14802);
xnor U15154 (N_15154,N_14984,N_14889);
nand U15155 (N_15155,N_14757,N_14951);
xnor U15156 (N_15156,N_14911,N_14780);
xor U15157 (N_15157,N_14999,N_14952);
nand U15158 (N_15158,N_14922,N_14940);
or U15159 (N_15159,N_14769,N_14799);
nor U15160 (N_15160,N_14910,N_14964);
xnor U15161 (N_15161,N_14795,N_14996);
nand U15162 (N_15162,N_14828,N_14793);
xor U15163 (N_15163,N_14860,N_14880);
and U15164 (N_15164,N_14976,N_14920);
nand U15165 (N_15165,N_14932,N_14773);
and U15166 (N_15166,N_14925,N_14862);
xnor U15167 (N_15167,N_14911,N_14824);
and U15168 (N_15168,N_14936,N_14853);
and U15169 (N_15169,N_14807,N_14800);
or U15170 (N_15170,N_14953,N_14883);
nand U15171 (N_15171,N_14970,N_14920);
nand U15172 (N_15172,N_14859,N_14768);
xnor U15173 (N_15173,N_14992,N_14833);
xor U15174 (N_15174,N_14980,N_14750);
nor U15175 (N_15175,N_14794,N_14848);
xnor U15176 (N_15176,N_14768,N_14850);
nand U15177 (N_15177,N_14967,N_14799);
and U15178 (N_15178,N_14788,N_14857);
xor U15179 (N_15179,N_14955,N_14853);
and U15180 (N_15180,N_14766,N_14828);
or U15181 (N_15181,N_14803,N_14923);
and U15182 (N_15182,N_14808,N_14774);
nand U15183 (N_15183,N_14934,N_14878);
nor U15184 (N_15184,N_14759,N_14901);
xnor U15185 (N_15185,N_14844,N_14856);
xnor U15186 (N_15186,N_14852,N_14891);
xor U15187 (N_15187,N_14854,N_14803);
nor U15188 (N_15188,N_14769,N_14998);
nand U15189 (N_15189,N_14763,N_14791);
nor U15190 (N_15190,N_14869,N_14819);
and U15191 (N_15191,N_14839,N_14996);
nor U15192 (N_15192,N_14964,N_14888);
or U15193 (N_15193,N_14877,N_14796);
or U15194 (N_15194,N_14800,N_14828);
nor U15195 (N_15195,N_14811,N_14764);
nand U15196 (N_15196,N_14916,N_14802);
nand U15197 (N_15197,N_14986,N_14849);
and U15198 (N_15198,N_14799,N_14772);
or U15199 (N_15199,N_14928,N_14960);
nand U15200 (N_15200,N_14848,N_14806);
or U15201 (N_15201,N_14829,N_14917);
xnor U15202 (N_15202,N_14783,N_14931);
nor U15203 (N_15203,N_14774,N_14891);
and U15204 (N_15204,N_14785,N_14756);
nor U15205 (N_15205,N_14902,N_14827);
nor U15206 (N_15206,N_14941,N_14965);
nor U15207 (N_15207,N_14991,N_14908);
xor U15208 (N_15208,N_14994,N_14982);
nand U15209 (N_15209,N_14802,N_14846);
and U15210 (N_15210,N_14989,N_14868);
nor U15211 (N_15211,N_14981,N_14973);
nand U15212 (N_15212,N_14933,N_14758);
nor U15213 (N_15213,N_14954,N_14991);
xor U15214 (N_15214,N_14959,N_14877);
or U15215 (N_15215,N_14943,N_14880);
or U15216 (N_15216,N_14757,N_14777);
nand U15217 (N_15217,N_14933,N_14904);
xor U15218 (N_15218,N_14928,N_14968);
or U15219 (N_15219,N_14764,N_14781);
nor U15220 (N_15220,N_14901,N_14839);
and U15221 (N_15221,N_14818,N_14883);
xor U15222 (N_15222,N_14835,N_14894);
or U15223 (N_15223,N_14958,N_14812);
nand U15224 (N_15224,N_14769,N_14814);
nand U15225 (N_15225,N_14997,N_14962);
and U15226 (N_15226,N_14802,N_14948);
nand U15227 (N_15227,N_14886,N_14958);
and U15228 (N_15228,N_14898,N_14821);
nor U15229 (N_15229,N_14850,N_14874);
or U15230 (N_15230,N_14958,N_14960);
xnor U15231 (N_15231,N_14952,N_14921);
nand U15232 (N_15232,N_14803,N_14754);
and U15233 (N_15233,N_14755,N_14996);
and U15234 (N_15234,N_14890,N_14917);
xor U15235 (N_15235,N_14989,N_14930);
and U15236 (N_15236,N_14917,N_14815);
nor U15237 (N_15237,N_14866,N_14963);
nand U15238 (N_15238,N_14857,N_14865);
and U15239 (N_15239,N_14767,N_14766);
xor U15240 (N_15240,N_14838,N_14931);
or U15241 (N_15241,N_14796,N_14886);
xor U15242 (N_15242,N_14995,N_14856);
nor U15243 (N_15243,N_14971,N_14808);
nor U15244 (N_15244,N_14916,N_14765);
and U15245 (N_15245,N_14907,N_14925);
nor U15246 (N_15246,N_14811,N_14867);
and U15247 (N_15247,N_14885,N_14921);
nand U15248 (N_15248,N_14893,N_14868);
nand U15249 (N_15249,N_14996,N_14902);
or U15250 (N_15250,N_15111,N_15185);
or U15251 (N_15251,N_15010,N_15049);
xnor U15252 (N_15252,N_15142,N_15071);
nand U15253 (N_15253,N_15220,N_15126);
xnor U15254 (N_15254,N_15044,N_15131);
and U15255 (N_15255,N_15163,N_15150);
nand U15256 (N_15256,N_15171,N_15029);
and U15257 (N_15257,N_15184,N_15034);
nor U15258 (N_15258,N_15036,N_15246);
or U15259 (N_15259,N_15221,N_15188);
or U15260 (N_15260,N_15177,N_15075);
nor U15261 (N_15261,N_15038,N_15240);
nor U15262 (N_15262,N_15170,N_15008);
xnor U15263 (N_15263,N_15067,N_15074);
and U15264 (N_15264,N_15080,N_15230);
or U15265 (N_15265,N_15066,N_15143);
nand U15266 (N_15266,N_15024,N_15238);
nand U15267 (N_15267,N_15204,N_15091);
nand U15268 (N_15268,N_15026,N_15200);
xnor U15269 (N_15269,N_15103,N_15187);
nand U15270 (N_15270,N_15181,N_15212);
nand U15271 (N_15271,N_15242,N_15249);
and U15272 (N_15272,N_15015,N_15082);
nand U15273 (N_15273,N_15206,N_15144);
and U15274 (N_15274,N_15118,N_15198);
or U15275 (N_15275,N_15194,N_15209);
xnor U15276 (N_15276,N_15175,N_15048);
nand U15277 (N_15277,N_15125,N_15215);
and U15278 (N_15278,N_15226,N_15234);
and U15279 (N_15279,N_15011,N_15006);
nand U15280 (N_15280,N_15179,N_15014);
xor U15281 (N_15281,N_15000,N_15173);
nand U15282 (N_15282,N_15197,N_15135);
or U15283 (N_15283,N_15040,N_15012);
or U15284 (N_15284,N_15065,N_15033);
or U15285 (N_15285,N_15155,N_15043);
or U15286 (N_15286,N_15133,N_15057);
nand U15287 (N_15287,N_15153,N_15207);
nand U15288 (N_15288,N_15019,N_15028);
and U15289 (N_15289,N_15132,N_15025);
or U15290 (N_15290,N_15104,N_15094);
and U15291 (N_15291,N_15076,N_15053);
nor U15292 (N_15292,N_15121,N_15102);
nor U15293 (N_15293,N_15077,N_15116);
xnor U15294 (N_15294,N_15004,N_15001);
xor U15295 (N_15295,N_15203,N_15083);
nand U15296 (N_15296,N_15223,N_15106);
and U15297 (N_15297,N_15139,N_15084);
or U15298 (N_15298,N_15162,N_15146);
nor U15299 (N_15299,N_15069,N_15086);
or U15300 (N_15300,N_15013,N_15101);
nand U15301 (N_15301,N_15037,N_15222);
nor U15302 (N_15302,N_15214,N_15055);
xnor U15303 (N_15303,N_15201,N_15031);
nor U15304 (N_15304,N_15191,N_15023);
or U15305 (N_15305,N_15039,N_15099);
xor U15306 (N_15306,N_15003,N_15231);
nand U15307 (N_15307,N_15138,N_15107);
xnor U15308 (N_15308,N_15156,N_15047);
nor U15309 (N_15309,N_15061,N_15169);
or U15310 (N_15310,N_15009,N_15159);
xnor U15311 (N_15311,N_15237,N_15167);
nor U15312 (N_15312,N_15202,N_15196);
nor U15313 (N_15313,N_15217,N_15152);
xor U15314 (N_15314,N_15161,N_15166);
nand U15315 (N_15315,N_15193,N_15064);
nor U15316 (N_15316,N_15241,N_15151);
xnor U15317 (N_15317,N_15149,N_15190);
xor U15318 (N_15318,N_15072,N_15136);
and U15319 (N_15319,N_15228,N_15005);
nand U15320 (N_15320,N_15141,N_15092);
xor U15321 (N_15321,N_15128,N_15002);
and U15322 (N_15322,N_15079,N_15225);
and U15323 (N_15323,N_15165,N_15060);
or U15324 (N_15324,N_15158,N_15090);
nor U15325 (N_15325,N_15120,N_15210);
or U15326 (N_15326,N_15195,N_15045);
or U15327 (N_15327,N_15063,N_15218);
and U15328 (N_15328,N_15227,N_15030);
and U15329 (N_15329,N_15224,N_15216);
nand U15330 (N_15330,N_15186,N_15088);
or U15331 (N_15331,N_15022,N_15042);
and U15332 (N_15332,N_15174,N_15095);
nor U15333 (N_15333,N_15148,N_15239);
nand U15334 (N_15334,N_15062,N_15050);
nand U15335 (N_15335,N_15105,N_15180);
and U15336 (N_15336,N_15233,N_15122);
nor U15337 (N_15337,N_15020,N_15130);
or U15338 (N_15338,N_15229,N_15017);
and U15339 (N_15339,N_15127,N_15245);
and U15340 (N_15340,N_15054,N_15182);
xnor U15341 (N_15341,N_15089,N_15124);
and U15342 (N_15342,N_15235,N_15056);
xor U15343 (N_15343,N_15093,N_15100);
or U15344 (N_15344,N_15113,N_15081);
and U15345 (N_15345,N_15244,N_15137);
xor U15346 (N_15346,N_15160,N_15032);
and U15347 (N_15347,N_15119,N_15157);
nor U15348 (N_15348,N_15108,N_15236);
nand U15349 (N_15349,N_15247,N_15018);
and U15350 (N_15350,N_15219,N_15147);
nand U15351 (N_15351,N_15097,N_15051);
and U15352 (N_15352,N_15058,N_15248);
or U15353 (N_15353,N_15211,N_15052);
xor U15354 (N_15354,N_15154,N_15199);
and U15355 (N_15355,N_15243,N_15007);
nand U15356 (N_15356,N_15232,N_15129);
nand U15357 (N_15357,N_15134,N_15046);
or U15358 (N_15358,N_15192,N_15145);
nand U15359 (N_15359,N_15183,N_15109);
nor U15360 (N_15360,N_15070,N_15016);
xor U15361 (N_15361,N_15176,N_15087);
nand U15362 (N_15362,N_15059,N_15085);
nand U15363 (N_15363,N_15027,N_15021);
xnor U15364 (N_15364,N_15168,N_15208);
and U15365 (N_15365,N_15073,N_15117);
xnor U15366 (N_15366,N_15035,N_15041);
or U15367 (N_15367,N_15112,N_15189);
and U15368 (N_15368,N_15096,N_15164);
nor U15369 (N_15369,N_15205,N_15178);
nand U15370 (N_15370,N_15068,N_15213);
xor U15371 (N_15371,N_15110,N_15115);
xnor U15372 (N_15372,N_15098,N_15078);
xor U15373 (N_15373,N_15123,N_15140);
or U15374 (N_15374,N_15114,N_15172);
nand U15375 (N_15375,N_15166,N_15125);
nor U15376 (N_15376,N_15240,N_15131);
or U15377 (N_15377,N_15012,N_15203);
xor U15378 (N_15378,N_15198,N_15019);
xnor U15379 (N_15379,N_15079,N_15092);
xnor U15380 (N_15380,N_15204,N_15026);
or U15381 (N_15381,N_15111,N_15196);
nand U15382 (N_15382,N_15181,N_15164);
xnor U15383 (N_15383,N_15014,N_15068);
nor U15384 (N_15384,N_15030,N_15100);
xnor U15385 (N_15385,N_15126,N_15005);
and U15386 (N_15386,N_15091,N_15070);
and U15387 (N_15387,N_15052,N_15036);
xnor U15388 (N_15388,N_15111,N_15166);
nor U15389 (N_15389,N_15079,N_15057);
nor U15390 (N_15390,N_15187,N_15102);
nand U15391 (N_15391,N_15127,N_15121);
or U15392 (N_15392,N_15091,N_15003);
nand U15393 (N_15393,N_15095,N_15043);
and U15394 (N_15394,N_15035,N_15050);
nor U15395 (N_15395,N_15219,N_15201);
and U15396 (N_15396,N_15109,N_15059);
xor U15397 (N_15397,N_15244,N_15061);
nand U15398 (N_15398,N_15137,N_15002);
and U15399 (N_15399,N_15176,N_15217);
and U15400 (N_15400,N_15173,N_15159);
nor U15401 (N_15401,N_15247,N_15243);
nor U15402 (N_15402,N_15178,N_15199);
and U15403 (N_15403,N_15153,N_15177);
and U15404 (N_15404,N_15056,N_15141);
nor U15405 (N_15405,N_15043,N_15188);
or U15406 (N_15406,N_15183,N_15021);
or U15407 (N_15407,N_15131,N_15170);
nor U15408 (N_15408,N_15140,N_15017);
xor U15409 (N_15409,N_15202,N_15229);
nand U15410 (N_15410,N_15207,N_15159);
xnor U15411 (N_15411,N_15044,N_15043);
xnor U15412 (N_15412,N_15119,N_15138);
xor U15413 (N_15413,N_15244,N_15184);
nor U15414 (N_15414,N_15206,N_15146);
and U15415 (N_15415,N_15102,N_15172);
nand U15416 (N_15416,N_15184,N_15131);
nand U15417 (N_15417,N_15203,N_15077);
or U15418 (N_15418,N_15002,N_15214);
or U15419 (N_15419,N_15086,N_15066);
xor U15420 (N_15420,N_15145,N_15101);
nand U15421 (N_15421,N_15006,N_15074);
nand U15422 (N_15422,N_15177,N_15004);
and U15423 (N_15423,N_15001,N_15211);
xor U15424 (N_15424,N_15245,N_15238);
and U15425 (N_15425,N_15156,N_15168);
nand U15426 (N_15426,N_15203,N_15141);
nor U15427 (N_15427,N_15193,N_15036);
nor U15428 (N_15428,N_15148,N_15039);
nor U15429 (N_15429,N_15056,N_15075);
or U15430 (N_15430,N_15142,N_15164);
xnor U15431 (N_15431,N_15122,N_15230);
xnor U15432 (N_15432,N_15007,N_15147);
nor U15433 (N_15433,N_15126,N_15195);
nand U15434 (N_15434,N_15109,N_15243);
xor U15435 (N_15435,N_15007,N_15013);
nand U15436 (N_15436,N_15115,N_15105);
xor U15437 (N_15437,N_15101,N_15135);
and U15438 (N_15438,N_15244,N_15038);
nand U15439 (N_15439,N_15113,N_15127);
nor U15440 (N_15440,N_15074,N_15126);
xor U15441 (N_15441,N_15107,N_15142);
nor U15442 (N_15442,N_15111,N_15079);
and U15443 (N_15443,N_15197,N_15107);
and U15444 (N_15444,N_15122,N_15100);
and U15445 (N_15445,N_15026,N_15016);
and U15446 (N_15446,N_15126,N_15072);
xor U15447 (N_15447,N_15182,N_15043);
or U15448 (N_15448,N_15113,N_15194);
xnor U15449 (N_15449,N_15078,N_15162);
xnor U15450 (N_15450,N_15194,N_15058);
nand U15451 (N_15451,N_15126,N_15208);
or U15452 (N_15452,N_15042,N_15019);
nand U15453 (N_15453,N_15128,N_15042);
nor U15454 (N_15454,N_15006,N_15099);
and U15455 (N_15455,N_15143,N_15086);
nand U15456 (N_15456,N_15249,N_15241);
nand U15457 (N_15457,N_15221,N_15025);
or U15458 (N_15458,N_15219,N_15082);
and U15459 (N_15459,N_15030,N_15138);
or U15460 (N_15460,N_15005,N_15212);
nor U15461 (N_15461,N_15240,N_15178);
nor U15462 (N_15462,N_15104,N_15162);
and U15463 (N_15463,N_15001,N_15108);
nand U15464 (N_15464,N_15186,N_15210);
xnor U15465 (N_15465,N_15012,N_15099);
and U15466 (N_15466,N_15247,N_15129);
and U15467 (N_15467,N_15005,N_15131);
or U15468 (N_15468,N_15016,N_15059);
nand U15469 (N_15469,N_15240,N_15170);
xnor U15470 (N_15470,N_15239,N_15105);
nand U15471 (N_15471,N_15248,N_15235);
nand U15472 (N_15472,N_15046,N_15245);
nand U15473 (N_15473,N_15023,N_15088);
and U15474 (N_15474,N_15114,N_15163);
nand U15475 (N_15475,N_15213,N_15007);
nand U15476 (N_15476,N_15148,N_15146);
nand U15477 (N_15477,N_15019,N_15066);
xnor U15478 (N_15478,N_15041,N_15047);
nor U15479 (N_15479,N_15012,N_15146);
nor U15480 (N_15480,N_15016,N_15160);
nand U15481 (N_15481,N_15126,N_15159);
nor U15482 (N_15482,N_15040,N_15179);
nand U15483 (N_15483,N_15003,N_15160);
nand U15484 (N_15484,N_15090,N_15191);
and U15485 (N_15485,N_15059,N_15180);
and U15486 (N_15486,N_15046,N_15158);
and U15487 (N_15487,N_15142,N_15037);
nand U15488 (N_15488,N_15018,N_15114);
xnor U15489 (N_15489,N_15120,N_15106);
xnor U15490 (N_15490,N_15095,N_15113);
or U15491 (N_15491,N_15112,N_15049);
xor U15492 (N_15492,N_15020,N_15183);
or U15493 (N_15493,N_15145,N_15164);
or U15494 (N_15494,N_15162,N_15053);
xor U15495 (N_15495,N_15006,N_15023);
nand U15496 (N_15496,N_15000,N_15091);
and U15497 (N_15497,N_15229,N_15081);
nand U15498 (N_15498,N_15019,N_15006);
nand U15499 (N_15499,N_15215,N_15037);
xnor U15500 (N_15500,N_15313,N_15298);
nand U15501 (N_15501,N_15427,N_15403);
xor U15502 (N_15502,N_15318,N_15417);
xnor U15503 (N_15503,N_15320,N_15344);
nor U15504 (N_15504,N_15434,N_15294);
nor U15505 (N_15505,N_15454,N_15285);
and U15506 (N_15506,N_15253,N_15306);
and U15507 (N_15507,N_15437,N_15472);
or U15508 (N_15508,N_15431,N_15464);
xor U15509 (N_15509,N_15351,N_15354);
xnor U15510 (N_15510,N_15453,N_15451);
and U15511 (N_15511,N_15268,N_15392);
xor U15512 (N_15512,N_15433,N_15394);
and U15513 (N_15513,N_15481,N_15442);
or U15514 (N_15514,N_15452,N_15468);
nor U15515 (N_15515,N_15339,N_15273);
and U15516 (N_15516,N_15415,N_15416);
and U15517 (N_15517,N_15422,N_15343);
or U15518 (N_15518,N_15301,N_15419);
or U15519 (N_15519,N_15488,N_15496);
nor U15520 (N_15520,N_15439,N_15372);
and U15521 (N_15521,N_15336,N_15328);
or U15522 (N_15522,N_15323,N_15347);
nand U15523 (N_15523,N_15400,N_15469);
nand U15524 (N_15524,N_15492,N_15293);
nand U15525 (N_15525,N_15305,N_15258);
or U15526 (N_15526,N_15438,N_15460);
nor U15527 (N_15527,N_15441,N_15310);
or U15528 (N_15528,N_15280,N_15383);
nand U15529 (N_15529,N_15399,N_15369);
nand U15530 (N_15530,N_15428,N_15477);
xnor U15531 (N_15531,N_15390,N_15282);
xnor U15532 (N_15532,N_15362,N_15319);
xor U15533 (N_15533,N_15283,N_15259);
nor U15534 (N_15534,N_15334,N_15317);
and U15535 (N_15535,N_15277,N_15395);
xor U15536 (N_15536,N_15377,N_15495);
nor U15537 (N_15537,N_15489,N_15482);
nor U15538 (N_15538,N_15291,N_15455);
or U15539 (N_15539,N_15288,N_15389);
or U15540 (N_15540,N_15474,N_15370);
nor U15541 (N_15541,N_15497,N_15411);
nor U15542 (N_15542,N_15420,N_15274);
and U15543 (N_15543,N_15322,N_15401);
nand U15544 (N_15544,N_15286,N_15467);
nand U15545 (N_15545,N_15487,N_15311);
and U15546 (N_15546,N_15486,N_15251);
nand U15547 (N_15547,N_15479,N_15379);
and U15548 (N_15548,N_15376,N_15295);
nor U15549 (N_15549,N_15314,N_15429);
xor U15550 (N_15550,N_15413,N_15375);
nand U15551 (N_15551,N_15360,N_15459);
or U15552 (N_15552,N_15367,N_15304);
and U15553 (N_15553,N_15350,N_15443);
nor U15554 (N_15554,N_15326,N_15255);
nor U15555 (N_15555,N_15475,N_15353);
and U15556 (N_15556,N_15287,N_15470);
or U15557 (N_15557,N_15358,N_15312);
and U15558 (N_15558,N_15348,N_15299);
nand U15559 (N_15559,N_15426,N_15483);
xor U15560 (N_15560,N_15393,N_15342);
or U15561 (N_15561,N_15478,N_15378);
and U15562 (N_15562,N_15466,N_15391);
nor U15563 (N_15563,N_15456,N_15352);
nor U15564 (N_15564,N_15254,N_15397);
xor U15565 (N_15565,N_15414,N_15361);
or U15566 (N_15566,N_15316,N_15335);
nand U15567 (N_15567,N_15292,N_15385);
xor U15568 (N_15568,N_15484,N_15345);
or U15569 (N_15569,N_15265,N_15386);
or U15570 (N_15570,N_15359,N_15449);
nand U15571 (N_15571,N_15333,N_15406);
xor U15572 (N_15572,N_15357,N_15279);
nand U15573 (N_15573,N_15337,N_15499);
xor U15574 (N_15574,N_15463,N_15398);
nand U15575 (N_15575,N_15424,N_15296);
nand U15576 (N_15576,N_15471,N_15410);
and U15577 (N_15577,N_15366,N_15260);
xnor U15578 (N_15578,N_15445,N_15480);
nand U15579 (N_15579,N_15261,N_15380);
or U15580 (N_15580,N_15269,N_15450);
nand U15581 (N_15581,N_15412,N_15373);
nand U15582 (N_15582,N_15325,N_15462);
xor U15583 (N_15583,N_15498,N_15284);
nand U15584 (N_15584,N_15270,N_15271);
nor U15585 (N_15585,N_15374,N_15331);
xnor U15586 (N_15586,N_15262,N_15368);
nor U15587 (N_15587,N_15307,N_15446);
and U15588 (N_15588,N_15256,N_15444);
xnor U15589 (N_15589,N_15384,N_15289);
and U15590 (N_15590,N_15266,N_15302);
or U15591 (N_15591,N_15447,N_15473);
xor U15592 (N_15592,N_15388,N_15272);
and U15593 (N_15593,N_15409,N_15290);
nand U15594 (N_15594,N_15494,N_15267);
xnor U15595 (N_15595,N_15332,N_15363);
or U15596 (N_15596,N_15341,N_15321);
nand U15597 (N_15597,N_15387,N_15457);
xor U15598 (N_15598,N_15476,N_15440);
or U15599 (N_15599,N_15327,N_15324);
nor U15600 (N_15600,N_15264,N_15381);
nor U15601 (N_15601,N_15418,N_15448);
nand U15602 (N_15602,N_15315,N_15408);
and U15603 (N_15603,N_15329,N_15465);
nor U15604 (N_15604,N_15300,N_15330);
nor U15605 (N_15605,N_15297,N_15309);
and U15606 (N_15606,N_15436,N_15461);
xnor U15607 (N_15607,N_15281,N_15491);
xor U15608 (N_15608,N_15364,N_15252);
nor U15609 (N_15609,N_15346,N_15430);
or U15610 (N_15610,N_15404,N_15250);
or U15611 (N_15611,N_15421,N_15355);
and U15612 (N_15612,N_15485,N_15425);
nor U15613 (N_15613,N_15371,N_15276);
nand U15614 (N_15614,N_15432,N_15458);
nor U15615 (N_15615,N_15338,N_15382);
xnor U15616 (N_15616,N_15490,N_15275);
xor U15617 (N_15617,N_15423,N_15303);
nor U15618 (N_15618,N_15435,N_15263);
xor U15619 (N_15619,N_15340,N_15349);
xnor U15620 (N_15620,N_15308,N_15356);
nor U15621 (N_15621,N_15365,N_15278);
nand U15622 (N_15622,N_15257,N_15405);
nand U15623 (N_15623,N_15493,N_15407);
and U15624 (N_15624,N_15402,N_15396);
xor U15625 (N_15625,N_15473,N_15407);
or U15626 (N_15626,N_15273,N_15498);
or U15627 (N_15627,N_15463,N_15387);
or U15628 (N_15628,N_15327,N_15286);
nor U15629 (N_15629,N_15377,N_15360);
or U15630 (N_15630,N_15451,N_15346);
or U15631 (N_15631,N_15350,N_15330);
nand U15632 (N_15632,N_15424,N_15313);
nor U15633 (N_15633,N_15473,N_15441);
nand U15634 (N_15634,N_15433,N_15369);
xnor U15635 (N_15635,N_15468,N_15483);
nor U15636 (N_15636,N_15263,N_15354);
nand U15637 (N_15637,N_15260,N_15307);
nand U15638 (N_15638,N_15291,N_15394);
nand U15639 (N_15639,N_15373,N_15331);
or U15640 (N_15640,N_15384,N_15370);
and U15641 (N_15641,N_15455,N_15420);
nand U15642 (N_15642,N_15321,N_15467);
or U15643 (N_15643,N_15485,N_15470);
nand U15644 (N_15644,N_15266,N_15314);
xor U15645 (N_15645,N_15333,N_15442);
and U15646 (N_15646,N_15307,N_15427);
nand U15647 (N_15647,N_15440,N_15306);
or U15648 (N_15648,N_15471,N_15252);
and U15649 (N_15649,N_15310,N_15445);
or U15650 (N_15650,N_15255,N_15452);
nor U15651 (N_15651,N_15261,N_15387);
and U15652 (N_15652,N_15496,N_15478);
xor U15653 (N_15653,N_15385,N_15300);
or U15654 (N_15654,N_15292,N_15400);
nor U15655 (N_15655,N_15271,N_15422);
and U15656 (N_15656,N_15281,N_15418);
or U15657 (N_15657,N_15324,N_15415);
xnor U15658 (N_15658,N_15268,N_15446);
nor U15659 (N_15659,N_15493,N_15390);
or U15660 (N_15660,N_15280,N_15419);
nand U15661 (N_15661,N_15366,N_15254);
or U15662 (N_15662,N_15301,N_15486);
nand U15663 (N_15663,N_15372,N_15262);
nor U15664 (N_15664,N_15302,N_15279);
or U15665 (N_15665,N_15258,N_15462);
nor U15666 (N_15666,N_15499,N_15455);
xnor U15667 (N_15667,N_15386,N_15429);
xor U15668 (N_15668,N_15409,N_15469);
or U15669 (N_15669,N_15315,N_15429);
and U15670 (N_15670,N_15394,N_15405);
or U15671 (N_15671,N_15429,N_15262);
nand U15672 (N_15672,N_15320,N_15473);
nor U15673 (N_15673,N_15290,N_15433);
nand U15674 (N_15674,N_15416,N_15291);
nor U15675 (N_15675,N_15392,N_15499);
nor U15676 (N_15676,N_15490,N_15312);
nand U15677 (N_15677,N_15270,N_15405);
nor U15678 (N_15678,N_15290,N_15370);
nor U15679 (N_15679,N_15357,N_15380);
nand U15680 (N_15680,N_15370,N_15472);
nand U15681 (N_15681,N_15490,N_15274);
nand U15682 (N_15682,N_15313,N_15289);
nand U15683 (N_15683,N_15365,N_15489);
nand U15684 (N_15684,N_15446,N_15350);
or U15685 (N_15685,N_15314,N_15492);
nand U15686 (N_15686,N_15372,N_15484);
and U15687 (N_15687,N_15476,N_15361);
and U15688 (N_15688,N_15496,N_15292);
xnor U15689 (N_15689,N_15272,N_15428);
and U15690 (N_15690,N_15289,N_15451);
and U15691 (N_15691,N_15445,N_15342);
nand U15692 (N_15692,N_15469,N_15453);
nor U15693 (N_15693,N_15302,N_15388);
or U15694 (N_15694,N_15373,N_15302);
xnor U15695 (N_15695,N_15401,N_15438);
or U15696 (N_15696,N_15352,N_15490);
nand U15697 (N_15697,N_15401,N_15286);
nand U15698 (N_15698,N_15448,N_15253);
or U15699 (N_15699,N_15463,N_15434);
or U15700 (N_15700,N_15253,N_15278);
nor U15701 (N_15701,N_15454,N_15442);
nor U15702 (N_15702,N_15354,N_15474);
xor U15703 (N_15703,N_15340,N_15391);
or U15704 (N_15704,N_15308,N_15448);
nand U15705 (N_15705,N_15443,N_15288);
nand U15706 (N_15706,N_15453,N_15391);
xor U15707 (N_15707,N_15350,N_15284);
and U15708 (N_15708,N_15332,N_15425);
and U15709 (N_15709,N_15475,N_15310);
xnor U15710 (N_15710,N_15453,N_15413);
nand U15711 (N_15711,N_15287,N_15478);
and U15712 (N_15712,N_15422,N_15341);
xnor U15713 (N_15713,N_15309,N_15286);
xnor U15714 (N_15714,N_15340,N_15264);
and U15715 (N_15715,N_15374,N_15327);
nor U15716 (N_15716,N_15438,N_15311);
nand U15717 (N_15717,N_15451,N_15434);
xnor U15718 (N_15718,N_15477,N_15269);
or U15719 (N_15719,N_15418,N_15292);
nor U15720 (N_15720,N_15487,N_15483);
nor U15721 (N_15721,N_15384,N_15394);
xor U15722 (N_15722,N_15266,N_15301);
nand U15723 (N_15723,N_15332,N_15253);
or U15724 (N_15724,N_15470,N_15312);
nand U15725 (N_15725,N_15340,N_15389);
xor U15726 (N_15726,N_15342,N_15366);
nand U15727 (N_15727,N_15329,N_15260);
or U15728 (N_15728,N_15273,N_15456);
nor U15729 (N_15729,N_15387,N_15360);
and U15730 (N_15730,N_15307,N_15335);
and U15731 (N_15731,N_15320,N_15319);
xor U15732 (N_15732,N_15401,N_15387);
xor U15733 (N_15733,N_15290,N_15484);
and U15734 (N_15734,N_15452,N_15471);
xnor U15735 (N_15735,N_15446,N_15324);
and U15736 (N_15736,N_15287,N_15385);
nor U15737 (N_15737,N_15432,N_15411);
nand U15738 (N_15738,N_15259,N_15491);
nor U15739 (N_15739,N_15349,N_15480);
xnor U15740 (N_15740,N_15467,N_15417);
and U15741 (N_15741,N_15434,N_15405);
or U15742 (N_15742,N_15319,N_15365);
or U15743 (N_15743,N_15429,N_15410);
nor U15744 (N_15744,N_15330,N_15321);
or U15745 (N_15745,N_15355,N_15318);
nand U15746 (N_15746,N_15339,N_15316);
or U15747 (N_15747,N_15346,N_15317);
nor U15748 (N_15748,N_15319,N_15490);
nand U15749 (N_15749,N_15282,N_15254);
nand U15750 (N_15750,N_15534,N_15595);
nor U15751 (N_15751,N_15728,N_15618);
and U15752 (N_15752,N_15518,N_15690);
nand U15753 (N_15753,N_15571,N_15606);
or U15754 (N_15754,N_15604,N_15747);
and U15755 (N_15755,N_15637,N_15726);
or U15756 (N_15756,N_15636,N_15742);
and U15757 (N_15757,N_15663,N_15525);
nand U15758 (N_15758,N_15650,N_15695);
and U15759 (N_15759,N_15531,N_15649);
or U15760 (N_15760,N_15641,N_15546);
xor U15761 (N_15761,N_15706,N_15743);
nand U15762 (N_15762,N_15514,N_15608);
nand U15763 (N_15763,N_15738,N_15727);
nor U15764 (N_15764,N_15607,N_15699);
xor U15765 (N_15765,N_15657,N_15533);
or U15766 (N_15766,N_15528,N_15716);
or U15767 (N_15767,N_15745,N_15611);
nor U15768 (N_15768,N_15577,N_15715);
or U15769 (N_15769,N_15732,N_15537);
and U15770 (N_15770,N_15741,N_15562);
nand U15771 (N_15771,N_15516,N_15730);
or U15772 (N_15772,N_15720,N_15513);
nor U15773 (N_15773,N_15683,N_15713);
nand U15774 (N_15774,N_15541,N_15647);
or U15775 (N_15775,N_15620,N_15504);
xnor U15776 (N_15776,N_15521,N_15666);
xor U15777 (N_15777,N_15687,N_15576);
nand U15778 (N_15778,N_15555,N_15633);
xor U15779 (N_15779,N_15526,N_15621);
and U15780 (N_15780,N_15554,N_15685);
or U15781 (N_15781,N_15565,N_15547);
and U15782 (N_15782,N_15567,N_15627);
and U15783 (N_15783,N_15731,N_15655);
nand U15784 (N_15784,N_15586,N_15639);
nor U15785 (N_15785,N_15563,N_15740);
nor U15786 (N_15786,N_15501,N_15626);
and U15787 (N_15787,N_15517,N_15509);
and U15788 (N_15788,N_15572,N_15550);
nor U15789 (N_15789,N_15612,N_15671);
or U15790 (N_15790,N_15506,N_15700);
or U15791 (N_15791,N_15508,N_15545);
or U15792 (N_15792,N_15592,N_15566);
nand U15793 (N_15793,N_15662,N_15529);
or U15794 (N_15794,N_15574,N_15634);
or U15795 (N_15795,N_15638,N_15603);
xor U15796 (N_15796,N_15629,N_15654);
or U15797 (N_15797,N_15581,N_15693);
and U15798 (N_15798,N_15536,N_15552);
nand U15799 (N_15799,N_15669,N_15510);
xor U15800 (N_15800,N_15703,N_15519);
nand U15801 (N_15801,N_15575,N_15553);
and U15802 (N_15802,N_15615,N_15587);
nor U15803 (N_15803,N_15594,N_15622);
xnor U15804 (N_15804,N_15535,N_15591);
xnor U15805 (N_15805,N_15551,N_15719);
and U15806 (N_15806,N_15590,N_15659);
and U15807 (N_15807,N_15646,N_15648);
xnor U15808 (N_15808,N_15684,N_15540);
nand U15809 (N_15809,N_15681,N_15569);
xnor U15810 (N_15810,N_15734,N_15682);
nor U15811 (N_15811,N_15714,N_15630);
nor U15812 (N_15812,N_15675,N_15711);
nand U15813 (N_15813,N_15524,N_15670);
nor U15814 (N_15814,N_15696,N_15692);
and U15815 (N_15815,N_15511,N_15739);
nor U15816 (N_15816,N_15705,N_15527);
nand U15817 (N_15817,N_15721,N_15593);
or U15818 (N_15818,N_15661,N_15584);
nand U15819 (N_15819,N_15616,N_15619);
nor U15820 (N_15820,N_15694,N_15532);
and U15821 (N_15821,N_15676,N_15631);
xnor U15822 (N_15822,N_15688,N_15539);
nand U15823 (N_15823,N_15725,N_15617);
nand U15824 (N_15824,N_15523,N_15573);
and U15825 (N_15825,N_15582,N_15672);
and U15826 (N_15826,N_15733,N_15689);
nand U15827 (N_15827,N_15673,N_15707);
and U15828 (N_15828,N_15512,N_15602);
nor U15829 (N_15829,N_15579,N_15644);
or U15830 (N_15830,N_15500,N_15601);
nand U15831 (N_15831,N_15667,N_15642);
xnor U15832 (N_15832,N_15645,N_15588);
or U15833 (N_15833,N_15589,N_15656);
nand U15834 (N_15834,N_15718,N_15598);
and U15835 (N_15835,N_15624,N_15580);
xor U15836 (N_15836,N_15559,N_15680);
or U15837 (N_15837,N_15708,N_15709);
or U15838 (N_15838,N_15724,N_15691);
or U15839 (N_15839,N_15674,N_15564);
or U15840 (N_15840,N_15686,N_15640);
nor U15841 (N_15841,N_15505,N_15613);
nand U15842 (N_15842,N_15600,N_15522);
nand U15843 (N_15843,N_15729,N_15749);
nand U15844 (N_15844,N_15548,N_15678);
nand U15845 (N_15845,N_15614,N_15543);
and U15846 (N_15846,N_15549,N_15717);
xnor U15847 (N_15847,N_15568,N_15651);
and U15848 (N_15848,N_15643,N_15596);
nand U15849 (N_15849,N_15625,N_15599);
xnor U15850 (N_15850,N_15710,N_15570);
xor U15851 (N_15851,N_15544,N_15558);
nand U15852 (N_15852,N_15701,N_15585);
nor U15853 (N_15853,N_15556,N_15583);
nor U15854 (N_15854,N_15538,N_15609);
xnor U15855 (N_15855,N_15723,N_15578);
or U15856 (N_15856,N_15665,N_15704);
xor U15857 (N_15857,N_15560,N_15597);
nand U15858 (N_15858,N_15744,N_15698);
xor U15859 (N_15859,N_15520,N_15530);
and U15860 (N_15860,N_15679,N_15735);
nor U15861 (N_15861,N_15610,N_15658);
or U15862 (N_15862,N_15722,N_15628);
xor U15863 (N_15863,N_15502,N_15737);
nand U15864 (N_15864,N_15668,N_15632);
xnor U15865 (N_15865,N_15653,N_15660);
nand U15866 (N_15866,N_15677,N_15557);
or U15867 (N_15867,N_15635,N_15702);
nor U15868 (N_15868,N_15503,N_15697);
or U15869 (N_15869,N_15623,N_15664);
nor U15870 (N_15870,N_15746,N_15605);
and U15871 (N_15871,N_15515,N_15748);
nor U15872 (N_15872,N_15542,N_15561);
nor U15873 (N_15873,N_15712,N_15507);
or U15874 (N_15874,N_15736,N_15652);
nor U15875 (N_15875,N_15543,N_15650);
xor U15876 (N_15876,N_15731,N_15638);
and U15877 (N_15877,N_15549,N_15735);
and U15878 (N_15878,N_15622,N_15537);
or U15879 (N_15879,N_15674,N_15535);
nor U15880 (N_15880,N_15695,N_15615);
nor U15881 (N_15881,N_15681,N_15604);
xor U15882 (N_15882,N_15595,N_15687);
xor U15883 (N_15883,N_15668,N_15516);
nand U15884 (N_15884,N_15748,N_15625);
or U15885 (N_15885,N_15541,N_15671);
nand U15886 (N_15886,N_15730,N_15696);
nand U15887 (N_15887,N_15625,N_15718);
nor U15888 (N_15888,N_15679,N_15687);
or U15889 (N_15889,N_15689,N_15704);
xor U15890 (N_15890,N_15745,N_15562);
or U15891 (N_15891,N_15615,N_15654);
xor U15892 (N_15892,N_15554,N_15513);
nand U15893 (N_15893,N_15601,N_15603);
nor U15894 (N_15894,N_15585,N_15511);
and U15895 (N_15895,N_15639,N_15558);
nor U15896 (N_15896,N_15715,N_15639);
nor U15897 (N_15897,N_15745,N_15546);
xnor U15898 (N_15898,N_15552,N_15528);
and U15899 (N_15899,N_15541,N_15702);
or U15900 (N_15900,N_15643,N_15592);
nand U15901 (N_15901,N_15611,N_15647);
or U15902 (N_15902,N_15579,N_15659);
xor U15903 (N_15903,N_15551,N_15728);
nand U15904 (N_15904,N_15514,N_15699);
xor U15905 (N_15905,N_15676,N_15652);
and U15906 (N_15906,N_15658,N_15521);
or U15907 (N_15907,N_15709,N_15591);
nor U15908 (N_15908,N_15612,N_15709);
xor U15909 (N_15909,N_15567,N_15580);
nand U15910 (N_15910,N_15608,N_15647);
nor U15911 (N_15911,N_15687,N_15585);
xnor U15912 (N_15912,N_15642,N_15717);
or U15913 (N_15913,N_15581,N_15500);
xor U15914 (N_15914,N_15528,N_15581);
and U15915 (N_15915,N_15572,N_15693);
xor U15916 (N_15916,N_15612,N_15573);
xor U15917 (N_15917,N_15557,N_15529);
nor U15918 (N_15918,N_15617,N_15530);
xor U15919 (N_15919,N_15538,N_15588);
nor U15920 (N_15920,N_15610,N_15556);
and U15921 (N_15921,N_15543,N_15740);
nor U15922 (N_15922,N_15605,N_15649);
nor U15923 (N_15923,N_15711,N_15672);
xnor U15924 (N_15924,N_15553,N_15540);
xnor U15925 (N_15925,N_15620,N_15733);
nor U15926 (N_15926,N_15558,N_15566);
and U15927 (N_15927,N_15509,N_15580);
nand U15928 (N_15928,N_15596,N_15532);
xnor U15929 (N_15929,N_15683,N_15531);
nand U15930 (N_15930,N_15657,N_15623);
xnor U15931 (N_15931,N_15706,N_15523);
and U15932 (N_15932,N_15719,N_15685);
nor U15933 (N_15933,N_15705,N_15639);
nor U15934 (N_15934,N_15591,N_15558);
xor U15935 (N_15935,N_15536,N_15641);
xor U15936 (N_15936,N_15675,N_15569);
nand U15937 (N_15937,N_15516,N_15688);
nand U15938 (N_15938,N_15596,N_15633);
nand U15939 (N_15939,N_15626,N_15534);
or U15940 (N_15940,N_15548,N_15658);
and U15941 (N_15941,N_15635,N_15608);
nor U15942 (N_15942,N_15689,N_15519);
xor U15943 (N_15943,N_15577,N_15603);
and U15944 (N_15944,N_15639,N_15701);
nand U15945 (N_15945,N_15634,N_15619);
nor U15946 (N_15946,N_15563,N_15608);
nand U15947 (N_15947,N_15585,N_15597);
and U15948 (N_15948,N_15731,N_15707);
nand U15949 (N_15949,N_15665,N_15554);
or U15950 (N_15950,N_15673,N_15655);
nand U15951 (N_15951,N_15694,N_15731);
nor U15952 (N_15952,N_15521,N_15581);
and U15953 (N_15953,N_15728,N_15576);
or U15954 (N_15954,N_15569,N_15608);
xor U15955 (N_15955,N_15579,N_15551);
nor U15956 (N_15956,N_15597,N_15686);
nor U15957 (N_15957,N_15553,N_15547);
and U15958 (N_15958,N_15728,N_15714);
xor U15959 (N_15959,N_15702,N_15587);
or U15960 (N_15960,N_15521,N_15673);
nor U15961 (N_15961,N_15634,N_15662);
nand U15962 (N_15962,N_15550,N_15747);
nor U15963 (N_15963,N_15645,N_15566);
xnor U15964 (N_15964,N_15528,N_15597);
and U15965 (N_15965,N_15615,N_15742);
xnor U15966 (N_15966,N_15719,N_15697);
or U15967 (N_15967,N_15573,N_15600);
nor U15968 (N_15968,N_15695,N_15584);
xnor U15969 (N_15969,N_15569,N_15692);
xnor U15970 (N_15970,N_15520,N_15735);
or U15971 (N_15971,N_15548,N_15597);
nor U15972 (N_15972,N_15747,N_15507);
nand U15973 (N_15973,N_15506,N_15680);
nor U15974 (N_15974,N_15747,N_15566);
xor U15975 (N_15975,N_15641,N_15595);
and U15976 (N_15976,N_15611,N_15559);
and U15977 (N_15977,N_15736,N_15562);
nand U15978 (N_15978,N_15718,N_15590);
and U15979 (N_15979,N_15527,N_15610);
or U15980 (N_15980,N_15686,N_15735);
nor U15981 (N_15981,N_15560,N_15641);
xnor U15982 (N_15982,N_15667,N_15590);
nand U15983 (N_15983,N_15509,N_15691);
and U15984 (N_15984,N_15716,N_15606);
and U15985 (N_15985,N_15538,N_15685);
or U15986 (N_15986,N_15505,N_15513);
or U15987 (N_15987,N_15545,N_15586);
and U15988 (N_15988,N_15689,N_15702);
nor U15989 (N_15989,N_15661,N_15629);
and U15990 (N_15990,N_15532,N_15626);
and U15991 (N_15991,N_15585,N_15742);
nand U15992 (N_15992,N_15638,N_15630);
and U15993 (N_15993,N_15588,N_15647);
nor U15994 (N_15994,N_15674,N_15529);
and U15995 (N_15995,N_15615,N_15566);
or U15996 (N_15996,N_15713,N_15581);
and U15997 (N_15997,N_15737,N_15559);
nand U15998 (N_15998,N_15698,N_15511);
xor U15999 (N_15999,N_15589,N_15644);
and U16000 (N_16000,N_15864,N_15993);
and U16001 (N_16001,N_15770,N_15807);
nor U16002 (N_16002,N_15900,N_15781);
nor U16003 (N_16003,N_15950,N_15765);
xor U16004 (N_16004,N_15788,N_15888);
nor U16005 (N_16005,N_15951,N_15894);
nor U16006 (N_16006,N_15969,N_15805);
and U16007 (N_16007,N_15970,N_15871);
and U16008 (N_16008,N_15922,N_15972);
xor U16009 (N_16009,N_15790,N_15806);
or U16010 (N_16010,N_15898,N_15776);
or U16011 (N_16011,N_15913,N_15884);
or U16012 (N_16012,N_15930,N_15800);
and U16013 (N_16013,N_15985,N_15809);
and U16014 (N_16014,N_15932,N_15971);
or U16015 (N_16015,N_15840,N_15846);
xor U16016 (N_16016,N_15915,N_15837);
or U16017 (N_16017,N_15940,N_15937);
nand U16018 (N_16018,N_15895,N_15870);
or U16019 (N_16019,N_15750,N_15916);
xnor U16020 (N_16020,N_15810,N_15883);
nand U16021 (N_16021,N_15908,N_15826);
and U16022 (N_16022,N_15816,N_15803);
and U16023 (N_16023,N_15785,N_15987);
or U16024 (N_16024,N_15757,N_15962);
xnor U16025 (N_16025,N_15943,N_15760);
xnor U16026 (N_16026,N_15899,N_15821);
xnor U16027 (N_16027,N_15959,N_15897);
or U16028 (N_16028,N_15945,N_15933);
nand U16029 (N_16029,N_15861,N_15793);
xnor U16030 (N_16030,N_15820,N_15801);
nand U16031 (N_16031,N_15852,N_15762);
and U16032 (N_16032,N_15795,N_15983);
nor U16033 (N_16033,N_15818,N_15956);
nor U16034 (N_16034,N_15882,N_15904);
xor U16035 (N_16035,N_15841,N_15981);
xnor U16036 (N_16036,N_15968,N_15921);
nand U16037 (N_16037,N_15942,N_15850);
nor U16038 (N_16038,N_15887,N_15825);
xnor U16039 (N_16039,N_15823,N_15768);
and U16040 (N_16040,N_15880,N_15999);
xnor U16041 (N_16041,N_15980,N_15901);
or U16042 (N_16042,N_15812,N_15777);
xnor U16043 (N_16043,N_15892,N_15960);
nand U16044 (N_16044,N_15996,N_15862);
xor U16045 (N_16045,N_15890,N_15856);
nor U16046 (N_16046,N_15799,N_15958);
or U16047 (N_16047,N_15863,N_15831);
and U16048 (N_16048,N_15752,N_15911);
xnor U16049 (N_16049,N_15905,N_15934);
nor U16050 (N_16050,N_15859,N_15941);
or U16051 (N_16051,N_15961,N_15796);
nor U16052 (N_16052,N_15875,N_15804);
xor U16053 (N_16053,N_15995,N_15784);
nand U16054 (N_16054,N_15955,N_15789);
nand U16055 (N_16055,N_15952,N_15792);
and U16056 (N_16056,N_15833,N_15967);
nor U16057 (N_16057,N_15978,N_15866);
or U16058 (N_16058,N_15872,N_15885);
nand U16059 (N_16059,N_15949,N_15979);
nand U16060 (N_16060,N_15926,N_15988);
xor U16061 (N_16061,N_15773,N_15822);
and U16062 (N_16062,N_15923,N_15779);
or U16063 (N_16063,N_15798,N_15868);
nor U16064 (N_16064,N_15860,N_15819);
xor U16065 (N_16065,N_15977,N_15997);
xor U16066 (N_16066,N_15891,N_15836);
and U16067 (N_16067,N_15853,N_15865);
or U16068 (N_16068,N_15858,N_15857);
xnor U16069 (N_16069,N_15756,N_15827);
and U16070 (N_16070,N_15964,N_15838);
and U16071 (N_16071,N_15808,N_15973);
xor U16072 (N_16072,N_15954,N_15786);
nand U16073 (N_16073,N_15953,N_15912);
or U16074 (N_16074,N_15948,N_15925);
or U16075 (N_16075,N_15855,N_15813);
nor U16076 (N_16076,N_15842,N_15817);
and U16077 (N_16077,N_15910,N_15767);
nor U16078 (N_16078,N_15989,N_15766);
or U16079 (N_16079,N_15917,N_15966);
and U16080 (N_16080,N_15787,N_15751);
and U16081 (N_16081,N_15893,N_15938);
nand U16082 (N_16082,N_15778,N_15909);
nor U16083 (N_16083,N_15919,N_15902);
xnor U16084 (N_16084,N_15811,N_15944);
or U16085 (N_16085,N_15845,N_15758);
nor U16086 (N_16086,N_15876,N_15772);
xor U16087 (N_16087,N_15947,N_15994);
or U16088 (N_16088,N_15931,N_15889);
nand U16089 (N_16089,N_15918,N_15847);
xnor U16090 (N_16090,N_15843,N_15984);
nor U16091 (N_16091,N_15764,N_15939);
nor U16092 (N_16092,N_15783,N_15769);
xor U16093 (N_16093,N_15755,N_15975);
nor U16094 (N_16094,N_15903,N_15771);
and U16095 (N_16095,N_15946,N_15832);
and U16096 (N_16096,N_15879,N_15814);
or U16097 (N_16097,N_15754,N_15867);
nor U16098 (N_16098,N_15802,N_15896);
nor U16099 (N_16099,N_15869,N_15775);
and U16100 (N_16100,N_15834,N_15844);
nor U16101 (N_16101,N_15936,N_15774);
nand U16102 (N_16102,N_15824,N_15974);
and U16103 (N_16103,N_15986,N_15914);
and U16104 (N_16104,N_15835,N_15992);
nand U16105 (N_16105,N_15957,N_15763);
xnor U16106 (N_16106,N_15851,N_15920);
nor U16107 (N_16107,N_15907,N_15991);
nor U16108 (N_16108,N_15854,N_15759);
nand U16109 (N_16109,N_15839,N_15849);
nand U16110 (N_16110,N_15906,N_15881);
nand U16111 (N_16111,N_15927,N_15815);
and U16112 (N_16112,N_15965,N_15886);
nor U16113 (N_16113,N_15782,N_15998);
or U16114 (N_16114,N_15829,N_15828);
xor U16115 (N_16115,N_15753,N_15982);
xnor U16116 (N_16116,N_15877,N_15990);
nor U16117 (N_16117,N_15976,N_15929);
xnor U16118 (N_16118,N_15830,N_15874);
nor U16119 (N_16119,N_15794,N_15780);
nor U16120 (N_16120,N_15963,N_15935);
nand U16121 (N_16121,N_15761,N_15878);
or U16122 (N_16122,N_15924,N_15848);
nand U16123 (N_16123,N_15928,N_15791);
or U16124 (N_16124,N_15873,N_15797);
nor U16125 (N_16125,N_15774,N_15781);
nor U16126 (N_16126,N_15945,N_15815);
or U16127 (N_16127,N_15987,N_15811);
and U16128 (N_16128,N_15962,N_15932);
nor U16129 (N_16129,N_15995,N_15899);
nand U16130 (N_16130,N_15824,N_15987);
or U16131 (N_16131,N_15967,N_15861);
xor U16132 (N_16132,N_15908,N_15804);
nand U16133 (N_16133,N_15813,N_15911);
nand U16134 (N_16134,N_15958,N_15977);
nand U16135 (N_16135,N_15953,N_15899);
xnor U16136 (N_16136,N_15870,N_15975);
and U16137 (N_16137,N_15981,N_15805);
nand U16138 (N_16138,N_15917,N_15899);
or U16139 (N_16139,N_15928,N_15770);
or U16140 (N_16140,N_15830,N_15903);
and U16141 (N_16141,N_15762,N_15782);
and U16142 (N_16142,N_15803,N_15798);
nand U16143 (N_16143,N_15857,N_15846);
or U16144 (N_16144,N_15836,N_15872);
nand U16145 (N_16145,N_15765,N_15935);
nor U16146 (N_16146,N_15907,N_15866);
and U16147 (N_16147,N_15962,N_15939);
and U16148 (N_16148,N_15993,N_15773);
or U16149 (N_16149,N_15989,N_15800);
nand U16150 (N_16150,N_15860,N_15778);
and U16151 (N_16151,N_15757,N_15780);
nor U16152 (N_16152,N_15875,N_15884);
or U16153 (N_16153,N_15752,N_15893);
and U16154 (N_16154,N_15897,N_15912);
xnor U16155 (N_16155,N_15794,N_15753);
and U16156 (N_16156,N_15972,N_15887);
nor U16157 (N_16157,N_15771,N_15940);
and U16158 (N_16158,N_15806,N_15816);
and U16159 (N_16159,N_15856,N_15977);
nor U16160 (N_16160,N_15843,N_15941);
xnor U16161 (N_16161,N_15816,N_15939);
or U16162 (N_16162,N_15966,N_15914);
xnor U16163 (N_16163,N_15840,N_15960);
nand U16164 (N_16164,N_15752,N_15995);
and U16165 (N_16165,N_15779,N_15752);
and U16166 (N_16166,N_15910,N_15996);
or U16167 (N_16167,N_15888,N_15967);
xor U16168 (N_16168,N_15796,N_15927);
xor U16169 (N_16169,N_15814,N_15860);
and U16170 (N_16170,N_15887,N_15776);
nand U16171 (N_16171,N_15930,N_15891);
or U16172 (N_16172,N_15968,N_15970);
xnor U16173 (N_16173,N_15904,N_15897);
or U16174 (N_16174,N_15877,N_15947);
nand U16175 (N_16175,N_15841,N_15848);
and U16176 (N_16176,N_15974,N_15780);
or U16177 (N_16177,N_15783,N_15849);
or U16178 (N_16178,N_15913,N_15798);
and U16179 (N_16179,N_15767,N_15930);
and U16180 (N_16180,N_15855,N_15945);
nand U16181 (N_16181,N_15967,N_15912);
and U16182 (N_16182,N_15985,N_15932);
and U16183 (N_16183,N_15770,N_15870);
nor U16184 (N_16184,N_15751,N_15794);
nand U16185 (N_16185,N_15786,N_15850);
xor U16186 (N_16186,N_15784,N_15983);
nand U16187 (N_16187,N_15797,N_15997);
nand U16188 (N_16188,N_15810,N_15824);
and U16189 (N_16189,N_15808,N_15797);
nand U16190 (N_16190,N_15818,N_15869);
and U16191 (N_16191,N_15906,N_15853);
and U16192 (N_16192,N_15864,N_15926);
and U16193 (N_16193,N_15810,N_15815);
or U16194 (N_16194,N_15809,N_15973);
nand U16195 (N_16195,N_15814,N_15812);
or U16196 (N_16196,N_15895,N_15876);
nand U16197 (N_16197,N_15752,N_15889);
or U16198 (N_16198,N_15822,N_15936);
xor U16199 (N_16199,N_15921,N_15790);
xor U16200 (N_16200,N_15795,N_15945);
xor U16201 (N_16201,N_15925,N_15858);
xor U16202 (N_16202,N_15752,N_15912);
nand U16203 (N_16203,N_15825,N_15867);
and U16204 (N_16204,N_15825,N_15790);
and U16205 (N_16205,N_15804,N_15753);
or U16206 (N_16206,N_15797,N_15755);
and U16207 (N_16207,N_15807,N_15986);
and U16208 (N_16208,N_15879,N_15905);
and U16209 (N_16209,N_15832,N_15926);
xnor U16210 (N_16210,N_15861,N_15937);
nand U16211 (N_16211,N_15769,N_15958);
and U16212 (N_16212,N_15815,N_15819);
nand U16213 (N_16213,N_15857,N_15954);
or U16214 (N_16214,N_15977,N_15986);
xor U16215 (N_16215,N_15803,N_15791);
nor U16216 (N_16216,N_15928,N_15837);
or U16217 (N_16217,N_15970,N_15999);
xnor U16218 (N_16218,N_15975,N_15938);
or U16219 (N_16219,N_15765,N_15842);
or U16220 (N_16220,N_15911,N_15980);
nor U16221 (N_16221,N_15888,N_15957);
xnor U16222 (N_16222,N_15968,N_15907);
nor U16223 (N_16223,N_15809,N_15918);
nand U16224 (N_16224,N_15791,N_15756);
nor U16225 (N_16225,N_15894,N_15869);
or U16226 (N_16226,N_15751,N_15819);
or U16227 (N_16227,N_15889,N_15784);
nand U16228 (N_16228,N_15810,N_15878);
nor U16229 (N_16229,N_15942,N_15797);
nand U16230 (N_16230,N_15904,N_15786);
and U16231 (N_16231,N_15787,N_15763);
nand U16232 (N_16232,N_15760,N_15807);
nor U16233 (N_16233,N_15915,N_15761);
xnor U16234 (N_16234,N_15831,N_15767);
xor U16235 (N_16235,N_15817,N_15874);
xor U16236 (N_16236,N_15895,N_15753);
or U16237 (N_16237,N_15766,N_15968);
and U16238 (N_16238,N_15803,N_15821);
or U16239 (N_16239,N_15859,N_15794);
and U16240 (N_16240,N_15891,N_15811);
nand U16241 (N_16241,N_15884,N_15827);
xnor U16242 (N_16242,N_15800,N_15857);
nor U16243 (N_16243,N_15767,N_15751);
nor U16244 (N_16244,N_15985,N_15962);
nor U16245 (N_16245,N_15784,N_15870);
xnor U16246 (N_16246,N_15990,N_15872);
nand U16247 (N_16247,N_15935,N_15902);
or U16248 (N_16248,N_15889,N_15952);
or U16249 (N_16249,N_15752,N_15799);
nor U16250 (N_16250,N_16175,N_16021);
xor U16251 (N_16251,N_16094,N_16138);
nor U16252 (N_16252,N_16073,N_16056);
xnor U16253 (N_16253,N_16212,N_16211);
xor U16254 (N_16254,N_16144,N_16182);
or U16255 (N_16255,N_16154,N_16107);
nand U16256 (N_16256,N_16204,N_16024);
xnor U16257 (N_16257,N_16159,N_16193);
xnor U16258 (N_16258,N_16033,N_16026);
and U16259 (N_16259,N_16040,N_16028);
nand U16260 (N_16260,N_16219,N_16174);
nand U16261 (N_16261,N_16049,N_16222);
and U16262 (N_16262,N_16196,N_16228);
nor U16263 (N_16263,N_16106,N_16079);
xnor U16264 (N_16264,N_16080,N_16189);
nand U16265 (N_16265,N_16194,N_16157);
nand U16266 (N_16266,N_16085,N_16229);
nand U16267 (N_16267,N_16132,N_16075);
nand U16268 (N_16268,N_16035,N_16198);
xnor U16269 (N_16269,N_16156,N_16060);
nand U16270 (N_16270,N_16004,N_16202);
nand U16271 (N_16271,N_16062,N_16235);
or U16272 (N_16272,N_16238,N_16183);
xnor U16273 (N_16273,N_16045,N_16249);
nor U16274 (N_16274,N_16129,N_16244);
xor U16275 (N_16275,N_16239,N_16207);
nor U16276 (N_16276,N_16008,N_16109);
nand U16277 (N_16277,N_16065,N_16227);
nand U16278 (N_16278,N_16027,N_16037);
or U16279 (N_16279,N_16124,N_16052);
xor U16280 (N_16280,N_16043,N_16117);
or U16281 (N_16281,N_16181,N_16000);
and U16282 (N_16282,N_16215,N_16187);
or U16283 (N_16283,N_16084,N_16083);
nor U16284 (N_16284,N_16150,N_16230);
and U16285 (N_16285,N_16088,N_16180);
and U16286 (N_16286,N_16039,N_16050);
nand U16287 (N_16287,N_16218,N_16205);
and U16288 (N_16288,N_16128,N_16126);
nor U16289 (N_16289,N_16010,N_16170);
or U16290 (N_16290,N_16165,N_16018);
and U16291 (N_16291,N_16042,N_16122);
xnor U16292 (N_16292,N_16208,N_16192);
xor U16293 (N_16293,N_16007,N_16153);
nor U16294 (N_16294,N_16086,N_16070);
or U16295 (N_16295,N_16186,N_16237);
xor U16296 (N_16296,N_16140,N_16214);
nand U16297 (N_16297,N_16006,N_16044);
and U16298 (N_16298,N_16179,N_16223);
xor U16299 (N_16299,N_16188,N_16016);
and U16300 (N_16300,N_16099,N_16226);
nor U16301 (N_16301,N_16151,N_16178);
nand U16302 (N_16302,N_16234,N_16142);
and U16303 (N_16303,N_16118,N_16091);
nor U16304 (N_16304,N_16082,N_16096);
xor U16305 (N_16305,N_16092,N_16145);
and U16306 (N_16306,N_16093,N_16169);
nor U16307 (N_16307,N_16216,N_16184);
and U16308 (N_16308,N_16095,N_16071);
xor U16309 (N_16309,N_16020,N_16241);
or U16310 (N_16310,N_16161,N_16197);
or U16311 (N_16311,N_16200,N_16149);
xor U16312 (N_16312,N_16139,N_16097);
xor U16313 (N_16313,N_16111,N_16101);
and U16314 (N_16314,N_16199,N_16100);
nand U16315 (N_16315,N_16248,N_16034);
nor U16316 (N_16316,N_16038,N_16233);
nand U16317 (N_16317,N_16110,N_16209);
and U16318 (N_16318,N_16242,N_16134);
or U16319 (N_16319,N_16177,N_16090);
xnor U16320 (N_16320,N_16166,N_16172);
xnor U16321 (N_16321,N_16001,N_16046);
nand U16322 (N_16322,N_16114,N_16168);
and U16323 (N_16323,N_16176,N_16002);
or U16324 (N_16324,N_16123,N_16055);
and U16325 (N_16325,N_16057,N_16011);
nor U16326 (N_16326,N_16120,N_16143);
xnor U16327 (N_16327,N_16069,N_16243);
and U16328 (N_16328,N_16108,N_16031);
or U16329 (N_16329,N_16068,N_16081);
nand U16330 (N_16330,N_16190,N_16032);
or U16331 (N_16331,N_16136,N_16163);
nor U16332 (N_16332,N_16224,N_16063);
and U16333 (N_16333,N_16012,N_16147);
or U16334 (N_16334,N_16148,N_16047);
nand U16335 (N_16335,N_16051,N_16029);
xnor U16336 (N_16336,N_16041,N_16087);
or U16337 (N_16337,N_16158,N_16206);
xnor U16338 (N_16338,N_16155,N_16231);
and U16339 (N_16339,N_16022,N_16221);
nand U16340 (N_16340,N_16210,N_16173);
xor U16341 (N_16341,N_16162,N_16059);
nand U16342 (N_16342,N_16003,N_16217);
nand U16343 (N_16343,N_16025,N_16121);
or U16344 (N_16344,N_16125,N_16135);
or U16345 (N_16345,N_16067,N_16089);
nand U16346 (N_16346,N_16246,N_16064);
and U16347 (N_16347,N_16076,N_16103);
xor U16348 (N_16348,N_16017,N_16164);
and U16349 (N_16349,N_16171,N_16232);
or U16350 (N_16350,N_16146,N_16201);
or U16351 (N_16351,N_16131,N_16009);
nand U16352 (N_16352,N_16116,N_16061);
and U16353 (N_16353,N_16113,N_16058);
and U16354 (N_16354,N_16098,N_16074);
nor U16355 (N_16355,N_16072,N_16112);
xnor U16356 (N_16356,N_16225,N_16127);
nor U16357 (N_16357,N_16141,N_16245);
and U16358 (N_16358,N_16220,N_16048);
nand U16359 (N_16359,N_16133,N_16130);
xor U16360 (N_16360,N_16213,N_16240);
nor U16361 (N_16361,N_16236,N_16054);
xor U16362 (N_16362,N_16203,N_16167);
or U16363 (N_16363,N_16104,N_16160);
and U16364 (N_16364,N_16105,N_16030);
nand U16365 (N_16365,N_16019,N_16115);
nand U16366 (N_16366,N_16015,N_16247);
nand U16367 (N_16367,N_16191,N_16078);
xnor U16368 (N_16368,N_16053,N_16077);
and U16369 (N_16369,N_16119,N_16102);
and U16370 (N_16370,N_16185,N_16013);
or U16371 (N_16371,N_16014,N_16195);
nor U16372 (N_16372,N_16005,N_16152);
or U16373 (N_16373,N_16023,N_16137);
nand U16374 (N_16374,N_16036,N_16066);
and U16375 (N_16375,N_16008,N_16037);
nand U16376 (N_16376,N_16068,N_16235);
or U16377 (N_16377,N_16234,N_16055);
xnor U16378 (N_16378,N_16216,N_16010);
or U16379 (N_16379,N_16145,N_16099);
xor U16380 (N_16380,N_16016,N_16212);
nand U16381 (N_16381,N_16044,N_16144);
or U16382 (N_16382,N_16120,N_16169);
xnor U16383 (N_16383,N_16160,N_16137);
and U16384 (N_16384,N_16113,N_16010);
or U16385 (N_16385,N_16182,N_16084);
nor U16386 (N_16386,N_16085,N_16093);
and U16387 (N_16387,N_16049,N_16043);
and U16388 (N_16388,N_16228,N_16188);
nand U16389 (N_16389,N_16054,N_16099);
xor U16390 (N_16390,N_16043,N_16031);
xor U16391 (N_16391,N_16049,N_16111);
nor U16392 (N_16392,N_16100,N_16112);
nor U16393 (N_16393,N_16119,N_16087);
and U16394 (N_16394,N_16018,N_16104);
nand U16395 (N_16395,N_16233,N_16244);
nand U16396 (N_16396,N_16083,N_16103);
xnor U16397 (N_16397,N_16229,N_16185);
or U16398 (N_16398,N_16074,N_16148);
or U16399 (N_16399,N_16087,N_16142);
nor U16400 (N_16400,N_16238,N_16045);
xnor U16401 (N_16401,N_16235,N_16118);
nor U16402 (N_16402,N_16149,N_16046);
and U16403 (N_16403,N_16176,N_16017);
nand U16404 (N_16404,N_16212,N_16181);
xnor U16405 (N_16405,N_16116,N_16187);
or U16406 (N_16406,N_16133,N_16026);
or U16407 (N_16407,N_16158,N_16211);
or U16408 (N_16408,N_16082,N_16107);
nor U16409 (N_16409,N_16166,N_16087);
or U16410 (N_16410,N_16103,N_16154);
or U16411 (N_16411,N_16137,N_16116);
xnor U16412 (N_16412,N_16079,N_16007);
and U16413 (N_16413,N_16097,N_16229);
xor U16414 (N_16414,N_16130,N_16194);
or U16415 (N_16415,N_16046,N_16204);
nor U16416 (N_16416,N_16231,N_16103);
nor U16417 (N_16417,N_16082,N_16130);
nor U16418 (N_16418,N_16164,N_16009);
nor U16419 (N_16419,N_16206,N_16095);
and U16420 (N_16420,N_16236,N_16118);
nor U16421 (N_16421,N_16200,N_16021);
xnor U16422 (N_16422,N_16125,N_16136);
xnor U16423 (N_16423,N_16166,N_16008);
nand U16424 (N_16424,N_16000,N_16172);
nor U16425 (N_16425,N_16061,N_16017);
and U16426 (N_16426,N_16162,N_16104);
nor U16427 (N_16427,N_16126,N_16098);
nor U16428 (N_16428,N_16029,N_16213);
nor U16429 (N_16429,N_16186,N_16218);
and U16430 (N_16430,N_16235,N_16225);
nand U16431 (N_16431,N_16167,N_16113);
and U16432 (N_16432,N_16163,N_16238);
xor U16433 (N_16433,N_16135,N_16019);
nor U16434 (N_16434,N_16165,N_16042);
or U16435 (N_16435,N_16055,N_16197);
and U16436 (N_16436,N_16002,N_16147);
or U16437 (N_16437,N_16230,N_16115);
and U16438 (N_16438,N_16167,N_16145);
nor U16439 (N_16439,N_16088,N_16092);
nor U16440 (N_16440,N_16227,N_16082);
or U16441 (N_16441,N_16134,N_16226);
xnor U16442 (N_16442,N_16012,N_16118);
nor U16443 (N_16443,N_16171,N_16226);
nor U16444 (N_16444,N_16069,N_16080);
nor U16445 (N_16445,N_16029,N_16131);
nor U16446 (N_16446,N_16037,N_16088);
xor U16447 (N_16447,N_16199,N_16173);
nand U16448 (N_16448,N_16060,N_16087);
and U16449 (N_16449,N_16125,N_16022);
or U16450 (N_16450,N_16052,N_16136);
and U16451 (N_16451,N_16165,N_16190);
nor U16452 (N_16452,N_16164,N_16072);
nor U16453 (N_16453,N_16107,N_16110);
xnor U16454 (N_16454,N_16090,N_16010);
nor U16455 (N_16455,N_16168,N_16249);
xnor U16456 (N_16456,N_16030,N_16192);
and U16457 (N_16457,N_16222,N_16070);
nor U16458 (N_16458,N_16104,N_16190);
nor U16459 (N_16459,N_16094,N_16089);
or U16460 (N_16460,N_16149,N_16207);
or U16461 (N_16461,N_16161,N_16207);
or U16462 (N_16462,N_16129,N_16056);
nor U16463 (N_16463,N_16005,N_16239);
nor U16464 (N_16464,N_16189,N_16233);
xor U16465 (N_16465,N_16157,N_16013);
nor U16466 (N_16466,N_16107,N_16001);
and U16467 (N_16467,N_16211,N_16021);
nor U16468 (N_16468,N_16139,N_16219);
nor U16469 (N_16469,N_16067,N_16088);
xor U16470 (N_16470,N_16114,N_16194);
xnor U16471 (N_16471,N_16241,N_16004);
and U16472 (N_16472,N_16018,N_16034);
xnor U16473 (N_16473,N_16116,N_16246);
and U16474 (N_16474,N_16200,N_16160);
or U16475 (N_16475,N_16197,N_16034);
nand U16476 (N_16476,N_16086,N_16199);
xnor U16477 (N_16477,N_16036,N_16204);
or U16478 (N_16478,N_16003,N_16043);
and U16479 (N_16479,N_16209,N_16211);
nor U16480 (N_16480,N_16245,N_16050);
and U16481 (N_16481,N_16204,N_16043);
nand U16482 (N_16482,N_16221,N_16086);
xor U16483 (N_16483,N_16142,N_16181);
nor U16484 (N_16484,N_16024,N_16080);
nand U16485 (N_16485,N_16010,N_16055);
and U16486 (N_16486,N_16093,N_16198);
xor U16487 (N_16487,N_16099,N_16223);
nand U16488 (N_16488,N_16030,N_16016);
nor U16489 (N_16489,N_16136,N_16239);
nand U16490 (N_16490,N_16053,N_16097);
and U16491 (N_16491,N_16129,N_16114);
xnor U16492 (N_16492,N_16059,N_16054);
and U16493 (N_16493,N_16042,N_16093);
nor U16494 (N_16494,N_16109,N_16183);
xor U16495 (N_16495,N_16091,N_16085);
xor U16496 (N_16496,N_16144,N_16010);
xnor U16497 (N_16497,N_16072,N_16209);
nor U16498 (N_16498,N_16082,N_16188);
nor U16499 (N_16499,N_16112,N_16001);
nand U16500 (N_16500,N_16458,N_16415);
and U16501 (N_16501,N_16459,N_16352);
and U16502 (N_16502,N_16495,N_16381);
xor U16503 (N_16503,N_16342,N_16369);
xor U16504 (N_16504,N_16480,N_16467);
nor U16505 (N_16505,N_16274,N_16396);
and U16506 (N_16506,N_16377,N_16428);
or U16507 (N_16507,N_16365,N_16367);
and U16508 (N_16508,N_16453,N_16384);
nand U16509 (N_16509,N_16498,N_16491);
and U16510 (N_16510,N_16436,N_16460);
nor U16511 (N_16511,N_16321,N_16486);
and U16512 (N_16512,N_16456,N_16475);
or U16513 (N_16513,N_16464,N_16316);
xnor U16514 (N_16514,N_16253,N_16287);
xnor U16515 (N_16515,N_16499,N_16437);
and U16516 (N_16516,N_16303,N_16344);
and U16517 (N_16517,N_16419,N_16356);
nand U16518 (N_16518,N_16382,N_16266);
and U16519 (N_16519,N_16429,N_16271);
or U16520 (N_16520,N_16434,N_16439);
and U16521 (N_16521,N_16264,N_16331);
nand U16522 (N_16522,N_16442,N_16485);
nor U16523 (N_16523,N_16282,N_16335);
nand U16524 (N_16524,N_16492,N_16490);
xor U16525 (N_16525,N_16279,N_16457);
nand U16526 (N_16526,N_16450,N_16405);
and U16527 (N_16527,N_16354,N_16447);
nand U16528 (N_16528,N_16478,N_16289);
and U16529 (N_16529,N_16257,N_16297);
xor U16530 (N_16530,N_16325,N_16416);
and U16531 (N_16531,N_16443,N_16411);
nand U16532 (N_16532,N_16280,N_16446);
nor U16533 (N_16533,N_16349,N_16433);
nand U16534 (N_16534,N_16291,N_16328);
nand U16535 (N_16535,N_16374,N_16292);
and U16536 (N_16536,N_16472,N_16401);
nor U16537 (N_16537,N_16296,N_16418);
nor U16538 (N_16538,N_16269,N_16340);
or U16539 (N_16539,N_16345,N_16399);
nand U16540 (N_16540,N_16307,N_16281);
or U16541 (N_16541,N_16390,N_16398);
and U16542 (N_16542,N_16394,N_16327);
or U16543 (N_16543,N_16387,N_16406);
and U16544 (N_16544,N_16404,N_16355);
and U16545 (N_16545,N_16422,N_16341);
nand U16546 (N_16546,N_16262,N_16427);
nand U16547 (N_16547,N_16333,N_16273);
nor U16548 (N_16548,N_16337,N_16250);
xor U16549 (N_16549,N_16285,N_16305);
nor U16550 (N_16550,N_16493,N_16421);
nand U16551 (N_16551,N_16484,N_16389);
nand U16552 (N_16552,N_16317,N_16283);
or U16553 (N_16553,N_16376,N_16397);
or U16554 (N_16554,N_16403,N_16330);
xor U16555 (N_16555,N_16483,N_16295);
nand U16556 (N_16556,N_16364,N_16375);
nand U16557 (N_16557,N_16290,N_16255);
or U16558 (N_16558,N_16449,N_16258);
or U16559 (N_16559,N_16420,N_16362);
xor U16560 (N_16560,N_16380,N_16313);
or U16561 (N_16561,N_16251,N_16476);
or U16562 (N_16562,N_16432,N_16276);
nand U16563 (N_16563,N_16310,N_16267);
or U16564 (N_16564,N_16494,N_16407);
and U16565 (N_16565,N_16360,N_16293);
nand U16566 (N_16566,N_16261,N_16254);
nor U16567 (N_16567,N_16431,N_16320);
xor U16568 (N_16568,N_16477,N_16358);
nor U16569 (N_16569,N_16470,N_16496);
and U16570 (N_16570,N_16466,N_16469);
and U16571 (N_16571,N_16277,N_16471);
nand U16572 (N_16572,N_16372,N_16309);
and U16573 (N_16573,N_16417,N_16489);
nand U16574 (N_16574,N_16265,N_16391);
nand U16575 (N_16575,N_16343,N_16497);
and U16576 (N_16576,N_16315,N_16286);
nor U16577 (N_16577,N_16298,N_16423);
nand U16578 (N_16578,N_16346,N_16388);
nor U16579 (N_16579,N_16252,N_16462);
or U16580 (N_16580,N_16339,N_16312);
and U16581 (N_16581,N_16412,N_16357);
nor U16582 (N_16582,N_16332,N_16448);
nor U16583 (N_16583,N_16299,N_16425);
nor U16584 (N_16584,N_16385,N_16474);
and U16585 (N_16585,N_16288,N_16413);
nand U16586 (N_16586,N_16334,N_16366);
xor U16587 (N_16587,N_16392,N_16256);
nand U16588 (N_16588,N_16359,N_16370);
xor U16589 (N_16589,N_16314,N_16426);
xnor U16590 (N_16590,N_16301,N_16414);
nor U16591 (N_16591,N_16302,N_16481);
and U16592 (N_16592,N_16393,N_16259);
and U16593 (N_16593,N_16348,N_16322);
and U16594 (N_16594,N_16378,N_16338);
xor U16595 (N_16595,N_16383,N_16488);
or U16596 (N_16596,N_16260,N_16465);
xor U16597 (N_16597,N_16351,N_16444);
xnor U16598 (N_16598,N_16278,N_16455);
nor U16599 (N_16599,N_16400,N_16440);
nand U16600 (N_16600,N_16371,N_16473);
and U16601 (N_16601,N_16373,N_16402);
or U16602 (N_16602,N_16487,N_16361);
xor U16603 (N_16603,N_16454,N_16445);
nor U16604 (N_16604,N_16294,N_16409);
nor U16605 (N_16605,N_16323,N_16410);
xnor U16606 (N_16606,N_16311,N_16284);
nor U16607 (N_16607,N_16386,N_16368);
or U16608 (N_16608,N_16430,N_16463);
nor U16609 (N_16609,N_16308,N_16326);
nor U16610 (N_16610,N_16461,N_16272);
xor U16611 (N_16611,N_16268,N_16438);
nand U16612 (N_16612,N_16408,N_16318);
or U16613 (N_16613,N_16270,N_16452);
and U16614 (N_16614,N_16324,N_16424);
and U16615 (N_16615,N_16329,N_16275);
and U16616 (N_16616,N_16379,N_16353);
and U16617 (N_16617,N_16347,N_16479);
nand U16618 (N_16618,N_16363,N_16468);
nand U16619 (N_16619,N_16350,N_16435);
nor U16620 (N_16620,N_16441,N_16451);
or U16621 (N_16621,N_16304,N_16395);
nor U16622 (N_16622,N_16482,N_16300);
nand U16623 (N_16623,N_16306,N_16319);
and U16624 (N_16624,N_16336,N_16263);
nand U16625 (N_16625,N_16300,N_16461);
xor U16626 (N_16626,N_16424,N_16443);
nand U16627 (N_16627,N_16399,N_16444);
nor U16628 (N_16628,N_16483,N_16462);
nor U16629 (N_16629,N_16268,N_16376);
nor U16630 (N_16630,N_16309,N_16258);
nor U16631 (N_16631,N_16492,N_16267);
xor U16632 (N_16632,N_16345,N_16321);
nor U16633 (N_16633,N_16294,N_16351);
nand U16634 (N_16634,N_16379,N_16291);
and U16635 (N_16635,N_16491,N_16393);
nor U16636 (N_16636,N_16305,N_16449);
nor U16637 (N_16637,N_16320,N_16339);
xnor U16638 (N_16638,N_16395,N_16449);
and U16639 (N_16639,N_16345,N_16333);
nand U16640 (N_16640,N_16410,N_16494);
and U16641 (N_16641,N_16296,N_16316);
or U16642 (N_16642,N_16457,N_16448);
nand U16643 (N_16643,N_16352,N_16479);
xor U16644 (N_16644,N_16260,N_16308);
xnor U16645 (N_16645,N_16454,N_16385);
or U16646 (N_16646,N_16371,N_16281);
or U16647 (N_16647,N_16302,N_16404);
xor U16648 (N_16648,N_16428,N_16473);
and U16649 (N_16649,N_16301,N_16474);
and U16650 (N_16650,N_16409,N_16436);
nand U16651 (N_16651,N_16416,N_16285);
or U16652 (N_16652,N_16490,N_16323);
nor U16653 (N_16653,N_16291,N_16344);
xnor U16654 (N_16654,N_16372,N_16340);
nor U16655 (N_16655,N_16301,N_16458);
or U16656 (N_16656,N_16364,N_16431);
nand U16657 (N_16657,N_16448,N_16250);
nand U16658 (N_16658,N_16457,N_16330);
nand U16659 (N_16659,N_16330,N_16321);
nand U16660 (N_16660,N_16251,N_16472);
xnor U16661 (N_16661,N_16327,N_16415);
xnor U16662 (N_16662,N_16251,N_16479);
nand U16663 (N_16663,N_16332,N_16441);
and U16664 (N_16664,N_16372,N_16398);
and U16665 (N_16665,N_16415,N_16484);
xnor U16666 (N_16666,N_16422,N_16446);
nand U16667 (N_16667,N_16368,N_16468);
xor U16668 (N_16668,N_16388,N_16429);
or U16669 (N_16669,N_16340,N_16440);
nand U16670 (N_16670,N_16382,N_16471);
nand U16671 (N_16671,N_16425,N_16443);
or U16672 (N_16672,N_16462,N_16414);
or U16673 (N_16673,N_16432,N_16471);
nor U16674 (N_16674,N_16347,N_16337);
nand U16675 (N_16675,N_16442,N_16255);
and U16676 (N_16676,N_16332,N_16391);
nor U16677 (N_16677,N_16302,N_16413);
nand U16678 (N_16678,N_16380,N_16357);
nand U16679 (N_16679,N_16417,N_16339);
xnor U16680 (N_16680,N_16358,N_16278);
or U16681 (N_16681,N_16471,N_16283);
or U16682 (N_16682,N_16410,N_16483);
and U16683 (N_16683,N_16339,N_16460);
xnor U16684 (N_16684,N_16284,N_16293);
or U16685 (N_16685,N_16420,N_16464);
xnor U16686 (N_16686,N_16323,N_16324);
and U16687 (N_16687,N_16269,N_16367);
xnor U16688 (N_16688,N_16430,N_16287);
and U16689 (N_16689,N_16466,N_16304);
xor U16690 (N_16690,N_16317,N_16465);
or U16691 (N_16691,N_16353,N_16411);
and U16692 (N_16692,N_16260,N_16272);
nand U16693 (N_16693,N_16281,N_16365);
or U16694 (N_16694,N_16393,N_16490);
or U16695 (N_16695,N_16386,N_16273);
xor U16696 (N_16696,N_16369,N_16413);
or U16697 (N_16697,N_16391,N_16397);
nor U16698 (N_16698,N_16380,N_16261);
nor U16699 (N_16699,N_16317,N_16444);
nor U16700 (N_16700,N_16468,N_16482);
nor U16701 (N_16701,N_16424,N_16259);
xnor U16702 (N_16702,N_16358,N_16491);
or U16703 (N_16703,N_16277,N_16344);
xnor U16704 (N_16704,N_16306,N_16370);
or U16705 (N_16705,N_16385,N_16325);
or U16706 (N_16706,N_16423,N_16289);
nand U16707 (N_16707,N_16271,N_16495);
xor U16708 (N_16708,N_16310,N_16475);
or U16709 (N_16709,N_16417,N_16395);
nand U16710 (N_16710,N_16372,N_16426);
xor U16711 (N_16711,N_16284,N_16445);
or U16712 (N_16712,N_16406,N_16304);
xnor U16713 (N_16713,N_16385,N_16269);
or U16714 (N_16714,N_16300,N_16420);
and U16715 (N_16715,N_16383,N_16386);
nand U16716 (N_16716,N_16272,N_16367);
and U16717 (N_16717,N_16440,N_16459);
or U16718 (N_16718,N_16348,N_16445);
nand U16719 (N_16719,N_16345,N_16416);
xor U16720 (N_16720,N_16346,N_16258);
nor U16721 (N_16721,N_16324,N_16280);
nor U16722 (N_16722,N_16479,N_16267);
nor U16723 (N_16723,N_16322,N_16328);
nor U16724 (N_16724,N_16437,N_16299);
xor U16725 (N_16725,N_16342,N_16457);
nor U16726 (N_16726,N_16380,N_16364);
nand U16727 (N_16727,N_16394,N_16497);
or U16728 (N_16728,N_16331,N_16368);
nor U16729 (N_16729,N_16472,N_16434);
xnor U16730 (N_16730,N_16439,N_16334);
nor U16731 (N_16731,N_16256,N_16283);
and U16732 (N_16732,N_16311,N_16261);
and U16733 (N_16733,N_16467,N_16452);
xor U16734 (N_16734,N_16336,N_16341);
and U16735 (N_16735,N_16270,N_16333);
nand U16736 (N_16736,N_16274,N_16378);
or U16737 (N_16737,N_16372,N_16370);
nor U16738 (N_16738,N_16307,N_16489);
nand U16739 (N_16739,N_16456,N_16350);
nand U16740 (N_16740,N_16453,N_16266);
and U16741 (N_16741,N_16375,N_16485);
xor U16742 (N_16742,N_16270,N_16338);
or U16743 (N_16743,N_16497,N_16345);
or U16744 (N_16744,N_16358,N_16454);
and U16745 (N_16745,N_16308,N_16437);
or U16746 (N_16746,N_16494,N_16342);
or U16747 (N_16747,N_16428,N_16291);
and U16748 (N_16748,N_16483,N_16445);
or U16749 (N_16749,N_16346,N_16321);
nand U16750 (N_16750,N_16612,N_16745);
and U16751 (N_16751,N_16639,N_16672);
xor U16752 (N_16752,N_16562,N_16656);
nor U16753 (N_16753,N_16552,N_16585);
xor U16754 (N_16754,N_16610,N_16593);
or U16755 (N_16755,N_16618,N_16643);
xor U16756 (N_16756,N_16511,N_16731);
and U16757 (N_16757,N_16685,N_16742);
nor U16758 (N_16758,N_16657,N_16586);
and U16759 (N_16759,N_16500,N_16524);
nand U16760 (N_16760,N_16730,N_16531);
or U16761 (N_16761,N_16702,N_16719);
or U16762 (N_16762,N_16665,N_16622);
nor U16763 (N_16763,N_16613,N_16740);
xor U16764 (N_16764,N_16519,N_16654);
nor U16765 (N_16765,N_16581,N_16725);
nor U16766 (N_16766,N_16735,N_16522);
or U16767 (N_16767,N_16583,N_16544);
nand U16768 (N_16768,N_16734,N_16576);
nand U16769 (N_16769,N_16599,N_16545);
or U16770 (N_16770,N_16688,N_16646);
and U16771 (N_16771,N_16591,N_16503);
and U16772 (N_16772,N_16549,N_16739);
nand U16773 (N_16773,N_16705,N_16594);
xor U16774 (N_16774,N_16523,N_16542);
nor U16775 (N_16775,N_16539,N_16700);
xnor U16776 (N_16776,N_16717,N_16575);
xnor U16777 (N_16777,N_16632,N_16543);
nor U16778 (N_16778,N_16670,N_16709);
xnor U16779 (N_16779,N_16556,N_16693);
or U16780 (N_16780,N_16713,N_16679);
nand U16781 (N_16781,N_16687,N_16720);
and U16782 (N_16782,N_16668,N_16578);
or U16783 (N_16783,N_16572,N_16708);
or U16784 (N_16784,N_16718,N_16736);
and U16785 (N_16785,N_16635,N_16529);
xnor U16786 (N_16786,N_16627,N_16620);
and U16787 (N_16787,N_16553,N_16608);
nand U16788 (N_16788,N_16567,N_16729);
nor U16789 (N_16789,N_16640,N_16642);
and U16790 (N_16790,N_16636,N_16727);
xnor U16791 (N_16791,N_16722,N_16714);
and U16792 (N_16792,N_16653,N_16664);
or U16793 (N_16793,N_16607,N_16507);
xnor U16794 (N_16794,N_16516,N_16631);
or U16795 (N_16795,N_16696,N_16692);
xnor U16796 (N_16796,N_16565,N_16561);
nand U16797 (N_16797,N_16596,N_16538);
nand U16798 (N_16798,N_16704,N_16595);
nor U16799 (N_16799,N_16655,N_16680);
nor U16800 (N_16800,N_16536,N_16728);
nor U16801 (N_16801,N_16744,N_16689);
nor U16802 (N_16802,N_16617,N_16710);
nor U16803 (N_16803,N_16647,N_16590);
nor U16804 (N_16804,N_16526,N_16588);
and U16805 (N_16805,N_16557,N_16533);
nand U16806 (N_16806,N_16724,N_16597);
xnor U16807 (N_16807,N_16648,N_16615);
nor U16808 (N_16808,N_16686,N_16611);
nor U16809 (N_16809,N_16673,N_16695);
or U16810 (N_16810,N_16589,N_16661);
xor U16811 (N_16811,N_16525,N_16569);
or U16812 (N_16812,N_16652,N_16662);
xor U16813 (N_16813,N_16509,N_16645);
nor U16814 (N_16814,N_16603,N_16512);
nor U16815 (N_16815,N_16520,N_16667);
nor U16816 (N_16816,N_16579,N_16532);
nor U16817 (N_16817,N_16733,N_16747);
and U16818 (N_16818,N_16624,N_16634);
nand U16819 (N_16819,N_16501,N_16721);
xnor U16820 (N_16820,N_16546,N_16649);
or U16821 (N_16821,N_16682,N_16726);
nor U16822 (N_16822,N_16605,N_16671);
xnor U16823 (N_16823,N_16570,N_16521);
nand U16824 (N_16824,N_16587,N_16601);
xnor U16825 (N_16825,N_16746,N_16609);
or U16826 (N_16826,N_16690,N_16582);
or U16827 (N_16827,N_16555,N_16681);
nand U16828 (N_16828,N_16505,N_16626);
or U16829 (N_16829,N_16616,N_16691);
nand U16830 (N_16830,N_16559,N_16514);
and U16831 (N_16831,N_16660,N_16659);
nand U16832 (N_16832,N_16614,N_16676);
xor U16833 (N_16833,N_16743,N_16698);
nand U16834 (N_16834,N_16706,N_16748);
xnor U16835 (N_16835,N_16592,N_16551);
nand U16836 (N_16836,N_16602,N_16684);
or U16837 (N_16837,N_16711,N_16629);
nand U16838 (N_16838,N_16644,N_16510);
xor U16839 (N_16839,N_16715,N_16502);
xor U16840 (N_16840,N_16574,N_16716);
nand U16841 (N_16841,N_16699,N_16677);
nand U16842 (N_16842,N_16666,N_16651);
xnor U16843 (N_16843,N_16694,N_16554);
xor U16844 (N_16844,N_16701,N_16628);
or U16845 (N_16845,N_16535,N_16564);
nor U16846 (N_16846,N_16530,N_16606);
or U16847 (N_16847,N_16604,N_16683);
and U16848 (N_16848,N_16633,N_16738);
nand U16849 (N_16849,N_16678,N_16504);
or U16850 (N_16850,N_16737,N_16550);
nor U16851 (N_16851,N_16560,N_16749);
or U16852 (N_16852,N_16537,N_16518);
and U16853 (N_16853,N_16638,N_16517);
xnor U16854 (N_16854,N_16513,N_16515);
nand U16855 (N_16855,N_16568,N_16558);
xnor U16856 (N_16856,N_16674,N_16508);
xnor U16857 (N_16857,N_16663,N_16703);
and U16858 (N_16858,N_16625,N_16548);
or U16859 (N_16859,N_16600,N_16584);
nand U16860 (N_16860,N_16641,N_16707);
xnor U16861 (N_16861,N_16741,N_16527);
nor U16862 (N_16862,N_16723,N_16675);
and U16863 (N_16863,N_16712,N_16580);
and U16864 (N_16864,N_16650,N_16563);
xnor U16865 (N_16865,N_16577,N_16571);
nand U16866 (N_16866,N_16540,N_16732);
and U16867 (N_16867,N_16534,N_16573);
nor U16868 (N_16868,N_16619,N_16637);
and U16869 (N_16869,N_16598,N_16566);
nand U16870 (N_16870,N_16697,N_16541);
xor U16871 (N_16871,N_16630,N_16623);
or U16872 (N_16872,N_16658,N_16506);
nand U16873 (N_16873,N_16528,N_16669);
nand U16874 (N_16874,N_16547,N_16621);
nor U16875 (N_16875,N_16543,N_16740);
and U16876 (N_16876,N_16501,N_16683);
and U16877 (N_16877,N_16562,N_16518);
and U16878 (N_16878,N_16742,N_16600);
or U16879 (N_16879,N_16610,N_16631);
nor U16880 (N_16880,N_16575,N_16518);
or U16881 (N_16881,N_16501,N_16714);
xnor U16882 (N_16882,N_16745,N_16697);
nor U16883 (N_16883,N_16528,N_16536);
xnor U16884 (N_16884,N_16655,N_16717);
nor U16885 (N_16885,N_16683,N_16694);
nor U16886 (N_16886,N_16543,N_16656);
nand U16887 (N_16887,N_16615,N_16638);
or U16888 (N_16888,N_16624,N_16708);
nand U16889 (N_16889,N_16675,N_16510);
xnor U16890 (N_16890,N_16625,N_16710);
xnor U16891 (N_16891,N_16545,N_16584);
and U16892 (N_16892,N_16587,N_16641);
xor U16893 (N_16893,N_16547,N_16542);
xor U16894 (N_16894,N_16611,N_16644);
nand U16895 (N_16895,N_16573,N_16668);
or U16896 (N_16896,N_16704,N_16706);
nor U16897 (N_16897,N_16561,N_16705);
xor U16898 (N_16898,N_16724,N_16573);
xnor U16899 (N_16899,N_16592,N_16552);
nand U16900 (N_16900,N_16585,N_16520);
xor U16901 (N_16901,N_16645,N_16585);
nand U16902 (N_16902,N_16500,N_16508);
nand U16903 (N_16903,N_16671,N_16680);
xnor U16904 (N_16904,N_16508,N_16746);
and U16905 (N_16905,N_16598,N_16505);
xnor U16906 (N_16906,N_16720,N_16718);
or U16907 (N_16907,N_16700,N_16576);
nand U16908 (N_16908,N_16599,N_16610);
nor U16909 (N_16909,N_16729,N_16704);
nand U16910 (N_16910,N_16556,N_16537);
and U16911 (N_16911,N_16727,N_16675);
and U16912 (N_16912,N_16648,N_16744);
xor U16913 (N_16913,N_16727,N_16538);
nor U16914 (N_16914,N_16726,N_16582);
xor U16915 (N_16915,N_16677,N_16718);
xnor U16916 (N_16916,N_16578,N_16534);
nor U16917 (N_16917,N_16512,N_16688);
or U16918 (N_16918,N_16587,N_16504);
or U16919 (N_16919,N_16555,N_16522);
and U16920 (N_16920,N_16680,N_16561);
xor U16921 (N_16921,N_16700,N_16671);
xor U16922 (N_16922,N_16629,N_16637);
xnor U16923 (N_16923,N_16537,N_16566);
xor U16924 (N_16924,N_16697,N_16525);
nor U16925 (N_16925,N_16595,N_16529);
or U16926 (N_16926,N_16560,N_16721);
xnor U16927 (N_16927,N_16633,N_16515);
xnor U16928 (N_16928,N_16685,N_16582);
nor U16929 (N_16929,N_16604,N_16748);
nor U16930 (N_16930,N_16685,N_16502);
xnor U16931 (N_16931,N_16538,N_16740);
and U16932 (N_16932,N_16557,N_16630);
and U16933 (N_16933,N_16717,N_16597);
and U16934 (N_16934,N_16749,N_16691);
nand U16935 (N_16935,N_16557,N_16749);
or U16936 (N_16936,N_16590,N_16681);
and U16937 (N_16937,N_16612,N_16600);
or U16938 (N_16938,N_16685,N_16536);
xnor U16939 (N_16939,N_16617,N_16588);
and U16940 (N_16940,N_16672,N_16744);
and U16941 (N_16941,N_16609,N_16600);
nand U16942 (N_16942,N_16718,N_16661);
xor U16943 (N_16943,N_16533,N_16596);
and U16944 (N_16944,N_16560,N_16530);
nand U16945 (N_16945,N_16689,N_16569);
or U16946 (N_16946,N_16593,N_16528);
xnor U16947 (N_16947,N_16605,N_16530);
and U16948 (N_16948,N_16719,N_16706);
nor U16949 (N_16949,N_16631,N_16685);
nor U16950 (N_16950,N_16549,N_16662);
or U16951 (N_16951,N_16681,N_16578);
or U16952 (N_16952,N_16535,N_16666);
nand U16953 (N_16953,N_16556,N_16744);
and U16954 (N_16954,N_16638,N_16607);
nand U16955 (N_16955,N_16637,N_16504);
and U16956 (N_16956,N_16578,N_16715);
xnor U16957 (N_16957,N_16651,N_16734);
nand U16958 (N_16958,N_16598,N_16535);
or U16959 (N_16959,N_16556,N_16722);
or U16960 (N_16960,N_16526,N_16627);
nand U16961 (N_16961,N_16632,N_16601);
nand U16962 (N_16962,N_16606,N_16660);
or U16963 (N_16963,N_16584,N_16593);
xnor U16964 (N_16964,N_16612,N_16500);
nand U16965 (N_16965,N_16507,N_16744);
xor U16966 (N_16966,N_16686,N_16540);
xnor U16967 (N_16967,N_16662,N_16605);
and U16968 (N_16968,N_16545,N_16655);
xor U16969 (N_16969,N_16571,N_16527);
or U16970 (N_16970,N_16695,N_16535);
nand U16971 (N_16971,N_16630,N_16508);
nand U16972 (N_16972,N_16728,N_16722);
xor U16973 (N_16973,N_16632,N_16619);
xnor U16974 (N_16974,N_16651,N_16619);
nor U16975 (N_16975,N_16746,N_16643);
nor U16976 (N_16976,N_16691,N_16609);
or U16977 (N_16977,N_16539,N_16748);
and U16978 (N_16978,N_16544,N_16638);
xor U16979 (N_16979,N_16668,N_16550);
or U16980 (N_16980,N_16667,N_16735);
nand U16981 (N_16981,N_16707,N_16689);
nor U16982 (N_16982,N_16679,N_16624);
xor U16983 (N_16983,N_16528,N_16503);
nor U16984 (N_16984,N_16694,N_16592);
nor U16985 (N_16985,N_16573,N_16749);
xor U16986 (N_16986,N_16532,N_16746);
or U16987 (N_16987,N_16644,N_16544);
xnor U16988 (N_16988,N_16616,N_16645);
xnor U16989 (N_16989,N_16719,N_16591);
xor U16990 (N_16990,N_16663,N_16742);
nand U16991 (N_16991,N_16627,N_16514);
nor U16992 (N_16992,N_16589,N_16638);
nor U16993 (N_16993,N_16683,N_16638);
and U16994 (N_16994,N_16708,N_16693);
nand U16995 (N_16995,N_16715,N_16535);
and U16996 (N_16996,N_16713,N_16667);
nand U16997 (N_16997,N_16518,N_16742);
nor U16998 (N_16998,N_16578,N_16508);
nand U16999 (N_16999,N_16663,N_16620);
nand U17000 (N_17000,N_16789,N_16886);
and U17001 (N_17001,N_16906,N_16910);
or U17002 (N_17002,N_16971,N_16979);
nand U17003 (N_17003,N_16922,N_16811);
and U17004 (N_17004,N_16919,N_16771);
or U17005 (N_17005,N_16907,N_16933);
xnor U17006 (N_17006,N_16778,N_16889);
nand U17007 (N_17007,N_16888,N_16961);
nand U17008 (N_17008,N_16801,N_16960);
nand U17009 (N_17009,N_16800,N_16904);
xnor U17010 (N_17010,N_16772,N_16903);
and U17011 (N_17011,N_16905,N_16926);
nor U17012 (N_17012,N_16970,N_16785);
xnor U17013 (N_17013,N_16947,N_16767);
nand U17014 (N_17014,N_16783,N_16917);
nand U17015 (N_17015,N_16898,N_16948);
or U17016 (N_17016,N_16795,N_16807);
and U17017 (N_17017,N_16844,N_16791);
nand U17018 (N_17018,N_16859,N_16794);
and U17019 (N_17019,N_16850,N_16851);
and U17020 (N_17020,N_16820,N_16892);
and U17021 (N_17021,N_16992,N_16923);
nor U17022 (N_17022,N_16842,N_16941);
or U17023 (N_17023,N_16880,N_16757);
nand U17024 (N_17024,N_16829,N_16884);
nand U17025 (N_17025,N_16848,N_16990);
nor U17026 (N_17026,N_16956,N_16949);
nand U17027 (N_17027,N_16838,N_16980);
and U17028 (N_17028,N_16847,N_16999);
xnor U17029 (N_17029,N_16901,N_16938);
nor U17030 (N_17030,N_16989,N_16890);
and U17031 (N_17031,N_16865,N_16802);
and U17032 (N_17032,N_16927,N_16997);
xor U17033 (N_17033,N_16774,N_16872);
nor U17034 (N_17034,N_16831,N_16840);
nand U17035 (N_17035,N_16944,N_16914);
and U17036 (N_17036,N_16895,N_16885);
or U17037 (N_17037,N_16845,N_16766);
nor U17038 (N_17038,N_16788,N_16962);
nand U17039 (N_17039,N_16937,N_16893);
xnor U17040 (N_17040,N_16856,N_16822);
or U17041 (N_17041,N_16902,N_16758);
and U17042 (N_17042,N_16854,N_16752);
and U17043 (N_17043,N_16994,N_16875);
or U17044 (N_17044,N_16899,N_16770);
and U17045 (N_17045,N_16755,N_16779);
nand U17046 (N_17046,N_16759,N_16821);
or U17047 (N_17047,N_16977,N_16803);
xnor U17048 (N_17048,N_16972,N_16943);
nand U17049 (N_17049,N_16853,N_16958);
or U17050 (N_17050,N_16866,N_16861);
and U17051 (N_17051,N_16756,N_16876);
nand U17052 (N_17052,N_16965,N_16868);
and U17053 (N_17053,N_16974,N_16978);
or U17054 (N_17054,N_16964,N_16998);
xor U17055 (N_17055,N_16753,N_16867);
or U17056 (N_17056,N_16928,N_16858);
nor U17057 (N_17057,N_16834,N_16967);
xnor U17058 (N_17058,N_16931,N_16874);
and U17059 (N_17059,N_16963,N_16839);
nand U17060 (N_17060,N_16894,N_16953);
and U17061 (N_17061,N_16780,N_16827);
nand U17062 (N_17062,N_16793,N_16835);
nand U17063 (N_17063,N_16814,N_16932);
nand U17064 (N_17064,N_16760,N_16878);
and U17065 (N_17065,N_16900,N_16776);
nor U17066 (N_17066,N_16934,N_16983);
xnor U17067 (N_17067,N_16855,N_16987);
or U17068 (N_17068,N_16764,N_16986);
nand U17069 (N_17069,N_16768,N_16891);
nand U17070 (N_17070,N_16818,N_16881);
nor U17071 (N_17071,N_16913,N_16995);
nor U17072 (N_17072,N_16750,N_16826);
nand U17073 (N_17073,N_16836,N_16897);
nand U17074 (N_17074,N_16832,N_16942);
nand U17075 (N_17075,N_16925,N_16911);
nor U17076 (N_17076,N_16815,N_16804);
xor U17077 (N_17077,N_16812,N_16796);
and U17078 (N_17078,N_16976,N_16823);
and U17079 (N_17079,N_16882,N_16981);
nand U17080 (N_17080,N_16765,N_16763);
nand U17081 (N_17081,N_16828,N_16860);
nand U17082 (N_17082,N_16887,N_16952);
nor U17083 (N_17083,N_16985,N_16769);
or U17084 (N_17084,N_16864,N_16936);
xor U17085 (N_17085,N_16806,N_16798);
and U17086 (N_17086,N_16915,N_16805);
nor U17087 (N_17087,N_16813,N_16852);
nand U17088 (N_17088,N_16773,N_16883);
nor U17089 (N_17089,N_16939,N_16973);
or U17090 (N_17090,N_16761,N_16825);
nor U17091 (N_17091,N_16879,N_16968);
and U17092 (N_17092,N_16975,N_16799);
xnor U17093 (N_17093,N_16817,N_16869);
nor U17094 (N_17094,N_16996,N_16993);
nand U17095 (N_17095,N_16966,N_16809);
nand U17096 (N_17096,N_16930,N_16863);
nor U17097 (N_17097,N_16870,N_16957);
nor U17098 (N_17098,N_16808,N_16918);
nor U17099 (N_17099,N_16754,N_16843);
and U17100 (N_17100,N_16777,N_16871);
nor U17101 (N_17101,N_16959,N_16792);
or U17102 (N_17102,N_16896,N_16955);
xor U17103 (N_17103,N_16797,N_16940);
xor U17104 (N_17104,N_16921,N_16916);
and U17105 (N_17105,N_16849,N_16857);
xor U17106 (N_17106,N_16837,N_16991);
or U17107 (N_17107,N_16846,N_16830);
nor U17108 (N_17108,N_16950,N_16984);
nand U17109 (N_17109,N_16969,N_16841);
xnor U17110 (N_17110,N_16946,N_16912);
or U17111 (N_17111,N_16945,N_16824);
nand U17112 (N_17112,N_16819,N_16762);
xnor U17113 (N_17113,N_16784,N_16951);
and U17114 (N_17114,N_16935,N_16924);
xnor U17115 (N_17115,N_16781,N_16862);
nand U17116 (N_17116,N_16787,N_16877);
xnor U17117 (N_17117,N_16982,N_16751);
nand U17118 (N_17118,N_16929,N_16873);
xnor U17119 (N_17119,N_16908,N_16816);
nand U17120 (N_17120,N_16786,N_16810);
nor U17121 (N_17121,N_16920,N_16790);
xnor U17122 (N_17122,N_16833,N_16775);
and U17123 (N_17123,N_16988,N_16909);
xor U17124 (N_17124,N_16782,N_16954);
or U17125 (N_17125,N_16899,N_16751);
or U17126 (N_17126,N_16983,N_16819);
and U17127 (N_17127,N_16984,N_16780);
and U17128 (N_17128,N_16895,N_16933);
nor U17129 (N_17129,N_16932,N_16788);
nand U17130 (N_17130,N_16841,N_16992);
nor U17131 (N_17131,N_16845,N_16850);
or U17132 (N_17132,N_16753,N_16896);
nand U17133 (N_17133,N_16964,N_16790);
nand U17134 (N_17134,N_16947,N_16883);
and U17135 (N_17135,N_16782,N_16880);
nor U17136 (N_17136,N_16905,N_16919);
nand U17137 (N_17137,N_16851,N_16931);
or U17138 (N_17138,N_16865,N_16788);
xnor U17139 (N_17139,N_16842,N_16916);
nand U17140 (N_17140,N_16903,N_16819);
xor U17141 (N_17141,N_16927,N_16773);
and U17142 (N_17142,N_16824,N_16993);
nand U17143 (N_17143,N_16837,N_16792);
and U17144 (N_17144,N_16898,N_16907);
or U17145 (N_17145,N_16873,N_16893);
nor U17146 (N_17146,N_16756,N_16965);
nand U17147 (N_17147,N_16797,N_16962);
or U17148 (N_17148,N_16946,N_16977);
or U17149 (N_17149,N_16922,N_16996);
nor U17150 (N_17150,N_16771,N_16992);
and U17151 (N_17151,N_16839,N_16928);
or U17152 (N_17152,N_16803,N_16972);
and U17153 (N_17153,N_16850,N_16800);
nand U17154 (N_17154,N_16906,N_16839);
and U17155 (N_17155,N_16750,N_16829);
xnor U17156 (N_17156,N_16944,N_16957);
xnor U17157 (N_17157,N_16959,N_16881);
nand U17158 (N_17158,N_16869,N_16931);
xor U17159 (N_17159,N_16750,N_16929);
nor U17160 (N_17160,N_16989,N_16764);
nor U17161 (N_17161,N_16845,N_16752);
nor U17162 (N_17162,N_16808,N_16997);
nand U17163 (N_17163,N_16787,N_16818);
xor U17164 (N_17164,N_16970,N_16969);
and U17165 (N_17165,N_16936,N_16859);
nor U17166 (N_17166,N_16944,N_16777);
nand U17167 (N_17167,N_16990,N_16817);
xor U17168 (N_17168,N_16997,N_16904);
xnor U17169 (N_17169,N_16810,N_16966);
and U17170 (N_17170,N_16775,N_16983);
xnor U17171 (N_17171,N_16766,N_16869);
nand U17172 (N_17172,N_16754,N_16859);
and U17173 (N_17173,N_16954,N_16929);
nor U17174 (N_17174,N_16792,N_16798);
or U17175 (N_17175,N_16986,N_16901);
nand U17176 (N_17176,N_16850,N_16823);
nor U17177 (N_17177,N_16931,N_16754);
xnor U17178 (N_17178,N_16979,N_16859);
xor U17179 (N_17179,N_16874,N_16925);
and U17180 (N_17180,N_16961,N_16882);
and U17181 (N_17181,N_16754,N_16862);
and U17182 (N_17182,N_16820,N_16815);
nor U17183 (N_17183,N_16770,N_16811);
nor U17184 (N_17184,N_16937,N_16923);
and U17185 (N_17185,N_16989,N_16765);
xnor U17186 (N_17186,N_16806,N_16871);
xor U17187 (N_17187,N_16815,N_16914);
xor U17188 (N_17188,N_16790,N_16915);
and U17189 (N_17189,N_16976,N_16951);
nor U17190 (N_17190,N_16839,N_16834);
and U17191 (N_17191,N_16850,N_16764);
or U17192 (N_17192,N_16999,N_16756);
or U17193 (N_17193,N_16900,N_16819);
xnor U17194 (N_17194,N_16839,N_16998);
xnor U17195 (N_17195,N_16791,N_16898);
and U17196 (N_17196,N_16803,N_16833);
nand U17197 (N_17197,N_16889,N_16867);
nand U17198 (N_17198,N_16944,N_16784);
xor U17199 (N_17199,N_16929,N_16968);
xnor U17200 (N_17200,N_16887,N_16918);
or U17201 (N_17201,N_16843,N_16839);
or U17202 (N_17202,N_16872,N_16911);
and U17203 (N_17203,N_16840,N_16841);
xor U17204 (N_17204,N_16987,N_16875);
nor U17205 (N_17205,N_16868,N_16799);
and U17206 (N_17206,N_16785,N_16798);
or U17207 (N_17207,N_16831,N_16957);
xnor U17208 (N_17208,N_16908,N_16807);
nand U17209 (N_17209,N_16920,N_16781);
nand U17210 (N_17210,N_16955,N_16986);
and U17211 (N_17211,N_16938,N_16935);
and U17212 (N_17212,N_16797,N_16941);
or U17213 (N_17213,N_16811,N_16768);
nand U17214 (N_17214,N_16822,N_16815);
nand U17215 (N_17215,N_16941,N_16944);
nor U17216 (N_17216,N_16760,N_16857);
and U17217 (N_17217,N_16978,N_16991);
nor U17218 (N_17218,N_16944,N_16816);
and U17219 (N_17219,N_16992,N_16849);
and U17220 (N_17220,N_16855,N_16998);
and U17221 (N_17221,N_16804,N_16844);
nor U17222 (N_17222,N_16889,N_16927);
xnor U17223 (N_17223,N_16829,N_16986);
and U17224 (N_17224,N_16994,N_16878);
and U17225 (N_17225,N_16931,N_16856);
xor U17226 (N_17226,N_16858,N_16871);
and U17227 (N_17227,N_16967,N_16774);
or U17228 (N_17228,N_16920,N_16937);
and U17229 (N_17229,N_16815,N_16842);
xnor U17230 (N_17230,N_16994,N_16800);
nor U17231 (N_17231,N_16845,N_16966);
nor U17232 (N_17232,N_16823,N_16939);
and U17233 (N_17233,N_16970,N_16870);
or U17234 (N_17234,N_16991,N_16823);
and U17235 (N_17235,N_16815,N_16785);
and U17236 (N_17236,N_16839,N_16970);
nor U17237 (N_17237,N_16897,N_16884);
or U17238 (N_17238,N_16911,N_16755);
and U17239 (N_17239,N_16906,N_16810);
nor U17240 (N_17240,N_16951,N_16806);
xor U17241 (N_17241,N_16997,N_16790);
xor U17242 (N_17242,N_16896,N_16887);
xor U17243 (N_17243,N_16759,N_16791);
and U17244 (N_17244,N_16812,N_16828);
xor U17245 (N_17245,N_16759,N_16822);
nor U17246 (N_17246,N_16975,N_16915);
nor U17247 (N_17247,N_16968,N_16851);
nand U17248 (N_17248,N_16758,N_16795);
or U17249 (N_17249,N_16766,N_16837);
or U17250 (N_17250,N_17112,N_17150);
nor U17251 (N_17251,N_17045,N_17046);
nand U17252 (N_17252,N_17179,N_17003);
nor U17253 (N_17253,N_17210,N_17165);
and U17254 (N_17254,N_17117,N_17017);
and U17255 (N_17255,N_17102,N_17122);
and U17256 (N_17256,N_17141,N_17224);
and U17257 (N_17257,N_17114,N_17175);
nor U17258 (N_17258,N_17158,N_17075);
and U17259 (N_17259,N_17015,N_17187);
xnor U17260 (N_17260,N_17007,N_17245);
xor U17261 (N_17261,N_17155,N_17092);
and U17262 (N_17262,N_17199,N_17218);
and U17263 (N_17263,N_17002,N_17244);
nor U17264 (N_17264,N_17048,N_17162);
nand U17265 (N_17265,N_17032,N_17108);
or U17266 (N_17266,N_17131,N_17088);
xnor U17267 (N_17267,N_17174,N_17226);
and U17268 (N_17268,N_17231,N_17191);
nand U17269 (N_17269,N_17043,N_17080);
and U17270 (N_17270,N_17180,N_17097);
xnor U17271 (N_17271,N_17010,N_17103);
or U17272 (N_17272,N_17056,N_17094);
nand U17273 (N_17273,N_17203,N_17125);
nor U17274 (N_17274,N_17026,N_17240);
xnor U17275 (N_17275,N_17055,N_17035);
nor U17276 (N_17276,N_17189,N_17115);
or U17277 (N_17277,N_17087,N_17182);
or U17278 (N_17278,N_17148,N_17246);
xnor U17279 (N_17279,N_17132,N_17042);
and U17280 (N_17280,N_17221,N_17028);
xor U17281 (N_17281,N_17215,N_17078);
or U17282 (N_17282,N_17000,N_17160);
nand U17283 (N_17283,N_17036,N_17128);
nor U17284 (N_17284,N_17070,N_17027);
or U17285 (N_17285,N_17213,N_17126);
xnor U17286 (N_17286,N_17152,N_17037);
nor U17287 (N_17287,N_17209,N_17201);
or U17288 (N_17288,N_17023,N_17001);
and U17289 (N_17289,N_17192,N_17107);
nor U17290 (N_17290,N_17237,N_17163);
or U17291 (N_17291,N_17133,N_17190);
xor U17292 (N_17292,N_17166,N_17071);
nor U17293 (N_17293,N_17137,N_17138);
xnor U17294 (N_17294,N_17156,N_17013);
and U17295 (N_17295,N_17247,N_17105);
xor U17296 (N_17296,N_17196,N_17177);
xnor U17297 (N_17297,N_17066,N_17211);
nor U17298 (N_17298,N_17044,N_17123);
nand U17299 (N_17299,N_17020,N_17142);
nor U17300 (N_17300,N_17079,N_17051);
xor U17301 (N_17301,N_17049,N_17034);
xor U17302 (N_17302,N_17081,N_17083);
or U17303 (N_17303,N_17157,N_17151);
xor U17304 (N_17304,N_17176,N_17171);
and U17305 (N_17305,N_17022,N_17031);
xor U17306 (N_17306,N_17161,N_17019);
or U17307 (N_17307,N_17145,N_17091);
or U17308 (N_17308,N_17005,N_17186);
and U17309 (N_17309,N_17129,N_17219);
xnor U17310 (N_17310,N_17134,N_17012);
nor U17311 (N_17311,N_17217,N_17225);
and U17312 (N_17312,N_17068,N_17135);
nand U17313 (N_17313,N_17111,N_17099);
or U17314 (N_17314,N_17062,N_17220);
xor U17315 (N_17315,N_17139,N_17104);
or U17316 (N_17316,N_17030,N_17033);
nor U17317 (N_17317,N_17052,N_17098);
and U17318 (N_17318,N_17127,N_17064);
xor U17319 (N_17319,N_17222,N_17106);
xnor U17320 (N_17320,N_17038,N_17058);
nor U17321 (N_17321,N_17119,N_17159);
and U17322 (N_17322,N_17193,N_17061);
nor U17323 (N_17323,N_17147,N_17248);
xnor U17324 (N_17324,N_17086,N_17149);
and U17325 (N_17325,N_17229,N_17095);
xnor U17326 (N_17326,N_17050,N_17183);
or U17327 (N_17327,N_17205,N_17168);
and U17328 (N_17328,N_17060,N_17207);
xor U17329 (N_17329,N_17188,N_17076);
or U17330 (N_17330,N_17195,N_17054);
and U17331 (N_17331,N_17082,N_17173);
xnor U17332 (N_17332,N_17185,N_17004);
and U17333 (N_17333,N_17072,N_17096);
xor U17334 (N_17334,N_17069,N_17235);
nor U17335 (N_17335,N_17109,N_17110);
and U17336 (N_17336,N_17241,N_17118);
and U17337 (N_17337,N_17090,N_17204);
and U17338 (N_17338,N_17197,N_17085);
nand U17339 (N_17339,N_17249,N_17074);
nand U17340 (N_17340,N_17011,N_17073);
and U17341 (N_17341,N_17198,N_17208);
xor U17342 (N_17342,N_17233,N_17093);
nand U17343 (N_17343,N_17113,N_17143);
or U17344 (N_17344,N_17154,N_17077);
or U17345 (N_17345,N_17018,N_17232);
nand U17346 (N_17346,N_17169,N_17057);
and U17347 (N_17347,N_17202,N_17178);
xnor U17348 (N_17348,N_17025,N_17167);
nand U17349 (N_17349,N_17243,N_17041);
nand U17350 (N_17350,N_17214,N_17172);
and U17351 (N_17351,N_17040,N_17029);
xnor U17352 (N_17352,N_17016,N_17238);
and U17353 (N_17353,N_17120,N_17227);
nor U17354 (N_17354,N_17206,N_17124);
xnor U17355 (N_17355,N_17053,N_17130);
nor U17356 (N_17356,N_17089,N_17212);
xor U17357 (N_17357,N_17216,N_17140);
nand U17358 (N_17358,N_17116,N_17047);
xnor U17359 (N_17359,N_17194,N_17234);
or U17360 (N_17360,N_17239,N_17236);
nor U17361 (N_17361,N_17200,N_17223);
and U17362 (N_17362,N_17121,N_17006);
nor U17363 (N_17363,N_17101,N_17067);
nor U17364 (N_17364,N_17039,N_17065);
or U17365 (N_17365,N_17228,N_17100);
and U17366 (N_17366,N_17153,N_17084);
or U17367 (N_17367,N_17009,N_17136);
or U17368 (N_17368,N_17230,N_17059);
xnor U17369 (N_17369,N_17164,N_17008);
xor U17370 (N_17370,N_17184,N_17063);
and U17371 (N_17371,N_17014,N_17144);
xor U17372 (N_17372,N_17021,N_17170);
nand U17373 (N_17373,N_17146,N_17024);
nand U17374 (N_17374,N_17181,N_17242);
and U17375 (N_17375,N_17190,N_17084);
nor U17376 (N_17376,N_17013,N_17057);
and U17377 (N_17377,N_17042,N_17241);
or U17378 (N_17378,N_17074,N_17178);
or U17379 (N_17379,N_17190,N_17157);
nor U17380 (N_17380,N_17008,N_17127);
nand U17381 (N_17381,N_17147,N_17172);
xnor U17382 (N_17382,N_17196,N_17090);
nor U17383 (N_17383,N_17036,N_17091);
or U17384 (N_17384,N_17042,N_17146);
nor U17385 (N_17385,N_17136,N_17010);
xnor U17386 (N_17386,N_17010,N_17053);
nand U17387 (N_17387,N_17150,N_17020);
nor U17388 (N_17388,N_17022,N_17060);
or U17389 (N_17389,N_17161,N_17220);
nand U17390 (N_17390,N_17055,N_17207);
nand U17391 (N_17391,N_17207,N_17219);
or U17392 (N_17392,N_17054,N_17044);
xor U17393 (N_17393,N_17138,N_17100);
or U17394 (N_17394,N_17079,N_17173);
nand U17395 (N_17395,N_17092,N_17179);
or U17396 (N_17396,N_17147,N_17083);
xor U17397 (N_17397,N_17099,N_17057);
and U17398 (N_17398,N_17200,N_17045);
and U17399 (N_17399,N_17053,N_17001);
xnor U17400 (N_17400,N_17190,N_17090);
and U17401 (N_17401,N_17164,N_17049);
and U17402 (N_17402,N_17169,N_17154);
nand U17403 (N_17403,N_17006,N_17179);
nand U17404 (N_17404,N_17116,N_17152);
nor U17405 (N_17405,N_17106,N_17162);
or U17406 (N_17406,N_17057,N_17149);
and U17407 (N_17407,N_17233,N_17043);
or U17408 (N_17408,N_17104,N_17214);
nand U17409 (N_17409,N_17141,N_17046);
and U17410 (N_17410,N_17130,N_17218);
or U17411 (N_17411,N_17050,N_17228);
nor U17412 (N_17412,N_17203,N_17159);
xnor U17413 (N_17413,N_17066,N_17117);
nand U17414 (N_17414,N_17156,N_17199);
or U17415 (N_17415,N_17036,N_17238);
or U17416 (N_17416,N_17162,N_17104);
xnor U17417 (N_17417,N_17119,N_17091);
or U17418 (N_17418,N_17068,N_17076);
nand U17419 (N_17419,N_17011,N_17111);
and U17420 (N_17420,N_17200,N_17084);
and U17421 (N_17421,N_17228,N_17197);
xnor U17422 (N_17422,N_17146,N_17099);
and U17423 (N_17423,N_17128,N_17054);
and U17424 (N_17424,N_17176,N_17059);
xor U17425 (N_17425,N_17071,N_17218);
nand U17426 (N_17426,N_17021,N_17000);
or U17427 (N_17427,N_17019,N_17169);
or U17428 (N_17428,N_17132,N_17195);
nand U17429 (N_17429,N_17068,N_17040);
nor U17430 (N_17430,N_17091,N_17126);
nor U17431 (N_17431,N_17225,N_17238);
or U17432 (N_17432,N_17166,N_17164);
and U17433 (N_17433,N_17175,N_17073);
nor U17434 (N_17434,N_17019,N_17136);
xnor U17435 (N_17435,N_17085,N_17067);
or U17436 (N_17436,N_17075,N_17157);
nand U17437 (N_17437,N_17245,N_17104);
xnor U17438 (N_17438,N_17099,N_17033);
or U17439 (N_17439,N_17130,N_17232);
and U17440 (N_17440,N_17198,N_17169);
xor U17441 (N_17441,N_17039,N_17004);
nor U17442 (N_17442,N_17067,N_17009);
nand U17443 (N_17443,N_17199,N_17109);
nand U17444 (N_17444,N_17097,N_17220);
and U17445 (N_17445,N_17248,N_17090);
or U17446 (N_17446,N_17058,N_17103);
xnor U17447 (N_17447,N_17139,N_17196);
nor U17448 (N_17448,N_17133,N_17154);
or U17449 (N_17449,N_17151,N_17093);
nand U17450 (N_17450,N_17217,N_17134);
nand U17451 (N_17451,N_17153,N_17189);
nand U17452 (N_17452,N_17051,N_17083);
or U17453 (N_17453,N_17061,N_17046);
xor U17454 (N_17454,N_17031,N_17169);
nor U17455 (N_17455,N_17057,N_17014);
nand U17456 (N_17456,N_17050,N_17164);
nand U17457 (N_17457,N_17177,N_17195);
nor U17458 (N_17458,N_17164,N_17153);
xor U17459 (N_17459,N_17015,N_17122);
xor U17460 (N_17460,N_17018,N_17145);
xnor U17461 (N_17461,N_17176,N_17184);
nand U17462 (N_17462,N_17038,N_17092);
nand U17463 (N_17463,N_17127,N_17104);
nor U17464 (N_17464,N_17147,N_17000);
nor U17465 (N_17465,N_17126,N_17216);
nor U17466 (N_17466,N_17196,N_17147);
and U17467 (N_17467,N_17220,N_17088);
nor U17468 (N_17468,N_17017,N_17094);
xnor U17469 (N_17469,N_17213,N_17159);
or U17470 (N_17470,N_17000,N_17237);
nand U17471 (N_17471,N_17133,N_17060);
or U17472 (N_17472,N_17103,N_17171);
xor U17473 (N_17473,N_17014,N_17145);
nor U17474 (N_17474,N_17232,N_17111);
nor U17475 (N_17475,N_17121,N_17044);
and U17476 (N_17476,N_17139,N_17040);
and U17477 (N_17477,N_17008,N_17204);
or U17478 (N_17478,N_17131,N_17056);
nand U17479 (N_17479,N_17216,N_17040);
nand U17480 (N_17480,N_17114,N_17089);
and U17481 (N_17481,N_17061,N_17197);
xnor U17482 (N_17482,N_17243,N_17009);
or U17483 (N_17483,N_17167,N_17234);
nor U17484 (N_17484,N_17227,N_17176);
and U17485 (N_17485,N_17208,N_17179);
xnor U17486 (N_17486,N_17050,N_17129);
xor U17487 (N_17487,N_17032,N_17147);
nor U17488 (N_17488,N_17211,N_17204);
xor U17489 (N_17489,N_17103,N_17167);
or U17490 (N_17490,N_17196,N_17048);
nand U17491 (N_17491,N_17168,N_17047);
and U17492 (N_17492,N_17159,N_17177);
nand U17493 (N_17493,N_17116,N_17139);
xnor U17494 (N_17494,N_17174,N_17239);
nand U17495 (N_17495,N_17249,N_17232);
or U17496 (N_17496,N_17192,N_17134);
nor U17497 (N_17497,N_17083,N_17142);
nor U17498 (N_17498,N_17208,N_17151);
or U17499 (N_17499,N_17085,N_17199);
or U17500 (N_17500,N_17344,N_17447);
xnor U17501 (N_17501,N_17375,N_17358);
xnor U17502 (N_17502,N_17263,N_17299);
nand U17503 (N_17503,N_17318,N_17330);
nor U17504 (N_17504,N_17311,N_17279);
nand U17505 (N_17505,N_17421,N_17469);
xnor U17506 (N_17506,N_17293,N_17496);
or U17507 (N_17507,N_17402,N_17345);
nand U17508 (N_17508,N_17270,N_17314);
xnor U17509 (N_17509,N_17442,N_17264);
and U17510 (N_17510,N_17266,N_17336);
or U17511 (N_17511,N_17269,N_17477);
nor U17512 (N_17512,N_17411,N_17438);
and U17513 (N_17513,N_17484,N_17453);
or U17514 (N_17514,N_17407,N_17403);
and U17515 (N_17515,N_17487,N_17347);
xnor U17516 (N_17516,N_17492,N_17388);
nor U17517 (N_17517,N_17291,N_17325);
nor U17518 (N_17518,N_17408,N_17425);
nand U17519 (N_17519,N_17301,N_17446);
or U17520 (N_17520,N_17437,N_17465);
and U17521 (N_17521,N_17267,N_17409);
nand U17522 (N_17522,N_17371,N_17294);
or U17523 (N_17523,N_17395,N_17404);
nand U17524 (N_17524,N_17374,N_17315);
or U17525 (N_17525,N_17420,N_17332);
nand U17526 (N_17526,N_17415,N_17365);
or U17527 (N_17527,N_17430,N_17457);
or U17528 (N_17528,N_17253,N_17423);
xor U17529 (N_17529,N_17275,N_17381);
and U17530 (N_17530,N_17312,N_17260);
nor U17531 (N_17531,N_17452,N_17460);
nor U17532 (N_17532,N_17431,N_17262);
and U17533 (N_17533,N_17254,N_17339);
xnor U17534 (N_17534,N_17351,N_17333);
xnor U17535 (N_17535,N_17359,N_17323);
or U17536 (N_17536,N_17448,N_17288);
xnor U17537 (N_17537,N_17272,N_17441);
or U17538 (N_17538,N_17474,N_17440);
nand U17539 (N_17539,N_17406,N_17385);
or U17540 (N_17540,N_17317,N_17372);
and U17541 (N_17541,N_17483,N_17256);
and U17542 (N_17542,N_17303,N_17429);
or U17543 (N_17543,N_17286,N_17445);
nor U17544 (N_17544,N_17384,N_17470);
xor U17545 (N_17545,N_17498,N_17418);
nand U17546 (N_17546,N_17324,N_17490);
nor U17547 (N_17547,N_17391,N_17265);
or U17548 (N_17548,N_17436,N_17433);
or U17549 (N_17549,N_17461,N_17252);
and U17550 (N_17550,N_17485,N_17458);
xnor U17551 (N_17551,N_17287,N_17309);
and U17552 (N_17552,N_17261,N_17481);
xnor U17553 (N_17553,N_17449,N_17302);
or U17554 (N_17554,N_17427,N_17422);
nand U17555 (N_17555,N_17328,N_17364);
nand U17556 (N_17556,N_17306,N_17462);
xor U17557 (N_17557,N_17439,N_17277);
and U17558 (N_17558,N_17471,N_17424);
nor U17559 (N_17559,N_17482,N_17259);
and U17560 (N_17560,N_17405,N_17392);
or U17561 (N_17561,N_17459,N_17435);
xnor U17562 (N_17562,N_17396,N_17456);
nor U17563 (N_17563,N_17466,N_17489);
and U17564 (N_17564,N_17290,N_17273);
xnor U17565 (N_17565,N_17285,N_17389);
nand U17566 (N_17566,N_17497,N_17444);
xnor U17567 (N_17567,N_17467,N_17282);
nand U17568 (N_17568,N_17274,N_17283);
or U17569 (N_17569,N_17486,N_17419);
or U17570 (N_17570,N_17295,N_17250);
xor U17571 (N_17571,N_17376,N_17463);
xnor U17572 (N_17572,N_17473,N_17348);
xnor U17573 (N_17573,N_17399,N_17284);
or U17574 (N_17574,N_17499,N_17305);
or U17575 (N_17575,N_17354,N_17493);
xnor U17576 (N_17576,N_17337,N_17367);
or U17577 (N_17577,N_17417,N_17401);
and U17578 (N_17578,N_17304,N_17412);
nor U17579 (N_17579,N_17338,N_17434);
nor U17580 (N_17580,N_17289,N_17327);
xor U17581 (N_17581,N_17432,N_17377);
and U17582 (N_17582,N_17494,N_17310);
nand U17583 (N_17583,N_17335,N_17394);
nor U17584 (N_17584,N_17390,N_17257);
or U17585 (N_17585,N_17292,N_17296);
nor U17586 (N_17586,N_17255,N_17281);
xor U17587 (N_17587,N_17455,N_17268);
or U17588 (N_17588,N_17329,N_17495);
nor U17589 (N_17589,N_17331,N_17413);
xor U17590 (N_17590,N_17361,N_17373);
nand U17591 (N_17591,N_17360,N_17297);
xnor U17592 (N_17592,N_17478,N_17350);
xnor U17593 (N_17593,N_17475,N_17451);
xnor U17594 (N_17594,N_17393,N_17379);
nand U17595 (N_17595,N_17349,N_17298);
nand U17596 (N_17596,N_17450,N_17313);
xnor U17597 (N_17597,N_17366,N_17380);
and U17598 (N_17598,N_17343,N_17491);
xor U17599 (N_17599,N_17382,N_17326);
and U17600 (N_17600,N_17480,N_17276);
or U17601 (N_17601,N_17464,N_17397);
nor U17602 (N_17602,N_17454,N_17271);
or U17603 (N_17603,N_17316,N_17363);
xor U17604 (N_17604,N_17414,N_17468);
nand U17605 (N_17605,N_17353,N_17472);
nor U17606 (N_17606,N_17476,N_17258);
nand U17607 (N_17607,N_17300,N_17251);
nand U17608 (N_17608,N_17321,N_17479);
or U17609 (N_17609,N_17320,N_17383);
nor U17610 (N_17610,N_17369,N_17488);
and U17611 (N_17611,N_17342,N_17307);
and U17612 (N_17612,N_17352,N_17386);
nor U17613 (N_17613,N_17443,N_17357);
and U17614 (N_17614,N_17426,N_17356);
xnor U17615 (N_17615,N_17340,N_17378);
and U17616 (N_17616,N_17322,N_17410);
and U17617 (N_17617,N_17428,N_17334);
or U17618 (N_17618,N_17416,N_17319);
xnor U17619 (N_17619,N_17368,N_17398);
xor U17620 (N_17620,N_17280,N_17346);
nor U17621 (N_17621,N_17355,N_17400);
or U17622 (N_17622,N_17278,N_17341);
nand U17623 (N_17623,N_17308,N_17362);
or U17624 (N_17624,N_17370,N_17387);
xor U17625 (N_17625,N_17364,N_17323);
and U17626 (N_17626,N_17483,N_17273);
xor U17627 (N_17627,N_17494,N_17255);
or U17628 (N_17628,N_17268,N_17307);
xnor U17629 (N_17629,N_17372,N_17275);
and U17630 (N_17630,N_17353,N_17385);
or U17631 (N_17631,N_17265,N_17383);
xnor U17632 (N_17632,N_17289,N_17419);
xor U17633 (N_17633,N_17397,N_17423);
nor U17634 (N_17634,N_17260,N_17359);
or U17635 (N_17635,N_17415,N_17320);
nand U17636 (N_17636,N_17278,N_17423);
and U17637 (N_17637,N_17418,N_17494);
nor U17638 (N_17638,N_17465,N_17329);
nor U17639 (N_17639,N_17341,N_17331);
nor U17640 (N_17640,N_17476,N_17323);
or U17641 (N_17641,N_17384,N_17427);
xor U17642 (N_17642,N_17323,N_17260);
or U17643 (N_17643,N_17293,N_17343);
nand U17644 (N_17644,N_17340,N_17260);
xnor U17645 (N_17645,N_17467,N_17406);
or U17646 (N_17646,N_17476,N_17453);
or U17647 (N_17647,N_17333,N_17408);
nor U17648 (N_17648,N_17375,N_17456);
nor U17649 (N_17649,N_17403,N_17377);
nand U17650 (N_17650,N_17386,N_17293);
xor U17651 (N_17651,N_17317,N_17322);
nand U17652 (N_17652,N_17400,N_17385);
nand U17653 (N_17653,N_17250,N_17267);
and U17654 (N_17654,N_17275,N_17493);
nor U17655 (N_17655,N_17337,N_17410);
xnor U17656 (N_17656,N_17265,N_17339);
xor U17657 (N_17657,N_17442,N_17449);
nor U17658 (N_17658,N_17275,N_17458);
or U17659 (N_17659,N_17254,N_17320);
xor U17660 (N_17660,N_17345,N_17461);
xnor U17661 (N_17661,N_17412,N_17272);
xor U17662 (N_17662,N_17291,N_17431);
or U17663 (N_17663,N_17336,N_17374);
nor U17664 (N_17664,N_17350,N_17421);
xnor U17665 (N_17665,N_17270,N_17441);
xnor U17666 (N_17666,N_17348,N_17336);
nor U17667 (N_17667,N_17357,N_17423);
xnor U17668 (N_17668,N_17376,N_17488);
xor U17669 (N_17669,N_17447,N_17330);
or U17670 (N_17670,N_17320,N_17425);
nor U17671 (N_17671,N_17282,N_17489);
nor U17672 (N_17672,N_17473,N_17316);
and U17673 (N_17673,N_17263,N_17498);
nor U17674 (N_17674,N_17322,N_17399);
and U17675 (N_17675,N_17281,N_17329);
nand U17676 (N_17676,N_17349,N_17360);
or U17677 (N_17677,N_17367,N_17355);
nand U17678 (N_17678,N_17395,N_17354);
nor U17679 (N_17679,N_17334,N_17489);
and U17680 (N_17680,N_17478,N_17286);
nor U17681 (N_17681,N_17316,N_17255);
or U17682 (N_17682,N_17394,N_17317);
xor U17683 (N_17683,N_17435,N_17395);
xnor U17684 (N_17684,N_17369,N_17467);
nor U17685 (N_17685,N_17415,N_17349);
nor U17686 (N_17686,N_17499,N_17420);
nand U17687 (N_17687,N_17256,N_17393);
xnor U17688 (N_17688,N_17286,N_17396);
nand U17689 (N_17689,N_17485,N_17320);
nand U17690 (N_17690,N_17383,N_17442);
xor U17691 (N_17691,N_17334,N_17422);
xnor U17692 (N_17692,N_17441,N_17417);
and U17693 (N_17693,N_17408,N_17316);
nand U17694 (N_17694,N_17286,N_17475);
nor U17695 (N_17695,N_17399,N_17326);
xnor U17696 (N_17696,N_17264,N_17493);
and U17697 (N_17697,N_17328,N_17287);
nand U17698 (N_17698,N_17463,N_17358);
or U17699 (N_17699,N_17464,N_17371);
xnor U17700 (N_17700,N_17332,N_17497);
nand U17701 (N_17701,N_17344,N_17267);
nand U17702 (N_17702,N_17339,N_17397);
and U17703 (N_17703,N_17434,N_17378);
xnor U17704 (N_17704,N_17280,N_17482);
nand U17705 (N_17705,N_17309,N_17484);
nor U17706 (N_17706,N_17431,N_17329);
xnor U17707 (N_17707,N_17420,N_17314);
nor U17708 (N_17708,N_17456,N_17441);
xnor U17709 (N_17709,N_17410,N_17482);
xnor U17710 (N_17710,N_17491,N_17291);
nand U17711 (N_17711,N_17435,N_17475);
and U17712 (N_17712,N_17438,N_17281);
nand U17713 (N_17713,N_17274,N_17356);
nor U17714 (N_17714,N_17387,N_17386);
or U17715 (N_17715,N_17371,N_17352);
and U17716 (N_17716,N_17277,N_17435);
and U17717 (N_17717,N_17465,N_17299);
or U17718 (N_17718,N_17429,N_17485);
or U17719 (N_17719,N_17255,N_17358);
nor U17720 (N_17720,N_17492,N_17301);
or U17721 (N_17721,N_17309,N_17342);
nor U17722 (N_17722,N_17303,N_17356);
or U17723 (N_17723,N_17410,N_17406);
xnor U17724 (N_17724,N_17449,N_17275);
xor U17725 (N_17725,N_17478,N_17447);
xor U17726 (N_17726,N_17272,N_17438);
and U17727 (N_17727,N_17328,N_17394);
nor U17728 (N_17728,N_17282,N_17465);
nor U17729 (N_17729,N_17462,N_17382);
and U17730 (N_17730,N_17304,N_17283);
and U17731 (N_17731,N_17416,N_17294);
xor U17732 (N_17732,N_17263,N_17280);
nand U17733 (N_17733,N_17455,N_17469);
nor U17734 (N_17734,N_17479,N_17325);
or U17735 (N_17735,N_17491,N_17403);
and U17736 (N_17736,N_17497,N_17347);
nand U17737 (N_17737,N_17337,N_17284);
or U17738 (N_17738,N_17279,N_17411);
xor U17739 (N_17739,N_17389,N_17443);
xor U17740 (N_17740,N_17284,N_17424);
xor U17741 (N_17741,N_17407,N_17400);
nor U17742 (N_17742,N_17297,N_17361);
nand U17743 (N_17743,N_17411,N_17358);
nand U17744 (N_17744,N_17268,N_17488);
or U17745 (N_17745,N_17372,N_17295);
nor U17746 (N_17746,N_17403,N_17481);
xor U17747 (N_17747,N_17438,N_17481);
xnor U17748 (N_17748,N_17463,N_17309);
nand U17749 (N_17749,N_17416,N_17428);
or U17750 (N_17750,N_17661,N_17598);
and U17751 (N_17751,N_17529,N_17715);
xor U17752 (N_17752,N_17698,N_17682);
or U17753 (N_17753,N_17747,N_17578);
nand U17754 (N_17754,N_17511,N_17500);
nand U17755 (N_17755,N_17561,N_17729);
nor U17756 (N_17756,N_17536,N_17604);
or U17757 (N_17757,N_17530,N_17683);
and U17758 (N_17758,N_17728,N_17641);
xnor U17759 (N_17759,N_17508,N_17717);
and U17760 (N_17760,N_17583,N_17581);
nand U17761 (N_17761,N_17606,N_17677);
or U17762 (N_17762,N_17587,N_17734);
xor U17763 (N_17763,N_17648,N_17691);
xnor U17764 (N_17764,N_17722,N_17611);
nand U17765 (N_17765,N_17615,N_17501);
xor U17766 (N_17766,N_17733,N_17541);
nor U17767 (N_17767,N_17674,N_17663);
nor U17768 (N_17768,N_17599,N_17547);
xor U17769 (N_17769,N_17580,N_17658);
nand U17770 (N_17770,N_17653,N_17689);
and U17771 (N_17771,N_17585,N_17656);
nor U17772 (N_17772,N_17708,N_17525);
and U17773 (N_17773,N_17667,N_17523);
nor U17774 (N_17774,N_17579,N_17589);
nand U17775 (N_17775,N_17614,N_17666);
xor U17776 (N_17776,N_17569,N_17694);
nor U17777 (N_17777,N_17506,N_17590);
or U17778 (N_17778,N_17636,N_17644);
or U17779 (N_17779,N_17533,N_17697);
and U17780 (N_17780,N_17515,N_17576);
xnor U17781 (N_17781,N_17516,N_17574);
or U17782 (N_17782,N_17588,N_17711);
or U17783 (N_17783,N_17625,N_17684);
nand U17784 (N_17784,N_17745,N_17713);
and U17785 (N_17785,N_17539,N_17612);
nand U17786 (N_17786,N_17730,N_17646);
or U17787 (N_17787,N_17743,N_17749);
xor U17788 (N_17788,N_17671,N_17584);
or U17789 (N_17789,N_17703,N_17701);
nor U17790 (N_17790,N_17527,N_17610);
and U17791 (N_17791,N_17563,N_17650);
nand U17792 (N_17792,N_17723,N_17744);
nand U17793 (N_17793,N_17595,N_17540);
xor U17794 (N_17794,N_17657,N_17572);
nor U17795 (N_17795,N_17522,N_17709);
and U17796 (N_17796,N_17686,N_17559);
nor U17797 (N_17797,N_17502,N_17637);
nor U17798 (N_17798,N_17738,N_17736);
or U17799 (N_17799,N_17554,N_17635);
nand U17800 (N_17800,N_17687,N_17543);
xor U17801 (N_17801,N_17514,N_17600);
and U17802 (N_17802,N_17647,N_17741);
nor U17803 (N_17803,N_17630,N_17685);
nor U17804 (N_17804,N_17654,N_17557);
nand U17805 (N_17805,N_17655,N_17725);
and U17806 (N_17806,N_17714,N_17603);
nor U17807 (N_17807,N_17699,N_17510);
xor U17808 (N_17808,N_17720,N_17532);
or U17809 (N_17809,N_17681,N_17621);
or U17810 (N_17810,N_17537,N_17593);
or U17811 (N_17811,N_17695,N_17690);
nor U17812 (N_17812,N_17732,N_17672);
xor U17813 (N_17813,N_17507,N_17705);
and U17814 (N_17814,N_17602,N_17716);
nor U17815 (N_17815,N_17545,N_17660);
and U17816 (N_17816,N_17740,N_17624);
or U17817 (N_17817,N_17575,N_17565);
and U17818 (N_17818,N_17638,N_17632);
nor U17819 (N_17819,N_17582,N_17634);
or U17820 (N_17820,N_17727,N_17601);
or U17821 (N_17821,N_17626,N_17577);
xor U17822 (N_17822,N_17618,N_17571);
nor U17823 (N_17823,N_17556,N_17519);
nand U17824 (N_17824,N_17718,N_17586);
nor U17825 (N_17825,N_17649,N_17668);
and U17826 (N_17826,N_17679,N_17700);
nor U17827 (N_17827,N_17573,N_17549);
and U17828 (N_17828,N_17550,N_17629);
nor U17829 (N_17829,N_17628,N_17704);
or U17830 (N_17830,N_17693,N_17617);
xor U17831 (N_17831,N_17662,N_17607);
or U17832 (N_17832,N_17568,N_17513);
nand U17833 (N_17833,N_17639,N_17521);
nand U17834 (N_17834,N_17702,N_17651);
and U17835 (N_17835,N_17596,N_17664);
or U17836 (N_17836,N_17517,N_17706);
or U17837 (N_17837,N_17564,N_17640);
xnor U17838 (N_17838,N_17562,N_17544);
nand U17839 (N_17839,N_17542,N_17742);
or U17840 (N_17840,N_17616,N_17567);
xor U17841 (N_17841,N_17594,N_17546);
and U17842 (N_17842,N_17528,N_17692);
xnor U17843 (N_17843,N_17707,N_17675);
nand U17844 (N_17844,N_17659,N_17620);
nand U17845 (N_17845,N_17652,N_17731);
nor U17846 (N_17846,N_17680,N_17538);
or U17847 (N_17847,N_17597,N_17710);
nor U17848 (N_17848,N_17552,N_17609);
or U17849 (N_17849,N_17592,N_17505);
nor U17850 (N_17850,N_17623,N_17670);
nand U17851 (N_17851,N_17534,N_17719);
nand U17852 (N_17852,N_17526,N_17643);
nand U17853 (N_17853,N_17746,N_17673);
or U17854 (N_17854,N_17535,N_17605);
xor U17855 (N_17855,N_17678,N_17608);
and U17856 (N_17856,N_17633,N_17551);
or U17857 (N_17857,N_17631,N_17553);
nor U17858 (N_17858,N_17665,N_17613);
xnor U17859 (N_17859,N_17555,N_17712);
xnor U17860 (N_17860,N_17627,N_17531);
nor U17861 (N_17861,N_17676,N_17558);
and U17862 (N_17862,N_17622,N_17509);
xor U17863 (N_17863,N_17520,N_17669);
and U17864 (N_17864,N_17726,N_17721);
xnor U17865 (N_17865,N_17696,N_17548);
xor U17866 (N_17866,N_17748,N_17504);
nand U17867 (N_17867,N_17619,N_17566);
nand U17868 (N_17868,N_17645,N_17560);
and U17869 (N_17869,N_17739,N_17518);
or U17870 (N_17870,N_17524,N_17503);
nand U17871 (N_17871,N_17737,N_17735);
nor U17872 (N_17872,N_17512,N_17591);
nor U17873 (N_17873,N_17724,N_17570);
nor U17874 (N_17874,N_17688,N_17642);
xor U17875 (N_17875,N_17657,N_17686);
xor U17876 (N_17876,N_17698,N_17723);
and U17877 (N_17877,N_17644,N_17589);
or U17878 (N_17878,N_17740,N_17647);
or U17879 (N_17879,N_17711,N_17528);
nor U17880 (N_17880,N_17510,N_17641);
or U17881 (N_17881,N_17659,N_17580);
xnor U17882 (N_17882,N_17665,N_17676);
nand U17883 (N_17883,N_17544,N_17532);
nand U17884 (N_17884,N_17709,N_17508);
nor U17885 (N_17885,N_17695,N_17617);
and U17886 (N_17886,N_17733,N_17745);
and U17887 (N_17887,N_17501,N_17559);
and U17888 (N_17888,N_17667,N_17647);
nor U17889 (N_17889,N_17703,N_17715);
and U17890 (N_17890,N_17592,N_17525);
and U17891 (N_17891,N_17639,N_17586);
nor U17892 (N_17892,N_17711,N_17559);
and U17893 (N_17893,N_17659,N_17598);
nand U17894 (N_17894,N_17716,N_17738);
or U17895 (N_17895,N_17700,N_17527);
nor U17896 (N_17896,N_17536,N_17724);
or U17897 (N_17897,N_17517,N_17685);
xnor U17898 (N_17898,N_17749,N_17554);
nor U17899 (N_17899,N_17685,N_17518);
nand U17900 (N_17900,N_17507,N_17517);
nand U17901 (N_17901,N_17658,N_17586);
nor U17902 (N_17902,N_17748,N_17626);
xnor U17903 (N_17903,N_17662,N_17521);
nor U17904 (N_17904,N_17509,N_17579);
nor U17905 (N_17905,N_17514,N_17615);
nor U17906 (N_17906,N_17672,N_17647);
or U17907 (N_17907,N_17677,N_17524);
xnor U17908 (N_17908,N_17536,N_17576);
xnor U17909 (N_17909,N_17739,N_17533);
xnor U17910 (N_17910,N_17709,N_17525);
xor U17911 (N_17911,N_17601,N_17593);
nor U17912 (N_17912,N_17716,N_17533);
or U17913 (N_17913,N_17507,N_17646);
or U17914 (N_17914,N_17705,N_17679);
xor U17915 (N_17915,N_17642,N_17527);
xor U17916 (N_17916,N_17623,N_17680);
nand U17917 (N_17917,N_17676,N_17528);
nand U17918 (N_17918,N_17702,N_17515);
xor U17919 (N_17919,N_17637,N_17515);
nor U17920 (N_17920,N_17574,N_17525);
and U17921 (N_17921,N_17631,N_17505);
nand U17922 (N_17922,N_17525,N_17502);
or U17923 (N_17923,N_17633,N_17734);
xnor U17924 (N_17924,N_17606,N_17549);
xnor U17925 (N_17925,N_17599,N_17677);
nor U17926 (N_17926,N_17581,N_17602);
xor U17927 (N_17927,N_17610,N_17526);
or U17928 (N_17928,N_17719,N_17562);
nor U17929 (N_17929,N_17738,N_17628);
or U17930 (N_17930,N_17725,N_17717);
xor U17931 (N_17931,N_17506,N_17725);
xnor U17932 (N_17932,N_17646,N_17662);
and U17933 (N_17933,N_17631,N_17524);
or U17934 (N_17934,N_17749,N_17596);
or U17935 (N_17935,N_17706,N_17586);
or U17936 (N_17936,N_17714,N_17575);
xnor U17937 (N_17937,N_17529,N_17709);
nor U17938 (N_17938,N_17743,N_17695);
or U17939 (N_17939,N_17578,N_17636);
nor U17940 (N_17940,N_17565,N_17647);
and U17941 (N_17941,N_17565,N_17705);
nor U17942 (N_17942,N_17562,N_17653);
nand U17943 (N_17943,N_17679,N_17589);
and U17944 (N_17944,N_17509,N_17643);
xor U17945 (N_17945,N_17507,N_17583);
nor U17946 (N_17946,N_17721,N_17567);
nor U17947 (N_17947,N_17522,N_17736);
and U17948 (N_17948,N_17552,N_17721);
or U17949 (N_17949,N_17629,N_17633);
and U17950 (N_17950,N_17747,N_17595);
or U17951 (N_17951,N_17508,N_17549);
and U17952 (N_17952,N_17682,N_17644);
nand U17953 (N_17953,N_17596,N_17673);
or U17954 (N_17954,N_17561,N_17548);
and U17955 (N_17955,N_17623,N_17581);
nor U17956 (N_17956,N_17692,N_17624);
nand U17957 (N_17957,N_17521,N_17527);
nor U17958 (N_17958,N_17522,N_17534);
xnor U17959 (N_17959,N_17713,N_17582);
or U17960 (N_17960,N_17583,N_17614);
nand U17961 (N_17961,N_17651,N_17681);
nor U17962 (N_17962,N_17608,N_17571);
nand U17963 (N_17963,N_17622,N_17582);
xnor U17964 (N_17964,N_17732,N_17706);
nor U17965 (N_17965,N_17652,N_17516);
nand U17966 (N_17966,N_17520,N_17745);
xnor U17967 (N_17967,N_17626,N_17677);
nand U17968 (N_17968,N_17566,N_17633);
xnor U17969 (N_17969,N_17653,N_17674);
nor U17970 (N_17970,N_17531,N_17520);
nand U17971 (N_17971,N_17593,N_17736);
and U17972 (N_17972,N_17701,N_17732);
and U17973 (N_17973,N_17534,N_17578);
and U17974 (N_17974,N_17653,N_17599);
nand U17975 (N_17975,N_17533,N_17522);
nor U17976 (N_17976,N_17529,N_17681);
nor U17977 (N_17977,N_17741,N_17702);
and U17978 (N_17978,N_17747,N_17562);
and U17979 (N_17979,N_17542,N_17520);
nor U17980 (N_17980,N_17659,N_17618);
nand U17981 (N_17981,N_17679,N_17548);
or U17982 (N_17982,N_17594,N_17593);
or U17983 (N_17983,N_17657,N_17518);
or U17984 (N_17984,N_17595,N_17745);
nand U17985 (N_17985,N_17681,N_17712);
and U17986 (N_17986,N_17521,N_17562);
and U17987 (N_17987,N_17604,N_17520);
or U17988 (N_17988,N_17733,N_17556);
xor U17989 (N_17989,N_17578,N_17731);
nand U17990 (N_17990,N_17740,N_17519);
xnor U17991 (N_17991,N_17643,N_17739);
and U17992 (N_17992,N_17601,N_17642);
or U17993 (N_17993,N_17677,N_17712);
nand U17994 (N_17994,N_17588,N_17539);
and U17995 (N_17995,N_17611,N_17550);
nand U17996 (N_17996,N_17562,N_17567);
xor U17997 (N_17997,N_17641,N_17559);
nor U17998 (N_17998,N_17500,N_17617);
or U17999 (N_17999,N_17559,N_17618);
or U18000 (N_18000,N_17812,N_17826);
xnor U18001 (N_18001,N_17926,N_17795);
nor U18002 (N_18002,N_17851,N_17901);
or U18003 (N_18003,N_17832,N_17854);
nand U18004 (N_18004,N_17923,N_17824);
xnor U18005 (N_18005,N_17968,N_17762);
nand U18006 (N_18006,N_17805,N_17966);
and U18007 (N_18007,N_17770,N_17972);
xor U18008 (N_18008,N_17889,N_17895);
nor U18009 (N_18009,N_17911,N_17856);
nor U18010 (N_18010,N_17767,N_17752);
xnor U18011 (N_18011,N_17891,N_17995);
xnor U18012 (N_18012,N_17804,N_17865);
nand U18013 (N_18013,N_17984,N_17783);
xnor U18014 (N_18014,N_17959,N_17753);
xor U18015 (N_18015,N_17806,N_17971);
nand U18016 (N_18016,N_17986,N_17949);
and U18017 (N_18017,N_17933,N_17834);
or U18018 (N_18018,N_17833,N_17827);
xnor U18019 (N_18019,N_17978,N_17788);
nor U18020 (N_18020,N_17758,N_17820);
nand U18021 (N_18021,N_17922,N_17957);
xor U18022 (N_18022,N_17835,N_17967);
or U18023 (N_18023,N_17792,N_17838);
xor U18024 (N_18024,N_17796,N_17886);
xor U18025 (N_18025,N_17987,N_17862);
nor U18026 (N_18026,N_17893,N_17840);
nor U18027 (N_18027,N_17777,N_17964);
xnor U18028 (N_18028,N_17844,N_17771);
nand U18029 (N_18029,N_17808,N_17936);
nor U18030 (N_18030,N_17831,N_17821);
xnor U18031 (N_18031,N_17800,N_17801);
xor U18032 (N_18032,N_17892,N_17845);
xnor U18033 (N_18033,N_17816,N_17785);
nor U18034 (N_18034,N_17823,N_17962);
nand U18035 (N_18035,N_17815,N_17946);
or U18036 (N_18036,N_17942,N_17861);
nor U18037 (N_18037,N_17905,N_17951);
or U18038 (N_18038,N_17909,N_17934);
and U18039 (N_18039,N_17954,N_17953);
nor U18040 (N_18040,N_17890,N_17996);
or U18041 (N_18041,N_17866,N_17882);
xor U18042 (N_18042,N_17784,N_17841);
nand U18043 (N_18043,N_17927,N_17880);
xor U18044 (N_18044,N_17774,N_17975);
or U18045 (N_18045,N_17868,N_17798);
nor U18046 (N_18046,N_17907,N_17988);
nor U18047 (N_18047,N_17791,N_17960);
xor U18048 (N_18048,N_17750,N_17813);
nand U18049 (N_18049,N_17846,N_17983);
and U18050 (N_18050,N_17903,N_17981);
xnor U18051 (N_18051,N_17908,N_17778);
nor U18052 (N_18052,N_17852,N_17755);
and U18053 (N_18053,N_17918,N_17974);
or U18054 (N_18054,N_17982,N_17764);
xnor U18055 (N_18055,N_17786,N_17828);
xnor U18056 (N_18056,N_17759,N_17937);
or U18057 (N_18057,N_17958,N_17754);
nand U18058 (N_18058,N_17929,N_17941);
xor U18059 (N_18059,N_17781,N_17979);
nand U18060 (N_18060,N_17789,N_17990);
nor U18061 (N_18061,N_17896,N_17775);
xnor U18062 (N_18062,N_17904,N_17883);
nor U18063 (N_18063,N_17760,N_17874);
xnor U18064 (N_18064,N_17939,N_17877);
nand U18065 (N_18065,N_17787,N_17894);
nand U18066 (N_18066,N_17859,N_17756);
nand U18067 (N_18067,N_17860,N_17961);
nor U18068 (N_18068,N_17999,N_17836);
nand U18069 (N_18069,N_17915,N_17963);
nor U18070 (N_18070,N_17769,N_17952);
and U18071 (N_18071,N_17849,N_17879);
xor U18072 (N_18072,N_17970,N_17873);
xnor U18073 (N_18073,N_17870,N_17817);
nor U18074 (N_18074,N_17766,N_17761);
nor U18075 (N_18075,N_17797,N_17980);
and U18076 (N_18076,N_17848,N_17869);
nand U18077 (N_18077,N_17768,N_17878);
nand U18078 (N_18078,N_17765,N_17940);
nand U18079 (N_18079,N_17921,N_17857);
xor U18080 (N_18080,N_17855,N_17867);
nand U18081 (N_18081,N_17803,N_17910);
nand U18082 (N_18082,N_17899,N_17898);
xor U18083 (N_18083,N_17998,N_17807);
nor U18084 (N_18084,N_17818,N_17794);
and U18085 (N_18085,N_17997,N_17948);
nand U18086 (N_18086,N_17914,N_17757);
and U18087 (N_18087,N_17779,N_17973);
xor U18088 (N_18088,N_17938,N_17932);
xor U18089 (N_18089,N_17843,N_17944);
nor U18090 (N_18090,N_17822,N_17994);
or U18091 (N_18091,N_17976,N_17943);
nor U18092 (N_18092,N_17811,N_17920);
nor U18093 (N_18093,N_17763,N_17989);
nor U18094 (N_18094,N_17993,N_17876);
or U18095 (N_18095,N_17965,N_17912);
or U18096 (N_18096,N_17888,N_17772);
nand U18097 (N_18097,N_17992,N_17985);
nand U18098 (N_18098,N_17925,N_17793);
nand U18099 (N_18099,N_17847,N_17881);
or U18100 (N_18100,N_17799,N_17819);
xnor U18101 (N_18101,N_17945,N_17842);
xnor U18102 (N_18102,N_17853,N_17947);
and U18103 (N_18103,N_17897,N_17825);
or U18104 (N_18104,N_17900,N_17935);
nor U18105 (N_18105,N_17928,N_17991);
nor U18106 (N_18106,N_17776,N_17885);
xnor U18107 (N_18107,N_17814,N_17875);
or U18108 (N_18108,N_17956,N_17858);
and U18109 (N_18109,N_17864,N_17751);
nor U18110 (N_18110,N_17837,N_17773);
or U18111 (N_18111,N_17780,N_17887);
or U18112 (N_18112,N_17863,N_17850);
nand U18113 (N_18113,N_17839,N_17913);
nor U18114 (N_18114,N_17810,N_17809);
xor U18115 (N_18115,N_17802,N_17902);
and U18116 (N_18116,N_17950,N_17977);
xnor U18117 (N_18117,N_17830,N_17916);
or U18118 (N_18118,N_17871,N_17955);
nor U18119 (N_18119,N_17829,N_17782);
and U18120 (N_18120,N_17924,N_17906);
and U18121 (N_18121,N_17969,N_17930);
nand U18122 (N_18122,N_17931,N_17872);
xnor U18123 (N_18123,N_17790,N_17917);
and U18124 (N_18124,N_17884,N_17919);
nor U18125 (N_18125,N_17915,N_17885);
and U18126 (N_18126,N_17854,N_17752);
nand U18127 (N_18127,N_17978,N_17905);
and U18128 (N_18128,N_17890,N_17851);
nor U18129 (N_18129,N_17818,N_17905);
and U18130 (N_18130,N_17934,N_17846);
nand U18131 (N_18131,N_17997,N_17797);
xnor U18132 (N_18132,N_17798,N_17872);
or U18133 (N_18133,N_17942,N_17953);
nor U18134 (N_18134,N_17970,N_17863);
and U18135 (N_18135,N_17830,N_17785);
nand U18136 (N_18136,N_17980,N_17822);
xnor U18137 (N_18137,N_17993,N_17883);
xnor U18138 (N_18138,N_17886,N_17982);
nand U18139 (N_18139,N_17979,N_17926);
nor U18140 (N_18140,N_17876,N_17770);
nand U18141 (N_18141,N_17769,N_17950);
nand U18142 (N_18142,N_17955,N_17965);
or U18143 (N_18143,N_17784,N_17754);
nor U18144 (N_18144,N_17880,N_17782);
xor U18145 (N_18145,N_17765,N_17905);
xnor U18146 (N_18146,N_17910,N_17835);
nor U18147 (N_18147,N_17886,N_17938);
nor U18148 (N_18148,N_17753,N_17868);
or U18149 (N_18149,N_17768,N_17865);
and U18150 (N_18150,N_17939,N_17797);
or U18151 (N_18151,N_17857,N_17953);
nor U18152 (N_18152,N_17808,N_17896);
nand U18153 (N_18153,N_17798,N_17847);
nor U18154 (N_18154,N_17813,N_17990);
xor U18155 (N_18155,N_17896,N_17852);
nand U18156 (N_18156,N_17773,N_17791);
nand U18157 (N_18157,N_17751,N_17898);
xor U18158 (N_18158,N_17772,N_17808);
nor U18159 (N_18159,N_17899,N_17808);
xnor U18160 (N_18160,N_17861,N_17975);
and U18161 (N_18161,N_17849,N_17912);
nand U18162 (N_18162,N_17812,N_17935);
nor U18163 (N_18163,N_17757,N_17763);
nand U18164 (N_18164,N_17861,N_17786);
xnor U18165 (N_18165,N_17792,N_17822);
and U18166 (N_18166,N_17984,N_17967);
xnor U18167 (N_18167,N_17815,N_17868);
nor U18168 (N_18168,N_17790,N_17871);
xor U18169 (N_18169,N_17991,N_17934);
and U18170 (N_18170,N_17814,N_17759);
and U18171 (N_18171,N_17918,N_17927);
nand U18172 (N_18172,N_17803,N_17989);
nand U18173 (N_18173,N_17904,N_17965);
nor U18174 (N_18174,N_17786,N_17962);
and U18175 (N_18175,N_17838,N_17979);
nor U18176 (N_18176,N_17773,N_17828);
and U18177 (N_18177,N_17924,N_17767);
and U18178 (N_18178,N_17781,N_17831);
nand U18179 (N_18179,N_17791,N_17814);
xor U18180 (N_18180,N_17905,N_17918);
nor U18181 (N_18181,N_17761,N_17776);
nand U18182 (N_18182,N_17867,N_17988);
xnor U18183 (N_18183,N_17773,N_17965);
nor U18184 (N_18184,N_17792,N_17953);
and U18185 (N_18185,N_17895,N_17920);
xnor U18186 (N_18186,N_17809,N_17895);
nand U18187 (N_18187,N_17895,N_17763);
nor U18188 (N_18188,N_17777,N_17915);
and U18189 (N_18189,N_17917,N_17882);
nor U18190 (N_18190,N_17985,N_17794);
or U18191 (N_18191,N_17929,N_17762);
nand U18192 (N_18192,N_17961,N_17854);
nor U18193 (N_18193,N_17802,N_17895);
and U18194 (N_18194,N_17811,N_17776);
nor U18195 (N_18195,N_17863,N_17833);
nor U18196 (N_18196,N_17831,N_17899);
or U18197 (N_18197,N_17873,N_17846);
nand U18198 (N_18198,N_17806,N_17956);
nand U18199 (N_18199,N_17973,N_17900);
xnor U18200 (N_18200,N_17764,N_17783);
nor U18201 (N_18201,N_17884,N_17815);
and U18202 (N_18202,N_17984,N_17989);
or U18203 (N_18203,N_17818,N_17826);
or U18204 (N_18204,N_17937,N_17830);
or U18205 (N_18205,N_17764,N_17919);
nand U18206 (N_18206,N_17941,N_17824);
nor U18207 (N_18207,N_17917,N_17929);
xnor U18208 (N_18208,N_17983,N_17807);
xor U18209 (N_18209,N_17760,N_17863);
nor U18210 (N_18210,N_17883,N_17803);
and U18211 (N_18211,N_17814,N_17855);
nand U18212 (N_18212,N_17851,N_17813);
or U18213 (N_18213,N_17929,N_17798);
nor U18214 (N_18214,N_17819,N_17927);
nor U18215 (N_18215,N_17790,N_17986);
and U18216 (N_18216,N_17964,N_17943);
nand U18217 (N_18217,N_17970,N_17929);
xor U18218 (N_18218,N_17880,N_17829);
nor U18219 (N_18219,N_17910,N_17793);
or U18220 (N_18220,N_17940,N_17995);
nor U18221 (N_18221,N_17793,N_17776);
nor U18222 (N_18222,N_17769,N_17940);
nand U18223 (N_18223,N_17767,N_17994);
xnor U18224 (N_18224,N_17831,N_17898);
or U18225 (N_18225,N_17866,N_17751);
nand U18226 (N_18226,N_17858,N_17874);
nand U18227 (N_18227,N_17934,N_17752);
nand U18228 (N_18228,N_17912,N_17945);
xor U18229 (N_18229,N_17818,N_17887);
nor U18230 (N_18230,N_17818,N_17892);
nand U18231 (N_18231,N_17815,N_17798);
or U18232 (N_18232,N_17796,N_17947);
and U18233 (N_18233,N_17907,N_17997);
and U18234 (N_18234,N_17770,N_17808);
and U18235 (N_18235,N_17847,N_17898);
and U18236 (N_18236,N_17920,N_17947);
nor U18237 (N_18237,N_17894,N_17982);
or U18238 (N_18238,N_17792,N_17955);
nand U18239 (N_18239,N_17808,N_17833);
and U18240 (N_18240,N_17873,N_17969);
or U18241 (N_18241,N_17909,N_17971);
nor U18242 (N_18242,N_17810,N_17756);
nor U18243 (N_18243,N_17901,N_17750);
or U18244 (N_18244,N_17914,N_17879);
and U18245 (N_18245,N_17760,N_17821);
xor U18246 (N_18246,N_17932,N_17889);
or U18247 (N_18247,N_17794,N_17979);
nand U18248 (N_18248,N_17919,N_17810);
nand U18249 (N_18249,N_17829,N_17940);
or U18250 (N_18250,N_18010,N_18044);
or U18251 (N_18251,N_18230,N_18110);
and U18252 (N_18252,N_18056,N_18029);
or U18253 (N_18253,N_18224,N_18014);
and U18254 (N_18254,N_18189,N_18012);
and U18255 (N_18255,N_18239,N_18125);
and U18256 (N_18256,N_18178,N_18211);
or U18257 (N_18257,N_18031,N_18115);
or U18258 (N_18258,N_18076,N_18111);
or U18259 (N_18259,N_18078,N_18164);
nor U18260 (N_18260,N_18204,N_18084);
xor U18261 (N_18261,N_18191,N_18124);
xor U18262 (N_18262,N_18062,N_18108);
or U18263 (N_18263,N_18158,N_18153);
xor U18264 (N_18264,N_18049,N_18024);
xnor U18265 (N_18265,N_18186,N_18120);
nand U18266 (N_18266,N_18068,N_18094);
nor U18267 (N_18267,N_18140,N_18098);
nand U18268 (N_18268,N_18074,N_18228);
or U18269 (N_18269,N_18244,N_18223);
xnor U18270 (N_18270,N_18053,N_18166);
nor U18271 (N_18271,N_18163,N_18090);
nand U18272 (N_18272,N_18041,N_18036);
nand U18273 (N_18273,N_18179,N_18018);
nand U18274 (N_18274,N_18180,N_18055);
nand U18275 (N_18275,N_18075,N_18217);
nand U18276 (N_18276,N_18088,N_18023);
or U18277 (N_18277,N_18019,N_18127);
or U18278 (N_18278,N_18071,N_18199);
xor U18279 (N_18279,N_18060,N_18025);
nand U18280 (N_18280,N_18006,N_18150);
nor U18281 (N_18281,N_18141,N_18231);
nor U18282 (N_18282,N_18149,N_18190);
nor U18283 (N_18283,N_18136,N_18194);
and U18284 (N_18284,N_18126,N_18181);
nand U18285 (N_18285,N_18128,N_18066);
xnor U18286 (N_18286,N_18214,N_18097);
xnor U18287 (N_18287,N_18184,N_18236);
and U18288 (N_18288,N_18045,N_18083);
and U18289 (N_18289,N_18104,N_18057);
xor U18290 (N_18290,N_18226,N_18048);
or U18291 (N_18291,N_18109,N_18095);
xor U18292 (N_18292,N_18210,N_18047);
nor U18293 (N_18293,N_18129,N_18195);
nor U18294 (N_18294,N_18234,N_18196);
xor U18295 (N_18295,N_18159,N_18064);
and U18296 (N_18296,N_18145,N_18119);
and U18297 (N_18297,N_18246,N_18212);
xor U18298 (N_18298,N_18034,N_18209);
and U18299 (N_18299,N_18201,N_18081);
nor U18300 (N_18300,N_18116,N_18219);
and U18301 (N_18301,N_18221,N_18156);
nor U18302 (N_18302,N_18168,N_18051);
nor U18303 (N_18303,N_18146,N_18027);
and U18304 (N_18304,N_18121,N_18114);
or U18305 (N_18305,N_18085,N_18225);
and U18306 (N_18306,N_18105,N_18122);
xnor U18307 (N_18307,N_18020,N_18142);
or U18308 (N_18308,N_18002,N_18192);
or U18309 (N_18309,N_18089,N_18144);
nor U18310 (N_18310,N_18235,N_18118);
nand U18311 (N_18311,N_18007,N_18046);
nor U18312 (N_18312,N_18132,N_18169);
or U18313 (N_18313,N_18175,N_18240);
and U18314 (N_18314,N_18011,N_18208);
xor U18315 (N_18315,N_18037,N_18233);
and U18316 (N_18316,N_18147,N_18038);
or U18317 (N_18317,N_18102,N_18004);
or U18318 (N_18318,N_18139,N_18193);
nor U18319 (N_18319,N_18131,N_18096);
nand U18320 (N_18320,N_18151,N_18107);
nor U18321 (N_18321,N_18069,N_18249);
nor U18322 (N_18322,N_18148,N_18173);
or U18323 (N_18323,N_18213,N_18200);
or U18324 (N_18324,N_18227,N_18216);
or U18325 (N_18325,N_18187,N_18022);
xor U18326 (N_18326,N_18242,N_18185);
nor U18327 (N_18327,N_18157,N_18106);
nor U18328 (N_18328,N_18167,N_18205);
xor U18329 (N_18329,N_18113,N_18206);
nand U18330 (N_18330,N_18170,N_18160);
and U18331 (N_18331,N_18035,N_18203);
or U18332 (N_18332,N_18188,N_18073);
nor U18333 (N_18333,N_18134,N_18032);
nor U18334 (N_18334,N_18198,N_18135);
or U18335 (N_18335,N_18220,N_18183);
nand U18336 (N_18336,N_18174,N_18082);
or U18337 (N_18337,N_18162,N_18177);
nor U18338 (N_18338,N_18067,N_18016);
and U18339 (N_18339,N_18101,N_18063);
nand U18340 (N_18340,N_18015,N_18172);
and U18341 (N_18341,N_18197,N_18238);
nor U18342 (N_18342,N_18017,N_18061);
nor U18343 (N_18343,N_18072,N_18059);
xor U18344 (N_18344,N_18091,N_18026);
and U18345 (N_18345,N_18001,N_18039);
nor U18346 (N_18346,N_18161,N_18237);
nand U18347 (N_18347,N_18154,N_18058);
or U18348 (N_18348,N_18232,N_18042);
and U18349 (N_18349,N_18171,N_18099);
nand U18350 (N_18350,N_18138,N_18052);
xor U18351 (N_18351,N_18008,N_18079);
or U18352 (N_18352,N_18241,N_18092);
and U18353 (N_18353,N_18207,N_18086);
nor U18354 (N_18354,N_18133,N_18054);
xor U18355 (N_18355,N_18021,N_18117);
and U18356 (N_18356,N_18103,N_18202);
nand U18357 (N_18357,N_18245,N_18033);
or U18358 (N_18358,N_18229,N_18070);
xnor U18359 (N_18359,N_18000,N_18218);
nor U18360 (N_18360,N_18155,N_18080);
xor U18361 (N_18361,N_18222,N_18005);
or U18362 (N_18362,N_18165,N_18040);
nor U18363 (N_18363,N_18143,N_18028);
and U18364 (N_18364,N_18152,N_18003);
or U18365 (N_18365,N_18182,N_18093);
nor U18366 (N_18366,N_18030,N_18065);
xor U18367 (N_18367,N_18009,N_18050);
nor U18368 (N_18368,N_18043,N_18247);
xnor U18369 (N_18369,N_18215,N_18123);
or U18370 (N_18370,N_18243,N_18077);
or U18371 (N_18371,N_18176,N_18248);
and U18372 (N_18372,N_18087,N_18130);
and U18373 (N_18373,N_18013,N_18100);
nor U18374 (N_18374,N_18137,N_18112);
and U18375 (N_18375,N_18062,N_18240);
xor U18376 (N_18376,N_18135,N_18042);
nor U18377 (N_18377,N_18005,N_18064);
nor U18378 (N_18378,N_18189,N_18211);
nand U18379 (N_18379,N_18110,N_18201);
nand U18380 (N_18380,N_18158,N_18034);
and U18381 (N_18381,N_18173,N_18150);
or U18382 (N_18382,N_18219,N_18246);
and U18383 (N_18383,N_18108,N_18022);
xor U18384 (N_18384,N_18092,N_18132);
nand U18385 (N_18385,N_18078,N_18009);
and U18386 (N_18386,N_18009,N_18236);
or U18387 (N_18387,N_18203,N_18169);
and U18388 (N_18388,N_18173,N_18012);
nor U18389 (N_18389,N_18093,N_18229);
nand U18390 (N_18390,N_18056,N_18011);
nand U18391 (N_18391,N_18072,N_18045);
or U18392 (N_18392,N_18099,N_18047);
nor U18393 (N_18393,N_18084,N_18225);
nor U18394 (N_18394,N_18156,N_18219);
nand U18395 (N_18395,N_18100,N_18176);
and U18396 (N_18396,N_18241,N_18187);
or U18397 (N_18397,N_18144,N_18005);
xor U18398 (N_18398,N_18116,N_18078);
nor U18399 (N_18399,N_18012,N_18239);
xnor U18400 (N_18400,N_18189,N_18011);
xor U18401 (N_18401,N_18113,N_18026);
nand U18402 (N_18402,N_18197,N_18235);
xor U18403 (N_18403,N_18023,N_18243);
nand U18404 (N_18404,N_18118,N_18165);
and U18405 (N_18405,N_18213,N_18227);
nor U18406 (N_18406,N_18118,N_18083);
and U18407 (N_18407,N_18233,N_18212);
nor U18408 (N_18408,N_18128,N_18165);
xnor U18409 (N_18409,N_18127,N_18050);
or U18410 (N_18410,N_18062,N_18023);
nor U18411 (N_18411,N_18203,N_18048);
nor U18412 (N_18412,N_18207,N_18217);
nand U18413 (N_18413,N_18206,N_18019);
nor U18414 (N_18414,N_18136,N_18066);
and U18415 (N_18415,N_18064,N_18156);
nor U18416 (N_18416,N_18026,N_18042);
and U18417 (N_18417,N_18164,N_18014);
xor U18418 (N_18418,N_18115,N_18218);
nor U18419 (N_18419,N_18087,N_18207);
and U18420 (N_18420,N_18220,N_18122);
nor U18421 (N_18421,N_18059,N_18068);
xor U18422 (N_18422,N_18068,N_18142);
nor U18423 (N_18423,N_18074,N_18006);
nand U18424 (N_18424,N_18066,N_18163);
xor U18425 (N_18425,N_18070,N_18194);
nand U18426 (N_18426,N_18136,N_18086);
nor U18427 (N_18427,N_18201,N_18109);
xnor U18428 (N_18428,N_18095,N_18172);
and U18429 (N_18429,N_18045,N_18094);
nand U18430 (N_18430,N_18005,N_18230);
xnor U18431 (N_18431,N_18130,N_18177);
or U18432 (N_18432,N_18231,N_18183);
and U18433 (N_18433,N_18175,N_18128);
or U18434 (N_18434,N_18016,N_18060);
or U18435 (N_18435,N_18213,N_18040);
nor U18436 (N_18436,N_18109,N_18044);
or U18437 (N_18437,N_18049,N_18044);
or U18438 (N_18438,N_18010,N_18165);
xnor U18439 (N_18439,N_18191,N_18143);
xnor U18440 (N_18440,N_18139,N_18074);
nor U18441 (N_18441,N_18168,N_18143);
nand U18442 (N_18442,N_18142,N_18053);
nor U18443 (N_18443,N_18183,N_18035);
nand U18444 (N_18444,N_18064,N_18155);
or U18445 (N_18445,N_18198,N_18125);
xnor U18446 (N_18446,N_18051,N_18050);
nor U18447 (N_18447,N_18147,N_18022);
and U18448 (N_18448,N_18089,N_18094);
or U18449 (N_18449,N_18186,N_18241);
nand U18450 (N_18450,N_18035,N_18130);
nand U18451 (N_18451,N_18154,N_18006);
xor U18452 (N_18452,N_18232,N_18208);
xor U18453 (N_18453,N_18011,N_18161);
xnor U18454 (N_18454,N_18001,N_18220);
and U18455 (N_18455,N_18172,N_18061);
and U18456 (N_18456,N_18196,N_18054);
and U18457 (N_18457,N_18004,N_18224);
nand U18458 (N_18458,N_18027,N_18003);
or U18459 (N_18459,N_18234,N_18215);
or U18460 (N_18460,N_18247,N_18105);
xor U18461 (N_18461,N_18228,N_18215);
xor U18462 (N_18462,N_18220,N_18217);
xor U18463 (N_18463,N_18125,N_18056);
nand U18464 (N_18464,N_18033,N_18076);
and U18465 (N_18465,N_18189,N_18099);
nand U18466 (N_18466,N_18167,N_18074);
xnor U18467 (N_18467,N_18182,N_18131);
and U18468 (N_18468,N_18104,N_18071);
nor U18469 (N_18469,N_18234,N_18057);
or U18470 (N_18470,N_18247,N_18191);
and U18471 (N_18471,N_18040,N_18075);
xor U18472 (N_18472,N_18051,N_18011);
and U18473 (N_18473,N_18145,N_18196);
nor U18474 (N_18474,N_18000,N_18245);
nand U18475 (N_18475,N_18197,N_18219);
nand U18476 (N_18476,N_18006,N_18240);
nor U18477 (N_18477,N_18188,N_18178);
xor U18478 (N_18478,N_18104,N_18079);
or U18479 (N_18479,N_18032,N_18229);
and U18480 (N_18480,N_18006,N_18030);
nor U18481 (N_18481,N_18147,N_18173);
and U18482 (N_18482,N_18010,N_18106);
or U18483 (N_18483,N_18244,N_18207);
xor U18484 (N_18484,N_18190,N_18139);
nand U18485 (N_18485,N_18203,N_18053);
xnor U18486 (N_18486,N_18127,N_18087);
or U18487 (N_18487,N_18195,N_18219);
and U18488 (N_18488,N_18181,N_18224);
xnor U18489 (N_18489,N_18107,N_18131);
nor U18490 (N_18490,N_18117,N_18160);
nor U18491 (N_18491,N_18064,N_18119);
nand U18492 (N_18492,N_18058,N_18195);
or U18493 (N_18493,N_18209,N_18232);
nand U18494 (N_18494,N_18046,N_18227);
or U18495 (N_18495,N_18134,N_18103);
nor U18496 (N_18496,N_18127,N_18001);
or U18497 (N_18497,N_18141,N_18234);
or U18498 (N_18498,N_18228,N_18199);
and U18499 (N_18499,N_18215,N_18131);
xor U18500 (N_18500,N_18257,N_18396);
or U18501 (N_18501,N_18341,N_18302);
or U18502 (N_18502,N_18392,N_18481);
nand U18503 (N_18503,N_18362,N_18387);
and U18504 (N_18504,N_18305,N_18471);
nor U18505 (N_18505,N_18403,N_18343);
xor U18506 (N_18506,N_18426,N_18280);
nand U18507 (N_18507,N_18442,N_18256);
nand U18508 (N_18508,N_18319,N_18320);
or U18509 (N_18509,N_18317,N_18309);
nor U18510 (N_18510,N_18447,N_18480);
xnor U18511 (N_18511,N_18338,N_18298);
nand U18512 (N_18512,N_18488,N_18325);
nor U18513 (N_18513,N_18301,N_18406);
or U18514 (N_18514,N_18457,N_18268);
xnor U18515 (N_18515,N_18398,N_18335);
or U18516 (N_18516,N_18294,N_18443);
xor U18517 (N_18517,N_18253,N_18349);
xnor U18518 (N_18518,N_18415,N_18371);
nand U18519 (N_18519,N_18353,N_18437);
or U18520 (N_18520,N_18283,N_18438);
xor U18521 (N_18521,N_18448,N_18327);
or U18522 (N_18522,N_18342,N_18446);
and U18523 (N_18523,N_18279,N_18436);
nand U18524 (N_18524,N_18485,N_18432);
or U18525 (N_18525,N_18478,N_18411);
and U18526 (N_18526,N_18422,N_18258);
xnor U18527 (N_18527,N_18308,N_18408);
xor U18528 (N_18528,N_18358,N_18296);
nor U18529 (N_18529,N_18297,N_18329);
and U18530 (N_18530,N_18374,N_18321);
and U18531 (N_18531,N_18334,N_18272);
and U18532 (N_18532,N_18351,N_18454);
nand U18533 (N_18533,N_18379,N_18372);
or U18534 (N_18534,N_18375,N_18449);
and U18535 (N_18535,N_18440,N_18355);
xnor U18536 (N_18536,N_18496,N_18427);
nor U18537 (N_18537,N_18441,N_18340);
xnor U18538 (N_18538,N_18475,N_18269);
xor U18539 (N_18539,N_18332,N_18425);
xor U18540 (N_18540,N_18393,N_18328);
nor U18541 (N_18541,N_18458,N_18430);
nor U18542 (N_18542,N_18336,N_18473);
nor U18543 (N_18543,N_18312,N_18397);
nand U18544 (N_18544,N_18368,N_18263);
nand U18545 (N_18545,N_18439,N_18260);
and U18546 (N_18546,N_18276,N_18450);
or U18547 (N_18547,N_18416,N_18453);
nand U18548 (N_18548,N_18483,N_18337);
or U18549 (N_18549,N_18391,N_18405);
xnor U18550 (N_18550,N_18431,N_18360);
xnor U18551 (N_18551,N_18267,N_18377);
and U18552 (N_18552,N_18487,N_18350);
nand U18553 (N_18553,N_18367,N_18266);
xor U18554 (N_18554,N_18363,N_18359);
or U18555 (N_18555,N_18383,N_18467);
xnor U18556 (N_18556,N_18490,N_18404);
xor U18557 (N_18557,N_18402,N_18281);
nand U18558 (N_18558,N_18300,N_18264);
and U18559 (N_18559,N_18369,N_18289);
nand U18560 (N_18560,N_18292,N_18385);
or U18561 (N_18561,N_18347,N_18290);
xnor U18562 (N_18562,N_18262,N_18315);
and U18563 (N_18563,N_18477,N_18252);
or U18564 (N_18564,N_18421,N_18282);
nor U18565 (N_18565,N_18434,N_18493);
or U18566 (N_18566,N_18459,N_18464);
nand U18567 (N_18567,N_18474,N_18330);
xor U18568 (N_18568,N_18318,N_18412);
and U18569 (N_18569,N_18251,N_18400);
nand U18570 (N_18570,N_18380,N_18420);
nand U18571 (N_18571,N_18401,N_18452);
xor U18572 (N_18572,N_18484,N_18295);
or U18573 (N_18573,N_18378,N_18313);
or U18574 (N_18574,N_18344,N_18451);
nand U18575 (N_18575,N_18288,N_18410);
or U18576 (N_18576,N_18462,N_18326);
and U18577 (N_18577,N_18435,N_18482);
or U18578 (N_18578,N_18407,N_18417);
xor U18579 (N_18579,N_18352,N_18495);
xor U18580 (N_18580,N_18419,N_18331);
or U18581 (N_18581,N_18428,N_18498);
nand U18582 (N_18582,N_18445,N_18348);
xor U18583 (N_18583,N_18271,N_18361);
nor U18584 (N_18584,N_18255,N_18499);
nand U18585 (N_18585,N_18366,N_18429);
and U18586 (N_18586,N_18414,N_18287);
nand U18587 (N_18587,N_18463,N_18382);
nor U18588 (N_18588,N_18461,N_18333);
nor U18589 (N_18589,N_18376,N_18497);
and U18590 (N_18590,N_18386,N_18423);
or U18591 (N_18591,N_18413,N_18479);
nand U18592 (N_18592,N_18261,N_18444);
nand U18593 (N_18593,N_18456,N_18395);
nand U18594 (N_18594,N_18291,N_18323);
or U18595 (N_18595,N_18311,N_18310);
nor U18596 (N_18596,N_18476,N_18286);
nand U18597 (N_18597,N_18373,N_18494);
nor U18598 (N_18598,N_18466,N_18424);
nor U18599 (N_18599,N_18486,N_18306);
nor U18600 (N_18600,N_18433,N_18270);
nand U18601 (N_18601,N_18274,N_18314);
nand U18602 (N_18602,N_18322,N_18307);
and U18603 (N_18603,N_18250,N_18339);
or U18604 (N_18604,N_18324,N_18278);
and U18605 (N_18605,N_18356,N_18389);
or U18606 (N_18606,N_18394,N_18465);
nor U18607 (N_18607,N_18345,N_18460);
nand U18608 (N_18608,N_18455,N_18381);
xnor U18609 (N_18609,N_18409,N_18418);
nor U18610 (N_18610,N_18265,N_18388);
and U18611 (N_18611,N_18469,N_18273);
nor U18612 (N_18612,N_18390,N_18293);
and U18613 (N_18613,N_18304,N_18259);
or U18614 (N_18614,N_18346,N_18468);
and U18615 (N_18615,N_18303,N_18285);
or U18616 (N_18616,N_18492,N_18491);
or U18617 (N_18617,N_18399,N_18472);
or U18618 (N_18618,N_18384,N_18284);
xnor U18619 (N_18619,N_18364,N_18354);
nand U18620 (N_18620,N_18254,N_18365);
nand U18621 (N_18621,N_18299,N_18357);
and U18622 (N_18622,N_18277,N_18275);
or U18623 (N_18623,N_18316,N_18470);
or U18624 (N_18624,N_18370,N_18489);
nor U18625 (N_18625,N_18419,N_18307);
nand U18626 (N_18626,N_18368,N_18480);
nor U18627 (N_18627,N_18305,N_18298);
or U18628 (N_18628,N_18256,N_18250);
xnor U18629 (N_18629,N_18361,N_18419);
or U18630 (N_18630,N_18476,N_18336);
or U18631 (N_18631,N_18405,N_18450);
xnor U18632 (N_18632,N_18305,N_18412);
nand U18633 (N_18633,N_18390,N_18494);
and U18634 (N_18634,N_18272,N_18322);
xor U18635 (N_18635,N_18334,N_18434);
xnor U18636 (N_18636,N_18384,N_18455);
nor U18637 (N_18637,N_18311,N_18276);
nand U18638 (N_18638,N_18333,N_18473);
or U18639 (N_18639,N_18384,N_18469);
nand U18640 (N_18640,N_18285,N_18393);
nand U18641 (N_18641,N_18378,N_18268);
nand U18642 (N_18642,N_18321,N_18365);
nand U18643 (N_18643,N_18336,N_18475);
or U18644 (N_18644,N_18428,N_18350);
and U18645 (N_18645,N_18432,N_18437);
and U18646 (N_18646,N_18469,N_18293);
nand U18647 (N_18647,N_18293,N_18497);
or U18648 (N_18648,N_18255,N_18423);
nor U18649 (N_18649,N_18427,N_18349);
or U18650 (N_18650,N_18351,N_18396);
nor U18651 (N_18651,N_18327,N_18306);
nor U18652 (N_18652,N_18429,N_18373);
nor U18653 (N_18653,N_18490,N_18305);
and U18654 (N_18654,N_18290,N_18486);
xnor U18655 (N_18655,N_18313,N_18262);
xnor U18656 (N_18656,N_18335,N_18432);
nor U18657 (N_18657,N_18320,N_18402);
or U18658 (N_18658,N_18426,N_18379);
and U18659 (N_18659,N_18255,N_18286);
xor U18660 (N_18660,N_18477,N_18427);
or U18661 (N_18661,N_18409,N_18361);
nor U18662 (N_18662,N_18294,N_18388);
xor U18663 (N_18663,N_18463,N_18388);
and U18664 (N_18664,N_18317,N_18331);
xor U18665 (N_18665,N_18478,N_18364);
xor U18666 (N_18666,N_18326,N_18339);
xor U18667 (N_18667,N_18305,N_18429);
nor U18668 (N_18668,N_18323,N_18478);
nand U18669 (N_18669,N_18320,N_18418);
nor U18670 (N_18670,N_18445,N_18481);
nand U18671 (N_18671,N_18425,N_18435);
or U18672 (N_18672,N_18357,N_18393);
and U18673 (N_18673,N_18404,N_18401);
nand U18674 (N_18674,N_18304,N_18379);
xor U18675 (N_18675,N_18279,N_18376);
and U18676 (N_18676,N_18357,N_18339);
and U18677 (N_18677,N_18403,N_18481);
xnor U18678 (N_18678,N_18261,N_18387);
and U18679 (N_18679,N_18449,N_18459);
and U18680 (N_18680,N_18460,N_18315);
nand U18681 (N_18681,N_18332,N_18256);
or U18682 (N_18682,N_18396,N_18465);
nor U18683 (N_18683,N_18470,N_18326);
xnor U18684 (N_18684,N_18284,N_18452);
nand U18685 (N_18685,N_18322,N_18251);
and U18686 (N_18686,N_18336,N_18331);
and U18687 (N_18687,N_18427,N_18369);
xor U18688 (N_18688,N_18272,N_18260);
xnor U18689 (N_18689,N_18332,N_18418);
or U18690 (N_18690,N_18460,N_18472);
nand U18691 (N_18691,N_18495,N_18325);
xor U18692 (N_18692,N_18464,N_18264);
xnor U18693 (N_18693,N_18305,N_18393);
nor U18694 (N_18694,N_18368,N_18304);
or U18695 (N_18695,N_18318,N_18383);
nor U18696 (N_18696,N_18373,N_18376);
nand U18697 (N_18697,N_18476,N_18317);
nand U18698 (N_18698,N_18284,N_18445);
or U18699 (N_18699,N_18370,N_18309);
and U18700 (N_18700,N_18314,N_18309);
or U18701 (N_18701,N_18401,N_18324);
nor U18702 (N_18702,N_18497,N_18257);
xnor U18703 (N_18703,N_18454,N_18262);
or U18704 (N_18704,N_18298,N_18443);
or U18705 (N_18705,N_18330,N_18406);
nand U18706 (N_18706,N_18254,N_18256);
and U18707 (N_18707,N_18412,N_18319);
nor U18708 (N_18708,N_18470,N_18466);
xor U18709 (N_18709,N_18465,N_18386);
xnor U18710 (N_18710,N_18415,N_18482);
nor U18711 (N_18711,N_18286,N_18402);
nand U18712 (N_18712,N_18466,N_18446);
xor U18713 (N_18713,N_18280,N_18406);
nor U18714 (N_18714,N_18364,N_18468);
and U18715 (N_18715,N_18370,N_18355);
or U18716 (N_18716,N_18325,N_18478);
xor U18717 (N_18717,N_18445,N_18460);
or U18718 (N_18718,N_18398,N_18425);
nor U18719 (N_18719,N_18410,N_18433);
or U18720 (N_18720,N_18489,N_18421);
xnor U18721 (N_18721,N_18373,N_18379);
nor U18722 (N_18722,N_18439,N_18276);
xnor U18723 (N_18723,N_18364,N_18342);
nand U18724 (N_18724,N_18393,N_18497);
nor U18725 (N_18725,N_18493,N_18483);
xor U18726 (N_18726,N_18491,N_18493);
xor U18727 (N_18727,N_18412,N_18276);
nor U18728 (N_18728,N_18442,N_18395);
nand U18729 (N_18729,N_18279,N_18358);
and U18730 (N_18730,N_18266,N_18308);
nand U18731 (N_18731,N_18395,N_18308);
nor U18732 (N_18732,N_18439,N_18358);
nor U18733 (N_18733,N_18442,N_18374);
nand U18734 (N_18734,N_18327,N_18284);
or U18735 (N_18735,N_18401,N_18306);
nand U18736 (N_18736,N_18360,N_18303);
xnor U18737 (N_18737,N_18415,N_18313);
xor U18738 (N_18738,N_18264,N_18447);
or U18739 (N_18739,N_18323,N_18263);
nor U18740 (N_18740,N_18405,N_18272);
nor U18741 (N_18741,N_18319,N_18257);
nor U18742 (N_18742,N_18368,N_18334);
nor U18743 (N_18743,N_18254,N_18472);
xor U18744 (N_18744,N_18444,N_18466);
and U18745 (N_18745,N_18466,N_18402);
xor U18746 (N_18746,N_18333,N_18359);
or U18747 (N_18747,N_18326,N_18374);
or U18748 (N_18748,N_18325,N_18384);
and U18749 (N_18749,N_18409,N_18322);
or U18750 (N_18750,N_18676,N_18507);
nor U18751 (N_18751,N_18678,N_18660);
xor U18752 (N_18752,N_18540,N_18627);
nor U18753 (N_18753,N_18656,N_18648);
nor U18754 (N_18754,N_18591,N_18748);
or U18755 (N_18755,N_18621,N_18577);
or U18756 (N_18756,N_18624,N_18585);
and U18757 (N_18757,N_18616,N_18604);
nor U18758 (N_18758,N_18610,N_18592);
or U18759 (N_18759,N_18552,N_18744);
xor U18760 (N_18760,N_18683,N_18694);
nor U18761 (N_18761,N_18566,N_18679);
xor U18762 (N_18762,N_18563,N_18546);
xnor U18763 (N_18763,N_18581,N_18729);
nand U18764 (N_18764,N_18518,N_18682);
or U18765 (N_18765,N_18722,N_18612);
or U18766 (N_18766,N_18614,N_18700);
and U18767 (N_18767,N_18559,N_18503);
and U18768 (N_18768,N_18630,N_18725);
nand U18769 (N_18769,N_18698,N_18705);
or U18770 (N_18770,N_18579,N_18655);
nor U18771 (N_18771,N_18590,N_18562);
xnor U18772 (N_18772,N_18586,N_18661);
nand U18773 (N_18773,N_18537,N_18525);
nand U18774 (N_18774,N_18513,N_18512);
nor U18775 (N_18775,N_18634,N_18565);
and U18776 (N_18776,N_18571,N_18524);
nor U18777 (N_18777,N_18506,N_18597);
xnor U18778 (N_18778,N_18721,N_18576);
nor U18779 (N_18779,N_18669,N_18693);
nor U18780 (N_18780,N_18690,N_18663);
or U18781 (N_18781,N_18681,N_18712);
or U18782 (N_18782,N_18548,N_18608);
and U18783 (N_18783,N_18715,N_18555);
nand U18784 (N_18784,N_18737,N_18732);
and U18785 (N_18785,N_18620,N_18743);
or U18786 (N_18786,N_18549,N_18501);
nand U18787 (N_18787,N_18739,N_18606);
nor U18788 (N_18788,N_18583,N_18684);
or U18789 (N_18789,N_18502,N_18557);
nor U18790 (N_18790,N_18633,N_18587);
or U18791 (N_18791,N_18645,N_18746);
or U18792 (N_18792,N_18658,N_18701);
nand U18793 (N_18793,N_18726,N_18711);
xor U18794 (N_18794,N_18596,N_18574);
or U18795 (N_18795,N_18723,N_18653);
nand U18796 (N_18796,N_18509,N_18717);
nand U18797 (N_18797,N_18742,N_18514);
or U18798 (N_18798,N_18593,N_18625);
nor U18799 (N_18799,N_18649,N_18622);
xor U18800 (N_18800,N_18735,N_18692);
or U18801 (N_18801,N_18522,N_18554);
or U18802 (N_18802,N_18561,N_18706);
or U18803 (N_18803,N_18703,N_18733);
nand U18804 (N_18804,N_18745,N_18582);
nand U18805 (N_18805,N_18638,N_18594);
xnor U18806 (N_18806,N_18618,N_18508);
nor U18807 (N_18807,N_18657,N_18516);
nor U18808 (N_18808,N_18728,N_18567);
xor U18809 (N_18809,N_18600,N_18564);
or U18810 (N_18810,N_18505,N_18504);
and U18811 (N_18811,N_18718,N_18652);
and U18812 (N_18812,N_18575,N_18521);
and U18813 (N_18813,N_18623,N_18500);
nand U18814 (N_18814,N_18714,N_18536);
nand U18815 (N_18815,N_18530,N_18719);
and U18816 (N_18816,N_18531,N_18670);
or U18817 (N_18817,N_18541,N_18523);
nor U18818 (N_18818,N_18617,N_18568);
and U18819 (N_18819,N_18687,N_18632);
xor U18820 (N_18820,N_18510,N_18560);
or U18821 (N_18821,N_18538,N_18511);
nand U18822 (N_18822,N_18727,N_18539);
or U18823 (N_18823,N_18527,N_18654);
nand U18824 (N_18824,N_18547,N_18664);
xor U18825 (N_18825,N_18680,N_18553);
and U18826 (N_18826,N_18686,N_18556);
and U18827 (N_18827,N_18674,N_18716);
xor U18828 (N_18828,N_18550,N_18607);
nand U18829 (N_18829,N_18668,N_18598);
and U18830 (N_18830,N_18710,N_18599);
nand U18831 (N_18831,N_18595,N_18666);
and U18832 (N_18832,N_18572,N_18529);
nand U18833 (N_18833,N_18584,N_18659);
nand U18834 (N_18834,N_18619,N_18672);
nand U18835 (N_18835,N_18738,N_18615);
nor U18836 (N_18836,N_18628,N_18677);
nand U18837 (N_18837,N_18626,N_18534);
nor U18838 (N_18838,N_18730,N_18588);
and U18839 (N_18839,N_18580,N_18709);
nor U18840 (N_18840,N_18697,N_18713);
and U18841 (N_18841,N_18665,N_18639);
xnor U18842 (N_18842,N_18558,N_18647);
nand U18843 (N_18843,N_18724,N_18695);
nand U18844 (N_18844,N_18611,N_18631);
nand U18845 (N_18845,N_18667,N_18573);
xnor U18846 (N_18846,N_18688,N_18543);
nand U18847 (N_18847,N_18702,N_18691);
nor U18848 (N_18848,N_18602,N_18731);
nor U18849 (N_18849,N_18551,N_18704);
nor U18850 (N_18850,N_18736,N_18570);
xnor U18851 (N_18851,N_18603,N_18734);
nor U18852 (N_18852,N_18640,N_18662);
nand U18853 (N_18853,N_18636,N_18578);
or U18854 (N_18854,N_18635,N_18685);
nand U18855 (N_18855,N_18696,N_18533);
nand U18856 (N_18856,N_18740,N_18747);
nor U18857 (N_18857,N_18720,N_18699);
or U18858 (N_18858,N_18605,N_18644);
nand U18859 (N_18859,N_18526,N_18517);
or U18860 (N_18860,N_18673,N_18749);
nand U18861 (N_18861,N_18589,N_18569);
nor U18862 (N_18862,N_18532,N_18675);
nor U18863 (N_18863,N_18613,N_18535);
nor U18864 (N_18864,N_18544,N_18689);
xnor U18865 (N_18865,N_18609,N_18528);
nand U18866 (N_18866,N_18708,N_18671);
nor U18867 (N_18867,N_18520,N_18651);
xnor U18868 (N_18868,N_18637,N_18519);
nor U18869 (N_18869,N_18629,N_18741);
nand U18870 (N_18870,N_18515,N_18707);
nand U18871 (N_18871,N_18642,N_18542);
and U18872 (N_18872,N_18650,N_18601);
and U18873 (N_18873,N_18643,N_18641);
and U18874 (N_18874,N_18545,N_18646);
or U18875 (N_18875,N_18705,N_18701);
nor U18876 (N_18876,N_18518,N_18678);
or U18877 (N_18877,N_18644,N_18657);
and U18878 (N_18878,N_18678,N_18583);
xor U18879 (N_18879,N_18512,N_18679);
nand U18880 (N_18880,N_18681,N_18582);
xnor U18881 (N_18881,N_18668,N_18747);
and U18882 (N_18882,N_18628,N_18528);
and U18883 (N_18883,N_18619,N_18659);
or U18884 (N_18884,N_18600,N_18677);
xnor U18885 (N_18885,N_18600,N_18674);
or U18886 (N_18886,N_18724,N_18660);
xnor U18887 (N_18887,N_18640,N_18611);
xnor U18888 (N_18888,N_18721,N_18507);
or U18889 (N_18889,N_18659,N_18571);
or U18890 (N_18890,N_18564,N_18502);
xor U18891 (N_18891,N_18682,N_18623);
xor U18892 (N_18892,N_18560,N_18646);
or U18893 (N_18893,N_18714,N_18658);
and U18894 (N_18894,N_18552,N_18547);
and U18895 (N_18895,N_18626,N_18740);
and U18896 (N_18896,N_18686,N_18693);
or U18897 (N_18897,N_18706,N_18741);
nor U18898 (N_18898,N_18637,N_18641);
nand U18899 (N_18899,N_18639,N_18627);
or U18900 (N_18900,N_18664,N_18670);
nand U18901 (N_18901,N_18538,N_18745);
nand U18902 (N_18902,N_18640,N_18602);
nand U18903 (N_18903,N_18698,N_18677);
nand U18904 (N_18904,N_18609,N_18666);
and U18905 (N_18905,N_18512,N_18609);
and U18906 (N_18906,N_18651,N_18552);
xor U18907 (N_18907,N_18595,N_18571);
nor U18908 (N_18908,N_18553,N_18552);
xnor U18909 (N_18909,N_18557,N_18735);
or U18910 (N_18910,N_18556,N_18670);
or U18911 (N_18911,N_18685,N_18648);
nand U18912 (N_18912,N_18662,N_18651);
nor U18913 (N_18913,N_18721,N_18567);
or U18914 (N_18914,N_18727,N_18748);
and U18915 (N_18915,N_18561,N_18666);
xnor U18916 (N_18916,N_18515,N_18547);
nand U18917 (N_18917,N_18697,N_18622);
or U18918 (N_18918,N_18532,N_18645);
nand U18919 (N_18919,N_18506,N_18707);
or U18920 (N_18920,N_18733,N_18511);
nor U18921 (N_18921,N_18537,N_18692);
nor U18922 (N_18922,N_18550,N_18738);
xnor U18923 (N_18923,N_18681,N_18558);
nand U18924 (N_18924,N_18516,N_18582);
xor U18925 (N_18925,N_18715,N_18671);
nor U18926 (N_18926,N_18708,N_18610);
nand U18927 (N_18927,N_18578,N_18567);
and U18928 (N_18928,N_18686,N_18666);
or U18929 (N_18929,N_18584,N_18704);
xor U18930 (N_18930,N_18672,N_18564);
nand U18931 (N_18931,N_18626,N_18716);
or U18932 (N_18932,N_18599,N_18677);
and U18933 (N_18933,N_18684,N_18687);
and U18934 (N_18934,N_18542,N_18524);
nand U18935 (N_18935,N_18607,N_18656);
nand U18936 (N_18936,N_18653,N_18738);
nand U18937 (N_18937,N_18561,N_18585);
xor U18938 (N_18938,N_18561,N_18646);
or U18939 (N_18939,N_18521,N_18693);
xnor U18940 (N_18940,N_18539,N_18655);
nand U18941 (N_18941,N_18597,N_18538);
and U18942 (N_18942,N_18621,N_18691);
xnor U18943 (N_18943,N_18746,N_18730);
or U18944 (N_18944,N_18560,N_18636);
nor U18945 (N_18945,N_18648,N_18531);
nand U18946 (N_18946,N_18713,N_18749);
nand U18947 (N_18947,N_18566,N_18677);
nor U18948 (N_18948,N_18583,N_18633);
xor U18949 (N_18949,N_18550,N_18710);
xor U18950 (N_18950,N_18708,N_18736);
nand U18951 (N_18951,N_18591,N_18512);
nor U18952 (N_18952,N_18524,N_18637);
nor U18953 (N_18953,N_18746,N_18650);
nand U18954 (N_18954,N_18698,N_18530);
nand U18955 (N_18955,N_18667,N_18506);
nor U18956 (N_18956,N_18610,N_18512);
or U18957 (N_18957,N_18501,N_18608);
nor U18958 (N_18958,N_18618,N_18507);
nor U18959 (N_18959,N_18698,N_18657);
nand U18960 (N_18960,N_18521,N_18656);
and U18961 (N_18961,N_18551,N_18745);
and U18962 (N_18962,N_18704,N_18711);
nand U18963 (N_18963,N_18577,N_18729);
and U18964 (N_18964,N_18749,N_18542);
and U18965 (N_18965,N_18572,N_18643);
or U18966 (N_18966,N_18614,N_18539);
xor U18967 (N_18967,N_18516,N_18709);
and U18968 (N_18968,N_18538,N_18714);
and U18969 (N_18969,N_18663,N_18725);
and U18970 (N_18970,N_18748,N_18509);
nand U18971 (N_18971,N_18686,N_18657);
xnor U18972 (N_18972,N_18547,N_18573);
nand U18973 (N_18973,N_18730,N_18512);
xnor U18974 (N_18974,N_18690,N_18711);
nor U18975 (N_18975,N_18749,N_18503);
or U18976 (N_18976,N_18619,N_18502);
or U18977 (N_18977,N_18503,N_18500);
or U18978 (N_18978,N_18693,N_18581);
and U18979 (N_18979,N_18652,N_18675);
or U18980 (N_18980,N_18501,N_18528);
or U18981 (N_18981,N_18506,N_18728);
nor U18982 (N_18982,N_18567,N_18680);
nor U18983 (N_18983,N_18565,N_18711);
or U18984 (N_18984,N_18540,N_18725);
or U18985 (N_18985,N_18689,N_18719);
nand U18986 (N_18986,N_18674,N_18588);
nand U18987 (N_18987,N_18747,N_18681);
xnor U18988 (N_18988,N_18618,N_18665);
xnor U18989 (N_18989,N_18610,N_18624);
nor U18990 (N_18990,N_18673,N_18543);
xor U18991 (N_18991,N_18705,N_18614);
or U18992 (N_18992,N_18650,N_18556);
and U18993 (N_18993,N_18586,N_18571);
nand U18994 (N_18994,N_18549,N_18618);
xor U18995 (N_18995,N_18631,N_18713);
or U18996 (N_18996,N_18602,N_18674);
nor U18997 (N_18997,N_18582,N_18688);
nand U18998 (N_18998,N_18517,N_18658);
and U18999 (N_18999,N_18526,N_18569);
nand U19000 (N_19000,N_18848,N_18863);
nand U19001 (N_19001,N_18867,N_18859);
nor U19002 (N_19002,N_18872,N_18801);
nor U19003 (N_19003,N_18906,N_18942);
or U19004 (N_19004,N_18963,N_18890);
nor U19005 (N_19005,N_18881,N_18773);
nand U19006 (N_19006,N_18896,N_18797);
nor U19007 (N_19007,N_18817,N_18922);
xnor U19008 (N_19008,N_18958,N_18913);
and U19009 (N_19009,N_18815,N_18956);
xor U19010 (N_19010,N_18768,N_18975);
nand U19011 (N_19011,N_18973,N_18766);
nor U19012 (N_19012,N_18826,N_18901);
nor U19013 (N_19013,N_18914,N_18789);
or U19014 (N_19014,N_18771,N_18823);
and U19015 (N_19015,N_18845,N_18920);
nor U19016 (N_19016,N_18853,N_18844);
xnor U19017 (N_19017,N_18992,N_18871);
or U19018 (N_19018,N_18761,N_18915);
xnor U19019 (N_19019,N_18880,N_18821);
and U19020 (N_19020,N_18990,N_18791);
or U19021 (N_19021,N_18833,N_18757);
nor U19022 (N_19022,N_18892,N_18957);
xor U19023 (N_19023,N_18910,N_18976);
or U19024 (N_19024,N_18861,N_18798);
xor U19025 (N_19025,N_18781,N_18796);
or U19026 (N_19026,N_18986,N_18782);
or U19027 (N_19027,N_18807,N_18926);
and U19028 (N_19028,N_18825,N_18783);
xor U19029 (N_19029,N_18932,N_18813);
nor U19030 (N_19030,N_18769,N_18944);
xor U19031 (N_19031,N_18857,N_18884);
xor U19032 (N_19032,N_18750,N_18804);
and U19033 (N_19033,N_18964,N_18893);
or U19034 (N_19034,N_18832,N_18984);
nand U19035 (N_19035,N_18888,N_18852);
xor U19036 (N_19036,N_18938,N_18868);
and U19037 (N_19037,N_18777,N_18754);
xnor U19038 (N_19038,N_18971,N_18997);
xor U19039 (N_19039,N_18836,N_18991);
or U19040 (N_19040,N_18847,N_18755);
nand U19041 (N_19041,N_18865,N_18827);
and U19042 (N_19042,N_18946,N_18787);
nor U19043 (N_19043,N_18940,N_18962);
xor U19044 (N_19044,N_18967,N_18993);
nor U19045 (N_19045,N_18972,N_18998);
nand U19046 (N_19046,N_18764,N_18904);
xnor U19047 (N_19047,N_18918,N_18824);
nand U19048 (N_19048,N_18995,N_18927);
nor U19049 (N_19049,N_18864,N_18941);
or U19050 (N_19050,N_18794,N_18921);
nand U19051 (N_19051,N_18855,N_18919);
xor U19052 (N_19052,N_18762,N_18961);
xor U19053 (N_19053,N_18834,N_18876);
and U19054 (N_19054,N_18923,N_18908);
or U19055 (N_19055,N_18811,N_18830);
nand U19056 (N_19056,N_18903,N_18945);
and U19057 (N_19057,N_18784,N_18900);
or U19058 (N_19058,N_18806,N_18959);
and U19059 (N_19059,N_18886,N_18862);
xnor U19060 (N_19060,N_18935,N_18786);
xor U19061 (N_19061,N_18842,N_18917);
and U19062 (N_19062,N_18816,N_18803);
or U19063 (N_19063,N_18778,N_18874);
xnor U19064 (N_19064,N_18854,N_18887);
nand U19065 (N_19065,N_18965,N_18882);
nor U19066 (N_19066,N_18828,N_18899);
or U19067 (N_19067,N_18799,N_18841);
and U19068 (N_19068,N_18902,N_18974);
xor U19069 (N_19069,N_18759,N_18858);
or U19070 (N_19070,N_18795,N_18793);
and U19071 (N_19071,N_18911,N_18883);
or U19072 (N_19072,N_18785,N_18994);
nand U19073 (N_19073,N_18969,N_18912);
and U19074 (N_19074,N_18928,N_18982);
nand U19075 (N_19075,N_18822,N_18758);
xor U19076 (N_19076,N_18837,N_18977);
nand U19077 (N_19077,N_18989,N_18838);
xor U19078 (N_19078,N_18996,N_18760);
xnor U19079 (N_19079,N_18951,N_18943);
nor U19080 (N_19080,N_18891,N_18790);
nand U19081 (N_19081,N_18851,N_18925);
or U19082 (N_19082,N_18763,N_18894);
and U19083 (N_19083,N_18788,N_18770);
nand U19084 (N_19084,N_18936,N_18756);
xor U19085 (N_19085,N_18879,N_18751);
nor U19086 (N_19086,N_18978,N_18999);
nand U19087 (N_19087,N_18981,N_18775);
xor U19088 (N_19088,N_18980,N_18869);
and U19089 (N_19089,N_18772,N_18929);
xor U19090 (N_19090,N_18860,N_18819);
or U19091 (N_19091,N_18934,N_18952);
or U19092 (N_19092,N_18765,N_18970);
nor U19093 (N_19093,N_18898,N_18953);
or U19094 (N_19094,N_18889,N_18829);
xnor U19095 (N_19095,N_18753,N_18987);
xnor U19096 (N_19096,N_18843,N_18839);
nand U19097 (N_19097,N_18774,N_18820);
or U19098 (N_19098,N_18950,N_18780);
xnor U19099 (N_19099,N_18776,N_18802);
nand U19100 (N_19100,N_18933,N_18968);
nor U19101 (N_19101,N_18810,N_18907);
xnor U19102 (N_19102,N_18916,N_18948);
and U19103 (N_19103,N_18870,N_18856);
nand U19104 (N_19104,N_18930,N_18931);
nand U19105 (N_19105,N_18960,N_18979);
and U19106 (N_19106,N_18947,N_18983);
and U19107 (N_19107,N_18966,N_18866);
and U19108 (N_19108,N_18835,N_18805);
nor U19109 (N_19109,N_18818,N_18767);
and U19110 (N_19110,N_18814,N_18812);
and U19111 (N_19111,N_18846,N_18800);
and U19112 (N_19112,N_18905,N_18937);
and U19113 (N_19113,N_18955,N_18924);
xor U19114 (N_19114,N_18885,N_18873);
nand U19115 (N_19115,N_18831,N_18752);
nor U19116 (N_19116,N_18897,N_18939);
xor U19117 (N_19117,N_18949,N_18877);
and U19118 (N_19118,N_18875,N_18954);
or U19119 (N_19119,N_18895,N_18792);
and U19120 (N_19120,N_18878,N_18850);
xor U19121 (N_19121,N_18779,N_18808);
or U19122 (N_19122,N_18840,N_18985);
nor U19123 (N_19123,N_18988,N_18809);
or U19124 (N_19124,N_18849,N_18909);
nand U19125 (N_19125,N_18882,N_18964);
and U19126 (N_19126,N_18776,N_18912);
xor U19127 (N_19127,N_18974,N_18946);
xnor U19128 (N_19128,N_18915,N_18835);
xnor U19129 (N_19129,N_18846,N_18827);
and U19130 (N_19130,N_18959,N_18821);
nand U19131 (N_19131,N_18814,N_18850);
and U19132 (N_19132,N_18969,N_18999);
and U19133 (N_19133,N_18871,N_18890);
nor U19134 (N_19134,N_18937,N_18990);
or U19135 (N_19135,N_18833,N_18916);
or U19136 (N_19136,N_18861,N_18996);
nand U19137 (N_19137,N_18919,N_18801);
or U19138 (N_19138,N_18971,N_18862);
or U19139 (N_19139,N_18878,N_18903);
and U19140 (N_19140,N_18827,N_18940);
xnor U19141 (N_19141,N_18837,N_18766);
or U19142 (N_19142,N_18817,N_18995);
xor U19143 (N_19143,N_18991,N_18751);
nor U19144 (N_19144,N_18995,N_18979);
nand U19145 (N_19145,N_18936,N_18836);
and U19146 (N_19146,N_18975,N_18762);
nor U19147 (N_19147,N_18846,N_18914);
nor U19148 (N_19148,N_18844,N_18958);
nand U19149 (N_19149,N_18750,N_18904);
nand U19150 (N_19150,N_18866,N_18875);
and U19151 (N_19151,N_18806,N_18967);
and U19152 (N_19152,N_18900,N_18813);
and U19153 (N_19153,N_18851,N_18858);
and U19154 (N_19154,N_18828,N_18877);
xnor U19155 (N_19155,N_18775,N_18852);
and U19156 (N_19156,N_18855,N_18823);
xnor U19157 (N_19157,N_18796,N_18883);
or U19158 (N_19158,N_18830,N_18900);
nand U19159 (N_19159,N_18829,N_18899);
nor U19160 (N_19160,N_18999,N_18982);
nand U19161 (N_19161,N_18976,N_18944);
and U19162 (N_19162,N_18981,N_18905);
and U19163 (N_19163,N_18772,N_18937);
or U19164 (N_19164,N_18973,N_18753);
nor U19165 (N_19165,N_18835,N_18783);
nand U19166 (N_19166,N_18877,N_18986);
nor U19167 (N_19167,N_18912,N_18867);
and U19168 (N_19168,N_18801,N_18932);
xor U19169 (N_19169,N_18807,N_18761);
and U19170 (N_19170,N_18809,N_18906);
nand U19171 (N_19171,N_18851,N_18975);
xor U19172 (N_19172,N_18809,N_18839);
and U19173 (N_19173,N_18879,N_18791);
nand U19174 (N_19174,N_18849,N_18987);
or U19175 (N_19175,N_18760,N_18978);
nand U19176 (N_19176,N_18761,N_18884);
or U19177 (N_19177,N_18787,N_18776);
or U19178 (N_19178,N_18975,N_18794);
nand U19179 (N_19179,N_18750,N_18761);
or U19180 (N_19180,N_18875,N_18885);
nand U19181 (N_19181,N_18780,N_18967);
and U19182 (N_19182,N_18789,N_18880);
and U19183 (N_19183,N_18968,N_18835);
nor U19184 (N_19184,N_18980,N_18981);
or U19185 (N_19185,N_18816,N_18837);
or U19186 (N_19186,N_18982,N_18856);
and U19187 (N_19187,N_18817,N_18980);
xor U19188 (N_19188,N_18975,N_18869);
nand U19189 (N_19189,N_18960,N_18951);
and U19190 (N_19190,N_18779,N_18971);
or U19191 (N_19191,N_18787,N_18866);
nor U19192 (N_19192,N_18998,N_18808);
or U19193 (N_19193,N_18915,N_18858);
nor U19194 (N_19194,N_18926,N_18880);
nor U19195 (N_19195,N_18796,N_18874);
nor U19196 (N_19196,N_18886,N_18900);
or U19197 (N_19197,N_18854,N_18777);
xnor U19198 (N_19198,N_18776,N_18773);
xor U19199 (N_19199,N_18942,N_18868);
xnor U19200 (N_19200,N_18994,N_18894);
or U19201 (N_19201,N_18926,N_18891);
nand U19202 (N_19202,N_18780,N_18984);
nand U19203 (N_19203,N_18992,N_18899);
and U19204 (N_19204,N_18895,N_18980);
or U19205 (N_19205,N_18790,N_18840);
xnor U19206 (N_19206,N_18852,N_18815);
nand U19207 (N_19207,N_18803,N_18887);
xnor U19208 (N_19208,N_18837,N_18770);
or U19209 (N_19209,N_18910,N_18972);
nand U19210 (N_19210,N_18757,N_18976);
nand U19211 (N_19211,N_18823,N_18903);
nor U19212 (N_19212,N_18819,N_18944);
nor U19213 (N_19213,N_18981,N_18876);
and U19214 (N_19214,N_18946,N_18936);
and U19215 (N_19215,N_18788,N_18976);
and U19216 (N_19216,N_18804,N_18888);
xnor U19217 (N_19217,N_18996,N_18982);
nand U19218 (N_19218,N_18850,N_18972);
and U19219 (N_19219,N_18798,N_18877);
nor U19220 (N_19220,N_18777,N_18779);
xor U19221 (N_19221,N_18763,N_18893);
nor U19222 (N_19222,N_18808,N_18811);
nand U19223 (N_19223,N_18958,N_18761);
nor U19224 (N_19224,N_18750,N_18995);
nor U19225 (N_19225,N_18848,N_18861);
or U19226 (N_19226,N_18773,N_18995);
nand U19227 (N_19227,N_18874,N_18936);
nor U19228 (N_19228,N_18843,N_18813);
and U19229 (N_19229,N_18916,N_18855);
nand U19230 (N_19230,N_18788,N_18894);
nand U19231 (N_19231,N_18794,N_18959);
nand U19232 (N_19232,N_18822,N_18782);
xnor U19233 (N_19233,N_18947,N_18948);
xnor U19234 (N_19234,N_18827,N_18852);
or U19235 (N_19235,N_18842,N_18968);
nand U19236 (N_19236,N_18925,N_18862);
xor U19237 (N_19237,N_18917,N_18810);
and U19238 (N_19238,N_18928,N_18879);
nand U19239 (N_19239,N_18807,N_18784);
xor U19240 (N_19240,N_18846,N_18927);
xnor U19241 (N_19241,N_18919,N_18782);
or U19242 (N_19242,N_18878,N_18914);
xnor U19243 (N_19243,N_18759,N_18980);
or U19244 (N_19244,N_18989,N_18860);
or U19245 (N_19245,N_18860,N_18883);
xor U19246 (N_19246,N_18844,N_18814);
or U19247 (N_19247,N_18874,N_18753);
nor U19248 (N_19248,N_18924,N_18788);
and U19249 (N_19249,N_18850,N_18967);
nor U19250 (N_19250,N_19079,N_19112);
nand U19251 (N_19251,N_19055,N_19046);
nand U19252 (N_19252,N_19192,N_19016);
and U19253 (N_19253,N_19098,N_19158);
and U19254 (N_19254,N_19196,N_19062);
and U19255 (N_19255,N_19164,N_19003);
or U19256 (N_19256,N_19049,N_19221);
nor U19257 (N_19257,N_19103,N_19228);
or U19258 (N_19258,N_19211,N_19172);
and U19259 (N_19259,N_19174,N_19037);
or U19260 (N_19260,N_19210,N_19249);
nand U19261 (N_19261,N_19073,N_19106);
nor U19262 (N_19262,N_19200,N_19147);
nor U19263 (N_19263,N_19244,N_19027);
nand U19264 (N_19264,N_19089,N_19092);
xor U19265 (N_19265,N_19214,N_19227);
xor U19266 (N_19266,N_19154,N_19233);
xnor U19267 (N_19267,N_19010,N_19189);
or U19268 (N_19268,N_19212,N_19095);
nand U19269 (N_19269,N_19063,N_19203);
xnor U19270 (N_19270,N_19176,N_19006);
nor U19271 (N_19271,N_19114,N_19122);
and U19272 (N_19272,N_19146,N_19240);
and U19273 (N_19273,N_19184,N_19173);
xor U19274 (N_19274,N_19008,N_19248);
xnor U19275 (N_19275,N_19126,N_19022);
nand U19276 (N_19276,N_19011,N_19129);
xnor U19277 (N_19277,N_19170,N_19130);
and U19278 (N_19278,N_19005,N_19155);
xor U19279 (N_19279,N_19071,N_19029);
and U19280 (N_19280,N_19216,N_19038);
nand U19281 (N_19281,N_19235,N_19209);
and U19282 (N_19282,N_19191,N_19243);
xor U19283 (N_19283,N_19230,N_19013);
nand U19284 (N_19284,N_19134,N_19224);
xnor U19285 (N_19285,N_19232,N_19034);
and U19286 (N_19286,N_19057,N_19099);
and U19287 (N_19287,N_19021,N_19125);
xnor U19288 (N_19288,N_19068,N_19028);
xnor U19289 (N_19289,N_19000,N_19111);
or U19290 (N_19290,N_19091,N_19165);
and U19291 (N_19291,N_19187,N_19035);
nand U19292 (N_19292,N_19199,N_19116);
nor U19293 (N_19293,N_19208,N_19054);
nand U19294 (N_19294,N_19004,N_19161);
or U19295 (N_19295,N_19058,N_19050);
and U19296 (N_19296,N_19171,N_19023);
nor U19297 (N_19297,N_19135,N_19094);
nor U19298 (N_19298,N_19198,N_19015);
or U19299 (N_19299,N_19145,N_19149);
xor U19300 (N_19300,N_19097,N_19065);
nor U19301 (N_19301,N_19012,N_19237);
xor U19302 (N_19302,N_19219,N_19084);
nor U19303 (N_19303,N_19117,N_19195);
xor U19304 (N_19304,N_19030,N_19059);
xor U19305 (N_19305,N_19064,N_19007);
nor U19306 (N_19306,N_19169,N_19040);
nor U19307 (N_19307,N_19247,N_19082);
or U19308 (N_19308,N_19078,N_19080);
or U19309 (N_19309,N_19014,N_19096);
and U19310 (N_19310,N_19143,N_19138);
and U19311 (N_19311,N_19140,N_19033);
or U19312 (N_19312,N_19047,N_19194);
nand U19313 (N_19313,N_19142,N_19115);
nor U19314 (N_19314,N_19137,N_19157);
or U19315 (N_19315,N_19204,N_19110);
xnor U19316 (N_19316,N_19223,N_19207);
nand U19317 (N_19317,N_19009,N_19231);
nor U19318 (N_19318,N_19226,N_19124);
and U19319 (N_19319,N_19156,N_19238);
nand U19320 (N_19320,N_19234,N_19236);
nand U19321 (N_19321,N_19002,N_19109);
and U19322 (N_19322,N_19090,N_19085);
or U19323 (N_19323,N_19118,N_19061);
and U19324 (N_19324,N_19018,N_19222);
or U19325 (N_19325,N_19019,N_19181);
nand U19326 (N_19326,N_19213,N_19148);
or U19327 (N_19327,N_19141,N_19105);
nand U19328 (N_19328,N_19075,N_19132);
or U19329 (N_19329,N_19093,N_19048);
nand U19330 (N_19330,N_19144,N_19104);
or U19331 (N_19331,N_19159,N_19175);
nand U19332 (N_19332,N_19024,N_19043);
or U19333 (N_19333,N_19039,N_19180);
xor U19334 (N_19334,N_19150,N_19139);
nand U19335 (N_19335,N_19152,N_19081);
nor U19336 (N_19336,N_19083,N_19190);
xnor U19337 (N_19337,N_19179,N_19026);
nand U19338 (N_19338,N_19215,N_19072);
or U19339 (N_19339,N_19121,N_19086);
and U19340 (N_19340,N_19202,N_19162);
and U19341 (N_19341,N_19045,N_19127);
nand U19342 (N_19342,N_19133,N_19206);
nor U19343 (N_19343,N_19101,N_19168);
nor U19344 (N_19344,N_19201,N_19119);
xnor U19345 (N_19345,N_19123,N_19107);
and U19346 (N_19346,N_19217,N_19074);
nor U19347 (N_19347,N_19205,N_19070);
nor U19348 (N_19348,N_19113,N_19041);
nand U19349 (N_19349,N_19100,N_19163);
nand U19350 (N_19350,N_19177,N_19131);
or U19351 (N_19351,N_19108,N_19239);
nand U19352 (N_19352,N_19020,N_19186);
and U19353 (N_19353,N_19188,N_19076);
and U19354 (N_19354,N_19167,N_19060);
xor U19355 (N_19355,N_19066,N_19242);
nand U19356 (N_19356,N_19102,N_19001);
or U19357 (N_19357,N_19151,N_19166);
and U19358 (N_19358,N_19183,N_19178);
xnor U19359 (N_19359,N_19087,N_19120);
nand U19360 (N_19360,N_19025,N_19128);
or U19361 (N_19361,N_19241,N_19246);
or U19362 (N_19362,N_19051,N_19056);
xnor U19363 (N_19363,N_19067,N_19052);
and U19364 (N_19364,N_19042,N_19153);
xnor U19365 (N_19365,N_19044,N_19077);
nand U19366 (N_19366,N_19031,N_19218);
or U19367 (N_19367,N_19225,N_19160);
or U19368 (N_19368,N_19182,N_19036);
xnor U19369 (N_19369,N_19229,N_19053);
or U19370 (N_19370,N_19136,N_19032);
nor U19371 (N_19371,N_19088,N_19220);
nor U19372 (N_19372,N_19069,N_19197);
nand U19373 (N_19373,N_19245,N_19193);
or U19374 (N_19374,N_19017,N_19185);
nand U19375 (N_19375,N_19182,N_19139);
or U19376 (N_19376,N_19079,N_19089);
xor U19377 (N_19377,N_19009,N_19138);
nor U19378 (N_19378,N_19153,N_19051);
nand U19379 (N_19379,N_19145,N_19228);
nand U19380 (N_19380,N_19245,N_19055);
xor U19381 (N_19381,N_19096,N_19104);
or U19382 (N_19382,N_19135,N_19128);
or U19383 (N_19383,N_19153,N_19028);
nand U19384 (N_19384,N_19091,N_19153);
nand U19385 (N_19385,N_19081,N_19012);
nand U19386 (N_19386,N_19033,N_19043);
nand U19387 (N_19387,N_19150,N_19200);
xor U19388 (N_19388,N_19142,N_19061);
or U19389 (N_19389,N_19017,N_19113);
and U19390 (N_19390,N_19169,N_19002);
or U19391 (N_19391,N_19181,N_19195);
nor U19392 (N_19392,N_19100,N_19158);
nor U19393 (N_19393,N_19096,N_19042);
nand U19394 (N_19394,N_19200,N_19076);
nand U19395 (N_19395,N_19176,N_19080);
nor U19396 (N_19396,N_19007,N_19053);
xnor U19397 (N_19397,N_19038,N_19095);
nor U19398 (N_19398,N_19235,N_19212);
xnor U19399 (N_19399,N_19007,N_19181);
or U19400 (N_19400,N_19111,N_19081);
or U19401 (N_19401,N_19207,N_19219);
xor U19402 (N_19402,N_19160,N_19102);
xnor U19403 (N_19403,N_19012,N_19123);
xor U19404 (N_19404,N_19187,N_19041);
and U19405 (N_19405,N_19104,N_19171);
and U19406 (N_19406,N_19211,N_19043);
nor U19407 (N_19407,N_19178,N_19166);
nand U19408 (N_19408,N_19148,N_19122);
nand U19409 (N_19409,N_19208,N_19002);
xor U19410 (N_19410,N_19221,N_19120);
or U19411 (N_19411,N_19030,N_19242);
xor U19412 (N_19412,N_19071,N_19200);
nor U19413 (N_19413,N_19208,N_19149);
or U19414 (N_19414,N_19212,N_19114);
nand U19415 (N_19415,N_19201,N_19038);
nand U19416 (N_19416,N_19197,N_19070);
and U19417 (N_19417,N_19156,N_19214);
nor U19418 (N_19418,N_19141,N_19099);
nor U19419 (N_19419,N_19177,N_19218);
nor U19420 (N_19420,N_19222,N_19051);
nand U19421 (N_19421,N_19205,N_19232);
nor U19422 (N_19422,N_19103,N_19045);
nand U19423 (N_19423,N_19000,N_19212);
nand U19424 (N_19424,N_19105,N_19072);
nand U19425 (N_19425,N_19085,N_19068);
nor U19426 (N_19426,N_19210,N_19136);
nor U19427 (N_19427,N_19193,N_19161);
xor U19428 (N_19428,N_19125,N_19080);
nor U19429 (N_19429,N_19183,N_19162);
nand U19430 (N_19430,N_19022,N_19209);
nor U19431 (N_19431,N_19011,N_19159);
and U19432 (N_19432,N_19114,N_19247);
or U19433 (N_19433,N_19188,N_19108);
xor U19434 (N_19434,N_19208,N_19038);
and U19435 (N_19435,N_19188,N_19040);
or U19436 (N_19436,N_19090,N_19190);
xnor U19437 (N_19437,N_19007,N_19065);
or U19438 (N_19438,N_19054,N_19244);
nor U19439 (N_19439,N_19235,N_19014);
xor U19440 (N_19440,N_19230,N_19249);
or U19441 (N_19441,N_19034,N_19106);
and U19442 (N_19442,N_19208,N_19089);
nor U19443 (N_19443,N_19016,N_19089);
xor U19444 (N_19444,N_19010,N_19135);
xor U19445 (N_19445,N_19237,N_19028);
or U19446 (N_19446,N_19242,N_19212);
xor U19447 (N_19447,N_19248,N_19109);
nand U19448 (N_19448,N_19147,N_19153);
and U19449 (N_19449,N_19066,N_19155);
nand U19450 (N_19450,N_19213,N_19136);
or U19451 (N_19451,N_19131,N_19121);
nand U19452 (N_19452,N_19143,N_19094);
xnor U19453 (N_19453,N_19215,N_19045);
and U19454 (N_19454,N_19213,N_19122);
xor U19455 (N_19455,N_19192,N_19043);
or U19456 (N_19456,N_19142,N_19184);
or U19457 (N_19457,N_19239,N_19067);
and U19458 (N_19458,N_19050,N_19075);
nor U19459 (N_19459,N_19107,N_19099);
nand U19460 (N_19460,N_19070,N_19235);
nand U19461 (N_19461,N_19133,N_19172);
and U19462 (N_19462,N_19195,N_19029);
nand U19463 (N_19463,N_19118,N_19221);
and U19464 (N_19464,N_19191,N_19212);
nor U19465 (N_19465,N_19020,N_19161);
nand U19466 (N_19466,N_19011,N_19119);
and U19467 (N_19467,N_19245,N_19083);
xor U19468 (N_19468,N_19139,N_19061);
nand U19469 (N_19469,N_19246,N_19203);
and U19470 (N_19470,N_19198,N_19008);
xnor U19471 (N_19471,N_19061,N_19117);
xnor U19472 (N_19472,N_19145,N_19059);
nand U19473 (N_19473,N_19041,N_19049);
nor U19474 (N_19474,N_19057,N_19051);
or U19475 (N_19475,N_19036,N_19220);
or U19476 (N_19476,N_19057,N_19058);
nor U19477 (N_19477,N_19060,N_19192);
xor U19478 (N_19478,N_19147,N_19152);
nor U19479 (N_19479,N_19064,N_19217);
nor U19480 (N_19480,N_19173,N_19087);
and U19481 (N_19481,N_19015,N_19226);
nor U19482 (N_19482,N_19242,N_19168);
xor U19483 (N_19483,N_19199,N_19014);
and U19484 (N_19484,N_19024,N_19062);
and U19485 (N_19485,N_19178,N_19173);
nand U19486 (N_19486,N_19113,N_19232);
or U19487 (N_19487,N_19220,N_19055);
or U19488 (N_19488,N_19108,N_19111);
xnor U19489 (N_19489,N_19133,N_19084);
or U19490 (N_19490,N_19188,N_19207);
xnor U19491 (N_19491,N_19049,N_19037);
or U19492 (N_19492,N_19186,N_19236);
or U19493 (N_19493,N_19193,N_19242);
xor U19494 (N_19494,N_19107,N_19095);
xnor U19495 (N_19495,N_19145,N_19131);
nand U19496 (N_19496,N_19074,N_19156);
and U19497 (N_19497,N_19131,N_19232);
nor U19498 (N_19498,N_19167,N_19049);
or U19499 (N_19499,N_19163,N_19006);
or U19500 (N_19500,N_19469,N_19358);
or U19501 (N_19501,N_19433,N_19266);
and U19502 (N_19502,N_19259,N_19462);
xnor U19503 (N_19503,N_19353,N_19456);
nand U19504 (N_19504,N_19264,N_19394);
or U19505 (N_19505,N_19306,N_19269);
xor U19506 (N_19506,N_19274,N_19432);
and U19507 (N_19507,N_19333,N_19477);
nor U19508 (N_19508,N_19430,N_19310);
or U19509 (N_19509,N_19389,N_19361);
and U19510 (N_19510,N_19287,N_19261);
nor U19511 (N_19511,N_19341,N_19263);
nor U19512 (N_19512,N_19258,N_19260);
or U19513 (N_19513,N_19444,N_19290);
or U19514 (N_19514,N_19450,N_19386);
nor U19515 (N_19515,N_19408,N_19443);
nor U19516 (N_19516,N_19422,N_19418);
and U19517 (N_19517,N_19344,N_19347);
nand U19518 (N_19518,N_19472,N_19338);
nor U19519 (N_19519,N_19385,N_19409);
or U19520 (N_19520,N_19465,N_19268);
and U19521 (N_19521,N_19334,N_19379);
nor U19522 (N_19522,N_19271,N_19357);
nand U19523 (N_19523,N_19425,N_19371);
nand U19524 (N_19524,N_19499,N_19359);
nor U19525 (N_19525,N_19317,N_19478);
nor U19526 (N_19526,N_19283,N_19404);
xnor U19527 (N_19527,N_19452,N_19281);
and U19528 (N_19528,N_19467,N_19415);
or U19529 (N_19529,N_19391,N_19336);
xor U19530 (N_19530,N_19479,N_19332);
and U19531 (N_19531,N_19284,N_19340);
and U19532 (N_19532,N_19364,N_19327);
and U19533 (N_19533,N_19449,N_19390);
nand U19534 (N_19534,N_19454,N_19460);
nand U19535 (N_19535,N_19368,N_19262);
xor U19536 (N_19536,N_19291,N_19400);
xnor U19537 (N_19537,N_19343,N_19459);
xor U19538 (N_19538,N_19257,N_19380);
nor U19539 (N_19539,N_19407,N_19303);
and U19540 (N_19540,N_19346,N_19267);
or U19541 (N_19541,N_19314,N_19481);
nand U19542 (N_19542,N_19475,N_19382);
or U19543 (N_19543,N_19277,N_19272);
and U19544 (N_19544,N_19435,N_19427);
and U19545 (N_19545,N_19419,N_19270);
nor U19546 (N_19546,N_19490,N_19378);
xnor U19547 (N_19547,N_19410,N_19292);
nor U19548 (N_19548,N_19365,N_19455);
and U19549 (N_19549,N_19484,N_19285);
or U19550 (N_19550,N_19253,N_19486);
or U19551 (N_19551,N_19476,N_19423);
and U19552 (N_19552,N_19383,N_19250);
nor U19553 (N_19553,N_19473,N_19316);
nor U19554 (N_19554,N_19335,N_19313);
xor U19555 (N_19555,N_19405,N_19298);
and U19556 (N_19556,N_19296,N_19331);
and U19557 (N_19557,N_19488,N_19416);
nand U19558 (N_19558,N_19437,N_19482);
and U19559 (N_19559,N_19480,N_19330);
and U19560 (N_19560,N_19373,N_19397);
nor U19561 (N_19561,N_19363,N_19273);
or U19562 (N_19562,N_19381,N_19497);
and U19563 (N_19563,N_19318,N_19302);
xnor U19564 (N_19564,N_19339,N_19375);
and U19565 (N_19565,N_19337,N_19352);
and U19566 (N_19566,N_19282,N_19278);
nand U19567 (N_19567,N_19300,N_19426);
or U19568 (N_19568,N_19288,N_19402);
or U19569 (N_19569,N_19436,N_19256);
xnor U19570 (N_19570,N_19320,N_19464);
nand U19571 (N_19571,N_19312,N_19401);
and U19572 (N_19572,N_19360,N_19463);
or U19573 (N_19573,N_19305,N_19376);
xnor U19574 (N_19574,N_19439,N_19275);
or U19575 (N_19575,N_19279,N_19398);
or U19576 (N_19576,N_19414,N_19325);
nor U19577 (N_19577,N_19498,N_19362);
nand U19578 (N_19578,N_19474,N_19252);
and U19579 (N_19579,N_19293,N_19417);
and U19580 (N_19580,N_19307,N_19280);
xnor U19581 (N_19581,N_19342,N_19495);
and U19582 (N_19582,N_19491,N_19461);
and U19583 (N_19583,N_19406,N_19424);
and U19584 (N_19584,N_19251,N_19388);
or U19585 (N_19585,N_19326,N_19384);
or U19586 (N_19586,N_19294,N_19276);
xnor U19587 (N_19587,N_19315,N_19483);
and U19588 (N_19588,N_19319,N_19489);
or U19589 (N_19589,N_19255,N_19487);
nand U19590 (N_19590,N_19457,N_19420);
and U19591 (N_19591,N_19345,N_19392);
xor U19592 (N_19592,N_19370,N_19369);
nand U19593 (N_19593,N_19468,N_19453);
or U19594 (N_19594,N_19458,N_19297);
and U19595 (N_19595,N_19299,N_19354);
nor U19596 (N_19596,N_19399,N_19393);
nand U19597 (N_19597,N_19309,N_19412);
nand U19598 (N_19598,N_19329,N_19441);
nor U19599 (N_19599,N_19289,N_19254);
and U19600 (N_19600,N_19366,N_19440);
nor U19601 (N_19601,N_19470,N_19311);
xor U19602 (N_19602,N_19321,N_19403);
or U19603 (N_19603,N_19367,N_19429);
xnor U19604 (N_19604,N_19411,N_19377);
nor U19605 (N_19605,N_19351,N_19348);
nor U19606 (N_19606,N_19421,N_19295);
nand U19607 (N_19607,N_19451,N_19355);
xnor U19608 (N_19608,N_19328,N_19356);
xor U19609 (N_19609,N_19349,N_19438);
and U19610 (N_19610,N_19304,N_19322);
xor U19611 (N_19611,N_19442,N_19485);
nand U19612 (N_19612,N_19471,N_19448);
or U19613 (N_19613,N_19350,N_19372);
xnor U19614 (N_19614,N_19323,N_19395);
nor U19615 (N_19615,N_19308,N_19413);
or U19616 (N_19616,N_19324,N_19374);
nor U19617 (N_19617,N_19446,N_19434);
xor U19618 (N_19618,N_19492,N_19431);
or U19619 (N_19619,N_19466,N_19286);
or U19620 (N_19620,N_19447,N_19493);
nand U19621 (N_19621,N_19445,N_19428);
xor U19622 (N_19622,N_19301,N_19496);
or U19623 (N_19623,N_19387,N_19265);
xnor U19624 (N_19624,N_19494,N_19396);
nand U19625 (N_19625,N_19388,N_19410);
xnor U19626 (N_19626,N_19404,N_19250);
xor U19627 (N_19627,N_19355,N_19438);
and U19628 (N_19628,N_19400,N_19499);
xnor U19629 (N_19629,N_19358,N_19309);
xnor U19630 (N_19630,N_19261,N_19443);
nand U19631 (N_19631,N_19289,N_19451);
or U19632 (N_19632,N_19293,N_19410);
nor U19633 (N_19633,N_19424,N_19366);
nor U19634 (N_19634,N_19450,N_19296);
xnor U19635 (N_19635,N_19454,N_19423);
xnor U19636 (N_19636,N_19375,N_19429);
nor U19637 (N_19637,N_19383,N_19313);
nand U19638 (N_19638,N_19455,N_19465);
nand U19639 (N_19639,N_19275,N_19265);
or U19640 (N_19640,N_19410,N_19489);
or U19641 (N_19641,N_19403,N_19417);
nor U19642 (N_19642,N_19251,N_19334);
nand U19643 (N_19643,N_19306,N_19377);
or U19644 (N_19644,N_19257,N_19365);
or U19645 (N_19645,N_19484,N_19345);
nand U19646 (N_19646,N_19463,N_19426);
and U19647 (N_19647,N_19399,N_19483);
nand U19648 (N_19648,N_19262,N_19302);
or U19649 (N_19649,N_19458,N_19251);
nand U19650 (N_19650,N_19289,N_19359);
or U19651 (N_19651,N_19428,N_19415);
or U19652 (N_19652,N_19371,N_19390);
or U19653 (N_19653,N_19489,N_19416);
nor U19654 (N_19654,N_19465,N_19351);
or U19655 (N_19655,N_19365,N_19252);
and U19656 (N_19656,N_19296,N_19447);
nor U19657 (N_19657,N_19380,N_19365);
nand U19658 (N_19658,N_19453,N_19263);
nor U19659 (N_19659,N_19351,N_19343);
nand U19660 (N_19660,N_19389,N_19445);
and U19661 (N_19661,N_19353,N_19281);
nor U19662 (N_19662,N_19368,N_19332);
or U19663 (N_19663,N_19256,N_19365);
and U19664 (N_19664,N_19466,N_19325);
xnor U19665 (N_19665,N_19261,N_19497);
xor U19666 (N_19666,N_19401,N_19345);
and U19667 (N_19667,N_19474,N_19380);
and U19668 (N_19668,N_19358,N_19333);
nor U19669 (N_19669,N_19459,N_19307);
or U19670 (N_19670,N_19263,N_19347);
xor U19671 (N_19671,N_19412,N_19361);
nor U19672 (N_19672,N_19429,N_19492);
and U19673 (N_19673,N_19366,N_19309);
nand U19674 (N_19674,N_19323,N_19259);
and U19675 (N_19675,N_19398,N_19456);
xor U19676 (N_19676,N_19304,N_19343);
xnor U19677 (N_19677,N_19314,N_19393);
xnor U19678 (N_19678,N_19379,N_19450);
or U19679 (N_19679,N_19266,N_19327);
or U19680 (N_19680,N_19278,N_19374);
or U19681 (N_19681,N_19333,N_19393);
or U19682 (N_19682,N_19321,N_19497);
nand U19683 (N_19683,N_19346,N_19261);
nor U19684 (N_19684,N_19437,N_19350);
nor U19685 (N_19685,N_19291,N_19369);
xnor U19686 (N_19686,N_19276,N_19260);
xnor U19687 (N_19687,N_19284,N_19348);
nand U19688 (N_19688,N_19436,N_19271);
or U19689 (N_19689,N_19483,N_19358);
and U19690 (N_19690,N_19339,N_19411);
nor U19691 (N_19691,N_19330,N_19297);
xor U19692 (N_19692,N_19343,N_19293);
nand U19693 (N_19693,N_19411,N_19458);
nand U19694 (N_19694,N_19443,N_19447);
xnor U19695 (N_19695,N_19315,N_19426);
xor U19696 (N_19696,N_19347,N_19314);
or U19697 (N_19697,N_19328,N_19363);
nor U19698 (N_19698,N_19329,N_19477);
xnor U19699 (N_19699,N_19337,N_19273);
and U19700 (N_19700,N_19283,N_19464);
and U19701 (N_19701,N_19499,N_19334);
and U19702 (N_19702,N_19498,N_19435);
and U19703 (N_19703,N_19270,N_19338);
xor U19704 (N_19704,N_19462,N_19407);
xor U19705 (N_19705,N_19254,N_19463);
nor U19706 (N_19706,N_19264,N_19453);
nand U19707 (N_19707,N_19429,N_19468);
or U19708 (N_19708,N_19282,N_19491);
and U19709 (N_19709,N_19264,N_19285);
nor U19710 (N_19710,N_19272,N_19257);
nand U19711 (N_19711,N_19256,N_19460);
or U19712 (N_19712,N_19287,N_19497);
and U19713 (N_19713,N_19473,N_19428);
or U19714 (N_19714,N_19423,N_19278);
xor U19715 (N_19715,N_19426,N_19475);
or U19716 (N_19716,N_19430,N_19452);
and U19717 (N_19717,N_19314,N_19475);
or U19718 (N_19718,N_19371,N_19356);
and U19719 (N_19719,N_19451,N_19479);
and U19720 (N_19720,N_19427,N_19297);
nor U19721 (N_19721,N_19466,N_19409);
nor U19722 (N_19722,N_19367,N_19423);
nor U19723 (N_19723,N_19381,N_19396);
and U19724 (N_19724,N_19277,N_19400);
nand U19725 (N_19725,N_19263,N_19340);
nand U19726 (N_19726,N_19452,N_19308);
nor U19727 (N_19727,N_19387,N_19394);
nand U19728 (N_19728,N_19371,N_19260);
xor U19729 (N_19729,N_19326,N_19405);
nor U19730 (N_19730,N_19340,N_19474);
xor U19731 (N_19731,N_19281,N_19330);
nor U19732 (N_19732,N_19343,N_19332);
xnor U19733 (N_19733,N_19442,N_19306);
xnor U19734 (N_19734,N_19345,N_19340);
or U19735 (N_19735,N_19397,N_19355);
and U19736 (N_19736,N_19384,N_19382);
nor U19737 (N_19737,N_19317,N_19499);
nand U19738 (N_19738,N_19409,N_19476);
or U19739 (N_19739,N_19454,N_19309);
and U19740 (N_19740,N_19441,N_19433);
xor U19741 (N_19741,N_19369,N_19386);
nor U19742 (N_19742,N_19255,N_19273);
and U19743 (N_19743,N_19419,N_19440);
nor U19744 (N_19744,N_19337,N_19264);
xnor U19745 (N_19745,N_19324,N_19298);
nand U19746 (N_19746,N_19434,N_19252);
nor U19747 (N_19747,N_19263,N_19267);
or U19748 (N_19748,N_19439,N_19324);
nor U19749 (N_19749,N_19285,N_19496);
xor U19750 (N_19750,N_19615,N_19524);
nor U19751 (N_19751,N_19613,N_19671);
xnor U19752 (N_19752,N_19656,N_19607);
nand U19753 (N_19753,N_19568,N_19601);
nor U19754 (N_19754,N_19534,N_19717);
and U19755 (N_19755,N_19580,N_19547);
and U19756 (N_19756,N_19542,N_19522);
and U19757 (N_19757,N_19558,N_19579);
or U19758 (N_19758,N_19609,N_19710);
and U19759 (N_19759,N_19508,N_19632);
or U19760 (N_19760,N_19606,N_19647);
or U19761 (N_19761,N_19749,N_19741);
nor U19762 (N_19762,N_19640,N_19659);
xor U19763 (N_19763,N_19564,N_19629);
nand U19764 (N_19764,N_19636,N_19748);
nor U19765 (N_19765,N_19502,N_19514);
and U19766 (N_19766,N_19589,N_19562);
or U19767 (N_19767,N_19718,N_19517);
xor U19768 (N_19768,N_19628,N_19667);
nor U19769 (N_19769,N_19618,N_19669);
or U19770 (N_19770,N_19592,N_19721);
and U19771 (N_19771,N_19588,N_19702);
nand U19772 (N_19772,N_19704,N_19708);
or U19773 (N_19773,N_19590,N_19673);
nor U19774 (N_19774,N_19712,N_19641);
nor U19775 (N_19775,N_19675,N_19544);
nor U19776 (N_19776,N_19674,N_19706);
xnor U19777 (N_19777,N_19739,N_19614);
nor U19778 (N_19778,N_19528,N_19696);
nand U19779 (N_19779,N_19596,N_19678);
xor U19780 (N_19780,N_19652,N_19597);
and U19781 (N_19781,N_19604,N_19620);
xor U19782 (N_19782,N_19593,N_19740);
nor U19783 (N_19783,N_19505,N_19716);
or U19784 (N_19784,N_19627,N_19500);
or U19785 (N_19785,N_19738,N_19693);
or U19786 (N_19786,N_19556,N_19577);
or U19787 (N_19787,N_19648,N_19503);
nor U19788 (N_19788,N_19680,N_19683);
and U19789 (N_19789,N_19668,N_19643);
and U19790 (N_19790,N_19713,N_19637);
or U19791 (N_19791,N_19584,N_19733);
nor U19792 (N_19792,N_19681,N_19504);
and U19793 (N_19793,N_19682,N_19638);
and U19794 (N_19794,N_19552,N_19545);
xor U19795 (N_19795,N_19605,N_19539);
nor U19796 (N_19796,N_19530,N_19676);
and U19797 (N_19797,N_19582,N_19744);
nor U19798 (N_19798,N_19662,N_19655);
or U19799 (N_19799,N_19536,N_19543);
nand U19800 (N_19800,N_19561,N_19714);
and U19801 (N_19801,N_19595,N_19688);
or U19802 (N_19802,N_19625,N_19623);
xor U19803 (N_19803,N_19571,N_19666);
and U19804 (N_19804,N_19583,N_19690);
and U19805 (N_19805,N_19694,N_19695);
nor U19806 (N_19806,N_19684,N_19569);
nor U19807 (N_19807,N_19722,N_19518);
xnor U19808 (N_19808,N_19521,N_19506);
nor U19809 (N_19809,N_19573,N_19730);
xnor U19810 (N_19810,N_19709,N_19723);
or U19811 (N_19811,N_19711,N_19520);
and U19812 (N_19812,N_19549,N_19516);
nand U19813 (N_19813,N_19698,N_19523);
nand U19814 (N_19814,N_19566,N_19649);
or U19815 (N_19815,N_19600,N_19519);
xor U19816 (N_19816,N_19617,N_19700);
nand U19817 (N_19817,N_19576,N_19670);
nand U19818 (N_19818,N_19715,N_19538);
xor U19819 (N_19819,N_19574,N_19554);
nor U19820 (N_19820,N_19575,N_19546);
nand U19821 (N_19821,N_19701,N_19586);
or U19822 (N_19822,N_19531,N_19642);
nand U19823 (N_19823,N_19626,N_19624);
and U19824 (N_19824,N_19509,N_19663);
nor U19825 (N_19825,N_19540,N_19705);
or U19826 (N_19826,N_19557,N_19731);
and U19827 (N_19827,N_19719,N_19634);
xor U19828 (N_19828,N_19532,N_19732);
nor U19829 (N_19829,N_19535,N_19687);
nand U19830 (N_19830,N_19707,N_19581);
and U19831 (N_19831,N_19631,N_19737);
and U19832 (N_19832,N_19585,N_19658);
and U19833 (N_19833,N_19570,N_19512);
and U19834 (N_19834,N_19720,N_19664);
nand U19835 (N_19835,N_19529,N_19622);
nor U19836 (N_19836,N_19507,N_19745);
nand U19837 (N_19837,N_19555,N_19699);
or U19838 (N_19838,N_19651,N_19677);
and U19839 (N_19839,N_19526,N_19525);
nor U19840 (N_19840,N_19563,N_19560);
xor U19841 (N_19841,N_19559,N_19728);
nor U19842 (N_19842,N_19515,N_19639);
xnor U19843 (N_19843,N_19567,N_19644);
nand U19844 (N_19844,N_19725,N_19510);
nand U19845 (N_19845,N_19550,N_19691);
nand U19846 (N_19846,N_19513,N_19729);
xor U19847 (N_19847,N_19501,N_19511);
xor U19848 (N_19848,N_19591,N_19686);
xor U19849 (N_19849,N_19742,N_19621);
nand U19850 (N_19850,N_19533,N_19735);
xnor U19851 (N_19851,N_19653,N_19743);
and U19852 (N_19852,N_19541,N_19726);
nand U19853 (N_19853,N_19602,N_19672);
or U19854 (N_19854,N_19608,N_19650);
and U19855 (N_19855,N_19635,N_19537);
nand U19856 (N_19856,N_19599,N_19610);
xnor U19857 (N_19857,N_19734,N_19685);
xnor U19858 (N_19858,N_19724,N_19689);
or U19859 (N_19859,N_19548,N_19603);
xor U19860 (N_19860,N_19616,N_19660);
and U19861 (N_19861,N_19594,N_19598);
xnor U19862 (N_19862,N_19697,N_19727);
or U19863 (N_19863,N_19527,N_19645);
xor U19864 (N_19864,N_19630,N_19612);
nand U19865 (N_19865,N_19587,N_19553);
nor U19866 (N_19866,N_19633,N_19747);
and U19867 (N_19867,N_19551,N_19565);
xnor U19868 (N_19868,N_19679,N_19746);
nor U19869 (N_19869,N_19665,N_19692);
xor U19870 (N_19870,N_19657,N_19703);
nor U19871 (N_19871,N_19654,N_19572);
nand U19872 (N_19872,N_19611,N_19578);
nand U19873 (N_19873,N_19661,N_19736);
nor U19874 (N_19874,N_19619,N_19646);
nor U19875 (N_19875,N_19600,N_19607);
or U19876 (N_19876,N_19649,N_19600);
nor U19877 (N_19877,N_19557,N_19746);
xnor U19878 (N_19878,N_19710,N_19701);
or U19879 (N_19879,N_19699,N_19626);
or U19880 (N_19880,N_19538,N_19601);
nor U19881 (N_19881,N_19560,N_19625);
and U19882 (N_19882,N_19712,N_19561);
xnor U19883 (N_19883,N_19701,N_19674);
or U19884 (N_19884,N_19739,N_19615);
nor U19885 (N_19885,N_19628,N_19676);
and U19886 (N_19886,N_19613,N_19743);
and U19887 (N_19887,N_19623,N_19645);
or U19888 (N_19888,N_19598,N_19722);
and U19889 (N_19889,N_19616,N_19651);
nor U19890 (N_19890,N_19634,N_19517);
and U19891 (N_19891,N_19671,N_19510);
and U19892 (N_19892,N_19657,N_19720);
nor U19893 (N_19893,N_19582,N_19623);
nor U19894 (N_19894,N_19636,N_19731);
nor U19895 (N_19895,N_19596,N_19654);
or U19896 (N_19896,N_19530,N_19660);
nor U19897 (N_19897,N_19585,N_19644);
and U19898 (N_19898,N_19613,N_19651);
or U19899 (N_19899,N_19501,N_19623);
xor U19900 (N_19900,N_19661,N_19618);
or U19901 (N_19901,N_19564,N_19725);
and U19902 (N_19902,N_19635,N_19693);
nor U19903 (N_19903,N_19601,N_19577);
or U19904 (N_19904,N_19646,N_19690);
or U19905 (N_19905,N_19606,N_19733);
and U19906 (N_19906,N_19649,N_19736);
and U19907 (N_19907,N_19519,N_19512);
and U19908 (N_19908,N_19648,N_19699);
and U19909 (N_19909,N_19672,N_19643);
nor U19910 (N_19910,N_19695,N_19701);
nor U19911 (N_19911,N_19539,N_19743);
nor U19912 (N_19912,N_19510,N_19656);
and U19913 (N_19913,N_19720,N_19691);
nand U19914 (N_19914,N_19576,N_19629);
or U19915 (N_19915,N_19674,N_19642);
or U19916 (N_19916,N_19602,N_19722);
nand U19917 (N_19917,N_19609,N_19605);
nand U19918 (N_19918,N_19669,N_19512);
and U19919 (N_19919,N_19506,N_19721);
xnor U19920 (N_19920,N_19694,N_19727);
nor U19921 (N_19921,N_19556,N_19571);
xor U19922 (N_19922,N_19637,N_19660);
xnor U19923 (N_19923,N_19527,N_19586);
and U19924 (N_19924,N_19707,N_19500);
or U19925 (N_19925,N_19708,N_19729);
nand U19926 (N_19926,N_19733,N_19682);
or U19927 (N_19927,N_19569,N_19561);
nor U19928 (N_19928,N_19736,N_19505);
nand U19929 (N_19929,N_19637,N_19721);
nor U19930 (N_19930,N_19646,N_19598);
nand U19931 (N_19931,N_19650,N_19687);
xnor U19932 (N_19932,N_19597,N_19704);
nand U19933 (N_19933,N_19656,N_19739);
nand U19934 (N_19934,N_19697,N_19544);
nand U19935 (N_19935,N_19645,N_19721);
or U19936 (N_19936,N_19509,N_19586);
nor U19937 (N_19937,N_19690,N_19660);
xnor U19938 (N_19938,N_19567,N_19594);
and U19939 (N_19939,N_19600,N_19642);
xnor U19940 (N_19940,N_19743,N_19710);
xor U19941 (N_19941,N_19731,N_19628);
nand U19942 (N_19942,N_19747,N_19514);
and U19943 (N_19943,N_19536,N_19597);
or U19944 (N_19944,N_19626,N_19704);
xor U19945 (N_19945,N_19737,N_19686);
nand U19946 (N_19946,N_19654,N_19653);
xor U19947 (N_19947,N_19531,N_19547);
nand U19948 (N_19948,N_19632,N_19665);
xnor U19949 (N_19949,N_19639,N_19503);
xor U19950 (N_19950,N_19542,N_19717);
and U19951 (N_19951,N_19658,N_19514);
xnor U19952 (N_19952,N_19743,N_19603);
nand U19953 (N_19953,N_19741,N_19713);
and U19954 (N_19954,N_19658,N_19531);
nand U19955 (N_19955,N_19699,N_19622);
and U19956 (N_19956,N_19555,N_19674);
and U19957 (N_19957,N_19681,N_19688);
nor U19958 (N_19958,N_19645,N_19637);
xnor U19959 (N_19959,N_19715,N_19689);
or U19960 (N_19960,N_19561,N_19653);
xor U19961 (N_19961,N_19738,N_19547);
xor U19962 (N_19962,N_19746,N_19550);
nand U19963 (N_19963,N_19663,N_19548);
xor U19964 (N_19964,N_19582,N_19636);
nor U19965 (N_19965,N_19586,N_19535);
nand U19966 (N_19966,N_19537,N_19731);
and U19967 (N_19967,N_19628,N_19641);
xnor U19968 (N_19968,N_19646,N_19604);
nand U19969 (N_19969,N_19603,N_19581);
nor U19970 (N_19970,N_19656,N_19665);
xnor U19971 (N_19971,N_19525,N_19646);
xnor U19972 (N_19972,N_19681,N_19544);
or U19973 (N_19973,N_19692,N_19660);
and U19974 (N_19974,N_19733,N_19533);
nor U19975 (N_19975,N_19546,N_19595);
xor U19976 (N_19976,N_19700,N_19717);
or U19977 (N_19977,N_19635,N_19625);
nor U19978 (N_19978,N_19548,N_19720);
or U19979 (N_19979,N_19638,N_19609);
or U19980 (N_19980,N_19624,N_19642);
nand U19981 (N_19981,N_19530,N_19687);
and U19982 (N_19982,N_19608,N_19660);
nand U19983 (N_19983,N_19609,N_19645);
xor U19984 (N_19984,N_19638,N_19670);
and U19985 (N_19985,N_19684,N_19681);
nor U19986 (N_19986,N_19731,N_19647);
and U19987 (N_19987,N_19679,N_19649);
xor U19988 (N_19988,N_19624,N_19693);
or U19989 (N_19989,N_19660,N_19667);
nor U19990 (N_19990,N_19509,N_19596);
and U19991 (N_19991,N_19729,N_19716);
nor U19992 (N_19992,N_19635,N_19741);
nor U19993 (N_19993,N_19575,N_19527);
nor U19994 (N_19994,N_19644,N_19624);
nand U19995 (N_19995,N_19749,N_19742);
nor U19996 (N_19996,N_19511,N_19508);
or U19997 (N_19997,N_19619,N_19548);
nor U19998 (N_19998,N_19553,N_19748);
and U19999 (N_19999,N_19737,N_19696);
or U20000 (N_20000,N_19908,N_19968);
xor U20001 (N_20001,N_19761,N_19927);
xnor U20002 (N_20002,N_19843,N_19881);
nor U20003 (N_20003,N_19943,N_19994);
nand U20004 (N_20004,N_19829,N_19816);
or U20005 (N_20005,N_19991,N_19999);
and U20006 (N_20006,N_19897,N_19872);
xor U20007 (N_20007,N_19988,N_19824);
or U20008 (N_20008,N_19993,N_19952);
nand U20009 (N_20009,N_19955,N_19808);
and U20010 (N_20010,N_19768,N_19800);
nand U20011 (N_20011,N_19982,N_19811);
and U20012 (N_20012,N_19856,N_19756);
or U20013 (N_20013,N_19951,N_19882);
or U20014 (N_20014,N_19821,N_19842);
and U20015 (N_20015,N_19967,N_19828);
nand U20016 (N_20016,N_19896,N_19774);
or U20017 (N_20017,N_19960,N_19849);
nor U20018 (N_20018,N_19794,N_19823);
xnor U20019 (N_20019,N_19846,N_19911);
and U20020 (N_20020,N_19876,N_19760);
nor U20021 (N_20021,N_19832,N_19889);
or U20022 (N_20022,N_19962,N_19932);
nand U20023 (N_20023,N_19797,N_19894);
or U20024 (N_20024,N_19961,N_19924);
or U20025 (N_20025,N_19840,N_19963);
and U20026 (N_20026,N_19783,N_19914);
or U20027 (N_20027,N_19959,N_19948);
xor U20028 (N_20028,N_19975,N_19771);
nor U20029 (N_20029,N_19877,N_19984);
nand U20030 (N_20030,N_19980,N_19901);
or U20031 (N_20031,N_19772,N_19930);
xnor U20032 (N_20032,N_19778,N_19874);
and U20033 (N_20033,N_19972,N_19921);
nand U20034 (N_20034,N_19766,N_19786);
or U20035 (N_20035,N_19986,N_19946);
nor U20036 (N_20036,N_19989,N_19825);
and U20037 (N_20037,N_19936,N_19998);
nor U20038 (N_20038,N_19933,N_19945);
nand U20039 (N_20039,N_19806,N_19868);
and U20040 (N_20040,N_19965,N_19789);
or U20041 (N_20041,N_19787,N_19848);
xnor U20042 (N_20042,N_19865,N_19983);
and U20043 (N_20043,N_19906,N_19819);
and U20044 (N_20044,N_19995,N_19807);
nor U20045 (N_20045,N_19770,N_19866);
and U20046 (N_20046,N_19922,N_19871);
nand U20047 (N_20047,N_19859,N_19754);
or U20048 (N_20048,N_19940,N_19979);
and U20049 (N_20049,N_19895,N_19903);
nand U20050 (N_20050,N_19854,N_19857);
xor U20051 (N_20051,N_19973,N_19785);
nand U20052 (N_20052,N_19947,N_19841);
or U20053 (N_20053,N_19827,N_19801);
nand U20054 (N_20054,N_19929,N_19904);
or U20055 (N_20055,N_19913,N_19822);
nand U20056 (N_20056,N_19831,N_19950);
and U20057 (N_20057,N_19835,N_19833);
and U20058 (N_20058,N_19905,N_19956);
nand U20059 (N_20059,N_19862,N_19870);
or U20060 (N_20060,N_19875,N_19753);
xnor U20061 (N_20061,N_19867,N_19869);
nor U20062 (N_20062,N_19757,N_19902);
nand U20063 (N_20063,N_19958,N_19817);
nand U20064 (N_20064,N_19907,N_19773);
nand U20065 (N_20065,N_19969,N_19939);
xnor U20066 (N_20066,N_19981,N_19977);
and U20067 (N_20067,N_19953,N_19751);
xor U20068 (N_20068,N_19917,N_19853);
or U20069 (N_20069,N_19971,N_19818);
or U20070 (N_20070,N_19750,N_19812);
nand U20071 (N_20071,N_19918,N_19762);
or U20072 (N_20072,N_19796,N_19851);
and U20073 (N_20073,N_19809,N_19777);
or U20074 (N_20074,N_19852,N_19855);
xnor U20075 (N_20075,N_19893,N_19931);
or U20076 (N_20076,N_19873,N_19863);
nor U20077 (N_20077,N_19949,N_19923);
nor U20078 (N_20078,N_19780,N_19944);
or U20079 (N_20079,N_19996,N_19891);
nand U20080 (N_20080,N_19820,N_19758);
xor U20081 (N_20081,N_19860,N_19966);
and U20082 (N_20082,N_19779,N_19810);
nor U20083 (N_20083,N_19784,N_19954);
and U20084 (N_20084,N_19805,N_19795);
nand U20085 (N_20085,N_19992,N_19765);
nor U20086 (N_20086,N_19976,N_19957);
nand U20087 (N_20087,N_19899,N_19888);
nor U20088 (N_20088,N_19916,N_19997);
and U20089 (N_20089,N_19826,N_19798);
and U20090 (N_20090,N_19781,N_19883);
nand U20091 (N_20091,N_19978,N_19964);
or U20092 (N_20092,N_19804,N_19799);
nand U20093 (N_20093,N_19892,N_19941);
xnor U20094 (N_20094,N_19878,N_19813);
nand U20095 (N_20095,N_19900,N_19792);
or U20096 (N_20096,N_19755,N_19884);
nand U20097 (N_20097,N_19938,N_19769);
nand U20098 (N_20098,N_19839,N_19858);
or U20099 (N_20099,N_19987,N_19887);
nand U20100 (N_20100,N_19844,N_19802);
nand U20101 (N_20101,N_19974,N_19898);
or U20102 (N_20102,N_19942,N_19788);
xnor U20103 (N_20103,N_19937,N_19886);
nand U20104 (N_20104,N_19838,N_19934);
nand U20105 (N_20105,N_19910,N_19880);
and U20106 (N_20106,N_19764,N_19850);
xnor U20107 (N_20107,N_19925,N_19912);
nand U20108 (N_20108,N_19836,N_19752);
or U20109 (N_20109,N_19763,N_19776);
nor U20110 (N_20110,N_19928,N_19885);
nand U20111 (N_20111,N_19775,N_19815);
and U20112 (N_20112,N_19935,N_19814);
and U20113 (N_20113,N_19845,N_19864);
xnor U20114 (N_20114,N_19834,N_19909);
nor U20115 (N_20115,N_19830,N_19879);
xnor U20116 (N_20116,N_19861,N_19890);
nand U20117 (N_20117,N_19985,N_19926);
nor U20118 (N_20118,N_19920,N_19759);
and U20119 (N_20119,N_19782,N_19990);
nor U20120 (N_20120,N_19791,N_19767);
nand U20121 (N_20121,N_19803,N_19790);
xor U20122 (N_20122,N_19837,N_19847);
or U20123 (N_20123,N_19915,N_19970);
nor U20124 (N_20124,N_19919,N_19793);
xor U20125 (N_20125,N_19906,N_19977);
nand U20126 (N_20126,N_19796,N_19974);
nor U20127 (N_20127,N_19776,N_19786);
xor U20128 (N_20128,N_19828,N_19790);
nand U20129 (N_20129,N_19930,N_19937);
and U20130 (N_20130,N_19991,N_19866);
xnor U20131 (N_20131,N_19873,N_19837);
nor U20132 (N_20132,N_19891,N_19826);
nor U20133 (N_20133,N_19901,N_19869);
nand U20134 (N_20134,N_19918,N_19959);
nor U20135 (N_20135,N_19810,N_19977);
nor U20136 (N_20136,N_19812,N_19803);
and U20137 (N_20137,N_19872,N_19963);
xor U20138 (N_20138,N_19900,N_19969);
or U20139 (N_20139,N_19816,N_19803);
or U20140 (N_20140,N_19828,N_19934);
or U20141 (N_20141,N_19795,N_19933);
xor U20142 (N_20142,N_19819,N_19915);
nor U20143 (N_20143,N_19797,N_19943);
and U20144 (N_20144,N_19791,N_19814);
and U20145 (N_20145,N_19870,N_19768);
nand U20146 (N_20146,N_19810,N_19812);
nor U20147 (N_20147,N_19832,N_19920);
or U20148 (N_20148,N_19939,N_19828);
or U20149 (N_20149,N_19791,N_19981);
or U20150 (N_20150,N_19848,N_19857);
nor U20151 (N_20151,N_19838,N_19926);
nor U20152 (N_20152,N_19978,N_19969);
xor U20153 (N_20153,N_19823,N_19879);
nand U20154 (N_20154,N_19943,N_19808);
xor U20155 (N_20155,N_19895,N_19781);
or U20156 (N_20156,N_19774,N_19939);
and U20157 (N_20157,N_19770,N_19956);
and U20158 (N_20158,N_19873,N_19812);
nor U20159 (N_20159,N_19801,N_19982);
xor U20160 (N_20160,N_19842,N_19956);
nor U20161 (N_20161,N_19958,N_19952);
nand U20162 (N_20162,N_19757,N_19810);
or U20163 (N_20163,N_19895,N_19815);
or U20164 (N_20164,N_19885,N_19940);
nor U20165 (N_20165,N_19778,N_19926);
nor U20166 (N_20166,N_19944,N_19952);
and U20167 (N_20167,N_19873,N_19885);
nor U20168 (N_20168,N_19793,N_19827);
and U20169 (N_20169,N_19988,N_19833);
nand U20170 (N_20170,N_19815,N_19983);
or U20171 (N_20171,N_19898,N_19767);
nand U20172 (N_20172,N_19856,N_19817);
or U20173 (N_20173,N_19901,N_19890);
and U20174 (N_20174,N_19884,N_19757);
xor U20175 (N_20175,N_19802,N_19919);
and U20176 (N_20176,N_19984,N_19947);
nand U20177 (N_20177,N_19831,N_19879);
xor U20178 (N_20178,N_19807,N_19952);
or U20179 (N_20179,N_19778,N_19875);
nand U20180 (N_20180,N_19965,N_19819);
or U20181 (N_20181,N_19823,N_19836);
nand U20182 (N_20182,N_19898,N_19999);
nor U20183 (N_20183,N_19807,N_19912);
nor U20184 (N_20184,N_19963,N_19982);
or U20185 (N_20185,N_19876,N_19768);
nand U20186 (N_20186,N_19876,N_19906);
xnor U20187 (N_20187,N_19844,N_19830);
xnor U20188 (N_20188,N_19817,N_19797);
xor U20189 (N_20189,N_19860,N_19929);
or U20190 (N_20190,N_19977,N_19952);
nand U20191 (N_20191,N_19970,N_19870);
or U20192 (N_20192,N_19777,N_19976);
xor U20193 (N_20193,N_19791,N_19816);
or U20194 (N_20194,N_19967,N_19791);
nor U20195 (N_20195,N_19949,N_19817);
nand U20196 (N_20196,N_19930,N_19818);
or U20197 (N_20197,N_19842,N_19886);
xnor U20198 (N_20198,N_19876,N_19964);
and U20199 (N_20199,N_19783,N_19791);
nor U20200 (N_20200,N_19769,N_19945);
nor U20201 (N_20201,N_19798,N_19934);
or U20202 (N_20202,N_19917,N_19859);
and U20203 (N_20203,N_19797,N_19923);
xnor U20204 (N_20204,N_19891,N_19761);
nand U20205 (N_20205,N_19902,N_19984);
nor U20206 (N_20206,N_19870,N_19930);
and U20207 (N_20207,N_19771,N_19932);
and U20208 (N_20208,N_19939,N_19836);
nor U20209 (N_20209,N_19814,N_19953);
nor U20210 (N_20210,N_19981,N_19934);
nor U20211 (N_20211,N_19963,N_19974);
nor U20212 (N_20212,N_19891,N_19854);
or U20213 (N_20213,N_19889,N_19972);
or U20214 (N_20214,N_19910,N_19821);
xor U20215 (N_20215,N_19894,N_19989);
xnor U20216 (N_20216,N_19890,N_19972);
nand U20217 (N_20217,N_19949,N_19947);
or U20218 (N_20218,N_19995,N_19951);
or U20219 (N_20219,N_19804,N_19877);
xnor U20220 (N_20220,N_19847,N_19862);
and U20221 (N_20221,N_19990,N_19915);
and U20222 (N_20222,N_19789,N_19855);
or U20223 (N_20223,N_19798,N_19988);
xor U20224 (N_20224,N_19965,N_19967);
nand U20225 (N_20225,N_19846,N_19929);
or U20226 (N_20226,N_19838,N_19866);
nor U20227 (N_20227,N_19843,N_19972);
nor U20228 (N_20228,N_19853,N_19887);
nor U20229 (N_20229,N_19833,N_19845);
and U20230 (N_20230,N_19884,N_19977);
or U20231 (N_20231,N_19807,N_19863);
xor U20232 (N_20232,N_19835,N_19899);
nand U20233 (N_20233,N_19881,N_19926);
or U20234 (N_20234,N_19859,N_19915);
and U20235 (N_20235,N_19869,N_19987);
xnor U20236 (N_20236,N_19902,N_19930);
and U20237 (N_20237,N_19889,N_19873);
and U20238 (N_20238,N_19785,N_19761);
and U20239 (N_20239,N_19798,N_19753);
nor U20240 (N_20240,N_19983,N_19852);
nor U20241 (N_20241,N_19750,N_19992);
or U20242 (N_20242,N_19987,N_19917);
nand U20243 (N_20243,N_19999,N_19907);
nor U20244 (N_20244,N_19934,N_19847);
or U20245 (N_20245,N_19960,N_19916);
and U20246 (N_20246,N_19779,N_19835);
or U20247 (N_20247,N_19846,N_19834);
nor U20248 (N_20248,N_19882,N_19917);
nor U20249 (N_20249,N_19880,N_19753);
or U20250 (N_20250,N_20078,N_20157);
nor U20251 (N_20251,N_20027,N_20053);
nor U20252 (N_20252,N_20141,N_20168);
xnor U20253 (N_20253,N_20148,N_20000);
nand U20254 (N_20254,N_20014,N_20108);
nor U20255 (N_20255,N_20020,N_20039);
xnor U20256 (N_20256,N_20209,N_20085);
or U20257 (N_20257,N_20084,N_20211);
nand U20258 (N_20258,N_20199,N_20128);
nand U20259 (N_20259,N_20190,N_20100);
xnor U20260 (N_20260,N_20069,N_20089);
nor U20261 (N_20261,N_20111,N_20215);
or U20262 (N_20262,N_20144,N_20042);
and U20263 (N_20263,N_20201,N_20193);
and U20264 (N_20264,N_20239,N_20140);
nor U20265 (N_20265,N_20101,N_20059);
and U20266 (N_20266,N_20159,N_20153);
nand U20267 (N_20267,N_20195,N_20230);
or U20268 (N_20268,N_20222,N_20246);
and U20269 (N_20269,N_20029,N_20189);
nor U20270 (N_20270,N_20238,N_20163);
nor U20271 (N_20271,N_20136,N_20207);
and U20272 (N_20272,N_20224,N_20142);
xor U20273 (N_20273,N_20156,N_20028);
xnor U20274 (N_20274,N_20048,N_20139);
and U20275 (N_20275,N_20040,N_20160);
xnor U20276 (N_20276,N_20013,N_20182);
and U20277 (N_20277,N_20206,N_20032);
and U20278 (N_20278,N_20158,N_20077);
nor U20279 (N_20279,N_20129,N_20073);
or U20280 (N_20280,N_20231,N_20060);
or U20281 (N_20281,N_20086,N_20093);
nor U20282 (N_20282,N_20019,N_20187);
nor U20283 (N_20283,N_20098,N_20102);
nor U20284 (N_20284,N_20165,N_20214);
nand U20285 (N_20285,N_20171,N_20050);
xnor U20286 (N_20286,N_20126,N_20143);
or U20287 (N_20287,N_20240,N_20072);
nand U20288 (N_20288,N_20055,N_20070);
xnor U20289 (N_20289,N_20200,N_20116);
xor U20290 (N_20290,N_20041,N_20067);
nand U20291 (N_20291,N_20091,N_20021);
xor U20292 (N_20292,N_20095,N_20226);
and U20293 (N_20293,N_20054,N_20058);
or U20294 (N_20294,N_20135,N_20012);
or U20295 (N_20295,N_20052,N_20096);
nand U20296 (N_20296,N_20161,N_20075);
nor U20297 (N_20297,N_20047,N_20225);
xor U20298 (N_20298,N_20104,N_20191);
or U20299 (N_20299,N_20249,N_20113);
xnor U20300 (N_20300,N_20074,N_20179);
or U20301 (N_20301,N_20245,N_20175);
nand U20302 (N_20302,N_20044,N_20205);
nor U20303 (N_20303,N_20026,N_20127);
xor U20304 (N_20304,N_20247,N_20164);
xnor U20305 (N_20305,N_20216,N_20004);
xnor U20306 (N_20306,N_20114,N_20071);
xnor U20307 (N_20307,N_20090,N_20131);
nor U20308 (N_20308,N_20137,N_20010);
nor U20309 (N_20309,N_20234,N_20066);
xnor U20310 (N_20310,N_20228,N_20123);
xnor U20311 (N_20311,N_20082,N_20197);
or U20312 (N_20312,N_20080,N_20018);
or U20313 (N_20313,N_20155,N_20223);
nand U20314 (N_20314,N_20196,N_20198);
xor U20315 (N_20315,N_20007,N_20138);
nand U20316 (N_20316,N_20130,N_20092);
and U20317 (N_20317,N_20051,N_20181);
xnor U20318 (N_20318,N_20124,N_20120);
or U20319 (N_20319,N_20030,N_20213);
nand U20320 (N_20320,N_20087,N_20049);
and U20321 (N_20321,N_20186,N_20210);
or U20322 (N_20322,N_20023,N_20045);
nor U20323 (N_20323,N_20167,N_20194);
nor U20324 (N_20324,N_20169,N_20064);
nor U20325 (N_20325,N_20003,N_20125);
nand U20326 (N_20326,N_20202,N_20145);
xor U20327 (N_20327,N_20097,N_20243);
nand U20328 (N_20328,N_20149,N_20033);
nand U20329 (N_20329,N_20152,N_20173);
xnor U20330 (N_20330,N_20036,N_20043);
xnor U20331 (N_20331,N_20134,N_20218);
nand U20332 (N_20332,N_20133,N_20180);
or U20333 (N_20333,N_20094,N_20068);
nand U20334 (N_20334,N_20248,N_20110);
nor U20335 (N_20335,N_20016,N_20154);
or U20336 (N_20336,N_20132,N_20022);
and U20337 (N_20337,N_20237,N_20172);
nand U20338 (N_20338,N_20221,N_20117);
or U20339 (N_20339,N_20217,N_20122);
and U20340 (N_20340,N_20121,N_20235);
or U20341 (N_20341,N_20185,N_20170);
and U20342 (N_20342,N_20119,N_20015);
xnor U20343 (N_20343,N_20046,N_20001);
and U20344 (N_20344,N_20166,N_20035);
and U20345 (N_20345,N_20109,N_20037);
xor U20346 (N_20346,N_20146,N_20083);
nand U20347 (N_20347,N_20203,N_20088);
nand U20348 (N_20348,N_20034,N_20229);
and U20349 (N_20349,N_20236,N_20204);
nor U20350 (N_20350,N_20174,N_20184);
and U20351 (N_20351,N_20147,N_20233);
nor U20352 (N_20352,N_20057,N_20025);
nor U20353 (N_20353,N_20038,N_20227);
or U20354 (N_20354,N_20188,N_20009);
xnor U20355 (N_20355,N_20005,N_20112);
nand U20356 (N_20356,N_20232,N_20212);
xnor U20357 (N_20357,N_20031,N_20061);
nand U20358 (N_20358,N_20002,N_20178);
and U20359 (N_20359,N_20244,N_20062);
xnor U20360 (N_20360,N_20079,N_20150);
or U20361 (N_20361,N_20220,N_20076);
xor U20362 (N_20362,N_20105,N_20017);
nor U20363 (N_20363,N_20099,N_20006);
nand U20364 (N_20364,N_20103,N_20192);
or U20365 (N_20365,N_20063,N_20115);
or U20366 (N_20366,N_20118,N_20177);
and U20367 (N_20367,N_20162,N_20008);
xnor U20368 (N_20368,N_20208,N_20011);
or U20369 (N_20369,N_20219,N_20081);
or U20370 (N_20370,N_20024,N_20183);
xnor U20371 (N_20371,N_20056,N_20241);
xor U20372 (N_20372,N_20242,N_20151);
nand U20373 (N_20373,N_20107,N_20065);
and U20374 (N_20374,N_20176,N_20106);
xor U20375 (N_20375,N_20032,N_20127);
or U20376 (N_20376,N_20056,N_20211);
xnor U20377 (N_20377,N_20018,N_20168);
nor U20378 (N_20378,N_20067,N_20163);
nor U20379 (N_20379,N_20135,N_20165);
nor U20380 (N_20380,N_20144,N_20098);
or U20381 (N_20381,N_20087,N_20240);
or U20382 (N_20382,N_20005,N_20155);
and U20383 (N_20383,N_20161,N_20157);
nand U20384 (N_20384,N_20148,N_20116);
or U20385 (N_20385,N_20182,N_20110);
nor U20386 (N_20386,N_20035,N_20161);
or U20387 (N_20387,N_20064,N_20018);
xnor U20388 (N_20388,N_20074,N_20198);
and U20389 (N_20389,N_20158,N_20197);
nand U20390 (N_20390,N_20089,N_20054);
and U20391 (N_20391,N_20222,N_20075);
nor U20392 (N_20392,N_20144,N_20134);
or U20393 (N_20393,N_20139,N_20076);
and U20394 (N_20394,N_20045,N_20089);
nor U20395 (N_20395,N_20212,N_20143);
nand U20396 (N_20396,N_20231,N_20036);
and U20397 (N_20397,N_20217,N_20213);
and U20398 (N_20398,N_20188,N_20210);
xnor U20399 (N_20399,N_20109,N_20082);
nor U20400 (N_20400,N_20235,N_20247);
and U20401 (N_20401,N_20237,N_20046);
and U20402 (N_20402,N_20190,N_20050);
nor U20403 (N_20403,N_20233,N_20070);
and U20404 (N_20404,N_20127,N_20090);
nor U20405 (N_20405,N_20025,N_20079);
xor U20406 (N_20406,N_20132,N_20236);
and U20407 (N_20407,N_20016,N_20196);
or U20408 (N_20408,N_20217,N_20220);
nor U20409 (N_20409,N_20191,N_20220);
and U20410 (N_20410,N_20236,N_20111);
nor U20411 (N_20411,N_20198,N_20112);
and U20412 (N_20412,N_20111,N_20155);
xnor U20413 (N_20413,N_20234,N_20049);
nor U20414 (N_20414,N_20018,N_20175);
or U20415 (N_20415,N_20019,N_20159);
nand U20416 (N_20416,N_20000,N_20232);
nor U20417 (N_20417,N_20096,N_20079);
and U20418 (N_20418,N_20233,N_20218);
or U20419 (N_20419,N_20243,N_20217);
or U20420 (N_20420,N_20217,N_20008);
nor U20421 (N_20421,N_20166,N_20165);
or U20422 (N_20422,N_20165,N_20134);
nor U20423 (N_20423,N_20222,N_20239);
and U20424 (N_20424,N_20010,N_20145);
and U20425 (N_20425,N_20180,N_20185);
or U20426 (N_20426,N_20000,N_20036);
nor U20427 (N_20427,N_20066,N_20043);
nand U20428 (N_20428,N_20047,N_20203);
nand U20429 (N_20429,N_20153,N_20076);
nand U20430 (N_20430,N_20204,N_20068);
and U20431 (N_20431,N_20120,N_20143);
xor U20432 (N_20432,N_20139,N_20023);
nand U20433 (N_20433,N_20054,N_20159);
and U20434 (N_20434,N_20074,N_20170);
and U20435 (N_20435,N_20118,N_20077);
or U20436 (N_20436,N_20049,N_20162);
xor U20437 (N_20437,N_20027,N_20141);
nand U20438 (N_20438,N_20204,N_20126);
or U20439 (N_20439,N_20197,N_20059);
xnor U20440 (N_20440,N_20029,N_20172);
or U20441 (N_20441,N_20068,N_20072);
nand U20442 (N_20442,N_20214,N_20126);
nor U20443 (N_20443,N_20117,N_20206);
or U20444 (N_20444,N_20222,N_20004);
or U20445 (N_20445,N_20059,N_20135);
or U20446 (N_20446,N_20081,N_20246);
nand U20447 (N_20447,N_20163,N_20173);
or U20448 (N_20448,N_20154,N_20097);
xnor U20449 (N_20449,N_20238,N_20184);
xnor U20450 (N_20450,N_20234,N_20231);
nand U20451 (N_20451,N_20187,N_20240);
and U20452 (N_20452,N_20129,N_20009);
xor U20453 (N_20453,N_20020,N_20074);
nand U20454 (N_20454,N_20052,N_20024);
and U20455 (N_20455,N_20046,N_20222);
and U20456 (N_20456,N_20242,N_20128);
xnor U20457 (N_20457,N_20211,N_20198);
xor U20458 (N_20458,N_20074,N_20132);
nand U20459 (N_20459,N_20242,N_20166);
and U20460 (N_20460,N_20216,N_20044);
nand U20461 (N_20461,N_20117,N_20007);
or U20462 (N_20462,N_20242,N_20150);
or U20463 (N_20463,N_20245,N_20064);
nand U20464 (N_20464,N_20087,N_20027);
xnor U20465 (N_20465,N_20077,N_20105);
and U20466 (N_20466,N_20241,N_20208);
nand U20467 (N_20467,N_20045,N_20189);
nand U20468 (N_20468,N_20062,N_20057);
nand U20469 (N_20469,N_20207,N_20081);
and U20470 (N_20470,N_20108,N_20122);
nor U20471 (N_20471,N_20169,N_20053);
nand U20472 (N_20472,N_20138,N_20008);
or U20473 (N_20473,N_20144,N_20226);
or U20474 (N_20474,N_20212,N_20199);
nand U20475 (N_20475,N_20008,N_20204);
nand U20476 (N_20476,N_20118,N_20005);
or U20477 (N_20477,N_20014,N_20207);
nor U20478 (N_20478,N_20134,N_20059);
and U20479 (N_20479,N_20011,N_20116);
xor U20480 (N_20480,N_20080,N_20017);
or U20481 (N_20481,N_20203,N_20232);
and U20482 (N_20482,N_20087,N_20075);
nor U20483 (N_20483,N_20212,N_20229);
and U20484 (N_20484,N_20156,N_20232);
nor U20485 (N_20485,N_20008,N_20029);
nor U20486 (N_20486,N_20246,N_20103);
nor U20487 (N_20487,N_20188,N_20137);
xor U20488 (N_20488,N_20132,N_20247);
nand U20489 (N_20489,N_20242,N_20210);
or U20490 (N_20490,N_20185,N_20013);
xnor U20491 (N_20491,N_20232,N_20074);
and U20492 (N_20492,N_20149,N_20197);
nor U20493 (N_20493,N_20246,N_20086);
and U20494 (N_20494,N_20014,N_20174);
and U20495 (N_20495,N_20244,N_20084);
nor U20496 (N_20496,N_20247,N_20234);
and U20497 (N_20497,N_20062,N_20031);
xor U20498 (N_20498,N_20169,N_20174);
xor U20499 (N_20499,N_20143,N_20152);
and U20500 (N_20500,N_20370,N_20479);
and U20501 (N_20501,N_20346,N_20389);
xnor U20502 (N_20502,N_20365,N_20472);
nand U20503 (N_20503,N_20279,N_20448);
xnor U20504 (N_20504,N_20436,N_20481);
xnor U20505 (N_20505,N_20492,N_20494);
nor U20506 (N_20506,N_20312,N_20344);
nand U20507 (N_20507,N_20496,N_20313);
xor U20508 (N_20508,N_20273,N_20367);
nor U20509 (N_20509,N_20468,N_20422);
xnor U20510 (N_20510,N_20420,N_20270);
xor U20511 (N_20511,N_20388,N_20325);
nor U20512 (N_20512,N_20363,N_20462);
and U20513 (N_20513,N_20441,N_20339);
xnor U20514 (N_20514,N_20392,N_20444);
nor U20515 (N_20515,N_20294,N_20330);
or U20516 (N_20516,N_20317,N_20401);
xnor U20517 (N_20517,N_20394,N_20355);
nor U20518 (N_20518,N_20275,N_20461);
and U20519 (N_20519,N_20369,N_20309);
nand U20520 (N_20520,N_20433,N_20299);
and U20521 (N_20521,N_20284,N_20482);
xnor U20522 (N_20522,N_20332,N_20435);
or U20523 (N_20523,N_20470,N_20424);
or U20524 (N_20524,N_20359,N_20301);
nand U20525 (N_20525,N_20447,N_20261);
and U20526 (N_20526,N_20327,N_20368);
and U20527 (N_20527,N_20310,N_20253);
nor U20528 (N_20528,N_20465,N_20374);
and U20529 (N_20529,N_20265,N_20425);
or U20530 (N_20530,N_20329,N_20377);
or U20531 (N_20531,N_20256,N_20338);
nand U20532 (N_20532,N_20259,N_20410);
and U20533 (N_20533,N_20271,N_20251);
nand U20534 (N_20534,N_20458,N_20356);
nor U20535 (N_20535,N_20416,N_20297);
or U20536 (N_20536,N_20342,N_20417);
or U20537 (N_20537,N_20335,N_20407);
nand U20538 (N_20538,N_20391,N_20408);
or U20539 (N_20539,N_20395,N_20292);
or U20540 (N_20540,N_20280,N_20400);
xor U20541 (N_20541,N_20489,N_20283);
or U20542 (N_20542,N_20498,N_20455);
or U20543 (N_20543,N_20304,N_20266);
nor U20544 (N_20544,N_20362,N_20257);
nor U20545 (N_20545,N_20398,N_20495);
or U20546 (N_20546,N_20477,N_20252);
or U20547 (N_20547,N_20484,N_20296);
and U20548 (N_20548,N_20318,N_20291);
xnor U20549 (N_20549,N_20396,N_20382);
nor U20550 (N_20550,N_20315,N_20326);
and U20551 (N_20551,N_20471,N_20314);
or U20552 (N_20552,N_20255,N_20258);
or U20553 (N_20553,N_20399,N_20403);
xor U20554 (N_20554,N_20336,N_20286);
xnor U20555 (N_20555,N_20405,N_20464);
or U20556 (N_20556,N_20449,N_20290);
nor U20557 (N_20557,N_20460,N_20347);
xnor U20558 (N_20558,N_20493,N_20285);
nor U20559 (N_20559,N_20340,N_20282);
nand U20560 (N_20560,N_20466,N_20307);
nor U20561 (N_20561,N_20413,N_20386);
and U20562 (N_20562,N_20333,N_20421);
xor U20563 (N_20563,N_20406,N_20260);
or U20564 (N_20564,N_20473,N_20404);
nand U20565 (N_20565,N_20293,N_20295);
or U20566 (N_20566,N_20381,N_20486);
nor U20567 (N_20567,N_20323,N_20480);
nor U20568 (N_20568,N_20298,N_20281);
xnor U20569 (N_20569,N_20430,N_20402);
nand U20570 (N_20570,N_20263,N_20262);
xor U20571 (N_20571,N_20278,N_20491);
xnor U20572 (N_20572,N_20384,N_20319);
xnor U20573 (N_20573,N_20437,N_20305);
nand U20574 (N_20574,N_20350,N_20415);
nor U20575 (N_20575,N_20328,N_20453);
nor U20576 (N_20576,N_20419,N_20373);
nor U20577 (N_20577,N_20276,N_20360);
or U20578 (N_20578,N_20375,N_20300);
or U20579 (N_20579,N_20371,N_20354);
nand U20580 (N_20580,N_20287,N_20478);
nand U20581 (N_20581,N_20390,N_20322);
xnor U20582 (N_20582,N_20269,N_20272);
nor U20583 (N_20583,N_20485,N_20467);
and U20584 (N_20584,N_20316,N_20418);
nor U20585 (N_20585,N_20277,N_20475);
xor U20586 (N_20586,N_20358,N_20412);
xnor U20587 (N_20587,N_20311,N_20443);
or U20588 (N_20588,N_20457,N_20331);
and U20589 (N_20589,N_20353,N_20343);
or U20590 (N_20590,N_20387,N_20483);
nor U20591 (N_20591,N_20463,N_20450);
and U20592 (N_20592,N_20308,N_20426);
and U20593 (N_20593,N_20439,N_20324);
and U20594 (N_20594,N_20454,N_20288);
nand U20595 (N_20595,N_20379,N_20372);
nand U20596 (N_20596,N_20334,N_20351);
nor U20597 (N_20597,N_20445,N_20497);
nand U20598 (N_20598,N_20431,N_20499);
nor U20599 (N_20599,N_20254,N_20423);
nor U20600 (N_20600,N_20432,N_20303);
nor U20601 (N_20601,N_20469,N_20440);
nand U20602 (N_20602,N_20456,N_20459);
and U20603 (N_20603,N_20352,N_20434);
nand U20604 (N_20604,N_20438,N_20345);
xnor U20605 (N_20605,N_20306,N_20302);
or U20606 (N_20606,N_20385,N_20361);
nand U20607 (N_20607,N_20268,N_20264);
or U20608 (N_20608,N_20274,N_20474);
nand U20609 (N_20609,N_20348,N_20488);
or U20610 (N_20610,N_20366,N_20250);
or U20611 (N_20611,N_20341,N_20349);
xnor U20612 (N_20612,N_20451,N_20321);
or U20613 (N_20613,N_20393,N_20409);
or U20614 (N_20614,N_20487,N_20383);
nor U20615 (N_20615,N_20442,N_20411);
nand U20616 (N_20616,N_20428,N_20357);
nand U20617 (N_20617,N_20427,N_20378);
or U20618 (N_20618,N_20289,N_20490);
nor U20619 (N_20619,N_20446,N_20397);
xor U20620 (N_20620,N_20376,N_20337);
nor U20621 (N_20621,N_20267,N_20380);
or U20622 (N_20622,N_20429,N_20476);
and U20623 (N_20623,N_20452,N_20364);
nor U20624 (N_20624,N_20414,N_20320);
and U20625 (N_20625,N_20289,N_20255);
nand U20626 (N_20626,N_20385,N_20439);
xor U20627 (N_20627,N_20402,N_20475);
and U20628 (N_20628,N_20497,N_20309);
nand U20629 (N_20629,N_20440,N_20273);
or U20630 (N_20630,N_20256,N_20368);
or U20631 (N_20631,N_20264,N_20289);
nand U20632 (N_20632,N_20495,N_20493);
or U20633 (N_20633,N_20412,N_20438);
xnor U20634 (N_20634,N_20318,N_20316);
and U20635 (N_20635,N_20485,N_20438);
xnor U20636 (N_20636,N_20376,N_20492);
or U20637 (N_20637,N_20374,N_20337);
nand U20638 (N_20638,N_20336,N_20477);
or U20639 (N_20639,N_20291,N_20273);
nor U20640 (N_20640,N_20372,N_20416);
or U20641 (N_20641,N_20474,N_20412);
or U20642 (N_20642,N_20289,N_20405);
nand U20643 (N_20643,N_20278,N_20391);
or U20644 (N_20644,N_20413,N_20473);
or U20645 (N_20645,N_20272,N_20323);
or U20646 (N_20646,N_20332,N_20484);
or U20647 (N_20647,N_20422,N_20272);
and U20648 (N_20648,N_20441,N_20364);
xnor U20649 (N_20649,N_20279,N_20263);
nor U20650 (N_20650,N_20496,N_20426);
xor U20651 (N_20651,N_20262,N_20374);
nor U20652 (N_20652,N_20356,N_20360);
or U20653 (N_20653,N_20348,N_20474);
and U20654 (N_20654,N_20389,N_20403);
or U20655 (N_20655,N_20406,N_20307);
xnor U20656 (N_20656,N_20374,N_20338);
xor U20657 (N_20657,N_20417,N_20374);
xnor U20658 (N_20658,N_20270,N_20278);
nand U20659 (N_20659,N_20365,N_20272);
xor U20660 (N_20660,N_20355,N_20250);
and U20661 (N_20661,N_20426,N_20402);
nand U20662 (N_20662,N_20353,N_20424);
nor U20663 (N_20663,N_20467,N_20301);
nand U20664 (N_20664,N_20268,N_20343);
and U20665 (N_20665,N_20319,N_20373);
xor U20666 (N_20666,N_20308,N_20452);
or U20667 (N_20667,N_20251,N_20359);
nand U20668 (N_20668,N_20281,N_20484);
nand U20669 (N_20669,N_20316,N_20257);
or U20670 (N_20670,N_20441,N_20289);
nor U20671 (N_20671,N_20438,N_20437);
nand U20672 (N_20672,N_20410,N_20464);
xor U20673 (N_20673,N_20404,N_20256);
and U20674 (N_20674,N_20319,N_20437);
nand U20675 (N_20675,N_20469,N_20493);
or U20676 (N_20676,N_20465,N_20360);
nor U20677 (N_20677,N_20472,N_20462);
nand U20678 (N_20678,N_20331,N_20444);
or U20679 (N_20679,N_20474,N_20289);
nand U20680 (N_20680,N_20350,N_20465);
xor U20681 (N_20681,N_20495,N_20261);
xor U20682 (N_20682,N_20450,N_20461);
nand U20683 (N_20683,N_20480,N_20413);
nor U20684 (N_20684,N_20444,N_20277);
or U20685 (N_20685,N_20274,N_20280);
nand U20686 (N_20686,N_20300,N_20327);
and U20687 (N_20687,N_20448,N_20468);
nand U20688 (N_20688,N_20253,N_20269);
or U20689 (N_20689,N_20394,N_20331);
nand U20690 (N_20690,N_20279,N_20438);
xor U20691 (N_20691,N_20334,N_20458);
and U20692 (N_20692,N_20299,N_20261);
nand U20693 (N_20693,N_20464,N_20399);
or U20694 (N_20694,N_20368,N_20291);
or U20695 (N_20695,N_20493,N_20435);
and U20696 (N_20696,N_20450,N_20257);
xor U20697 (N_20697,N_20411,N_20374);
nand U20698 (N_20698,N_20332,N_20426);
and U20699 (N_20699,N_20271,N_20280);
nor U20700 (N_20700,N_20314,N_20278);
xor U20701 (N_20701,N_20479,N_20492);
xnor U20702 (N_20702,N_20385,N_20457);
and U20703 (N_20703,N_20421,N_20281);
nor U20704 (N_20704,N_20477,N_20368);
and U20705 (N_20705,N_20458,N_20449);
or U20706 (N_20706,N_20452,N_20365);
xnor U20707 (N_20707,N_20406,N_20280);
nand U20708 (N_20708,N_20498,N_20264);
and U20709 (N_20709,N_20409,N_20436);
and U20710 (N_20710,N_20484,N_20433);
nor U20711 (N_20711,N_20314,N_20434);
and U20712 (N_20712,N_20418,N_20498);
nand U20713 (N_20713,N_20359,N_20429);
xor U20714 (N_20714,N_20352,N_20435);
xor U20715 (N_20715,N_20270,N_20467);
nor U20716 (N_20716,N_20493,N_20444);
nor U20717 (N_20717,N_20374,N_20364);
nand U20718 (N_20718,N_20283,N_20439);
xnor U20719 (N_20719,N_20255,N_20423);
nor U20720 (N_20720,N_20422,N_20348);
xnor U20721 (N_20721,N_20306,N_20396);
xor U20722 (N_20722,N_20321,N_20253);
xor U20723 (N_20723,N_20498,N_20312);
xnor U20724 (N_20724,N_20380,N_20296);
or U20725 (N_20725,N_20423,N_20469);
nand U20726 (N_20726,N_20256,N_20495);
or U20727 (N_20727,N_20456,N_20373);
xnor U20728 (N_20728,N_20457,N_20466);
and U20729 (N_20729,N_20334,N_20255);
and U20730 (N_20730,N_20446,N_20407);
or U20731 (N_20731,N_20410,N_20401);
nand U20732 (N_20732,N_20385,N_20440);
and U20733 (N_20733,N_20456,N_20425);
nor U20734 (N_20734,N_20398,N_20354);
and U20735 (N_20735,N_20257,N_20353);
or U20736 (N_20736,N_20435,N_20489);
or U20737 (N_20737,N_20341,N_20284);
nor U20738 (N_20738,N_20491,N_20326);
or U20739 (N_20739,N_20441,N_20287);
nor U20740 (N_20740,N_20380,N_20375);
nor U20741 (N_20741,N_20367,N_20490);
and U20742 (N_20742,N_20309,N_20410);
or U20743 (N_20743,N_20310,N_20254);
nand U20744 (N_20744,N_20344,N_20265);
xnor U20745 (N_20745,N_20483,N_20339);
xor U20746 (N_20746,N_20362,N_20332);
and U20747 (N_20747,N_20415,N_20400);
nor U20748 (N_20748,N_20447,N_20457);
nand U20749 (N_20749,N_20404,N_20494);
and U20750 (N_20750,N_20613,N_20540);
and U20751 (N_20751,N_20504,N_20621);
nand U20752 (N_20752,N_20618,N_20671);
or U20753 (N_20753,N_20636,N_20538);
nand U20754 (N_20754,N_20701,N_20668);
and U20755 (N_20755,N_20608,N_20650);
and U20756 (N_20756,N_20694,N_20577);
xnor U20757 (N_20757,N_20583,N_20556);
nand U20758 (N_20758,N_20574,N_20705);
nand U20759 (N_20759,N_20676,N_20601);
or U20760 (N_20760,N_20579,N_20689);
or U20761 (N_20761,N_20539,N_20542);
nor U20762 (N_20762,N_20634,N_20731);
or U20763 (N_20763,N_20728,N_20506);
or U20764 (N_20764,N_20704,N_20647);
and U20765 (N_20765,N_20683,N_20652);
nor U20766 (N_20766,N_20727,N_20721);
nor U20767 (N_20767,N_20588,N_20596);
or U20768 (N_20768,N_20706,N_20546);
or U20769 (N_20769,N_20663,N_20559);
nor U20770 (N_20770,N_20557,N_20572);
xnor U20771 (N_20771,N_20606,N_20598);
nor U20772 (N_20772,N_20656,N_20635);
or U20773 (N_20773,N_20669,N_20664);
and U20774 (N_20774,N_20591,N_20628);
nand U20775 (N_20775,N_20695,N_20672);
xor U20776 (N_20776,N_20551,N_20512);
nor U20777 (N_20777,N_20584,N_20600);
and U20778 (N_20778,N_20673,N_20674);
nor U20779 (N_20779,N_20722,N_20702);
nand U20780 (N_20780,N_20605,N_20681);
nand U20781 (N_20781,N_20528,N_20544);
or U20782 (N_20782,N_20717,N_20505);
nand U20783 (N_20783,N_20723,N_20675);
xor U20784 (N_20784,N_20517,N_20678);
and U20785 (N_20785,N_20644,N_20500);
nand U20786 (N_20786,N_20633,N_20548);
nor U20787 (N_20787,N_20733,N_20665);
nand U20788 (N_20788,N_20744,N_20549);
and U20789 (N_20789,N_20724,N_20738);
nor U20790 (N_20790,N_20575,N_20726);
xnor U20791 (N_20791,N_20629,N_20554);
or U20792 (N_20792,N_20576,N_20643);
or U20793 (N_20793,N_20581,N_20501);
nor U20794 (N_20794,N_20642,N_20699);
or U20795 (N_20795,N_20626,N_20565);
xor U20796 (N_20796,N_20735,N_20516);
nor U20797 (N_20797,N_20612,N_20703);
nor U20798 (N_20798,N_20578,N_20742);
xnor U20799 (N_20799,N_20533,N_20631);
xor U20800 (N_20800,N_20594,N_20716);
and U20801 (N_20801,N_20707,N_20573);
or U20802 (N_20802,N_20570,N_20743);
nand U20803 (N_20803,N_20590,N_20566);
nor U20804 (N_20804,N_20649,N_20526);
xor U20805 (N_20805,N_20611,N_20525);
nor U20806 (N_20806,N_20585,N_20690);
and U20807 (N_20807,N_20550,N_20749);
or U20808 (N_20808,N_20713,N_20688);
nor U20809 (N_20809,N_20641,N_20560);
nand U20810 (N_20810,N_20691,N_20615);
nand U20811 (N_20811,N_20680,N_20521);
xor U20812 (N_20812,N_20655,N_20592);
xor U20813 (N_20813,N_20604,N_20527);
or U20814 (N_20814,N_20692,N_20684);
xnor U20815 (N_20815,N_20593,N_20696);
or U20816 (N_20816,N_20536,N_20561);
xor U20817 (N_20817,N_20700,N_20653);
nor U20818 (N_20818,N_20730,N_20514);
nand U20819 (N_20819,N_20646,N_20503);
and U20820 (N_20820,N_20741,N_20509);
nor U20821 (N_20821,N_20622,N_20718);
or U20822 (N_20822,N_20543,N_20555);
xnor U20823 (N_20823,N_20545,N_20511);
or U20824 (N_20824,N_20697,N_20745);
nor U20825 (N_20825,N_20639,N_20589);
nor U20826 (N_20826,N_20667,N_20637);
nor U20827 (N_20827,N_20685,N_20710);
or U20828 (N_20828,N_20571,N_20720);
xnor U20829 (N_20829,N_20616,N_20693);
and U20830 (N_20830,N_20739,N_20518);
or U20831 (N_20831,N_20587,N_20607);
nor U20832 (N_20832,N_20719,N_20619);
nor U20833 (N_20833,N_20623,N_20659);
or U20834 (N_20834,N_20537,N_20507);
xor U20835 (N_20835,N_20638,N_20709);
and U20836 (N_20836,N_20515,N_20597);
nand U20837 (N_20837,N_20564,N_20679);
xor U20838 (N_20838,N_20519,N_20715);
xor U20839 (N_20839,N_20534,N_20531);
nand U20840 (N_20840,N_20582,N_20603);
and U20841 (N_20841,N_20734,N_20662);
nor U20842 (N_20842,N_20620,N_20609);
or U20843 (N_20843,N_20670,N_20625);
nand U20844 (N_20844,N_20522,N_20599);
xnor U20845 (N_20845,N_20740,N_20748);
and U20846 (N_20846,N_20654,N_20558);
or U20847 (N_20847,N_20529,N_20586);
and U20848 (N_20848,N_20523,N_20712);
or U20849 (N_20849,N_20502,N_20640);
or U20850 (N_20850,N_20714,N_20563);
or U20851 (N_20851,N_20732,N_20666);
nor U20852 (N_20852,N_20682,N_20569);
nor U20853 (N_20853,N_20708,N_20510);
nand U20854 (N_20854,N_20645,N_20541);
nand U20855 (N_20855,N_20630,N_20725);
or U20856 (N_20856,N_20627,N_20698);
xnor U20857 (N_20857,N_20736,N_20513);
nand U20858 (N_20858,N_20562,N_20677);
or U20859 (N_20859,N_20520,N_20660);
and U20860 (N_20860,N_20610,N_20651);
nor U20861 (N_20861,N_20648,N_20624);
xor U20862 (N_20862,N_20729,N_20746);
or U20863 (N_20863,N_20535,N_20595);
xor U20864 (N_20864,N_20532,N_20687);
xnor U20865 (N_20865,N_20524,N_20530);
nor U20866 (N_20866,N_20617,N_20657);
and U20867 (N_20867,N_20553,N_20737);
or U20868 (N_20868,N_20632,N_20508);
and U20869 (N_20869,N_20614,N_20552);
and U20870 (N_20870,N_20686,N_20658);
nand U20871 (N_20871,N_20547,N_20602);
or U20872 (N_20872,N_20711,N_20567);
nand U20873 (N_20873,N_20661,N_20747);
and U20874 (N_20874,N_20568,N_20580);
xnor U20875 (N_20875,N_20503,N_20642);
and U20876 (N_20876,N_20665,N_20584);
nor U20877 (N_20877,N_20624,N_20665);
nand U20878 (N_20878,N_20598,N_20682);
and U20879 (N_20879,N_20588,N_20611);
nand U20880 (N_20880,N_20724,N_20525);
xnor U20881 (N_20881,N_20536,N_20560);
xnor U20882 (N_20882,N_20624,N_20592);
xnor U20883 (N_20883,N_20580,N_20625);
nor U20884 (N_20884,N_20532,N_20738);
and U20885 (N_20885,N_20528,N_20504);
xor U20886 (N_20886,N_20646,N_20687);
nand U20887 (N_20887,N_20720,N_20652);
and U20888 (N_20888,N_20574,N_20696);
nand U20889 (N_20889,N_20648,N_20629);
nor U20890 (N_20890,N_20618,N_20611);
xor U20891 (N_20891,N_20726,N_20703);
nand U20892 (N_20892,N_20663,N_20650);
xnor U20893 (N_20893,N_20738,N_20745);
or U20894 (N_20894,N_20704,N_20562);
or U20895 (N_20895,N_20720,N_20527);
and U20896 (N_20896,N_20567,N_20577);
and U20897 (N_20897,N_20630,N_20577);
or U20898 (N_20898,N_20546,N_20580);
and U20899 (N_20899,N_20665,N_20521);
nand U20900 (N_20900,N_20579,N_20568);
nand U20901 (N_20901,N_20519,N_20739);
nand U20902 (N_20902,N_20574,N_20634);
and U20903 (N_20903,N_20728,N_20658);
xnor U20904 (N_20904,N_20510,N_20501);
nor U20905 (N_20905,N_20657,N_20573);
xnor U20906 (N_20906,N_20575,N_20580);
and U20907 (N_20907,N_20710,N_20728);
or U20908 (N_20908,N_20566,N_20592);
xor U20909 (N_20909,N_20530,N_20699);
nand U20910 (N_20910,N_20609,N_20731);
and U20911 (N_20911,N_20501,N_20543);
nand U20912 (N_20912,N_20546,N_20711);
nand U20913 (N_20913,N_20674,N_20517);
or U20914 (N_20914,N_20696,N_20737);
nand U20915 (N_20915,N_20726,N_20543);
or U20916 (N_20916,N_20510,N_20609);
xor U20917 (N_20917,N_20588,N_20648);
or U20918 (N_20918,N_20510,N_20575);
and U20919 (N_20919,N_20560,N_20581);
nand U20920 (N_20920,N_20536,N_20601);
nand U20921 (N_20921,N_20537,N_20595);
xor U20922 (N_20922,N_20739,N_20517);
nor U20923 (N_20923,N_20561,N_20683);
or U20924 (N_20924,N_20564,N_20587);
or U20925 (N_20925,N_20551,N_20574);
nor U20926 (N_20926,N_20578,N_20731);
nor U20927 (N_20927,N_20517,N_20566);
or U20928 (N_20928,N_20667,N_20734);
nand U20929 (N_20929,N_20686,N_20583);
nand U20930 (N_20930,N_20693,N_20503);
or U20931 (N_20931,N_20666,N_20596);
and U20932 (N_20932,N_20604,N_20658);
or U20933 (N_20933,N_20647,N_20748);
or U20934 (N_20934,N_20717,N_20598);
xor U20935 (N_20935,N_20558,N_20660);
nand U20936 (N_20936,N_20556,N_20508);
nand U20937 (N_20937,N_20610,N_20655);
nor U20938 (N_20938,N_20524,N_20620);
nand U20939 (N_20939,N_20518,N_20663);
and U20940 (N_20940,N_20536,N_20656);
and U20941 (N_20941,N_20749,N_20593);
or U20942 (N_20942,N_20713,N_20728);
nor U20943 (N_20943,N_20611,N_20661);
xor U20944 (N_20944,N_20663,N_20516);
nor U20945 (N_20945,N_20689,N_20742);
and U20946 (N_20946,N_20578,N_20705);
nor U20947 (N_20947,N_20742,N_20609);
nand U20948 (N_20948,N_20663,N_20645);
nor U20949 (N_20949,N_20574,N_20685);
nor U20950 (N_20950,N_20598,N_20583);
nand U20951 (N_20951,N_20743,N_20541);
nor U20952 (N_20952,N_20735,N_20554);
or U20953 (N_20953,N_20693,N_20537);
nor U20954 (N_20954,N_20568,N_20644);
nand U20955 (N_20955,N_20670,N_20668);
and U20956 (N_20956,N_20571,N_20697);
or U20957 (N_20957,N_20526,N_20572);
nand U20958 (N_20958,N_20569,N_20652);
and U20959 (N_20959,N_20588,N_20727);
xor U20960 (N_20960,N_20691,N_20689);
and U20961 (N_20961,N_20645,N_20534);
and U20962 (N_20962,N_20682,N_20587);
nand U20963 (N_20963,N_20589,N_20648);
or U20964 (N_20964,N_20605,N_20572);
nor U20965 (N_20965,N_20695,N_20680);
xnor U20966 (N_20966,N_20645,N_20512);
nand U20967 (N_20967,N_20640,N_20662);
nand U20968 (N_20968,N_20557,N_20669);
or U20969 (N_20969,N_20622,N_20703);
or U20970 (N_20970,N_20576,N_20612);
and U20971 (N_20971,N_20638,N_20642);
xnor U20972 (N_20972,N_20687,N_20679);
xnor U20973 (N_20973,N_20605,N_20571);
nor U20974 (N_20974,N_20582,N_20554);
or U20975 (N_20975,N_20669,N_20749);
nand U20976 (N_20976,N_20703,N_20519);
and U20977 (N_20977,N_20539,N_20597);
xnor U20978 (N_20978,N_20587,N_20716);
nand U20979 (N_20979,N_20708,N_20736);
and U20980 (N_20980,N_20690,N_20596);
or U20981 (N_20981,N_20737,N_20687);
nand U20982 (N_20982,N_20623,N_20622);
nand U20983 (N_20983,N_20577,N_20655);
and U20984 (N_20984,N_20670,N_20532);
or U20985 (N_20985,N_20690,N_20675);
or U20986 (N_20986,N_20691,N_20709);
or U20987 (N_20987,N_20577,N_20668);
xor U20988 (N_20988,N_20616,N_20700);
or U20989 (N_20989,N_20623,N_20553);
and U20990 (N_20990,N_20652,N_20621);
nor U20991 (N_20991,N_20632,N_20672);
nand U20992 (N_20992,N_20600,N_20519);
nand U20993 (N_20993,N_20678,N_20520);
nand U20994 (N_20994,N_20650,N_20569);
nand U20995 (N_20995,N_20644,N_20705);
or U20996 (N_20996,N_20593,N_20539);
or U20997 (N_20997,N_20672,N_20525);
xor U20998 (N_20998,N_20727,N_20505);
nand U20999 (N_20999,N_20618,N_20621);
nor U21000 (N_21000,N_20952,N_20950);
nand U21001 (N_21001,N_20764,N_20752);
xor U21002 (N_21002,N_20848,N_20795);
xnor U21003 (N_21003,N_20841,N_20948);
and U21004 (N_21004,N_20977,N_20807);
or U21005 (N_21005,N_20829,N_20883);
or U21006 (N_21006,N_20909,N_20904);
nor U21007 (N_21007,N_20990,N_20842);
nand U21008 (N_21008,N_20989,N_20801);
xor U21009 (N_21009,N_20938,N_20811);
and U21010 (N_21010,N_20789,N_20982);
nor U21011 (N_21011,N_20864,N_20913);
and U21012 (N_21012,N_20999,N_20939);
xnor U21013 (N_21013,N_20914,N_20884);
and U21014 (N_21014,N_20783,N_20954);
nand U21015 (N_21015,N_20784,N_20858);
xnor U21016 (N_21016,N_20959,N_20851);
nand U21017 (N_21017,N_20826,N_20926);
xnor U21018 (N_21018,N_20958,N_20855);
nor U21019 (N_21019,N_20768,N_20910);
nand U21020 (N_21020,N_20902,N_20906);
or U21021 (N_21021,N_20907,N_20928);
nor U21022 (N_21022,N_20940,N_20992);
nand U21023 (N_21023,N_20937,N_20885);
and U21024 (N_21024,N_20755,N_20837);
nor U21025 (N_21025,N_20993,N_20908);
or U21026 (N_21026,N_20896,N_20765);
xnor U21027 (N_21027,N_20818,N_20815);
and U21028 (N_21028,N_20934,N_20767);
or U21029 (N_21029,N_20964,N_20936);
xor U21030 (N_21030,N_20812,N_20780);
and U21031 (N_21031,N_20750,N_20875);
nor U21032 (N_21032,N_20856,N_20984);
xnor U21033 (N_21033,N_20862,N_20941);
or U21034 (N_21034,N_20873,N_20911);
and U21035 (N_21035,N_20876,N_20898);
nor U21036 (N_21036,N_20772,N_20854);
or U21037 (N_21037,N_20785,N_20878);
and U21038 (N_21038,N_20869,N_20790);
and U21039 (N_21039,N_20766,N_20979);
nor U21040 (N_21040,N_20761,N_20827);
and U21041 (N_21041,N_20857,N_20927);
or U21042 (N_21042,N_20974,N_20978);
nand U21043 (N_21043,N_20920,N_20887);
nor U21044 (N_21044,N_20833,N_20985);
xor U21045 (N_21045,N_20998,N_20921);
xor U21046 (N_21046,N_20882,N_20880);
or U21047 (N_21047,N_20915,N_20987);
and U21048 (N_21048,N_20966,N_20912);
nor U21049 (N_21049,N_20782,N_20774);
or U21050 (N_21050,N_20892,N_20751);
nor U21051 (N_21051,N_20968,N_20886);
nand U21052 (N_21052,N_20786,N_20753);
nor U21053 (N_21053,N_20961,N_20861);
nand U21054 (N_21054,N_20953,N_20770);
or U21055 (N_21055,N_20868,N_20895);
xnor U21056 (N_21056,N_20963,N_20798);
and U21057 (N_21057,N_20973,N_20943);
xor U21058 (N_21058,N_20757,N_20894);
nand U21059 (N_21059,N_20828,N_20891);
and U21060 (N_21060,N_20877,N_20781);
or U21061 (N_21061,N_20890,N_20849);
or U21062 (N_21062,N_20942,N_20771);
nor U21063 (N_21063,N_20946,N_20971);
nor U21064 (N_21064,N_20793,N_20778);
and U21065 (N_21065,N_20792,N_20756);
nor U21066 (N_21066,N_20922,N_20986);
nand U21067 (N_21067,N_20962,N_20846);
xnor U21068 (N_21068,N_20775,N_20867);
nor U21069 (N_21069,N_20802,N_20831);
xor U21070 (N_21070,N_20899,N_20860);
or U21071 (N_21071,N_20893,N_20845);
or U21072 (N_21072,N_20832,N_20931);
and U21073 (N_21073,N_20810,N_20835);
or U21074 (N_21074,N_20917,N_20859);
nor U21075 (N_21075,N_20866,N_20844);
or U21076 (N_21076,N_20944,N_20997);
and U21077 (N_21077,N_20821,N_20872);
xnor U21078 (N_21078,N_20791,N_20949);
xnor U21079 (N_21079,N_20769,N_20809);
nand U21080 (N_21080,N_20945,N_20776);
nor U21081 (N_21081,N_20988,N_20759);
and U21082 (N_21082,N_20779,N_20787);
or U21083 (N_21083,N_20897,N_20758);
and U21084 (N_21084,N_20960,N_20955);
or U21085 (N_21085,N_20799,N_20923);
xnor U21086 (N_21086,N_20918,N_20863);
nor U21087 (N_21087,N_20840,N_20814);
and U21088 (N_21088,N_20951,N_20889);
and U21089 (N_21089,N_20762,N_20817);
nand U21090 (N_21090,N_20773,N_20850);
xor U21091 (N_21091,N_20843,N_20975);
and U21092 (N_21092,N_20916,N_20800);
xnor U21093 (N_21093,N_20888,N_20839);
xor U21094 (N_21094,N_20870,N_20929);
or U21095 (N_21095,N_20957,N_20777);
and U21096 (N_21096,N_20794,N_20822);
nand U21097 (N_21097,N_20763,N_20865);
xnor U21098 (N_21098,N_20976,N_20819);
nand U21099 (N_21099,N_20806,N_20823);
nand U21100 (N_21100,N_20980,N_20919);
and U21101 (N_21101,N_20965,N_20830);
xnor U21102 (N_21102,N_20901,N_20797);
xnor U21103 (N_21103,N_20805,N_20788);
xnor U21104 (N_21104,N_20925,N_20760);
nand U21105 (N_21105,N_20838,N_20834);
nand U21106 (N_21106,N_20825,N_20852);
or U21107 (N_21107,N_20903,N_20900);
nand U21108 (N_21108,N_20932,N_20881);
nand U21109 (N_21109,N_20956,N_20947);
or U21110 (N_21110,N_20803,N_20995);
nor U21111 (N_21111,N_20935,N_20836);
nand U21112 (N_21112,N_20824,N_20991);
nand U21113 (N_21113,N_20933,N_20924);
nor U21114 (N_21114,N_20853,N_20871);
or U21115 (N_21115,N_20874,N_20970);
nor U21116 (N_21116,N_20905,N_20808);
nor U21117 (N_21117,N_20967,N_20804);
and U21118 (N_21118,N_20754,N_20969);
xnor U21119 (N_21119,N_20996,N_20972);
or U21120 (N_21120,N_20994,N_20796);
and U21121 (N_21121,N_20981,N_20847);
or U21122 (N_21122,N_20820,N_20983);
or U21123 (N_21123,N_20816,N_20813);
nand U21124 (N_21124,N_20879,N_20930);
xor U21125 (N_21125,N_20849,N_20907);
nand U21126 (N_21126,N_20932,N_20938);
or U21127 (N_21127,N_20929,N_20952);
xnor U21128 (N_21128,N_20905,N_20871);
nor U21129 (N_21129,N_20809,N_20983);
nand U21130 (N_21130,N_20953,N_20797);
nor U21131 (N_21131,N_20787,N_20780);
nand U21132 (N_21132,N_20914,N_20979);
nand U21133 (N_21133,N_20981,N_20820);
xnor U21134 (N_21134,N_20790,N_20988);
xnor U21135 (N_21135,N_20946,N_20855);
xnor U21136 (N_21136,N_20776,N_20988);
and U21137 (N_21137,N_20877,N_20902);
and U21138 (N_21138,N_20848,N_20850);
and U21139 (N_21139,N_20791,N_20919);
nand U21140 (N_21140,N_20947,N_20898);
or U21141 (N_21141,N_20859,N_20824);
nor U21142 (N_21142,N_20880,N_20949);
nor U21143 (N_21143,N_20814,N_20763);
nand U21144 (N_21144,N_20993,N_20845);
xnor U21145 (N_21145,N_20920,N_20910);
nand U21146 (N_21146,N_20841,N_20891);
nand U21147 (N_21147,N_20823,N_20845);
nand U21148 (N_21148,N_20887,N_20792);
or U21149 (N_21149,N_20941,N_20762);
xor U21150 (N_21150,N_20886,N_20751);
nand U21151 (N_21151,N_20957,N_20924);
nand U21152 (N_21152,N_20773,N_20759);
or U21153 (N_21153,N_20941,N_20866);
or U21154 (N_21154,N_20797,N_20781);
xnor U21155 (N_21155,N_20766,N_20892);
and U21156 (N_21156,N_20845,N_20797);
or U21157 (N_21157,N_20778,N_20887);
or U21158 (N_21158,N_20872,N_20953);
or U21159 (N_21159,N_20783,N_20832);
xnor U21160 (N_21160,N_20915,N_20990);
nor U21161 (N_21161,N_20767,N_20940);
nor U21162 (N_21162,N_20766,N_20860);
or U21163 (N_21163,N_20966,N_20821);
and U21164 (N_21164,N_20859,N_20963);
xor U21165 (N_21165,N_20891,N_20899);
xor U21166 (N_21166,N_20967,N_20784);
nor U21167 (N_21167,N_20962,N_20767);
nand U21168 (N_21168,N_20833,N_20764);
and U21169 (N_21169,N_20760,N_20970);
and U21170 (N_21170,N_20889,N_20924);
xor U21171 (N_21171,N_20951,N_20922);
nand U21172 (N_21172,N_20888,N_20894);
and U21173 (N_21173,N_20855,N_20898);
nand U21174 (N_21174,N_20968,N_20957);
nor U21175 (N_21175,N_20938,N_20864);
and U21176 (N_21176,N_20768,N_20801);
and U21177 (N_21177,N_20922,N_20969);
xnor U21178 (N_21178,N_20775,N_20955);
nand U21179 (N_21179,N_20895,N_20894);
nand U21180 (N_21180,N_20953,N_20914);
nor U21181 (N_21181,N_20806,N_20779);
or U21182 (N_21182,N_20812,N_20962);
and U21183 (N_21183,N_20954,N_20772);
nor U21184 (N_21184,N_20933,N_20860);
nor U21185 (N_21185,N_20999,N_20958);
xnor U21186 (N_21186,N_20825,N_20865);
nand U21187 (N_21187,N_20866,N_20901);
nor U21188 (N_21188,N_20927,N_20998);
or U21189 (N_21189,N_20856,N_20900);
xor U21190 (N_21190,N_20751,N_20783);
or U21191 (N_21191,N_20980,N_20815);
xor U21192 (N_21192,N_20847,N_20979);
or U21193 (N_21193,N_20804,N_20752);
and U21194 (N_21194,N_20970,N_20777);
nand U21195 (N_21195,N_20991,N_20861);
nor U21196 (N_21196,N_20869,N_20811);
or U21197 (N_21197,N_20842,N_20950);
and U21198 (N_21198,N_20771,N_20979);
xor U21199 (N_21199,N_20882,N_20818);
or U21200 (N_21200,N_20902,N_20858);
xor U21201 (N_21201,N_20772,N_20866);
nand U21202 (N_21202,N_20823,N_20966);
nor U21203 (N_21203,N_20990,N_20936);
nand U21204 (N_21204,N_20840,N_20888);
or U21205 (N_21205,N_20894,N_20843);
or U21206 (N_21206,N_20765,N_20809);
nand U21207 (N_21207,N_20894,N_20791);
nand U21208 (N_21208,N_20930,N_20858);
xnor U21209 (N_21209,N_20815,N_20811);
nand U21210 (N_21210,N_20981,N_20859);
and U21211 (N_21211,N_20784,N_20854);
nand U21212 (N_21212,N_20918,N_20888);
xnor U21213 (N_21213,N_20991,N_20759);
or U21214 (N_21214,N_20964,N_20866);
and U21215 (N_21215,N_20979,N_20951);
nand U21216 (N_21216,N_20847,N_20805);
or U21217 (N_21217,N_20961,N_20965);
nand U21218 (N_21218,N_20754,N_20915);
and U21219 (N_21219,N_20994,N_20841);
or U21220 (N_21220,N_20793,N_20856);
or U21221 (N_21221,N_20926,N_20800);
and U21222 (N_21222,N_20821,N_20931);
nor U21223 (N_21223,N_20961,N_20818);
xnor U21224 (N_21224,N_20927,N_20808);
xor U21225 (N_21225,N_20754,N_20781);
xor U21226 (N_21226,N_20888,N_20838);
xor U21227 (N_21227,N_20822,N_20796);
or U21228 (N_21228,N_20887,N_20900);
nand U21229 (N_21229,N_20971,N_20796);
or U21230 (N_21230,N_20803,N_20927);
or U21231 (N_21231,N_20752,N_20798);
xor U21232 (N_21232,N_20799,N_20901);
nand U21233 (N_21233,N_20816,N_20826);
or U21234 (N_21234,N_20957,N_20844);
xor U21235 (N_21235,N_20946,N_20982);
or U21236 (N_21236,N_20970,N_20794);
nor U21237 (N_21237,N_20784,N_20935);
and U21238 (N_21238,N_20925,N_20954);
nor U21239 (N_21239,N_20823,N_20910);
or U21240 (N_21240,N_20992,N_20789);
nor U21241 (N_21241,N_20845,N_20885);
and U21242 (N_21242,N_20755,N_20921);
nor U21243 (N_21243,N_20839,N_20936);
or U21244 (N_21244,N_20781,N_20911);
nand U21245 (N_21245,N_20983,N_20828);
xor U21246 (N_21246,N_20962,N_20798);
nor U21247 (N_21247,N_20814,N_20801);
or U21248 (N_21248,N_20976,N_20788);
and U21249 (N_21249,N_20926,N_20933);
and U21250 (N_21250,N_21238,N_21166);
or U21251 (N_21251,N_21157,N_21162);
xnor U21252 (N_21252,N_21116,N_21120);
nor U21253 (N_21253,N_21058,N_21081);
and U21254 (N_21254,N_21046,N_21193);
or U21255 (N_21255,N_21156,N_21073);
nand U21256 (N_21256,N_21104,N_21095);
nor U21257 (N_21257,N_21235,N_21054);
xnor U21258 (N_21258,N_21138,N_21124);
nor U21259 (N_21259,N_21152,N_21018);
and U21260 (N_21260,N_21014,N_21128);
nor U21261 (N_21261,N_21146,N_21107);
nor U21262 (N_21262,N_21165,N_21100);
xor U21263 (N_21263,N_21143,N_21249);
nand U21264 (N_21264,N_21209,N_21180);
nand U21265 (N_21265,N_21139,N_21178);
nor U21266 (N_21266,N_21030,N_21201);
or U21267 (N_21267,N_21223,N_21111);
or U21268 (N_21268,N_21089,N_21169);
and U21269 (N_21269,N_21174,N_21145);
nor U21270 (N_21270,N_21133,N_21117);
nand U21271 (N_21271,N_21024,N_21130);
nand U21272 (N_21272,N_21034,N_21211);
or U21273 (N_21273,N_21028,N_21083);
xnor U21274 (N_21274,N_21237,N_21096);
nand U21275 (N_21275,N_21017,N_21231);
or U21276 (N_21276,N_21086,N_21079);
or U21277 (N_21277,N_21112,N_21230);
xnor U21278 (N_21278,N_21021,N_21229);
and U21279 (N_21279,N_21233,N_21093);
or U21280 (N_21280,N_21189,N_21177);
and U21281 (N_21281,N_21052,N_21232);
and U21282 (N_21282,N_21023,N_21241);
xnor U21283 (N_21283,N_21234,N_21218);
or U21284 (N_21284,N_21029,N_21153);
or U21285 (N_21285,N_21142,N_21092);
nor U21286 (N_21286,N_21216,N_21125);
nor U21287 (N_21287,N_21063,N_21057);
and U21288 (N_21288,N_21248,N_21160);
nand U21289 (N_21289,N_21167,N_21186);
nor U21290 (N_21290,N_21147,N_21008);
nor U21291 (N_21291,N_21072,N_21042);
nor U21292 (N_21292,N_21069,N_21078);
xor U21293 (N_21293,N_21199,N_21219);
xnor U21294 (N_21294,N_21048,N_21011);
nor U21295 (N_21295,N_21002,N_21194);
xnor U21296 (N_21296,N_21026,N_21141);
nor U21297 (N_21297,N_21051,N_21094);
or U21298 (N_21298,N_21053,N_21135);
xor U21299 (N_21299,N_21105,N_21070);
nand U21300 (N_21300,N_21032,N_21010);
nor U21301 (N_21301,N_21164,N_21060);
xor U21302 (N_21302,N_21190,N_21119);
or U21303 (N_21303,N_21181,N_21213);
nand U21304 (N_21304,N_21087,N_21085);
nand U21305 (N_21305,N_21038,N_21245);
xnor U21306 (N_21306,N_21061,N_21033);
xnor U21307 (N_21307,N_21197,N_21025);
and U21308 (N_21308,N_21227,N_21084);
and U21309 (N_21309,N_21191,N_21000);
or U21310 (N_21310,N_21110,N_21236);
or U21311 (N_21311,N_21102,N_21071);
or U21312 (N_21312,N_21019,N_21035);
nand U21313 (N_21313,N_21240,N_21168);
and U21314 (N_21314,N_21013,N_21088);
xor U21315 (N_21315,N_21055,N_21045);
nand U21316 (N_21316,N_21243,N_21212);
nor U21317 (N_21317,N_21108,N_21208);
and U21318 (N_21318,N_21115,N_21132);
xnor U21319 (N_21319,N_21082,N_21012);
and U21320 (N_21320,N_21161,N_21150);
and U21321 (N_21321,N_21202,N_21056);
and U21322 (N_21322,N_21050,N_21144);
or U21323 (N_21323,N_21170,N_21151);
and U21324 (N_21324,N_21247,N_21159);
xor U21325 (N_21325,N_21003,N_21076);
xnor U21326 (N_21326,N_21196,N_21204);
nor U21327 (N_21327,N_21106,N_21068);
or U21328 (N_21328,N_21109,N_21040);
xor U21329 (N_21329,N_21075,N_21155);
nor U21330 (N_21330,N_21136,N_21210);
or U21331 (N_21331,N_21039,N_21121);
nor U21332 (N_21332,N_21214,N_21066);
nor U21333 (N_21333,N_21239,N_21200);
nand U21334 (N_21334,N_21185,N_21036);
nand U21335 (N_21335,N_21044,N_21059);
xor U21336 (N_21336,N_21226,N_21148);
or U21337 (N_21337,N_21001,N_21080);
and U21338 (N_21338,N_21015,N_21022);
xnor U21339 (N_21339,N_21221,N_21005);
nor U21340 (N_21340,N_21224,N_21041);
nor U21341 (N_21341,N_21004,N_21103);
nand U21342 (N_21342,N_21244,N_21172);
nor U21343 (N_21343,N_21043,N_21198);
xnor U21344 (N_21344,N_21016,N_21182);
nor U21345 (N_21345,N_21126,N_21077);
and U21346 (N_21346,N_21175,N_21009);
xnor U21347 (N_21347,N_21206,N_21207);
or U21348 (N_21348,N_21065,N_21074);
xnor U21349 (N_21349,N_21154,N_21027);
nand U21350 (N_21350,N_21064,N_21140);
and U21351 (N_21351,N_21137,N_21228);
and U21352 (N_21352,N_21099,N_21183);
xnor U21353 (N_21353,N_21006,N_21203);
xor U21354 (N_21354,N_21134,N_21188);
and U21355 (N_21355,N_21158,N_21215);
and U21356 (N_21356,N_21205,N_21222);
and U21357 (N_21357,N_21176,N_21163);
or U21358 (N_21358,N_21217,N_21114);
or U21359 (N_21359,N_21220,N_21122);
or U21360 (N_21360,N_21127,N_21020);
nand U21361 (N_21361,N_21242,N_21131);
or U21362 (N_21362,N_21225,N_21179);
nand U21363 (N_21363,N_21062,N_21187);
and U21364 (N_21364,N_21173,N_21101);
nor U21365 (N_21365,N_21192,N_21123);
xor U21366 (N_21366,N_21097,N_21246);
nor U21367 (N_21367,N_21184,N_21047);
or U21368 (N_21368,N_21195,N_21091);
and U21369 (N_21369,N_21113,N_21067);
or U21370 (N_21370,N_21049,N_21031);
nand U21371 (N_21371,N_21118,N_21171);
xnor U21372 (N_21372,N_21129,N_21007);
xor U21373 (N_21373,N_21149,N_21037);
nor U21374 (N_21374,N_21090,N_21098);
nor U21375 (N_21375,N_21243,N_21027);
nand U21376 (N_21376,N_21105,N_21133);
xnor U21377 (N_21377,N_21047,N_21229);
nor U21378 (N_21378,N_21017,N_21010);
nor U21379 (N_21379,N_21024,N_21083);
or U21380 (N_21380,N_21234,N_21023);
and U21381 (N_21381,N_21203,N_21157);
or U21382 (N_21382,N_21040,N_21159);
nand U21383 (N_21383,N_21115,N_21162);
xor U21384 (N_21384,N_21075,N_21056);
or U21385 (N_21385,N_21090,N_21081);
or U21386 (N_21386,N_21216,N_21051);
nand U21387 (N_21387,N_21179,N_21000);
xnor U21388 (N_21388,N_21098,N_21209);
and U21389 (N_21389,N_21171,N_21205);
or U21390 (N_21390,N_21032,N_21047);
and U21391 (N_21391,N_21246,N_21249);
nor U21392 (N_21392,N_21011,N_21173);
nand U21393 (N_21393,N_21086,N_21141);
xnor U21394 (N_21394,N_21214,N_21161);
and U21395 (N_21395,N_21037,N_21019);
xnor U21396 (N_21396,N_21100,N_21109);
nand U21397 (N_21397,N_21165,N_21120);
xor U21398 (N_21398,N_21142,N_21164);
and U21399 (N_21399,N_21016,N_21174);
nor U21400 (N_21400,N_21124,N_21226);
nand U21401 (N_21401,N_21158,N_21140);
nand U21402 (N_21402,N_21140,N_21226);
or U21403 (N_21403,N_21204,N_21005);
nand U21404 (N_21404,N_21010,N_21245);
xnor U21405 (N_21405,N_21219,N_21104);
or U21406 (N_21406,N_21083,N_21051);
nor U21407 (N_21407,N_21003,N_21043);
nor U21408 (N_21408,N_21079,N_21012);
and U21409 (N_21409,N_21222,N_21033);
nor U21410 (N_21410,N_21170,N_21046);
and U21411 (N_21411,N_21127,N_21225);
nor U21412 (N_21412,N_21191,N_21005);
nand U21413 (N_21413,N_21215,N_21087);
nor U21414 (N_21414,N_21130,N_21245);
xor U21415 (N_21415,N_21188,N_21185);
and U21416 (N_21416,N_21218,N_21146);
xor U21417 (N_21417,N_21014,N_21078);
xnor U21418 (N_21418,N_21149,N_21027);
nand U21419 (N_21419,N_21192,N_21127);
xor U21420 (N_21420,N_21054,N_21138);
and U21421 (N_21421,N_21155,N_21228);
and U21422 (N_21422,N_21116,N_21012);
and U21423 (N_21423,N_21215,N_21130);
nand U21424 (N_21424,N_21200,N_21128);
nor U21425 (N_21425,N_21192,N_21175);
nor U21426 (N_21426,N_21034,N_21075);
xnor U21427 (N_21427,N_21161,N_21009);
nor U21428 (N_21428,N_21232,N_21118);
xor U21429 (N_21429,N_21191,N_21050);
nor U21430 (N_21430,N_21156,N_21181);
or U21431 (N_21431,N_21125,N_21001);
nand U21432 (N_21432,N_21134,N_21215);
and U21433 (N_21433,N_21107,N_21240);
xnor U21434 (N_21434,N_21120,N_21089);
xor U21435 (N_21435,N_21219,N_21214);
nor U21436 (N_21436,N_21083,N_21184);
nor U21437 (N_21437,N_21095,N_21040);
xnor U21438 (N_21438,N_21214,N_21043);
or U21439 (N_21439,N_21072,N_21151);
nor U21440 (N_21440,N_21236,N_21228);
or U21441 (N_21441,N_21133,N_21008);
xnor U21442 (N_21442,N_21007,N_21239);
or U21443 (N_21443,N_21057,N_21014);
nand U21444 (N_21444,N_21219,N_21184);
nand U21445 (N_21445,N_21248,N_21096);
and U21446 (N_21446,N_21211,N_21145);
and U21447 (N_21447,N_21236,N_21073);
xor U21448 (N_21448,N_21038,N_21092);
nand U21449 (N_21449,N_21172,N_21170);
nor U21450 (N_21450,N_21167,N_21045);
and U21451 (N_21451,N_21115,N_21247);
or U21452 (N_21452,N_21123,N_21080);
and U21453 (N_21453,N_21163,N_21178);
nor U21454 (N_21454,N_21174,N_21108);
or U21455 (N_21455,N_21109,N_21021);
and U21456 (N_21456,N_21007,N_21131);
and U21457 (N_21457,N_21219,N_21044);
or U21458 (N_21458,N_21194,N_21127);
nor U21459 (N_21459,N_21054,N_21106);
xor U21460 (N_21460,N_21109,N_21081);
or U21461 (N_21461,N_21046,N_21103);
or U21462 (N_21462,N_21084,N_21140);
nand U21463 (N_21463,N_21000,N_21031);
nand U21464 (N_21464,N_21241,N_21032);
or U21465 (N_21465,N_21225,N_21211);
xor U21466 (N_21466,N_21067,N_21029);
nor U21467 (N_21467,N_21235,N_21169);
nor U21468 (N_21468,N_21181,N_21138);
nand U21469 (N_21469,N_21219,N_21175);
and U21470 (N_21470,N_21133,N_21076);
xnor U21471 (N_21471,N_21125,N_21188);
or U21472 (N_21472,N_21181,N_21220);
or U21473 (N_21473,N_21004,N_21245);
xnor U21474 (N_21474,N_21012,N_21094);
and U21475 (N_21475,N_21060,N_21101);
xnor U21476 (N_21476,N_21220,N_21173);
nor U21477 (N_21477,N_21048,N_21216);
nor U21478 (N_21478,N_21219,N_21119);
nand U21479 (N_21479,N_21042,N_21044);
nand U21480 (N_21480,N_21150,N_21022);
nor U21481 (N_21481,N_21210,N_21215);
nor U21482 (N_21482,N_21245,N_21111);
or U21483 (N_21483,N_21082,N_21121);
xnor U21484 (N_21484,N_21047,N_21044);
xnor U21485 (N_21485,N_21056,N_21234);
and U21486 (N_21486,N_21067,N_21183);
nor U21487 (N_21487,N_21171,N_21165);
xnor U21488 (N_21488,N_21223,N_21069);
nand U21489 (N_21489,N_21204,N_21000);
nor U21490 (N_21490,N_21153,N_21217);
nand U21491 (N_21491,N_21207,N_21040);
nand U21492 (N_21492,N_21057,N_21128);
nor U21493 (N_21493,N_21174,N_21075);
and U21494 (N_21494,N_21146,N_21249);
xnor U21495 (N_21495,N_21029,N_21050);
or U21496 (N_21496,N_21081,N_21201);
or U21497 (N_21497,N_21221,N_21146);
and U21498 (N_21498,N_21050,N_21172);
xnor U21499 (N_21499,N_21160,N_21096);
xor U21500 (N_21500,N_21281,N_21304);
or U21501 (N_21501,N_21292,N_21453);
and U21502 (N_21502,N_21349,N_21339);
nand U21503 (N_21503,N_21340,N_21479);
xor U21504 (N_21504,N_21498,N_21378);
and U21505 (N_21505,N_21363,N_21345);
xor U21506 (N_21506,N_21254,N_21399);
xor U21507 (N_21507,N_21491,N_21468);
and U21508 (N_21508,N_21428,N_21497);
nand U21509 (N_21509,N_21300,N_21402);
nor U21510 (N_21510,N_21429,N_21407);
or U21511 (N_21511,N_21320,N_21411);
or U21512 (N_21512,N_21288,N_21344);
nand U21513 (N_21513,N_21482,N_21371);
xnor U21514 (N_21514,N_21357,N_21303);
or U21515 (N_21515,N_21393,N_21256);
xor U21516 (N_21516,N_21440,N_21492);
nor U21517 (N_21517,N_21406,N_21298);
xor U21518 (N_21518,N_21352,N_21255);
nor U21519 (N_21519,N_21251,N_21365);
and U21520 (N_21520,N_21471,N_21457);
and U21521 (N_21521,N_21328,N_21469);
or U21522 (N_21522,N_21348,N_21419);
xor U21523 (N_21523,N_21416,N_21262);
or U21524 (N_21524,N_21435,N_21350);
nor U21525 (N_21525,N_21316,N_21494);
xnor U21526 (N_21526,N_21372,N_21408);
nor U21527 (N_21527,N_21327,N_21282);
xnor U21528 (N_21528,N_21370,N_21484);
and U21529 (N_21529,N_21276,N_21272);
or U21530 (N_21530,N_21331,N_21455);
nand U21531 (N_21531,N_21477,N_21286);
xor U21532 (N_21532,N_21376,N_21444);
or U21533 (N_21533,N_21330,N_21431);
nand U21534 (N_21534,N_21325,N_21369);
nor U21535 (N_21535,N_21436,N_21391);
nor U21536 (N_21536,N_21359,N_21480);
nand U21537 (N_21537,N_21441,N_21293);
and U21538 (N_21538,N_21258,N_21485);
or U21539 (N_21539,N_21317,N_21486);
nand U21540 (N_21540,N_21499,N_21319);
or U21541 (N_21541,N_21366,N_21358);
and U21542 (N_21542,N_21367,N_21297);
and U21543 (N_21543,N_21261,N_21489);
nor U21544 (N_21544,N_21334,N_21470);
nand U21545 (N_21545,N_21379,N_21315);
xnor U21546 (N_21546,N_21375,N_21259);
nor U21547 (N_21547,N_21437,N_21373);
or U21548 (N_21548,N_21301,N_21314);
nor U21549 (N_21549,N_21417,N_21487);
and U21550 (N_21550,N_21267,N_21451);
nand U21551 (N_21551,N_21380,N_21287);
xnor U21552 (N_21552,N_21253,N_21302);
and U21553 (N_21553,N_21414,N_21341);
xnor U21554 (N_21554,N_21274,N_21461);
nor U21555 (N_21555,N_21332,N_21462);
xor U21556 (N_21556,N_21443,N_21432);
nor U21557 (N_21557,N_21454,N_21335);
and U21558 (N_21558,N_21280,N_21450);
or U21559 (N_21559,N_21475,N_21313);
nand U21560 (N_21560,N_21397,N_21275);
nand U21561 (N_21561,N_21270,N_21488);
nand U21562 (N_21562,N_21307,N_21438);
xnor U21563 (N_21563,N_21377,N_21420);
nor U21564 (N_21564,N_21427,N_21278);
and U21565 (N_21565,N_21310,N_21362);
nor U21566 (N_21566,N_21329,N_21311);
xor U21567 (N_21567,N_21333,N_21264);
xor U21568 (N_21568,N_21446,N_21291);
or U21569 (N_21569,N_21347,N_21382);
nand U21570 (N_21570,N_21252,N_21257);
and U21571 (N_21571,N_21424,N_21434);
xor U21572 (N_21572,N_21495,N_21452);
and U21573 (N_21573,N_21422,N_21405);
xor U21574 (N_21574,N_21390,N_21456);
nor U21575 (N_21575,N_21409,N_21263);
xor U21576 (N_21576,N_21442,N_21290);
nor U21577 (N_21577,N_21386,N_21396);
nor U21578 (N_21578,N_21299,N_21439);
nand U21579 (N_21579,N_21460,N_21318);
and U21580 (N_21580,N_21490,N_21426);
or U21581 (N_21581,N_21351,N_21392);
nor U21582 (N_21582,N_21463,N_21493);
or U21583 (N_21583,N_21284,N_21295);
xor U21584 (N_21584,N_21354,N_21445);
xor U21585 (N_21585,N_21364,N_21472);
or U21586 (N_21586,N_21296,N_21374);
or U21587 (N_21587,N_21476,N_21277);
nor U21588 (N_21588,N_21342,N_21459);
nand U21589 (N_21589,N_21400,N_21273);
nand U21590 (N_21590,N_21271,N_21323);
xor U21591 (N_21591,N_21404,N_21324);
or U21592 (N_21592,N_21421,N_21337);
nor U21593 (N_21593,N_21388,N_21481);
xnor U21594 (N_21594,N_21321,N_21448);
nor U21595 (N_21595,N_21285,N_21410);
xnor U21596 (N_21596,N_21346,N_21464);
nor U21597 (N_21597,N_21389,N_21355);
or U21598 (N_21598,N_21343,N_21353);
xnor U21599 (N_21599,N_21401,N_21360);
xnor U21600 (N_21600,N_21467,N_21423);
xnor U21601 (N_21601,N_21425,N_21387);
or U21602 (N_21602,N_21415,N_21356);
xnor U21603 (N_21603,N_21458,N_21403);
nor U21604 (N_21604,N_21381,N_21473);
nor U21605 (N_21605,N_21308,N_21398);
xnor U21606 (N_21606,N_21266,N_21269);
nor U21607 (N_21607,N_21412,N_21326);
or U21608 (N_21608,N_21433,N_21368);
xnor U21609 (N_21609,N_21361,N_21250);
nor U21610 (N_21610,N_21395,N_21265);
nor U21611 (N_21611,N_21283,N_21384);
or U21612 (N_21612,N_21394,N_21336);
nand U21613 (N_21613,N_21385,N_21418);
xor U21614 (N_21614,N_21483,N_21322);
nand U21615 (N_21615,N_21447,N_21306);
nand U21616 (N_21616,N_21466,N_21449);
nor U21617 (N_21617,N_21338,N_21496);
and U21618 (N_21618,N_21279,N_21305);
nor U21619 (N_21619,N_21474,N_21268);
nor U21620 (N_21620,N_21294,N_21260);
xnor U21621 (N_21621,N_21478,N_21383);
and U21622 (N_21622,N_21413,N_21430);
nor U21623 (N_21623,N_21465,N_21289);
and U21624 (N_21624,N_21309,N_21312);
nor U21625 (N_21625,N_21467,N_21295);
nand U21626 (N_21626,N_21347,N_21409);
nor U21627 (N_21627,N_21314,N_21402);
xnor U21628 (N_21628,N_21492,N_21359);
xnor U21629 (N_21629,N_21364,N_21478);
or U21630 (N_21630,N_21488,N_21311);
nand U21631 (N_21631,N_21252,N_21312);
and U21632 (N_21632,N_21331,N_21394);
nor U21633 (N_21633,N_21307,N_21385);
or U21634 (N_21634,N_21392,N_21491);
and U21635 (N_21635,N_21263,N_21387);
or U21636 (N_21636,N_21369,N_21451);
and U21637 (N_21637,N_21467,N_21339);
and U21638 (N_21638,N_21296,N_21301);
nor U21639 (N_21639,N_21282,N_21289);
or U21640 (N_21640,N_21440,N_21351);
or U21641 (N_21641,N_21255,N_21432);
and U21642 (N_21642,N_21418,N_21478);
nor U21643 (N_21643,N_21274,N_21389);
and U21644 (N_21644,N_21470,N_21294);
and U21645 (N_21645,N_21464,N_21425);
nand U21646 (N_21646,N_21388,N_21469);
xnor U21647 (N_21647,N_21278,N_21377);
nor U21648 (N_21648,N_21275,N_21282);
nand U21649 (N_21649,N_21259,N_21438);
and U21650 (N_21650,N_21486,N_21424);
xor U21651 (N_21651,N_21263,N_21463);
nand U21652 (N_21652,N_21463,N_21308);
and U21653 (N_21653,N_21394,N_21431);
and U21654 (N_21654,N_21357,N_21374);
nand U21655 (N_21655,N_21302,N_21460);
xnor U21656 (N_21656,N_21439,N_21415);
and U21657 (N_21657,N_21386,N_21271);
or U21658 (N_21658,N_21254,N_21482);
nor U21659 (N_21659,N_21340,N_21465);
and U21660 (N_21660,N_21401,N_21481);
xor U21661 (N_21661,N_21270,N_21403);
nor U21662 (N_21662,N_21329,N_21438);
xor U21663 (N_21663,N_21443,N_21445);
and U21664 (N_21664,N_21446,N_21346);
xor U21665 (N_21665,N_21483,N_21330);
and U21666 (N_21666,N_21272,N_21356);
nor U21667 (N_21667,N_21458,N_21417);
nor U21668 (N_21668,N_21447,N_21261);
nand U21669 (N_21669,N_21361,N_21253);
and U21670 (N_21670,N_21368,N_21333);
nand U21671 (N_21671,N_21433,N_21439);
xor U21672 (N_21672,N_21387,N_21473);
xnor U21673 (N_21673,N_21421,N_21268);
nor U21674 (N_21674,N_21452,N_21326);
xnor U21675 (N_21675,N_21447,N_21369);
nor U21676 (N_21676,N_21331,N_21453);
xor U21677 (N_21677,N_21271,N_21446);
and U21678 (N_21678,N_21352,N_21333);
nor U21679 (N_21679,N_21320,N_21254);
nand U21680 (N_21680,N_21312,N_21429);
nand U21681 (N_21681,N_21473,N_21362);
or U21682 (N_21682,N_21496,N_21386);
nand U21683 (N_21683,N_21273,N_21337);
xnor U21684 (N_21684,N_21404,N_21325);
or U21685 (N_21685,N_21275,N_21377);
xnor U21686 (N_21686,N_21374,N_21290);
nand U21687 (N_21687,N_21499,N_21397);
xor U21688 (N_21688,N_21305,N_21446);
nand U21689 (N_21689,N_21284,N_21420);
or U21690 (N_21690,N_21420,N_21270);
xor U21691 (N_21691,N_21405,N_21453);
and U21692 (N_21692,N_21475,N_21406);
nor U21693 (N_21693,N_21464,N_21419);
nand U21694 (N_21694,N_21405,N_21318);
nor U21695 (N_21695,N_21422,N_21292);
nand U21696 (N_21696,N_21445,N_21447);
and U21697 (N_21697,N_21416,N_21276);
and U21698 (N_21698,N_21287,N_21294);
xnor U21699 (N_21699,N_21293,N_21490);
or U21700 (N_21700,N_21361,N_21445);
nand U21701 (N_21701,N_21463,N_21452);
or U21702 (N_21702,N_21414,N_21477);
nor U21703 (N_21703,N_21424,N_21451);
and U21704 (N_21704,N_21331,N_21277);
and U21705 (N_21705,N_21327,N_21376);
nor U21706 (N_21706,N_21341,N_21359);
nand U21707 (N_21707,N_21342,N_21373);
nor U21708 (N_21708,N_21288,N_21364);
or U21709 (N_21709,N_21382,N_21251);
xnor U21710 (N_21710,N_21263,N_21383);
nor U21711 (N_21711,N_21383,N_21447);
or U21712 (N_21712,N_21256,N_21478);
or U21713 (N_21713,N_21285,N_21413);
nor U21714 (N_21714,N_21484,N_21302);
nor U21715 (N_21715,N_21415,N_21291);
nor U21716 (N_21716,N_21312,N_21392);
nand U21717 (N_21717,N_21303,N_21285);
nand U21718 (N_21718,N_21377,N_21424);
nand U21719 (N_21719,N_21320,N_21481);
nand U21720 (N_21720,N_21250,N_21471);
xnor U21721 (N_21721,N_21345,N_21269);
or U21722 (N_21722,N_21488,N_21437);
xor U21723 (N_21723,N_21402,N_21471);
or U21724 (N_21724,N_21454,N_21387);
xor U21725 (N_21725,N_21320,N_21425);
and U21726 (N_21726,N_21421,N_21485);
or U21727 (N_21727,N_21296,N_21263);
or U21728 (N_21728,N_21304,N_21375);
or U21729 (N_21729,N_21402,N_21455);
or U21730 (N_21730,N_21408,N_21486);
or U21731 (N_21731,N_21467,N_21293);
xnor U21732 (N_21732,N_21458,N_21309);
nor U21733 (N_21733,N_21252,N_21411);
and U21734 (N_21734,N_21340,N_21323);
nand U21735 (N_21735,N_21329,N_21340);
and U21736 (N_21736,N_21489,N_21349);
or U21737 (N_21737,N_21273,N_21387);
nand U21738 (N_21738,N_21292,N_21309);
nor U21739 (N_21739,N_21373,N_21273);
nor U21740 (N_21740,N_21279,N_21324);
or U21741 (N_21741,N_21316,N_21492);
nor U21742 (N_21742,N_21442,N_21418);
and U21743 (N_21743,N_21498,N_21258);
and U21744 (N_21744,N_21390,N_21337);
nand U21745 (N_21745,N_21328,N_21343);
or U21746 (N_21746,N_21488,N_21445);
nand U21747 (N_21747,N_21425,N_21311);
nand U21748 (N_21748,N_21420,N_21308);
xor U21749 (N_21749,N_21363,N_21288);
nor U21750 (N_21750,N_21747,N_21518);
nand U21751 (N_21751,N_21500,N_21511);
nand U21752 (N_21752,N_21633,N_21584);
or U21753 (N_21753,N_21550,N_21555);
nor U21754 (N_21754,N_21706,N_21577);
xor U21755 (N_21755,N_21733,N_21531);
nor U21756 (N_21756,N_21696,N_21582);
xnor U21757 (N_21757,N_21667,N_21662);
or U21758 (N_21758,N_21722,N_21532);
and U21759 (N_21759,N_21638,N_21612);
xor U21760 (N_21760,N_21716,N_21668);
nor U21761 (N_21761,N_21519,N_21514);
nor U21762 (N_21762,N_21601,N_21598);
nor U21763 (N_21763,N_21656,N_21501);
and U21764 (N_21764,N_21551,N_21536);
nor U21765 (N_21765,N_21544,N_21527);
nor U21766 (N_21766,N_21558,N_21541);
and U21767 (N_21767,N_21507,N_21505);
nand U21768 (N_21768,N_21708,N_21520);
nor U21769 (N_21769,N_21607,N_21628);
xnor U21770 (N_21770,N_21659,N_21560);
and U21771 (N_21771,N_21545,N_21744);
xnor U21772 (N_21772,N_21661,N_21743);
nand U21773 (N_21773,N_21583,N_21516);
and U21774 (N_21774,N_21569,N_21637);
nor U21775 (N_21775,N_21735,N_21634);
xor U21776 (N_21776,N_21554,N_21515);
xnor U21777 (N_21777,N_21508,N_21564);
or U21778 (N_21778,N_21680,N_21692);
nor U21779 (N_21779,N_21713,N_21586);
nor U21780 (N_21780,N_21610,N_21710);
and U21781 (N_21781,N_21619,N_21618);
nand U21782 (N_21782,N_21694,N_21709);
or U21783 (N_21783,N_21512,N_21556);
xnor U21784 (N_21784,N_21526,N_21746);
or U21785 (N_21785,N_21685,N_21537);
nand U21786 (N_21786,N_21630,N_21721);
and U21787 (N_21787,N_21543,N_21566);
xnor U21788 (N_21788,N_21681,N_21734);
or U21789 (N_21789,N_21533,N_21621);
nor U21790 (N_21790,N_21625,N_21687);
nor U21791 (N_21791,N_21711,N_21671);
or U21792 (N_21792,N_21674,N_21645);
xor U21793 (N_21793,N_21652,N_21684);
and U21794 (N_21794,N_21732,N_21540);
and U21795 (N_21795,N_21641,N_21592);
nor U21796 (N_21796,N_21563,N_21657);
or U21797 (N_21797,N_21655,N_21615);
or U21798 (N_21798,N_21702,N_21594);
xor U21799 (N_21799,N_21620,N_21595);
or U21800 (N_21800,N_21679,N_21600);
nor U21801 (N_21801,N_21596,N_21683);
and U21802 (N_21802,N_21712,N_21725);
nand U21803 (N_21803,N_21559,N_21640);
xnor U21804 (N_21804,N_21742,N_21572);
xor U21805 (N_21805,N_21636,N_21647);
xnor U21806 (N_21806,N_21728,N_21593);
nand U21807 (N_21807,N_21573,N_21547);
nand U21808 (N_21808,N_21529,N_21650);
xnor U21809 (N_21809,N_21642,N_21521);
xnor U21810 (N_21810,N_21729,N_21691);
nand U21811 (N_21811,N_21718,N_21568);
nand U21812 (N_21812,N_21609,N_21654);
and U21813 (N_21813,N_21737,N_21749);
and U21814 (N_21814,N_21567,N_21597);
xor U21815 (N_21815,N_21693,N_21602);
and U21816 (N_21816,N_21688,N_21528);
and U21817 (N_21817,N_21736,N_21522);
and U21818 (N_21818,N_21686,N_21627);
xnor U21819 (N_21819,N_21579,N_21666);
xor U21820 (N_21820,N_21703,N_21726);
and U21821 (N_21821,N_21606,N_21631);
nand U21822 (N_21822,N_21727,N_21665);
nand U21823 (N_21823,N_21689,N_21523);
nor U21824 (N_21824,N_21715,N_21701);
or U21825 (N_21825,N_21614,N_21678);
and U21826 (N_21826,N_21739,N_21629);
or U21827 (N_21827,N_21660,N_21509);
xnor U21828 (N_21828,N_21599,N_21622);
or U21829 (N_21829,N_21644,N_21730);
or U21830 (N_21830,N_21670,N_21605);
nand U21831 (N_21831,N_21731,N_21570);
nand U21832 (N_21832,N_21672,N_21546);
and U21833 (N_21833,N_21651,N_21695);
and U21834 (N_21834,N_21676,N_21574);
xnor U21835 (N_21835,N_21603,N_21571);
nor U21836 (N_21836,N_21530,N_21673);
nand U21837 (N_21837,N_21617,N_21604);
or U21838 (N_21838,N_21517,N_21538);
and U21839 (N_21839,N_21646,N_21669);
and U21840 (N_21840,N_21704,N_21707);
nand U21841 (N_21841,N_21626,N_21697);
nand U21842 (N_21842,N_21675,N_21575);
or U21843 (N_21843,N_21717,N_21504);
and U21844 (N_21844,N_21677,N_21714);
xor U21845 (N_21845,N_21513,N_21542);
xnor U21846 (N_21846,N_21525,N_21553);
nand U21847 (N_21847,N_21585,N_21719);
or U21848 (N_21848,N_21549,N_21616);
nand U21849 (N_21849,N_21653,N_21534);
xor U21850 (N_21850,N_21548,N_21524);
and U21851 (N_21851,N_21591,N_21658);
nand U21852 (N_21852,N_21562,N_21748);
xor U21853 (N_21853,N_21503,N_21682);
and U21854 (N_21854,N_21506,N_21581);
or U21855 (N_21855,N_21565,N_21587);
or U21856 (N_21856,N_21700,N_21690);
or U21857 (N_21857,N_21623,N_21741);
or U21858 (N_21858,N_21723,N_21552);
xnor U21859 (N_21859,N_21578,N_21608);
or U21860 (N_21860,N_21632,N_21535);
nor U21861 (N_21861,N_21649,N_21699);
or U21862 (N_21862,N_21510,N_21724);
and U21863 (N_21863,N_21580,N_21576);
nor U21864 (N_21864,N_21738,N_21740);
and U21865 (N_21865,N_21648,N_21561);
and U21866 (N_21866,N_21590,N_21720);
nor U21867 (N_21867,N_21588,N_21745);
or U21868 (N_21868,N_21663,N_21698);
nand U21869 (N_21869,N_21539,N_21639);
nor U21870 (N_21870,N_21635,N_21611);
xnor U21871 (N_21871,N_21624,N_21502);
xor U21872 (N_21872,N_21613,N_21705);
or U21873 (N_21873,N_21589,N_21664);
and U21874 (N_21874,N_21643,N_21557);
xor U21875 (N_21875,N_21601,N_21529);
and U21876 (N_21876,N_21528,N_21610);
and U21877 (N_21877,N_21638,N_21654);
or U21878 (N_21878,N_21570,N_21719);
or U21879 (N_21879,N_21550,N_21505);
nand U21880 (N_21880,N_21591,N_21551);
or U21881 (N_21881,N_21723,N_21566);
nor U21882 (N_21882,N_21660,N_21519);
and U21883 (N_21883,N_21553,N_21686);
or U21884 (N_21884,N_21740,N_21522);
xnor U21885 (N_21885,N_21703,N_21637);
nor U21886 (N_21886,N_21500,N_21517);
or U21887 (N_21887,N_21569,N_21533);
and U21888 (N_21888,N_21594,N_21507);
and U21889 (N_21889,N_21525,N_21740);
or U21890 (N_21890,N_21539,N_21614);
and U21891 (N_21891,N_21626,N_21513);
and U21892 (N_21892,N_21653,N_21714);
xor U21893 (N_21893,N_21634,N_21553);
and U21894 (N_21894,N_21637,N_21691);
or U21895 (N_21895,N_21729,N_21703);
xnor U21896 (N_21896,N_21689,N_21514);
xnor U21897 (N_21897,N_21541,N_21628);
or U21898 (N_21898,N_21548,N_21690);
nor U21899 (N_21899,N_21514,N_21665);
nor U21900 (N_21900,N_21701,N_21697);
xor U21901 (N_21901,N_21566,N_21561);
xnor U21902 (N_21902,N_21678,N_21670);
nor U21903 (N_21903,N_21590,N_21664);
or U21904 (N_21904,N_21658,N_21527);
or U21905 (N_21905,N_21610,N_21616);
and U21906 (N_21906,N_21611,N_21515);
and U21907 (N_21907,N_21745,N_21637);
nor U21908 (N_21908,N_21670,N_21660);
nand U21909 (N_21909,N_21539,N_21599);
nand U21910 (N_21910,N_21543,N_21652);
and U21911 (N_21911,N_21704,N_21711);
and U21912 (N_21912,N_21663,N_21658);
or U21913 (N_21913,N_21736,N_21551);
nor U21914 (N_21914,N_21529,N_21737);
xor U21915 (N_21915,N_21524,N_21551);
nor U21916 (N_21916,N_21500,N_21575);
nor U21917 (N_21917,N_21646,N_21519);
and U21918 (N_21918,N_21712,N_21532);
nand U21919 (N_21919,N_21539,N_21709);
nand U21920 (N_21920,N_21510,N_21549);
nor U21921 (N_21921,N_21561,N_21700);
nor U21922 (N_21922,N_21722,N_21515);
or U21923 (N_21923,N_21593,N_21746);
and U21924 (N_21924,N_21577,N_21734);
xnor U21925 (N_21925,N_21581,N_21735);
nand U21926 (N_21926,N_21703,N_21573);
nor U21927 (N_21927,N_21565,N_21548);
nand U21928 (N_21928,N_21651,N_21696);
xor U21929 (N_21929,N_21746,N_21658);
and U21930 (N_21930,N_21628,N_21731);
xor U21931 (N_21931,N_21610,N_21602);
and U21932 (N_21932,N_21531,N_21748);
and U21933 (N_21933,N_21684,N_21688);
and U21934 (N_21934,N_21717,N_21626);
nand U21935 (N_21935,N_21636,N_21679);
or U21936 (N_21936,N_21725,N_21717);
nor U21937 (N_21937,N_21668,N_21505);
or U21938 (N_21938,N_21738,N_21642);
and U21939 (N_21939,N_21651,N_21653);
or U21940 (N_21940,N_21725,N_21671);
nor U21941 (N_21941,N_21524,N_21645);
xor U21942 (N_21942,N_21718,N_21582);
xor U21943 (N_21943,N_21740,N_21574);
nor U21944 (N_21944,N_21621,N_21571);
and U21945 (N_21945,N_21602,N_21725);
nor U21946 (N_21946,N_21676,N_21525);
nand U21947 (N_21947,N_21533,N_21546);
nor U21948 (N_21948,N_21627,N_21661);
xnor U21949 (N_21949,N_21662,N_21696);
and U21950 (N_21950,N_21737,N_21724);
xnor U21951 (N_21951,N_21517,N_21616);
nor U21952 (N_21952,N_21543,N_21584);
xnor U21953 (N_21953,N_21517,N_21533);
nand U21954 (N_21954,N_21682,N_21593);
nor U21955 (N_21955,N_21594,N_21662);
nand U21956 (N_21956,N_21573,N_21676);
nor U21957 (N_21957,N_21511,N_21740);
nor U21958 (N_21958,N_21513,N_21514);
xnor U21959 (N_21959,N_21564,N_21659);
xnor U21960 (N_21960,N_21504,N_21651);
nor U21961 (N_21961,N_21736,N_21561);
or U21962 (N_21962,N_21667,N_21614);
xnor U21963 (N_21963,N_21501,N_21657);
and U21964 (N_21964,N_21558,N_21745);
and U21965 (N_21965,N_21609,N_21634);
or U21966 (N_21966,N_21563,N_21624);
nand U21967 (N_21967,N_21521,N_21720);
nor U21968 (N_21968,N_21673,N_21653);
xnor U21969 (N_21969,N_21744,N_21647);
nor U21970 (N_21970,N_21572,N_21722);
xnor U21971 (N_21971,N_21600,N_21571);
and U21972 (N_21972,N_21624,N_21732);
nor U21973 (N_21973,N_21617,N_21555);
and U21974 (N_21974,N_21647,N_21522);
nor U21975 (N_21975,N_21577,N_21726);
nand U21976 (N_21976,N_21679,N_21563);
or U21977 (N_21977,N_21526,N_21747);
or U21978 (N_21978,N_21506,N_21583);
xor U21979 (N_21979,N_21558,N_21555);
xnor U21980 (N_21980,N_21658,N_21563);
and U21981 (N_21981,N_21587,N_21548);
and U21982 (N_21982,N_21679,N_21613);
nand U21983 (N_21983,N_21500,N_21610);
nor U21984 (N_21984,N_21684,N_21673);
and U21985 (N_21985,N_21698,N_21740);
nor U21986 (N_21986,N_21642,N_21650);
or U21987 (N_21987,N_21735,N_21505);
nand U21988 (N_21988,N_21665,N_21502);
nand U21989 (N_21989,N_21592,N_21576);
nor U21990 (N_21990,N_21647,N_21598);
or U21991 (N_21991,N_21625,N_21716);
and U21992 (N_21992,N_21715,N_21662);
and U21993 (N_21993,N_21725,N_21542);
or U21994 (N_21994,N_21640,N_21654);
and U21995 (N_21995,N_21558,N_21722);
nor U21996 (N_21996,N_21735,N_21716);
or U21997 (N_21997,N_21630,N_21535);
xor U21998 (N_21998,N_21695,N_21549);
xnor U21999 (N_21999,N_21644,N_21551);
and U22000 (N_22000,N_21888,N_21892);
xnor U22001 (N_22001,N_21899,N_21920);
and U22002 (N_22002,N_21806,N_21994);
nor U22003 (N_22003,N_21857,N_21969);
or U22004 (N_22004,N_21757,N_21887);
or U22005 (N_22005,N_21764,N_21786);
and U22006 (N_22006,N_21964,N_21762);
nand U22007 (N_22007,N_21987,N_21914);
nand U22008 (N_22008,N_21946,N_21897);
xnor U22009 (N_22009,N_21944,N_21945);
or U22010 (N_22010,N_21922,N_21751);
xor U22011 (N_22011,N_21942,N_21816);
and U22012 (N_22012,N_21884,N_21877);
or U22013 (N_22013,N_21825,N_21872);
nand U22014 (N_22014,N_21807,N_21900);
nor U22015 (N_22015,N_21866,N_21931);
or U22016 (N_22016,N_21809,N_21896);
or U22017 (N_22017,N_21775,N_21752);
and U22018 (N_22018,N_21871,N_21779);
or U22019 (N_22019,N_21902,N_21859);
nor U22020 (N_22020,N_21916,N_21975);
nor U22021 (N_22021,N_21974,N_21928);
xor U22022 (N_22022,N_21901,N_21970);
and U22023 (N_22023,N_21958,N_21771);
xnor U22024 (N_22024,N_21878,N_21938);
or U22025 (N_22025,N_21956,N_21962);
and U22026 (N_22026,N_21939,N_21963);
and U22027 (N_22027,N_21924,N_21915);
nand U22028 (N_22028,N_21820,N_21972);
or U22029 (N_22029,N_21908,N_21790);
and U22030 (N_22030,N_21918,N_21991);
nand U22031 (N_22031,N_21907,N_21805);
and U22032 (N_22032,N_21849,N_21865);
nand U22033 (N_22033,N_21980,N_21829);
nand U22034 (N_22034,N_21812,N_21833);
nor U22035 (N_22035,N_21759,N_21983);
and U22036 (N_22036,N_21875,N_21986);
and U22037 (N_22037,N_21995,N_21836);
nand U22038 (N_22038,N_21799,N_21760);
xnor U22039 (N_22039,N_21832,N_21934);
nor U22040 (N_22040,N_21834,N_21977);
xor U22041 (N_22041,N_21870,N_21767);
xor U22042 (N_22042,N_21936,N_21784);
and U22043 (N_22043,N_21840,N_21971);
and U22044 (N_22044,N_21993,N_21772);
or U22045 (N_22045,N_21842,N_21848);
xnor U22046 (N_22046,N_21826,N_21860);
xnor U22047 (N_22047,N_21981,N_21881);
xnor U22048 (N_22048,N_21879,N_21948);
or U22049 (N_22049,N_21808,N_21800);
and U22050 (N_22050,N_21817,N_21804);
xnor U22051 (N_22051,N_21852,N_21932);
xnor U22052 (N_22052,N_21839,N_21856);
nand U22053 (N_22053,N_21750,N_21814);
nor U22054 (N_22054,N_21935,N_21927);
or U22055 (N_22055,N_21867,N_21973);
nor U22056 (N_22056,N_21874,N_21880);
nand U22057 (N_22057,N_21824,N_21998);
nand U22058 (N_22058,N_21855,N_21768);
nand U22059 (N_22059,N_21845,N_21844);
or U22060 (N_22060,N_21780,N_21929);
and U22061 (N_22061,N_21850,N_21827);
xor U22062 (N_22062,N_21992,N_21885);
and U22063 (N_22063,N_21894,N_21947);
nor U22064 (N_22064,N_21959,N_21838);
or U22065 (N_22065,N_21854,N_21803);
and U22066 (N_22066,N_21882,N_21841);
xor U22067 (N_22067,N_21996,N_21797);
xor U22068 (N_22068,N_21766,N_21796);
or U22069 (N_22069,N_21949,N_21802);
and U22070 (N_22070,N_21769,N_21773);
nor U22071 (N_22071,N_21837,N_21965);
nand U22072 (N_22072,N_21989,N_21821);
xor U22073 (N_22073,N_21940,N_21910);
nor U22074 (N_22074,N_21919,N_21777);
xor U22075 (N_22075,N_21781,N_21787);
nor U22076 (N_22076,N_21813,N_21776);
xor U22077 (N_22077,N_21861,N_21886);
nor U22078 (N_22078,N_21794,N_21990);
nor U22079 (N_22079,N_21765,N_21778);
nand U22080 (N_22080,N_21864,N_21761);
xnor U22081 (N_22081,N_21823,N_21831);
and U22082 (N_22082,N_21955,N_21869);
nand U22083 (N_22083,N_21984,N_21953);
and U22084 (N_22084,N_21951,N_21801);
nand U22085 (N_22085,N_21876,N_21952);
nand U22086 (N_22086,N_21795,N_21883);
xor U22087 (N_22087,N_21830,N_21782);
or U22088 (N_22088,N_21811,N_21997);
or U22089 (N_22089,N_21893,N_21933);
xnor U22090 (N_22090,N_21968,N_21793);
xor U22091 (N_22091,N_21906,N_21966);
xnor U22092 (N_22092,N_21976,N_21756);
or U22093 (N_22093,N_21754,N_21783);
nand U22094 (N_22094,N_21930,N_21758);
or U22095 (N_22095,N_21755,N_21898);
nor U22096 (N_22096,N_21985,N_21921);
nor U22097 (N_22097,N_21911,N_21815);
xor U22098 (N_22098,N_21789,N_21982);
nor U22099 (N_22099,N_21999,N_21873);
nor U22100 (N_22100,N_21913,N_21943);
nand U22101 (N_22101,N_21862,N_21822);
or U22102 (N_22102,N_21912,N_21858);
nand U22103 (N_22103,N_21903,N_21979);
and U22104 (N_22104,N_21863,N_21846);
and U22105 (N_22105,N_21798,N_21763);
and U22106 (N_22106,N_21791,N_21828);
xnor U22107 (N_22107,N_21835,N_21954);
xnor U22108 (N_22108,N_21917,N_21810);
xor U22109 (N_22109,N_21960,N_21978);
nand U22110 (N_22110,N_21853,N_21941);
nand U22111 (N_22111,N_21847,N_21891);
nand U22112 (N_22112,N_21753,N_21909);
xnor U22113 (N_22113,N_21785,N_21818);
nor U22114 (N_22114,N_21843,N_21890);
xnor U22115 (N_22115,N_21895,N_21788);
xor U22116 (N_22116,N_21957,N_21961);
and U22117 (N_22117,N_21950,N_21792);
nand U22118 (N_22118,N_21988,N_21889);
nor U22119 (N_22119,N_21770,N_21923);
nor U22120 (N_22120,N_21925,N_21851);
xnor U22121 (N_22121,N_21904,N_21926);
and U22122 (N_22122,N_21819,N_21967);
or U22123 (N_22123,N_21937,N_21774);
and U22124 (N_22124,N_21905,N_21868);
nor U22125 (N_22125,N_21969,N_21817);
or U22126 (N_22126,N_21912,N_21822);
or U22127 (N_22127,N_21901,N_21884);
and U22128 (N_22128,N_21841,N_21870);
and U22129 (N_22129,N_21999,N_21987);
or U22130 (N_22130,N_21919,N_21924);
or U22131 (N_22131,N_21786,N_21755);
or U22132 (N_22132,N_21938,N_21884);
xor U22133 (N_22133,N_21999,N_21976);
or U22134 (N_22134,N_21857,N_21772);
nor U22135 (N_22135,N_21977,N_21960);
xnor U22136 (N_22136,N_21782,N_21799);
and U22137 (N_22137,N_21820,N_21919);
and U22138 (N_22138,N_21952,N_21961);
nor U22139 (N_22139,N_21797,N_21873);
nor U22140 (N_22140,N_21937,N_21930);
nand U22141 (N_22141,N_21779,N_21981);
or U22142 (N_22142,N_21827,N_21807);
nand U22143 (N_22143,N_21989,N_21757);
or U22144 (N_22144,N_21973,N_21813);
nand U22145 (N_22145,N_21756,N_21890);
and U22146 (N_22146,N_21825,N_21953);
nor U22147 (N_22147,N_21877,N_21958);
xnor U22148 (N_22148,N_21819,N_21771);
and U22149 (N_22149,N_21752,N_21801);
nand U22150 (N_22150,N_21863,N_21917);
xor U22151 (N_22151,N_21754,N_21799);
xor U22152 (N_22152,N_21815,N_21949);
or U22153 (N_22153,N_21993,N_21903);
xnor U22154 (N_22154,N_21974,N_21966);
nor U22155 (N_22155,N_21844,N_21864);
and U22156 (N_22156,N_21806,N_21825);
nor U22157 (N_22157,N_21949,N_21805);
nand U22158 (N_22158,N_21894,N_21811);
nand U22159 (N_22159,N_21942,N_21982);
nand U22160 (N_22160,N_21972,N_21841);
or U22161 (N_22161,N_21807,N_21803);
or U22162 (N_22162,N_21757,N_21980);
nor U22163 (N_22163,N_21800,N_21926);
xnor U22164 (N_22164,N_21916,N_21974);
and U22165 (N_22165,N_21919,N_21947);
nor U22166 (N_22166,N_21847,N_21856);
xnor U22167 (N_22167,N_21988,N_21837);
xnor U22168 (N_22168,N_21764,N_21929);
nand U22169 (N_22169,N_21993,N_21760);
nor U22170 (N_22170,N_21995,N_21936);
or U22171 (N_22171,N_21929,N_21804);
or U22172 (N_22172,N_21908,N_21832);
nand U22173 (N_22173,N_21887,N_21980);
nor U22174 (N_22174,N_21807,N_21850);
nand U22175 (N_22175,N_21818,N_21918);
xnor U22176 (N_22176,N_21914,N_21926);
nor U22177 (N_22177,N_21953,N_21778);
nor U22178 (N_22178,N_21807,N_21928);
nor U22179 (N_22179,N_21810,N_21841);
xor U22180 (N_22180,N_21810,N_21865);
xnor U22181 (N_22181,N_21863,N_21924);
and U22182 (N_22182,N_21816,N_21772);
nand U22183 (N_22183,N_21805,N_21789);
and U22184 (N_22184,N_21756,N_21848);
and U22185 (N_22185,N_21857,N_21811);
nand U22186 (N_22186,N_21953,N_21990);
or U22187 (N_22187,N_21782,N_21775);
nor U22188 (N_22188,N_21835,N_21974);
nor U22189 (N_22189,N_21855,N_21888);
nand U22190 (N_22190,N_21884,N_21939);
and U22191 (N_22191,N_21816,N_21976);
nand U22192 (N_22192,N_21918,N_21910);
nor U22193 (N_22193,N_21971,N_21918);
and U22194 (N_22194,N_21804,N_21921);
xnor U22195 (N_22195,N_21850,N_21935);
xor U22196 (N_22196,N_21956,N_21948);
or U22197 (N_22197,N_21834,N_21825);
nor U22198 (N_22198,N_21986,N_21959);
nand U22199 (N_22199,N_21972,N_21908);
and U22200 (N_22200,N_21905,N_21854);
nor U22201 (N_22201,N_21918,N_21878);
and U22202 (N_22202,N_21951,N_21784);
and U22203 (N_22203,N_21973,N_21901);
xor U22204 (N_22204,N_21860,N_21975);
nor U22205 (N_22205,N_21805,N_21892);
and U22206 (N_22206,N_21852,N_21817);
nor U22207 (N_22207,N_21878,N_21788);
nor U22208 (N_22208,N_21802,N_21848);
or U22209 (N_22209,N_21972,N_21986);
or U22210 (N_22210,N_21857,N_21956);
or U22211 (N_22211,N_21921,N_21772);
xor U22212 (N_22212,N_21902,N_21847);
nor U22213 (N_22213,N_21964,N_21818);
and U22214 (N_22214,N_21843,N_21829);
or U22215 (N_22215,N_21935,N_21986);
nor U22216 (N_22216,N_21928,N_21893);
or U22217 (N_22217,N_21916,N_21810);
or U22218 (N_22218,N_21896,N_21838);
nor U22219 (N_22219,N_21906,N_21858);
nand U22220 (N_22220,N_21979,N_21860);
nor U22221 (N_22221,N_21960,N_21955);
or U22222 (N_22222,N_21799,N_21807);
nor U22223 (N_22223,N_21987,N_21822);
nand U22224 (N_22224,N_21925,N_21832);
nand U22225 (N_22225,N_21942,N_21779);
nand U22226 (N_22226,N_21973,N_21866);
xor U22227 (N_22227,N_21983,N_21755);
and U22228 (N_22228,N_21812,N_21978);
nor U22229 (N_22229,N_21939,N_21971);
xnor U22230 (N_22230,N_21814,N_21930);
nand U22231 (N_22231,N_21979,N_21823);
nor U22232 (N_22232,N_21948,N_21979);
nor U22233 (N_22233,N_21884,N_21935);
xnor U22234 (N_22234,N_21851,N_21908);
and U22235 (N_22235,N_21915,N_21809);
xnor U22236 (N_22236,N_21900,N_21975);
xor U22237 (N_22237,N_21875,N_21818);
nand U22238 (N_22238,N_21936,N_21762);
nand U22239 (N_22239,N_21803,N_21964);
nor U22240 (N_22240,N_21853,N_21953);
xor U22241 (N_22241,N_21914,N_21906);
nand U22242 (N_22242,N_21976,N_21750);
or U22243 (N_22243,N_21771,N_21917);
or U22244 (N_22244,N_21860,N_21837);
xor U22245 (N_22245,N_21971,N_21848);
or U22246 (N_22246,N_21813,N_21881);
xor U22247 (N_22247,N_21773,N_21982);
xor U22248 (N_22248,N_21829,N_21987);
or U22249 (N_22249,N_21998,N_21910);
nor U22250 (N_22250,N_22165,N_22217);
or U22251 (N_22251,N_22208,N_22057);
xnor U22252 (N_22252,N_22173,N_22187);
and U22253 (N_22253,N_22190,N_22064);
xor U22254 (N_22254,N_22119,N_22035);
or U22255 (N_22255,N_22195,N_22104);
nand U22256 (N_22256,N_22101,N_22009);
nor U22257 (N_22257,N_22046,N_22180);
or U22258 (N_22258,N_22248,N_22003);
xor U22259 (N_22259,N_22047,N_22201);
xor U22260 (N_22260,N_22044,N_22055);
xnor U22261 (N_22261,N_22125,N_22108);
nor U22262 (N_22262,N_22154,N_22162);
nand U22263 (N_22263,N_22206,N_22218);
and U22264 (N_22264,N_22075,N_22139);
nor U22265 (N_22265,N_22028,N_22110);
xnor U22266 (N_22266,N_22065,N_22233);
nand U22267 (N_22267,N_22024,N_22086);
nand U22268 (N_22268,N_22213,N_22211);
and U22269 (N_22269,N_22242,N_22069);
and U22270 (N_22270,N_22018,N_22023);
nor U22271 (N_22271,N_22156,N_22168);
nand U22272 (N_22272,N_22058,N_22192);
or U22273 (N_22273,N_22137,N_22060);
xnor U22274 (N_22274,N_22177,N_22151);
nand U22275 (N_22275,N_22198,N_22045);
nor U22276 (N_22276,N_22053,N_22080);
nand U22277 (N_22277,N_22091,N_22226);
or U22278 (N_22278,N_22088,N_22081);
and U22279 (N_22279,N_22048,N_22114);
or U22280 (N_22280,N_22234,N_22004);
and U22281 (N_22281,N_22246,N_22228);
nor U22282 (N_22282,N_22161,N_22116);
nor U22283 (N_22283,N_22202,N_22050);
nor U22284 (N_22284,N_22230,N_22209);
xnor U22285 (N_22285,N_22164,N_22025);
and U22286 (N_22286,N_22127,N_22207);
xnor U22287 (N_22287,N_22094,N_22016);
nand U22288 (N_22288,N_22068,N_22073);
and U22289 (N_22289,N_22186,N_22197);
or U22290 (N_22290,N_22030,N_22232);
nor U22291 (N_22291,N_22077,N_22227);
or U22292 (N_22292,N_22184,N_22189);
nor U22293 (N_22293,N_22015,N_22146);
or U22294 (N_22294,N_22049,N_22224);
or U22295 (N_22295,N_22097,N_22111);
xor U22296 (N_22296,N_22200,N_22089);
nand U22297 (N_22297,N_22033,N_22013);
xor U22298 (N_22298,N_22056,N_22196);
nor U22299 (N_22299,N_22054,N_22225);
and U22300 (N_22300,N_22229,N_22038);
nor U22301 (N_22301,N_22012,N_22134);
or U22302 (N_22302,N_22221,N_22244);
nand U22303 (N_22303,N_22093,N_22002);
nor U22304 (N_22304,N_22131,N_22032);
xnor U22305 (N_22305,N_22092,N_22243);
xor U22306 (N_22306,N_22063,N_22102);
xor U22307 (N_22307,N_22193,N_22126);
xnor U22308 (N_22308,N_22084,N_22099);
or U22309 (N_22309,N_22214,N_22039);
and U22310 (N_22310,N_22183,N_22235);
and U22311 (N_22311,N_22090,N_22001);
and U22312 (N_22312,N_22174,N_22017);
and U22313 (N_22313,N_22117,N_22005);
nand U22314 (N_22314,N_22062,N_22239);
nor U22315 (N_22315,N_22199,N_22098);
nand U22316 (N_22316,N_22149,N_22113);
or U22317 (N_22317,N_22014,N_22059);
or U22318 (N_22318,N_22027,N_22191);
nand U22319 (N_22319,N_22115,N_22181);
xnor U22320 (N_22320,N_22067,N_22103);
and U22321 (N_22321,N_22170,N_22082);
or U22322 (N_22322,N_22140,N_22022);
xor U22323 (N_22323,N_22153,N_22241);
or U22324 (N_22324,N_22167,N_22031);
or U22325 (N_22325,N_22085,N_22122);
and U22326 (N_22326,N_22194,N_22247);
and U22327 (N_22327,N_22128,N_22188);
and U22328 (N_22328,N_22236,N_22071);
nand U22329 (N_22329,N_22147,N_22155);
nor U22330 (N_22330,N_22141,N_22112);
or U22331 (N_22331,N_22096,N_22204);
or U22332 (N_22332,N_22036,N_22124);
xnor U22333 (N_22333,N_22223,N_22105);
and U22334 (N_22334,N_22210,N_22171);
xnor U22335 (N_22335,N_22135,N_22034);
and U22336 (N_22336,N_22106,N_22220);
xor U22337 (N_22337,N_22160,N_22176);
xnor U22338 (N_22338,N_22219,N_22172);
or U22339 (N_22339,N_22007,N_22182);
and U22340 (N_22340,N_22152,N_22240);
nor U22341 (N_22341,N_22169,N_22010);
and U22342 (N_22342,N_22043,N_22166);
nand U22343 (N_22343,N_22066,N_22150);
nand U22344 (N_22344,N_22132,N_22205);
and U22345 (N_22345,N_22136,N_22040);
or U22346 (N_22346,N_22185,N_22238);
and U22347 (N_22347,N_22087,N_22051);
xnor U22348 (N_22348,N_22006,N_22212);
and U22349 (N_22349,N_22011,N_22061);
or U22350 (N_22350,N_22138,N_22245);
nor U22351 (N_22351,N_22179,N_22079);
nand U22352 (N_22352,N_22123,N_22095);
nand U22353 (N_22353,N_22020,N_22109);
nor U22354 (N_22354,N_22158,N_22121);
and U22355 (N_22355,N_22000,N_22107);
xor U22356 (N_22356,N_22144,N_22072);
nand U22357 (N_22357,N_22019,N_22129);
and U22358 (N_22358,N_22052,N_22120);
xnor U22359 (N_22359,N_22157,N_22175);
xor U22360 (N_22360,N_22100,N_22078);
and U22361 (N_22361,N_22130,N_22008);
and U22362 (N_22362,N_22021,N_22026);
xor U22363 (N_22363,N_22042,N_22074);
nor U22364 (N_22364,N_22037,N_22178);
nor U22365 (N_22365,N_22145,N_22237);
and U22366 (N_22366,N_22249,N_22029);
or U22367 (N_22367,N_22222,N_22159);
xor U22368 (N_22368,N_22070,N_22041);
or U22369 (N_22369,N_22143,N_22133);
nor U22370 (N_22370,N_22083,N_22142);
and U22371 (N_22371,N_22148,N_22231);
nor U22372 (N_22372,N_22076,N_22118);
nor U22373 (N_22373,N_22203,N_22216);
xor U22374 (N_22374,N_22163,N_22215);
or U22375 (N_22375,N_22006,N_22020);
nor U22376 (N_22376,N_22239,N_22054);
xnor U22377 (N_22377,N_22216,N_22108);
nor U22378 (N_22378,N_22235,N_22223);
xor U22379 (N_22379,N_22012,N_22148);
or U22380 (N_22380,N_22036,N_22077);
nand U22381 (N_22381,N_22060,N_22029);
and U22382 (N_22382,N_22165,N_22132);
and U22383 (N_22383,N_22059,N_22147);
and U22384 (N_22384,N_22034,N_22117);
or U22385 (N_22385,N_22207,N_22099);
nand U22386 (N_22386,N_22008,N_22058);
or U22387 (N_22387,N_22169,N_22192);
xor U22388 (N_22388,N_22058,N_22024);
or U22389 (N_22389,N_22046,N_22191);
xor U22390 (N_22390,N_22246,N_22123);
or U22391 (N_22391,N_22050,N_22089);
nand U22392 (N_22392,N_22170,N_22199);
and U22393 (N_22393,N_22140,N_22246);
nand U22394 (N_22394,N_22031,N_22142);
xor U22395 (N_22395,N_22140,N_22194);
xnor U22396 (N_22396,N_22153,N_22231);
and U22397 (N_22397,N_22119,N_22158);
or U22398 (N_22398,N_22117,N_22171);
and U22399 (N_22399,N_22086,N_22081);
nand U22400 (N_22400,N_22040,N_22246);
nand U22401 (N_22401,N_22055,N_22140);
nand U22402 (N_22402,N_22173,N_22018);
xnor U22403 (N_22403,N_22236,N_22168);
xnor U22404 (N_22404,N_22140,N_22174);
xor U22405 (N_22405,N_22032,N_22050);
and U22406 (N_22406,N_22206,N_22045);
xor U22407 (N_22407,N_22137,N_22113);
nand U22408 (N_22408,N_22068,N_22192);
xnor U22409 (N_22409,N_22137,N_22182);
nand U22410 (N_22410,N_22212,N_22136);
and U22411 (N_22411,N_22097,N_22070);
nor U22412 (N_22412,N_22210,N_22162);
nor U22413 (N_22413,N_22031,N_22067);
or U22414 (N_22414,N_22040,N_22209);
and U22415 (N_22415,N_22065,N_22080);
nand U22416 (N_22416,N_22033,N_22004);
nand U22417 (N_22417,N_22148,N_22110);
xnor U22418 (N_22418,N_22165,N_22023);
nand U22419 (N_22419,N_22197,N_22102);
nor U22420 (N_22420,N_22156,N_22006);
or U22421 (N_22421,N_22192,N_22189);
and U22422 (N_22422,N_22072,N_22215);
nand U22423 (N_22423,N_22230,N_22155);
nor U22424 (N_22424,N_22227,N_22159);
xor U22425 (N_22425,N_22010,N_22062);
nand U22426 (N_22426,N_22091,N_22156);
or U22427 (N_22427,N_22226,N_22077);
nor U22428 (N_22428,N_22185,N_22158);
or U22429 (N_22429,N_22149,N_22125);
and U22430 (N_22430,N_22120,N_22014);
nor U22431 (N_22431,N_22027,N_22015);
and U22432 (N_22432,N_22077,N_22082);
nand U22433 (N_22433,N_22185,N_22107);
nor U22434 (N_22434,N_22006,N_22077);
nor U22435 (N_22435,N_22076,N_22244);
xnor U22436 (N_22436,N_22068,N_22131);
nor U22437 (N_22437,N_22028,N_22179);
nand U22438 (N_22438,N_22240,N_22049);
nand U22439 (N_22439,N_22234,N_22195);
xnor U22440 (N_22440,N_22222,N_22120);
nor U22441 (N_22441,N_22119,N_22224);
xnor U22442 (N_22442,N_22069,N_22112);
nor U22443 (N_22443,N_22101,N_22151);
nor U22444 (N_22444,N_22230,N_22170);
and U22445 (N_22445,N_22136,N_22054);
xor U22446 (N_22446,N_22176,N_22212);
nor U22447 (N_22447,N_22234,N_22089);
xor U22448 (N_22448,N_22101,N_22232);
xor U22449 (N_22449,N_22161,N_22124);
nand U22450 (N_22450,N_22043,N_22002);
or U22451 (N_22451,N_22179,N_22091);
and U22452 (N_22452,N_22034,N_22160);
or U22453 (N_22453,N_22063,N_22147);
or U22454 (N_22454,N_22116,N_22145);
or U22455 (N_22455,N_22097,N_22081);
or U22456 (N_22456,N_22191,N_22177);
nand U22457 (N_22457,N_22078,N_22000);
and U22458 (N_22458,N_22202,N_22203);
nor U22459 (N_22459,N_22117,N_22212);
nand U22460 (N_22460,N_22170,N_22212);
xnor U22461 (N_22461,N_22205,N_22092);
nand U22462 (N_22462,N_22048,N_22054);
and U22463 (N_22463,N_22165,N_22233);
nor U22464 (N_22464,N_22044,N_22093);
nor U22465 (N_22465,N_22032,N_22207);
xnor U22466 (N_22466,N_22122,N_22112);
or U22467 (N_22467,N_22026,N_22133);
xnor U22468 (N_22468,N_22159,N_22204);
xor U22469 (N_22469,N_22036,N_22001);
and U22470 (N_22470,N_22026,N_22027);
nand U22471 (N_22471,N_22142,N_22155);
or U22472 (N_22472,N_22140,N_22227);
and U22473 (N_22473,N_22234,N_22010);
nor U22474 (N_22474,N_22217,N_22109);
nor U22475 (N_22475,N_22118,N_22147);
nor U22476 (N_22476,N_22189,N_22146);
nor U22477 (N_22477,N_22098,N_22200);
nor U22478 (N_22478,N_22079,N_22163);
nand U22479 (N_22479,N_22140,N_22080);
and U22480 (N_22480,N_22002,N_22216);
and U22481 (N_22481,N_22061,N_22047);
or U22482 (N_22482,N_22051,N_22015);
or U22483 (N_22483,N_22218,N_22115);
nor U22484 (N_22484,N_22046,N_22094);
nand U22485 (N_22485,N_22085,N_22158);
or U22486 (N_22486,N_22036,N_22175);
nand U22487 (N_22487,N_22181,N_22229);
xor U22488 (N_22488,N_22124,N_22080);
xor U22489 (N_22489,N_22086,N_22080);
nor U22490 (N_22490,N_22117,N_22151);
xnor U22491 (N_22491,N_22193,N_22008);
and U22492 (N_22492,N_22162,N_22104);
xnor U22493 (N_22493,N_22178,N_22068);
xnor U22494 (N_22494,N_22215,N_22070);
or U22495 (N_22495,N_22004,N_22158);
nor U22496 (N_22496,N_22033,N_22131);
or U22497 (N_22497,N_22140,N_22167);
and U22498 (N_22498,N_22059,N_22213);
xor U22499 (N_22499,N_22049,N_22025);
xnor U22500 (N_22500,N_22452,N_22308);
and U22501 (N_22501,N_22437,N_22319);
nand U22502 (N_22502,N_22335,N_22315);
and U22503 (N_22503,N_22374,N_22286);
nor U22504 (N_22504,N_22403,N_22376);
nor U22505 (N_22505,N_22334,N_22389);
or U22506 (N_22506,N_22326,N_22343);
and U22507 (N_22507,N_22383,N_22401);
xor U22508 (N_22508,N_22378,N_22350);
and U22509 (N_22509,N_22283,N_22414);
nand U22510 (N_22510,N_22313,N_22311);
or U22511 (N_22511,N_22348,N_22304);
nor U22512 (N_22512,N_22475,N_22309);
xnor U22513 (N_22513,N_22296,N_22418);
nor U22514 (N_22514,N_22497,N_22337);
and U22515 (N_22515,N_22275,N_22307);
xnor U22516 (N_22516,N_22386,N_22458);
nor U22517 (N_22517,N_22290,N_22456);
nand U22518 (N_22518,N_22448,N_22255);
nor U22519 (N_22519,N_22372,N_22453);
nor U22520 (N_22520,N_22382,N_22274);
and U22521 (N_22521,N_22263,N_22393);
or U22522 (N_22522,N_22384,N_22366);
xnor U22523 (N_22523,N_22292,N_22422);
or U22524 (N_22524,N_22446,N_22339);
xnor U22525 (N_22525,N_22294,N_22287);
nand U22526 (N_22526,N_22415,N_22471);
nor U22527 (N_22527,N_22492,N_22370);
and U22528 (N_22528,N_22430,N_22439);
nand U22529 (N_22529,N_22289,N_22268);
nand U22530 (N_22530,N_22302,N_22429);
nand U22531 (N_22531,N_22481,N_22441);
nor U22532 (N_22532,N_22327,N_22493);
nor U22533 (N_22533,N_22463,N_22431);
nor U22534 (N_22534,N_22428,N_22336);
nand U22535 (N_22535,N_22388,N_22465);
xor U22536 (N_22536,N_22312,N_22279);
xor U22537 (N_22537,N_22257,N_22434);
and U22538 (N_22538,N_22278,N_22300);
or U22539 (N_22539,N_22375,N_22398);
nor U22540 (N_22540,N_22342,N_22485);
xnor U22541 (N_22541,N_22489,N_22399);
xor U22542 (N_22542,N_22272,N_22484);
or U22543 (N_22543,N_22397,N_22277);
nand U22544 (N_22544,N_22261,N_22267);
nor U22545 (N_22545,N_22461,N_22297);
xnor U22546 (N_22546,N_22394,N_22498);
or U22547 (N_22547,N_22412,N_22328);
xor U22548 (N_22548,N_22488,N_22347);
xor U22549 (N_22549,N_22251,N_22436);
or U22550 (N_22550,N_22404,N_22365);
xor U22551 (N_22551,N_22285,N_22413);
or U22552 (N_22552,N_22454,N_22340);
nor U22553 (N_22553,N_22432,N_22468);
nand U22554 (N_22554,N_22466,N_22318);
and U22555 (N_22555,N_22258,N_22259);
or U22556 (N_22556,N_22387,N_22361);
nor U22557 (N_22557,N_22435,N_22469);
or U22558 (N_22558,N_22360,N_22368);
nor U22559 (N_22559,N_22421,N_22451);
or U22560 (N_22560,N_22495,N_22345);
and U22561 (N_22561,N_22464,N_22472);
nor U22562 (N_22562,N_22344,N_22496);
and U22563 (N_22563,N_22280,N_22320);
xor U22564 (N_22564,N_22351,N_22322);
xnor U22565 (N_22565,N_22379,N_22395);
nor U22566 (N_22566,N_22396,N_22442);
xnor U22567 (N_22567,N_22349,N_22305);
or U22568 (N_22568,N_22405,N_22253);
xnor U22569 (N_22569,N_22447,N_22491);
nand U22570 (N_22570,N_22459,N_22332);
nor U22571 (N_22571,N_22407,N_22377);
xnor U22572 (N_22572,N_22449,N_22476);
nand U22573 (N_22573,N_22482,N_22462);
or U22574 (N_22574,N_22353,N_22420);
and U22575 (N_22575,N_22254,N_22390);
or U22576 (N_22576,N_22474,N_22486);
nand U22577 (N_22577,N_22444,N_22250);
nor U22578 (N_22578,N_22324,N_22298);
or U22579 (N_22579,N_22381,N_22359);
or U22580 (N_22580,N_22310,N_22271);
nor U22581 (N_22581,N_22358,N_22262);
nor U22582 (N_22582,N_22288,N_22424);
nand U22583 (N_22583,N_22417,N_22355);
or U22584 (N_22584,N_22356,N_22291);
xnor U22585 (N_22585,N_22426,N_22467);
and U22586 (N_22586,N_22338,N_22252);
nor U22587 (N_22587,N_22427,N_22385);
and U22588 (N_22588,N_22457,N_22478);
nand U22589 (N_22589,N_22443,N_22293);
xor U22590 (N_22590,N_22281,N_22408);
xor U22591 (N_22591,N_22490,N_22406);
and U22592 (N_22592,N_22265,N_22410);
xnor U22593 (N_22593,N_22364,N_22367);
xor U22594 (N_22594,N_22301,N_22477);
and U22595 (N_22595,N_22316,N_22499);
and U22596 (N_22596,N_22380,N_22330);
and U22597 (N_22597,N_22419,N_22480);
or U22598 (N_22598,N_22479,N_22440);
nor U22599 (N_22599,N_22346,N_22314);
nor U22600 (N_22600,N_22303,N_22341);
xnor U22601 (N_22601,N_22282,N_22362);
or U22602 (N_22602,N_22483,N_22276);
or U22603 (N_22603,N_22357,N_22306);
and U22604 (N_22604,N_22295,N_22354);
or U22605 (N_22605,N_22392,N_22450);
nand U22606 (N_22606,N_22445,N_22487);
xor U22607 (N_22607,N_22363,N_22331);
and U22608 (N_22608,N_22371,N_22317);
and U22609 (N_22609,N_22473,N_22409);
nand U22610 (N_22610,N_22352,N_22270);
or U22611 (N_22611,N_22256,N_22460);
nand U22612 (N_22612,N_22438,N_22269);
xnor U22613 (N_22613,N_22369,N_22494);
and U22614 (N_22614,N_22373,N_22273);
or U22615 (N_22615,N_22455,N_22416);
nand U22616 (N_22616,N_22323,N_22266);
nand U22617 (N_22617,N_22425,N_22433);
nand U22618 (N_22618,N_22411,N_22321);
nor U22619 (N_22619,N_22284,N_22470);
and U22620 (N_22620,N_22325,N_22260);
nor U22621 (N_22621,N_22423,N_22400);
or U22622 (N_22622,N_22264,N_22299);
nor U22623 (N_22623,N_22391,N_22333);
nor U22624 (N_22624,N_22402,N_22329);
nand U22625 (N_22625,N_22485,N_22495);
nand U22626 (N_22626,N_22370,N_22261);
and U22627 (N_22627,N_22495,N_22396);
nand U22628 (N_22628,N_22260,N_22333);
nand U22629 (N_22629,N_22489,N_22265);
or U22630 (N_22630,N_22449,N_22306);
nand U22631 (N_22631,N_22491,N_22441);
and U22632 (N_22632,N_22445,N_22292);
xor U22633 (N_22633,N_22263,N_22271);
or U22634 (N_22634,N_22366,N_22282);
nand U22635 (N_22635,N_22453,N_22468);
nor U22636 (N_22636,N_22300,N_22389);
and U22637 (N_22637,N_22397,N_22404);
xor U22638 (N_22638,N_22431,N_22373);
and U22639 (N_22639,N_22291,N_22329);
or U22640 (N_22640,N_22250,N_22459);
or U22641 (N_22641,N_22254,N_22267);
and U22642 (N_22642,N_22374,N_22284);
xnor U22643 (N_22643,N_22370,N_22459);
nand U22644 (N_22644,N_22445,N_22369);
nor U22645 (N_22645,N_22453,N_22301);
or U22646 (N_22646,N_22290,N_22375);
nor U22647 (N_22647,N_22361,N_22424);
and U22648 (N_22648,N_22390,N_22283);
nand U22649 (N_22649,N_22406,N_22438);
xnor U22650 (N_22650,N_22390,N_22320);
nand U22651 (N_22651,N_22433,N_22415);
nor U22652 (N_22652,N_22288,N_22381);
nor U22653 (N_22653,N_22405,N_22384);
and U22654 (N_22654,N_22390,N_22340);
and U22655 (N_22655,N_22260,N_22309);
and U22656 (N_22656,N_22484,N_22294);
or U22657 (N_22657,N_22444,N_22309);
xor U22658 (N_22658,N_22380,N_22423);
xor U22659 (N_22659,N_22320,N_22423);
nor U22660 (N_22660,N_22488,N_22282);
and U22661 (N_22661,N_22275,N_22406);
nand U22662 (N_22662,N_22425,N_22317);
nand U22663 (N_22663,N_22435,N_22305);
nand U22664 (N_22664,N_22308,N_22433);
nor U22665 (N_22665,N_22267,N_22465);
or U22666 (N_22666,N_22385,N_22392);
nand U22667 (N_22667,N_22269,N_22251);
nor U22668 (N_22668,N_22438,N_22422);
or U22669 (N_22669,N_22494,N_22454);
nor U22670 (N_22670,N_22288,N_22435);
xnor U22671 (N_22671,N_22294,N_22302);
or U22672 (N_22672,N_22367,N_22415);
nand U22673 (N_22673,N_22265,N_22412);
nand U22674 (N_22674,N_22448,N_22427);
and U22675 (N_22675,N_22413,N_22408);
and U22676 (N_22676,N_22259,N_22255);
and U22677 (N_22677,N_22468,N_22295);
xor U22678 (N_22678,N_22318,N_22396);
xnor U22679 (N_22679,N_22461,N_22289);
and U22680 (N_22680,N_22386,N_22407);
or U22681 (N_22681,N_22308,N_22272);
nand U22682 (N_22682,N_22411,N_22469);
nor U22683 (N_22683,N_22309,N_22418);
xnor U22684 (N_22684,N_22408,N_22459);
nand U22685 (N_22685,N_22270,N_22408);
nor U22686 (N_22686,N_22337,N_22294);
xor U22687 (N_22687,N_22301,N_22459);
and U22688 (N_22688,N_22435,N_22486);
nand U22689 (N_22689,N_22260,N_22353);
nor U22690 (N_22690,N_22353,N_22443);
nand U22691 (N_22691,N_22486,N_22414);
xnor U22692 (N_22692,N_22359,N_22351);
nor U22693 (N_22693,N_22424,N_22488);
xnor U22694 (N_22694,N_22334,N_22463);
nand U22695 (N_22695,N_22423,N_22352);
and U22696 (N_22696,N_22354,N_22349);
nand U22697 (N_22697,N_22498,N_22263);
nand U22698 (N_22698,N_22478,N_22415);
and U22699 (N_22699,N_22278,N_22250);
nor U22700 (N_22700,N_22461,N_22346);
or U22701 (N_22701,N_22393,N_22431);
nand U22702 (N_22702,N_22277,N_22402);
xnor U22703 (N_22703,N_22381,N_22316);
and U22704 (N_22704,N_22282,N_22490);
xnor U22705 (N_22705,N_22332,N_22342);
and U22706 (N_22706,N_22388,N_22385);
xnor U22707 (N_22707,N_22331,N_22267);
or U22708 (N_22708,N_22284,N_22468);
nand U22709 (N_22709,N_22387,N_22311);
nor U22710 (N_22710,N_22306,N_22343);
or U22711 (N_22711,N_22262,N_22485);
xnor U22712 (N_22712,N_22329,N_22325);
or U22713 (N_22713,N_22402,N_22419);
nor U22714 (N_22714,N_22402,N_22317);
nor U22715 (N_22715,N_22268,N_22435);
or U22716 (N_22716,N_22261,N_22456);
or U22717 (N_22717,N_22279,N_22256);
and U22718 (N_22718,N_22437,N_22341);
and U22719 (N_22719,N_22272,N_22318);
xor U22720 (N_22720,N_22368,N_22471);
or U22721 (N_22721,N_22309,N_22479);
xor U22722 (N_22722,N_22259,N_22467);
or U22723 (N_22723,N_22282,N_22387);
nand U22724 (N_22724,N_22444,N_22386);
nand U22725 (N_22725,N_22392,N_22497);
and U22726 (N_22726,N_22470,N_22481);
xnor U22727 (N_22727,N_22322,N_22432);
xor U22728 (N_22728,N_22306,N_22398);
xnor U22729 (N_22729,N_22485,N_22411);
nand U22730 (N_22730,N_22321,N_22414);
and U22731 (N_22731,N_22269,N_22443);
xnor U22732 (N_22732,N_22424,N_22317);
and U22733 (N_22733,N_22410,N_22323);
nand U22734 (N_22734,N_22370,N_22382);
xor U22735 (N_22735,N_22434,N_22422);
nor U22736 (N_22736,N_22470,N_22283);
or U22737 (N_22737,N_22396,N_22430);
xnor U22738 (N_22738,N_22314,N_22452);
or U22739 (N_22739,N_22349,N_22304);
or U22740 (N_22740,N_22266,N_22398);
or U22741 (N_22741,N_22414,N_22344);
or U22742 (N_22742,N_22299,N_22477);
nand U22743 (N_22743,N_22387,N_22460);
and U22744 (N_22744,N_22480,N_22272);
or U22745 (N_22745,N_22263,N_22298);
nand U22746 (N_22746,N_22441,N_22404);
or U22747 (N_22747,N_22295,N_22266);
or U22748 (N_22748,N_22392,N_22458);
and U22749 (N_22749,N_22419,N_22477);
or U22750 (N_22750,N_22623,N_22724);
nand U22751 (N_22751,N_22590,N_22725);
or U22752 (N_22752,N_22529,N_22729);
and U22753 (N_22753,N_22710,N_22594);
and U22754 (N_22754,N_22514,N_22584);
and U22755 (N_22755,N_22622,N_22748);
nand U22756 (N_22756,N_22632,N_22631);
or U22757 (N_22757,N_22621,N_22721);
and U22758 (N_22758,N_22676,N_22624);
or U22759 (N_22759,N_22570,N_22741);
nor U22760 (N_22760,N_22677,N_22638);
or U22761 (N_22761,N_22599,N_22609);
nor U22762 (N_22762,N_22597,N_22591);
nand U22763 (N_22763,N_22668,N_22582);
or U22764 (N_22764,N_22617,N_22580);
and U22765 (N_22765,N_22626,N_22516);
and U22766 (N_22766,N_22685,N_22527);
or U22767 (N_22767,N_22512,N_22720);
nand U22768 (N_22768,N_22630,N_22726);
nand U22769 (N_22769,N_22505,N_22614);
nand U22770 (N_22770,N_22517,N_22712);
nand U22771 (N_22771,N_22523,N_22678);
and U22772 (N_22772,N_22501,N_22684);
xor U22773 (N_22773,N_22544,N_22589);
xnor U22774 (N_22774,N_22672,N_22603);
or U22775 (N_22775,N_22694,N_22716);
and U22776 (N_22776,N_22649,N_22522);
or U22777 (N_22777,N_22576,N_22616);
nand U22778 (N_22778,N_22502,N_22648);
nor U22779 (N_22779,N_22572,N_22690);
nand U22780 (N_22780,N_22722,N_22506);
nand U22781 (N_22781,N_22607,N_22604);
and U22782 (N_22782,N_22535,N_22679);
nor U22783 (N_22783,N_22697,N_22655);
xor U22784 (N_22784,N_22504,N_22541);
nand U22785 (N_22785,N_22733,N_22736);
xnor U22786 (N_22786,N_22521,N_22548);
nor U22787 (N_22787,N_22605,N_22565);
xnor U22788 (N_22788,N_22536,N_22513);
and U22789 (N_22789,N_22564,N_22593);
xor U22790 (N_22790,N_22666,N_22634);
and U22791 (N_22791,N_22637,N_22503);
xor U22792 (N_22792,N_22670,N_22552);
xnor U22793 (N_22793,N_22742,N_22569);
nor U22794 (N_22794,N_22680,N_22731);
xnor U22795 (N_22795,N_22518,N_22538);
or U22796 (N_22796,N_22619,N_22539);
nor U22797 (N_22797,N_22573,N_22625);
and U22798 (N_22798,N_22732,N_22525);
xor U22799 (N_22799,N_22559,N_22654);
and U22800 (N_22800,N_22709,N_22557);
xor U22801 (N_22801,N_22553,N_22683);
nand U22802 (N_22802,N_22574,N_22739);
and U22803 (N_22803,N_22602,N_22660);
nor U22804 (N_22804,N_22515,N_22700);
xor U22805 (N_22805,N_22592,N_22727);
nand U22806 (N_22806,N_22508,N_22618);
nor U22807 (N_22807,N_22558,N_22601);
and U22808 (N_22808,N_22644,N_22674);
or U22809 (N_22809,N_22545,N_22629);
xnor U22810 (N_22810,N_22509,N_22526);
nand U22811 (N_22811,N_22665,N_22563);
or U22812 (N_22812,N_22714,N_22500);
or U22813 (N_22813,N_22585,N_22600);
and U22814 (N_22814,N_22735,N_22640);
nor U22815 (N_22815,N_22745,N_22659);
or U22816 (N_22816,N_22613,N_22596);
or U22817 (N_22817,N_22667,N_22708);
or U22818 (N_22818,N_22528,N_22531);
and U22819 (N_22819,N_22661,N_22702);
and U22820 (N_22820,N_22693,N_22575);
xor U22821 (N_22821,N_22717,N_22627);
xnor U22822 (N_22822,N_22636,N_22658);
nand U22823 (N_22823,N_22682,N_22519);
or U22824 (N_22824,N_22588,N_22587);
nor U22825 (N_22825,N_22562,N_22567);
and U22826 (N_22826,N_22639,N_22738);
xnor U22827 (N_22827,N_22686,N_22542);
or U22828 (N_22828,N_22704,N_22691);
and U22829 (N_22829,N_22663,N_22706);
and U22830 (N_22830,N_22635,N_22652);
xor U22831 (N_22831,N_22550,N_22740);
or U22832 (N_22832,N_22520,N_22507);
and U22833 (N_22833,N_22543,N_22687);
nor U22834 (N_22834,N_22681,N_22662);
nor U22835 (N_22835,N_22671,N_22696);
nor U22836 (N_22836,N_22610,N_22556);
and U22837 (N_22837,N_22524,N_22641);
or U22838 (N_22838,N_22581,N_22719);
or U22839 (N_22839,N_22718,N_22579);
nand U22840 (N_22840,N_22737,N_22749);
and U22841 (N_22841,N_22578,N_22695);
xnor U22842 (N_22842,N_22730,N_22656);
or U22843 (N_22843,N_22747,N_22643);
nand U22844 (N_22844,N_22540,N_22560);
nor U22845 (N_22845,N_22705,N_22651);
xnor U22846 (N_22846,N_22688,N_22547);
xor U22847 (N_22847,N_22692,N_22746);
or U22848 (N_22848,N_22650,N_22510);
nor U22849 (N_22849,N_22669,N_22628);
nand U22850 (N_22850,N_22642,N_22657);
or U22851 (N_22851,N_22549,N_22554);
nand U22852 (N_22852,N_22595,N_22703);
and U22853 (N_22853,N_22675,N_22571);
and U22854 (N_22854,N_22612,N_22664);
nor U22855 (N_22855,N_22606,N_22715);
nor U22856 (N_22856,N_22583,N_22673);
or U22857 (N_22857,N_22701,N_22653);
nand U22858 (N_22858,N_22555,N_22699);
and U22859 (N_22859,N_22633,N_22586);
xnor U22860 (N_22860,N_22689,N_22698);
nand U22861 (N_22861,N_22537,N_22530);
or U22862 (N_22862,N_22568,N_22546);
and U22863 (N_22863,N_22646,N_22728);
and U22864 (N_22864,N_22532,N_22647);
and U22865 (N_22865,N_22511,N_22645);
xnor U22866 (N_22866,N_22713,N_22743);
and U22867 (N_22867,N_22734,N_22551);
nand U22868 (N_22868,N_22534,N_22533);
nand U22869 (N_22869,N_22611,N_22598);
xnor U22870 (N_22870,N_22615,N_22707);
nand U22871 (N_22871,N_22608,N_22620);
or U22872 (N_22872,N_22744,N_22577);
nand U22873 (N_22873,N_22561,N_22711);
or U22874 (N_22874,N_22566,N_22723);
nor U22875 (N_22875,N_22534,N_22692);
and U22876 (N_22876,N_22550,N_22672);
and U22877 (N_22877,N_22749,N_22550);
nand U22878 (N_22878,N_22662,N_22505);
or U22879 (N_22879,N_22509,N_22510);
nand U22880 (N_22880,N_22597,N_22513);
nor U22881 (N_22881,N_22541,N_22651);
nor U22882 (N_22882,N_22573,N_22661);
nand U22883 (N_22883,N_22568,N_22571);
or U22884 (N_22884,N_22720,N_22539);
nor U22885 (N_22885,N_22725,N_22573);
or U22886 (N_22886,N_22696,N_22639);
nand U22887 (N_22887,N_22687,N_22690);
or U22888 (N_22888,N_22731,N_22611);
nand U22889 (N_22889,N_22531,N_22508);
xnor U22890 (N_22890,N_22548,N_22722);
and U22891 (N_22891,N_22573,N_22637);
and U22892 (N_22892,N_22559,N_22506);
or U22893 (N_22893,N_22509,N_22585);
nor U22894 (N_22894,N_22668,N_22548);
or U22895 (N_22895,N_22617,N_22536);
or U22896 (N_22896,N_22728,N_22734);
nor U22897 (N_22897,N_22653,N_22540);
or U22898 (N_22898,N_22558,N_22602);
nor U22899 (N_22899,N_22682,N_22522);
nor U22900 (N_22900,N_22637,N_22574);
or U22901 (N_22901,N_22512,N_22504);
nor U22902 (N_22902,N_22663,N_22732);
nor U22903 (N_22903,N_22647,N_22581);
or U22904 (N_22904,N_22580,N_22529);
nand U22905 (N_22905,N_22742,N_22665);
nand U22906 (N_22906,N_22685,N_22556);
and U22907 (N_22907,N_22654,N_22684);
and U22908 (N_22908,N_22695,N_22568);
xnor U22909 (N_22909,N_22660,N_22617);
nand U22910 (N_22910,N_22649,N_22637);
xnor U22911 (N_22911,N_22664,N_22699);
and U22912 (N_22912,N_22685,N_22722);
and U22913 (N_22913,N_22743,N_22616);
nand U22914 (N_22914,N_22605,N_22591);
nor U22915 (N_22915,N_22509,N_22524);
nor U22916 (N_22916,N_22513,N_22629);
or U22917 (N_22917,N_22522,N_22667);
nand U22918 (N_22918,N_22613,N_22623);
and U22919 (N_22919,N_22544,N_22538);
and U22920 (N_22920,N_22589,N_22549);
xnor U22921 (N_22921,N_22733,N_22550);
nor U22922 (N_22922,N_22749,N_22733);
xnor U22923 (N_22923,N_22742,N_22559);
nor U22924 (N_22924,N_22501,N_22505);
and U22925 (N_22925,N_22540,N_22543);
nor U22926 (N_22926,N_22655,N_22724);
nand U22927 (N_22927,N_22619,N_22583);
and U22928 (N_22928,N_22575,N_22527);
or U22929 (N_22929,N_22500,N_22712);
nor U22930 (N_22930,N_22680,N_22617);
or U22931 (N_22931,N_22609,N_22563);
nor U22932 (N_22932,N_22506,N_22669);
nor U22933 (N_22933,N_22510,N_22575);
nand U22934 (N_22934,N_22662,N_22550);
and U22935 (N_22935,N_22611,N_22687);
nor U22936 (N_22936,N_22636,N_22677);
and U22937 (N_22937,N_22543,N_22707);
nor U22938 (N_22938,N_22600,N_22598);
nand U22939 (N_22939,N_22598,N_22502);
or U22940 (N_22940,N_22704,N_22690);
and U22941 (N_22941,N_22607,N_22566);
xor U22942 (N_22942,N_22679,N_22721);
xor U22943 (N_22943,N_22714,N_22703);
and U22944 (N_22944,N_22731,N_22580);
nor U22945 (N_22945,N_22733,N_22679);
or U22946 (N_22946,N_22673,N_22549);
and U22947 (N_22947,N_22589,N_22723);
or U22948 (N_22948,N_22672,N_22606);
nand U22949 (N_22949,N_22668,N_22725);
nand U22950 (N_22950,N_22505,N_22527);
nor U22951 (N_22951,N_22745,N_22625);
nor U22952 (N_22952,N_22584,N_22710);
or U22953 (N_22953,N_22640,N_22693);
or U22954 (N_22954,N_22687,N_22572);
nor U22955 (N_22955,N_22635,N_22584);
and U22956 (N_22956,N_22505,N_22548);
xnor U22957 (N_22957,N_22670,N_22705);
nand U22958 (N_22958,N_22558,N_22551);
or U22959 (N_22959,N_22529,N_22682);
nand U22960 (N_22960,N_22520,N_22653);
xnor U22961 (N_22961,N_22716,N_22592);
or U22962 (N_22962,N_22572,N_22704);
or U22963 (N_22963,N_22574,N_22724);
xnor U22964 (N_22964,N_22579,N_22717);
and U22965 (N_22965,N_22602,N_22507);
and U22966 (N_22966,N_22644,N_22552);
and U22967 (N_22967,N_22708,N_22642);
xor U22968 (N_22968,N_22581,N_22721);
or U22969 (N_22969,N_22701,N_22593);
nand U22970 (N_22970,N_22550,N_22579);
or U22971 (N_22971,N_22645,N_22602);
xor U22972 (N_22972,N_22704,N_22503);
xnor U22973 (N_22973,N_22557,N_22500);
xor U22974 (N_22974,N_22728,N_22660);
xor U22975 (N_22975,N_22508,N_22645);
nand U22976 (N_22976,N_22592,N_22745);
and U22977 (N_22977,N_22623,N_22637);
nor U22978 (N_22978,N_22705,N_22678);
xor U22979 (N_22979,N_22567,N_22677);
or U22980 (N_22980,N_22698,N_22546);
and U22981 (N_22981,N_22575,N_22667);
or U22982 (N_22982,N_22729,N_22635);
and U22983 (N_22983,N_22534,N_22512);
nand U22984 (N_22984,N_22503,N_22663);
nor U22985 (N_22985,N_22688,N_22555);
xnor U22986 (N_22986,N_22708,N_22663);
or U22987 (N_22987,N_22722,N_22588);
and U22988 (N_22988,N_22638,N_22622);
and U22989 (N_22989,N_22518,N_22531);
xor U22990 (N_22990,N_22531,N_22547);
and U22991 (N_22991,N_22743,N_22524);
and U22992 (N_22992,N_22640,N_22523);
and U22993 (N_22993,N_22745,N_22500);
xnor U22994 (N_22994,N_22630,N_22627);
or U22995 (N_22995,N_22543,N_22550);
and U22996 (N_22996,N_22521,N_22581);
nand U22997 (N_22997,N_22535,N_22514);
or U22998 (N_22998,N_22508,N_22583);
or U22999 (N_22999,N_22592,N_22629);
nor U23000 (N_23000,N_22865,N_22833);
nand U23001 (N_23001,N_22799,N_22887);
nand U23002 (N_23002,N_22800,N_22776);
or U23003 (N_23003,N_22936,N_22972);
or U23004 (N_23004,N_22761,N_22870);
nor U23005 (N_23005,N_22931,N_22991);
or U23006 (N_23006,N_22933,N_22874);
and U23007 (N_23007,N_22946,N_22967);
or U23008 (N_23008,N_22823,N_22829);
xnor U23009 (N_23009,N_22994,N_22818);
and U23010 (N_23010,N_22753,N_22948);
and U23011 (N_23011,N_22786,N_22839);
or U23012 (N_23012,N_22847,N_22883);
or U23013 (N_23013,N_22889,N_22898);
and U23014 (N_23014,N_22860,N_22770);
nand U23015 (N_23015,N_22825,N_22767);
or U23016 (N_23016,N_22861,N_22805);
nor U23017 (N_23017,N_22755,N_22966);
nor U23018 (N_23018,N_22928,N_22962);
and U23019 (N_23019,N_22932,N_22848);
and U23020 (N_23020,N_22896,N_22945);
nand U23021 (N_23021,N_22846,N_22797);
xnor U23022 (N_23022,N_22939,N_22777);
or U23023 (N_23023,N_22866,N_22989);
nand U23024 (N_23024,N_22971,N_22924);
or U23025 (N_23025,N_22869,N_22765);
and U23026 (N_23026,N_22804,N_22910);
nand U23027 (N_23027,N_22844,N_22852);
or U23028 (N_23028,N_22750,N_22773);
nor U23029 (N_23029,N_22787,N_22978);
nor U23030 (N_23030,N_22842,N_22892);
or U23031 (N_23031,N_22851,N_22821);
or U23032 (N_23032,N_22993,N_22768);
or U23033 (N_23033,N_22969,N_22778);
nor U23034 (N_23034,N_22999,N_22819);
or U23035 (N_23035,N_22888,N_22794);
nor U23036 (N_23036,N_22957,N_22783);
nor U23037 (N_23037,N_22752,N_22877);
xor U23038 (N_23038,N_22762,N_22836);
or U23039 (N_23039,N_22813,N_22830);
nor U23040 (N_23040,N_22902,N_22795);
xor U23041 (N_23041,N_22878,N_22769);
and U23042 (N_23042,N_22824,N_22873);
xnor U23043 (N_23043,N_22900,N_22827);
nor U23044 (N_23044,N_22816,N_22756);
or U23045 (N_23045,N_22970,N_22938);
or U23046 (N_23046,N_22868,N_22992);
xnor U23047 (N_23047,N_22879,N_22922);
or U23048 (N_23048,N_22942,N_22929);
or U23049 (N_23049,N_22781,N_22838);
and U23050 (N_23050,N_22858,N_22801);
and U23051 (N_23051,N_22990,N_22895);
and U23052 (N_23052,N_22826,N_22803);
or U23053 (N_23053,N_22906,N_22760);
nor U23054 (N_23054,N_22832,N_22996);
nor U23055 (N_23055,N_22940,N_22894);
nor U23056 (N_23056,N_22763,N_22817);
nand U23057 (N_23057,N_22974,N_22986);
or U23058 (N_23058,N_22925,N_22959);
nand U23059 (N_23059,N_22856,N_22893);
and U23060 (N_23060,N_22943,N_22960);
or U23061 (N_23061,N_22834,N_22855);
and U23062 (N_23062,N_22904,N_22984);
or U23063 (N_23063,N_22872,N_22798);
nor U23064 (N_23064,N_22909,N_22901);
nor U23065 (N_23065,N_22784,N_22771);
xnor U23066 (N_23066,N_22880,N_22806);
nand U23067 (N_23067,N_22837,N_22796);
or U23068 (N_23068,N_22905,N_22980);
or U23069 (N_23069,N_22863,N_22956);
xnor U23070 (N_23070,N_22754,N_22791);
xnor U23071 (N_23071,N_22897,N_22937);
or U23072 (N_23072,N_22881,N_22782);
nor U23073 (N_23073,N_22965,N_22914);
and U23074 (N_23074,N_22774,N_22891);
xor U23075 (N_23075,N_22822,N_22812);
or U23076 (N_23076,N_22814,N_22958);
or U23077 (N_23077,N_22841,N_22947);
nand U23078 (N_23078,N_22975,N_22859);
or U23079 (N_23079,N_22845,N_22964);
nand U23080 (N_23080,N_22950,N_22961);
nor U23081 (N_23081,N_22916,N_22785);
and U23082 (N_23082,N_22927,N_22998);
nor U23083 (N_23083,N_22985,N_22995);
xor U23084 (N_23084,N_22864,N_22923);
or U23085 (N_23085,N_22867,N_22875);
xor U23086 (N_23086,N_22831,N_22751);
nand U23087 (N_23087,N_22828,N_22807);
nand U23088 (N_23088,N_22772,N_22876);
and U23089 (N_23089,N_22759,N_22973);
xor U23090 (N_23090,N_22955,N_22857);
and U23091 (N_23091,N_22802,N_22780);
or U23092 (N_23092,N_22944,N_22913);
nand U23093 (N_23093,N_22885,N_22840);
and U23094 (N_23094,N_22911,N_22882);
or U23095 (N_23095,N_22890,N_22934);
and U23096 (N_23096,N_22951,N_22775);
nand U23097 (N_23097,N_22982,N_22757);
and U23098 (N_23098,N_22850,N_22997);
or U23099 (N_23099,N_22820,N_22835);
nand U23100 (N_23100,N_22808,N_22792);
nand U23101 (N_23101,N_22790,N_22983);
and U23102 (N_23102,N_22949,N_22917);
or U23103 (N_23103,N_22809,N_22968);
nand U23104 (N_23104,N_22912,N_22849);
and U23105 (N_23105,N_22854,N_22884);
xnor U23106 (N_23106,N_22953,N_22779);
or U23107 (N_23107,N_22811,N_22915);
and U23108 (N_23108,N_22899,N_22935);
xnor U23109 (N_23109,N_22976,N_22954);
and U23110 (N_23110,N_22871,N_22930);
xor U23111 (N_23111,N_22766,N_22764);
nor U23112 (N_23112,N_22988,N_22977);
nand U23113 (N_23113,N_22981,N_22903);
and U23114 (N_23114,N_22987,N_22919);
nor U23115 (N_23115,N_22788,N_22963);
nor U23116 (N_23116,N_22941,N_22758);
nand U23117 (N_23117,N_22862,N_22789);
or U23118 (N_23118,N_22810,N_22979);
or U23119 (N_23119,N_22815,N_22908);
xnor U23120 (N_23120,N_22793,N_22907);
nor U23121 (N_23121,N_22920,N_22926);
xor U23122 (N_23122,N_22843,N_22886);
nor U23123 (N_23123,N_22921,N_22853);
nor U23124 (N_23124,N_22918,N_22952);
xor U23125 (N_23125,N_22754,N_22887);
and U23126 (N_23126,N_22939,N_22923);
and U23127 (N_23127,N_22992,N_22759);
nor U23128 (N_23128,N_22808,N_22785);
xnor U23129 (N_23129,N_22893,N_22909);
or U23130 (N_23130,N_22866,N_22937);
and U23131 (N_23131,N_22944,N_22960);
nand U23132 (N_23132,N_22920,N_22940);
nand U23133 (N_23133,N_22790,N_22875);
nand U23134 (N_23134,N_22777,N_22840);
or U23135 (N_23135,N_22964,N_22887);
nor U23136 (N_23136,N_22780,N_22853);
xnor U23137 (N_23137,N_22990,N_22767);
or U23138 (N_23138,N_22833,N_22939);
or U23139 (N_23139,N_22947,N_22768);
and U23140 (N_23140,N_22802,N_22836);
xor U23141 (N_23141,N_22846,N_22757);
nand U23142 (N_23142,N_22989,N_22817);
or U23143 (N_23143,N_22871,N_22985);
nand U23144 (N_23144,N_22888,N_22973);
or U23145 (N_23145,N_22891,N_22921);
xnor U23146 (N_23146,N_22865,N_22916);
or U23147 (N_23147,N_22780,N_22879);
or U23148 (N_23148,N_22862,N_22778);
nor U23149 (N_23149,N_22871,N_22811);
nand U23150 (N_23150,N_22756,N_22825);
nand U23151 (N_23151,N_22936,N_22845);
xnor U23152 (N_23152,N_22982,N_22925);
xnor U23153 (N_23153,N_22819,N_22900);
and U23154 (N_23154,N_22834,N_22888);
or U23155 (N_23155,N_22962,N_22870);
and U23156 (N_23156,N_22910,N_22775);
or U23157 (N_23157,N_22773,N_22928);
nand U23158 (N_23158,N_22973,N_22848);
xor U23159 (N_23159,N_22927,N_22942);
and U23160 (N_23160,N_22865,N_22989);
and U23161 (N_23161,N_22881,N_22857);
or U23162 (N_23162,N_22922,N_22832);
xnor U23163 (N_23163,N_22924,N_22860);
xnor U23164 (N_23164,N_22990,N_22872);
nand U23165 (N_23165,N_22873,N_22763);
xor U23166 (N_23166,N_22957,N_22981);
xor U23167 (N_23167,N_22947,N_22925);
nand U23168 (N_23168,N_22999,N_22787);
nand U23169 (N_23169,N_22973,N_22783);
nor U23170 (N_23170,N_22807,N_22817);
nand U23171 (N_23171,N_22816,N_22762);
nor U23172 (N_23172,N_22865,N_22994);
nor U23173 (N_23173,N_22805,N_22753);
and U23174 (N_23174,N_22785,N_22948);
nand U23175 (N_23175,N_22827,N_22788);
nor U23176 (N_23176,N_22768,N_22793);
and U23177 (N_23177,N_22859,N_22767);
nand U23178 (N_23178,N_22915,N_22920);
nand U23179 (N_23179,N_22997,N_22991);
nand U23180 (N_23180,N_22772,N_22909);
nor U23181 (N_23181,N_22861,N_22937);
nor U23182 (N_23182,N_22896,N_22943);
or U23183 (N_23183,N_22770,N_22941);
xnor U23184 (N_23184,N_22771,N_22875);
or U23185 (N_23185,N_22813,N_22918);
nor U23186 (N_23186,N_22759,N_22901);
nor U23187 (N_23187,N_22806,N_22764);
or U23188 (N_23188,N_22915,N_22989);
and U23189 (N_23189,N_22771,N_22947);
xnor U23190 (N_23190,N_22885,N_22926);
or U23191 (N_23191,N_22979,N_22816);
xnor U23192 (N_23192,N_22820,N_22773);
and U23193 (N_23193,N_22781,N_22797);
nand U23194 (N_23194,N_22996,N_22844);
nor U23195 (N_23195,N_22922,N_22798);
nand U23196 (N_23196,N_22852,N_22907);
or U23197 (N_23197,N_22929,N_22827);
nand U23198 (N_23198,N_22957,N_22788);
and U23199 (N_23199,N_22873,N_22842);
xor U23200 (N_23200,N_22922,N_22781);
nand U23201 (N_23201,N_22776,N_22936);
xor U23202 (N_23202,N_22758,N_22887);
or U23203 (N_23203,N_22950,N_22979);
nand U23204 (N_23204,N_22871,N_22969);
or U23205 (N_23205,N_22835,N_22799);
xor U23206 (N_23206,N_22769,N_22948);
nor U23207 (N_23207,N_22978,N_22877);
xnor U23208 (N_23208,N_22829,N_22753);
and U23209 (N_23209,N_22980,N_22927);
and U23210 (N_23210,N_22810,N_22768);
nor U23211 (N_23211,N_22793,N_22893);
nand U23212 (N_23212,N_22783,N_22902);
or U23213 (N_23213,N_22996,N_22985);
or U23214 (N_23214,N_22909,N_22884);
and U23215 (N_23215,N_22925,N_22779);
nand U23216 (N_23216,N_22758,N_22892);
and U23217 (N_23217,N_22978,N_22915);
and U23218 (N_23218,N_22812,N_22762);
xor U23219 (N_23219,N_22907,N_22986);
nor U23220 (N_23220,N_22885,N_22812);
xor U23221 (N_23221,N_22887,N_22941);
xnor U23222 (N_23222,N_22808,N_22791);
nor U23223 (N_23223,N_22917,N_22845);
xnor U23224 (N_23224,N_22762,N_22909);
nor U23225 (N_23225,N_22993,N_22761);
nor U23226 (N_23226,N_22844,N_22870);
xor U23227 (N_23227,N_22973,N_22822);
nand U23228 (N_23228,N_22896,N_22968);
nor U23229 (N_23229,N_22950,N_22895);
xor U23230 (N_23230,N_22912,N_22798);
nand U23231 (N_23231,N_22958,N_22808);
nand U23232 (N_23232,N_22913,N_22979);
and U23233 (N_23233,N_22802,N_22774);
nand U23234 (N_23234,N_22806,N_22770);
nor U23235 (N_23235,N_22890,N_22881);
xor U23236 (N_23236,N_22815,N_22786);
nand U23237 (N_23237,N_22803,N_22939);
nor U23238 (N_23238,N_22888,N_22806);
nor U23239 (N_23239,N_22999,N_22941);
nor U23240 (N_23240,N_22871,N_22967);
xnor U23241 (N_23241,N_22947,N_22772);
xor U23242 (N_23242,N_22993,N_22885);
or U23243 (N_23243,N_22991,N_22962);
xnor U23244 (N_23244,N_22769,N_22788);
xor U23245 (N_23245,N_22908,N_22793);
and U23246 (N_23246,N_22934,N_22852);
and U23247 (N_23247,N_22846,N_22979);
nand U23248 (N_23248,N_22951,N_22970);
or U23249 (N_23249,N_22905,N_22997);
nor U23250 (N_23250,N_23101,N_23075);
or U23251 (N_23251,N_23192,N_23174);
xor U23252 (N_23252,N_23133,N_23023);
and U23253 (N_23253,N_23082,N_23145);
xnor U23254 (N_23254,N_23084,N_23178);
and U23255 (N_23255,N_23067,N_23048);
xnor U23256 (N_23256,N_23008,N_23236);
nand U23257 (N_23257,N_23244,N_23181);
or U23258 (N_23258,N_23005,N_23168);
xnor U23259 (N_23259,N_23165,N_23053);
nor U23260 (N_23260,N_23016,N_23017);
nand U23261 (N_23261,N_23211,N_23117);
and U23262 (N_23262,N_23076,N_23202);
nand U23263 (N_23263,N_23201,N_23109);
nand U23264 (N_23264,N_23136,N_23043);
or U23265 (N_23265,N_23175,N_23121);
xnor U23266 (N_23266,N_23152,N_23128);
xnor U23267 (N_23267,N_23034,N_23057);
or U23268 (N_23268,N_23242,N_23006);
xnor U23269 (N_23269,N_23146,N_23170);
nor U23270 (N_23270,N_23234,N_23130);
nand U23271 (N_23271,N_23229,N_23065);
nand U23272 (N_23272,N_23206,N_23245);
and U23273 (N_23273,N_23177,N_23194);
nand U23274 (N_23274,N_23155,N_23191);
nor U23275 (N_23275,N_23169,N_23135);
and U23276 (N_23276,N_23064,N_23077);
or U23277 (N_23277,N_23239,N_23100);
nand U23278 (N_23278,N_23197,N_23086);
xor U23279 (N_23279,N_23156,N_23096);
nand U23280 (N_23280,N_23089,N_23013);
nand U23281 (N_23281,N_23238,N_23209);
or U23282 (N_23282,N_23226,N_23220);
and U23283 (N_23283,N_23161,N_23088);
and U23284 (N_23284,N_23148,N_23102);
or U23285 (N_23285,N_23228,N_23003);
nand U23286 (N_23286,N_23176,N_23112);
and U23287 (N_23287,N_23036,N_23164);
nor U23288 (N_23288,N_23007,N_23137);
or U23289 (N_23289,N_23231,N_23074);
xor U23290 (N_23290,N_23200,N_23113);
and U23291 (N_23291,N_23040,N_23061);
or U23292 (N_23292,N_23166,N_23223);
xor U23293 (N_23293,N_23087,N_23103);
xnor U23294 (N_23294,N_23157,N_23217);
nor U23295 (N_23295,N_23190,N_23021);
nor U23296 (N_23296,N_23237,N_23111);
nor U23297 (N_23297,N_23131,N_23218);
or U23298 (N_23298,N_23095,N_23104);
xor U23299 (N_23299,N_23062,N_23119);
or U23300 (N_23300,N_23060,N_23026);
or U23301 (N_23301,N_23204,N_23120);
xnor U23302 (N_23302,N_23031,N_23068);
nor U23303 (N_23303,N_23207,N_23247);
xor U23304 (N_23304,N_23212,N_23085);
and U23305 (N_23305,N_23230,N_23147);
and U23306 (N_23306,N_23173,N_23032);
and U23307 (N_23307,N_23159,N_23000);
and U23308 (N_23308,N_23183,N_23070);
or U23309 (N_23309,N_23078,N_23210);
xor U23310 (N_23310,N_23019,N_23222);
xor U23311 (N_23311,N_23184,N_23105);
and U23312 (N_23312,N_23205,N_23213);
and U23313 (N_23313,N_23083,N_23046);
and U23314 (N_23314,N_23134,N_23091);
nor U23315 (N_23315,N_23153,N_23129);
or U23316 (N_23316,N_23160,N_23058);
and U23317 (N_23317,N_23122,N_23246);
or U23318 (N_23318,N_23193,N_23187);
and U23319 (N_23319,N_23047,N_23241);
or U23320 (N_23320,N_23052,N_23004);
nand U23321 (N_23321,N_23009,N_23158);
nor U23322 (N_23322,N_23185,N_23198);
nor U23323 (N_23323,N_23069,N_23195);
and U23324 (N_23324,N_23029,N_23154);
xnor U23325 (N_23325,N_23215,N_23056);
or U23326 (N_23326,N_23039,N_23033);
nor U23327 (N_23327,N_23010,N_23038);
xor U23328 (N_23328,N_23214,N_23240);
xor U23329 (N_23329,N_23115,N_23015);
xnor U23330 (N_23330,N_23225,N_23232);
nor U23331 (N_23331,N_23167,N_23024);
or U23332 (N_23332,N_23118,N_23149);
xnor U23333 (N_23333,N_23059,N_23142);
and U23334 (N_23334,N_23203,N_23186);
and U23335 (N_23335,N_23182,N_23051);
nand U23336 (N_23336,N_23018,N_23138);
nor U23337 (N_23337,N_23106,N_23248);
and U23338 (N_23338,N_23045,N_23126);
and U23339 (N_23339,N_23072,N_23014);
xnor U23340 (N_23340,N_23063,N_23093);
nor U23341 (N_23341,N_23243,N_23127);
xor U23342 (N_23342,N_23125,N_23073);
nand U23343 (N_23343,N_23216,N_23180);
xnor U23344 (N_23344,N_23199,N_23108);
nand U23345 (N_23345,N_23141,N_23172);
nor U23346 (N_23346,N_23219,N_23163);
and U23347 (N_23347,N_23114,N_23233);
nor U23348 (N_23348,N_23099,N_23150);
or U23349 (N_23349,N_23079,N_23124);
and U23350 (N_23350,N_23035,N_23151);
nor U23351 (N_23351,N_23097,N_23042);
or U23352 (N_23352,N_23143,N_23110);
nand U23353 (N_23353,N_23139,N_23144);
and U23354 (N_23354,N_23249,N_23049);
nand U23355 (N_23355,N_23041,N_23066);
and U23356 (N_23356,N_23054,N_23094);
nor U23357 (N_23357,N_23171,N_23080);
nand U23358 (N_23358,N_23055,N_23235);
or U23359 (N_23359,N_23027,N_23179);
nand U23360 (N_23360,N_23107,N_23123);
nor U23361 (N_23361,N_23071,N_23011);
or U23362 (N_23362,N_23116,N_23098);
xor U23363 (N_23363,N_23092,N_23001);
xnor U23364 (N_23364,N_23221,N_23012);
and U23365 (N_23365,N_23028,N_23224);
or U23366 (N_23366,N_23090,N_23037);
or U23367 (N_23367,N_23081,N_23022);
xor U23368 (N_23368,N_23227,N_23162);
xor U23369 (N_23369,N_23140,N_23188);
or U23370 (N_23370,N_23025,N_23002);
nand U23371 (N_23371,N_23196,N_23208);
xor U23372 (N_23372,N_23030,N_23050);
nand U23373 (N_23373,N_23044,N_23020);
nand U23374 (N_23374,N_23132,N_23189);
or U23375 (N_23375,N_23247,N_23049);
nor U23376 (N_23376,N_23164,N_23073);
xor U23377 (N_23377,N_23216,N_23217);
or U23378 (N_23378,N_23208,N_23226);
nor U23379 (N_23379,N_23059,N_23099);
nor U23380 (N_23380,N_23232,N_23079);
and U23381 (N_23381,N_23092,N_23027);
or U23382 (N_23382,N_23054,N_23068);
nor U23383 (N_23383,N_23082,N_23029);
and U23384 (N_23384,N_23125,N_23058);
nand U23385 (N_23385,N_23249,N_23088);
and U23386 (N_23386,N_23028,N_23208);
or U23387 (N_23387,N_23117,N_23049);
xor U23388 (N_23388,N_23228,N_23164);
xor U23389 (N_23389,N_23041,N_23046);
nand U23390 (N_23390,N_23118,N_23013);
nor U23391 (N_23391,N_23188,N_23205);
nand U23392 (N_23392,N_23191,N_23144);
or U23393 (N_23393,N_23135,N_23207);
xnor U23394 (N_23394,N_23043,N_23012);
and U23395 (N_23395,N_23036,N_23236);
and U23396 (N_23396,N_23158,N_23143);
nand U23397 (N_23397,N_23066,N_23032);
and U23398 (N_23398,N_23120,N_23241);
and U23399 (N_23399,N_23098,N_23192);
or U23400 (N_23400,N_23091,N_23236);
nand U23401 (N_23401,N_23207,N_23116);
nand U23402 (N_23402,N_23120,N_23178);
or U23403 (N_23403,N_23208,N_23030);
or U23404 (N_23404,N_23129,N_23235);
and U23405 (N_23405,N_23083,N_23015);
nand U23406 (N_23406,N_23084,N_23093);
or U23407 (N_23407,N_23058,N_23000);
xor U23408 (N_23408,N_23126,N_23173);
xor U23409 (N_23409,N_23119,N_23143);
nor U23410 (N_23410,N_23069,N_23060);
nor U23411 (N_23411,N_23214,N_23101);
and U23412 (N_23412,N_23155,N_23146);
nor U23413 (N_23413,N_23071,N_23109);
nor U23414 (N_23414,N_23104,N_23018);
and U23415 (N_23415,N_23213,N_23226);
xor U23416 (N_23416,N_23002,N_23107);
and U23417 (N_23417,N_23034,N_23211);
nand U23418 (N_23418,N_23166,N_23182);
or U23419 (N_23419,N_23006,N_23129);
and U23420 (N_23420,N_23205,N_23144);
nand U23421 (N_23421,N_23206,N_23127);
nand U23422 (N_23422,N_23160,N_23095);
xnor U23423 (N_23423,N_23214,N_23187);
nand U23424 (N_23424,N_23139,N_23120);
or U23425 (N_23425,N_23134,N_23059);
or U23426 (N_23426,N_23146,N_23207);
nand U23427 (N_23427,N_23186,N_23228);
nor U23428 (N_23428,N_23065,N_23116);
nor U23429 (N_23429,N_23197,N_23196);
or U23430 (N_23430,N_23182,N_23004);
xnor U23431 (N_23431,N_23076,N_23142);
or U23432 (N_23432,N_23061,N_23098);
xnor U23433 (N_23433,N_23139,N_23110);
and U23434 (N_23434,N_23002,N_23137);
nor U23435 (N_23435,N_23020,N_23167);
xor U23436 (N_23436,N_23148,N_23091);
nor U23437 (N_23437,N_23175,N_23189);
nor U23438 (N_23438,N_23080,N_23224);
nand U23439 (N_23439,N_23047,N_23167);
nand U23440 (N_23440,N_23152,N_23201);
nor U23441 (N_23441,N_23122,N_23066);
or U23442 (N_23442,N_23220,N_23210);
nor U23443 (N_23443,N_23018,N_23123);
xor U23444 (N_23444,N_23153,N_23126);
and U23445 (N_23445,N_23199,N_23243);
nand U23446 (N_23446,N_23135,N_23096);
and U23447 (N_23447,N_23031,N_23070);
xor U23448 (N_23448,N_23096,N_23125);
xnor U23449 (N_23449,N_23077,N_23031);
and U23450 (N_23450,N_23156,N_23059);
xor U23451 (N_23451,N_23164,N_23015);
nand U23452 (N_23452,N_23031,N_23148);
and U23453 (N_23453,N_23122,N_23112);
and U23454 (N_23454,N_23044,N_23139);
or U23455 (N_23455,N_23187,N_23170);
and U23456 (N_23456,N_23226,N_23246);
or U23457 (N_23457,N_23196,N_23012);
nand U23458 (N_23458,N_23206,N_23090);
xnor U23459 (N_23459,N_23042,N_23178);
nand U23460 (N_23460,N_23132,N_23015);
xnor U23461 (N_23461,N_23108,N_23035);
xnor U23462 (N_23462,N_23184,N_23155);
and U23463 (N_23463,N_23128,N_23155);
or U23464 (N_23464,N_23056,N_23207);
or U23465 (N_23465,N_23146,N_23005);
and U23466 (N_23466,N_23108,N_23197);
or U23467 (N_23467,N_23233,N_23050);
nand U23468 (N_23468,N_23212,N_23138);
or U23469 (N_23469,N_23051,N_23197);
xor U23470 (N_23470,N_23132,N_23160);
nand U23471 (N_23471,N_23004,N_23070);
or U23472 (N_23472,N_23057,N_23231);
nor U23473 (N_23473,N_23214,N_23242);
nor U23474 (N_23474,N_23130,N_23203);
nor U23475 (N_23475,N_23122,N_23009);
nand U23476 (N_23476,N_23225,N_23077);
xnor U23477 (N_23477,N_23157,N_23079);
nor U23478 (N_23478,N_23232,N_23054);
or U23479 (N_23479,N_23043,N_23218);
xor U23480 (N_23480,N_23113,N_23127);
or U23481 (N_23481,N_23193,N_23184);
or U23482 (N_23482,N_23013,N_23235);
and U23483 (N_23483,N_23076,N_23010);
or U23484 (N_23484,N_23129,N_23240);
nor U23485 (N_23485,N_23020,N_23134);
nor U23486 (N_23486,N_23123,N_23030);
and U23487 (N_23487,N_23018,N_23022);
xor U23488 (N_23488,N_23203,N_23094);
nor U23489 (N_23489,N_23179,N_23162);
xor U23490 (N_23490,N_23220,N_23194);
nand U23491 (N_23491,N_23170,N_23218);
or U23492 (N_23492,N_23069,N_23198);
xnor U23493 (N_23493,N_23228,N_23107);
or U23494 (N_23494,N_23126,N_23092);
or U23495 (N_23495,N_23072,N_23109);
nor U23496 (N_23496,N_23020,N_23068);
nand U23497 (N_23497,N_23212,N_23147);
nor U23498 (N_23498,N_23114,N_23177);
nor U23499 (N_23499,N_23165,N_23204);
or U23500 (N_23500,N_23318,N_23466);
or U23501 (N_23501,N_23262,N_23345);
nand U23502 (N_23502,N_23255,N_23475);
xor U23503 (N_23503,N_23461,N_23264);
or U23504 (N_23504,N_23292,N_23270);
and U23505 (N_23505,N_23320,N_23409);
and U23506 (N_23506,N_23263,N_23400);
nand U23507 (N_23507,N_23381,N_23382);
xnor U23508 (N_23508,N_23251,N_23361);
xor U23509 (N_23509,N_23302,N_23453);
xor U23510 (N_23510,N_23498,N_23285);
and U23511 (N_23511,N_23380,N_23434);
nor U23512 (N_23512,N_23317,N_23405);
nand U23513 (N_23513,N_23481,N_23343);
xnor U23514 (N_23514,N_23399,N_23493);
xnor U23515 (N_23515,N_23342,N_23269);
or U23516 (N_23516,N_23406,N_23344);
xor U23517 (N_23517,N_23412,N_23433);
and U23518 (N_23518,N_23467,N_23408);
nor U23519 (N_23519,N_23303,N_23259);
or U23520 (N_23520,N_23415,N_23458);
nand U23521 (N_23521,N_23266,N_23418);
xor U23522 (N_23522,N_23425,N_23328);
and U23523 (N_23523,N_23252,N_23474);
or U23524 (N_23524,N_23265,N_23478);
xnor U23525 (N_23525,N_23393,N_23451);
nor U23526 (N_23526,N_23330,N_23295);
xor U23527 (N_23527,N_23485,N_23395);
nor U23528 (N_23528,N_23438,N_23437);
nor U23529 (N_23529,N_23424,N_23482);
nor U23530 (N_23530,N_23370,N_23309);
nand U23531 (N_23531,N_23427,N_23294);
nor U23532 (N_23532,N_23304,N_23281);
nor U23533 (N_23533,N_23457,N_23348);
and U23534 (N_23534,N_23279,N_23416);
nand U23535 (N_23535,N_23488,N_23456);
and U23536 (N_23536,N_23316,N_23460);
or U23537 (N_23537,N_23315,N_23258);
nor U23538 (N_23538,N_23256,N_23273);
nand U23539 (N_23539,N_23301,N_23374);
or U23540 (N_23540,N_23357,N_23383);
xor U23541 (N_23541,N_23404,N_23337);
nor U23542 (N_23542,N_23336,N_23463);
nor U23543 (N_23543,N_23402,N_23452);
nand U23544 (N_23544,N_23355,N_23277);
and U23545 (N_23545,N_23496,N_23486);
xor U23546 (N_23546,N_23378,N_23322);
nand U23547 (N_23547,N_23310,N_23396);
xor U23548 (N_23548,N_23254,N_23299);
and U23549 (N_23549,N_23275,N_23298);
or U23550 (N_23550,N_23468,N_23426);
nand U23551 (N_23551,N_23489,N_23454);
xnor U23552 (N_23552,N_23379,N_23449);
xnor U23553 (N_23553,N_23366,N_23494);
and U23554 (N_23554,N_23436,N_23432);
or U23555 (N_23555,N_23308,N_23313);
or U23556 (N_23556,N_23441,N_23431);
and U23557 (N_23557,N_23423,N_23284);
and U23558 (N_23558,N_23377,N_23483);
and U23559 (N_23559,N_23332,N_23398);
nor U23560 (N_23560,N_23392,N_23338);
or U23561 (N_23561,N_23329,N_23492);
nor U23562 (N_23562,N_23397,N_23479);
or U23563 (N_23563,N_23368,N_23359);
or U23564 (N_23564,N_23472,N_23282);
and U23565 (N_23565,N_23495,N_23356);
xor U23566 (N_23566,N_23365,N_23323);
nor U23567 (N_23567,N_23363,N_23499);
and U23568 (N_23568,N_23417,N_23307);
nor U23569 (N_23569,N_23290,N_23419);
xnor U23570 (N_23570,N_23455,N_23459);
nor U23571 (N_23571,N_23387,N_23391);
nand U23572 (N_23572,N_23354,N_23369);
and U23573 (N_23573,N_23278,N_23465);
xnor U23574 (N_23574,N_23422,N_23326);
or U23575 (N_23575,N_23325,N_23420);
nand U23576 (N_23576,N_23407,N_23351);
or U23577 (N_23577,N_23293,N_23352);
nand U23578 (N_23578,N_23257,N_23261);
or U23579 (N_23579,N_23267,N_23471);
xor U23580 (N_23580,N_23291,N_23401);
or U23581 (N_23581,N_23447,N_23477);
xnor U23582 (N_23582,N_23339,N_23312);
nand U23583 (N_23583,N_23413,N_23464);
and U23584 (N_23584,N_23296,N_23271);
and U23585 (N_23585,N_23372,N_23444);
nand U23586 (N_23586,N_23314,N_23272);
nor U23587 (N_23587,N_23414,N_23428);
and U23588 (N_23588,N_23394,N_23390);
nand U23589 (N_23589,N_23327,N_23403);
nand U23590 (N_23590,N_23324,N_23435);
xnor U23591 (N_23591,N_23491,N_23353);
or U23592 (N_23592,N_23469,N_23311);
and U23593 (N_23593,N_23333,N_23376);
xnor U23594 (N_23594,N_23490,N_23331);
nand U23595 (N_23595,N_23288,N_23410);
and U23596 (N_23596,N_23286,N_23283);
nand U23597 (N_23597,N_23470,N_23364);
nor U23598 (N_23598,N_23446,N_23442);
xnor U23599 (N_23599,N_23276,N_23289);
xnor U23600 (N_23600,N_23385,N_23305);
xor U23601 (N_23601,N_23487,N_23450);
xor U23602 (N_23602,N_23268,N_23300);
nor U23603 (N_23603,N_23462,N_23362);
nand U23604 (N_23604,N_23253,N_23389);
nand U23605 (N_23605,N_23384,N_23448);
nor U23606 (N_23606,N_23360,N_23430);
xnor U23607 (N_23607,N_23476,N_23334);
nand U23608 (N_23608,N_23497,N_23473);
or U23609 (N_23609,N_23274,N_23250);
nor U23610 (N_23610,N_23480,N_23297);
or U23611 (N_23611,N_23340,N_23287);
nand U23612 (N_23612,N_23440,N_23349);
or U23613 (N_23613,N_23371,N_23341);
xnor U23614 (N_23614,N_23421,N_23319);
or U23615 (N_23615,N_23346,N_23439);
nand U23616 (N_23616,N_23367,N_23373);
and U23617 (N_23617,N_23350,N_23347);
nand U23618 (N_23618,N_23386,N_23260);
xnor U23619 (N_23619,N_23375,N_23443);
xnor U23620 (N_23620,N_23445,N_23429);
and U23621 (N_23621,N_23411,N_23358);
nand U23622 (N_23622,N_23306,N_23280);
nand U23623 (N_23623,N_23335,N_23484);
or U23624 (N_23624,N_23321,N_23388);
nand U23625 (N_23625,N_23408,N_23317);
or U23626 (N_23626,N_23289,N_23361);
and U23627 (N_23627,N_23420,N_23372);
nand U23628 (N_23628,N_23369,N_23323);
nor U23629 (N_23629,N_23408,N_23406);
nor U23630 (N_23630,N_23251,N_23454);
xor U23631 (N_23631,N_23380,N_23414);
nor U23632 (N_23632,N_23477,N_23387);
xor U23633 (N_23633,N_23286,N_23252);
nor U23634 (N_23634,N_23485,N_23464);
or U23635 (N_23635,N_23340,N_23364);
and U23636 (N_23636,N_23405,N_23497);
nor U23637 (N_23637,N_23490,N_23261);
nor U23638 (N_23638,N_23424,N_23467);
xor U23639 (N_23639,N_23259,N_23352);
and U23640 (N_23640,N_23462,N_23347);
nand U23641 (N_23641,N_23458,N_23495);
or U23642 (N_23642,N_23374,N_23256);
and U23643 (N_23643,N_23314,N_23495);
or U23644 (N_23644,N_23479,N_23354);
or U23645 (N_23645,N_23255,N_23300);
and U23646 (N_23646,N_23460,N_23452);
nand U23647 (N_23647,N_23344,N_23302);
xnor U23648 (N_23648,N_23495,N_23258);
nor U23649 (N_23649,N_23267,N_23354);
or U23650 (N_23650,N_23478,N_23481);
nand U23651 (N_23651,N_23445,N_23449);
or U23652 (N_23652,N_23410,N_23470);
or U23653 (N_23653,N_23441,N_23418);
nand U23654 (N_23654,N_23255,N_23447);
nor U23655 (N_23655,N_23373,N_23433);
or U23656 (N_23656,N_23408,N_23490);
nand U23657 (N_23657,N_23375,N_23418);
or U23658 (N_23658,N_23471,N_23338);
or U23659 (N_23659,N_23479,N_23266);
or U23660 (N_23660,N_23395,N_23397);
xnor U23661 (N_23661,N_23418,N_23434);
or U23662 (N_23662,N_23471,N_23475);
xnor U23663 (N_23663,N_23469,N_23268);
and U23664 (N_23664,N_23272,N_23251);
nand U23665 (N_23665,N_23405,N_23332);
nor U23666 (N_23666,N_23300,N_23422);
nor U23667 (N_23667,N_23438,N_23279);
nand U23668 (N_23668,N_23456,N_23264);
xnor U23669 (N_23669,N_23445,N_23328);
or U23670 (N_23670,N_23334,N_23289);
or U23671 (N_23671,N_23492,N_23282);
nor U23672 (N_23672,N_23387,N_23328);
nor U23673 (N_23673,N_23326,N_23300);
and U23674 (N_23674,N_23421,N_23402);
nor U23675 (N_23675,N_23353,N_23478);
xnor U23676 (N_23676,N_23311,N_23420);
nor U23677 (N_23677,N_23352,N_23429);
or U23678 (N_23678,N_23423,N_23458);
nor U23679 (N_23679,N_23355,N_23377);
xnor U23680 (N_23680,N_23441,N_23319);
or U23681 (N_23681,N_23278,N_23393);
and U23682 (N_23682,N_23376,N_23352);
and U23683 (N_23683,N_23382,N_23279);
or U23684 (N_23684,N_23373,N_23435);
nand U23685 (N_23685,N_23275,N_23440);
or U23686 (N_23686,N_23271,N_23334);
or U23687 (N_23687,N_23262,N_23267);
xor U23688 (N_23688,N_23323,N_23401);
and U23689 (N_23689,N_23462,N_23483);
xnor U23690 (N_23690,N_23300,N_23256);
and U23691 (N_23691,N_23371,N_23264);
nand U23692 (N_23692,N_23270,N_23269);
nand U23693 (N_23693,N_23257,N_23476);
and U23694 (N_23694,N_23375,N_23278);
or U23695 (N_23695,N_23497,N_23495);
nor U23696 (N_23696,N_23265,N_23426);
nor U23697 (N_23697,N_23292,N_23353);
and U23698 (N_23698,N_23439,N_23326);
or U23699 (N_23699,N_23356,N_23264);
xnor U23700 (N_23700,N_23271,N_23405);
nand U23701 (N_23701,N_23457,N_23286);
xnor U23702 (N_23702,N_23479,N_23311);
xnor U23703 (N_23703,N_23429,N_23488);
nand U23704 (N_23704,N_23310,N_23350);
nor U23705 (N_23705,N_23466,N_23474);
xor U23706 (N_23706,N_23498,N_23334);
nor U23707 (N_23707,N_23418,N_23278);
nor U23708 (N_23708,N_23462,N_23427);
and U23709 (N_23709,N_23430,N_23395);
nand U23710 (N_23710,N_23452,N_23266);
nand U23711 (N_23711,N_23280,N_23286);
xnor U23712 (N_23712,N_23407,N_23291);
or U23713 (N_23713,N_23311,N_23419);
or U23714 (N_23714,N_23467,N_23402);
and U23715 (N_23715,N_23313,N_23357);
or U23716 (N_23716,N_23457,N_23365);
nor U23717 (N_23717,N_23335,N_23336);
and U23718 (N_23718,N_23343,N_23332);
and U23719 (N_23719,N_23279,N_23474);
and U23720 (N_23720,N_23298,N_23384);
xor U23721 (N_23721,N_23305,N_23459);
nand U23722 (N_23722,N_23487,N_23363);
and U23723 (N_23723,N_23487,N_23486);
or U23724 (N_23724,N_23498,N_23469);
nor U23725 (N_23725,N_23276,N_23277);
nor U23726 (N_23726,N_23309,N_23444);
nor U23727 (N_23727,N_23326,N_23260);
and U23728 (N_23728,N_23355,N_23382);
xor U23729 (N_23729,N_23286,N_23473);
nand U23730 (N_23730,N_23318,N_23496);
nand U23731 (N_23731,N_23272,N_23302);
and U23732 (N_23732,N_23282,N_23493);
xnor U23733 (N_23733,N_23293,N_23309);
or U23734 (N_23734,N_23356,N_23270);
xor U23735 (N_23735,N_23314,N_23318);
nand U23736 (N_23736,N_23271,N_23483);
or U23737 (N_23737,N_23370,N_23266);
or U23738 (N_23738,N_23346,N_23365);
nor U23739 (N_23739,N_23339,N_23306);
and U23740 (N_23740,N_23478,N_23376);
nand U23741 (N_23741,N_23436,N_23332);
or U23742 (N_23742,N_23431,N_23255);
xor U23743 (N_23743,N_23319,N_23384);
and U23744 (N_23744,N_23453,N_23422);
xnor U23745 (N_23745,N_23418,N_23280);
and U23746 (N_23746,N_23406,N_23319);
xor U23747 (N_23747,N_23463,N_23408);
xor U23748 (N_23748,N_23485,N_23291);
nor U23749 (N_23749,N_23282,N_23270);
or U23750 (N_23750,N_23502,N_23621);
xnor U23751 (N_23751,N_23639,N_23721);
and U23752 (N_23752,N_23746,N_23553);
and U23753 (N_23753,N_23535,N_23573);
or U23754 (N_23754,N_23522,N_23557);
nand U23755 (N_23755,N_23723,N_23541);
nor U23756 (N_23756,N_23585,N_23577);
or U23757 (N_23757,N_23580,N_23685);
nor U23758 (N_23758,N_23520,N_23665);
nor U23759 (N_23759,N_23538,N_23513);
nor U23760 (N_23760,N_23567,N_23619);
nor U23761 (N_23761,N_23725,N_23674);
xnor U23762 (N_23762,N_23652,N_23667);
or U23763 (N_23763,N_23632,N_23681);
xnor U23764 (N_23764,N_23518,N_23542);
or U23765 (N_23765,N_23612,N_23544);
nand U23766 (N_23766,N_23673,N_23747);
nor U23767 (N_23767,N_23514,N_23593);
xor U23768 (N_23768,N_23555,N_23688);
or U23769 (N_23769,N_23635,N_23734);
nand U23770 (N_23770,N_23724,N_23562);
nor U23771 (N_23771,N_23702,N_23661);
or U23772 (N_23772,N_23568,N_23708);
nor U23773 (N_23773,N_23655,N_23602);
xor U23774 (N_23774,N_23715,N_23503);
nand U23775 (N_23775,N_23537,N_23556);
and U23776 (N_23776,N_23682,N_23578);
or U23777 (N_23777,N_23710,N_23588);
nor U23778 (N_23778,N_23605,N_23699);
nand U23779 (N_23779,N_23560,N_23575);
nor U23780 (N_23780,N_23533,N_23552);
or U23781 (N_23781,N_23579,N_23517);
or U23782 (N_23782,N_23549,N_23510);
and U23783 (N_23783,N_23569,N_23660);
xnor U23784 (N_23784,N_23664,N_23519);
xor U23785 (N_23785,N_23689,N_23611);
or U23786 (N_23786,N_23730,N_23618);
nor U23787 (N_23787,N_23629,N_23550);
and U23788 (N_23788,N_23693,N_23726);
nand U23789 (N_23789,N_23515,N_23532);
xor U23790 (N_23790,N_23500,N_23528);
or U23791 (N_23791,N_23564,N_23608);
nand U23792 (N_23792,N_23590,N_23703);
nor U23793 (N_23793,N_23624,N_23679);
and U23794 (N_23794,N_23543,N_23672);
nor U23795 (N_23795,N_23701,N_23646);
xnor U23796 (N_23796,N_23582,N_23627);
and U23797 (N_23797,N_23743,N_23698);
xor U23798 (N_23798,N_23524,N_23576);
or U23799 (N_23799,N_23650,N_23606);
and U23800 (N_23800,N_23668,N_23600);
nor U23801 (N_23801,N_23675,N_23731);
xnor U23802 (N_23802,N_23539,N_23735);
or U23803 (N_23803,N_23589,N_23643);
nor U23804 (N_23804,N_23738,N_23603);
nor U23805 (N_23805,N_23531,N_23604);
or U23806 (N_23806,N_23653,N_23545);
nor U23807 (N_23807,N_23598,N_23656);
and U23808 (N_23808,N_23565,N_23687);
nor U23809 (N_23809,N_23613,N_23663);
nand U23810 (N_23810,N_23647,N_23622);
xnor U23811 (N_23811,N_23530,N_23529);
nand U23812 (N_23812,N_23718,N_23620);
nand U23813 (N_23813,N_23527,N_23601);
nand U23814 (N_23814,N_23630,N_23677);
xor U23815 (N_23815,N_23511,N_23691);
or U23816 (N_23816,N_23709,N_23516);
or U23817 (N_23817,N_23645,N_23566);
or U23818 (N_23818,N_23628,N_23716);
nand U23819 (N_23819,N_23626,N_23637);
nand U23820 (N_23820,N_23540,N_23594);
nand U23821 (N_23821,N_23700,N_23648);
nand U23822 (N_23822,N_23587,N_23658);
or U23823 (N_23823,N_23633,N_23631);
and U23824 (N_23824,N_23615,N_23670);
xor U23825 (N_23825,N_23680,N_23742);
and U23826 (N_23826,N_23739,N_23683);
or U23827 (N_23827,N_23662,N_23625);
or U23828 (N_23828,N_23748,N_23642);
and U23829 (N_23829,N_23737,N_23728);
nand U23830 (N_23830,N_23581,N_23671);
or U23831 (N_23831,N_23546,N_23690);
or U23832 (N_23832,N_23644,N_23504);
xor U23833 (N_23833,N_23634,N_23706);
and U23834 (N_23834,N_23714,N_23696);
xnor U23835 (N_23835,N_23583,N_23526);
nor U23836 (N_23836,N_23720,N_23676);
or U23837 (N_23837,N_23554,N_23505);
nor U23838 (N_23838,N_23512,N_23744);
nand U23839 (N_23839,N_23669,N_23713);
nand U23840 (N_23840,N_23607,N_23741);
nand U23841 (N_23841,N_23745,N_23610);
nand U23842 (N_23842,N_23599,N_23616);
and U23843 (N_23843,N_23561,N_23609);
or U23844 (N_23844,N_23595,N_23570);
nand U23845 (N_23845,N_23558,N_23727);
or U23846 (N_23846,N_23684,N_23749);
nand U23847 (N_23847,N_23641,N_23551);
xor U23848 (N_23848,N_23509,N_23719);
nor U23849 (N_23849,N_23572,N_23640);
nor U23850 (N_23850,N_23678,N_23584);
nand U23851 (N_23851,N_23695,N_23636);
or U23852 (N_23852,N_23597,N_23506);
nand U23853 (N_23853,N_23548,N_23722);
or U23854 (N_23854,N_23717,N_23586);
nand U23855 (N_23855,N_23571,N_23536);
nor U23856 (N_23856,N_23574,N_23501);
nand U23857 (N_23857,N_23712,N_23657);
nand U23858 (N_23858,N_23638,N_23596);
and U23859 (N_23859,N_23736,N_23623);
nand U23860 (N_23860,N_23704,N_23694);
nor U23861 (N_23861,N_23521,N_23666);
nand U23862 (N_23862,N_23707,N_23559);
xnor U23863 (N_23863,N_23733,N_23654);
or U23864 (N_23864,N_23697,N_23523);
and U23865 (N_23865,N_23686,N_23547);
and U23866 (N_23866,N_23740,N_23711);
xnor U23867 (N_23867,N_23508,N_23591);
and U23868 (N_23868,N_23692,N_23659);
or U23869 (N_23869,N_23563,N_23729);
nor U23870 (N_23870,N_23649,N_23651);
xnor U23871 (N_23871,N_23534,N_23507);
nand U23872 (N_23872,N_23614,N_23732);
xnor U23873 (N_23873,N_23617,N_23705);
or U23874 (N_23874,N_23525,N_23592);
xnor U23875 (N_23875,N_23559,N_23712);
or U23876 (N_23876,N_23739,N_23736);
nand U23877 (N_23877,N_23564,N_23616);
and U23878 (N_23878,N_23600,N_23692);
and U23879 (N_23879,N_23549,N_23711);
or U23880 (N_23880,N_23570,N_23641);
or U23881 (N_23881,N_23514,N_23529);
nor U23882 (N_23882,N_23564,N_23647);
nand U23883 (N_23883,N_23736,N_23595);
nand U23884 (N_23884,N_23553,N_23640);
or U23885 (N_23885,N_23546,N_23619);
and U23886 (N_23886,N_23647,N_23603);
and U23887 (N_23887,N_23541,N_23679);
nor U23888 (N_23888,N_23621,N_23539);
xor U23889 (N_23889,N_23538,N_23666);
nor U23890 (N_23890,N_23624,N_23533);
nand U23891 (N_23891,N_23657,N_23638);
nor U23892 (N_23892,N_23670,N_23606);
nand U23893 (N_23893,N_23508,N_23531);
nand U23894 (N_23894,N_23581,N_23585);
nand U23895 (N_23895,N_23501,N_23537);
nand U23896 (N_23896,N_23706,N_23571);
and U23897 (N_23897,N_23534,N_23719);
or U23898 (N_23898,N_23618,N_23585);
or U23899 (N_23899,N_23617,N_23650);
xor U23900 (N_23900,N_23730,N_23544);
nand U23901 (N_23901,N_23734,N_23594);
nand U23902 (N_23902,N_23722,N_23737);
or U23903 (N_23903,N_23639,N_23508);
or U23904 (N_23904,N_23732,N_23646);
and U23905 (N_23905,N_23630,N_23697);
or U23906 (N_23906,N_23726,N_23645);
or U23907 (N_23907,N_23740,N_23560);
and U23908 (N_23908,N_23535,N_23615);
and U23909 (N_23909,N_23505,N_23704);
or U23910 (N_23910,N_23533,N_23598);
xor U23911 (N_23911,N_23606,N_23548);
xor U23912 (N_23912,N_23712,N_23569);
xnor U23913 (N_23913,N_23739,N_23710);
nor U23914 (N_23914,N_23654,N_23729);
and U23915 (N_23915,N_23526,N_23562);
xnor U23916 (N_23916,N_23590,N_23631);
or U23917 (N_23917,N_23731,N_23566);
xnor U23918 (N_23918,N_23692,N_23596);
or U23919 (N_23919,N_23693,N_23603);
nor U23920 (N_23920,N_23518,N_23669);
and U23921 (N_23921,N_23556,N_23554);
nand U23922 (N_23922,N_23634,N_23584);
nand U23923 (N_23923,N_23746,N_23697);
and U23924 (N_23924,N_23645,N_23552);
nand U23925 (N_23925,N_23538,N_23510);
and U23926 (N_23926,N_23569,N_23542);
nor U23927 (N_23927,N_23721,N_23590);
xnor U23928 (N_23928,N_23731,N_23644);
or U23929 (N_23929,N_23590,N_23686);
or U23930 (N_23930,N_23640,N_23741);
or U23931 (N_23931,N_23739,N_23729);
nor U23932 (N_23932,N_23617,N_23532);
xnor U23933 (N_23933,N_23528,N_23670);
nor U23934 (N_23934,N_23551,N_23601);
xnor U23935 (N_23935,N_23746,N_23524);
xor U23936 (N_23936,N_23537,N_23532);
or U23937 (N_23937,N_23640,N_23675);
or U23938 (N_23938,N_23658,N_23717);
nand U23939 (N_23939,N_23548,N_23523);
and U23940 (N_23940,N_23505,N_23606);
nand U23941 (N_23941,N_23700,N_23735);
or U23942 (N_23942,N_23705,N_23517);
nand U23943 (N_23943,N_23530,N_23622);
xnor U23944 (N_23944,N_23735,N_23644);
or U23945 (N_23945,N_23718,N_23576);
xnor U23946 (N_23946,N_23731,N_23625);
or U23947 (N_23947,N_23543,N_23671);
nand U23948 (N_23948,N_23661,N_23617);
xnor U23949 (N_23949,N_23543,N_23724);
or U23950 (N_23950,N_23614,N_23608);
and U23951 (N_23951,N_23675,N_23570);
nand U23952 (N_23952,N_23625,N_23556);
and U23953 (N_23953,N_23748,N_23741);
nor U23954 (N_23954,N_23723,N_23738);
or U23955 (N_23955,N_23714,N_23504);
nor U23956 (N_23956,N_23547,N_23552);
nor U23957 (N_23957,N_23637,N_23570);
or U23958 (N_23958,N_23663,N_23731);
nor U23959 (N_23959,N_23664,N_23732);
xor U23960 (N_23960,N_23544,N_23650);
nor U23961 (N_23961,N_23612,N_23533);
nor U23962 (N_23962,N_23638,N_23695);
and U23963 (N_23963,N_23561,N_23563);
and U23964 (N_23964,N_23744,N_23632);
xor U23965 (N_23965,N_23519,N_23560);
nor U23966 (N_23966,N_23680,N_23632);
xnor U23967 (N_23967,N_23709,N_23668);
and U23968 (N_23968,N_23734,N_23502);
nor U23969 (N_23969,N_23624,N_23599);
nand U23970 (N_23970,N_23575,N_23723);
nand U23971 (N_23971,N_23651,N_23637);
or U23972 (N_23972,N_23506,N_23655);
xnor U23973 (N_23973,N_23668,N_23529);
nor U23974 (N_23974,N_23729,N_23514);
and U23975 (N_23975,N_23559,N_23604);
and U23976 (N_23976,N_23643,N_23717);
nor U23977 (N_23977,N_23553,N_23508);
or U23978 (N_23978,N_23599,N_23523);
nor U23979 (N_23979,N_23722,N_23618);
or U23980 (N_23980,N_23737,N_23502);
or U23981 (N_23981,N_23744,N_23634);
and U23982 (N_23982,N_23507,N_23663);
or U23983 (N_23983,N_23655,N_23569);
xnor U23984 (N_23984,N_23618,N_23514);
and U23985 (N_23985,N_23624,N_23550);
nor U23986 (N_23986,N_23549,N_23555);
nor U23987 (N_23987,N_23721,N_23694);
and U23988 (N_23988,N_23682,N_23508);
and U23989 (N_23989,N_23678,N_23728);
nand U23990 (N_23990,N_23646,N_23689);
nor U23991 (N_23991,N_23536,N_23550);
nor U23992 (N_23992,N_23724,N_23561);
nor U23993 (N_23993,N_23574,N_23522);
nand U23994 (N_23994,N_23700,N_23605);
nor U23995 (N_23995,N_23694,N_23503);
nand U23996 (N_23996,N_23589,N_23542);
xor U23997 (N_23997,N_23710,N_23655);
nand U23998 (N_23998,N_23661,N_23536);
or U23999 (N_23999,N_23608,N_23723);
nand U24000 (N_24000,N_23805,N_23752);
xnor U24001 (N_24001,N_23767,N_23867);
and U24002 (N_24002,N_23913,N_23911);
and U24003 (N_24003,N_23807,N_23923);
nor U24004 (N_24004,N_23966,N_23936);
and U24005 (N_24005,N_23991,N_23922);
or U24006 (N_24006,N_23789,N_23770);
and U24007 (N_24007,N_23829,N_23916);
or U24008 (N_24008,N_23880,N_23924);
xor U24009 (N_24009,N_23802,N_23878);
and U24010 (N_24010,N_23840,N_23946);
or U24011 (N_24011,N_23845,N_23952);
nor U24012 (N_24012,N_23915,N_23876);
nor U24013 (N_24013,N_23885,N_23989);
and U24014 (N_24014,N_23831,N_23959);
nand U24015 (N_24015,N_23781,N_23926);
nand U24016 (N_24016,N_23943,N_23983);
and U24017 (N_24017,N_23753,N_23996);
xnor U24018 (N_24018,N_23920,N_23758);
and U24019 (N_24019,N_23814,N_23759);
xor U24020 (N_24020,N_23775,N_23875);
or U24021 (N_24021,N_23799,N_23750);
or U24022 (N_24022,N_23882,N_23955);
nor U24023 (N_24023,N_23999,N_23965);
or U24024 (N_24024,N_23854,N_23801);
nor U24025 (N_24025,N_23968,N_23891);
or U24026 (N_24026,N_23818,N_23815);
xor U24027 (N_24027,N_23768,N_23905);
nor U24028 (N_24028,N_23763,N_23974);
nor U24029 (N_24029,N_23964,N_23914);
and U24030 (N_24030,N_23994,N_23844);
nand U24031 (N_24031,N_23798,N_23860);
nand U24032 (N_24032,N_23884,N_23949);
nor U24033 (N_24033,N_23843,N_23997);
nand U24034 (N_24034,N_23881,N_23821);
xor U24035 (N_24035,N_23765,N_23907);
nor U24036 (N_24036,N_23836,N_23795);
xnor U24037 (N_24037,N_23823,N_23981);
and U24038 (N_24038,N_23896,N_23998);
nor U24039 (N_24039,N_23898,N_23866);
xnor U24040 (N_24040,N_23925,N_23755);
xor U24041 (N_24041,N_23954,N_23837);
and U24042 (N_24042,N_23816,N_23901);
and U24043 (N_24043,N_23903,N_23848);
or U24044 (N_24044,N_23811,N_23899);
xnor U24045 (N_24045,N_23838,N_23892);
or U24046 (N_24046,N_23963,N_23842);
xnor U24047 (N_24047,N_23919,N_23774);
nand U24048 (N_24048,N_23872,N_23921);
xor U24049 (N_24049,N_23810,N_23786);
xor U24050 (N_24050,N_23904,N_23857);
xor U24051 (N_24051,N_23850,N_23822);
nand U24052 (N_24052,N_23797,N_23819);
or U24053 (N_24053,N_23883,N_23825);
nor U24054 (N_24054,N_23993,N_23820);
xnor U24055 (N_24055,N_23900,N_23785);
and U24056 (N_24056,N_23947,N_23769);
nor U24057 (N_24057,N_23957,N_23894);
xnor U24058 (N_24058,N_23986,N_23934);
nor U24059 (N_24059,N_23929,N_23931);
nand U24060 (N_24060,N_23958,N_23933);
nor U24061 (N_24061,N_23912,N_23779);
nand U24062 (N_24062,N_23791,N_23794);
or U24063 (N_24063,N_23942,N_23841);
or U24064 (N_24064,N_23826,N_23897);
nand U24065 (N_24065,N_23908,N_23978);
and U24066 (N_24066,N_23888,N_23972);
and U24067 (N_24067,N_23887,N_23889);
nor U24068 (N_24068,N_23773,N_23960);
nor U24069 (N_24069,N_23839,N_23828);
and U24070 (N_24070,N_23856,N_23778);
nor U24071 (N_24071,N_23893,N_23944);
xnor U24072 (N_24072,N_23868,N_23865);
nor U24073 (N_24073,N_23935,N_23995);
and U24074 (N_24074,N_23890,N_23772);
xnor U24075 (N_24075,N_23754,N_23776);
nor U24076 (N_24076,N_23762,N_23792);
xor U24077 (N_24077,N_23852,N_23832);
nor U24078 (N_24078,N_23800,N_23777);
nor U24079 (N_24079,N_23979,N_23855);
xnor U24080 (N_24080,N_23862,N_23962);
nand U24081 (N_24081,N_23859,N_23910);
or U24082 (N_24082,N_23938,N_23809);
xor U24083 (N_24083,N_23967,N_23812);
nor U24084 (N_24084,N_23847,N_23956);
and U24085 (N_24085,N_23757,N_23756);
and U24086 (N_24086,N_23760,N_23951);
nor U24087 (N_24087,N_23858,N_23988);
and U24088 (N_24088,N_23793,N_23917);
xor U24089 (N_24089,N_23784,N_23782);
nand U24090 (N_24090,N_23930,N_23751);
or U24091 (N_24091,N_23873,N_23813);
and U24092 (N_24092,N_23928,N_23830);
xnor U24093 (N_24093,N_23940,N_23853);
xnor U24094 (N_24094,N_23980,N_23824);
nor U24095 (N_24095,N_23970,N_23804);
and U24096 (N_24096,N_23817,N_23941);
and U24097 (N_24097,N_23953,N_23864);
or U24098 (N_24098,N_23909,N_23886);
nor U24099 (N_24099,N_23990,N_23937);
and U24100 (N_24100,N_23877,N_23796);
xnor U24101 (N_24101,N_23992,N_23808);
and U24102 (N_24102,N_23846,N_23788);
xnor U24103 (N_24103,N_23803,N_23871);
xor U24104 (N_24104,N_23835,N_23787);
nor U24105 (N_24105,N_23948,N_23961);
and U24106 (N_24106,N_23870,N_23827);
nand U24107 (N_24107,N_23780,N_23764);
nor U24108 (N_24108,N_23977,N_23761);
nor U24109 (N_24109,N_23976,N_23879);
or U24110 (N_24110,N_23790,N_23973);
or U24111 (N_24111,N_23895,N_23971);
or U24112 (N_24112,N_23939,N_23918);
and U24113 (N_24113,N_23833,N_23834);
and U24114 (N_24114,N_23861,N_23975);
nor U24115 (N_24115,N_23984,N_23927);
xor U24116 (N_24116,N_23906,N_23982);
nor U24117 (N_24117,N_23771,N_23985);
xor U24118 (N_24118,N_23863,N_23987);
or U24119 (N_24119,N_23945,N_23950);
or U24120 (N_24120,N_23932,N_23902);
nand U24121 (N_24121,N_23806,N_23969);
nand U24122 (N_24122,N_23849,N_23869);
xnor U24123 (N_24123,N_23783,N_23766);
or U24124 (N_24124,N_23874,N_23851);
nand U24125 (N_24125,N_23975,N_23787);
xnor U24126 (N_24126,N_23987,N_23866);
xnor U24127 (N_24127,N_23766,N_23934);
and U24128 (N_24128,N_23941,N_23795);
or U24129 (N_24129,N_23963,N_23856);
and U24130 (N_24130,N_23803,N_23983);
and U24131 (N_24131,N_23867,N_23832);
xor U24132 (N_24132,N_23808,N_23987);
xor U24133 (N_24133,N_23973,N_23990);
and U24134 (N_24134,N_23775,N_23876);
nand U24135 (N_24135,N_23944,N_23920);
xnor U24136 (N_24136,N_23845,N_23935);
nand U24137 (N_24137,N_23785,N_23853);
xor U24138 (N_24138,N_23957,N_23757);
or U24139 (N_24139,N_23815,N_23788);
nand U24140 (N_24140,N_23851,N_23961);
nand U24141 (N_24141,N_23906,N_23940);
and U24142 (N_24142,N_23958,N_23989);
nor U24143 (N_24143,N_23856,N_23802);
nand U24144 (N_24144,N_23893,N_23964);
or U24145 (N_24145,N_23993,N_23882);
xor U24146 (N_24146,N_23950,N_23784);
nand U24147 (N_24147,N_23839,N_23988);
xnor U24148 (N_24148,N_23868,N_23871);
or U24149 (N_24149,N_23851,N_23981);
nand U24150 (N_24150,N_23969,N_23893);
nor U24151 (N_24151,N_23978,N_23861);
and U24152 (N_24152,N_23784,N_23958);
nor U24153 (N_24153,N_23945,N_23924);
or U24154 (N_24154,N_23803,N_23787);
nand U24155 (N_24155,N_23862,N_23808);
nand U24156 (N_24156,N_23856,N_23982);
and U24157 (N_24157,N_23910,N_23893);
xor U24158 (N_24158,N_23833,N_23777);
or U24159 (N_24159,N_23994,N_23961);
or U24160 (N_24160,N_23906,N_23763);
nor U24161 (N_24161,N_23945,N_23898);
nor U24162 (N_24162,N_23834,N_23827);
nor U24163 (N_24163,N_23839,N_23915);
xor U24164 (N_24164,N_23825,N_23765);
xnor U24165 (N_24165,N_23971,N_23813);
nor U24166 (N_24166,N_23861,N_23784);
nor U24167 (N_24167,N_23978,N_23761);
and U24168 (N_24168,N_23859,N_23922);
nor U24169 (N_24169,N_23768,N_23981);
nor U24170 (N_24170,N_23939,N_23805);
xnor U24171 (N_24171,N_23776,N_23923);
nor U24172 (N_24172,N_23831,N_23995);
nand U24173 (N_24173,N_23768,N_23791);
nand U24174 (N_24174,N_23982,N_23821);
nor U24175 (N_24175,N_23768,N_23771);
nand U24176 (N_24176,N_23871,N_23988);
nand U24177 (N_24177,N_23806,N_23785);
xor U24178 (N_24178,N_23914,N_23872);
nor U24179 (N_24179,N_23962,N_23863);
or U24180 (N_24180,N_23809,N_23936);
nand U24181 (N_24181,N_23802,N_23860);
nor U24182 (N_24182,N_23766,N_23994);
or U24183 (N_24183,N_23827,N_23957);
and U24184 (N_24184,N_23845,N_23775);
or U24185 (N_24185,N_23967,N_23847);
nand U24186 (N_24186,N_23771,N_23904);
or U24187 (N_24187,N_23864,N_23942);
or U24188 (N_24188,N_23956,N_23860);
and U24189 (N_24189,N_23791,N_23786);
nand U24190 (N_24190,N_23849,N_23848);
or U24191 (N_24191,N_23805,N_23975);
or U24192 (N_24192,N_23840,N_23992);
nor U24193 (N_24193,N_23937,N_23944);
or U24194 (N_24194,N_23988,N_23867);
or U24195 (N_24195,N_23807,N_23817);
nand U24196 (N_24196,N_23778,N_23849);
or U24197 (N_24197,N_23800,N_23776);
or U24198 (N_24198,N_23761,N_23773);
nor U24199 (N_24199,N_23956,N_23906);
xnor U24200 (N_24200,N_23768,N_23909);
nor U24201 (N_24201,N_23923,N_23813);
or U24202 (N_24202,N_23955,N_23789);
xnor U24203 (N_24203,N_23795,N_23991);
or U24204 (N_24204,N_23787,N_23938);
xor U24205 (N_24205,N_23796,N_23960);
nor U24206 (N_24206,N_23970,N_23805);
xnor U24207 (N_24207,N_23847,N_23825);
nor U24208 (N_24208,N_23857,N_23823);
and U24209 (N_24209,N_23985,N_23890);
and U24210 (N_24210,N_23889,N_23876);
nand U24211 (N_24211,N_23795,N_23756);
xnor U24212 (N_24212,N_23867,N_23774);
nor U24213 (N_24213,N_23802,N_23828);
xor U24214 (N_24214,N_23933,N_23988);
nor U24215 (N_24215,N_23933,N_23801);
and U24216 (N_24216,N_23815,N_23843);
nor U24217 (N_24217,N_23759,N_23945);
xor U24218 (N_24218,N_23799,N_23873);
nand U24219 (N_24219,N_23812,N_23871);
xor U24220 (N_24220,N_23922,N_23805);
nor U24221 (N_24221,N_23979,N_23947);
xor U24222 (N_24222,N_23901,N_23977);
xnor U24223 (N_24223,N_23997,N_23770);
or U24224 (N_24224,N_23847,N_23856);
nor U24225 (N_24225,N_23820,N_23758);
or U24226 (N_24226,N_23934,N_23867);
or U24227 (N_24227,N_23862,N_23795);
xnor U24228 (N_24228,N_23826,N_23822);
and U24229 (N_24229,N_23935,N_23801);
or U24230 (N_24230,N_23986,N_23985);
nor U24231 (N_24231,N_23851,N_23963);
and U24232 (N_24232,N_23867,N_23993);
xnor U24233 (N_24233,N_23969,N_23910);
nand U24234 (N_24234,N_23927,N_23921);
or U24235 (N_24235,N_23754,N_23857);
nor U24236 (N_24236,N_23767,N_23928);
and U24237 (N_24237,N_23938,N_23765);
and U24238 (N_24238,N_23978,N_23896);
or U24239 (N_24239,N_23896,N_23968);
nand U24240 (N_24240,N_23800,N_23851);
or U24241 (N_24241,N_23751,N_23939);
and U24242 (N_24242,N_23923,N_23868);
or U24243 (N_24243,N_23891,N_23959);
nand U24244 (N_24244,N_23857,N_23756);
nor U24245 (N_24245,N_23795,N_23958);
xnor U24246 (N_24246,N_23769,N_23973);
and U24247 (N_24247,N_23798,N_23942);
nor U24248 (N_24248,N_23813,N_23927);
xnor U24249 (N_24249,N_23930,N_23928);
and U24250 (N_24250,N_24188,N_24238);
or U24251 (N_24251,N_24209,N_24096);
nor U24252 (N_24252,N_24142,N_24053);
xnor U24253 (N_24253,N_24134,N_24018);
and U24254 (N_24254,N_24163,N_24225);
and U24255 (N_24255,N_24130,N_24110);
nand U24256 (N_24256,N_24167,N_24005);
and U24257 (N_24257,N_24204,N_24194);
nand U24258 (N_24258,N_24003,N_24056);
nor U24259 (N_24259,N_24216,N_24229);
nand U24260 (N_24260,N_24081,N_24201);
nand U24261 (N_24261,N_24135,N_24121);
nor U24262 (N_24262,N_24128,N_24249);
nor U24263 (N_24263,N_24217,N_24078);
and U24264 (N_24264,N_24024,N_24234);
or U24265 (N_24265,N_24035,N_24191);
nand U24266 (N_24266,N_24155,N_24162);
and U24267 (N_24267,N_24073,N_24231);
or U24268 (N_24268,N_24021,N_24176);
or U24269 (N_24269,N_24108,N_24222);
nand U24270 (N_24270,N_24186,N_24020);
nand U24271 (N_24271,N_24170,N_24182);
nand U24272 (N_24272,N_24175,N_24232);
xnor U24273 (N_24273,N_24092,N_24240);
and U24274 (N_24274,N_24242,N_24164);
or U24275 (N_24275,N_24178,N_24214);
nor U24276 (N_24276,N_24193,N_24016);
and U24277 (N_24277,N_24027,N_24028);
and U24278 (N_24278,N_24051,N_24014);
and U24279 (N_24279,N_24023,N_24116);
xor U24280 (N_24280,N_24086,N_24091);
xor U24281 (N_24281,N_24082,N_24127);
or U24282 (N_24282,N_24105,N_24239);
or U24283 (N_24283,N_24143,N_24150);
xor U24284 (N_24284,N_24034,N_24006);
nand U24285 (N_24285,N_24007,N_24022);
and U24286 (N_24286,N_24075,N_24119);
and U24287 (N_24287,N_24100,N_24058);
nand U24288 (N_24288,N_24198,N_24112);
nand U24289 (N_24289,N_24079,N_24185);
or U24290 (N_24290,N_24159,N_24227);
xnor U24291 (N_24291,N_24236,N_24087);
and U24292 (N_24292,N_24126,N_24088);
xnor U24293 (N_24293,N_24102,N_24174);
nand U24294 (N_24294,N_24084,N_24235);
or U24295 (N_24295,N_24136,N_24030);
nand U24296 (N_24296,N_24202,N_24036);
xor U24297 (N_24297,N_24077,N_24224);
xnor U24298 (N_24298,N_24161,N_24095);
and U24299 (N_24299,N_24085,N_24042);
and U24300 (N_24300,N_24248,N_24109);
xnor U24301 (N_24301,N_24173,N_24017);
and U24302 (N_24302,N_24057,N_24200);
nand U24303 (N_24303,N_24213,N_24152);
and U24304 (N_24304,N_24101,N_24179);
nand U24305 (N_24305,N_24004,N_24187);
nor U24306 (N_24306,N_24097,N_24064);
nor U24307 (N_24307,N_24207,N_24048);
xor U24308 (N_24308,N_24068,N_24212);
xnor U24309 (N_24309,N_24243,N_24066);
nor U24310 (N_24310,N_24197,N_24148);
and U24311 (N_24311,N_24065,N_24046);
and U24312 (N_24312,N_24153,N_24118);
nand U24313 (N_24313,N_24089,N_24050);
xnor U24314 (N_24314,N_24098,N_24129);
or U24315 (N_24315,N_24203,N_24008);
nor U24316 (N_24316,N_24009,N_24210);
and U24317 (N_24317,N_24059,N_24138);
xnor U24318 (N_24318,N_24049,N_24094);
and U24319 (N_24319,N_24149,N_24169);
and U24320 (N_24320,N_24172,N_24010);
xor U24321 (N_24321,N_24141,N_24195);
nand U24322 (N_24322,N_24183,N_24165);
nand U24323 (N_24323,N_24111,N_24133);
or U24324 (N_24324,N_24072,N_24223);
nor U24325 (N_24325,N_24060,N_24147);
and U24326 (N_24326,N_24052,N_24026);
and U24327 (N_24327,N_24139,N_24039);
xor U24328 (N_24328,N_24074,N_24171);
nor U24329 (N_24329,N_24192,N_24033);
nor U24330 (N_24330,N_24221,N_24124);
xnor U24331 (N_24331,N_24043,N_24069);
or U24332 (N_24332,N_24241,N_24038);
nand U24333 (N_24333,N_24137,N_24206);
or U24334 (N_24334,N_24047,N_24146);
nand U24335 (N_24335,N_24032,N_24168);
nand U24336 (N_24336,N_24166,N_24011);
xnor U24337 (N_24337,N_24040,N_24113);
nor U24338 (N_24338,N_24031,N_24237);
nor U24339 (N_24339,N_24070,N_24189);
nand U24340 (N_24340,N_24067,N_24123);
nor U24341 (N_24341,N_24120,N_24117);
nor U24342 (N_24342,N_24199,N_24080);
nand U24343 (N_24343,N_24157,N_24054);
nand U24344 (N_24344,N_24103,N_24190);
nand U24345 (N_24345,N_24037,N_24158);
nor U24346 (N_24346,N_24132,N_24001);
nor U24347 (N_24347,N_24041,N_24145);
and U24348 (N_24348,N_24228,N_24215);
xor U24349 (N_24349,N_24083,N_24012);
xnor U24350 (N_24350,N_24205,N_24226);
or U24351 (N_24351,N_24002,N_24115);
xor U24352 (N_24352,N_24044,N_24093);
nor U24353 (N_24353,N_24076,N_24090);
xnor U24354 (N_24354,N_24230,N_24099);
or U24355 (N_24355,N_24131,N_24208);
nor U24356 (N_24356,N_24061,N_24140);
nor U24357 (N_24357,N_24196,N_24063);
and U24358 (N_24358,N_24246,N_24154);
nand U24359 (N_24359,N_24122,N_24156);
nand U24360 (N_24360,N_24181,N_24114);
xor U24361 (N_24361,N_24045,N_24144);
xnor U24362 (N_24362,N_24125,N_24071);
and U24363 (N_24363,N_24211,N_24245);
xnor U24364 (N_24364,N_24180,N_24019);
nand U24365 (N_24365,N_24029,N_24160);
and U24366 (N_24366,N_24218,N_24000);
nor U24367 (N_24367,N_24184,N_24219);
and U24368 (N_24368,N_24247,N_24220);
nor U24369 (N_24369,N_24244,N_24015);
and U24370 (N_24370,N_24055,N_24062);
and U24371 (N_24371,N_24233,N_24106);
or U24372 (N_24372,N_24151,N_24025);
or U24373 (N_24373,N_24104,N_24107);
and U24374 (N_24374,N_24177,N_24013);
and U24375 (N_24375,N_24218,N_24220);
and U24376 (N_24376,N_24199,N_24060);
nor U24377 (N_24377,N_24247,N_24107);
or U24378 (N_24378,N_24025,N_24198);
or U24379 (N_24379,N_24044,N_24159);
xnor U24380 (N_24380,N_24158,N_24040);
or U24381 (N_24381,N_24097,N_24153);
or U24382 (N_24382,N_24107,N_24166);
and U24383 (N_24383,N_24120,N_24159);
nand U24384 (N_24384,N_24186,N_24168);
and U24385 (N_24385,N_24248,N_24110);
xnor U24386 (N_24386,N_24193,N_24062);
nand U24387 (N_24387,N_24131,N_24231);
xor U24388 (N_24388,N_24060,N_24208);
nand U24389 (N_24389,N_24196,N_24152);
nor U24390 (N_24390,N_24114,N_24167);
nand U24391 (N_24391,N_24003,N_24241);
or U24392 (N_24392,N_24241,N_24121);
xor U24393 (N_24393,N_24072,N_24070);
nand U24394 (N_24394,N_24191,N_24112);
nand U24395 (N_24395,N_24027,N_24208);
xor U24396 (N_24396,N_24188,N_24024);
nand U24397 (N_24397,N_24118,N_24103);
xor U24398 (N_24398,N_24126,N_24112);
xor U24399 (N_24399,N_24099,N_24014);
and U24400 (N_24400,N_24162,N_24085);
and U24401 (N_24401,N_24233,N_24172);
nor U24402 (N_24402,N_24108,N_24188);
and U24403 (N_24403,N_24187,N_24155);
nor U24404 (N_24404,N_24015,N_24068);
or U24405 (N_24405,N_24184,N_24122);
and U24406 (N_24406,N_24242,N_24073);
or U24407 (N_24407,N_24051,N_24176);
nand U24408 (N_24408,N_24148,N_24006);
xnor U24409 (N_24409,N_24074,N_24234);
or U24410 (N_24410,N_24164,N_24122);
nand U24411 (N_24411,N_24018,N_24078);
nand U24412 (N_24412,N_24139,N_24031);
xor U24413 (N_24413,N_24096,N_24065);
xor U24414 (N_24414,N_24057,N_24076);
and U24415 (N_24415,N_24092,N_24180);
xor U24416 (N_24416,N_24205,N_24123);
and U24417 (N_24417,N_24032,N_24166);
and U24418 (N_24418,N_24126,N_24037);
nor U24419 (N_24419,N_24181,N_24069);
xor U24420 (N_24420,N_24249,N_24065);
or U24421 (N_24421,N_24078,N_24191);
nor U24422 (N_24422,N_24082,N_24003);
nand U24423 (N_24423,N_24231,N_24158);
or U24424 (N_24424,N_24062,N_24088);
nand U24425 (N_24425,N_24104,N_24125);
nor U24426 (N_24426,N_24196,N_24025);
and U24427 (N_24427,N_24168,N_24088);
and U24428 (N_24428,N_24219,N_24096);
or U24429 (N_24429,N_24117,N_24235);
xnor U24430 (N_24430,N_24071,N_24219);
xnor U24431 (N_24431,N_24081,N_24203);
nand U24432 (N_24432,N_24249,N_24237);
and U24433 (N_24433,N_24118,N_24002);
nand U24434 (N_24434,N_24156,N_24113);
or U24435 (N_24435,N_24007,N_24241);
xnor U24436 (N_24436,N_24245,N_24141);
and U24437 (N_24437,N_24249,N_24043);
xor U24438 (N_24438,N_24068,N_24000);
and U24439 (N_24439,N_24105,N_24224);
xor U24440 (N_24440,N_24044,N_24014);
nand U24441 (N_24441,N_24209,N_24147);
and U24442 (N_24442,N_24066,N_24072);
nand U24443 (N_24443,N_24066,N_24247);
xor U24444 (N_24444,N_24008,N_24089);
nand U24445 (N_24445,N_24122,N_24224);
nor U24446 (N_24446,N_24031,N_24183);
nand U24447 (N_24447,N_24030,N_24230);
xnor U24448 (N_24448,N_24201,N_24204);
and U24449 (N_24449,N_24071,N_24119);
or U24450 (N_24450,N_24007,N_24018);
and U24451 (N_24451,N_24218,N_24150);
and U24452 (N_24452,N_24157,N_24218);
or U24453 (N_24453,N_24123,N_24001);
and U24454 (N_24454,N_24133,N_24088);
nand U24455 (N_24455,N_24012,N_24118);
and U24456 (N_24456,N_24003,N_24169);
nand U24457 (N_24457,N_24225,N_24191);
xnor U24458 (N_24458,N_24232,N_24160);
nand U24459 (N_24459,N_24082,N_24166);
or U24460 (N_24460,N_24221,N_24174);
nor U24461 (N_24461,N_24100,N_24218);
and U24462 (N_24462,N_24132,N_24049);
xnor U24463 (N_24463,N_24059,N_24151);
nand U24464 (N_24464,N_24105,N_24146);
and U24465 (N_24465,N_24151,N_24004);
nand U24466 (N_24466,N_24031,N_24103);
and U24467 (N_24467,N_24221,N_24095);
nor U24468 (N_24468,N_24049,N_24110);
nor U24469 (N_24469,N_24126,N_24169);
and U24470 (N_24470,N_24067,N_24120);
and U24471 (N_24471,N_24239,N_24015);
and U24472 (N_24472,N_24229,N_24196);
or U24473 (N_24473,N_24189,N_24123);
xnor U24474 (N_24474,N_24113,N_24124);
xor U24475 (N_24475,N_24195,N_24112);
xor U24476 (N_24476,N_24235,N_24197);
and U24477 (N_24477,N_24088,N_24218);
and U24478 (N_24478,N_24152,N_24083);
xor U24479 (N_24479,N_24109,N_24066);
xnor U24480 (N_24480,N_24146,N_24244);
nor U24481 (N_24481,N_24225,N_24229);
nor U24482 (N_24482,N_24009,N_24241);
and U24483 (N_24483,N_24125,N_24004);
nor U24484 (N_24484,N_24071,N_24012);
xor U24485 (N_24485,N_24170,N_24103);
and U24486 (N_24486,N_24208,N_24124);
nand U24487 (N_24487,N_24053,N_24170);
or U24488 (N_24488,N_24194,N_24008);
xor U24489 (N_24489,N_24234,N_24071);
and U24490 (N_24490,N_24093,N_24102);
or U24491 (N_24491,N_24028,N_24070);
or U24492 (N_24492,N_24232,N_24130);
or U24493 (N_24493,N_24034,N_24195);
or U24494 (N_24494,N_24115,N_24193);
xnor U24495 (N_24495,N_24099,N_24036);
xor U24496 (N_24496,N_24090,N_24029);
and U24497 (N_24497,N_24156,N_24079);
xnor U24498 (N_24498,N_24102,N_24159);
nor U24499 (N_24499,N_24104,N_24142);
xor U24500 (N_24500,N_24278,N_24390);
nand U24501 (N_24501,N_24446,N_24294);
or U24502 (N_24502,N_24256,N_24462);
xnor U24503 (N_24503,N_24250,N_24347);
nand U24504 (N_24504,N_24405,N_24366);
nand U24505 (N_24505,N_24438,N_24391);
nor U24506 (N_24506,N_24287,N_24422);
and U24507 (N_24507,N_24376,N_24400);
nor U24508 (N_24508,N_24404,N_24309);
xor U24509 (N_24509,N_24358,N_24341);
or U24510 (N_24510,N_24316,N_24328);
xor U24511 (N_24511,N_24477,N_24353);
or U24512 (N_24512,N_24291,N_24401);
nor U24513 (N_24513,N_24361,N_24421);
nand U24514 (N_24514,N_24416,N_24420);
nor U24515 (N_24515,N_24425,N_24266);
xor U24516 (N_24516,N_24465,N_24355);
nor U24517 (N_24517,N_24293,N_24498);
xor U24518 (N_24518,N_24299,N_24359);
and U24519 (N_24519,N_24327,N_24488);
nor U24520 (N_24520,N_24267,N_24490);
nor U24521 (N_24521,N_24472,N_24264);
nand U24522 (N_24522,N_24298,N_24292);
nor U24523 (N_24523,N_24460,N_24286);
nand U24524 (N_24524,N_24356,N_24411);
xor U24525 (N_24525,N_24285,N_24354);
nor U24526 (N_24526,N_24445,N_24275);
and U24527 (N_24527,N_24379,N_24423);
xor U24528 (N_24528,N_24461,N_24373);
nor U24529 (N_24529,N_24319,N_24324);
xor U24530 (N_24530,N_24305,N_24268);
xnor U24531 (N_24531,N_24351,N_24381);
or U24532 (N_24532,N_24413,N_24282);
and U24533 (N_24533,N_24451,N_24474);
and U24534 (N_24534,N_24393,N_24463);
nor U24535 (N_24535,N_24396,N_24295);
and U24536 (N_24536,N_24442,N_24457);
or U24537 (N_24537,N_24310,N_24435);
or U24538 (N_24538,N_24406,N_24473);
and U24539 (N_24539,N_24350,N_24377);
nand U24540 (N_24540,N_24434,N_24251);
nand U24541 (N_24541,N_24408,N_24453);
nor U24542 (N_24542,N_24270,N_24260);
nand U24543 (N_24543,N_24429,N_24253);
xnor U24544 (N_24544,N_24397,N_24357);
or U24545 (N_24545,N_24458,N_24304);
or U24546 (N_24546,N_24367,N_24449);
xor U24547 (N_24547,N_24448,N_24279);
nand U24548 (N_24548,N_24384,N_24482);
or U24549 (N_24549,N_24339,N_24492);
xnor U24550 (N_24550,N_24255,N_24283);
xnor U24551 (N_24551,N_24464,N_24430);
nand U24552 (N_24552,N_24409,N_24300);
nand U24553 (N_24553,N_24315,N_24261);
nand U24554 (N_24554,N_24440,N_24265);
and U24555 (N_24555,N_24415,N_24399);
or U24556 (N_24556,N_24385,N_24494);
nor U24557 (N_24557,N_24343,N_24439);
or U24558 (N_24558,N_24491,N_24314);
nand U24559 (N_24559,N_24468,N_24378);
nor U24560 (N_24560,N_24333,N_24431);
nand U24561 (N_24561,N_24290,N_24368);
or U24562 (N_24562,N_24369,N_24301);
nor U24563 (N_24563,N_24363,N_24487);
and U24564 (N_24564,N_24476,N_24475);
nor U24565 (N_24565,N_24273,N_24318);
xor U24566 (N_24566,N_24447,N_24412);
and U24567 (N_24567,N_24387,N_24436);
nor U24568 (N_24568,N_24312,N_24280);
nand U24569 (N_24569,N_24484,N_24395);
nand U24570 (N_24570,N_24272,N_24276);
or U24571 (N_24571,N_24388,N_24302);
and U24572 (N_24572,N_24426,N_24394);
or U24573 (N_24573,N_24496,N_24459);
nor U24574 (N_24574,N_24345,N_24495);
or U24575 (N_24575,N_24325,N_24259);
xnor U24576 (N_24576,N_24322,N_24489);
nor U24577 (N_24577,N_24414,N_24258);
nor U24578 (N_24578,N_24284,N_24403);
nand U24579 (N_24579,N_24323,N_24469);
or U24580 (N_24580,N_24375,N_24274);
nor U24581 (N_24581,N_24340,N_24254);
or U24582 (N_24582,N_24386,N_24321);
or U24583 (N_24583,N_24263,N_24432);
xnor U24584 (N_24584,N_24452,N_24346);
and U24585 (N_24585,N_24252,N_24307);
or U24586 (N_24586,N_24437,N_24433);
or U24587 (N_24587,N_24479,N_24311);
and U24588 (N_24588,N_24398,N_24419);
and U24589 (N_24589,N_24392,N_24344);
or U24590 (N_24590,N_24456,N_24454);
and U24591 (N_24591,N_24372,N_24320);
nand U24592 (N_24592,N_24478,N_24289);
nor U24593 (N_24593,N_24360,N_24481);
and U24594 (N_24594,N_24499,N_24466);
and U24595 (N_24595,N_24296,N_24428);
nand U24596 (N_24596,N_24443,N_24371);
or U24597 (N_24597,N_24308,N_24383);
xnor U24598 (N_24598,N_24338,N_24402);
nor U24599 (N_24599,N_24483,N_24370);
nor U24600 (N_24600,N_24336,N_24332);
and U24601 (N_24601,N_24262,N_24427);
or U24602 (N_24602,N_24467,N_24329);
xnor U24603 (N_24603,N_24444,N_24364);
nand U24604 (N_24604,N_24497,N_24288);
and U24605 (N_24605,N_24257,N_24424);
or U24606 (N_24606,N_24334,N_24331);
xor U24607 (N_24607,N_24306,N_24441);
nor U24608 (N_24608,N_24493,N_24418);
nor U24609 (N_24609,N_24410,N_24389);
nand U24610 (N_24610,N_24471,N_24365);
nor U24611 (N_24611,N_24303,N_24317);
nor U24612 (N_24612,N_24271,N_24352);
nor U24613 (N_24613,N_24313,N_24337);
or U24614 (N_24614,N_24485,N_24417);
xnor U24615 (N_24615,N_24335,N_24382);
and U24616 (N_24616,N_24281,N_24269);
or U24617 (N_24617,N_24450,N_24349);
or U24618 (N_24618,N_24277,N_24362);
or U24619 (N_24619,N_24455,N_24486);
xnor U24620 (N_24620,N_24380,N_24470);
or U24621 (N_24621,N_24374,N_24407);
nor U24622 (N_24622,N_24297,N_24330);
nor U24623 (N_24623,N_24480,N_24326);
or U24624 (N_24624,N_24342,N_24348);
xnor U24625 (N_24625,N_24340,N_24380);
nor U24626 (N_24626,N_24277,N_24265);
nand U24627 (N_24627,N_24271,N_24449);
xor U24628 (N_24628,N_24433,N_24405);
or U24629 (N_24629,N_24337,N_24319);
and U24630 (N_24630,N_24338,N_24421);
xnor U24631 (N_24631,N_24438,N_24250);
nor U24632 (N_24632,N_24374,N_24494);
xor U24633 (N_24633,N_24363,N_24271);
xnor U24634 (N_24634,N_24324,N_24300);
xnor U24635 (N_24635,N_24271,N_24390);
and U24636 (N_24636,N_24360,N_24412);
or U24637 (N_24637,N_24359,N_24306);
nor U24638 (N_24638,N_24354,N_24297);
nor U24639 (N_24639,N_24321,N_24289);
nand U24640 (N_24640,N_24408,N_24311);
nor U24641 (N_24641,N_24267,N_24394);
or U24642 (N_24642,N_24456,N_24368);
xnor U24643 (N_24643,N_24438,N_24375);
nor U24644 (N_24644,N_24423,N_24358);
xor U24645 (N_24645,N_24350,N_24277);
nor U24646 (N_24646,N_24287,N_24284);
xor U24647 (N_24647,N_24454,N_24363);
nor U24648 (N_24648,N_24384,N_24418);
and U24649 (N_24649,N_24417,N_24424);
nor U24650 (N_24650,N_24436,N_24320);
nand U24651 (N_24651,N_24439,N_24304);
xnor U24652 (N_24652,N_24342,N_24391);
nor U24653 (N_24653,N_24437,N_24367);
nand U24654 (N_24654,N_24473,N_24400);
nand U24655 (N_24655,N_24471,N_24278);
nor U24656 (N_24656,N_24485,N_24388);
nand U24657 (N_24657,N_24284,N_24358);
or U24658 (N_24658,N_24441,N_24277);
nor U24659 (N_24659,N_24417,N_24395);
or U24660 (N_24660,N_24488,N_24420);
or U24661 (N_24661,N_24341,N_24277);
nor U24662 (N_24662,N_24273,N_24411);
or U24663 (N_24663,N_24297,N_24498);
xnor U24664 (N_24664,N_24408,N_24435);
nor U24665 (N_24665,N_24351,N_24378);
nand U24666 (N_24666,N_24280,N_24454);
xor U24667 (N_24667,N_24431,N_24449);
xnor U24668 (N_24668,N_24300,N_24452);
and U24669 (N_24669,N_24443,N_24457);
xnor U24670 (N_24670,N_24263,N_24304);
or U24671 (N_24671,N_24287,N_24257);
xor U24672 (N_24672,N_24457,N_24400);
nor U24673 (N_24673,N_24250,N_24444);
or U24674 (N_24674,N_24272,N_24428);
and U24675 (N_24675,N_24346,N_24353);
or U24676 (N_24676,N_24327,N_24373);
or U24677 (N_24677,N_24319,N_24461);
and U24678 (N_24678,N_24313,N_24391);
and U24679 (N_24679,N_24443,N_24259);
or U24680 (N_24680,N_24407,N_24252);
nand U24681 (N_24681,N_24453,N_24373);
nand U24682 (N_24682,N_24386,N_24363);
nand U24683 (N_24683,N_24410,N_24309);
xor U24684 (N_24684,N_24425,N_24495);
nand U24685 (N_24685,N_24383,N_24296);
or U24686 (N_24686,N_24271,N_24497);
and U24687 (N_24687,N_24370,N_24291);
nor U24688 (N_24688,N_24260,N_24344);
nor U24689 (N_24689,N_24349,N_24424);
nand U24690 (N_24690,N_24499,N_24477);
xor U24691 (N_24691,N_24481,N_24445);
xnor U24692 (N_24692,N_24496,N_24465);
nor U24693 (N_24693,N_24311,N_24494);
nor U24694 (N_24694,N_24344,N_24456);
and U24695 (N_24695,N_24346,N_24260);
and U24696 (N_24696,N_24438,N_24471);
nand U24697 (N_24697,N_24355,N_24468);
or U24698 (N_24698,N_24334,N_24326);
or U24699 (N_24699,N_24428,N_24479);
nand U24700 (N_24700,N_24361,N_24463);
nand U24701 (N_24701,N_24260,N_24250);
xnor U24702 (N_24702,N_24413,N_24378);
nand U24703 (N_24703,N_24320,N_24308);
or U24704 (N_24704,N_24266,N_24321);
xor U24705 (N_24705,N_24362,N_24356);
xor U24706 (N_24706,N_24271,N_24398);
or U24707 (N_24707,N_24440,N_24320);
or U24708 (N_24708,N_24315,N_24268);
and U24709 (N_24709,N_24440,N_24254);
nand U24710 (N_24710,N_24307,N_24427);
nand U24711 (N_24711,N_24465,N_24256);
or U24712 (N_24712,N_24312,N_24491);
nor U24713 (N_24713,N_24284,N_24312);
nand U24714 (N_24714,N_24290,N_24316);
nand U24715 (N_24715,N_24413,N_24480);
and U24716 (N_24716,N_24298,N_24383);
or U24717 (N_24717,N_24471,N_24260);
xnor U24718 (N_24718,N_24476,N_24469);
and U24719 (N_24719,N_24426,N_24332);
and U24720 (N_24720,N_24470,N_24462);
xnor U24721 (N_24721,N_24257,N_24438);
nand U24722 (N_24722,N_24470,N_24498);
and U24723 (N_24723,N_24287,N_24472);
and U24724 (N_24724,N_24490,N_24340);
and U24725 (N_24725,N_24359,N_24479);
nor U24726 (N_24726,N_24386,N_24452);
nand U24727 (N_24727,N_24430,N_24499);
and U24728 (N_24728,N_24435,N_24297);
xor U24729 (N_24729,N_24391,N_24363);
nor U24730 (N_24730,N_24499,N_24420);
or U24731 (N_24731,N_24385,N_24488);
nand U24732 (N_24732,N_24351,N_24279);
or U24733 (N_24733,N_24465,N_24477);
nor U24734 (N_24734,N_24378,N_24318);
nand U24735 (N_24735,N_24261,N_24279);
nor U24736 (N_24736,N_24441,N_24259);
xor U24737 (N_24737,N_24345,N_24356);
nand U24738 (N_24738,N_24478,N_24264);
xor U24739 (N_24739,N_24444,N_24411);
and U24740 (N_24740,N_24283,N_24370);
and U24741 (N_24741,N_24280,N_24278);
nand U24742 (N_24742,N_24283,N_24458);
or U24743 (N_24743,N_24314,N_24355);
xor U24744 (N_24744,N_24293,N_24290);
xor U24745 (N_24745,N_24347,N_24440);
nand U24746 (N_24746,N_24342,N_24311);
and U24747 (N_24747,N_24491,N_24333);
xor U24748 (N_24748,N_24385,N_24434);
nor U24749 (N_24749,N_24393,N_24477);
nand U24750 (N_24750,N_24637,N_24535);
nand U24751 (N_24751,N_24687,N_24507);
nor U24752 (N_24752,N_24677,N_24573);
nand U24753 (N_24753,N_24723,N_24736);
or U24754 (N_24754,N_24529,N_24706);
or U24755 (N_24755,N_24639,N_24608);
or U24756 (N_24756,N_24672,N_24605);
and U24757 (N_24757,N_24695,N_24577);
or U24758 (N_24758,N_24621,N_24634);
and U24759 (N_24759,N_24720,N_24597);
nor U24760 (N_24760,N_24673,N_24707);
xnor U24761 (N_24761,N_24557,N_24580);
and U24762 (N_24762,N_24700,N_24518);
xor U24763 (N_24763,N_24711,N_24603);
nand U24764 (N_24764,N_24680,N_24564);
nand U24765 (N_24765,N_24614,N_24578);
or U24766 (N_24766,N_24598,N_24519);
nand U24767 (N_24767,N_24686,N_24622);
and U24768 (N_24768,N_24737,N_24701);
and U24769 (N_24769,N_24696,N_24693);
and U24770 (N_24770,N_24531,N_24501);
or U24771 (N_24771,N_24521,N_24624);
and U24772 (N_24772,N_24604,N_24527);
and U24773 (N_24773,N_24562,N_24626);
xnor U24774 (N_24774,N_24619,N_24512);
or U24775 (N_24775,N_24589,N_24552);
nand U24776 (N_24776,N_24613,N_24666);
nor U24777 (N_24777,N_24617,N_24583);
or U24778 (N_24778,N_24620,N_24630);
nand U24779 (N_24779,N_24508,N_24709);
or U24780 (N_24780,N_24543,N_24599);
and U24781 (N_24781,N_24749,N_24533);
or U24782 (N_24782,N_24625,N_24545);
nand U24783 (N_24783,N_24675,N_24669);
and U24784 (N_24784,N_24633,N_24502);
nand U24785 (N_24785,N_24538,N_24595);
nor U24786 (N_24786,N_24635,N_24646);
or U24787 (N_24787,N_24575,N_24615);
or U24788 (N_24788,N_24593,N_24611);
nor U24789 (N_24789,N_24732,N_24657);
or U24790 (N_24790,N_24738,N_24678);
or U24791 (N_24791,N_24655,N_24641);
xnor U24792 (N_24792,N_24728,N_24618);
nor U24793 (N_24793,N_24705,N_24559);
and U24794 (N_24794,N_24713,N_24511);
nor U24795 (N_24795,N_24648,N_24550);
nand U24796 (N_24796,N_24742,N_24600);
or U24797 (N_24797,N_24532,N_24612);
and U24798 (N_24798,N_24590,N_24730);
xnor U24799 (N_24799,N_24509,N_24667);
or U24800 (N_24800,N_24747,N_24743);
or U24801 (N_24801,N_24610,N_24537);
nand U24802 (N_24802,N_24724,N_24676);
nor U24803 (N_24803,N_24722,N_24729);
xnor U24804 (N_24804,N_24748,N_24522);
xor U24805 (N_24805,N_24572,N_24636);
or U24806 (N_24806,N_24530,N_24704);
or U24807 (N_24807,N_24689,N_24524);
nand U24808 (N_24808,N_24503,N_24571);
nand U24809 (N_24809,N_24645,N_24546);
nor U24810 (N_24810,N_24607,N_24548);
xor U24811 (N_24811,N_24638,N_24744);
or U24812 (N_24812,N_24569,N_24581);
xnor U24813 (N_24813,N_24654,N_24640);
nor U24814 (N_24814,N_24682,N_24623);
xnor U24815 (N_24815,N_24651,N_24712);
xnor U24816 (N_24816,N_24555,N_24725);
nand U24817 (N_24817,N_24631,N_24733);
xor U24818 (N_24818,N_24592,N_24629);
nor U24819 (N_24819,N_24539,N_24525);
and U24820 (N_24820,N_24661,N_24544);
and U24821 (N_24821,N_24647,N_24567);
nor U24822 (N_24822,N_24560,N_24536);
nor U24823 (N_24823,N_24515,N_24591);
nor U24824 (N_24824,N_24649,N_24558);
and U24825 (N_24825,N_24516,N_24710);
and U24826 (N_24826,N_24585,N_24643);
xnor U24827 (N_24827,N_24727,N_24719);
nor U24828 (N_24828,N_24534,N_24683);
and U24829 (N_24829,N_24556,N_24684);
nand U24830 (N_24830,N_24685,N_24505);
and U24831 (N_24831,N_24692,N_24721);
nor U24832 (N_24832,N_24596,N_24734);
nor U24833 (N_24833,N_24500,N_24632);
nor U24834 (N_24834,N_24674,N_24602);
or U24835 (N_24835,N_24694,N_24691);
nor U24836 (N_24836,N_24526,N_24513);
or U24837 (N_24837,N_24670,N_24579);
and U24838 (N_24838,N_24716,N_24520);
xor U24839 (N_24839,N_24587,N_24697);
and U24840 (N_24840,N_24628,N_24627);
xnor U24841 (N_24841,N_24584,N_24594);
nor U24842 (N_24842,N_24642,N_24653);
and U24843 (N_24843,N_24745,N_24708);
nand U24844 (N_24844,N_24561,N_24662);
xnor U24845 (N_24845,N_24664,N_24650);
nand U24846 (N_24846,N_24679,N_24576);
nand U24847 (N_24847,N_24568,N_24663);
and U24848 (N_24848,N_24563,N_24659);
nand U24849 (N_24849,N_24671,N_24542);
or U24850 (N_24850,N_24735,N_24570);
nor U24851 (N_24851,N_24717,N_24616);
xnor U24852 (N_24852,N_24731,N_24718);
xnor U24853 (N_24853,N_24586,N_24681);
and U24854 (N_24854,N_24566,N_24574);
and U24855 (N_24855,N_24554,N_24739);
and U24856 (N_24856,N_24523,N_24703);
or U24857 (N_24857,N_24541,N_24652);
and U24858 (N_24858,N_24510,N_24549);
xor U24859 (N_24859,N_24506,N_24699);
nand U24860 (N_24860,N_24665,N_24702);
nand U24861 (N_24861,N_24553,N_24528);
or U24862 (N_24862,N_24658,N_24601);
xnor U24863 (N_24863,N_24565,N_24690);
xnor U24864 (N_24864,N_24540,N_24726);
nand U24865 (N_24865,N_24741,N_24668);
or U24866 (N_24866,N_24514,N_24660);
or U24867 (N_24867,N_24714,N_24746);
nor U24868 (N_24868,N_24606,N_24688);
xnor U24869 (N_24869,N_24715,N_24609);
nor U24870 (N_24870,N_24551,N_24582);
nand U24871 (N_24871,N_24644,N_24547);
nor U24872 (N_24872,N_24517,N_24504);
or U24873 (N_24873,N_24740,N_24698);
xor U24874 (N_24874,N_24656,N_24588);
nor U24875 (N_24875,N_24648,N_24682);
or U24876 (N_24876,N_24621,N_24564);
nor U24877 (N_24877,N_24624,N_24743);
xnor U24878 (N_24878,N_24535,N_24513);
nand U24879 (N_24879,N_24704,N_24730);
nor U24880 (N_24880,N_24646,N_24630);
nor U24881 (N_24881,N_24676,N_24731);
and U24882 (N_24882,N_24721,N_24578);
nand U24883 (N_24883,N_24573,N_24553);
or U24884 (N_24884,N_24623,N_24589);
or U24885 (N_24885,N_24687,N_24735);
nor U24886 (N_24886,N_24631,N_24722);
or U24887 (N_24887,N_24656,N_24643);
or U24888 (N_24888,N_24639,N_24500);
nand U24889 (N_24889,N_24656,N_24556);
and U24890 (N_24890,N_24580,N_24592);
nor U24891 (N_24891,N_24726,N_24541);
nor U24892 (N_24892,N_24505,N_24620);
nand U24893 (N_24893,N_24739,N_24683);
and U24894 (N_24894,N_24502,N_24612);
xnor U24895 (N_24895,N_24716,N_24511);
xor U24896 (N_24896,N_24531,N_24663);
nor U24897 (N_24897,N_24589,N_24616);
xnor U24898 (N_24898,N_24628,N_24563);
nor U24899 (N_24899,N_24634,N_24605);
nand U24900 (N_24900,N_24620,N_24534);
nand U24901 (N_24901,N_24689,N_24661);
xnor U24902 (N_24902,N_24570,N_24719);
nor U24903 (N_24903,N_24687,N_24682);
or U24904 (N_24904,N_24712,N_24593);
or U24905 (N_24905,N_24530,N_24674);
xnor U24906 (N_24906,N_24676,N_24684);
nand U24907 (N_24907,N_24701,N_24643);
xor U24908 (N_24908,N_24564,N_24515);
nor U24909 (N_24909,N_24556,N_24508);
and U24910 (N_24910,N_24516,N_24690);
nand U24911 (N_24911,N_24539,N_24651);
or U24912 (N_24912,N_24700,N_24717);
xor U24913 (N_24913,N_24594,N_24749);
nor U24914 (N_24914,N_24674,N_24573);
xor U24915 (N_24915,N_24668,N_24701);
nand U24916 (N_24916,N_24622,N_24711);
xnor U24917 (N_24917,N_24627,N_24705);
nor U24918 (N_24918,N_24546,N_24720);
or U24919 (N_24919,N_24699,N_24567);
nand U24920 (N_24920,N_24592,N_24577);
and U24921 (N_24921,N_24681,N_24590);
or U24922 (N_24922,N_24501,N_24743);
nand U24923 (N_24923,N_24669,N_24579);
nand U24924 (N_24924,N_24523,N_24502);
nand U24925 (N_24925,N_24722,N_24636);
xor U24926 (N_24926,N_24554,N_24556);
nand U24927 (N_24927,N_24613,N_24598);
and U24928 (N_24928,N_24674,N_24584);
and U24929 (N_24929,N_24655,N_24702);
or U24930 (N_24930,N_24593,N_24566);
xnor U24931 (N_24931,N_24518,N_24741);
nor U24932 (N_24932,N_24586,N_24650);
nand U24933 (N_24933,N_24604,N_24615);
and U24934 (N_24934,N_24571,N_24526);
or U24935 (N_24935,N_24557,N_24671);
xor U24936 (N_24936,N_24571,N_24537);
or U24937 (N_24937,N_24660,N_24501);
or U24938 (N_24938,N_24731,N_24663);
or U24939 (N_24939,N_24545,N_24626);
and U24940 (N_24940,N_24681,N_24742);
nor U24941 (N_24941,N_24681,N_24595);
xnor U24942 (N_24942,N_24534,N_24724);
and U24943 (N_24943,N_24738,N_24663);
or U24944 (N_24944,N_24568,N_24672);
nor U24945 (N_24945,N_24598,N_24540);
nor U24946 (N_24946,N_24519,N_24725);
nor U24947 (N_24947,N_24683,N_24719);
nor U24948 (N_24948,N_24735,N_24561);
nor U24949 (N_24949,N_24572,N_24573);
and U24950 (N_24950,N_24501,N_24561);
or U24951 (N_24951,N_24629,N_24748);
nand U24952 (N_24952,N_24501,N_24723);
xnor U24953 (N_24953,N_24691,N_24688);
or U24954 (N_24954,N_24718,N_24710);
nand U24955 (N_24955,N_24693,N_24638);
nand U24956 (N_24956,N_24516,N_24740);
xnor U24957 (N_24957,N_24555,N_24536);
xnor U24958 (N_24958,N_24746,N_24636);
and U24959 (N_24959,N_24716,N_24572);
or U24960 (N_24960,N_24630,N_24557);
and U24961 (N_24961,N_24549,N_24611);
or U24962 (N_24962,N_24690,N_24692);
and U24963 (N_24963,N_24629,N_24560);
nand U24964 (N_24964,N_24635,N_24691);
xor U24965 (N_24965,N_24601,N_24721);
and U24966 (N_24966,N_24505,N_24596);
nand U24967 (N_24967,N_24670,N_24729);
and U24968 (N_24968,N_24672,N_24536);
nand U24969 (N_24969,N_24577,N_24594);
xor U24970 (N_24970,N_24644,N_24555);
nand U24971 (N_24971,N_24502,N_24700);
xor U24972 (N_24972,N_24720,N_24664);
or U24973 (N_24973,N_24557,N_24704);
or U24974 (N_24974,N_24735,N_24647);
or U24975 (N_24975,N_24578,N_24620);
xor U24976 (N_24976,N_24640,N_24736);
xor U24977 (N_24977,N_24648,N_24546);
nand U24978 (N_24978,N_24713,N_24585);
nor U24979 (N_24979,N_24501,N_24711);
and U24980 (N_24980,N_24715,N_24592);
nand U24981 (N_24981,N_24711,N_24667);
or U24982 (N_24982,N_24583,N_24518);
and U24983 (N_24983,N_24562,N_24662);
nor U24984 (N_24984,N_24529,N_24745);
nor U24985 (N_24985,N_24671,N_24693);
and U24986 (N_24986,N_24726,N_24571);
nor U24987 (N_24987,N_24690,N_24688);
nand U24988 (N_24988,N_24649,N_24683);
nor U24989 (N_24989,N_24516,N_24619);
and U24990 (N_24990,N_24600,N_24644);
or U24991 (N_24991,N_24532,N_24719);
nand U24992 (N_24992,N_24550,N_24583);
xnor U24993 (N_24993,N_24703,N_24673);
xor U24994 (N_24994,N_24690,N_24705);
or U24995 (N_24995,N_24568,N_24697);
xor U24996 (N_24996,N_24689,N_24742);
xor U24997 (N_24997,N_24743,N_24701);
nor U24998 (N_24998,N_24644,N_24511);
nor U24999 (N_24999,N_24675,N_24652);
or UO_0 (O_0,N_24991,N_24764);
and UO_1 (O_1,N_24880,N_24860);
xor UO_2 (O_2,N_24870,N_24781);
nor UO_3 (O_3,N_24858,N_24840);
or UO_4 (O_4,N_24789,N_24893);
nand UO_5 (O_5,N_24927,N_24946);
and UO_6 (O_6,N_24957,N_24850);
or UO_7 (O_7,N_24940,N_24819);
nand UO_8 (O_8,N_24836,N_24871);
nor UO_9 (O_9,N_24924,N_24908);
and UO_10 (O_10,N_24759,N_24841);
xor UO_11 (O_11,N_24766,N_24797);
or UO_12 (O_12,N_24967,N_24996);
or UO_13 (O_13,N_24867,N_24821);
or UO_14 (O_14,N_24817,N_24943);
nor UO_15 (O_15,N_24892,N_24997);
nor UO_16 (O_16,N_24888,N_24909);
nand UO_17 (O_17,N_24823,N_24798);
or UO_18 (O_18,N_24779,N_24906);
nor UO_19 (O_19,N_24780,N_24785);
xnor UO_20 (O_20,N_24810,N_24921);
nand UO_21 (O_21,N_24869,N_24885);
and UO_22 (O_22,N_24993,N_24975);
or UO_23 (O_23,N_24775,N_24942);
nand UO_24 (O_24,N_24983,N_24790);
nand UO_25 (O_25,N_24904,N_24769);
nor UO_26 (O_26,N_24808,N_24941);
nand UO_27 (O_27,N_24799,N_24831);
nand UO_28 (O_28,N_24986,N_24917);
nor UO_29 (O_29,N_24838,N_24879);
xnor UO_30 (O_30,N_24820,N_24796);
and UO_31 (O_31,N_24762,N_24757);
and UO_32 (O_32,N_24899,N_24752);
nor UO_33 (O_33,N_24777,N_24883);
nor UO_34 (O_34,N_24771,N_24911);
nand UO_35 (O_35,N_24786,N_24890);
nand UO_36 (O_36,N_24832,N_24852);
nand UO_37 (O_37,N_24963,N_24964);
or UO_38 (O_38,N_24998,N_24804);
nor UO_39 (O_39,N_24788,N_24994);
nor UO_40 (O_40,N_24966,N_24970);
nand UO_41 (O_41,N_24876,N_24928);
or UO_42 (O_42,N_24894,N_24981);
nand UO_43 (O_43,N_24952,N_24811);
nor UO_44 (O_44,N_24837,N_24969);
nand UO_45 (O_45,N_24767,N_24770);
and UO_46 (O_46,N_24953,N_24873);
nor UO_47 (O_47,N_24972,N_24945);
and UO_48 (O_48,N_24816,N_24829);
nand UO_49 (O_49,N_24968,N_24980);
or UO_50 (O_50,N_24863,N_24987);
or UO_51 (O_51,N_24750,N_24918);
xnor UO_52 (O_52,N_24973,N_24874);
and UO_53 (O_53,N_24793,N_24910);
nor UO_54 (O_54,N_24857,N_24897);
or UO_55 (O_55,N_24854,N_24926);
nor UO_56 (O_56,N_24791,N_24826);
or UO_57 (O_57,N_24795,N_24809);
nand UO_58 (O_58,N_24828,N_24824);
and UO_59 (O_59,N_24903,N_24955);
nand UO_60 (O_60,N_24847,N_24774);
and UO_61 (O_61,N_24822,N_24988);
nor UO_62 (O_62,N_24751,N_24979);
or UO_63 (O_63,N_24835,N_24976);
xor UO_64 (O_64,N_24803,N_24959);
xnor UO_65 (O_65,N_24982,N_24882);
xnor UO_66 (O_66,N_24755,N_24827);
or UO_67 (O_67,N_24891,N_24920);
nand UO_68 (O_68,N_24855,N_24784);
nor UO_69 (O_69,N_24872,N_24801);
nor UO_70 (O_70,N_24938,N_24949);
xnor UO_71 (O_71,N_24778,N_24758);
and UO_72 (O_72,N_24990,N_24802);
xor UO_73 (O_73,N_24901,N_24765);
nand UO_74 (O_74,N_24815,N_24846);
xnor UO_75 (O_75,N_24776,N_24935);
or UO_76 (O_76,N_24944,N_24977);
nor UO_77 (O_77,N_24830,N_24761);
nor UO_78 (O_78,N_24754,N_24962);
nand UO_79 (O_79,N_24884,N_24922);
nand UO_80 (O_80,N_24834,N_24999);
or UO_81 (O_81,N_24805,N_24851);
or UO_82 (O_82,N_24807,N_24881);
and UO_83 (O_83,N_24933,N_24868);
nor UO_84 (O_84,N_24814,N_24954);
xor UO_85 (O_85,N_24813,N_24848);
or UO_86 (O_86,N_24773,N_24947);
nor UO_87 (O_87,N_24974,N_24960);
or UO_88 (O_88,N_24756,N_24956);
xnor UO_89 (O_89,N_24958,N_24948);
xnor UO_90 (O_90,N_24875,N_24812);
nand UO_91 (O_91,N_24862,N_24915);
or UO_92 (O_92,N_24985,N_24900);
nand UO_93 (O_93,N_24833,N_24889);
nor UO_94 (O_94,N_24806,N_24772);
nand UO_95 (O_95,N_24753,N_24886);
nand UO_96 (O_96,N_24787,N_24929);
xnor UO_97 (O_97,N_24923,N_24853);
and UO_98 (O_98,N_24989,N_24961);
and UO_99 (O_99,N_24800,N_24768);
or UO_100 (O_100,N_24849,N_24783);
xor UO_101 (O_101,N_24913,N_24782);
nor UO_102 (O_102,N_24825,N_24984);
nand UO_103 (O_103,N_24843,N_24877);
or UO_104 (O_104,N_24878,N_24794);
xnor UO_105 (O_105,N_24939,N_24895);
or UO_106 (O_106,N_24950,N_24931);
or UO_107 (O_107,N_24914,N_24919);
nand UO_108 (O_108,N_24844,N_24763);
or UO_109 (O_109,N_24861,N_24845);
nor UO_110 (O_110,N_24760,N_24818);
and UO_111 (O_111,N_24792,N_24839);
and UO_112 (O_112,N_24916,N_24905);
and UO_113 (O_113,N_24856,N_24907);
nand UO_114 (O_114,N_24912,N_24902);
nand UO_115 (O_115,N_24934,N_24896);
nand UO_116 (O_116,N_24859,N_24992);
xor UO_117 (O_117,N_24887,N_24930);
or UO_118 (O_118,N_24937,N_24936);
nand UO_119 (O_119,N_24864,N_24925);
nor UO_120 (O_120,N_24971,N_24842);
or UO_121 (O_121,N_24866,N_24898);
or UO_122 (O_122,N_24978,N_24965);
xor UO_123 (O_123,N_24951,N_24865);
or UO_124 (O_124,N_24995,N_24932);
nand UO_125 (O_125,N_24821,N_24761);
nor UO_126 (O_126,N_24873,N_24997);
nand UO_127 (O_127,N_24847,N_24891);
and UO_128 (O_128,N_24996,N_24775);
nor UO_129 (O_129,N_24812,N_24791);
nor UO_130 (O_130,N_24977,N_24960);
and UO_131 (O_131,N_24904,N_24775);
nor UO_132 (O_132,N_24969,N_24860);
nor UO_133 (O_133,N_24898,N_24948);
and UO_134 (O_134,N_24852,N_24785);
or UO_135 (O_135,N_24762,N_24826);
or UO_136 (O_136,N_24887,N_24845);
nand UO_137 (O_137,N_24762,N_24973);
or UO_138 (O_138,N_24817,N_24868);
and UO_139 (O_139,N_24906,N_24913);
or UO_140 (O_140,N_24891,N_24751);
xnor UO_141 (O_141,N_24874,N_24832);
xor UO_142 (O_142,N_24962,N_24770);
or UO_143 (O_143,N_24815,N_24989);
nor UO_144 (O_144,N_24901,N_24966);
or UO_145 (O_145,N_24818,N_24889);
nand UO_146 (O_146,N_24823,N_24994);
or UO_147 (O_147,N_24858,N_24989);
or UO_148 (O_148,N_24880,N_24891);
nor UO_149 (O_149,N_24936,N_24852);
or UO_150 (O_150,N_24992,N_24952);
or UO_151 (O_151,N_24846,N_24893);
or UO_152 (O_152,N_24807,N_24759);
and UO_153 (O_153,N_24882,N_24751);
or UO_154 (O_154,N_24830,N_24993);
and UO_155 (O_155,N_24868,N_24946);
or UO_156 (O_156,N_24765,N_24891);
and UO_157 (O_157,N_24971,N_24805);
nor UO_158 (O_158,N_24950,N_24842);
and UO_159 (O_159,N_24845,N_24891);
nor UO_160 (O_160,N_24775,N_24750);
nor UO_161 (O_161,N_24899,N_24768);
nand UO_162 (O_162,N_24963,N_24810);
nand UO_163 (O_163,N_24879,N_24954);
and UO_164 (O_164,N_24827,N_24936);
xnor UO_165 (O_165,N_24776,N_24817);
and UO_166 (O_166,N_24842,N_24955);
nor UO_167 (O_167,N_24911,N_24997);
and UO_168 (O_168,N_24976,N_24796);
nand UO_169 (O_169,N_24994,N_24842);
nand UO_170 (O_170,N_24756,N_24761);
or UO_171 (O_171,N_24850,N_24768);
xnor UO_172 (O_172,N_24903,N_24966);
nand UO_173 (O_173,N_24920,N_24881);
nand UO_174 (O_174,N_24884,N_24833);
nand UO_175 (O_175,N_24842,N_24848);
nor UO_176 (O_176,N_24977,N_24825);
xnor UO_177 (O_177,N_24777,N_24830);
nor UO_178 (O_178,N_24993,N_24976);
and UO_179 (O_179,N_24769,N_24955);
nor UO_180 (O_180,N_24976,N_24766);
and UO_181 (O_181,N_24950,N_24947);
or UO_182 (O_182,N_24791,N_24981);
xor UO_183 (O_183,N_24854,N_24778);
or UO_184 (O_184,N_24935,N_24950);
xor UO_185 (O_185,N_24811,N_24992);
or UO_186 (O_186,N_24958,N_24985);
or UO_187 (O_187,N_24752,N_24814);
and UO_188 (O_188,N_24984,N_24888);
or UO_189 (O_189,N_24965,N_24866);
nor UO_190 (O_190,N_24803,N_24971);
xor UO_191 (O_191,N_24904,N_24984);
nor UO_192 (O_192,N_24868,N_24911);
xor UO_193 (O_193,N_24821,N_24936);
xor UO_194 (O_194,N_24863,N_24765);
or UO_195 (O_195,N_24901,N_24830);
nand UO_196 (O_196,N_24895,N_24830);
xor UO_197 (O_197,N_24800,N_24750);
and UO_198 (O_198,N_24900,N_24793);
nand UO_199 (O_199,N_24847,N_24940);
xor UO_200 (O_200,N_24868,N_24919);
xor UO_201 (O_201,N_24750,N_24752);
nand UO_202 (O_202,N_24948,N_24927);
xor UO_203 (O_203,N_24873,N_24937);
and UO_204 (O_204,N_24885,N_24909);
nor UO_205 (O_205,N_24968,N_24778);
nor UO_206 (O_206,N_24852,N_24904);
nand UO_207 (O_207,N_24788,N_24843);
nand UO_208 (O_208,N_24876,N_24967);
xor UO_209 (O_209,N_24904,N_24960);
or UO_210 (O_210,N_24891,N_24938);
or UO_211 (O_211,N_24906,N_24851);
xnor UO_212 (O_212,N_24932,N_24765);
and UO_213 (O_213,N_24778,N_24959);
nor UO_214 (O_214,N_24791,N_24811);
nor UO_215 (O_215,N_24916,N_24789);
or UO_216 (O_216,N_24888,N_24849);
and UO_217 (O_217,N_24860,N_24864);
nor UO_218 (O_218,N_24853,N_24871);
xnor UO_219 (O_219,N_24793,N_24938);
xnor UO_220 (O_220,N_24801,N_24930);
nor UO_221 (O_221,N_24769,N_24902);
nor UO_222 (O_222,N_24864,N_24872);
and UO_223 (O_223,N_24953,N_24932);
nand UO_224 (O_224,N_24856,N_24853);
nand UO_225 (O_225,N_24941,N_24817);
or UO_226 (O_226,N_24940,N_24906);
and UO_227 (O_227,N_24806,N_24779);
nand UO_228 (O_228,N_24994,N_24833);
nor UO_229 (O_229,N_24943,N_24784);
xnor UO_230 (O_230,N_24820,N_24927);
nor UO_231 (O_231,N_24860,N_24899);
and UO_232 (O_232,N_24878,N_24968);
nor UO_233 (O_233,N_24995,N_24788);
nand UO_234 (O_234,N_24811,N_24817);
nor UO_235 (O_235,N_24969,N_24864);
nand UO_236 (O_236,N_24833,N_24752);
nor UO_237 (O_237,N_24985,N_24974);
nor UO_238 (O_238,N_24918,N_24796);
nor UO_239 (O_239,N_24945,N_24999);
xnor UO_240 (O_240,N_24853,N_24873);
nor UO_241 (O_241,N_24787,N_24801);
or UO_242 (O_242,N_24786,N_24828);
and UO_243 (O_243,N_24896,N_24995);
nor UO_244 (O_244,N_24873,N_24839);
and UO_245 (O_245,N_24777,N_24762);
nor UO_246 (O_246,N_24814,N_24777);
xnor UO_247 (O_247,N_24839,N_24925);
xnor UO_248 (O_248,N_24968,N_24897);
and UO_249 (O_249,N_24926,N_24966);
nand UO_250 (O_250,N_24941,N_24958);
and UO_251 (O_251,N_24860,N_24872);
xor UO_252 (O_252,N_24759,N_24870);
or UO_253 (O_253,N_24916,N_24906);
nor UO_254 (O_254,N_24923,N_24991);
or UO_255 (O_255,N_24938,N_24785);
and UO_256 (O_256,N_24894,N_24807);
or UO_257 (O_257,N_24754,N_24793);
xnor UO_258 (O_258,N_24913,N_24890);
xor UO_259 (O_259,N_24894,N_24814);
nand UO_260 (O_260,N_24918,N_24757);
nand UO_261 (O_261,N_24976,N_24983);
nand UO_262 (O_262,N_24765,N_24981);
nor UO_263 (O_263,N_24847,N_24980);
nand UO_264 (O_264,N_24954,N_24788);
and UO_265 (O_265,N_24937,N_24855);
nor UO_266 (O_266,N_24781,N_24913);
nor UO_267 (O_267,N_24754,N_24988);
or UO_268 (O_268,N_24825,N_24998);
nand UO_269 (O_269,N_24823,N_24921);
and UO_270 (O_270,N_24887,N_24851);
nand UO_271 (O_271,N_24810,N_24809);
nand UO_272 (O_272,N_24890,N_24880);
and UO_273 (O_273,N_24762,N_24983);
xnor UO_274 (O_274,N_24906,N_24862);
nand UO_275 (O_275,N_24885,N_24894);
or UO_276 (O_276,N_24781,N_24874);
xor UO_277 (O_277,N_24782,N_24880);
and UO_278 (O_278,N_24932,N_24825);
or UO_279 (O_279,N_24817,N_24887);
xnor UO_280 (O_280,N_24918,N_24883);
xor UO_281 (O_281,N_24914,N_24938);
and UO_282 (O_282,N_24896,N_24925);
xor UO_283 (O_283,N_24985,N_24970);
or UO_284 (O_284,N_24845,N_24968);
nor UO_285 (O_285,N_24935,N_24856);
nor UO_286 (O_286,N_24879,N_24782);
xnor UO_287 (O_287,N_24874,N_24856);
nand UO_288 (O_288,N_24797,N_24948);
nand UO_289 (O_289,N_24894,N_24750);
nor UO_290 (O_290,N_24781,N_24871);
nor UO_291 (O_291,N_24934,N_24944);
or UO_292 (O_292,N_24976,N_24786);
nand UO_293 (O_293,N_24900,N_24938);
xnor UO_294 (O_294,N_24905,N_24759);
nor UO_295 (O_295,N_24903,N_24921);
or UO_296 (O_296,N_24780,N_24996);
nor UO_297 (O_297,N_24842,N_24875);
xnor UO_298 (O_298,N_24922,N_24814);
nand UO_299 (O_299,N_24785,N_24814);
or UO_300 (O_300,N_24900,N_24894);
or UO_301 (O_301,N_24846,N_24940);
xor UO_302 (O_302,N_24968,N_24798);
nand UO_303 (O_303,N_24764,N_24920);
nand UO_304 (O_304,N_24915,N_24922);
xnor UO_305 (O_305,N_24985,N_24819);
or UO_306 (O_306,N_24843,N_24762);
nor UO_307 (O_307,N_24770,N_24889);
and UO_308 (O_308,N_24759,N_24874);
or UO_309 (O_309,N_24794,N_24975);
nand UO_310 (O_310,N_24930,N_24868);
or UO_311 (O_311,N_24919,N_24788);
or UO_312 (O_312,N_24936,N_24920);
xnor UO_313 (O_313,N_24948,N_24955);
nor UO_314 (O_314,N_24916,N_24802);
nand UO_315 (O_315,N_24933,N_24896);
and UO_316 (O_316,N_24785,N_24804);
xnor UO_317 (O_317,N_24967,N_24837);
or UO_318 (O_318,N_24874,N_24938);
and UO_319 (O_319,N_24996,N_24979);
or UO_320 (O_320,N_24956,N_24844);
nor UO_321 (O_321,N_24968,N_24805);
nor UO_322 (O_322,N_24894,N_24761);
or UO_323 (O_323,N_24780,N_24957);
and UO_324 (O_324,N_24978,N_24932);
nor UO_325 (O_325,N_24893,N_24875);
and UO_326 (O_326,N_24755,N_24909);
or UO_327 (O_327,N_24833,N_24841);
and UO_328 (O_328,N_24949,N_24995);
and UO_329 (O_329,N_24754,N_24800);
and UO_330 (O_330,N_24763,N_24961);
or UO_331 (O_331,N_24773,N_24910);
nor UO_332 (O_332,N_24897,N_24759);
xnor UO_333 (O_333,N_24914,N_24974);
and UO_334 (O_334,N_24772,N_24863);
or UO_335 (O_335,N_24954,N_24844);
nand UO_336 (O_336,N_24857,N_24761);
nor UO_337 (O_337,N_24905,N_24937);
or UO_338 (O_338,N_24832,N_24922);
nand UO_339 (O_339,N_24834,N_24801);
xnor UO_340 (O_340,N_24779,N_24853);
or UO_341 (O_341,N_24984,N_24956);
or UO_342 (O_342,N_24923,N_24932);
xnor UO_343 (O_343,N_24925,N_24760);
and UO_344 (O_344,N_24825,N_24902);
nand UO_345 (O_345,N_24765,N_24971);
or UO_346 (O_346,N_24825,N_24909);
nand UO_347 (O_347,N_24933,N_24842);
nand UO_348 (O_348,N_24941,N_24810);
and UO_349 (O_349,N_24927,N_24897);
xnor UO_350 (O_350,N_24816,N_24782);
and UO_351 (O_351,N_24984,N_24808);
or UO_352 (O_352,N_24922,N_24752);
nand UO_353 (O_353,N_24797,N_24871);
or UO_354 (O_354,N_24777,N_24973);
nand UO_355 (O_355,N_24861,N_24924);
and UO_356 (O_356,N_24890,N_24886);
or UO_357 (O_357,N_24752,N_24904);
xnor UO_358 (O_358,N_24973,N_24781);
or UO_359 (O_359,N_24893,N_24773);
nand UO_360 (O_360,N_24829,N_24981);
xor UO_361 (O_361,N_24883,N_24780);
xnor UO_362 (O_362,N_24934,N_24830);
nor UO_363 (O_363,N_24907,N_24963);
and UO_364 (O_364,N_24864,N_24826);
nor UO_365 (O_365,N_24906,N_24945);
nor UO_366 (O_366,N_24752,N_24825);
nand UO_367 (O_367,N_24773,N_24852);
nand UO_368 (O_368,N_24864,N_24970);
xnor UO_369 (O_369,N_24866,N_24928);
or UO_370 (O_370,N_24802,N_24978);
and UO_371 (O_371,N_24779,N_24902);
nor UO_372 (O_372,N_24797,N_24954);
and UO_373 (O_373,N_24982,N_24935);
nand UO_374 (O_374,N_24993,N_24832);
and UO_375 (O_375,N_24766,N_24868);
and UO_376 (O_376,N_24950,N_24886);
and UO_377 (O_377,N_24762,N_24756);
nand UO_378 (O_378,N_24927,N_24958);
nand UO_379 (O_379,N_24967,N_24893);
nor UO_380 (O_380,N_24995,N_24960);
and UO_381 (O_381,N_24773,N_24837);
or UO_382 (O_382,N_24825,N_24764);
xor UO_383 (O_383,N_24926,N_24937);
and UO_384 (O_384,N_24945,N_24979);
xor UO_385 (O_385,N_24875,N_24943);
nor UO_386 (O_386,N_24891,N_24982);
xnor UO_387 (O_387,N_24981,N_24872);
nor UO_388 (O_388,N_24833,N_24914);
nand UO_389 (O_389,N_24981,N_24985);
nor UO_390 (O_390,N_24877,N_24905);
xor UO_391 (O_391,N_24933,N_24963);
nand UO_392 (O_392,N_24901,N_24775);
nand UO_393 (O_393,N_24922,N_24806);
and UO_394 (O_394,N_24940,N_24849);
or UO_395 (O_395,N_24951,N_24969);
nand UO_396 (O_396,N_24801,N_24961);
xor UO_397 (O_397,N_24882,N_24826);
or UO_398 (O_398,N_24957,N_24995);
nor UO_399 (O_399,N_24942,N_24845);
and UO_400 (O_400,N_24967,N_24878);
nand UO_401 (O_401,N_24837,N_24891);
or UO_402 (O_402,N_24897,N_24918);
and UO_403 (O_403,N_24898,N_24771);
or UO_404 (O_404,N_24908,N_24917);
and UO_405 (O_405,N_24854,N_24996);
and UO_406 (O_406,N_24880,N_24763);
nor UO_407 (O_407,N_24957,N_24779);
or UO_408 (O_408,N_24753,N_24870);
nand UO_409 (O_409,N_24808,N_24900);
and UO_410 (O_410,N_24831,N_24801);
or UO_411 (O_411,N_24868,N_24755);
xnor UO_412 (O_412,N_24813,N_24753);
or UO_413 (O_413,N_24822,N_24868);
nor UO_414 (O_414,N_24857,N_24997);
or UO_415 (O_415,N_24778,N_24779);
nand UO_416 (O_416,N_24784,N_24942);
nor UO_417 (O_417,N_24848,N_24883);
nand UO_418 (O_418,N_24849,N_24824);
or UO_419 (O_419,N_24912,N_24989);
nor UO_420 (O_420,N_24854,N_24809);
nor UO_421 (O_421,N_24877,N_24788);
nand UO_422 (O_422,N_24800,N_24942);
and UO_423 (O_423,N_24877,N_24847);
or UO_424 (O_424,N_24843,N_24771);
and UO_425 (O_425,N_24897,N_24871);
and UO_426 (O_426,N_24989,N_24916);
and UO_427 (O_427,N_24849,N_24789);
nor UO_428 (O_428,N_24966,N_24898);
xnor UO_429 (O_429,N_24843,N_24933);
and UO_430 (O_430,N_24934,N_24969);
or UO_431 (O_431,N_24951,N_24844);
nor UO_432 (O_432,N_24801,N_24861);
or UO_433 (O_433,N_24947,N_24820);
nand UO_434 (O_434,N_24804,N_24764);
nand UO_435 (O_435,N_24850,N_24929);
or UO_436 (O_436,N_24918,N_24923);
nand UO_437 (O_437,N_24786,N_24766);
or UO_438 (O_438,N_24969,N_24985);
and UO_439 (O_439,N_24892,N_24790);
nor UO_440 (O_440,N_24885,N_24902);
xnor UO_441 (O_441,N_24991,N_24783);
and UO_442 (O_442,N_24937,N_24983);
nor UO_443 (O_443,N_24979,N_24875);
xnor UO_444 (O_444,N_24923,N_24815);
nand UO_445 (O_445,N_24859,N_24988);
xor UO_446 (O_446,N_24947,N_24999);
and UO_447 (O_447,N_24755,N_24752);
xnor UO_448 (O_448,N_24935,N_24770);
or UO_449 (O_449,N_24806,N_24869);
xor UO_450 (O_450,N_24913,N_24900);
and UO_451 (O_451,N_24842,N_24830);
xor UO_452 (O_452,N_24750,N_24793);
nand UO_453 (O_453,N_24929,N_24789);
nor UO_454 (O_454,N_24872,N_24794);
or UO_455 (O_455,N_24868,N_24965);
nand UO_456 (O_456,N_24990,N_24888);
and UO_457 (O_457,N_24965,N_24835);
nand UO_458 (O_458,N_24784,N_24968);
xor UO_459 (O_459,N_24891,N_24852);
and UO_460 (O_460,N_24973,N_24818);
nor UO_461 (O_461,N_24932,N_24785);
or UO_462 (O_462,N_24923,N_24978);
xnor UO_463 (O_463,N_24803,N_24927);
and UO_464 (O_464,N_24874,N_24923);
nand UO_465 (O_465,N_24964,N_24867);
xnor UO_466 (O_466,N_24773,N_24830);
nand UO_467 (O_467,N_24755,N_24846);
or UO_468 (O_468,N_24911,N_24933);
or UO_469 (O_469,N_24987,N_24998);
nor UO_470 (O_470,N_24790,N_24768);
nand UO_471 (O_471,N_24927,N_24795);
nand UO_472 (O_472,N_24886,N_24940);
and UO_473 (O_473,N_24854,N_24823);
nor UO_474 (O_474,N_24843,N_24809);
and UO_475 (O_475,N_24777,N_24885);
nand UO_476 (O_476,N_24878,N_24915);
and UO_477 (O_477,N_24993,N_24824);
nand UO_478 (O_478,N_24786,N_24836);
nor UO_479 (O_479,N_24864,N_24898);
xor UO_480 (O_480,N_24926,N_24947);
nand UO_481 (O_481,N_24968,N_24961);
nand UO_482 (O_482,N_24804,N_24809);
xnor UO_483 (O_483,N_24940,N_24787);
xnor UO_484 (O_484,N_24935,N_24756);
and UO_485 (O_485,N_24761,N_24828);
and UO_486 (O_486,N_24970,N_24887);
or UO_487 (O_487,N_24897,N_24903);
or UO_488 (O_488,N_24841,N_24804);
nor UO_489 (O_489,N_24902,N_24998);
xnor UO_490 (O_490,N_24830,N_24956);
or UO_491 (O_491,N_24790,N_24834);
nand UO_492 (O_492,N_24904,N_24776);
nand UO_493 (O_493,N_24814,N_24800);
or UO_494 (O_494,N_24960,N_24907);
and UO_495 (O_495,N_24869,N_24940);
or UO_496 (O_496,N_24897,N_24889);
and UO_497 (O_497,N_24970,N_24854);
nor UO_498 (O_498,N_24966,N_24858);
and UO_499 (O_499,N_24834,N_24755);
nand UO_500 (O_500,N_24887,N_24973);
or UO_501 (O_501,N_24762,N_24910);
xnor UO_502 (O_502,N_24856,N_24839);
or UO_503 (O_503,N_24995,N_24968);
nor UO_504 (O_504,N_24878,N_24851);
nor UO_505 (O_505,N_24994,N_24794);
or UO_506 (O_506,N_24781,N_24861);
nor UO_507 (O_507,N_24966,N_24925);
nor UO_508 (O_508,N_24858,N_24784);
or UO_509 (O_509,N_24902,N_24792);
and UO_510 (O_510,N_24981,N_24835);
nor UO_511 (O_511,N_24752,N_24931);
and UO_512 (O_512,N_24832,N_24918);
and UO_513 (O_513,N_24948,N_24906);
nor UO_514 (O_514,N_24849,N_24970);
xor UO_515 (O_515,N_24925,N_24761);
and UO_516 (O_516,N_24945,N_24899);
or UO_517 (O_517,N_24761,N_24785);
or UO_518 (O_518,N_24781,N_24805);
nand UO_519 (O_519,N_24811,N_24913);
xor UO_520 (O_520,N_24962,N_24987);
and UO_521 (O_521,N_24853,N_24935);
nand UO_522 (O_522,N_24835,N_24810);
nand UO_523 (O_523,N_24927,N_24921);
and UO_524 (O_524,N_24857,N_24771);
nand UO_525 (O_525,N_24864,N_24873);
nand UO_526 (O_526,N_24827,N_24798);
or UO_527 (O_527,N_24988,N_24764);
or UO_528 (O_528,N_24828,N_24997);
xnor UO_529 (O_529,N_24761,N_24787);
nor UO_530 (O_530,N_24993,N_24764);
and UO_531 (O_531,N_24828,N_24879);
or UO_532 (O_532,N_24802,N_24786);
or UO_533 (O_533,N_24897,N_24785);
xor UO_534 (O_534,N_24904,N_24878);
nand UO_535 (O_535,N_24753,N_24817);
and UO_536 (O_536,N_24883,N_24923);
xor UO_537 (O_537,N_24946,N_24825);
xor UO_538 (O_538,N_24933,N_24886);
and UO_539 (O_539,N_24929,N_24958);
nand UO_540 (O_540,N_24908,N_24827);
or UO_541 (O_541,N_24998,N_24886);
nor UO_542 (O_542,N_24974,N_24825);
and UO_543 (O_543,N_24762,N_24808);
and UO_544 (O_544,N_24831,N_24764);
nor UO_545 (O_545,N_24772,N_24822);
nand UO_546 (O_546,N_24758,N_24841);
or UO_547 (O_547,N_24770,N_24976);
nand UO_548 (O_548,N_24870,N_24839);
nor UO_549 (O_549,N_24952,N_24841);
xor UO_550 (O_550,N_24769,N_24778);
xnor UO_551 (O_551,N_24764,N_24907);
nor UO_552 (O_552,N_24987,N_24919);
nand UO_553 (O_553,N_24770,N_24823);
nor UO_554 (O_554,N_24953,N_24833);
nor UO_555 (O_555,N_24951,N_24932);
nor UO_556 (O_556,N_24898,N_24897);
and UO_557 (O_557,N_24843,N_24863);
and UO_558 (O_558,N_24897,N_24986);
xnor UO_559 (O_559,N_24904,N_24798);
nand UO_560 (O_560,N_24932,N_24937);
xnor UO_561 (O_561,N_24757,N_24892);
and UO_562 (O_562,N_24869,N_24859);
and UO_563 (O_563,N_24781,N_24788);
xnor UO_564 (O_564,N_24751,N_24959);
xor UO_565 (O_565,N_24831,N_24984);
and UO_566 (O_566,N_24926,N_24794);
and UO_567 (O_567,N_24809,N_24911);
or UO_568 (O_568,N_24762,N_24953);
nor UO_569 (O_569,N_24805,N_24797);
nor UO_570 (O_570,N_24999,N_24953);
nand UO_571 (O_571,N_24995,N_24984);
xnor UO_572 (O_572,N_24878,N_24830);
and UO_573 (O_573,N_24941,N_24836);
xnor UO_574 (O_574,N_24955,N_24809);
nand UO_575 (O_575,N_24761,N_24904);
nand UO_576 (O_576,N_24818,N_24787);
nand UO_577 (O_577,N_24828,N_24969);
or UO_578 (O_578,N_24774,N_24965);
or UO_579 (O_579,N_24889,N_24844);
or UO_580 (O_580,N_24805,N_24867);
and UO_581 (O_581,N_24831,N_24872);
or UO_582 (O_582,N_24877,N_24925);
and UO_583 (O_583,N_24959,N_24805);
nor UO_584 (O_584,N_24975,N_24983);
xor UO_585 (O_585,N_24917,N_24975);
nand UO_586 (O_586,N_24961,N_24777);
or UO_587 (O_587,N_24943,N_24972);
and UO_588 (O_588,N_24837,N_24848);
nor UO_589 (O_589,N_24917,N_24832);
xor UO_590 (O_590,N_24879,N_24997);
nor UO_591 (O_591,N_24915,N_24777);
and UO_592 (O_592,N_24974,N_24761);
nand UO_593 (O_593,N_24950,N_24937);
xor UO_594 (O_594,N_24774,N_24840);
xor UO_595 (O_595,N_24969,N_24822);
xor UO_596 (O_596,N_24859,N_24998);
and UO_597 (O_597,N_24887,N_24868);
xnor UO_598 (O_598,N_24998,N_24979);
nand UO_599 (O_599,N_24792,N_24834);
and UO_600 (O_600,N_24898,N_24757);
nor UO_601 (O_601,N_24933,N_24917);
and UO_602 (O_602,N_24849,N_24973);
xnor UO_603 (O_603,N_24807,N_24814);
and UO_604 (O_604,N_24975,N_24856);
xor UO_605 (O_605,N_24851,N_24888);
and UO_606 (O_606,N_24832,N_24873);
nand UO_607 (O_607,N_24918,N_24880);
or UO_608 (O_608,N_24999,N_24836);
nor UO_609 (O_609,N_24803,N_24840);
or UO_610 (O_610,N_24829,N_24889);
nor UO_611 (O_611,N_24770,N_24988);
and UO_612 (O_612,N_24994,N_24930);
xnor UO_613 (O_613,N_24770,N_24787);
nand UO_614 (O_614,N_24958,N_24770);
xor UO_615 (O_615,N_24754,N_24948);
nor UO_616 (O_616,N_24848,N_24982);
and UO_617 (O_617,N_24824,N_24990);
xor UO_618 (O_618,N_24840,N_24863);
nor UO_619 (O_619,N_24994,N_24849);
xor UO_620 (O_620,N_24823,N_24785);
xnor UO_621 (O_621,N_24938,N_24980);
nand UO_622 (O_622,N_24863,N_24906);
xnor UO_623 (O_623,N_24904,N_24997);
and UO_624 (O_624,N_24785,N_24770);
nand UO_625 (O_625,N_24950,N_24943);
or UO_626 (O_626,N_24834,N_24774);
xor UO_627 (O_627,N_24825,N_24842);
nand UO_628 (O_628,N_24926,N_24915);
nor UO_629 (O_629,N_24998,N_24842);
nand UO_630 (O_630,N_24865,N_24883);
and UO_631 (O_631,N_24870,N_24790);
xnor UO_632 (O_632,N_24818,N_24965);
and UO_633 (O_633,N_24767,N_24901);
or UO_634 (O_634,N_24856,N_24828);
nand UO_635 (O_635,N_24870,N_24993);
nor UO_636 (O_636,N_24996,N_24953);
xor UO_637 (O_637,N_24816,N_24986);
and UO_638 (O_638,N_24783,N_24820);
nand UO_639 (O_639,N_24778,N_24751);
or UO_640 (O_640,N_24785,N_24765);
nor UO_641 (O_641,N_24923,N_24947);
and UO_642 (O_642,N_24871,N_24852);
nor UO_643 (O_643,N_24913,N_24891);
nand UO_644 (O_644,N_24806,N_24788);
nor UO_645 (O_645,N_24920,N_24996);
and UO_646 (O_646,N_24990,N_24952);
or UO_647 (O_647,N_24927,N_24836);
nor UO_648 (O_648,N_24870,N_24812);
nor UO_649 (O_649,N_24760,N_24830);
nand UO_650 (O_650,N_24754,N_24971);
xor UO_651 (O_651,N_24888,N_24893);
and UO_652 (O_652,N_24860,N_24901);
xnor UO_653 (O_653,N_24900,N_24762);
or UO_654 (O_654,N_24851,N_24849);
nor UO_655 (O_655,N_24766,N_24930);
or UO_656 (O_656,N_24754,N_24952);
and UO_657 (O_657,N_24790,N_24860);
nand UO_658 (O_658,N_24770,N_24870);
xor UO_659 (O_659,N_24932,N_24930);
nor UO_660 (O_660,N_24879,N_24836);
xnor UO_661 (O_661,N_24828,N_24854);
and UO_662 (O_662,N_24878,N_24922);
and UO_663 (O_663,N_24934,N_24915);
and UO_664 (O_664,N_24880,N_24935);
and UO_665 (O_665,N_24766,N_24893);
or UO_666 (O_666,N_24793,N_24885);
and UO_667 (O_667,N_24931,N_24912);
xor UO_668 (O_668,N_24864,N_24884);
and UO_669 (O_669,N_24884,N_24825);
xnor UO_670 (O_670,N_24921,N_24999);
or UO_671 (O_671,N_24962,N_24759);
nand UO_672 (O_672,N_24804,N_24780);
nor UO_673 (O_673,N_24832,N_24868);
nand UO_674 (O_674,N_24867,N_24837);
or UO_675 (O_675,N_24926,N_24858);
nand UO_676 (O_676,N_24986,N_24824);
nor UO_677 (O_677,N_24769,N_24848);
or UO_678 (O_678,N_24972,N_24792);
xor UO_679 (O_679,N_24953,N_24981);
xor UO_680 (O_680,N_24828,N_24762);
or UO_681 (O_681,N_24840,N_24833);
or UO_682 (O_682,N_24885,N_24836);
or UO_683 (O_683,N_24791,N_24914);
or UO_684 (O_684,N_24956,N_24853);
and UO_685 (O_685,N_24832,N_24856);
nor UO_686 (O_686,N_24959,N_24864);
or UO_687 (O_687,N_24905,N_24787);
nand UO_688 (O_688,N_24853,N_24917);
and UO_689 (O_689,N_24779,N_24889);
xor UO_690 (O_690,N_24839,N_24986);
or UO_691 (O_691,N_24880,N_24960);
nand UO_692 (O_692,N_24879,N_24858);
nand UO_693 (O_693,N_24753,N_24847);
nand UO_694 (O_694,N_24987,N_24797);
xnor UO_695 (O_695,N_24940,N_24979);
and UO_696 (O_696,N_24847,N_24913);
or UO_697 (O_697,N_24936,N_24832);
nand UO_698 (O_698,N_24888,N_24793);
or UO_699 (O_699,N_24859,N_24816);
nand UO_700 (O_700,N_24945,N_24909);
xnor UO_701 (O_701,N_24751,N_24964);
nand UO_702 (O_702,N_24916,N_24854);
xnor UO_703 (O_703,N_24997,N_24773);
or UO_704 (O_704,N_24801,N_24962);
xnor UO_705 (O_705,N_24951,N_24962);
nor UO_706 (O_706,N_24795,N_24923);
xnor UO_707 (O_707,N_24763,N_24901);
or UO_708 (O_708,N_24832,N_24862);
and UO_709 (O_709,N_24804,N_24985);
nand UO_710 (O_710,N_24844,N_24853);
nor UO_711 (O_711,N_24798,N_24885);
and UO_712 (O_712,N_24826,N_24902);
or UO_713 (O_713,N_24983,N_24799);
and UO_714 (O_714,N_24984,N_24920);
and UO_715 (O_715,N_24752,N_24819);
xnor UO_716 (O_716,N_24798,N_24787);
and UO_717 (O_717,N_24922,N_24917);
xnor UO_718 (O_718,N_24773,N_24783);
and UO_719 (O_719,N_24777,N_24838);
nand UO_720 (O_720,N_24759,N_24974);
xor UO_721 (O_721,N_24860,N_24842);
xnor UO_722 (O_722,N_24941,N_24940);
and UO_723 (O_723,N_24891,N_24860);
xor UO_724 (O_724,N_24887,N_24804);
nor UO_725 (O_725,N_24994,N_24821);
and UO_726 (O_726,N_24946,N_24866);
xor UO_727 (O_727,N_24994,N_24811);
and UO_728 (O_728,N_24896,N_24993);
xor UO_729 (O_729,N_24916,N_24998);
xor UO_730 (O_730,N_24952,N_24771);
or UO_731 (O_731,N_24942,N_24987);
xnor UO_732 (O_732,N_24843,N_24805);
nor UO_733 (O_733,N_24820,N_24760);
xnor UO_734 (O_734,N_24941,N_24912);
nand UO_735 (O_735,N_24950,N_24844);
nand UO_736 (O_736,N_24931,N_24923);
nand UO_737 (O_737,N_24928,N_24953);
and UO_738 (O_738,N_24918,N_24855);
or UO_739 (O_739,N_24833,N_24831);
nand UO_740 (O_740,N_24902,N_24849);
or UO_741 (O_741,N_24897,N_24977);
xnor UO_742 (O_742,N_24771,N_24801);
xor UO_743 (O_743,N_24869,N_24840);
xnor UO_744 (O_744,N_24910,N_24997);
or UO_745 (O_745,N_24834,N_24933);
nand UO_746 (O_746,N_24784,N_24893);
nor UO_747 (O_747,N_24904,N_24793);
xor UO_748 (O_748,N_24998,N_24969);
or UO_749 (O_749,N_24930,N_24863);
xor UO_750 (O_750,N_24865,N_24848);
nor UO_751 (O_751,N_24919,N_24915);
nor UO_752 (O_752,N_24947,N_24827);
nand UO_753 (O_753,N_24771,N_24909);
or UO_754 (O_754,N_24803,N_24824);
nand UO_755 (O_755,N_24867,N_24751);
or UO_756 (O_756,N_24803,N_24950);
xnor UO_757 (O_757,N_24817,N_24815);
or UO_758 (O_758,N_24867,N_24760);
xnor UO_759 (O_759,N_24866,N_24907);
nand UO_760 (O_760,N_24993,N_24866);
xnor UO_761 (O_761,N_24977,N_24831);
and UO_762 (O_762,N_24985,N_24815);
nand UO_763 (O_763,N_24798,N_24760);
xnor UO_764 (O_764,N_24788,N_24929);
nand UO_765 (O_765,N_24829,N_24901);
or UO_766 (O_766,N_24851,N_24903);
nand UO_767 (O_767,N_24785,N_24917);
or UO_768 (O_768,N_24791,N_24762);
xor UO_769 (O_769,N_24890,N_24891);
xnor UO_770 (O_770,N_24778,N_24966);
nor UO_771 (O_771,N_24878,N_24770);
nor UO_772 (O_772,N_24804,N_24939);
nand UO_773 (O_773,N_24978,N_24891);
and UO_774 (O_774,N_24849,N_24758);
and UO_775 (O_775,N_24870,N_24913);
xor UO_776 (O_776,N_24807,N_24933);
and UO_777 (O_777,N_24888,N_24936);
nand UO_778 (O_778,N_24946,N_24962);
xnor UO_779 (O_779,N_24855,N_24853);
nor UO_780 (O_780,N_24959,N_24995);
or UO_781 (O_781,N_24915,N_24771);
xor UO_782 (O_782,N_24981,N_24768);
nor UO_783 (O_783,N_24929,N_24918);
nor UO_784 (O_784,N_24991,N_24957);
and UO_785 (O_785,N_24803,N_24967);
and UO_786 (O_786,N_24868,N_24750);
xor UO_787 (O_787,N_24843,N_24810);
nor UO_788 (O_788,N_24870,N_24806);
nand UO_789 (O_789,N_24872,N_24752);
or UO_790 (O_790,N_24881,N_24850);
or UO_791 (O_791,N_24831,N_24815);
nand UO_792 (O_792,N_24878,N_24862);
nand UO_793 (O_793,N_24974,N_24943);
nand UO_794 (O_794,N_24937,N_24788);
or UO_795 (O_795,N_24759,N_24871);
nor UO_796 (O_796,N_24789,N_24976);
or UO_797 (O_797,N_24995,N_24847);
xor UO_798 (O_798,N_24856,N_24909);
xnor UO_799 (O_799,N_24854,N_24909);
or UO_800 (O_800,N_24755,N_24751);
nor UO_801 (O_801,N_24816,N_24791);
and UO_802 (O_802,N_24846,N_24955);
or UO_803 (O_803,N_24836,N_24757);
xor UO_804 (O_804,N_24850,N_24781);
nand UO_805 (O_805,N_24964,N_24930);
or UO_806 (O_806,N_24976,N_24928);
nor UO_807 (O_807,N_24919,N_24772);
and UO_808 (O_808,N_24785,N_24799);
nor UO_809 (O_809,N_24961,N_24950);
xnor UO_810 (O_810,N_24753,N_24937);
nor UO_811 (O_811,N_24901,N_24802);
nor UO_812 (O_812,N_24871,N_24867);
nand UO_813 (O_813,N_24957,N_24775);
nor UO_814 (O_814,N_24904,N_24865);
nor UO_815 (O_815,N_24867,N_24998);
and UO_816 (O_816,N_24969,N_24859);
nor UO_817 (O_817,N_24782,N_24997);
nand UO_818 (O_818,N_24921,N_24995);
or UO_819 (O_819,N_24803,N_24790);
and UO_820 (O_820,N_24786,N_24850);
and UO_821 (O_821,N_24880,N_24954);
nor UO_822 (O_822,N_24845,N_24874);
and UO_823 (O_823,N_24838,N_24875);
xor UO_824 (O_824,N_24792,N_24955);
or UO_825 (O_825,N_24907,N_24772);
and UO_826 (O_826,N_24920,N_24834);
xor UO_827 (O_827,N_24973,N_24907);
or UO_828 (O_828,N_24851,N_24943);
and UO_829 (O_829,N_24754,N_24978);
xnor UO_830 (O_830,N_24922,N_24950);
nor UO_831 (O_831,N_24795,N_24853);
and UO_832 (O_832,N_24821,N_24860);
nand UO_833 (O_833,N_24971,N_24872);
nand UO_834 (O_834,N_24904,N_24760);
nor UO_835 (O_835,N_24872,N_24803);
nor UO_836 (O_836,N_24753,N_24811);
or UO_837 (O_837,N_24884,N_24915);
or UO_838 (O_838,N_24873,N_24787);
or UO_839 (O_839,N_24784,N_24925);
nor UO_840 (O_840,N_24982,N_24986);
and UO_841 (O_841,N_24753,N_24810);
and UO_842 (O_842,N_24995,N_24766);
or UO_843 (O_843,N_24806,N_24758);
or UO_844 (O_844,N_24815,N_24873);
nand UO_845 (O_845,N_24814,N_24804);
and UO_846 (O_846,N_24763,N_24847);
xor UO_847 (O_847,N_24757,N_24990);
nor UO_848 (O_848,N_24892,N_24928);
nand UO_849 (O_849,N_24949,N_24803);
or UO_850 (O_850,N_24895,N_24917);
and UO_851 (O_851,N_24780,N_24903);
or UO_852 (O_852,N_24903,N_24870);
nand UO_853 (O_853,N_24765,N_24846);
xor UO_854 (O_854,N_24862,N_24998);
xnor UO_855 (O_855,N_24784,N_24769);
nand UO_856 (O_856,N_24948,N_24990);
or UO_857 (O_857,N_24989,N_24801);
nor UO_858 (O_858,N_24869,N_24947);
nand UO_859 (O_859,N_24948,N_24976);
or UO_860 (O_860,N_24779,N_24820);
or UO_861 (O_861,N_24931,N_24859);
xor UO_862 (O_862,N_24761,N_24900);
nand UO_863 (O_863,N_24769,N_24858);
and UO_864 (O_864,N_24798,N_24877);
nand UO_865 (O_865,N_24758,N_24903);
and UO_866 (O_866,N_24890,N_24923);
nor UO_867 (O_867,N_24850,N_24842);
nor UO_868 (O_868,N_24954,N_24972);
nor UO_869 (O_869,N_24773,N_24966);
nand UO_870 (O_870,N_24911,N_24950);
or UO_871 (O_871,N_24934,N_24981);
xor UO_872 (O_872,N_24864,N_24944);
or UO_873 (O_873,N_24765,N_24967);
nor UO_874 (O_874,N_24844,N_24972);
xnor UO_875 (O_875,N_24846,N_24896);
nand UO_876 (O_876,N_24856,N_24952);
xor UO_877 (O_877,N_24767,N_24992);
nand UO_878 (O_878,N_24959,N_24845);
nand UO_879 (O_879,N_24994,N_24790);
or UO_880 (O_880,N_24901,N_24883);
and UO_881 (O_881,N_24891,N_24940);
and UO_882 (O_882,N_24882,N_24884);
nor UO_883 (O_883,N_24769,N_24833);
xnor UO_884 (O_884,N_24784,N_24924);
nor UO_885 (O_885,N_24854,N_24984);
nor UO_886 (O_886,N_24917,N_24935);
xnor UO_887 (O_887,N_24753,N_24798);
nand UO_888 (O_888,N_24837,N_24760);
nand UO_889 (O_889,N_24997,N_24962);
xnor UO_890 (O_890,N_24890,N_24976);
and UO_891 (O_891,N_24766,N_24987);
nor UO_892 (O_892,N_24839,N_24806);
and UO_893 (O_893,N_24848,N_24853);
nor UO_894 (O_894,N_24798,N_24952);
or UO_895 (O_895,N_24837,N_24790);
and UO_896 (O_896,N_24859,N_24759);
or UO_897 (O_897,N_24969,N_24996);
xnor UO_898 (O_898,N_24871,N_24914);
nand UO_899 (O_899,N_24966,N_24978);
or UO_900 (O_900,N_24805,N_24941);
xnor UO_901 (O_901,N_24882,N_24948);
and UO_902 (O_902,N_24892,N_24806);
nand UO_903 (O_903,N_24982,N_24887);
and UO_904 (O_904,N_24991,N_24998);
or UO_905 (O_905,N_24907,N_24859);
or UO_906 (O_906,N_24780,N_24874);
nand UO_907 (O_907,N_24884,N_24962);
nand UO_908 (O_908,N_24958,N_24809);
nand UO_909 (O_909,N_24903,N_24941);
nor UO_910 (O_910,N_24758,N_24961);
nor UO_911 (O_911,N_24885,N_24771);
nand UO_912 (O_912,N_24924,N_24776);
or UO_913 (O_913,N_24815,N_24786);
and UO_914 (O_914,N_24798,N_24931);
nand UO_915 (O_915,N_24982,N_24859);
and UO_916 (O_916,N_24844,N_24760);
nor UO_917 (O_917,N_24780,N_24854);
or UO_918 (O_918,N_24854,N_24779);
nand UO_919 (O_919,N_24780,N_24994);
nor UO_920 (O_920,N_24882,N_24790);
xnor UO_921 (O_921,N_24897,N_24830);
nor UO_922 (O_922,N_24787,N_24760);
nor UO_923 (O_923,N_24988,N_24871);
and UO_924 (O_924,N_24805,N_24923);
or UO_925 (O_925,N_24988,N_24955);
and UO_926 (O_926,N_24942,N_24905);
nand UO_927 (O_927,N_24977,N_24837);
xnor UO_928 (O_928,N_24858,N_24821);
and UO_929 (O_929,N_24983,N_24886);
nor UO_930 (O_930,N_24926,N_24948);
nand UO_931 (O_931,N_24986,N_24777);
or UO_932 (O_932,N_24755,N_24882);
nand UO_933 (O_933,N_24995,N_24868);
or UO_934 (O_934,N_24982,N_24863);
or UO_935 (O_935,N_24805,N_24999);
and UO_936 (O_936,N_24965,N_24881);
or UO_937 (O_937,N_24764,N_24811);
nor UO_938 (O_938,N_24773,N_24976);
and UO_939 (O_939,N_24841,N_24894);
nand UO_940 (O_940,N_24943,N_24781);
nor UO_941 (O_941,N_24962,N_24758);
nor UO_942 (O_942,N_24953,N_24758);
xor UO_943 (O_943,N_24892,N_24776);
nand UO_944 (O_944,N_24847,N_24959);
xor UO_945 (O_945,N_24764,N_24960);
nor UO_946 (O_946,N_24919,N_24834);
nand UO_947 (O_947,N_24821,N_24764);
xor UO_948 (O_948,N_24840,N_24923);
xor UO_949 (O_949,N_24766,N_24904);
xor UO_950 (O_950,N_24931,N_24895);
nor UO_951 (O_951,N_24842,N_24910);
nor UO_952 (O_952,N_24784,N_24969);
and UO_953 (O_953,N_24763,N_24998);
nor UO_954 (O_954,N_24790,N_24852);
and UO_955 (O_955,N_24913,N_24848);
nand UO_956 (O_956,N_24976,N_24965);
or UO_957 (O_957,N_24808,N_24799);
xnor UO_958 (O_958,N_24785,N_24773);
nor UO_959 (O_959,N_24854,N_24786);
nand UO_960 (O_960,N_24880,N_24873);
nand UO_961 (O_961,N_24803,N_24997);
xor UO_962 (O_962,N_24827,N_24960);
and UO_963 (O_963,N_24937,N_24992);
or UO_964 (O_964,N_24847,N_24832);
nand UO_965 (O_965,N_24986,N_24885);
nor UO_966 (O_966,N_24980,N_24810);
or UO_967 (O_967,N_24786,N_24889);
nand UO_968 (O_968,N_24833,N_24843);
or UO_969 (O_969,N_24878,N_24781);
or UO_970 (O_970,N_24863,N_24873);
and UO_971 (O_971,N_24942,N_24788);
and UO_972 (O_972,N_24791,N_24939);
nor UO_973 (O_973,N_24921,N_24804);
nor UO_974 (O_974,N_24948,N_24819);
nand UO_975 (O_975,N_24845,N_24926);
nor UO_976 (O_976,N_24887,N_24774);
xnor UO_977 (O_977,N_24767,N_24900);
nor UO_978 (O_978,N_24977,N_24817);
xnor UO_979 (O_979,N_24903,N_24776);
xnor UO_980 (O_980,N_24870,N_24957);
or UO_981 (O_981,N_24838,N_24889);
nor UO_982 (O_982,N_24913,N_24858);
nor UO_983 (O_983,N_24935,N_24775);
and UO_984 (O_984,N_24967,N_24830);
and UO_985 (O_985,N_24874,N_24928);
xor UO_986 (O_986,N_24985,N_24784);
nor UO_987 (O_987,N_24966,N_24999);
or UO_988 (O_988,N_24820,N_24865);
nor UO_989 (O_989,N_24836,N_24938);
nor UO_990 (O_990,N_24822,N_24833);
xnor UO_991 (O_991,N_24774,N_24838);
or UO_992 (O_992,N_24920,N_24966);
nor UO_993 (O_993,N_24933,N_24765);
xnor UO_994 (O_994,N_24897,N_24980);
and UO_995 (O_995,N_24833,N_24929);
nor UO_996 (O_996,N_24832,N_24859);
nor UO_997 (O_997,N_24796,N_24850);
and UO_998 (O_998,N_24759,N_24825);
xnor UO_999 (O_999,N_24933,N_24810);
and UO_1000 (O_1000,N_24795,N_24947);
xor UO_1001 (O_1001,N_24966,N_24882);
or UO_1002 (O_1002,N_24864,N_24913);
and UO_1003 (O_1003,N_24909,N_24752);
and UO_1004 (O_1004,N_24819,N_24872);
nand UO_1005 (O_1005,N_24972,N_24846);
nand UO_1006 (O_1006,N_24887,N_24881);
and UO_1007 (O_1007,N_24758,N_24965);
and UO_1008 (O_1008,N_24962,N_24942);
xnor UO_1009 (O_1009,N_24955,N_24850);
nor UO_1010 (O_1010,N_24864,N_24760);
nand UO_1011 (O_1011,N_24799,N_24943);
xnor UO_1012 (O_1012,N_24970,N_24968);
nor UO_1013 (O_1013,N_24972,N_24997);
and UO_1014 (O_1014,N_24839,N_24975);
nand UO_1015 (O_1015,N_24818,N_24861);
xor UO_1016 (O_1016,N_24772,N_24861);
xnor UO_1017 (O_1017,N_24879,N_24793);
or UO_1018 (O_1018,N_24879,N_24823);
xor UO_1019 (O_1019,N_24959,N_24762);
nand UO_1020 (O_1020,N_24929,N_24883);
or UO_1021 (O_1021,N_24835,N_24855);
xnor UO_1022 (O_1022,N_24762,N_24830);
nand UO_1023 (O_1023,N_24995,N_24819);
nand UO_1024 (O_1024,N_24982,N_24866);
and UO_1025 (O_1025,N_24754,N_24847);
xor UO_1026 (O_1026,N_24822,N_24952);
nand UO_1027 (O_1027,N_24932,N_24952);
nor UO_1028 (O_1028,N_24844,N_24995);
nand UO_1029 (O_1029,N_24771,N_24786);
and UO_1030 (O_1030,N_24980,N_24887);
nand UO_1031 (O_1031,N_24905,N_24959);
nand UO_1032 (O_1032,N_24941,N_24977);
nor UO_1033 (O_1033,N_24787,N_24837);
xnor UO_1034 (O_1034,N_24844,N_24976);
or UO_1035 (O_1035,N_24959,N_24966);
nor UO_1036 (O_1036,N_24792,N_24769);
or UO_1037 (O_1037,N_24813,N_24972);
and UO_1038 (O_1038,N_24878,N_24852);
nor UO_1039 (O_1039,N_24786,N_24806);
nand UO_1040 (O_1040,N_24955,N_24944);
and UO_1041 (O_1041,N_24803,N_24786);
and UO_1042 (O_1042,N_24779,N_24836);
and UO_1043 (O_1043,N_24917,N_24847);
nor UO_1044 (O_1044,N_24826,N_24981);
nor UO_1045 (O_1045,N_24914,N_24783);
nor UO_1046 (O_1046,N_24905,N_24855);
and UO_1047 (O_1047,N_24888,N_24916);
xor UO_1048 (O_1048,N_24932,N_24939);
and UO_1049 (O_1049,N_24934,N_24821);
nand UO_1050 (O_1050,N_24929,N_24928);
and UO_1051 (O_1051,N_24819,N_24900);
nand UO_1052 (O_1052,N_24863,N_24934);
nor UO_1053 (O_1053,N_24886,N_24980);
xnor UO_1054 (O_1054,N_24904,N_24887);
xnor UO_1055 (O_1055,N_24893,N_24908);
xnor UO_1056 (O_1056,N_24985,N_24863);
nand UO_1057 (O_1057,N_24912,N_24926);
xnor UO_1058 (O_1058,N_24851,N_24848);
xor UO_1059 (O_1059,N_24782,N_24768);
nand UO_1060 (O_1060,N_24774,N_24801);
and UO_1061 (O_1061,N_24818,N_24765);
or UO_1062 (O_1062,N_24867,N_24893);
and UO_1063 (O_1063,N_24933,N_24952);
nand UO_1064 (O_1064,N_24866,N_24766);
or UO_1065 (O_1065,N_24788,N_24775);
nor UO_1066 (O_1066,N_24797,N_24804);
or UO_1067 (O_1067,N_24760,N_24900);
nand UO_1068 (O_1068,N_24992,N_24772);
xnor UO_1069 (O_1069,N_24885,N_24872);
and UO_1070 (O_1070,N_24803,N_24804);
or UO_1071 (O_1071,N_24949,N_24977);
xor UO_1072 (O_1072,N_24962,N_24979);
or UO_1073 (O_1073,N_24899,N_24916);
nand UO_1074 (O_1074,N_24905,N_24875);
nor UO_1075 (O_1075,N_24953,N_24903);
or UO_1076 (O_1076,N_24991,N_24885);
nor UO_1077 (O_1077,N_24853,N_24985);
nor UO_1078 (O_1078,N_24753,N_24980);
and UO_1079 (O_1079,N_24940,N_24910);
xor UO_1080 (O_1080,N_24798,N_24788);
nor UO_1081 (O_1081,N_24805,N_24877);
and UO_1082 (O_1082,N_24761,N_24913);
nand UO_1083 (O_1083,N_24754,N_24920);
nor UO_1084 (O_1084,N_24846,N_24800);
xnor UO_1085 (O_1085,N_24781,N_24772);
xnor UO_1086 (O_1086,N_24912,N_24760);
xor UO_1087 (O_1087,N_24816,N_24812);
xor UO_1088 (O_1088,N_24888,N_24832);
nor UO_1089 (O_1089,N_24993,N_24895);
nand UO_1090 (O_1090,N_24992,N_24877);
nor UO_1091 (O_1091,N_24792,N_24907);
nand UO_1092 (O_1092,N_24928,N_24758);
or UO_1093 (O_1093,N_24950,N_24975);
nor UO_1094 (O_1094,N_24968,N_24771);
xnor UO_1095 (O_1095,N_24752,N_24812);
nor UO_1096 (O_1096,N_24827,N_24951);
nand UO_1097 (O_1097,N_24938,N_24780);
nand UO_1098 (O_1098,N_24947,N_24990);
and UO_1099 (O_1099,N_24797,N_24998);
nand UO_1100 (O_1100,N_24817,N_24810);
nor UO_1101 (O_1101,N_24807,N_24940);
xnor UO_1102 (O_1102,N_24813,N_24984);
xor UO_1103 (O_1103,N_24902,N_24758);
or UO_1104 (O_1104,N_24922,N_24891);
or UO_1105 (O_1105,N_24961,N_24988);
nand UO_1106 (O_1106,N_24935,N_24925);
and UO_1107 (O_1107,N_24873,N_24883);
nor UO_1108 (O_1108,N_24911,N_24923);
and UO_1109 (O_1109,N_24869,N_24754);
xor UO_1110 (O_1110,N_24940,N_24963);
nor UO_1111 (O_1111,N_24910,N_24833);
nor UO_1112 (O_1112,N_24799,N_24985);
nor UO_1113 (O_1113,N_24775,N_24839);
nand UO_1114 (O_1114,N_24751,N_24833);
nand UO_1115 (O_1115,N_24950,N_24805);
and UO_1116 (O_1116,N_24962,N_24910);
and UO_1117 (O_1117,N_24886,N_24797);
or UO_1118 (O_1118,N_24882,N_24834);
and UO_1119 (O_1119,N_24954,N_24881);
nand UO_1120 (O_1120,N_24781,N_24765);
nand UO_1121 (O_1121,N_24856,N_24960);
or UO_1122 (O_1122,N_24809,N_24980);
nor UO_1123 (O_1123,N_24870,N_24868);
and UO_1124 (O_1124,N_24908,N_24838);
and UO_1125 (O_1125,N_24921,N_24928);
and UO_1126 (O_1126,N_24774,N_24809);
or UO_1127 (O_1127,N_24826,N_24789);
nand UO_1128 (O_1128,N_24954,N_24812);
or UO_1129 (O_1129,N_24857,N_24926);
or UO_1130 (O_1130,N_24789,N_24847);
xor UO_1131 (O_1131,N_24832,N_24970);
and UO_1132 (O_1132,N_24876,N_24852);
xnor UO_1133 (O_1133,N_24901,N_24844);
xnor UO_1134 (O_1134,N_24857,N_24879);
nand UO_1135 (O_1135,N_24880,N_24920);
and UO_1136 (O_1136,N_24877,N_24962);
or UO_1137 (O_1137,N_24878,N_24924);
and UO_1138 (O_1138,N_24878,N_24775);
nand UO_1139 (O_1139,N_24893,N_24960);
xor UO_1140 (O_1140,N_24970,N_24790);
nand UO_1141 (O_1141,N_24792,N_24911);
or UO_1142 (O_1142,N_24962,N_24820);
or UO_1143 (O_1143,N_24849,N_24805);
and UO_1144 (O_1144,N_24949,N_24885);
or UO_1145 (O_1145,N_24857,N_24844);
nand UO_1146 (O_1146,N_24914,N_24765);
nand UO_1147 (O_1147,N_24990,N_24851);
and UO_1148 (O_1148,N_24857,N_24790);
nor UO_1149 (O_1149,N_24883,N_24979);
or UO_1150 (O_1150,N_24896,N_24861);
or UO_1151 (O_1151,N_24767,N_24766);
nand UO_1152 (O_1152,N_24983,N_24977);
xnor UO_1153 (O_1153,N_24871,N_24851);
nand UO_1154 (O_1154,N_24839,N_24831);
or UO_1155 (O_1155,N_24893,N_24870);
or UO_1156 (O_1156,N_24971,N_24942);
nor UO_1157 (O_1157,N_24994,N_24908);
xnor UO_1158 (O_1158,N_24751,N_24911);
nand UO_1159 (O_1159,N_24955,N_24861);
or UO_1160 (O_1160,N_24914,N_24963);
or UO_1161 (O_1161,N_24843,N_24914);
and UO_1162 (O_1162,N_24951,N_24766);
or UO_1163 (O_1163,N_24759,N_24916);
xnor UO_1164 (O_1164,N_24924,N_24953);
xor UO_1165 (O_1165,N_24755,N_24785);
or UO_1166 (O_1166,N_24809,N_24858);
and UO_1167 (O_1167,N_24883,N_24919);
xor UO_1168 (O_1168,N_24853,N_24944);
xor UO_1169 (O_1169,N_24842,N_24871);
nand UO_1170 (O_1170,N_24790,N_24998);
or UO_1171 (O_1171,N_24832,N_24768);
nor UO_1172 (O_1172,N_24810,N_24813);
xor UO_1173 (O_1173,N_24829,N_24812);
nor UO_1174 (O_1174,N_24804,N_24766);
xor UO_1175 (O_1175,N_24763,N_24799);
and UO_1176 (O_1176,N_24880,N_24813);
or UO_1177 (O_1177,N_24889,N_24768);
and UO_1178 (O_1178,N_24899,N_24843);
nand UO_1179 (O_1179,N_24753,N_24866);
nor UO_1180 (O_1180,N_24997,N_24826);
nor UO_1181 (O_1181,N_24861,N_24920);
and UO_1182 (O_1182,N_24929,N_24880);
or UO_1183 (O_1183,N_24864,N_24842);
xnor UO_1184 (O_1184,N_24894,N_24919);
nand UO_1185 (O_1185,N_24832,N_24943);
xor UO_1186 (O_1186,N_24838,N_24929);
or UO_1187 (O_1187,N_24959,N_24938);
xor UO_1188 (O_1188,N_24777,N_24862);
nand UO_1189 (O_1189,N_24941,N_24857);
or UO_1190 (O_1190,N_24867,N_24820);
and UO_1191 (O_1191,N_24871,N_24875);
nand UO_1192 (O_1192,N_24893,N_24964);
nor UO_1193 (O_1193,N_24752,N_24785);
or UO_1194 (O_1194,N_24820,N_24920);
xnor UO_1195 (O_1195,N_24752,N_24788);
and UO_1196 (O_1196,N_24922,N_24850);
and UO_1197 (O_1197,N_24950,N_24949);
and UO_1198 (O_1198,N_24903,N_24993);
or UO_1199 (O_1199,N_24877,N_24967);
nand UO_1200 (O_1200,N_24909,N_24797);
nand UO_1201 (O_1201,N_24811,N_24909);
nor UO_1202 (O_1202,N_24775,N_24889);
nand UO_1203 (O_1203,N_24967,N_24925);
and UO_1204 (O_1204,N_24892,N_24924);
nand UO_1205 (O_1205,N_24809,N_24944);
xor UO_1206 (O_1206,N_24856,N_24767);
or UO_1207 (O_1207,N_24850,N_24825);
xor UO_1208 (O_1208,N_24901,N_24755);
nor UO_1209 (O_1209,N_24781,N_24945);
or UO_1210 (O_1210,N_24864,N_24857);
or UO_1211 (O_1211,N_24765,N_24966);
xor UO_1212 (O_1212,N_24922,N_24994);
nand UO_1213 (O_1213,N_24755,N_24825);
and UO_1214 (O_1214,N_24821,N_24964);
and UO_1215 (O_1215,N_24767,N_24961);
xor UO_1216 (O_1216,N_24807,N_24947);
xnor UO_1217 (O_1217,N_24992,N_24998);
nand UO_1218 (O_1218,N_24968,N_24770);
xnor UO_1219 (O_1219,N_24772,N_24886);
nor UO_1220 (O_1220,N_24799,N_24814);
or UO_1221 (O_1221,N_24890,N_24757);
or UO_1222 (O_1222,N_24961,N_24896);
xnor UO_1223 (O_1223,N_24965,N_24962);
xnor UO_1224 (O_1224,N_24944,N_24903);
or UO_1225 (O_1225,N_24797,N_24812);
and UO_1226 (O_1226,N_24987,N_24941);
nand UO_1227 (O_1227,N_24824,N_24964);
or UO_1228 (O_1228,N_24877,N_24799);
and UO_1229 (O_1229,N_24773,N_24808);
nand UO_1230 (O_1230,N_24938,N_24819);
nand UO_1231 (O_1231,N_24765,N_24927);
or UO_1232 (O_1232,N_24828,N_24974);
nand UO_1233 (O_1233,N_24929,N_24865);
nand UO_1234 (O_1234,N_24849,N_24924);
and UO_1235 (O_1235,N_24966,N_24919);
nor UO_1236 (O_1236,N_24782,N_24773);
nor UO_1237 (O_1237,N_24869,N_24879);
nor UO_1238 (O_1238,N_24753,N_24835);
and UO_1239 (O_1239,N_24948,N_24859);
and UO_1240 (O_1240,N_24808,N_24819);
xnor UO_1241 (O_1241,N_24840,N_24926);
nand UO_1242 (O_1242,N_24989,N_24776);
nand UO_1243 (O_1243,N_24865,N_24853);
nor UO_1244 (O_1244,N_24903,N_24974);
nand UO_1245 (O_1245,N_24976,N_24769);
or UO_1246 (O_1246,N_24976,N_24939);
nand UO_1247 (O_1247,N_24806,N_24990);
or UO_1248 (O_1248,N_24862,N_24908);
nand UO_1249 (O_1249,N_24832,N_24900);
xnor UO_1250 (O_1250,N_24883,N_24944);
xor UO_1251 (O_1251,N_24866,N_24925);
nand UO_1252 (O_1252,N_24985,N_24931);
and UO_1253 (O_1253,N_24914,N_24927);
nand UO_1254 (O_1254,N_24889,N_24970);
xor UO_1255 (O_1255,N_24925,N_24811);
nand UO_1256 (O_1256,N_24791,N_24757);
and UO_1257 (O_1257,N_24885,N_24768);
xor UO_1258 (O_1258,N_24847,N_24873);
nor UO_1259 (O_1259,N_24889,N_24957);
nand UO_1260 (O_1260,N_24814,N_24939);
or UO_1261 (O_1261,N_24888,N_24907);
xor UO_1262 (O_1262,N_24952,N_24779);
nor UO_1263 (O_1263,N_24891,N_24867);
nand UO_1264 (O_1264,N_24802,N_24963);
or UO_1265 (O_1265,N_24961,N_24965);
nand UO_1266 (O_1266,N_24841,N_24887);
or UO_1267 (O_1267,N_24954,N_24829);
nand UO_1268 (O_1268,N_24772,N_24983);
nand UO_1269 (O_1269,N_24805,N_24818);
nand UO_1270 (O_1270,N_24916,N_24757);
or UO_1271 (O_1271,N_24990,N_24854);
xnor UO_1272 (O_1272,N_24814,N_24958);
xnor UO_1273 (O_1273,N_24856,N_24949);
xor UO_1274 (O_1274,N_24851,N_24869);
nor UO_1275 (O_1275,N_24963,N_24908);
xnor UO_1276 (O_1276,N_24948,N_24807);
or UO_1277 (O_1277,N_24980,N_24918);
and UO_1278 (O_1278,N_24774,N_24778);
or UO_1279 (O_1279,N_24823,N_24807);
xnor UO_1280 (O_1280,N_24996,N_24947);
nor UO_1281 (O_1281,N_24929,N_24761);
nand UO_1282 (O_1282,N_24894,N_24895);
xor UO_1283 (O_1283,N_24872,N_24843);
xor UO_1284 (O_1284,N_24972,N_24959);
nand UO_1285 (O_1285,N_24917,N_24938);
nor UO_1286 (O_1286,N_24852,N_24944);
or UO_1287 (O_1287,N_24836,N_24993);
xnor UO_1288 (O_1288,N_24796,N_24786);
or UO_1289 (O_1289,N_24852,N_24848);
xor UO_1290 (O_1290,N_24886,N_24885);
nor UO_1291 (O_1291,N_24805,N_24760);
nand UO_1292 (O_1292,N_24951,N_24772);
xor UO_1293 (O_1293,N_24987,N_24794);
nand UO_1294 (O_1294,N_24875,N_24960);
or UO_1295 (O_1295,N_24775,N_24858);
or UO_1296 (O_1296,N_24962,N_24830);
and UO_1297 (O_1297,N_24917,N_24823);
nand UO_1298 (O_1298,N_24978,N_24958);
and UO_1299 (O_1299,N_24819,N_24917);
nor UO_1300 (O_1300,N_24997,N_24750);
and UO_1301 (O_1301,N_24926,N_24914);
or UO_1302 (O_1302,N_24978,N_24866);
xor UO_1303 (O_1303,N_24936,N_24830);
nand UO_1304 (O_1304,N_24873,N_24817);
and UO_1305 (O_1305,N_24783,N_24806);
xnor UO_1306 (O_1306,N_24760,N_24921);
nor UO_1307 (O_1307,N_24934,N_24859);
or UO_1308 (O_1308,N_24802,N_24874);
nor UO_1309 (O_1309,N_24935,N_24941);
and UO_1310 (O_1310,N_24764,N_24961);
nand UO_1311 (O_1311,N_24847,N_24989);
xnor UO_1312 (O_1312,N_24813,N_24902);
or UO_1313 (O_1313,N_24793,N_24883);
or UO_1314 (O_1314,N_24956,N_24888);
nor UO_1315 (O_1315,N_24942,N_24866);
or UO_1316 (O_1316,N_24892,N_24869);
nor UO_1317 (O_1317,N_24943,N_24878);
or UO_1318 (O_1318,N_24990,N_24789);
nand UO_1319 (O_1319,N_24995,N_24962);
xor UO_1320 (O_1320,N_24906,N_24905);
nand UO_1321 (O_1321,N_24978,N_24976);
or UO_1322 (O_1322,N_24933,N_24752);
or UO_1323 (O_1323,N_24856,N_24850);
xor UO_1324 (O_1324,N_24886,N_24949);
nor UO_1325 (O_1325,N_24957,N_24909);
or UO_1326 (O_1326,N_24962,N_24760);
xnor UO_1327 (O_1327,N_24968,N_24811);
nand UO_1328 (O_1328,N_24905,N_24930);
xnor UO_1329 (O_1329,N_24988,N_24858);
or UO_1330 (O_1330,N_24817,N_24801);
and UO_1331 (O_1331,N_24833,N_24893);
and UO_1332 (O_1332,N_24762,N_24974);
xnor UO_1333 (O_1333,N_24878,N_24751);
nor UO_1334 (O_1334,N_24799,N_24788);
and UO_1335 (O_1335,N_24818,N_24931);
or UO_1336 (O_1336,N_24983,N_24761);
nor UO_1337 (O_1337,N_24751,N_24797);
nand UO_1338 (O_1338,N_24952,N_24833);
nor UO_1339 (O_1339,N_24798,N_24870);
xor UO_1340 (O_1340,N_24851,N_24949);
xor UO_1341 (O_1341,N_24960,N_24973);
nor UO_1342 (O_1342,N_24878,N_24898);
or UO_1343 (O_1343,N_24918,N_24802);
nor UO_1344 (O_1344,N_24978,N_24893);
and UO_1345 (O_1345,N_24799,N_24795);
or UO_1346 (O_1346,N_24975,N_24796);
xnor UO_1347 (O_1347,N_24905,N_24867);
nand UO_1348 (O_1348,N_24875,N_24789);
xor UO_1349 (O_1349,N_24877,N_24893);
xor UO_1350 (O_1350,N_24966,N_24941);
xnor UO_1351 (O_1351,N_24859,N_24810);
or UO_1352 (O_1352,N_24879,N_24958);
xnor UO_1353 (O_1353,N_24781,N_24886);
nor UO_1354 (O_1354,N_24873,N_24833);
and UO_1355 (O_1355,N_24848,N_24969);
xnor UO_1356 (O_1356,N_24832,N_24919);
and UO_1357 (O_1357,N_24759,N_24928);
and UO_1358 (O_1358,N_24780,N_24766);
nand UO_1359 (O_1359,N_24835,N_24971);
or UO_1360 (O_1360,N_24829,N_24915);
nand UO_1361 (O_1361,N_24966,N_24894);
nor UO_1362 (O_1362,N_24926,N_24942);
xor UO_1363 (O_1363,N_24947,N_24852);
and UO_1364 (O_1364,N_24772,N_24821);
xor UO_1365 (O_1365,N_24957,N_24783);
nand UO_1366 (O_1366,N_24927,N_24892);
or UO_1367 (O_1367,N_24807,N_24783);
and UO_1368 (O_1368,N_24821,N_24794);
xnor UO_1369 (O_1369,N_24779,N_24845);
or UO_1370 (O_1370,N_24957,N_24916);
and UO_1371 (O_1371,N_24865,N_24983);
nor UO_1372 (O_1372,N_24799,N_24946);
nand UO_1373 (O_1373,N_24852,N_24925);
nor UO_1374 (O_1374,N_24807,N_24765);
and UO_1375 (O_1375,N_24766,N_24865);
and UO_1376 (O_1376,N_24935,N_24779);
and UO_1377 (O_1377,N_24879,N_24980);
xnor UO_1378 (O_1378,N_24918,N_24903);
xnor UO_1379 (O_1379,N_24974,N_24889);
xnor UO_1380 (O_1380,N_24820,N_24998);
or UO_1381 (O_1381,N_24769,N_24915);
xnor UO_1382 (O_1382,N_24928,N_24791);
and UO_1383 (O_1383,N_24768,N_24814);
nand UO_1384 (O_1384,N_24786,N_24757);
or UO_1385 (O_1385,N_24894,N_24816);
or UO_1386 (O_1386,N_24870,N_24898);
and UO_1387 (O_1387,N_24842,N_24783);
and UO_1388 (O_1388,N_24952,N_24790);
nand UO_1389 (O_1389,N_24870,N_24862);
nor UO_1390 (O_1390,N_24896,N_24763);
or UO_1391 (O_1391,N_24795,N_24977);
xnor UO_1392 (O_1392,N_24756,N_24967);
nor UO_1393 (O_1393,N_24926,N_24755);
and UO_1394 (O_1394,N_24806,N_24814);
and UO_1395 (O_1395,N_24911,N_24870);
nand UO_1396 (O_1396,N_24834,N_24915);
nor UO_1397 (O_1397,N_24824,N_24922);
xnor UO_1398 (O_1398,N_24803,N_24890);
nor UO_1399 (O_1399,N_24897,N_24852);
or UO_1400 (O_1400,N_24841,N_24822);
nand UO_1401 (O_1401,N_24765,N_24928);
xor UO_1402 (O_1402,N_24982,N_24804);
xor UO_1403 (O_1403,N_24920,N_24943);
xnor UO_1404 (O_1404,N_24884,N_24965);
and UO_1405 (O_1405,N_24904,N_24859);
xor UO_1406 (O_1406,N_24848,N_24838);
nand UO_1407 (O_1407,N_24862,N_24880);
nor UO_1408 (O_1408,N_24867,N_24843);
and UO_1409 (O_1409,N_24772,N_24775);
xor UO_1410 (O_1410,N_24836,N_24926);
or UO_1411 (O_1411,N_24979,N_24814);
and UO_1412 (O_1412,N_24795,N_24872);
and UO_1413 (O_1413,N_24762,N_24772);
nor UO_1414 (O_1414,N_24856,N_24808);
and UO_1415 (O_1415,N_24813,N_24985);
xor UO_1416 (O_1416,N_24957,N_24848);
or UO_1417 (O_1417,N_24788,N_24883);
xnor UO_1418 (O_1418,N_24921,N_24886);
or UO_1419 (O_1419,N_24758,N_24970);
xnor UO_1420 (O_1420,N_24885,N_24954);
or UO_1421 (O_1421,N_24947,N_24899);
xor UO_1422 (O_1422,N_24950,N_24917);
or UO_1423 (O_1423,N_24969,N_24914);
nand UO_1424 (O_1424,N_24891,N_24898);
or UO_1425 (O_1425,N_24805,N_24939);
or UO_1426 (O_1426,N_24794,N_24929);
nand UO_1427 (O_1427,N_24952,N_24861);
or UO_1428 (O_1428,N_24871,N_24848);
xor UO_1429 (O_1429,N_24997,N_24755);
or UO_1430 (O_1430,N_24819,N_24779);
or UO_1431 (O_1431,N_24752,N_24925);
or UO_1432 (O_1432,N_24865,N_24872);
or UO_1433 (O_1433,N_24880,N_24994);
or UO_1434 (O_1434,N_24936,N_24887);
nand UO_1435 (O_1435,N_24847,N_24982);
or UO_1436 (O_1436,N_24971,N_24751);
or UO_1437 (O_1437,N_24820,N_24871);
and UO_1438 (O_1438,N_24897,N_24949);
nand UO_1439 (O_1439,N_24766,N_24790);
nor UO_1440 (O_1440,N_24867,N_24754);
xor UO_1441 (O_1441,N_24870,N_24912);
xnor UO_1442 (O_1442,N_24863,N_24861);
or UO_1443 (O_1443,N_24832,N_24842);
xor UO_1444 (O_1444,N_24837,N_24850);
and UO_1445 (O_1445,N_24863,N_24838);
and UO_1446 (O_1446,N_24981,N_24936);
and UO_1447 (O_1447,N_24859,N_24840);
xor UO_1448 (O_1448,N_24918,N_24959);
xor UO_1449 (O_1449,N_24777,N_24848);
and UO_1450 (O_1450,N_24982,N_24938);
nor UO_1451 (O_1451,N_24859,N_24936);
nor UO_1452 (O_1452,N_24811,N_24914);
nor UO_1453 (O_1453,N_24999,N_24827);
nand UO_1454 (O_1454,N_24938,N_24761);
or UO_1455 (O_1455,N_24862,N_24846);
nand UO_1456 (O_1456,N_24781,N_24995);
or UO_1457 (O_1457,N_24782,N_24862);
nand UO_1458 (O_1458,N_24996,N_24987);
or UO_1459 (O_1459,N_24829,N_24822);
and UO_1460 (O_1460,N_24955,N_24868);
and UO_1461 (O_1461,N_24816,N_24964);
nand UO_1462 (O_1462,N_24947,N_24972);
nand UO_1463 (O_1463,N_24932,N_24859);
and UO_1464 (O_1464,N_24996,N_24830);
or UO_1465 (O_1465,N_24925,N_24846);
or UO_1466 (O_1466,N_24875,N_24864);
or UO_1467 (O_1467,N_24834,N_24921);
and UO_1468 (O_1468,N_24820,N_24854);
xor UO_1469 (O_1469,N_24928,N_24775);
xnor UO_1470 (O_1470,N_24968,N_24975);
or UO_1471 (O_1471,N_24962,N_24890);
and UO_1472 (O_1472,N_24949,N_24859);
xor UO_1473 (O_1473,N_24790,N_24977);
xnor UO_1474 (O_1474,N_24826,N_24958);
and UO_1475 (O_1475,N_24801,N_24929);
nand UO_1476 (O_1476,N_24997,N_24825);
nor UO_1477 (O_1477,N_24983,N_24995);
nor UO_1478 (O_1478,N_24903,N_24890);
nor UO_1479 (O_1479,N_24809,N_24750);
xor UO_1480 (O_1480,N_24935,N_24976);
nor UO_1481 (O_1481,N_24800,N_24781);
xnor UO_1482 (O_1482,N_24861,N_24919);
and UO_1483 (O_1483,N_24950,N_24882);
xnor UO_1484 (O_1484,N_24756,N_24923);
and UO_1485 (O_1485,N_24939,N_24914);
nand UO_1486 (O_1486,N_24951,N_24952);
and UO_1487 (O_1487,N_24941,N_24962);
nor UO_1488 (O_1488,N_24975,N_24824);
or UO_1489 (O_1489,N_24951,N_24759);
nor UO_1490 (O_1490,N_24980,N_24864);
xor UO_1491 (O_1491,N_24826,N_24810);
or UO_1492 (O_1492,N_24757,N_24834);
and UO_1493 (O_1493,N_24934,N_24758);
or UO_1494 (O_1494,N_24936,N_24774);
xor UO_1495 (O_1495,N_24968,N_24760);
or UO_1496 (O_1496,N_24986,N_24895);
nand UO_1497 (O_1497,N_24821,N_24785);
nand UO_1498 (O_1498,N_24822,N_24869);
xor UO_1499 (O_1499,N_24951,N_24866);
xnor UO_1500 (O_1500,N_24863,N_24761);
nor UO_1501 (O_1501,N_24767,N_24848);
and UO_1502 (O_1502,N_24896,N_24780);
nor UO_1503 (O_1503,N_24906,N_24976);
and UO_1504 (O_1504,N_24995,N_24895);
nand UO_1505 (O_1505,N_24956,N_24880);
xor UO_1506 (O_1506,N_24804,N_24941);
xor UO_1507 (O_1507,N_24841,N_24939);
nand UO_1508 (O_1508,N_24885,N_24940);
xor UO_1509 (O_1509,N_24841,N_24875);
and UO_1510 (O_1510,N_24970,N_24942);
nor UO_1511 (O_1511,N_24947,N_24750);
nand UO_1512 (O_1512,N_24892,N_24837);
nor UO_1513 (O_1513,N_24978,N_24872);
and UO_1514 (O_1514,N_24842,N_24886);
nand UO_1515 (O_1515,N_24799,N_24897);
xnor UO_1516 (O_1516,N_24899,N_24901);
nor UO_1517 (O_1517,N_24985,N_24926);
and UO_1518 (O_1518,N_24884,N_24798);
nor UO_1519 (O_1519,N_24981,N_24860);
or UO_1520 (O_1520,N_24915,N_24882);
xor UO_1521 (O_1521,N_24947,N_24850);
nand UO_1522 (O_1522,N_24864,N_24839);
xor UO_1523 (O_1523,N_24980,N_24861);
nor UO_1524 (O_1524,N_24794,N_24817);
or UO_1525 (O_1525,N_24882,N_24952);
nor UO_1526 (O_1526,N_24773,N_24918);
nand UO_1527 (O_1527,N_24891,N_24994);
nor UO_1528 (O_1528,N_24996,N_24883);
xor UO_1529 (O_1529,N_24870,N_24782);
xor UO_1530 (O_1530,N_24988,N_24775);
and UO_1531 (O_1531,N_24851,N_24780);
nor UO_1532 (O_1532,N_24995,N_24860);
xnor UO_1533 (O_1533,N_24762,N_24854);
nor UO_1534 (O_1534,N_24891,N_24774);
nor UO_1535 (O_1535,N_24952,N_24934);
xnor UO_1536 (O_1536,N_24981,N_24762);
or UO_1537 (O_1537,N_24832,N_24808);
and UO_1538 (O_1538,N_24894,N_24902);
and UO_1539 (O_1539,N_24821,N_24848);
xnor UO_1540 (O_1540,N_24940,N_24995);
nand UO_1541 (O_1541,N_24846,N_24997);
xnor UO_1542 (O_1542,N_24756,N_24953);
nor UO_1543 (O_1543,N_24764,N_24784);
or UO_1544 (O_1544,N_24807,N_24986);
nor UO_1545 (O_1545,N_24995,N_24925);
xnor UO_1546 (O_1546,N_24984,N_24837);
nand UO_1547 (O_1547,N_24834,N_24828);
or UO_1548 (O_1548,N_24976,N_24790);
xor UO_1549 (O_1549,N_24777,N_24932);
nand UO_1550 (O_1550,N_24989,N_24963);
xor UO_1551 (O_1551,N_24959,N_24870);
or UO_1552 (O_1552,N_24753,N_24918);
and UO_1553 (O_1553,N_24898,N_24973);
or UO_1554 (O_1554,N_24888,N_24753);
nor UO_1555 (O_1555,N_24848,N_24789);
or UO_1556 (O_1556,N_24880,N_24753);
nor UO_1557 (O_1557,N_24807,N_24811);
xor UO_1558 (O_1558,N_24932,N_24940);
and UO_1559 (O_1559,N_24872,N_24901);
or UO_1560 (O_1560,N_24986,N_24981);
xor UO_1561 (O_1561,N_24970,N_24752);
nand UO_1562 (O_1562,N_24994,N_24874);
nor UO_1563 (O_1563,N_24814,N_24895);
xor UO_1564 (O_1564,N_24838,N_24991);
xor UO_1565 (O_1565,N_24858,N_24963);
nand UO_1566 (O_1566,N_24947,N_24759);
or UO_1567 (O_1567,N_24926,N_24783);
and UO_1568 (O_1568,N_24812,N_24815);
or UO_1569 (O_1569,N_24947,N_24862);
xnor UO_1570 (O_1570,N_24792,N_24952);
and UO_1571 (O_1571,N_24977,N_24842);
xnor UO_1572 (O_1572,N_24841,N_24802);
and UO_1573 (O_1573,N_24962,N_24986);
or UO_1574 (O_1574,N_24976,N_24998);
xor UO_1575 (O_1575,N_24760,N_24774);
or UO_1576 (O_1576,N_24783,N_24915);
nand UO_1577 (O_1577,N_24891,N_24780);
nor UO_1578 (O_1578,N_24955,N_24805);
or UO_1579 (O_1579,N_24977,N_24930);
xnor UO_1580 (O_1580,N_24856,N_24757);
and UO_1581 (O_1581,N_24823,N_24910);
nor UO_1582 (O_1582,N_24800,N_24806);
or UO_1583 (O_1583,N_24958,N_24759);
nand UO_1584 (O_1584,N_24910,N_24895);
or UO_1585 (O_1585,N_24820,N_24893);
nand UO_1586 (O_1586,N_24910,N_24952);
xor UO_1587 (O_1587,N_24967,N_24938);
nor UO_1588 (O_1588,N_24855,N_24949);
or UO_1589 (O_1589,N_24828,N_24800);
or UO_1590 (O_1590,N_24918,N_24794);
nor UO_1591 (O_1591,N_24766,N_24910);
nand UO_1592 (O_1592,N_24778,N_24766);
or UO_1593 (O_1593,N_24789,N_24873);
nor UO_1594 (O_1594,N_24809,N_24921);
and UO_1595 (O_1595,N_24909,N_24998);
and UO_1596 (O_1596,N_24789,N_24928);
xor UO_1597 (O_1597,N_24909,N_24836);
and UO_1598 (O_1598,N_24819,N_24927);
nor UO_1599 (O_1599,N_24956,N_24847);
xor UO_1600 (O_1600,N_24893,N_24984);
and UO_1601 (O_1601,N_24985,N_24793);
and UO_1602 (O_1602,N_24931,N_24848);
and UO_1603 (O_1603,N_24787,N_24823);
nand UO_1604 (O_1604,N_24989,N_24950);
nor UO_1605 (O_1605,N_24856,N_24970);
and UO_1606 (O_1606,N_24957,N_24921);
and UO_1607 (O_1607,N_24832,N_24795);
xnor UO_1608 (O_1608,N_24761,N_24970);
xor UO_1609 (O_1609,N_24969,N_24851);
and UO_1610 (O_1610,N_24997,N_24790);
xnor UO_1611 (O_1611,N_24897,N_24922);
nand UO_1612 (O_1612,N_24860,N_24902);
nand UO_1613 (O_1613,N_24762,N_24996);
and UO_1614 (O_1614,N_24835,N_24819);
xnor UO_1615 (O_1615,N_24941,N_24802);
xor UO_1616 (O_1616,N_24846,N_24961);
nand UO_1617 (O_1617,N_24906,N_24788);
nor UO_1618 (O_1618,N_24934,N_24814);
and UO_1619 (O_1619,N_24779,N_24910);
nor UO_1620 (O_1620,N_24825,N_24936);
nor UO_1621 (O_1621,N_24986,N_24766);
or UO_1622 (O_1622,N_24956,N_24959);
nand UO_1623 (O_1623,N_24782,N_24942);
and UO_1624 (O_1624,N_24895,N_24893);
or UO_1625 (O_1625,N_24836,N_24825);
nor UO_1626 (O_1626,N_24834,N_24990);
and UO_1627 (O_1627,N_24829,N_24926);
nand UO_1628 (O_1628,N_24757,N_24785);
nand UO_1629 (O_1629,N_24984,N_24935);
nand UO_1630 (O_1630,N_24766,N_24971);
xor UO_1631 (O_1631,N_24930,N_24761);
or UO_1632 (O_1632,N_24923,N_24936);
xor UO_1633 (O_1633,N_24984,N_24782);
or UO_1634 (O_1634,N_24873,N_24776);
and UO_1635 (O_1635,N_24788,N_24999);
and UO_1636 (O_1636,N_24987,N_24961);
nor UO_1637 (O_1637,N_24778,N_24888);
and UO_1638 (O_1638,N_24933,N_24758);
xor UO_1639 (O_1639,N_24812,N_24981);
or UO_1640 (O_1640,N_24796,N_24963);
and UO_1641 (O_1641,N_24772,N_24780);
or UO_1642 (O_1642,N_24801,N_24792);
or UO_1643 (O_1643,N_24751,N_24935);
and UO_1644 (O_1644,N_24855,N_24881);
nand UO_1645 (O_1645,N_24977,N_24865);
nor UO_1646 (O_1646,N_24956,N_24789);
and UO_1647 (O_1647,N_24995,N_24923);
nand UO_1648 (O_1648,N_24894,N_24934);
or UO_1649 (O_1649,N_24774,N_24895);
nor UO_1650 (O_1650,N_24753,N_24874);
xnor UO_1651 (O_1651,N_24906,N_24764);
nand UO_1652 (O_1652,N_24910,N_24988);
and UO_1653 (O_1653,N_24985,N_24854);
nand UO_1654 (O_1654,N_24904,N_24942);
nand UO_1655 (O_1655,N_24809,N_24783);
nand UO_1656 (O_1656,N_24878,N_24763);
nor UO_1657 (O_1657,N_24856,N_24987);
and UO_1658 (O_1658,N_24911,N_24823);
and UO_1659 (O_1659,N_24935,N_24992);
nand UO_1660 (O_1660,N_24875,N_24974);
nand UO_1661 (O_1661,N_24876,N_24799);
xnor UO_1662 (O_1662,N_24900,N_24854);
xnor UO_1663 (O_1663,N_24932,N_24862);
xor UO_1664 (O_1664,N_24913,N_24836);
nand UO_1665 (O_1665,N_24981,N_24758);
nor UO_1666 (O_1666,N_24793,N_24860);
nor UO_1667 (O_1667,N_24762,N_24915);
nand UO_1668 (O_1668,N_24970,N_24759);
and UO_1669 (O_1669,N_24843,N_24849);
or UO_1670 (O_1670,N_24873,N_24786);
and UO_1671 (O_1671,N_24991,N_24928);
xnor UO_1672 (O_1672,N_24802,N_24927);
and UO_1673 (O_1673,N_24808,N_24820);
nor UO_1674 (O_1674,N_24958,N_24993);
or UO_1675 (O_1675,N_24986,N_24939);
nand UO_1676 (O_1676,N_24866,N_24954);
xor UO_1677 (O_1677,N_24871,N_24783);
or UO_1678 (O_1678,N_24948,N_24895);
and UO_1679 (O_1679,N_24960,N_24763);
nor UO_1680 (O_1680,N_24852,N_24863);
nand UO_1681 (O_1681,N_24866,N_24884);
nand UO_1682 (O_1682,N_24797,N_24961);
and UO_1683 (O_1683,N_24987,N_24833);
or UO_1684 (O_1684,N_24778,N_24868);
nor UO_1685 (O_1685,N_24895,N_24963);
or UO_1686 (O_1686,N_24921,N_24950);
nor UO_1687 (O_1687,N_24870,N_24856);
and UO_1688 (O_1688,N_24770,N_24936);
xor UO_1689 (O_1689,N_24776,N_24784);
nand UO_1690 (O_1690,N_24917,N_24765);
or UO_1691 (O_1691,N_24916,N_24992);
or UO_1692 (O_1692,N_24767,N_24948);
or UO_1693 (O_1693,N_24800,N_24788);
xnor UO_1694 (O_1694,N_24948,N_24790);
or UO_1695 (O_1695,N_24817,N_24965);
and UO_1696 (O_1696,N_24900,N_24766);
nand UO_1697 (O_1697,N_24922,N_24769);
xor UO_1698 (O_1698,N_24763,N_24884);
or UO_1699 (O_1699,N_24770,N_24945);
nand UO_1700 (O_1700,N_24959,N_24757);
xnor UO_1701 (O_1701,N_24796,N_24753);
nor UO_1702 (O_1702,N_24935,N_24812);
or UO_1703 (O_1703,N_24935,N_24863);
or UO_1704 (O_1704,N_24772,N_24921);
and UO_1705 (O_1705,N_24967,N_24886);
nand UO_1706 (O_1706,N_24934,N_24801);
nor UO_1707 (O_1707,N_24835,N_24802);
xor UO_1708 (O_1708,N_24791,N_24788);
or UO_1709 (O_1709,N_24838,N_24988);
or UO_1710 (O_1710,N_24831,N_24844);
nor UO_1711 (O_1711,N_24913,N_24775);
or UO_1712 (O_1712,N_24844,N_24943);
nand UO_1713 (O_1713,N_24776,N_24864);
nor UO_1714 (O_1714,N_24828,N_24789);
or UO_1715 (O_1715,N_24936,N_24849);
nor UO_1716 (O_1716,N_24802,N_24922);
nor UO_1717 (O_1717,N_24991,N_24762);
nand UO_1718 (O_1718,N_24851,N_24900);
or UO_1719 (O_1719,N_24872,N_24800);
and UO_1720 (O_1720,N_24790,N_24909);
and UO_1721 (O_1721,N_24984,N_24996);
and UO_1722 (O_1722,N_24951,N_24828);
xnor UO_1723 (O_1723,N_24904,N_24928);
or UO_1724 (O_1724,N_24933,N_24968);
and UO_1725 (O_1725,N_24806,N_24799);
or UO_1726 (O_1726,N_24775,N_24840);
and UO_1727 (O_1727,N_24966,N_24889);
xnor UO_1728 (O_1728,N_24958,N_24865);
nand UO_1729 (O_1729,N_24990,N_24800);
and UO_1730 (O_1730,N_24901,N_24874);
nor UO_1731 (O_1731,N_24892,N_24958);
xnor UO_1732 (O_1732,N_24995,N_24769);
nand UO_1733 (O_1733,N_24823,N_24832);
xor UO_1734 (O_1734,N_24881,N_24811);
xor UO_1735 (O_1735,N_24937,N_24964);
or UO_1736 (O_1736,N_24755,N_24960);
and UO_1737 (O_1737,N_24760,N_24842);
nand UO_1738 (O_1738,N_24967,N_24810);
and UO_1739 (O_1739,N_24878,N_24908);
and UO_1740 (O_1740,N_24783,N_24837);
or UO_1741 (O_1741,N_24870,N_24963);
and UO_1742 (O_1742,N_24866,N_24763);
and UO_1743 (O_1743,N_24804,N_24913);
or UO_1744 (O_1744,N_24994,N_24822);
or UO_1745 (O_1745,N_24960,N_24831);
and UO_1746 (O_1746,N_24864,N_24997);
or UO_1747 (O_1747,N_24753,N_24930);
and UO_1748 (O_1748,N_24828,N_24753);
and UO_1749 (O_1749,N_24981,N_24969);
xor UO_1750 (O_1750,N_24950,N_24859);
nor UO_1751 (O_1751,N_24962,N_24827);
or UO_1752 (O_1752,N_24868,N_24881);
or UO_1753 (O_1753,N_24865,N_24757);
xnor UO_1754 (O_1754,N_24855,N_24904);
nand UO_1755 (O_1755,N_24754,N_24966);
and UO_1756 (O_1756,N_24821,N_24880);
and UO_1757 (O_1757,N_24975,N_24936);
nor UO_1758 (O_1758,N_24888,N_24752);
or UO_1759 (O_1759,N_24795,N_24888);
nor UO_1760 (O_1760,N_24889,N_24935);
nand UO_1761 (O_1761,N_24999,N_24998);
xor UO_1762 (O_1762,N_24792,N_24751);
nand UO_1763 (O_1763,N_24939,N_24912);
xnor UO_1764 (O_1764,N_24805,N_24912);
or UO_1765 (O_1765,N_24850,N_24942);
nand UO_1766 (O_1766,N_24762,N_24902);
xnor UO_1767 (O_1767,N_24990,N_24872);
xor UO_1768 (O_1768,N_24926,N_24900);
nand UO_1769 (O_1769,N_24904,N_24944);
nand UO_1770 (O_1770,N_24773,N_24814);
nor UO_1771 (O_1771,N_24880,N_24972);
xnor UO_1772 (O_1772,N_24876,N_24939);
nor UO_1773 (O_1773,N_24777,N_24783);
xnor UO_1774 (O_1774,N_24795,N_24897);
xor UO_1775 (O_1775,N_24952,N_24881);
nand UO_1776 (O_1776,N_24757,N_24849);
xnor UO_1777 (O_1777,N_24910,N_24979);
or UO_1778 (O_1778,N_24856,N_24830);
and UO_1779 (O_1779,N_24940,N_24937);
nand UO_1780 (O_1780,N_24910,N_24805);
and UO_1781 (O_1781,N_24802,N_24836);
xor UO_1782 (O_1782,N_24822,N_24954);
nand UO_1783 (O_1783,N_24910,N_24981);
nor UO_1784 (O_1784,N_24851,N_24827);
nor UO_1785 (O_1785,N_24935,N_24846);
nor UO_1786 (O_1786,N_24851,N_24824);
or UO_1787 (O_1787,N_24860,N_24892);
or UO_1788 (O_1788,N_24806,N_24877);
and UO_1789 (O_1789,N_24763,N_24792);
and UO_1790 (O_1790,N_24868,N_24937);
nor UO_1791 (O_1791,N_24892,N_24952);
nor UO_1792 (O_1792,N_24881,N_24960);
or UO_1793 (O_1793,N_24819,N_24868);
and UO_1794 (O_1794,N_24978,N_24819);
nor UO_1795 (O_1795,N_24824,N_24889);
nor UO_1796 (O_1796,N_24827,N_24995);
nand UO_1797 (O_1797,N_24942,N_24790);
nor UO_1798 (O_1798,N_24919,N_24979);
nor UO_1799 (O_1799,N_24984,N_24841);
and UO_1800 (O_1800,N_24784,N_24892);
and UO_1801 (O_1801,N_24919,N_24755);
and UO_1802 (O_1802,N_24831,N_24789);
or UO_1803 (O_1803,N_24754,N_24973);
nor UO_1804 (O_1804,N_24861,N_24770);
nand UO_1805 (O_1805,N_24930,N_24931);
and UO_1806 (O_1806,N_24941,N_24984);
nor UO_1807 (O_1807,N_24860,N_24795);
and UO_1808 (O_1808,N_24893,N_24914);
nor UO_1809 (O_1809,N_24896,N_24970);
nor UO_1810 (O_1810,N_24752,N_24910);
nand UO_1811 (O_1811,N_24870,N_24948);
or UO_1812 (O_1812,N_24763,N_24804);
nand UO_1813 (O_1813,N_24762,N_24782);
nand UO_1814 (O_1814,N_24781,N_24869);
xor UO_1815 (O_1815,N_24822,N_24921);
nand UO_1816 (O_1816,N_24854,N_24871);
and UO_1817 (O_1817,N_24920,N_24819);
and UO_1818 (O_1818,N_24922,N_24782);
nor UO_1819 (O_1819,N_24807,N_24917);
nor UO_1820 (O_1820,N_24938,N_24772);
and UO_1821 (O_1821,N_24852,N_24756);
nand UO_1822 (O_1822,N_24956,N_24964);
and UO_1823 (O_1823,N_24919,N_24929);
nor UO_1824 (O_1824,N_24925,N_24827);
nor UO_1825 (O_1825,N_24767,N_24972);
xnor UO_1826 (O_1826,N_24777,N_24898);
or UO_1827 (O_1827,N_24910,N_24867);
nor UO_1828 (O_1828,N_24798,N_24792);
nor UO_1829 (O_1829,N_24946,N_24802);
xnor UO_1830 (O_1830,N_24858,N_24917);
xnor UO_1831 (O_1831,N_24922,N_24919);
nand UO_1832 (O_1832,N_24832,N_24885);
xnor UO_1833 (O_1833,N_24770,N_24949);
nand UO_1834 (O_1834,N_24896,N_24950);
or UO_1835 (O_1835,N_24967,N_24927);
nand UO_1836 (O_1836,N_24959,N_24986);
nand UO_1837 (O_1837,N_24899,N_24924);
nand UO_1838 (O_1838,N_24777,N_24959);
nor UO_1839 (O_1839,N_24913,N_24933);
and UO_1840 (O_1840,N_24768,N_24922);
nor UO_1841 (O_1841,N_24866,N_24915);
nor UO_1842 (O_1842,N_24853,N_24976);
nand UO_1843 (O_1843,N_24976,N_24839);
nand UO_1844 (O_1844,N_24998,N_24898);
nand UO_1845 (O_1845,N_24981,N_24757);
nand UO_1846 (O_1846,N_24935,N_24891);
and UO_1847 (O_1847,N_24974,N_24789);
or UO_1848 (O_1848,N_24968,N_24908);
nor UO_1849 (O_1849,N_24770,N_24892);
nand UO_1850 (O_1850,N_24895,N_24971);
or UO_1851 (O_1851,N_24881,N_24827);
xnor UO_1852 (O_1852,N_24947,N_24905);
xor UO_1853 (O_1853,N_24929,N_24977);
nor UO_1854 (O_1854,N_24891,N_24998);
xnor UO_1855 (O_1855,N_24809,N_24919);
nand UO_1856 (O_1856,N_24952,N_24756);
nor UO_1857 (O_1857,N_24885,N_24818);
xor UO_1858 (O_1858,N_24875,N_24941);
or UO_1859 (O_1859,N_24824,N_24845);
and UO_1860 (O_1860,N_24961,N_24963);
nand UO_1861 (O_1861,N_24858,N_24943);
nor UO_1862 (O_1862,N_24986,N_24922);
nand UO_1863 (O_1863,N_24771,N_24914);
or UO_1864 (O_1864,N_24799,N_24862);
xnor UO_1865 (O_1865,N_24837,N_24778);
nand UO_1866 (O_1866,N_24980,N_24788);
nand UO_1867 (O_1867,N_24807,N_24928);
nand UO_1868 (O_1868,N_24924,N_24778);
and UO_1869 (O_1869,N_24876,N_24805);
and UO_1870 (O_1870,N_24946,N_24850);
or UO_1871 (O_1871,N_24766,N_24887);
xor UO_1872 (O_1872,N_24796,N_24890);
or UO_1873 (O_1873,N_24782,N_24826);
nand UO_1874 (O_1874,N_24820,N_24879);
nand UO_1875 (O_1875,N_24916,N_24882);
xnor UO_1876 (O_1876,N_24858,N_24912);
or UO_1877 (O_1877,N_24932,N_24922);
or UO_1878 (O_1878,N_24911,N_24790);
xor UO_1879 (O_1879,N_24960,N_24819);
nand UO_1880 (O_1880,N_24769,N_24882);
or UO_1881 (O_1881,N_24835,N_24975);
nor UO_1882 (O_1882,N_24777,N_24788);
nand UO_1883 (O_1883,N_24915,N_24874);
nand UO_1884 (O_1884,N_24801,N_24948);
nand UO_1885 (O_1885,N_24950,N_24847);
nor UO_1886 (O_1886,N_24828,N_24792);
nor UO_1887 (O_1887,N_24829,N_24995);
nor UO_1888 (O_1888,N_24795,N_24807);
nor UO_1889 (O_1889,N_24820,N_24786);
nand UO_1890 (O_1890,N_24946,N_24824);
nand UO_1891 (O_1891,N_24784,N_24816);
nor UO_1892 (O_1892,N_24976,N_24815);
nand UO_1893 (O_1893,N_24848,N_24891);
xnor UO_1894 (O_1894,N_24813,N_24814);
or UO_1895 (O_1895,N_24862,N_24779);
xnor UO_1896 (O_1896,N_24960,N_24845);
and UO_1897 (O_1897,N_24847,N_24963);
xnor UO_1898 (O_1898,N_24790,N_24859);
nand UO_1899 (O_1899,N_24814,N_24945);
and UO_1900 (O_1900,N_24753,N_24777);
and UO_1901 (O_1901,N_24940,N_24829);
and UO_1902 (O_1902,N_24811,N_24841);
xnor UO_1903 (O_1903,N_24819,N_24842);
and UO_1904 (O_1904,N_24930,N_24807);
xor UO_1905 (O_1905,N_24852,N_24913);
or UO_1906 (O_1906,N_24791,N_24937);
xor UO_1907 (O_1907,N_24788,N_24887);
nand UO_1908 (O_1908,N_24886,N_24754);
nor UO_1909 (O_1909,N_24922,N_24794);
xor UO_1910 (O_1910,N_24766,N_24754);
or UO_1911 (O_1911,N_24882,N_24867);
nor UO_1912 (O_1912,N_24851,N_24985);
or UO_1913 (O_1913,N_24783,N_24903);
and UO_1914 (O_1914,N_24921,N_24968);
nor UO_1915 (O_1915,N_24891,N_24901);
or UO_1916 (O_1916,N_24845,N_24984);
nand UO_1917 (O_1917,N_24838,N_24845);
nor UO_1918 (O_1918,N_24814,N_24783);
nor UO_1919 (O_1919,N_24889,N_24887);
xor UO_1920 (O_1920,N_24789,N_24750);
nand UO_1921 (O_1921,N_24931,N_24807);
xor UO_1922 (O_1922,N_24897,N_24931);
or UO_1923 (O_1923,N_24927,N_24770);
nand UO_1924 (O_1924,N_24949,N_24881);
nor UO_1925 (O_1925,N_24888,N_24798);
nor UO_1926 (O_1926,N_24919,N_24841);
nand UO_1927 (O_1927,N_24933,N_24848);
nor UO_1928 (O_1928,N_24851,N_24866);
and UO_1929 (O_1929,N_24774,N_24793);
nand UO_1930 (O_1930,N_24773,N_24761);
and UO_1931 (O_1931,N_24867,N_24845);
and UO_1932 (O_1932,N_24836,N_24957);
or UO_1933 (O_1933,N_24891,N_24959);
nor UO_1934 (O_1934,N_24988,N_24997);
nor UO_1935 (O_1935,N_24820,N_24758);
and UO_1936 (O_1936,N_24958,N_24792);
and UO_1937 (O_1937,N_24866,N_24875);
nor UO_1938 (O_1938,N_24881,N_24824);
xnor UO_1939 (O_1939,N_24762,N_24823);
or UO_1940 (O_1940,N_24887,N_24914);
nand UO_1941 (O_1941,N_24980,N_24921);
or UO_1942 (O_1942,N_24816,N_24757);
and UO_1943 (O_1943,N_24942,N_24843);
nor UO_1944 (O_1944,N_24946,N_24750);
nor UO_1945 (O_1945,N_24984,N_24982);
nor UO_1946 (O_1946,N_24968,N_24750);
xnor UO_1947 (O_1947,N_24777,N_24874);
xor UO_1948 (O_1948,N_24956,N_24977);
nor UO_1949 (O_1949,N_24974,N_24932);
and UO_1950 (O_1950,N_24906,N_24803);
nor UO_1951 (O_1951,N_24790,N_24929);
nor UO_1952 (O_1952,N_24850,N_24961);
xor UO_1953 (O_1953,N_24773,N_24809);
and UO_1954 (O_1954,N_24961,N_24981);
or UO_1955 (O_1955,N_24930,N_24995);
and UO_1956 (O_1956,N_24992,N_24846);
nor UO_1957 (O_1957,N_24812,N_24810);
xnor UO_1958 (O_1958,N_24921,N_24918);
nor UO_1959 (O_1959,N_24854,N_24947);
and UO_1960 (O_1960,N_24807,N_24874);
xor UO_1961 (O_1961,N_24821,N_24805);
nor UO_1962 (O_1962,N_24957,N_24934);
xnor UO_1963 (O_1963,N_24793,N_24968);
or UO_1964 (O_1964,N_24985,N_24882);
nor UO_1965 (O_1965,N_24993,N_24863);
and UO_1966 (O_1966,N_24969,N_24839);
and UO_1967 (O_1967,N_24886,N_24938);
or UO_1968 (O_1968,N_24948,N_24820);
nor UO_1969 (O_1969,N_24948,N_24845);
nor UO_1970 (O_1970,N_24930,N_24842);
nor UO_1971 (O_1971,N_24881,N_24776);
or UO_1972 (O_1972,N_24948,N_24889);
and UO_1973 (O_1973,N_24793,N_24875);
and UO_1974 (O_1974,N_24771,N_24795);
or UO_1975 (O_1975,N_24943,N_24825);
xnor UO_1976 (O_1976,N_24859,N_24754);
xnor UO_1977 (O_1977,N_24885,N_24984);
nand UO_1978 (O_1978,N_24816,N_24930);
and UO_1979 (O_1979,N_24903,N_24816);
or UO_1980 (O_1980,N_24810,N_24920);
or UO_1981 (O_1981,N_24853,N_24941);
or UO_1982 (O_1982,N_24810,N_24796);
nand UO_1983 (O_1983,N_24814,N_24771);
and UO_1984 (O_1984,N_24810,N_24966);
xnor UO_1985 (O_1985,N_24930,N_24850);
xor UO_1986 (O_1986,N_24885,N_24778);
and UO_1987 (O_1987,N_24951,N_24817);
or UO_1988 (O_1988,N_24928,N_24911);
or UO_1989 (O_1989,N_24753,N_24827);
nand UO_1990 (O_1990,N_24868,N_24813);
nand UO_1991 (O_1991,N_24868,N_24830);
xor UO_1992 (O_1992,N_24869,N_24820);
and UO_1993 (O_1993,N_24845,N_24849);
and UO_1994 (O_1994,N_24801,N_24979);
or UO_1995 (O_1995,N_24956,N_24836);
xnor UO_1996 (O_1996,N_24816,N_24850);
nor UO_1997 (O_1997,N_24981,N_24844);
and UO_1998 (O_1998,N_24766,N_24847);
and UO_1999 (O_1999,N_24762,N_24907);
or UO_2000 (O_2000,N_24787,N_24920);
xor UO_2001 (O_2001,N_24866,N_24775);
nand UO_2002 (O_2002,N_24760,N_24762);
nand UO_2003 (O_2003,N_24944,N_24813);
xnor UO_2004 (O_2004,N_24812,N_24983);
xnor UO_2005 (O_2005,N_24860,N_24942);
or UO_2006 (O_2006,N_24962,N_24851);
xor UO_2007 (O_2007,N_24829,N_24959);
nor UO_2008 (O_2008,N_24897,N_24848);
nand UO_2009 (O_2009,N_24950,N_24787);
nor UO_2010 (O_2010,N_24810,N_24959);
xnor UO_2011 (O_2011,N_24817,N_24886);
nor UO_2012 (O_2012,N_24932,N_24854);
and UO_2013 (O_2013,N_24794,N_24991);
nand UO_2014 (O_2014,N_24755,N_24817);
and UO_2015 (O_2015,N_24920,N_24898);
nor UO_2016 (O_2016,N_24851,N_24820);
or UO_2017 (O_2017,N_24757,N_24925);
and UO_2018 (O_2018,N_24922,N_24834);
xnor UO_2019 (O_2019,N_24897,N_24831);
xor UO_2020 (O_2020,N_24751,N_24787);
xor UO_2021 (O_2021,N_24920,N_24860);
nand UO_2022 (O_2022,N_24861,N_24757);
and UO_2023 (O_2023,N_24766,N_24801);
nor UO_2024 (O_2024,N_24996,N_24810);
nor UO_2025 (O_2025,N_24751,N_24810);
and UO_2026 (O_2026,N_24767,N_24962);
and UO_2027 (O_2027,N_24948,N_24937);
nor UO_2028 (O_2028,N_24794,N_24884);
nand UO_2029 (O_2029,N_24975,N_24768);
nor UO_2030 (O_2030,N_24997,N_24981);
or UO_2031 (O_2031,N_24985,N_24968);
and UO_2032 (O_2032,N_24928,N_24831);
nand UO_2033 (O_2033,N_24922,N_24833);
and UO_2034 (O_2034,N_24843,N_24986);
nand UO_2035 (O_2035,N_24954,N_24872);
nand UO_2036 (O_2036,N_24905,N_24848);
and UO_2037 (O_2037,N_24797,N_24901);
nand UO_2038 (O_2038,N_24772,N_24820);
or UO_2039 (O_2039,N_24951,N_24757);
or UO_2040 (O_2040,N_24777,N_24826);
and UO_2041 (O_2041,N_24924,N_24888);
and UO_2042 (O_2042,N_24998,N_24868);
nor UO_2043 (O_2043,N_24836,N_24795);
xor UO_2044 (O_2044,N_24896,N_24850);
nor UO_2045 (O_2045,N_24893,N_24972);
nor UO_2046 (O_2046,N_24879,N_24956);
nand UO_2047 (O_2047,N_24913,N_24955);
nor UO_2048 (O_2048,N_24759,N_24965);
and UO_2049 (O_2049,N_24841,N_24924);
nor UO_2050 (O_2050,N_24837,N_24952);
or UO_2051 (O_2051,N_24955,N_24752);
nand UO_2052 (O_2052,N_24997,N_24799);
nand UO_2053 (O_2053,N_24999,N_24828);
or UO_2054 (O_2054,N_24967,N_24885);
xnor UO_2055 (O_2055,N_24907,N_24890);
or UO_2056 (O_2056,N_24915,N_24975);
or UO_2057 (O_2057,N_24859,N_24981);
and UO_2058 (O_2058,N_24779,N_24942);
nand UO_2059 (O_2059,N_24885,N_24938);
xnor UO_2060 (O_2060,N_24823,N_24942);
or UO_2061 (O_2061,N_24839,N_24950);
or UO_2062 (O_2062,N_24818,N_24848);
or UO_2063 (O_2063,N_24965,N_24837);
or UO_2064 (O_2064,N_24808,N_24875);
or UO_2065 (O_2065,N_24916,N_24758);
nand UO_2066 (O_2066,N_24930,N_24921);
xnor UO_2067 (O_2067,N_24923,N_24779);
xnor UO_2068 (O_2068,N_24868,N_24906);
nor UO_2069 (O_2069,N_24922,N_24933);
or UO_2070 (O_2070,N_24794,N_24775);
or UO_2071 (O_2071,N_24780,N_24764);
nor UO_2072 (O_2072,N_24754,N_24751);
xor UO_2073 (O_2073,N_24880,N_24760);
and UO_2074 (O_2074,N_24841,N_24843);
nor UO_2075 (O_2075,N_24942,N_24955);
xnor UO_2076 (O_2076,N_24961,N_24892);
and UO_2077 (O_2077,N_24778,N_24819);
nor UO_2078 (O_2078,N_24966,N_24995);
or UO_2079 (O_2079,N_24753,N_24996);
and UO_2080 (O_2080,N_24908,N_24814);
and UO_2081 (O_2081,N_24848,N_24899);
and UO_2082 (O_2082,N_24861,N_24799);
or UO_2083 (O_2083,N_24976,N_24988);
nor UO_2084 (O_2084,N_24772,N_24844);
nand UO_2085 (O_2085,N_24808,N_24755);
or UO_2086 (O_2086,N_24891,N_24952);
and UO_2087 (O_2087,N_24914,N_24950);
nor UO_2088 (O_2088,N_24872,N_24988);
nor UO_2089 (O_2089,N_24829,N_24815);
nor UO_2090 (O_2090,N_24937,N_24887);
xor UO_2091 (O_2091,N_24979,N_24770);
nand UO_2092 (O_2092,N_24830,N_24948);
xnor UO_2093 (O_2093,N_24855,N_24773);
nand UO_2094 (O_2094,N_24753,N_24820);
nor UO_2095 (O_2095,N_24988,N_24831);
or UO_2096 (O_2096,N_24967,N_24835);
nand UO_2097 (O_2097,N_24985,N_24951);
nand UO_2098 (O_2098,N_24813,N_24871);
or UO_2099 (O_2099,N_24864,N_24824);
xor UO_2100 (O_2100,N_24944,N_24857);
nand UO_2101 (O_2101,N_24859,N_24814);
nor UO_2102 (O_2102,N_24955,N_24817);
and UO_2103 (O_2103,N_24754,N_24926);
nand UO_2104 (O_2104,N_24829,N_24884);
xor UO_2105 (O_2105,N_24971,N_24825);
nand UO_2106 (O_2106,N_24765,N_24861);
nor UO_2107 (O_2107,N_24837,N_24895);
nor UO_2108 (O_2108,N_24983,N_24978);
nor UO_2109 (O_2109,N_24801,N_24810);
or UO_2110 (O_2110,N_24821,N_24828);
and UO_2111 (O_2111,N_24926,N_24940);
xnor UO_2112 (O_2112,N_24784,N_24822);
xnor UO_2113 (O_2113,N_24801,N_24758);
nand UO_2114 (O_2114,N_24975,N_24932);
nor UO_2115 (O_2115,N_24887,N_24838);
and UO_2116 (O_2116,N_24851,N_24996);
and UO_2117 (O_2117,N_24889,N_24822);
nor UO_2118 (O_2118,N_24920,N_24776);
nor UO_2119 (O_2119,N_24908,N_24791);
xnor UO_2120 (O_2120,N_24751,N_24758);
or UO_2121 (O_2121,N_24901,N_24854);
xnor UO_2122 (O_2122,N_24911,N_24785);
or UO_2123 (O_2123,N_24958,N_24757);
nor UO_2124 (O_2124,N_24949,N_24902);
nor UO_2125 (O_2125,N_24777,N_24945);
xnor UO_2126 (O_2126,N_24858,N_24868);
and UO_2127 (O_2127,N_24795,N_24933);
or UO_2128 (O_2128,N_24965,N_24851);
xor UO_2129 (O_2129,N_24793,N_24917);
nor UO_2130 (O_2130,N_24923,N_24802);
nand UO_2131 (O_2131,N_24750,N_24770);
and UO_2132 (O_2132,N_24829,N_24809);
and UO_2133 (O_2133,N_24844,N_24910);
and UO_2134 (O_2134,N_24903,N_24797);
and UO_2135 (O_2135,N_24853,N_24781);
and UO_2136 (O_2136,N_24929,N_24791);
and UO_2137 (O_2137,N_24792,N_24796);
or UO_2138 (O_2138,N_24831,N_24892);
nor UO_2139 (O_2139,N_24885,N_24882);
or UO_2140 (O_2140,N_24912,N_24955);
xnor UO_2141 (O_2141,N_24770,N_24913);
or UO_2142 (O_2142,N_24750,N_24869);
or UO_2143 (O_2143,N_24838,N_24813);
and UO_2144 (O_2144,N_24950,N_24862);
or UO_2145 (O_2145,N_24996,N_24819);
and UO_2146 (O_2146,N_24775,N_24884);
or UO_2147 (O_2147,N_24999,N_24853);
nor UO_2148 (O_2148,N_24981,N_24858);
xnor UO_2149 (O_2149,N_24811,N_24849);
and UO_2150 (O_2150,N_24902,N_24821);
nor UO_2151 (O_2151,N_24926,N_24951);
xor UO_2152 (O_2152,N_24892,N_24867);
and UO_2153 (O_2153,N_24971,N_24817);
or UO_2154 (O_2154,N_24787,N_24765);
nor UO_2155 (O_2155,N_24831,N_24863);
nor UO_2156 (O_2156,N_24975,N_24906);
and UO_2157 (O_2157,N_24754,N_24936);
xnor UO_2158 (O_2158,N_24860,N_24840);
or UO_2159 (O_2159,N_24866,N_24997);
xnor UO_2160 (O_2160,N_24905,N_24935);
or UO_2161 (O_2161,N_24884,N_24917);
and UO_2162 (O_2162,N_24846,N_24921);
and UO_2163 (O_2163,N_24821,N_24949);
nor UO_2164 (O_2164,N_24918,N_24894);
nor UO_2165 (O_2165,N_24861,N_24877);
and UO_2166 (O_2166,N_24922,N_24786);
nand UO_2167 (O_2167,N_24825,N_24864);
or UO_2168 (O_2168,N_24974,N_24804);
nor UO_2169 (O_2169,N_24908,N_24888);
or UO_2170 (O_2170,N_24860,N_24786);
xnor UO_2171 (O_2171,N_24913,N_24875);
xor UO_2172 (O_2172,N_24878,N_24907);
nand UO_2173 (O_2173,N_24794,N_24948);
nand UO_2174 (O_2174,N_24797,N_24960);
nor UO_2175 (O_2175,N_24993,N_24995);
or UO_2176 (O_2176,N_24945,N_24848);
nor UO_2177 (O_2177,N_24923,N_24837);
and UO_2178 (O_2178,N_24874,N_24859);
nand UO_2179 (O_2179,N_24977,N_24967);
or UO_2180 (O_2180,N_24902,N_24970);
and UO_2181 (O_2181,N_24770,N_24925);
or UO_2182 (O_2182,N_24780,N_24767);
or UO_2183 (O_2183,N_24993,N_24795);
xor UO_2184 (O_2184,N_24784,N_24894);
xor UO_2185 (O_2185,N_24755,N_24788);
and UO_2186 (O_2186,N_24819,N_24846);
or UO_2187 (O_2187,N_24786,N_24998);
nor UO_2188 (O_2188,N_24821,N_24775);
nand UO_2189 (O_2189,N_24907,N_24999);
xor UO_2190 (O_2190,N_24948,N_24791);
nor UO_2191 (O_2191,N_24894,N_24780);
nand UO_2192 (O_2192,N_24782,N_24948);
or UO_2193 (O_2193,N_24920,N_24827);
or UO_2194 (O_2194,N_24909,N_24971);
or UO_2195 (O_2195,N_24965,N_24968);
nand UO_2196 (O_2196,N_24951,N_24891);
nor UO_2197 (O_2197,N_24788,N_24918);
nand UO_2198 (O_2198,N_24870,N_24955);
xor UO_2199 (O_2199,N_24940,N_24953);
nor UO_2200 (O_2200,N_24793,N_24949);
or UO_2201 (O_2201,N_24807,N_24837);
xor UO_2202 (O_2202,N_24764,N_24805);
xnor UO_2203 (O_2203,N_24906,N_24860);
xnor UO_2204 (O_2204,N_24941,N_24813);
and UO_2205 (O_2205,N_24875,N_24939);
and UO_2206 (O_2206,N_24760,N_24941);
or UO_2207 (O_2207,N_24799,N_24762);
and UO_2208 (O_2208,N_24796,N_24825);
nor UO_2209 (O_2209,N_24915,N_24828);
nand UO_2210 (O_2210,N_24880,N_24848);
and UO_2211 (O_2211,N_24923,N_24904);
nor UO_2212 (O_2212,N_24828,N_24945);
xnor UO_2213 (O_2213,N_24867,N_24872);
nor UO_2214 (O_2214,N_24981,N_24856);
and UO_2215 (O_2215,N_24958,N_24808);
xnor UO_2216 (O_2216,N_24798,N_24980);
nor UO_2217 (O_2217,N_24981,N_24975);
nand UO_2218 (O_2218,N_24884,N_24933);
and UO_2219 (O_2219,N_24806,N_24866);
nor UO_2220 (O_2220,N_24831,N_24903);
or UO_2221 (O_2221,N_24927,N_24828);
xor UO_2222 (O_2222,N_24796,N_24882);
nand UO_2223 (O_2223,N_24882,N_24880);
or UO_2224 (O_2224,N_24839,N_24851);
nand UO_2225 (O_2225,N_24980,N_24926);
nor UO_2226 (O_2226,N_24972,N_24847);
nor UO_2227 (O_2227,N_24905,N_24856);
xor UO_2228 (O_2228,N_24976,N_24919);
and UO_2229 (O_2229,N_24835,N_24933);
or UO_2230 (O_2230,N_24795,N_24796);
or UO_2231 (O_2231,N_24942,N_24758);
or UO_2232 (O_2232,N_24922,N_24910);
or UO_2233 (O_2233,N_24996,N_24900);
xor UO_2234 (O_2234,N_24910,N_24754);
and UO_2235 (O_2235,N_24903,N_24895);
xor UO_2236 (O_2236,N_24829,N_24849);
nand UO_2237 (O_2237,N_24787,N_24911);
nor UO_2238 (O_2238,N_24990,N_24887);
xor UO_2239 (O_2239,N_24873,N_24766);
nor UO_2240 (O_2240,N_24764,N_24972);
nand UO_2241 (O_2241,N_24952,N_24871);
or UO_2242 (O_2242,N_24816,N_24906);
and UO_2243 (O_2243,N_24920,N_24797);
or UO_2244 (O_2244,N_24968,N_24924);
nor UO_2245 (O_2245,N_24918,N_24943);
xnor UO_2246 (O_2246,N_24947,N_24940);
or UO_2247 (O_2247,N_24844,N_24752);
and UO_2248 (O_2248,N_24990,N_24817);
and UO_2249 (O_2249,N_24910,N_24816);
and UO_2250 (O_2250,N_24955,N_24862);
nand UO_2251 (O_2251,N_24824,N_24985);
or UO_2252 (O_2252,N_24965,N_24895);
nor UO_2253 (O_2253,N_24895,N_24888);
and UO_2254 (O_2254,N_24995,N_24780);
and UO_2255 (O_2255,N_24787,N_24912);
or UO_2256 (O_2256,N_24859,N_24967);
or UO_2257 (O_2257,N_24900,N_24977);
and UO_2258 (O_2258,N_24757,N_24945);
and UO_2259 (O_2259,N_24923,N_24867);
or UO_2260 (O_2260,N_24935,N_24931);
or UO_2261 (O_2261,N_24993,N_24997);
or UO_2262 (O_2262,N_24844,N_24944);
nor UO_2263 (O_2263,N_24924,N_24825);
and UO_2264 (O_2264,N_24894,N_24973);
xnor UO_2265 (O_2265,N_24855,N_24956);
nand UO_2266 (O_2266,N_24921,N_24951);
and UO_2267 (O_2267,N_24785,N_24805);
nor UO_2268 (O_2268,N_24782,N_24967);
or UO_2269 (O_2269,N_24757,N_24991);
xnor UO_2270 (O_2270,N_24759,N_24767);
or UO_2271 (O_2271,N_24982,N_24763);
or UO_2272 (O_2272,N_24823,N_24871);
and UO_2273 (O_2273,N_24972,N_24843);
and UO_2274 (O_2274,N_24993,N_24802);
and UO_2275 (O_2275,N_24892,N_24844);
xnor UO_2276 (O_2276,N_24926,N_24850);
nor UO_2277 (O_2277,N_24964,N_24786);
nand UO_2278 (O_2278,N_24992,N_24847);
or UO_2279 (O_2279,N_24751,N_24912);
or UO_2280 (O_2280,N_24884,N_24830);
nand UO_2281 (O_2281,N_24831,N_24945);
nor UO_2282 (O_2282,N_24998,N_24968);
nand UO_2283 (O_2283,N_24753,N_24782);
and UO_2284 (O_2284,N_24819,N_24983);
xor UO_2285 (O_2285,N_24874,N_24891);
and UO_2286 (O_2286,N_24802,N_24930);
xnor UO_2287 (O_2287,N_24946,N_24905);
and UO_2288 (O_2288,N_24938,N_24832);
and UO_2289 (O_2289,N_24945,N_24872);
nor UO_2290 (O_2290,N_24988,N_24845);
or UO_2291 (O_2291,N_24974,N_24888);
or UO_2292 (O_2292,N_24948,N_24996);
nor UO_2293 (O_2293,N_24868,N_24860);
and UO_2294 (O_2294,N_24953,N_24825);
xnor UO_2295 (O_2295,N_24851,N_24979);
nor UO_2296 (O_2296,N_24990,N_24801);
nand UO_2297 (O_2297,N_24897,N_24774);
or UO_2298 (O_2298,N_24820,N_24821);
nand UO_2299 (O_2299,N_24890,N_24843);
xnor UO_2300 (O_2300,N_24788,N_24968);
xor UO_2301 (O_2301,N_24940,N_24875);
or UO_2302 (O_2302,N_24996,N_24905);
and UO_2303 (O_2303,N_24891,N_24965);
nor UO_2304 (O_2304,N_24811,N_24963);
or UO_2305 (O_2305,N_24751,N_24942);
or UO_2306 (O_2306,N_24870,N_24919);
or UO_2307 (O_2307,N_24947,N_24954);
and UO_2308 (O_2308,N_24911,N_24914);
or UO_2309 (O_2309,N_24783,N_24851);
xnor UO_2310 (O_2310,N_24836,N_24915);
or UO_2311 (O_2311,N_24940,N_24914);
or UO_2312 (O_2312,N_24846,N_24951);
nand UO_2313 (O_2313,N_24919,N_24918);
or UO_2314 (O_2314,N_24795,N_24822);
or UO_2315 (O_2315,N_24963,N_24965);
xnor UO_2316 (O_2316,N_24838,N_24849);
nand UO_2317 (O_2317,N_24862,N_24885);
and UO_2318 (O_2318,N_24926,N_24967);
or UO_2319 (O_2319,N_24846,N_24903);
and UO_2320 (O_2320,N_24870,N_24791);
nor UO_2321 (O_2321,N_24922,N_24912);
or UO_2322 (O_2322,N_24936,N_24787);
nor UO_2323 (O_2323,N_24953,N_24950);
and UO_2324 (O_2324,N_24843,N_24917);
xor UO_2325 (O_2325,N_24861,N_24873);
or UO_2326 (O_2326,N_24969,N_24989);
nor UO_2327 (O_2327,N_24807,N_24936);
or UO_2328 (O_2328,N_24899,N_24757);
nand UO_2329 (O_2329,N_24891,N_24977);
or UO_2330 (O_2330,N_24776,N_24916);
or UO_2331 (O_2331,N_24947,N_24919);
or UO_2332 (O_2332,N_24968,N_24936);
and UO_2333 (O_2333,N_24906,N_24853);
xnor UO_2334 (O_2334,N_24832,N_24798);
nand UO_2335 (O_2335,N_24948,N_24965);
xnor UO_2336 (O_2336,N_24811,N_24820);
xnor UO_2337 (O_2337,N_24894,N_24987);
or UO_2338 (O_2338,N_24928,N_24926);
or UO_2339 (O_2339,N_24752,N_24842);
xor UO_2340 (O_2340,N_24863,N_24959);
xor UO_2341 (O_2341,N_24807,N_24895);
and UO_2342 (O_2342,N_24841,N_24865);
nor UO_2343 (O_2343,N_24918,N_24806);
or UO_2344 (O_2344,N_24864,N_24880);
nor UO_2345 (O_2345,N_24873,N_24954);
nor UO_2346 (O_2346,N_24858,N_24975);
nor UO_2347 (O_2347,N_24900,N_24951);
nand UO_2348 (O_2348,N_24845,N_24815);
xor UO_2349 (O_2349,N_24807,N_24938);
nand UO_2350 (O_2350,N_24925,N_24861);
and UO_2351 (O_2351,N_24886,N_24896);
or UO_2352 (O_2352,N_24958,N_24953);
and UO_2353 (O_2353,N_24956,N_24790);
and UO_2354 (O_2354,N_24854,N_24840);
nor UO_2355 (O_2355,N_24789,N_24751);
and UO_2356 (O_2356,N_24849,N_24826);
or UO_2357 (O_2357,N_24874,N_24816);
xor UO_2358 (O_2358,N_24854,N_24821);
nor UO_2359 (O_2359,N_24840,N_24895);
nor UO_2360 (O_2360,N_24965,N_24823);
and UO_2361 (O_2361,N_24812,N_24910);
or UO_2362 (O_2362,N_24888,N_24844);
and UO_2363 (O_2363,N_24924,N_24931);
xnor UO_2364 (O_2364,N_24920,N_24839);
or UO_2365 (O_2365,N_24991,N_24834);
or UO_2366 (O_2366,N_24883,N_24886);
nand UO_2367 (O_2367,N_24852,N_24994);
xor UO_2368 (O_2368,N_24979,N_24912);
nand UO_2369 (O_2369,N_24755,N_24771);
xnor UO_2370 (O_2370,N_24821,N_24992);
xor UO_2371 (O_2371,N_24976,N_24781);
or UO_2372 (O_2372,N_24912,N_24826);
nand UO_2373 (O_2373,N_24871,N_24839);
xnor UO_2374 (O_2374,N_24858,N_24844);
nor UO_2375 (O_2375,N_24798,N_24996);
nor UO_2376 (O_2376,N_24812,N_24950);
or UO_2377 (O_2377,N_24791,N_24909);
xnor UO_2378 (O_2378,N_24822,N_24878);
or UO_2379 (O_2379,N_24775,N_24849);
and UO_2380 (O_2380,N_24759,N_24786);
nand UO_2381 (O_2381,N_24789,N_24794);
xnor UO_2382 (O_2382,N_24867,N_24940);
nand UO_2383 (O_2383,N_24992,N_24829);
nand UO_2384 (O_2384,N_24936,N_24886);
or UO_2385 (O_2385,N_24907,N_24829);
and UO_2386 (O_2386,N_24884,N_24761);
and UO_2387 (O_2387,N_24915,N_24765);
nor UO_2388 (O_2388,N_24867,N_24803);
and UO_2389 (O_2389,N_24752,N_24771);
and UO_2390 (O_2390,N_24790,N_24821);
and UO_2391 (O_2391,N_24968,N_24780);
and UO_2392 (O_2392,N_24976,N_24816);
and UO_2393 (O_2393,N_24772,N_24817);
or UO_2394 (O_2394,N_24772,N_24999);
xnor UO_2395 (O_2395,N_24890,N_24920);
or UO_2396 (O_2396,N_24760,N_24796);
or UO_2397 (O_2397,N_24868,N_24799);
and UO_2398 (O_2398,N_24947,N_24895);
and UO_2399 (O_2399,N_24996,N_24842);
or UO_2400 (O_2400,N_24889,N_24780);
nor UO_2401 (O_2401,N_24938,N_24934);
or UO_2402 (O_2402,N_24836,N_24863);
and UO_2403 (O_2403,N_24773,N_24869);
or UO_2404 (O_2404,N_24839,N_24909);
nand UO_2405 (O_2405,N_24980,N_24895);
nor UO_2406 (O_2406,N_24909,N_24989);
xnor UO_2407 (O_2407,N_24774,N_24810);
and UO_2408 (O_2408,N_24929,N_24777);
or UO_2409 (O_2409,N_24812,N_24908);
xnor UO_2410 (O_2410,N_24971,N_24752);
or UO_2411 (O_2411,N_24905,N_24901);
nor UO_2412 (O_2412,N_24994,N_24993);
nand UO_2413 (O_2413,N_24893,N_24995);
nor UO_2414 (O_2414,N_24969,N_24854);
and UO_2415 (O_2415,N_24932,N_24762);
nor UO_2416 (O_2416,N_24924,N_24920);
and UO_2417 (O_2417,N_24799,N_24781);
or UO_2418 (O_2418,N_24878,N_24988);
nor UO_2419 (O_2419,N_24878,N_24846);
nor UO_2420 (O_2420,N_24761,N_24866);
nand UO_2421 (O_2421,N_24801,N_24920);
nand UO_2422 (O_2422,N_24816,N_24801);
nor UO_2423 (O_2423,N_24867,N_24978);
nand UO_2424 (O_2424,N_24815,N_24778);
xnor UO_2425 (O_2425,N_24952,N_24853);
nand UO_2426 (O_2426,N_24783,N_24857);
xnor UO_2427 (O_2427,N_24819,N_24830);
nor UO_2428 (O_2428,N_24906,N_24866);
and UO_2429 (O_2429,N_24906,N_24985);
xor UO_2430 (O_2430,N_24959,N_24880);
nor UO_2431 (O_2431,N_24754,N_24955);
or UO_2432 (O_2432,N_24801,N_24850);
or UO_2433 (O_2433,N_24805,N_24880);
xor UO_2434 (O_2434,N_24872,N_24899);
xnor UO_2435 (O_2435,N_24952,N_24862);
xnor UO_2436 (O_2436,N_24798,N_24922);
nand UO_2437 (O_2437,N_24904,N_24794);
xor UO_2438 (O_2438,N_24761,N_24764);
nor UO_2439 (O_2439,N_24764,N_24866);
nor UO_2440 (O_2440,N_24809,N_24994);
xor UO_2441 (O_2441,N_24856,N_24789);
or UO_2442 (O_2442,N_24798,N_24855);
or UO_2443 (O_2443,N_24817,N_24885);
and UO_2444 (O_2444,N_24848,N_24752);
or UO_2445 (O_2445,N_24875,N_24956);
or UO_2446 (O_2446,N_24798,N_24990);
or UO_2447 (O_2447,N_24899,N_24867);
and UO_2448 (O_2448,N_24938,N_24881);
and UO_2449 (O_2449,N_24997,N_24829);
xor UO_2450 (O_2450,N_24905,N_24814);
and UO_2451 (O_2451,N_24804,N_24819);
and UO_2452 (O_2452,N_24900,N_24921);
xor UO_2453 (O_2453,N_24792,N_24760);
nor UO_2454 (O_2454,N_24794,N_24791);
and UO_2455 (O_2455,N_24865,N_24981);
nor UO_2456 (O_2456,N_24851,N_24987);
nand UO_2457 (O_2457,N_24768,N_24759);
nand UO_2458 (O_2458,N_24779,N_24759);
or UO_2459 (O_2459,N_24981,N_24820);
nor UO_2460 (O_2460,N_24841,N_24874);
and UO_2461 (O_2461,N_24863,N_24757);
nor UO_2462 (O_2462,N_24788,N_24891);
or UO_2463 (O_2463,N_24791,N_24808);
nor UO_2464 (O_2464,N_24939,N_24794);
or UO_2465 (O_2465,N_24820,N_24773);
nor UO_2466 (O_2466,N_24850,N_24887);
and UO_2467 (O_2467,N_24875,N_24828);
nand UO_2468 (O_2468,N_24993,N_24949);
and UO_2469 (O_2469,N_24750,N_24982);
xnor UO_2470 (O_2470,N_24779,N_24992);
or UO_2471 (O_2471,N_24817,N_24925);
nand UO_2472 (O_2472,N_24945,N_24970);
xor UO_2473 (O_2473,N_24933,N_24907);
or UO_2474 (O_2474,N_24912,N_24880);
nor UO_2475 (O_2475,N_24779,N_24979);
or UO_2476 (O_2476,N_24924,N_24773);
or UO_2477 (O_2477,N_24959,N_24927);
xnor UO_2478 (O_2478,N_24989,N_24906);
nor UO_2479 (O_2479,N_24795,N_24892);
and UO_2480 (O_2480,N_24781,N_24938);
or UO_2481 (O_2481,N_24812,N_24852);
nor UO_2482 (O_2482,N_24961,N_24905);
xor UO_2483 (O_2483,N_24854,N_24768);
xnor UO_2484 (O_2484,N_24848,N_24986);
or UO_2485 (O_2485,N_24846,N_24968);
and UO_2486 (O_2486,N_24937,N_24889);
nor UO_2487 (O_2487,N_24915,N_24824);
and UO_2488 (O_2488,N_24825,N_24756);
and UO_2489 (O_2489,N_24958,N_24810);
xnor UO_2490 (O_2490,N_24889,N_24840);
nand UO_2491 (O_2491,N_24860,N_24823);
nand UO_2492 (O_2492,N_24804,N_24793);
xor UO_2493 (O_2493,N_24813,N_24932);
xnor UO_2494 (O_2494,N_24823,N_24926);
nor UO_2495 (O_2495,N_24802,N_24863);
and UO_2496 (O_2496,N_24992,N_24987);
or UO_2497 (O_2497,N_24766,N_24811);
nand UO_2498 (O_2498,N_24792,N_24818);
and UO_2499 (O_2499,N_24878,N_24882);
nor UO_2500 (O_2500,N_24888,N_24840);
or UO_2501 (O_2501,N_24859,N_24956);
nand UO_2502 (O_2502,N_24809,N_24761);
nor UO_2503 (O_2503,N_24843,N_24987);
and UO_2504 (O_2504,N_24945,N_24843);
xor UO_2505 (O_2505,N_24881,N_24918);
nor UO_2506 (O_2506,N_24818,N_24879);
xor UO_2507 (O_2507,N_24852,N_24838);
nand UO_2508 (O_2508,N_24936,N_24836);
and UO_2509 (O_2509,N_24974,N_24951);
and UO_2510 (O_2510,N_24910,N_24840);
nand UO_2511 (O_2511,N_24907,N_24978);
xor UO_2512 (O_2512,N_24857,N_24759);
xor UO_2513 (O_2513,N_24841,N_24768);
or UO_2514 (O_2514,N_24829,N_24796);
nand UO_2515 (O_2515,N_24892,N_24758);
nand UO_2516 (O_2516,N_24838,N_24847);
and UO_2517 (O_2517,N_24924,N_24847);
and UO_2518 (O_2518,N_24894,N_24828);
nor UO_2519 (O_2519,N_24990,N_24775);
or UO_2520 (O_2520,N_24938,N_24763);
or UO_2521 (O_2521,N_24911,N_24828);
or UO_2522 (O_2522,N_24975,N_24803);
and UO_2523 (O_2523,N_24900,N_24777);
nand UO_2524 (O_2524,N_24961,N_24789);
nor UO_2525 (O_2525,N_24874,N_24768);
xnor UO_2526 (O_2526,N_24911,N_24966);
nor UO_2527 (O_2527,N_24947,N_24824);
and UO_2528 (O_2528,N_24849,N_24752);
xor UO_2529 (O_2529,N_24805,N_24857);
nand UO_2530 (O_2530,N_24775,N_24798);
xor UO_2531 (O_2531,N_24751,N_24852);
nand UO_2532 (O_2532,N_24813,N_24799);
xor UO_2533 (O_2533,N_24980,N_24775);
and UO_2534 (O_2534,N_24948,N_24910);
and UO_2535 (O_2535,N_24762,N_24923);
and UO_2536 (O_2536,N_24896,N_24798);
xnor UO_2537 (O_2537,N_24752,N_24917);
nand UO_2538 (O_2538,N_24873,N_24842);
or UO_2539 (O_2539,N_24825,N_24970);
xnor UO_2540 (O_2540,N_24937,N_24975);
xor UO_2541 (O_2541,N_24827,N_24802);
xnor UO_2542 (O_2542,N_24802,N_24983);
and UO_2543 (O_2543,N_24977,N_24819);
or UO_2544 (O_2544,N_24844,N_24996);
xnor UO_2545 (O_2545,N_24908,N_24761);
or UO_2546 (O_2546,N_24754,N_24951);
nand UO_2547 (O_2547,N_24902,N_24816);
and UO_2548 (O_2548,N_24859,N_24937);
or UO_2549 (O_2549,N_24867,N_24767);
and UO_2550 (O_2550,N_24944,N_24939);
or UO_2551 (O_2551,N_24889,N_24967);
nor UO_2552 (O_2552,N_24909,N_24793);
xnor UO_2553 (O_2553,N_24879,N_24859);
or UO_2554 (O_2554,N_24912,N_24909);
and UO_2555 (O_2555,N_24919,N_24990);
and UO_2556 (O_2556,N_24916,N_24915);
nor UO_2557 (O_2557,N_24785,N_24956);
nand UO_2558 (O_2558,N_24875,N_24769);
nand UO_2559 (O_2559,N_24758,N_24842);
and UO_2560 (O_2560,N_24871,N_24785);
nand UO_2561 (O_2561,N_24919,N_24771);
nor UO_2562 (O_2562,N_24995,N_24973);
xor UO_2563 (O_2563,N_24901,N_24903);
nor UO_2564 (O_2564,N_24799,N_24778);
nor UO_2565 (O_2565,N_24873,N_24769);
or UO_2566 (O_2566,N_24754,N_24807);
and UO_2567 (O_2567,N_24934,N_24787);
or UO_2568 (O_2568,N_24847,N_24785);
or UO_2569 (O_2569,N_24885,N_24937);
nand UO_2570 (O_2570,N_24950,N_24895);
and UO_2571 (O_2571,N_24893,N_24810);
or UO_2572 (O_2572,N_24751,N_24805);
nor UO_2573 (O_2573,N_24813,N_24840);
nand UO_2574 (O_2574,N_24882,N_24973);
nand UO_2575 (O_2575,N_24843,N_24804);
nand UO_2576 (O_2576,N_24825,N_24778);
and UO_2577 (O_2577,N_24981,N_24955);
or UO_2578 (O_2578,N_24889,N_24846);
or UO_2579 (O_2579,N_24899,N_24920);
and UO_2580 (O_2580,N_24929,N_24962);
xor UO_2581 (O_2581,N_24911,N_24922);
and UO_2582 (O_2582,N_24816,N_24937);
nor UO_2583 (O_2583,N_24801,N_24905);
nor UO_2584 (O_2584,N_24998,N_24906);
nor UO_2585 (O_2585,N_24873,N_24932);
and UO_2586 (O_2586,N_24970,N_24901);
and UO_2587 (O_2587,N_24936,N_24819);
nor UO_2588 (O_2588,N_24798,N_24865);
nand UO_2589 (O_2589,N_24971,N_24892);
xor UO_2590 (O_2590,N_24875,N_24973);
and UO_2591 (O_2591,N_24857,N_24863);
and UO_2592 (O_2592,N_24860,N_24757);
xnor UO_2593 (O_2593,N_24980,N_24959);
and UO_2594 (O_2594,N_24933,N_24904);
nand UO_2595 (O_2595,N_24751,N_24817);
and UO_2596 (O_2596,N_24891,N_24916);
or UO_2597 (O_2597,N_24901,N_24939);
xor UO_2598 (O_2598,N_24829,N_24939);
and UO_2599 (O_2599,N_24846,N_24915);
and UO_2600 (O_2600,N_24971,N_24925);
and UO_2601 (O_2601,N_24995,N_24862);
nand UO_2602 (O_2602,N_24891,N_24981);
xor UO_2603 (O_2603,N_24957,N_24986);
xnor UO_2604 (O_2604,N_24868,N_24935);
and UO_2605 (O_2605,N_24877,N_24884);
xnor UO_2606 (O_2606,N_24813,N_24885);
xnor UO_2607 (O_2607,N_24886,N_24913);
nand UO_2608 (O_2608,N_24872,N_24787);
nor UO_2609 (O_2609,N_24906,N_24795);
or UO_2610 (O_2610,N_24876,N_24808);
nand UO_2611 (O_2611,N_24816,N_24956);
nand UO_2612 (O_2612,N_24925,N_24750);
xnor UO_2613 (O_2613,N_24782,N_24941);
nor UO_2614 (O_2614,N_24891,N_24950);
or UO_2615 (O_2615,N_24830,N_24791);
and UO_2616 (O_2616,N_24885,N_24792);
or UO_2617 (O_2617,N_24880,N_24903);
or UO_2618 (O_2618,N_24910,N_24797);
and UO_2619 (O_2619,N_24788,N_24907);
xor UO_2620 (O_2620,N_24869,N_24813);
or UO_2621 (O_2621,N_24997,N_24885);
nand UO_2622 (O_2622,N_24966,N_24833);
xor UO_2623 (O_2623,N_24954,N_24786);
and UO_2624 (O_2624,N_24784,N_24981);
nor UO_2625 (O_2625,N_24958,N_24982);
and UO_2626 (O_2626,N_24864,N_24762);
nor UO_2627 (O_2627,N_24809,N_24848);
nor UO_2628 (O_2628,N_24819,N_24969);
xor UO_2629 (O_2629,N_24843,N_24921);
nand UO_2630 (O_2630,N_24915,N_24853);
and UO_2631 (O_2631,N_24938,N_24852);
and UO_2632 (O_2632,N_24794,N_24907);
or UO_2633 (O_2633,N_24755,N_24819);
or UO_2634 (O_2634,N_24815,N_24858);
or UO_2635 (O_2635,N_24817,N_24979);
nand UO_2636 (O_2636,N_24882,N_24934);
or UO_2637 (O_2637,N_24992,N_24986);
and UO_2638 (O_2638,N_24926,N_24848);
nand UO_2639 (O_2639,N_24938,N_24841);
and UO_2640 (O_2640,N_24786,N_24896);
nand UO_2641 (O_2641,N_24881,N_24966);
and UO_2642 (O_2642,N_24933,N_24854);
and UO_2643 (O_2643,N_24966,N_24885);
xor UO_2644 (O_2644,N_24893,N_24847);
nor UO_2645 (O_2645,N_24993,N_24887);
nor UO_2646 (O_2646,N_24759,N_24852);
xnor UO_2647 (O_2647,N_24956,N_24784);
or UO_2648 (O_2648,N_24974,N_24890);
xor UO_2649 (O_2649,N_24890,N_24908);
and UO_2650 (O_2650,N_24755,N_24840);
xor UO_2651 (O_2651,N_24910,N_24817);
or UO_2652 (O_2652,N_24777,N_24992);
nand UO_2653 (O_2653,N_24895,N_24763);
xor UO_2654 (O_2654,N_24843,N_24806);
xor UO_2655 (O_2655,N_24805,N_24943);
xor UO_2656 (O_2656,N_24888,N_24951);
nand UO_2657 (O_2657,N_24999,N_24780);
and UO_2658 (O_2658,N_24877,N_24999);
nand UO_2659 (O_2659,N_24934,N_24965);
nor UO_2660 (O_2660,N_24792,N_24863);
nand UO_2661 (O_2661,N_24952,N_24939);
and UO_2662 (O_2662,N_24946,N_24967);
xnor UO_2663 (O_2663,N_24847,N_24779);
or UO_2664 (O_2664,N_24842,N_24818);
xnor UO_2665 (O_2665,N_24891,N_24816);
nor UO_2666 (O_2666,N_24847,N_24864);
nand UO_2667 (O_2667,N_24858,N_24839);
xnor UO_2668 (O_2668,N_24853,N_24766);
nand UO_2669 (O_2669,N_24985,N_24929);
and UO_2670 (O_2670,N_24985,N_24865);
or UO_2671 (O_2671,N_24945,N_24913);
nand UO_2672 (O_2672,N_24877,N_24870);
or UO_2673 (O_2673,N_24950,N_24929);
nor UO_2674 (O_2674,N_24818,N_24834);
nor UO_2675 (O_2675,N_24885,N_24961);
nor UO_2676 (O_2676,N_24842,N_24962);
and UO_2677 (O_2677,N_24779,N_24770);
nand UO_2678 (O_2678,N_24975,N_24930);
or UO_2679 (O_2679,N_24806,N_24886);
xnor UO_2680 (O_2680,N_24756,N_24993);
nor UO_2681 (O_2681,N_24884,N_24809);
and UO_2682 (O_2682,N_24938,N_24942);
nand UO_2683 (O_2683,N_24825,N_24808);
xor UO_2684 (O_2684,N_24994,N_24967);
and UO_2685 (O_2685,N_24967,N_24961);
nor UO_2686 (O_2686,N_24794,N_24958);
or UO_2687 (O_2687,N_24974,N_24973);
xor UO_2688 (O_2688,N_24945,N_24850);
nand UO_2689 (O_2689,N_24842,N_24908);
nand UO_2690 (O_2690,N_24813,N_24786);
or UO_2691 (O_2691,N_24889,N_24797);
and UO_2692 (O_2692,N_24863,N_24869);
or UO_2693 (O_2693,N_24826,N_24750);
xnor UO_2694 (O_2694,N_24902,N_24990);
and UO_2695 (O_2695,N_24979,N_24942);
or UO_2696 (O_2696,N_24920,N_24830);
nand UO_2697 (O_2697,N_24958,N_24781);
or UO_2698 (O_2698,N_24750,N_24971);
nor UO_2699 (O_2699,N_24979,N_24773);
xnor UO_2700 (O_2700,N_24868,N_24957);
nor UO_2701 (O_2701,N_24910,N_24882);
nand UO_2702 (O_2702,N_24902,N_24952);
or UO_2703 (O_2703,N_24911,N_24756);
nor UO_2704 (O_2704,N_24901,N_24836);
or UO_2705 (O_2705,N_24812,N_24854);
nor UO_2706 (O_2706,N_24772,N_24928);
or UO_2707 (O_2707,N_24914,N_24800);
nand UO_2708 (O_2708,N_24974,N_24953);
nand UO_2709 (O_2709,N_24876,N_24811);
xnor UO_2710 (O_2710,N_24778,N_24970);
or UO_2711 (O_2711,N_24992,N_24761);
nor UO_2712 (O_2712,N_24970,N_24879);
or UO_2713 (O_2713,N_24776,N_24909);
nand UO_2714 (O_2714,N_24900,N_24853);
nand UO_2715 (O_2715,N_24900,N_24919);
or UO_2716 (O_2716,N_24963,N_24970);
or UO_2717 (O_2717,N_24942,N_24933);
nand UO_2718 (O_2718,N_24983,N_24818);
nor UO_2719 (O_2719,N_24963,N_24797);
and UO_2720 (O_2720,N_24843,N_24758);
nor UO_2721 (O_2721,N_24984,N_24800);
nor UO_2722 (O_2722,N_24946,N_24763);
nor UO_2723 (O_2723,N_24938,N_24862);
nand UO_2724 (O_2724,N_24960,N_24758);
nor UO_2725 (O_2725,N_24910,N_24938);
nand UO_2726 (O_2726,N_24917,N_24875);
or UO_2727 (O_2727,N_24981,N_24884);
xor UO_2728 (O_2728,N_24977,N_24840);
nand UO_2729 (O_2729,N_24916,N_24938);
nand UO_2730 (O_2730,N_24803,N_24785);
nand UO_2731 (O_2731,N_24863,N_24800);
nor UO_2732 (O_2732,N_24886,N_24848);
and UO_2733 (O_2733,N_24815,N_24861);
or UO_2734 (O_2734,N_24949,N_24954);
nand UO_2735 (O_2735,N_24921,N_24888);
and UO_2736 (O_2736,N_24979,N_24781);
nor UO_2737 (O_2737,N_24750,N_24757);
or UO_2738 (O_2738,N_24905,N_24914);
nand UO_2739 (O_2739,N_24833,N_24947);
and UO_2740 (O_2740,N_24864,N_24978);
or UO_2741 (O_2741,N_24904,N_24991);
nand UO_2742 (O_2742,N_24791,N_24793);
nand UO_2743 (O_2743,N_24892,N_24825);
or UO_2744 (O_2744,N_24836,N_24894);
and UO_2745 (O_2745,N_24976,N_24811);
and UO_2746 (O_2746,N_24795,N_24995);
nor UO_2747 (O_2747,N_24894,N_24854);
and UO_2748 (O_2748,N_24822,N_24839);
nor UO_2749 (O_2749,N_24970,N_24891);
nor UO_2750 (O_2750,N_24847,N_24904);
nor UO_2751 (O_2751,N_24983,N_24868);
and UO_2752 (O_2752,N_24818,N_24932);
and UO_2753 (O_2753,N_24975,N_24777);
nor UO_2754 (O_2754,N_24967,N_24854);
nor UO_2755 (O_2755,N_24776,N_24965);
and UO_2756 (O_2756,N_24887,N_24952);
and UO_2757 (O_2757,N_24996,N_24812);
or UO_2758 (O_2758,N_24971,N_24819);
or UO_2759 (O_2759,N_24874,N_24900);
xnor UO_2760 (O_2760,N_24895,N_24785);
or UO_2761 (O_2761,N_24847,N_24958);
nand UO_2762 (O_2762,N_24883,N_24764);
or UO_2763 (O_2763,N_24923,N_24861);
xor UO_2764 (O_2764,N_24891,N_24917);
or UO_2765 (O_2765,N_24866,N_24848);
nand UO_2766 (O_2766,N_24903,N_24906);
and UO_2767 (O_2767,N_24883,N_24908);
or UO_2768 (O_2768,N_24961,N_24770);
xnor UO_2769 (O_2769,N_24874,N_24790);
nand UO_2770 (O_2770,N_24992,N_24818);
nand UO_2771 (O_2771,N_24901,N_24922);
or UO_2772 (O_2772,N_24890,N_24760);
or UO_2773 (O_2773,N_24935,N_24804);
or UO_2774 (O_2774,N_24974,N_24972);
nor UO_2775 (O_2775,N_24810,N_24871);
and UO_2776 (O_2776,N_24860,N_24760);
and UO_2777 (O_2777,N_24846,N_24977);
or UO_2778 (O_2778,N_24811,N_24774);
nor UO_2779 (O_2779,N_24977,N_24775);
and UO_2780 (O_2780,N_24990,N_24869);
xor UO_2781 (O_2781,N_24857,N_24830);
xor UO_2782 (O_2782,N_24990,N_24848);
or UO_2783 (O_2783,N_24770,N_24773);
nand UO_2784 (O_2784,N_24799,N_24899);
or UO_2785 (O_2785,N_24918,N_24913);
nor UO_2786 (O_2786,N_24761,N_24926);
nor UO_2787 (O_2787,N_24850,N_24966);
xor UO_2788 (O_2788,N_24779,N_24976);
or UO_2789 (O_2789,N_24776,N_24765);
and UO_2790 (O_2790,N_24972,N_24990);
nor UO_2791 (O_2791,N_24848,N_24942);
nor UO_2792 (O_2792,N_24968,N_24916);
nand UO_2793 (O_2793,N_24926,N_24815);
xnor UO_2794 (O_2794,N_24821,N_24835);
nand UO_2795 (O_2795,N_24929,N_24942);
nor UO_2796 (O_2796,N_24776,N_24782);
and UO_2797 (O_2797,N_24770,N_24778);
and UO_2798 (O_2798,N_24995,N_24832);
or UO_2799 (O_2799,N_24916,N_24811);
xor UO_2800 (O_2800,N_24768,N_24962);
or UO_2801 (O_2801,N_24943,N_24788);
nor UO_2802 (O_2802,N_24786,N_24937);
or UO_2803 (O_2803,N_24938,N_24922);
nor UO_2804 (O_2804,N_24790,N_24774);
nor UO_2805 (O_2805,N_24819,N_24769);
nand UO_2806 (O_2806,N_24977,N_24955);
xor UO_2807 (O_2807,N_24973,N_24821);
and UO_2808 (O_2808,N_24855,N_24799);
nor UO_2809 (O_2809,N_24812,N_24963);
nand UO_2810 (O_2810,N_24853,N_24799);
or UO_2811 (O_2811,N_24899,N_24854);
xor UO_2812 (O_2812,N_24869,N_24902);
and UO_2813 (O_2813,N_24912,N_24967);
nand UO_2814 (O_2814,N_24765,N_24838);
nand UO_2815 (O_2815,N_24933,N_24847);
or UO_2816 (O_2816,N_24851,N_24768);
nor UO_2817 (O_2817,N_24991,N_24952);
nand UO_2818 (O_2818,N_24920,N_24750);
nor UO_2819 (O_2819,N_24755,N_24863);
and UO_2820 (O_2820,N_24764,N_24953);
and UO_2821 (O_2821,N_24897,N_24982);
xor UO_2822 (O_2822,N_24976,N_24751);
and UO_2823 (O_2823,N_24778,N_24953);
xor UO_2824 (O_2824,N_24999,N_24872);
or UO_2825 (O_2825,N_24918,N_24907);
nor UO_2826 (O_2826,N_24761,N_24948);
or UO_2827 (O_2827,N_24932,N_24895);
or UO_2828 (O_2828,N_24836,N_24759);
nand UO_2829 (O_2829,N_24928,N_24999);
nor UO_2830 (O_2830,N_24957,N_24795);
and UO_2831 (O_2831,N_24876,N_24772);
nand UO_2832 (O_2832,N_24918,N_24812);
nand UO_2833 (O_2833,N_24779,N_24989);
or UO_2834 (O_2834,N_24863,N_24999);
and UO_2835 (O_2835,N_24815,N_24801);
or UO_2836 (O_2836,N_24782,N_24824);
nand UO_2837 (O_2837,N_24888,N_24801);
and UO_2838 (O_2838,N_24899,N_24782);
and UO_2839 (O_2839,N_24979,N_24789);
or UO_2840 (O_2840,N_24956,N_24797);
or UO_2841 (O_2841,N_24885,N_24828);
or UO_2842 (O_2842,N_24894,N_24972);
and UO_2843 (O_2843,N_24774,N_24952);
and UO_2844 (O_2844,N_24779,N_24915);
nand UO_2845 (O_2845,N_24928,N_24769);
or UO_2846 (O_2846,N_24891,N_24839);
or UO_2847 (O_2847,N_24902,N_24857);
nor UO_2848 (O_2848,N_24901,N_24908);
or UO_2849 (O_2849,N_24843,N_24803);
xor UO_2850 (O_2850,N_24983,N_24915);
or UO_2851 (O_2851,N_24756,N_24822);
nand UO_2852 (O_2852,N_24802,N_24996);
nand UO_2853 (O_2853,N_24820,N_24848);
and UO_2854 (O_2854,N_24824,N_24941);
nor UO_2855 (O_2855,N_24898,N_24810);
nand UO_2856 (O_2856,N_24825,N_24812);
nor UO_2857 (O_2857,N_24818,N_24862);
and UO_2858 (O_2858,N_24854,N_24897);
or UO_2859 (O_2859,N_24935,N_24798);
or UO_2860 (O_2860,N_24941,N_24774);
nor UO_2861 (O_2861,N_24768,N_24757);
xnor UO_2862 (O_2862,N_24989,N_24770);
and UO_2863 (O_2863,N_24945,N_24826);
xnor UO_2864 (O_2864,N_24903,N_24790);
and UO_2865 (O_2865,N_24974,N_24879);
xnor UO_2866 (O_2866,N_24911,N_24780);
xor UO_2867 (O_2867,N_24850,N_24830);
and UO_2868 (O_2868,N_24860,N_24944);
and UO_2869 (O_2869,N_24926,N_24818);
nand UO_2870 (O_2870,N_24979,N_24902);
and UO_2871 (O_2871,N_24936,N_24812);
xnor UO_2872 (O_2872,N_24810,N_24887);
and UO_2873 (O_2873,N_24825,N_24800);
or UO_2874 (O_2874,N_24757,N_24774);
and UO_2875 (O_2875,N_24786,N_24955);
nand UO_2876 (O_2876,N_24762,N_24883);
nor UO_2877 (O_2877,N_24830,N_24924);
or UO_2878 (O_2878,N_24939,N_24825);
nand UO_2879 (O_2879,N_24981,N_24794);
nand UO_2880 (O_2880,N_24839,N_24860);
nor UO_2881 (O_2881,N_24798,N_24901);
and UO_2882 (O_2882,N_24786,N_24783);
nor UO_2883 (O_2883,N_24766,N_24826);
or UO_2884 (O_2884,N_24853,N_24965);
nor UO_2885 (O_2885,N_24962,N_24876);
nor UO_2886 (O_2886,N_24908,N_24933);
nor UO_2887 (O_2887,N_24992,N_24890);
and UO_2888 (O_2888,N_24846,N_24927);
nor UO_2889 (O_2889,N_24759,N_24983);
nand UO_2890 (O_2890,N_24894,N_24935);
and UO_2891 (O_2891,N_24988,N_24874);
and UO_2892 (O_2892,N_24780,N_24935);
nand UO_2893 (O_2893,N_24835,N_24999);
nor UO_2894 (O_2894,N_24801,N_24973);
nand UO_2895 (O_2895,N_24817,N_24915);
xnor UO_2896 (O_2896,N_24768,N_24987);
xor UO_2897 (O_2897,N_24967,N_24958);
xor UO_2898 (O_2898,N_24874,N_24943);
or UO_2899 (O_2899,N_24922,N_24859);
and UO_2900 (O_2900,N_24903,N_24784);
and UO_2901 (O_2901,N_24995,N_24986);
or UO_2902 (O_2902,N_24967,N_24863);
nor UO_2903 (O_2903,N_24901,N_24850);
or UO_2904 (O_2904,N_24804,N_24975);
or UO_2905 (O_2905,N_24979,N_24873);
xnor UO_2906 (O_2906,N_24943,N_24806);
nor UO_2907 (O_2907,N_24955,N_24976);
nor UO_2908 (O_2908,N_24983,N_24847);
xnor UO_2909 (O_2909,N_24927,N_24936);
and UO_2910 (O_2910,N_24937,N_24913);
nand UO_2911 (O_2911,N_24891,N_24797);
and UO_2912 (O_2912,N_24949,N_24955);
and UO_2913 (O_2913,N_24993,N_24915);
nand UO_2914 (O_2914,N_24776,N_24779);
or UO_2915 (O_2915,N_24753,N_24995);
and UO_2916 (O_2916,N_24989,N_24917);
or UO_2917 (O_2917,N_24961,N_24933);
nand UO_2918 (O_2918,N_24986,N_24821);
and UO_2919 (O_2919,N_24876,N_24856);
and UO_2920 (O_2920,N_24824,N_24933);
nand UO_2921 (O_2921,N_24882,N_24964);
or UO_2922 (O_2922,N_24996,N_24992);
nand UO_2923 (O_2923,N_24854,N_24912);
xnor UO_2924 (O_2924,N_24752,N_24956);
or UO_2925 (O_2925,N_24819,N_24897);
xnor UO_2926 (O_2926,N_24856,N_24802);
and UO_2927 (O_2927,N_24935,N_24821);
nor UO_2928 (O_2928,N_24979,N_24870);
nor UO_2929 (O_2929,N_24997,N_24887);
nor UO_2930 (O_2930,N_24867,N_24780);
or UO_2931 (O_2931,N_24764,N_24815);
nor UO_2932 (O_2932,N_24990,N_24804);
xor UO_2933 (O_2933,N_24889,N_24951);
xnor UO_2934 (O_2934,N_24760,N_24886);
and UO_2935 (O_2935,N_24999,N_24885);
or UO_2936 (O_2936,N_24991,N_24809);
nand UO_2937 (O_2937,N_24900,N_24809);
or UO_2938 (O_2938,N_24820,N_24798);
xnor UO_2939 (O_2939,N_24768,N_24845);
nand UO_2940 (O_2940,N_24994,N_24918);
nand UO_2941 (O_2941,N_24971,N_24967);
xor UO_2942 (O_2942,N_24830,N_24807);
nor UO_2943 (O_2943,N_24918,N_24932);
or UO_2944 (O_2944,N_24900,N_24914);
nand UO_2945 (O_2945,N_24824,N_24860);
xnor UO_2946 (O_2946,N_24841,N_24762);
or UO_2947 (O_2947,N_24897,N_24970);
nor UO_2948 (O_2948,N_24926,N_24979);
and UO_2949 (O_2949,N_24987,N_24757);
and UO_2950 (O_2950,N_24813,N_24824);
nor UO_2951 (O_2951,N_24940,N_24998);
xnor UO_2952 (O_2952,N_24894,N_24965);
nand UO_2953 (O_2953,N_24772,N_24836);
xor UO_2954 (O_2954,N_24791,N_24842);
nor UO_2955 (O_2955,N_24848,N_24958);
or UO_2956 (O_2956,N_24845,N_24851);
or UO_2957 (O_2957,N_24781,N_24757);
xnor UO_2958 (O_2958,N_24991,N_24867);
and UO_2959 (O_2959,N_24969,N_24956);
nor UO_2960 (O_2960,N_24894,N_24890);
nand UO_2961 (O_2961,N_24908,N_24877);
nand UO_2962 (O_2962,N_24781,N_24790);
nor UO_2963 (O_2963,N_24829,N_24851);
and UO_2964 (O_2964,N_24964,N_24970);
or UO_2965 (O_2965,N_24859,N_24979);
xor UO_2966 (O_2966,N_24905,N_24854);
xor UO_2967 (O_2967,N_24767,N_24829);
nor UO_2968 (O_2968,N_24988,N_24944);
or UO_2969 (O_2969,N_24804,N_24789);
nand UO_2970 (O_2970,N_24878,N_24839);
xor UO_2971 (O_2971,N_24878,N_24801);
xnor UO_2972 (O_2972,N_24977,N_24808);
xor UO_2973 (O_2973,N_24998,N_24803);
nor UO_2974 (O_2974,N_24894,N_24781);
or UO_2975 (O_2975,N_24943,N_24926);
xor UO_2976 (O_2976,N_24955,N_24796);
xor UO_2977 (O_2977,N_24974,N_24904);
xor UO_2978 (O_2978,N_24988,N_24945);
nor UO_2979 (O_2979,N_24996,N_24962);
xor UO_2980 (O_2980,N_24815,N_24819);
and UO_2981 (O_2981,N_24969,N_24901);
or UO_2982 (O_2982,N_24996,N_24861);
or UO_2983 (O_2983,N_24763,N_24873);
and UO_2984 (O_2984,N_24874,N_24815);
or UO_2985 (O_2985,N_24750,N_24965);
nor UO_2986 (O_2986,N_24763,N_24781);
and UO_2987 (O_2987,N_24767,N_24798);
xor UO_2988 (O_2988,N_24776,N_24888);
or UO_2989 (O_2989,N_24934,N_24958);
xnor UO_2990 (O_2990,N_24849,N_24840);
xor UO_2991 (O_2991,N_24856,N_24914);
and UO_2992 (O_2992,N_24875,N_24762);
nand UO_2993 (O_2993,N_24860,N_24947);
xor UO_2994 (O_2994,N_24920,N_24849);
nand UO_2995 (O_2995,N_24801,N_24919);
or UO_2996 (O_2996,N_24871,N_24945);
nand UO_2997 (O_2997,N_24976,N_24787);
and UO_2998 (O_2998,N_24853,N_24946);
nor UO_2999 (O_2999,N_24805,N_24995);
endmodule