module basic_2000_20000_2500_125_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
nor U0 (N_0,In_1371,In_668);
nor U1 (N_1,In_1580,In_1286);
and U2 (N_2,In_705,In_1213);
and U3 (N_3,In_1464,In_683);
nor U4 (N_4,In_731,In_717);
or U5 (N_5,In_52,In_579);
xnor U6 (N_6,In_1832,In_167);
nand U7 (N_7,In_1396,In_1664);
or U8 (N_8,In_1723,In_664);
xnor U9 (N_9,In_532,In_126);
or U10 (N_10,In_1555,In_736);
nand U11 (N_11,In_85,In_342);
xor U12 (N_12,In_985,In_1673);
nor U13 (N_13,In_135,In_442);
nor U14 (N_14,In_6,In_1403);
nor U15 (N_15,In_1692,In_1310);
or U16 (N_16,In_1769,In_1375);
or U17 (N_17,In_1005,In_124);
xor U18 (N_18,In_217,In_1646);
and U19 (N_19,In_339,In_1971);
and U20 (N_20,In_498,In_1461);
and U21 (N_21,In_114,In_1475);
nand U22 (N_22,In_318,In_346);
nand U23 (N_23,In_1495,In_604);
xnor U24 (N_24,In_1168,In_711);
nand U25 (N_25,In_1939,In_870);
nor U26 (N_26,In_1276,In_1428);
or U27 (N_27,In_1257,In_64);
or U28 (N_28,In_1037,In_443);
and U29 (N_29,In_1797,In_817);
nand U30 (N_30,In_207,In_1894);
nor U31 (N_31,In_280,In_239);
xnor U32 (N_32,In_480,In_1914);
and U33 (N_33,In_413,In_1424);
and U34 (N_34,In_1741,In_1415);
or U35 (N_35,In_1657,In_1849);
nor U36 (N_36,In_1576,In_1943);
and U37 (N_37,In_1185,In_1134);
nor U38 (N_38,In_1116,In_1566);
and U39 (N_39,In_1903,In_1637);
nor U40 (N_40,In_1110,In_1523);
and U41 (N_41,In_566,In_249);
nor U42 (N_42,In_1485,In_991);
nand U43 (N_43,In_208,In_308);
nor U44 (N_44,In_1680,In_1079);
or U45 (N_45,In_620,In_1545);
nor U46 (N_46,In_1395,In_1277);
or U47 (N_47,In_1742,In_1011);
or U48 (N_48,In_844,In_1450);
or U49 (N_49,In_891,In_1196);
and U50 (N_50,In_675,In_700);
xnor U51 (N_51,In_1798,In_1136);
or U52 (N_52,In_487,In_1574);
nor U53 (N_53,In_586,In_344);
nor U54 (N_54,In_868,In_1223);
or U55 (N_55,In_1006,In_984);
or U56 (N_56,In_440,In_655);
and U57 (N_57,In_1416,In_1844);
or U58 (N_58,In_1009,In_1447);
nor U59 (N_59,In_1719,In_990);
nor U60 (N_60,In_1345,In_1237);
nor U61 (N_61,In_1486,In_1766);
and U62 (N_62,In_1000,In_323);
xnor U63 (N_63,In_1459,In_80);
xor U64 (N_64,In_1833,In_352);
nand U65 (N_65,In_543,In_1306);
or U66 (N_66,In_219,In_631);
nand U67 (N_67,In_1996,In_1171);
or U68 (N_68,In_1437,In_1929);
xor U69 (N_69,In_1684,In_792);
nor U70 (N_70,In_1367,In_530);
or U71 (N_71,In_131,In_647);
and U72 (N_72,In_1122,In_523);
and U73 (N_73,In_120,In_1278);
nand U74 (N_74,In_1467,In_1270);
xnor U75 (N_75,In_1454,In_1720);
nor U76 (N_76,In_583,In_992);
xor U77 (N_77,In_889,In_1198);
and U78 (N_78,In_412,In_69);
nor U79 (N_79,In_835,In_1210);
nand U80 (N_80,In_646,In_10);
or U81 (N_81,In_634,In_836);
and U82 (N_82,In_1259,In_1757);
nor U83 (N_83,In_197,In_71);
nor U84 (N_84,In_842,In_355);
and U85 (N_85,In_685,In_658);
and U86 (N_86,In_1627,In_562);
nand U87 (N_87,In_1650,In_1814);
nand U88 (N_88,In_1466,In_534);
and U89 (N_89,In_1651,In_356);
nand U90 (N_90,In_1618,In_1392);
xnor U91 (N_91,In_1207,In_212);
xnor U92 (N_92,In_17,In_1826);
nand U93 (N_93,In_1224,In_1861);
xor U94 (N_94,In_1955,In_1750);
and U95 (N_95,In_1705,In_788);
and U96 (N_96,In_1228,In_1801);
xor U97 (N_97,In_964,In_1496);
and U98 (N_98,In_1544,In_89);
nor U99 (N_99,In_1183,In_773);
nor U100 (N_100,In_977,In_1529);
or U101 (N_101,In_353,In_527);
or U102 (N_102,In_814,In_1030);
nand U103 (N_103,In_1036,In_1928);
xnor U104 (N_104,In_1509,In_1101);
nor U105 (N_105,In_1262,In_234);
and U106 (N_106,In_614,In_1867);
and U107 (N_107,In_763,In_809);
and U108 (N_108,In_259,In_1951);
and U109 (N_109,In_591,In_84);
xnor U110 (N_110,In_1655,In_53);
and U111 (N_111,In_1084,In_472);
and U112 (N_112,In_419,In_1409);
xnor U113 (N_113,In_752,In_494);
nor U114 (N_114,In_365,In_1194);
nor U115 (N_115,In_260,In_1290);
or U116 (N_116,In_629,In_1080);
nand U117 (N_117,In_1166,In_1180);
xnor U118 (N_118,In_1942,In_1812);
xnor U119 (N_119,In_1209,In_1035);
nor U120 (N_120,In_423,In_361);
and U121 (N_121,In_1232,In_929);
or U122 (N_122,In_238,In_580);
or U123 (N_123,In_1714,In_32);
and U124 (N_124,In_1519,In_1791);
and U125 (N_125,In_1315,In_1019);
xnor U126 (N_126,In_971,In_1795);
or U127 (N_127,In_186,In_1156);
xor U128 (N_128,In_1104,In_316);
nand U129 (N_129,In_1799,In_1856);
nand U130 (N_130,In_248,In_1387);
nor U131 (N_131,In_903,In_741);
and U132 (N_132,In_254,In_267);
nand U133 (N_133,In_815,In_1350);
or U134 (N_134,In_163,In_1220);
nor U135 (N_135,In_1384,In_58);
nand U136 (N_136,In_188,In_347);
and U137 (N_137,In_1900,In_210);
and U138 (N_138,In_1755,In_1758);
or U139 (N_139,In_805,In_1267);
xnor U140 (N_140,In_1328,In_552);
nor U141 (N_141,In_1398,In_1953);
nand U142 (N_142,In_1091,In_1882);
nor U143 (N_143,In_1029,In_1457);
nor U144 (N_144,In_912,In_955);
nor U145 (N_145,In_682,In_1252);
or U146 (N_146,In_112,In_825);
or U147 (N_147,In_1568,In_886);
nand U148 (N_148,In_652,In_1640);
nand U149 (N_149,In_1600,In_688);
and U150 (N_150,In_1992,In_1821);
and U151 (N_151,In_1569,In_1050);
and U152 (N_152,In_690,In_625);
nor U153 (N_153,In_505,In_1558);
and U154 (N_154,In_1153,In_1634);
xor U155 (N_155,In_1608,In_432);
and U156 (N_156,In_187,In_1342);
or U157 (N_157,In_1690,In_483);
and U158 (N_158,In_345,In_831);
nand U159 (N_159,In_1417,In_203);
xnor U160 (N_160,In_1526,In_1253);
xnor U161 (N_161,In_1382,In_1700);
nor U162 (N_162,In_235,In_1060);
xor U163 (N_163,In_698,In_531);
and U164 (N_164,In_1984,In_1255);
nand U165 (N_165,In_1099,In_136);
and U166 (N_166,N_130,N_20);
or U167 (N_167,In_828,In_1560);
and U168 (N_168,In_1347,N_52);
nor U169 (N_169,In_1133,In_284);
or U170 (N_170,In_1385,In_981);
xnor U171 (N_171,In_1291,In_1279);
and U172 (N_172,In_1327,In_1747);
and U173 (N_173,In_1443,In_734);
xor U174 (N_174,N_124,In_1932);
nand U175 (N_175,In_165,In_1408);
xnor U176 (N_176,In_500,In_29);
nor U177 (N_177,N_63,N_43);
and U178 (N_178,In_27,In_781);
or U179 (N_179,In_1445,In_1884);
nand U180 (N_180,In_1704,In_38);
and U181 (N_181,In_1179,In_541);
and U182 (N_182,In_1314,In_528);
and U183 (N_183,In_1172,In_1685);
nor U184 (N_184,In_1689,In_771);
and U185 (N_185,In_143,In_947);
xnor U186 (N_186,In_876,In_75);
and U187 (N_187,In_1546,In_1192);
or U188 (N_188,In_1629,In_28);
and U189 (N_189,In_1404,N_45);
nand U190 (N_190,N_62,In_198);
or U191 (N_191,In_1025,In_1401);
xnor U192 (N_192,In_657,In_291);
nor U193 (N_193,In_776,In_1659);
nor U194 (N_194,In_1683,In_901);
nand U195 (N_195,In_1046,In_986);
or U196 (N_196,In_846,In_996);
xnor U197 (N_197,In_1112,In_1191);
and U198 (N_198,In_521,In_1373);
nor U199 (N_199,In_457,In_1610);
nand U200 (N_200,In_926,In_1121);
and U201 (N_201,N_65,In_160);
and U202 (N_202,In_348,N_67);
nor U203 (N_203,In_304,In_1938);
xnor U204 (N_204,In_1540,In_1376);
and U205 (N_205,In_1752,In_770);
xnor U206 (N_206,In_1227,In_1785);
or U207 (N_207,In_1377,In_1021);
nand U208 (N_208,In_415,In_1451);
nand U209 (N_209,In_1311,In_74);
or U210 (N_210,In_908,In_1432);
xor U211 (N_211,In_1425,In_1258);
or U212 (N_212,In_1743,In_1418);
and U213 (N_213,In_204,In_502);
nor U214 (N_214,In_1499,In_818);
and U215 (N_215,In_1937,In_1835);
nor U216 (N_216,In_290,In_1400);
or U217 (N_217,In_738,In_1118);
or U218 (N_218,In_41,In_1246);
nor U219 (N_219,In_594,In_713);
nand U220 (N_220,In_1599,In_507);
xor U221 (N_221,In_1587,In_686);
xnor U222 (N_222,In_7,In_1312);
nand U223 (N_223,In_837,In_904);
nand U224 (N_224,In_549,In_179);
nor U225 (N_225,In_748,In_1893);
nor U226 (N_226,In_1807,In_1729);
xnor U227 (N_227,In_1825,In_1819);
and U228 (N_228,In_601,In_1904);
and U229 (N_229,In_966,In_1567);
nand U230 (N_230,In_125,In_1910);
nand U231 (N_231,In_873,In_1359);
and U232 (N_232,In_938,In_1950);
or U233 (N_233,In_1675,In_1200);
nand U234 (N_234,In_1438,In_1779);
xnor U235 (N_235,N_114,In_696);
and U236 (N_236,In_1641,In_1193);
and U237 (N_237,In_571,In_1887);
nor U238 (N_238,In_599,In_1563);
nand U239 (N_239,In_1820,In_722);
nand U240 (N_240,In_57,In_728);
and U241 (N_241,In_1841,In_376);
or U242 (N_242,In_1883,In_1788);
xnor U243 (N_243,In_1872,In_1733);
or U244 (N_244,In_175,In_590);
nor U245 (N_245,In_8,In_1973);
and U246 (N_246,In_402,In_24);
xnor U247 (N_247,In_1615,In_1749);
nand U248 (N_248,In_956,In_1732);
nor U249 (N_249,In_1614,In_492);
or U250 (N_250,N_85,In_1589);
and U251 (N_251,In_1987,In_1525);
and U252 (N_252,In_890,In_1473);
nor U253 (N_253,In_1537,In_1947);
nand U254 (N_254,N_39,In_1762);
nor U255 (N_255,In_1578,In_649);
or U256 (N_256,In_182,In_1869);
nor U257 (N_257,In_439,In_1096);
nand U258 (N_258,N_96,In_1239);
nor U259 (N_259,In_1763,In_1522);
or U260 (N_260,In_1759,In_917);
or U261 (N_261,In_482,In_597);
nor U262 (N_262,In_1508,In_177);
or U263 (N_263,In_1031,In_123);
nand U264 (N_264,In_1727,In_1287);
nand U265 (N_265,In_1282,In_1840);
nor U266 (N_266,In_87,In_1500);
or U267 (N_267,In_1871,In_1140);
and U268 (N_268,In_1137,In_1977);
or U269 (N_269,In_906,In_1751);
or U270 (N_270,In_319,In_397);
nor U271 (N_271,In_303,In_384);
nor U272 (N_272,In_1803,In_1958);
and U273 (N_273,In_1058,N_53);
and U274 (N_274,In_1076,In_1549);
and U275 (N_275,In_758,In_1520);
nor U276 (N_276,In_169,In_377);
and U277 (N_277,In_1303,In_619);
nand U278 (N_278,In_542,In_1730);
and U279 (N_279,In_1502,In_875);
nor U280 (N_280,In_775,In_1721);
xor U281 (N_281,In_1383,In_669);
nand U282 (N_282,In_621,In_885);
xor U283 (N_283,In_1745,In_1585);
or U284 (N_284,In_372,In_301);
nor U285 (N_285,N_139,In_1712);
nor U286 (N_286,In_1235,In_1441);
nor U287 (N_287,N_78,In_764);
xor U288 (N_288,In_573,In_1483);
xnor U289 (N_289,In_1676,In_1083);
or U290 (N_290,In_745,In_272);
nor U291 (N_291,In_367,In_1022);
or U292 (N_292,In_407,In_1389);
xnor U293 (N_293,In_1123,In_178);
or U294 (N_294,In_1902,In_164);
or U295 (N_295,N_31,In_952);
xor U296 (N_296,In_1407,In_859);
xnor U297 (N_297,In_398,In_1241);
xnor U298 (N_298,In_477,N_84);
nor U299 (N_299,In_559,In_1211);
xor U300 (N_300,In_845,In_1911);
or U301 (N_301,In_663,In_1264);
xor U302 (N_302,In_335,In_1838);
nand U303 (N_303,In_834,In_242);
nand U304 (N_304,In_1980,In_1127);
or U305 (N_305,In_45,In_1125);
nand U306 (N_306,N_121,In_974);
and U307 (N_307,In_1666,In_183);
nor U308 (N_308,In_750,In_998);
xnor U309 (N_309,In_360,In_1628);
or U310 (N_310,In_1656,In_735);
or U311 (N_311,In_1085,In_216);
or U312 (N_312,In_1420,N_88);
nor U313 (N_313,N_0,In_1460);
or U314 (N_314,In_1013,In_1090);
nand U315 (N_315,In_1806,In_1711);
and U316 (N_316,In_1471,In_759);
and U317 (N_317,In_269,In_281);
and U318 (N_318,In_1419,In_1511);
xnor U319 (N_319,N_137,In_861);
nor U320 (N_320,N_249,In_1824);
or U321 (N_321,In_1452,N_206);
nand U322 (N_322,N_184,In_1594);
or U323 (N_323,In_1131,In_1301);
and U324 (N_324,N_160,In_603);
nor U325 (N_325,In_306,In_765);
or U326 (N_326,In_694,In_681);
and U327 (N_327,In_840,In_99);
nor U328 (N_328,In_462,In_1805);
nand U329 (N_329,In_1412,In_812);
and U330 (N_330,In_1190,In_435);
nor U331 (N_331,In_895,In_1271);
nor U332 (N_332,In_1935,In_1480);
nor U333 (N_333,In_157,In_1899);
xnor U334 (N_334,In_1098,In_1173);
or U335 (N_335,In_830,In_411);
or U336 (N_336,In_1957,In_756);
and U337 (N_337,N_296,In_670);
nor U338 (N_338,In_394,In_278);
xnor U339 (N_339,In_554,In_1870);
nor U340 (N_340,In_958,N_21);
nand U341 (N_341,N_236,N_74);
nor U342 (N_342,N_1,In_1591);
or U343 (N_343,In_1538,In_545);
xor U344 (N_344,In_1514,In_899);
nor U345 (N_345,In_1411,In_1064);
nor U346 (N_346,In_1768,In_105);
and U347 (N_347,In_915,In_379);
nor U348 (N_348,In_1571,In_980);
nand U349 (N_349,In_1790,N_37);
and U350 (N_350,In_790,In_779);
nor U351 (N_351,In_1669,In_1603);
and U352 (N_352,In_1912,In_1468);
or U353 (N_353,In_1949,N_105);
xor U354 (N_354,In_226,In_1517);
nor U355 (N_355,In_612,In_1570);
and U356 (N_356,In_1174,In_12);
and U357 (N_357,In_223,In_36);
and U358 (N_358,In_643,In_1107);
nor U359 (N_359,In_1708,In_218);
nand U360 (N_360,In_170,In_1434);
xor U361 (N_361,N_248,In_496);
xor U362 (N_362,In_1126,N_77);
and U363 (N_363,In_1897,N_165);
and U364 (N_364,In_720,N_220);
xnor U365 (N_365,In_1962,In_1256);
nand U366 (N_366,In_707,In_1736);
or U367 (N_367,In_1501,In_1081);
and U368 (N_368,N_232,In_1828);
xor U369 (N_369,In_921,N_309);
and U370 (N_370,In_13,In_277);
nand U371 (N_371,In_733,N_292);
and U372 (N_372,In_548,N_169);
or U373 (N_373,In_957,In_563);
and U374 (N_374,In_1782,In_326);
or U375 (N_375,In_894,N_280);
and U376 (N_376,In_1405,N_34);
or U377 (N_377,In_61,In_689);
nand U378 (N_378,In_626,In_475);
and U379 (N_379,In_727,In_328);
xor U380 (N_380,In_1744,In_1890);
or U381 (N_381,In_710,N_100);
and U382 (N_382,In_181,N_101);
nor U383 (N_383,In_168,In_536);
nand U384 (N_384,N_228,In_1611);
and U385 (N_385,N_97,N_59);
nand U386 (N_386,In_1638,In_409);
nor U387 (N_387,In_778,N_193);
nand U388 (N_388,N_271,N_4);
nand U389 (N_389,In_428,In_111);
nand U390 (N_390,In_486,In_162);
nand U391 (N_391,In_1691,In_715);
nand U392 (N_392,In_1320,N_219);
nor U393 (N_393,In_1850,In_749);
nand U394 (N_394,N_94,In_684);
nand U395 (N_395,In_330,In_1654);
nor U396 (N_396,In_877,In_1907);
nor U397 (N_397,In_1152,In_538);
nor U398 (N_398,In_431,In_940);
and U399 (N_399,In_196,N_201);
nor U400 (N_400,In_1049,N_128);
and U401 (N_401,In_334,In_1874);
nand U402 (N_402,In_1491,In_332);
or U403 (N_403,In_102,In_1699);
xor U404 (N_404,N_24,In_458);
or U405 (N_405,In_185,N_92);
nor U406 (N_406,In_1448,N_268);
xor U407 (N_407,N_56,In_1672);
nand U408 (N_408,In_1891,In_1386);
xor U409 (N_409,N_27,In_98);
nand U410 (N_410,In_240,N_125);
nor U411 (N_411,N_261,In_489);
nor U412 (N_412,In_515,In_1913);
or U413 (N_413,In_953,N_35);
nor U414 (N_414,In_1189,In_1696);
or U415 (N_415,In_121,In_307);
nor U416 (N_416,In_1658,In_116);
and U417 (N_417,In_1007,In_1598);
or U418 (N_418,In_247,In_905);
and U419 (N_419,In_1332,In_774);
xor U420 (N_420,In_1510,In_1145);
xor U421 (N_421,In_82,In_995);
and U422 (N_422,In_1800,In_233);
xor U423 (N_423,In_806,In_86);
nor U424 (N_424,In_576,In_518);
nand U425 (N_425,In_1026,In_882);
nor U426 (N_426,In_390,In_300);
nor U427 (N_427,N_115,In_1815);
xnor U428 (N_428,N_194,In_418);
or U429 (N_429,In_40,In_471);
or U430 (N_430,N_278,In_195);
and U431 (N_431,In_1878,In_1718);
nand U432 (N_432,In_292,N_235);
nor U433 (N_433,In_931,In_789);
nor U434 (N_434,In_127,In_1433);
nor U435 (N_435,In_1487,In_1507);
and U436 (N_436,In_424,In_656);
xnor U437 (N_437,In_288,N_54);
nand U438 (N_438,In_1039,In_925);
or U439 (N_439,In_1340,N_216);
nor U440 (N_440,N_302,N_138);
nor U441 (N_441,N_245,In_769);
or U442 (N_442,In_1868,N_264);
and U443 (N_443,In_1885,In_1349);
nor U444 (N_444,N_303,In_1094);
nor U445 (N_445,In_537,In_1505);
or U446 (N_446,In_936,In_1956);
nand U447 (N_447,In_960,In_678);
or U448 (N_448,In_1606,In_1015);
nor U449 (N_449,In_176,In_967);
nor U450 (N_450,N_226,In_90);
or U451 (N_451,In_1754,In_461);
xnor U452 (N_452,In_589,N_181);
nand U453 (N_453,In_628,In_627);
nand U454 (N_454,In_1709,N_233);
or U455 (N_455,N_269,In_1042);
and U456 (N_456,In_857,In_374);
nor U457 (N_457,In_21,In_37);
nor U458 (N_458,In_1681,In_810);
and U459 (N_459,In_385,In_1695);
nor U460 (N_460,N_266,In_172);
or U461 (N_461,In_585,In_1863);
nand U462 (N_462,N_150,In_92);
nor U463 (N_463,In_1698,In_56);
or U464 (N_464,In_1242,In_1921);
or U465 (N_465,In_1177,N_11);
or U466 (N_466,In_119,In_1170);
and U467 (N_467,In_466,In_1045);
xor U468 (N_468,In_1852,In_595);
or U469 (N_469,In_732,In_30);
xnor U470 (N_470,N_319,In_1143);
nand U471 (N_471,In_1249,In_1933);
and U472 (N_472,In_555,In_305);
nor U473 (N_473,N_301,N_277);
or U474 (N_474,In_1061,In_1206);
nand U475 (N_475,In_1901,N_32);
or U476 (N_476,In_874,In_110);
or U477 (N_477,In_211,In_975);
nand U478 (N_478,In_1740,In_130);
nor U479 (N_479,In_222,In_1369);
nand U480 (N_480,N_472,In_946);
nor U481 (N_481,In_618,In_1186);
xnor U482 (N_482,N_287,In_1338);
and U483 (N_483,In_1917,N_87);
or U484 (N_484,In_31,In_315);
and U485 (N_485,In_1679,In_645);
and U486 (N_486,In_1023,N_200);
or U487 (N_487,In_1506,N_13);
nand U488 (N_488,In_1364,In_525);
xnor U489 (N_489,In_386,In_693);
or U490 (N_490,In_404,N_282);
nor U491 (N_491,In_753,In_979);
or U492 (N_492,In_1086,In_950);
or U493 (N_493,In_109,In_0);
and U494 (N_494,In_1588,In_1151);
xor U495 (N_495,In_73,In_863);
nor U496 (N_496,In_285,In_616);
xnor U497 (N_497,In_526,In_1216);
xnor U498 (N_498,In_1248,In_1251);
and U499 (N_499,In_1573,In_529);
xnor U500 (N_500,N_381,N_279);
xnor U501 (N_501,In_1556,In_481);
xor U502 (N_502,N_391,N_119);
or U503 (N_503,In_871,N_444);
nor U504 (N_504,In_1613,N_393);
and U505 (N_505,N_224,In_854);
nor U506 (N_506,In_1830,In_448);
and U507 (N_507,In_128,In_839);
and U508 (N_508,In_1339,In_144);
or U509 (N_509,In_644,N_8);
xnor U510 (N_510,N_196,N_172);
nand U511 (N_511,In_302,In_46);
or U512 (N_512,N_283,In_1786);
or U513 (N_513,N_338,In_230);
nor U514 (N_514,In_671,N_255);
nand U515 (N_515,In_1296,In_1427);
nand U516 (N_516,N_46,In_67);
nand U517 (N_517,In_1226,N_382);
or U518 (N_518,N_149,In_460);
xnor U519 (N_519,In_287,In_1582);
nand U520 (N_520,N_26,In_610);
or U521 (N_521,In_363,N_211);
xor U522 (N_522,In_1490,In_797);
and U523 (N_523,In_1357,In_1717);
and U524 (N_524,In_375,N_439);
nor U525 (N_525,In_1372,In_772);
nand U526 (N_526,In_1020,In_1584);
nand U527 (N_527,In_1968,N_234);
nor U528 (N_528,In_399,In_1682);
xnor U529 (N_529,In_615,In_1034);
and U530 (N_530,N_373,In_1041);
or U531 (N_531,In_336,In_1051);
xor U532 (N_532,In_1358,In_142);
or U533 (N_533,N_461,N_422);
xnor U534 (N_534,In_706,N_6);
nor U535 (N_535,N_142,N_449);
nand U536 (N_536,N_240,N_229);
or U537 (N_537,In_427,In_1920);
xor U538 (N_538,In_298,In_148);
or U539 (N_539,N_436,N_348);
nand U540 (N_540,In_1108,N_244);
nor U541 (N_541,In_994,In_1972);
nand U542 (N_542,In_1952,In_171);
xor U543 (N_543,In_426,N_346);
nand U544 (N_544,In_641,In_286);
or U545 (N_545,In_1756,In_1843);
and U546 (N_546,N_420,N_102);
or U547 (N_547,In_730,In_1111);
xnor U548 (N_548,N_202,In_550);
and U549 (N_549,In_1138,In_244);
xnor U550 (N_550,In_762,In_1150);
nand U551 (N_551,In_329,In_572);
nor U552 (N_552,In_1355,N_425);
xor U553 (N_553,In_1713,In_1981);
xor U554 (N_554,In_864,In_941);
nor U555 (N_555,N_259,In_1266);
xnor U556 (N_556,N_286,In_237);
nand U557 (N_557,In_847,In_463);
nor U558 (N_558,In_1990,In_495);
or U559 (N_559,N_49,In_1631);
nor U560 (N_560,In_703,In_1074);
and U561 (N_561,In_91,In_271);
and U562 (N_562,In_506,In_1289);
xor U563 (N_563,In_147,N_12);
or U564 (N_564,N_429,In_253);
nor U565 (N_565,N_431,N_392);
or U566 (N_566,In_565,In_295);
or U567 (N_567,In_1204,In_1132);
xnor U568 (N_568,In_1157,In_1866);
nor U569 (N_569,N_71,In_209);
xor U570 (N_570,In_1965,N_344);
and U571 (N_571,N_183,In_1668);
nand U572 (N_572,N_458,In_246);
nor U573 (N_573,In_1208,In_1865);
nand U574 (N_574,In_1836,N_366);
xor U575 (N_575,In_1100,In_1619);
nand U576 (N_576,In_1536,In_1528);
and U577 (N_577,In_808,N_3);
nand U578 (N_578,N_325,In_1504);
nor U579 (N_579,In_1834,In_1429);
or U580 (N_580,In_1141,In_948);
xnor U581 (N_581,In_1961,N_446);
xor U582 (N_582,In_1653,In_1954);
nand U583 (N_583,In_1781,In_129);
or U584 (N_584,N_270,N_129);
nand U585 (N_585,In_744,In_76);
and U586 (N_586,In_932,N_199);
xnor U587 (N_587,In_934,In_1738);
or U588 (N_588,In_1353,In_1829);
nand U589 (N_589,In_1097,In_1272);
nor U590 (N_590,In_416,N_146);
or U591 (N_591,N_433,In_1772);
nor U592 (N_592,In_1304,In_132);
nor U593 (N_593,N_17,In_910);
nor U594 (N_594,In_1557,N_442);
nand U595 (N_595,In_933,In_893);
and U596 (N_596,In_920,N_267);
or U597 (N_597,N_157,N_51);
and U598 (N_598,N_463,In_161);
nor U599 (N_599,In_1979,In_1380);
and U600 (N_600,In_1859,In_63);
nand U601 (N_601,In_1710,In_1813);
nand U602 (N_602,In_503,In_1916);
or U603 (N_603,N_343,In_1793);
and U604 (N_604,In_1877,In_1406);
nor U605 (N_605,In_1077,In_373);
nand U606 (N_606,In_189,In_635);
nor U607 (N_607,In_354,In_1985);
nand U608 (N_608,In_1970,In_473);
nor U609 (N_609,N_411,In_867);
or U610 (N_610,N_210,In_1356);
or U611 (N_611,In_1624,In_987);
nand U612 (N_612,N_400,N_322);
xor U613 (N_613,N_155,N_222);
and U614 (N_614,In_1817,In_62);
xnor U615 (N_615,In_252,In_16);
nor U616 (N_616,In_2,In_575);
nand U617 (N_617,In_767,In_802);
nor U618 (N_618,N_154,In_1784);
nor U619 (N_619,In_1661,In_1321);
nor U620 (N_620,In_725,In_1465);
or U621 (N_621,In_1048,In_632);
xnor U622 (N_622,In_1930,In_1188);
nor U623 (N_623,In_1532,In_1161);
xor U624 (N_624,In_659,In_746);
and U625 (N_625,In_1998,In_1374);
nor U626 (N_626,N_133,In_103);
nand U627 (N_627,In_1823,In_1966);
or U628 (N_628,In_1593,In_245);
or U629 (N_629,In_999,N_362);
xor U630 (N_630,N_151,In_520);
nor U631 (N_631,N_247,In_1853);
nor U632 (N_632,In_1012,In_1018);
or U633 (N_633,N_258,N_246);
nand U634 (N_634,In_1999,In_508);
nand U635 (N_635,In_1787,In_596);
nand U636 (N_636,In_721,In_517);
xnor U637 (N_637,N_300,In_1789);
and U638 (N_638,In_137,In_451);
nand U639 (N_639,In_1534,N_23);
xnor U640 (N_640,In_872,In_570);
nor U641 (N_641,N_437,N_495);
and U642 (N_642,In_1446,N_298);
or U643 (N_643,In_1044,In_1426);
and U644 (N_644,In_228,In_567);
nand U645 (N_645,N_47,In_97);
xnor U646 (N_646,In_609,N_498);
or U647 (N_647,N_380,N_89);
nand U648 (N_648,N_90,N_19);
nand U649 (N_649,N_5,In_973);
nor U650 (N_650,In_1215,In_1212);
nor U651 (N_651,In_1530,In_1731);
nand U652 (N_652,N_487,N_383);
or U653 (N_653,In_268,In_1335);
or U654 (N_654,In_70,N_600);
xnor U655 (N_655,N_186,N_48);
xnor U656 (N_656,In_184,In_1295);
nor U657 (N_657,In_1363,In_1440);
and U658 (N_658,N_409,N_104);
or U659 (N_659,In_1105,N_541);
or U660 (N_660,In_1305,In_799);
and U661 (N_661,N_311,N_326);
xnor U662 (N_662,In_1735,In_851);
xor U663 (N_663,In_742,In_1344);
xor U664 (N_664,In_1609,In_1182);
or U665 (N_665,N_132,In_944);
and U666 (N_666,In_968,N_76);
and U667 (N_667,In_1503,N_511);
and U668 (N_668,In_1366,N_335);
or U669 (N_669,In_553,In_833);
xor U670 (N_670,N_636,N_441);
xnor U671 (N_671,In_916,In_1095);
and U672 (N_672,In_918,In_606);
nand U673 (N_673,N_453,N_118);
or U674 (N_674,In_1895,In_1547);
xnor U675 (N_675,In_1994,In_314);
nand U676 (N_676,In_1436,N_2);
or U677 (N_677,In_1767,In_350);
nand U678 (N_678,N_95,In_1028);
xor U679 (N_679,In_602,In_154);
and U680 (N_680,In_650,N_83);
nand U681 (N_681,N_106,In_743);
xnor U682 (N_682,N_605,N_447);
nand U683 (N_683,In_1293,In_1792);
and U684 (N_684,In_898,In_937);
nand U685 (N_685,In_965,N_615);
nand U686 (N_686,In_1284,In_491);
nand U687 (N_687,N_469,In_478);
nand U688 (N_688,N_624,N_550);
and U689 (N_689,N_445,In_1038);
xnor U690 (N_690,In_983,N_73);
nand U691 (N_691,In_1178,N_408);
nor U692 (N_692,In_1146,N_179);
nor U693 (N_693,N_403,In_761);
or U694 (N_694,In_333,N_508);
nand U695 (N_695,In_1113,N_412);
nor U696 (N_696,In_383,In_194);
nand U697 (N_697,In_1351,In_1088);
or U698 (N_698,N_520,N_599);
xnor U699 (N_699,In_159,N_398);
xor U700 (N_700,N_460,In_1082);
nand U701 (N_701,N_33,In_438);
and U702 (N_702,In_1326,N_215);
and U703 (N_703,In_1581,In_214);
nor U704 (N_704,N_273,N_378);
nand U705 (N_705,N_521,In_737);
or U706 (N_706,N_333,In_106);
xor U707 (N_707,In_115,N_170);
xnor U708 (N_708,In_1810,In_878);
nand U709 (N_709,In_139,In_850);
nand U710 (N_710,In_909,In_648);
and U711 (N_711,In_1746,In_716);
nand U712 (N_712,N_103,N_355);
nor U713 (N_713,N_450,In_3);
xor U714 (N_714,N_167,N_585);
and U715 (N_715,In_569,In_1670);
and U716 (N_716,N_620,In_900);
nand U717 (N_717,N_597,In_803);
nor U718 (N_718,In_1936,In_444);
and U719 (N_719,N_416,In_1541);
nand U720 (N_720,In_540,In_1169);
nor U721 (N_721,In_270,In_55);
nor U722 (N_722,N_543,In_832);
or U723 (N_723,N_361,In_77);
or U724 (N_724,N_581,In_49);
or U725 (N_725,In_1488,In_1089);
nand U726 (N_726,In_1783,In_1275);
nand U727 (N_727,N_134,N_263);
or U728 (N_728,N_590,In_785);
nor U729 (N_729,In_1163,In_782);
or U730 (N_730,In_454,In_841);
nand U731 (N_731,In_1626,N_38);
nor U732 (N_732,N_257,In_1552);
xor U733 (N_733,N_528,N_432);
xor U734 (N_734,In_1273,In_1621);
and U735 (N_735,In_838,In_1822);
nor U736 (N_736,In_823,In_5);
nand U737 (N_737,In_1167,In_949);
nor U738 (N_738,In_317,N_285);
xor U739 (N_739,In_1201,In_1453);
nor U740 (N_740,In_1231,In_568);
nand U741 (N_741,N_136,N_58);
nand U742 (N_742,In_1765,In_257);
nand U743 (N_743,In_1093,In_429);
nand U744 (N_744,N_388,In_1632);
and U745 (N_745,N_152,N_345);
nor U746 (N_746,In_1413,N_284);
xnor U747 (N_747,In_1991,N_140);
nor U748 (N_748,In_1652,N_175);
nand U749 (N_749,In_1431,In_450);
nor U750 (N_750,In_989,N_608);
xor U751 (N_751,N_518,In_250);
or U752 (N_752,In_1724,N_616);
or U753 (N_753,In_997,N_327);
nor U754 (N_754,In_988,In_22);
xnor U755 (N_755,In_1770,N_542);
or U756 (N_756,In_816,In_642);
and U757 (N_757,N_162,In_1639);
or U758 (N_758,N_482,In_400);
nand U759 (N_759,In_624,N_353);
xnor U760 (N_760,In_1017,N_221);
nand U761 (N_761,N_504,In_1362);
xor U762 (N_762,In_1254,N_93);
and U763 (N_763,In_1230,In_1325);
nand U764 (N_764,In_1864,In_1737);
nand U765 (N_765,N_471,N_253);
nand U766 (N_766,In_674,In_47);
and U767 (N_767,N_318,N_478);
xor U768 (N_768,In_1024,N_15);
and U769 (N_769,In_945,In_464);
nand U770 (N_770,N_565,In_1442);
and U771 (N_771,In_1565,In_1135);
xnor U772 (N_772,In_665,In_470);
and U773 (N_773,In_1976,In_19);
and U774 (N_774,In_156,N_457);
nor U775 (N_775,In_1753,In_1458);
nand U776 (N_776,In_1922,In_1988);
and U777 (N_777,In_1625,In_1687);
or U778 (N_778,In_1268,In_1561);
xnor U779 (N_779,In_519,In_1583);
nor U780 (N_780,In_1313,In_1601);
or U781 (N_781,N_497,In_640);
nor U782 (N_782,In_558,In_14);
xor U783 (N_783,In_1707,In_392);
xnor U784 (N_784,N_569,In_513);
nand U785 (N_785,In_791,N_342);
or U786 (N_786,N_568,N_591);
xor U787 (N_787,N_143,In_113);
nor U788 (N_788,In_20,N_549);
and U789 (N_789,N_506,In_1489);
or U790 (N_790,In_1330,In_943);
and U791 (N_791,N_527,In_469);
nand U792 (N_792,N_40,In_23);
or U793 (N_793,N_22,N_69);
nor U794 (N_794,N_209,N_110);
xor U795 (N_795,In_1842,In_1181);
nand U796 (N_796,N_390,In_1165);
nor U797 (N_797,N_571,N_596);
xnor U798 (N_798,In_1635,N_36);
xnor U799 (N_799,In_370,In_1261);
xor U800 (N_800,N_176,In_784);
or U801 (N_801,N_650,N_307);
xnor U802 (N_802,In_449,N_480);
xor U803 (N_803,In_786,N_651);
nand U804 (N_804,In_1391,N_653);
nand U805 (N_805,N_767,In_1302);
xor U806 (N_806,N_628,In_1474);
and U807 (N_807,In_11,In_1300);
nor U808 (N_808,In_754,In_1128);
nand U809 (N_809,N_540,N_531);
nor U810 (N_810,In_83,In_343);
and U811 (N_811,In_1119,In_501);
nand U812 (N_812,In_856,N_242);
nor U813 (N_813,In_1027,In_1245);
and U814 (N_814,In_633,In_39);
nor U815 (N_815,In_153,In_320);
nand U816 (N_816,In_220,In_359);
and U817 (N_817,N_168,N_198);
and U818 (N_818,In_1142,In_1665);
xnor U819 (N_819,In_849,In_539);
or U820 (N_820,In_1773,N_697);
nor U821 (N_821,In_510,N_354);
nor U822 (N_822,N_159,N_336);
nand U823 (N_823,In_490,In_1463);
xor U824 (N_824,N_660,In_1063);
and U825 (N_825,In_852,N_602);
xnor U826 (N_826,In_855,N_195);
xor U827 (N_827,N_189,In_608);
nand U828 (N_828,In_497,N_281);
or U829 (N_829,N_276,In_1221);
nor U830 (N_830,N_368,In_813);
and U831 (N_831,In_794,In_1616);
nor U832 (N_832,N_739,In_1597);
nand U833 (N_833,In_18,N_538);
and U834 (N_834,N_328,N_55);
and U835 (N_835,N_718,N_779);
nor U836 (N_836,N_414,In_1130);
or U837 (N_837,N_791,In_1219);
nand U838 (N_838,In_1294,In_430);
or U839 (N_839,In_1059,N_639);
or U840 (N_840,N_481,N_117);
and U841 (N_841,In_1851,N_424);
nand U842 (N_842,In_1577,In_1430);
or U843 (N_843,In_173,In_341);
and U844 (N_844,N_737,In_1043);
nor U845 (N_845,N_668,In_1247);
and U846 (N_846,In_1388,In_299);
xnor U847 (N_847,N_158,In_433);
xor U848 (N_848,In_1775,In_1535);
nand U849 (N_849,In_1292,N_427);
or U850 (N_850,N_413,N_44);
or U851 (N_851,In_564,In_441);
xnor U852 (N_852,N_314,In_1423);
or U853 (N_853,In_1205,N_217);
or U854 (N_854,N_359,In_1155);
and U855 (N_855,In_1065,N_156);
nand U856 (N_856,N_293,In_96);
xnor U857 (N_857,In_1222,In_1776);
nand U858 (N_858,In_44,N_477);
or U859 (N_859,N_81,N_163);
nor U860 (N_860,N_363,In_993);
or U861 (N_861,N_288,In_1260);
nor U862 (N_862,In_1233,N_443);
or U863 (N_863,In_972,N_113);
nand U864 (N_864,In_766,In_456);
nor U865 (N_865,In_255,In_578);
or U866 (N_866,In_1667,In_843);
nor U867 (N_867,In_256,N_750);
and U868 (N_868,In_59,In_26);
nand U869 (N_869,In_1524,In_862);
or U870 (N_870,N_552,In_231);
nand U871 (N_871,In_1644,In_1439);
xnor U872 (N_872,In_297,N_644);
or U873 (N_873,In_1927,N_30);
and U874 (N_874,In_1092,In_1760);
or U875 (N_875,N_397,In_511);
or U876 (N_876,In_312,N_316);
or U877 (N_877,N_225,N_371);
or U878 (N_878,N_360,In_637);
and U879 (N_879,N_771,In_1482);
xor U880 (N_880,N_663,In_961);
nand U881 (N_881,N_323,N_402);
and U882 (N_882,In_747,In_798);
and U883 (N_883,In_969,N_440);
or U884 (N_884,In_313,In_476);
nand U885 (N_885,In_1831,N_684);
xnor U886 (N_886,N_70,In_1004);
nor U887 (N_887,In_829,In_1896);
nor U888 (N_888,N_499,In_321);
nand U889 (N_889,In_724,In_34);
and U890 (N_890,N_630,In_1343);
nand U891 (N_891,In_1915,In_1924);
nor U892 (N_892,In_1478,N_208);
or U893 (N_893,In_446,In_942);
nor U894 (N_894,N_395,N_352);
nor U895 (N_895,In_1308,In_293);
xor U896 (N_896,N_669,In_436);
xnor U897 (N_897,In_712,In_1804);
or U898 (N_898,N_317,In_1604);
nor U899 (N_899,N_265,In_1944);
xor U900 (N_900,N_557,In_1348);
or U901 (N_901,In_560,N_418);
nand U902 (N_902,In_202,N_732);
nand U903 (N_903,N_710,In_1);
or U904 (N_904,In_1494,N_213);
nand U905 (N_905,N_759,N_131);
nor U906 (N_906,In_1244,In_389);
xor U907 (N_907,N_634,N_312);
and U908 (N_908,N_680,In_499);
xor U909 (N_909,N_721,N_187);
and U910 (N_910,In_584,N_99);
or U911 (N_911,N_254,N_430);
or U912 (N_912,In_1726,In_465);
xor U913 (N_913,In_406,In_414);
and U914 (N_914,In_922,In_437);
nand U915 (N_915,N_582,In_1516);
xor U916 (N_916,In_780,In_141);
nor U917 (N_917,In_1964,N_785);
nor U918 (N_918,In_1857,In_381);
nor U919 (N_919,In_866,N_329);
xnor U920 (N_920,N_762,N_262);
xor U921 (N_921,N_313,N_786);
or U922 (N_922,In_118,In_296);
or U923 (N_923,In_1469,In_1886);
nor U924 (N_924,In_1539,In_1001);
nand U925 (N_925,N_407,N_656);
nor U926 (N_926,N_789,In_1010);
nand U927 (N_927,N_241,N_42);
nand U928 (N_928,In_1521,In_1553);
xor U929 (N_929,In_930,N_387);
and U930 (N_930,In_1562,N_61);
nor U931 (N_931,In_273,In_1630);
xor U932 (N_932,In_265,In_848);
nor U933 (N_933,In_1677,In_1346);
or U934 (N_934,N_410,In_1693);
nor U935 (N_935,N_613,In_205);
or U936 (N_936,N_577,N_14);
nor U937 (N_937,N_713,In_896);
and U938 (N_938,N_406,In_380);
nor U939 (N_939,In_1617,In_687);
xnor U940 (N_940,N_523,N_64);
and U941 (N_941,In_1809,In_236);
xor U942 (N_942,N_589,N_545);
nor U943 (N_943,N_753,In_913);
nand U944 (N_944,N_204,In_1960);
and U945 (N_945,In_1195,N_729);
and U946 (N_946,In_1764,In_1808);
xor U947 (N_947,In_1703,N_760);
xor U948 (N_948,N_448,N_231);
and U949 (N_949,In_677,In_1860);
nand U950 (N_950,In_145,In_283);
or U951 (N_951,In_1550,In_593);
or U952 (N_952,In_907,N_522);
nor U953 (N_953,N_107,In_1323);
and U954 (N_954,In_577,N_768);
nor U955 (N_955,In_1379,N_28);
nor U956 (N_956,In_1774,In_1197);
and U957 (N_957,In_1905,N_178);
or U958 (N_958,N_503,N_698);
and U959 (N_959,In_1336,In_192);
xnor U960 (N_960,N_188,In_729);
or U961 (N_961,N_875,N_116);
xnor U962 (N_962,In_1848,N_517);
xnor U963 (N_963,In_279,N_733);
xor U964 (N_964,In_533,In_227);
nand U965 (N_965,N_803,N_641);
and U966 (N_966,In_504,In_630);
nor U967 (N_967,In_1297,N_720);
and U968 (N_968,N_320,In_1069);
nand U969 (N_969,N_526,In_822);
nand U970 (N_970,N_917,In_611);
nand U971 (N_971,N_337,N_305);
or U972 (N_972,N_843,In_1414);
or U973 (N_973,N_857,N_844);
nor U974 (N_974,N_839,In_1662);
nor U975 (N_975,N_929,In_1109);
xor U976 (N_976,In_662,In_410);
xor U977 (N_977,In_405,N_784);
nor U978 (N_978,N_938,N_883);
nand U979 (N_979,N_717,In_1175);
and U980 (N_980,In_1995,In_1435);
nand U981 (N_981,In_134,N_609);
nor U982 (N_982,In_151,In_88);
and U983 (N_983,In_1686,In_1931);
xnor U984 (N_984,In_1926,In_1054);
xor U985 (N_985,In_493,In_425);
or U986 (N_986,In_714,In_1694);
nor U987 (N_987,In_1240,In_391);
or U988 (N_988,N_763,In_65);
or U989 (N_989,In_1879,In_1263);
nand U990 (N_990,N_858,In_892);
and U991 (N_991,N_643,N_510);
nor U992 (N_992,N_147,In_927);
nand U993 (N_993,In_820,In_1422);
nor U994 (N_994,N_570,In_1780);
nor U995 (N_995,In_1492,N_946);
or U996 (N_996,In_676,N_695);
or U997 (N_997,N_474,In_1002);
xor U998 (N_998,In_43,N_127);
xnor U999 (N_999,In_1410,N_428);
nand U1000 (N_1000,N_385,N_776);
nand U1001 (N_1001,N_793,N_743);
and U1002 (N_1002,N_678,N_256);
or U1003 (N_1003,In_258,In_1298);
nor U1004 (N_1004,N_770,In_581);
or U1005 (N_1005,In_1818,N_558);
xor U1006 (N_1006,In_1989,N_551);
nor U1007 (N_1007,N_866,In_880);
xnor U1008 (N_1008,In_262,N_544);
and U1009 (N_1009,N_340,In_364);
or U1010 (N_1010,In_1542,N_475);
nand U1011 (N_1011,In_1393,In_420);
and U1012 (N_1012,In_310,In_1909);
xor U1013 (N_1013,N_892,In_138);
or U1014 (N_1014,N_227,In_679);
or U1015 (N_1015,N_109,N_635);
xnor U1016 (N_1016,N_815,N_934);
nand U1017 (N_1017,In_1299,In_467);
nand U1018 (N_1018,In_691,N_349);
nand U1019 (N_1019,In_963,N_860);
nor U1020 (N_1020,N_889,N_374);
xor U1021 (N_1021,In_923,N_676);
nand U1022 (N_1022,N_888,N_848);
nand U1023 (N_1023,N_853,N_719);
nand U1024 (N_1024,N_766,N_949);
nor U1025 (N_1025,N_862,In_232);
nor U1026 (N_1026,In_1967,N_901);
nor U1027 (N_1027,N_726,N_675);
xor U1028 (N_1028,N_559,N_805);
nand U1029 (N_1029,In_309,N_741);
or U1030 (N_1030,In_60,N_810);
xnor U1031 (N_1031,In_1368,In_1543);
xor U1032 (N_1032,N_871,In_1203);
nor U1033 (N_1033,In_768,N_386);
xnor U1034 (N_1034,N_714,N_72);
and U1035 (N_1035,N_868,N_722);
xnor U1036 (N_1036,N_792,N_734);
xor U1037 (N_1037,N_752,N_494);
and U1038 (N_1038,N_819,In_327);
and U1039 (N_1039,In_795,In_1898);
nand U1040 (N_1040,N_646,In_1148);
xnor U1041 (N_1041,In_811,N_932);
xor U1042 (N_1042,N_603,N_884);
nand U1043 (N_1043,N_473,N_532);
nor U1044 (N_1044,N_488,In_1986);
nor U1045 (N_1045,N_704,In_1997);
xnor U1046 (N_1046,N_190,N_575);
and U1047 (N_1047,In_755,N_555);
nor U1048 (N_1048,In_1771,In_827);
nand U1049 (N_1049,N_816,In_911);
or U1050 (N_1050,In_826,N_821);
or U1051 (N_1051,In_881,In_821);
or U1052 (N_1052,N_872,In_1660);
nor U1053 (N_1053,In_1337,In_1068);
or U1054 (N_1054,N_18,N_626);
nand U1055 (N_1055,In_1236,N_959);
or U1056 (N_1056,N_958,N_813);
and U1057 (N_1057,N_703,N_665);
xor U1058 (N_1058,N_405,N_112);
xor U1059 (N_1059,In_1923,N_174);
nor U1060 (N_1060,N_631,N_560);
and U1061 (N_1061,In_479,In_206);
nor U1062 (N_1062,N_951,In_617);
xnor U1063 (N_1063,In_331,In_1993);
nor U1064 (N_1064,In_146,N_736);
or U1065 (N_1065,In_1225,In_1855);
and U1066 (N_1066,N_645,N_855);
nor U1067 (N_1067,N_715,N_324);
or U1068 (N_1068,N_914,N_735);
or U1069 (N_1069,N_859,N_180);
and U1070 (N_1070,N_619,In_1564);
xnor U1071 (N_1071,In_653,N_579);
or U1072 (N_1072,N_607,In_757);
or U1073 (N_1073,In_1974,In_401);
nand U1074 (N_1074,N_913,N_764);
xor U1075 (N_1075,In_1462,In_1839);
and U1076 (N_1076,N_10,In_1052);
xnor U1077 (N_1077,N_807,N_911);
or U1078 (N_1078,N_880,N_252);
or U1079 (N_1079,N_850,N_369);
or U1080 (N_1080,N_330,N_41);
nand U1081 (N_1081,In_382,N_809);
and U1082 (N_1082,N_700,In_1154);
nand U1083 (N_1083,In_883,In_1234);
xnor U1084 (N_1084,N_667,N_707);
xnor U1085 (N_1085,N_182,In_152);
nand U1086 (N_1086,N_584,In_266);
and U1087 (N_1087,In_1319,In_1238);
nor U1088 (N_1088,N_572,N_465);
nor U1089 (N_1089,N_384,In_1636);
and U1090 (N_1090,N_563,N_950);
nor U1091 (N_1091,In_1381,N_291);
nor U1092 (N_1092,In_522,In_1115);
nor U1093 (N_1093,In_25,In_970);
and U1094 (N_1094,N_837,In_1055);
or U1095 (N_1095,N_212,In_1217);
and U1096 (N_1096,In_282,N_7);
nor U1097 (N_1097,N_567,N_903);
nand U1098 (N_1098,N_250,N_484);
nand U1099 (N_1099,N_185,N_598);
nand U1100 (N_1100,In_1948,N_419);
xor U1101 (N_1101,In_1605,N_203);
nand U1102 (N_1102,In_587,N_434);
and U1103 (N_1103,N_524,N_794);
and U1104 (N_1104,In_1455,N_505);
nor U1105 (N_1105,In_561,N_823);
and U1106 (N_1106,N_812,In_708);
or U1107 (N_1107,In_1250,N_126);
nand U1108 (N_1108,N_761,N_207);
and U1109 (N_1109,In_322,In_1283);
and U1110 (N_1110,N_456,In_1796);
xor U1111 (N_1111,In_1678,N_490);
nand U1112 (N_1112,In_191,In_174);
and U1113 (N_1113,In_605,In_1725);
or U1114 (N_1114,N_899,N_674);
nor U1115 (N_1115,In_897,N_80);
nor U1116 (N_1116,In_807,N_829);
xor U1117 (N_1117,In_224,In_651);
xor U1118 (N_1118,In_455,N_748);
and U1119 (N_1119,In_104,N_956);
nor U1120 (N_1120,N_1026,In_623);
and U1121 (N_1121,N_746,N_1054);
nand U1122 (N_1122,In_1341,N_574);
xor U1123 (N_1123,N_197,In_1316);
nand U1124 (N_1124,N_612,N_404);
or U1125 (N_1125,N_982,N_205);
nor U1126 (N_1126,In_1269,N_1030);
nor U1127 (N_1127,In_393,N_924);
and U1128 (N_1128,N_1041,N_1070);
nor U1129 (N_1129,N_546,In_1706);
nand U1130 (N_1130,N_192,In_1397);
or U1131 (N_1131,N_930,In_54);
xor U1132 (N_1132,In_122,In_673);
nor U1133 (N_1133,In_887,N_561);
nand U1134 (N_1134,N_454,N_942);
and U1135 (N_1135,In_1940,N_830);
and U1136 (N_1136,In_1590,In_241);
and U1137 (N_1137,N_725,N_811);
nor U1138 (N_1138,N_765,N_466);
and U1139 (N_1139,In_800,N_509);
nor U1140 (N_1140,In_371,In_1575);
xor U1141 (N_1141,In_546,In_697);
and U1142 (N_1142,N_968,N_908);
nand U1143 (N_1143,In_1739,In_1969);
nor U1144 (N_1144,N_1015,N_820);
xor U1145 (N_1145,N_890,In_4);
and U1146 (N_1146,In_1158,N_1072);
nand U1147 (N_1147,In_1003,N_1001);
xnor U1148 (N_1148,In_600,In_557);
or U1149 (N_1149,N_1025,N_1085);
or U1150 (N_1150,N_981,In_1087);
nand U1151 (N_1151,N_375,N_1110);
or U1152 (N_1152,N_943,N_1053);
and U1153 (N_1153,N_389,N_1028);
xnor U1154 (N_1154,In_215,In_1449);
nor U1155 (N_1155,N_1105,N_966);
xnor U1156 (N_1156,In_1394,In_190);
or U1157 (N_1157,N_879,In_1072);
nor U1158 (N_1158,In_824,N_1111);
xnor U1159 (N_1159,N_781,In_357);
nor U1160 (N_1160,N_1008,In_1033);
or U1161 (N_1161,N_947,N_840);
nor U1162 (N_1162,N_238,N_516);
nand U1163 (N_1163,In_1671,In_1199);
or U1164 (N_1164,In_1497,N_841);
nor U1165 (N_1165,N_939,N_367);
or U1166 (N_1166,In_1378,In_777);
and U1167 (N_1167,In_275,N_796);
and U1168 (N_1168,N_898,N_690);
xnor U1169 (N_1169,N_894,N_1052);
xor U1170 (N_1170,In_574,N_1003);
nand U1171 (N_1171,In_902,N_514);
nand U1172 (N_1172,In_1531,N_778);
xnor U1173 (N_1173,N_214,N_679);
or U1174 (N_1174,N_907,In_660);
nand U1175 (N_1175,N_945,In_547);
xor U1176 (N_1176,In_1016,In_1053);
and U1177 (N_1177,N_1004,N_1113);
or U1178 (N_1178,N_1104,N_1095);
and U1179 (N_1179,N_1109,N_492);
xnor U1180 (N_1180,N_1023,N_919);
or U1181 (N_1181,N_476,N_16);
nand U1182 (N_1182,N_491,In_1147);
xor U1183 (N_1183,In_588,In_1307);
and U1184 (N_1184,In_488,N_637);
and U1185 (N_1185,N_464,In_453);
and U1186 (N_1186,In_403,N_145);
nand U1187 (N_1187,In_117,N_799);
nand U1188 (N_1188,In_607,In_1513);
or U1189 (N_1189,N_687,N_999);
nand U1190 (N_1190,In_1493,N_874);
xor U1191 (N_1191,In_101,N_588);
nor U1192 (N_1192,N_642,N_120);
nor U1193 (N_1193,N_638,In_1322);
nor U1194 (N_1194,N_906,N_462);
nor U1195 (N_1195,In_1070,N_1103);
nand U1196 (N_1196,N_399,N_1006);
nor U1197 (N_1197,In_516,N_171);
and U1198 (N_1198,In_180,In_387);
nor U1199 (N_1199,N_623,In_666);
nor U1200 (N_1200,N_161,In_695);
or U1201 (N_1201,In_48,N_417);
and U1202 (N_1202,N_1087,N_912);
xnor U1203 (N_1203,In_1880,In_535);
or U1204 (N_1204,N_594,In_740);
nand U1205 (N_1205,N_1014,In_1331);
nand U1206 (N_1206,N_832,N_486);
nand U1207 (N_1207,In_924,N_576);
and U1208 (N_1208,In_702,N_108);
and U1209 (N_1209,N_459,N_769);
nor U1210 (N_1210,N_960,N_990);
or U1211 (N_1211,In_1421,N_712);
or U1212 (N_1212,N_1042,In_726);
and U1213 (N_1213,In_1559,In_1456);
nand U1214 (N_1214,In_1073,N_940);
nor U1215 (N_1215,N_896,N_1108);
xor U1216 (N_1216,N_979,N_808);
xnor U1217 (N_1217,N_997,In_1317);
nand U1218 (N_1218,In_213,N_845);
and U1219 (N_1219,In_1324,In_1479);
or U1220 (N_1220,N_802,N_173);
and U1221 (N_1221,N_1017,In_760);
and U1222 (N_1222,N_747,In_1106);
nand U1223 (N_1223,N_239,N_742);
nor U1224 (N_1224,In_485,N_304);
or U1225 (N_1225,N_502,In_1117);
and U1226 (N_1226,In_1918,N_806);
or U1227 (N_1227,N_583,N_525);
or U1228 (N_1228,N_935,In_1975);
nor U1229 (N_1229,N_496,N_1045);
nor U1230 (N_1230,In_1982,N_922);
nand U1231 (N_1231,In_879,N_988);
and U1232 (N_1232,N_1115,In_95);
nor U1233 (N_1233,In_551,N_962);
xor U1234 (N_1234,N_122,N_798);
or U1235 (N_1235,N_611,In_819);
or U1236 (N_1236,N_833,N_451);
nand U1237 (N_1237,N_936,N_831);
or U1238 (N_1238,N_804,In_133);
xnor U1239 (N_1239,N_847,In_1643);
nor U1240 (N_1240,In_445,In_311);
or U1241 (N_1241,N_501,N_774);
nor U1242 (N_1242,N_728,In_193);
xnor U1243 (N_1243,In_976,N_694);
nor U1244 (N_1244,N_321,In_338);
nand U1245 (N_1245,In_718,N_671);
xor U1246 (N_1246,N_877,In_1889);
nor U1247 (N_1247,N_955,N_921);
nor U1248 (N_1248,N_1051,In_598);
nand U1249 (N_1249,In_1390,N_586);
or U1250 (N_1250,N_1119,In_959);
nand U1251 (N_1251,In_1722,N_500);
xor U1252 (N_1252,In_1586,N_627);
nor U1253 (N_1253,N_57,In_261);
nand U1254 (N_1254,N_954,N_553);
and U1255 (N_1255,In_1854,N_773);
xor U1256 (N_1256,N_606,N_537);
nand U1257 (N_1257,N_937,N_468);
or U1258 (N_1258,In_1945,N_601);
or U1259 (N_1259,In_853,N_587);
nand U1260 (N_1260,N_564,N_1074);
or U1261 (N_1261,In_951,N_964);
or U1262 (N_1262,N_854,N_976);
xnor U1263 (N_1263,In_860,In_199);
and U1264 (N_1264,N_692,N_29);
or U1265 (N_1265,N_1000,N_566);
nand U1266 (N_1266,N_918,N_944);
xor U1267 (N_1267,In_709,In_514);
and U1268 (N_1268,In_723,In_858);
nor U1269 (N_1269,N_1056,In_1623);
nand U1270 (N_1270,In_1103,In_1365);
nand U1271 (N_1271,N_356,N_237);
or U1272 (N_1272,In_459,In_1946);
or U1273 (N_1273,N_856,In_919);
nand U1274 (N_1274,N_479,N_144);
nand U1275 (N_1275,N_817,N_666);
nand U1276 (N_1276,In_1120,N_985);
and U1277 (N_1277,N_556,N_485);
nor U1278 (N_1278,N_274,N_148);
nand U1279 (N_1279,N_299,In_1941);
and U1280 (N_1280,N_1172,In_1214);
or U1281 (N_1281,N_1202,N_512);
nand U1282 (N_1282,N_617,N_562);
nor U1283 (N_1283,N_1185,N_1178);
and U1284 (N_1284,N_863,N_275);
and U1285 (N_1285,In_667,N_1277);
and U1286 (N_1286,N_1116,N_1204);
nor U1287 (N_1287,In_661,In_1919);
or U1288 (N_1288,N_455,In_149);
and U1289 (N_1289,In_1875,In_107);
nor U1290 (N_1290,N_659,N_995);
nor U1291 (N_1291,In_751,N_931);
xnor U1292 (N_1292,N_677,N_961);
nor U1293 (N_1293,N_1044,N_230);
xnor U1294 (N_1294,N_1150,N_1263);
xnor U1295 (N_1295,In_1845,N_1273);
nor U1296 (N_1296,In_1827,N_825);
or U1297 (N_1297,N_1226,In_51);
xor U1298 (N_1298,N_1118,In_1533);
nand U1299 (N_1299,N_614,In_1056);
and U1300 (N_1300,In_592,In_1159);
nor U1301 (N_1301,N_1222,N_315);
nor U1302 (N_1302,N_957,In_1444);
xnor U1303 (N_1303,N_923,N_1132);
nand U1304 (N_1304,N_849,N_1123);
xor U1305 (N_1305,N_1078,N_1252);
nor U1306 (N_1306,N_1011,N_1265);
or U1307 (N_1307,In_1280,N_164);
nor U1308 (N_1308,N_1084,N_426);
nor U1309 (N_1309,In_408,N_1093);
xor U1310 (N_1310,In_1187,N_79);
or U1311 (N_1311,N_851,In_914);
xor U1312 (N_1312,N_1022,In_1802);
and U1313 (N_1313,In_1008,N_1027);
nand U1314 (N_1314,N_1244,N_1144);
nand U1315 (N_1315,N_1050,N_654);
nor U1316 (N_1316,N_1158,N_1018);
nand U1317 (N_1317,In_276,N_310);
xnor U1318 (N_1318,In_793,N_716);
or U1319 (N_1319,N_1207,In_1663);
and U1320 (N_1320,N_640,In_81);
or U1321 (N_1321,N_1199,N_1164);
xnor U1322 (N_1322,N_891,N_1081);
xnor U1323 (N_1323,In_978,In_229);
or U1324 (N_1324,N_1157,N_513);
xnor U1325 (N_1325,In_1071,In_1164);
or U1326 (N_1326,N_996,In_447);
nor U1327 (N_1327,N_519,N_1020);
nor U1328 (N_1328,N_693,In_1688);
nor U1329 (N_1329,In_672,N_1089);
xnor U1330 (N_1330,N_795,N_394);
nor U1331 (N_1331,In_1329,N_893);
and U1332 (N_1332,N_243,In_1873);
nor U1333 (N_1333,N_1055,N_648);
or U1334 (N_1334,N_1002,N_755);
or U1335 (N_1335,In_78,N_933);
nor U1336 (N_1336,N_1129,N_657);
xnor U1337 (N_1337,N_1166,N_1241);
and U1338 (N_1338,N_1163,N_1194);
xor U1339 (N_1339,N_1068,In_1648);
nor U1340 (N_1340,N_1149,In_66);
nor U1341 (N_1341,N_967,N_1189);
nand U1342 (N_1342,N_1235,N_1203);
and U1343 (N_1343,N_777,N_1029);
nand U1344 (N_1344,N_800,N_983);
nand U1345 (N_1345,In_783,N_1083);
or U1346 (N_1346,In_1078,N_632);
nor U1347 (N_1347,N_123,N_1248);
xnor U1348 (N_1348,N_948,N_50);
or U1349 (N_1349,N_870,In_582);
nor U1350 (N_1350,N_1217,N_1279);
and U1351 (N_1351,N_1255,N_1160);
nand U1352 (N_1352,N_1007,N_909);
or U1353 (N_1353,N_1162,N_1013);
or U1354 (N_1354,In_512,In_1139);
and U1355 (N_1355,In_1734,N_1278);
nor U1356 (N_1356,In_1716,In_1032);
and U1357 (N_1357,N_691,In_1274);
or U1358 (N_1358,N_1032,In_340);
nand U1359 (N_1359,N_1156,N_370);
or U1360 (N_1360,N_842,N_372);
nand U1361 (N_1361,In_701,N_578);
nand U1362 (N_1362,N_1234,In_1160);
xor U1363 (N_1363,In_1402,N_533);
nor U1364 (N_1364,In_1176,N_66);
nand U1365 (N_1365,N_452,N_1237);
xnor U1366 (N_1366,N_885,N_882);
and U1367 (N_1367,N_1066,N_1256);
or U1368 (N_1368,N_1098,N_1031);
nand U1369 (N_1369,In_1602,In_395);
nand U1370 (N_1370,In_1470,N_1137);
and U1371 (N_1371,N_60,N_1173);
nor U1372 (N_1372,In_468,N_86);
xor U1373 (N_1373,In_351,N_365);
xnor U1374 (N_1374,N_438,N_886);
and U1375 (N_1375,N_780,In_1243);
xnor U1376 (N_1376,In_1620,In_358);
nand U1377 (N_1377,N_1169,N_1179);
or U1378 (N_1378,N_423,N_846);
and U1379 (N_1379,N_978,N_1106);
nor U1380 (N_1380,N_1262,In_1702);
xor U1381 (N_1381,N_1214,N_867);
xor U1382 (N_1382,N_1216,N_1100);
or U1383 (N_1383,N_1099,N_1246);
nor U1384 (N_1384,N_1219,In_1701);
and U1385 (N_1385,N_757,N_1121);
or U1386 (N_1386,In_452,N_339);
or U1387 (N_1387,N_25,N_701);
or U1388 (N_1388,N_9,N_347);
nor U1389 (N_1389,N_515,In_622);
nand U1390 (N_1390,In_1014,N_177);
and U1391 (N_1391,N_724,N_925);
and U1392 (N_1392,In_1612,N_740);
or U1393 (N_1393,N_1071,N_986);
xnor U1394 (N_1394,N_971,In_225);
nand U1395 (N_1395,N_824,In_1816);
or U1396 (N_1396,In_1352,N_534);
nand U1397 (N_1397,In_638,In_50);
xnor U1398 (N_1398,In_1162,N_1171);
nor U1399 (N_1399,In_100,N_1155);
xor U1400 (N_1400,N_289,N_295);
nor U1401 (N_1401,N_673,N_797);
nor U1402 (N_1402,In_524,In_1318);
and U1403 (N_1403,N_1210,N_1161);
or U1404 (N_1404,N_1201,N_1208);
nand U1405 (N_1405,N_306,N_536);
nand U1406 (N_1406,In_1748,N_974);
or U1407 (N_1407,N_332,N_916);
or U1408 (N_1408,N_467,In_1645);
or U1409 (N_1409,N_1046,N_788);
nand U1410 (N_1410,N_1272,In_79);
xor U1411 (N_1411,In_509,In_1647);
xor U1412 (N_1412,N_790,N_91);
or U1413 (N_1413,N_987,N_1251);
xor U1414 (N_1414,In_982,N_900);
nand U1415 (N_1415,N_1128,In_1472);
nor U1416 (N_1416,N_507,N_688);
nor U1417 (N_1417,In_544,N_350);
xor U1418 (N_1418,In_422,N_290);
nand U1419 (N_1419,N_984,N_548);
and U1420 (N_1420,N_664,N_649);
xnor U1421 (N_1421,N_1220,N_1154);
and U1422 (N_1422,N_754,N_364);
and U1423 (N_1423,In_140,In_1309);
nor U1424 (N_1424,N_965,In_72);
or U1425 (N_1425,N_625,N_1253);
nand U1426 (N_1426,N_401,N_1139);
and U1427 (N_1427,In_1881,N_910);
nand U1428 (N_1428,N_1091,In_378);
xor U1429 (N_1429,N_647,N_260);
nand U1430 (N_1430,N_135,In_1066);
or U1431 (N_1431,In_1674,N_98);
xor U1432 (N_1432,N_1125,N_869);
nand U1433 (N_1433,In_1477,In_1906);
or U1434 (N_1434,In_928,In_739);
and U1435 (N_1435,N_991,N_1079);
and U1436 (N_1436,N_1200,N_1101);
nor U1437 (N_1437,N_1141,N_1259);
or U1438 (N_1438,N_547,In_434);
or U1439 (N_1439,N_1225,N_1238);
nand U1440 (N_1440,In_1607,N_969);
nor U1441 (N_1441,In_251,N_878);
nor U1442 (N_1442,N_941,In_1361);
and U1443 (N_1443,In_1837,N_652);
nand U1444 (N_1444,N_1390,N_1260);
or U1445 (N_1445,N_1344,N_1288);
nor U1446 (N_1446,In_1811,N_493);
or U1447 (N_1447,N_580,N_1375);
nor U1448 (N_1448,In_613,N_1384);
and U1449 (N_1449,N_1389,N_836);
nand U1450 (N_1450,In_1794,N_1307);
xnor U1451 (N_1451,N_1348,N_1124);
nand U1452 (N_1452,N_953,In_263);
or U1453 (N_1453,N_1430,N_711);
nand U1454 (N_1454,N_1190,In_1697);
nor U1455 (N_1455,N_1414,N_1254);
nand U1456 (N_1456,N_1410,N_68);
nand U1457 (N_1457,N_1245,N_1309);
or U1458 (N_1458,N_685,N_655);
or U1459 (N_1459,In_396,In_1360);
and U1460 (N_1460,N_1406,N_928);
and U1461 (N_1461,N_1126,N_1140);
nor U1462 (N_1462,N_1133,In_1281);
nand U1463 (N_1463,N_530,N_1360);
nand U1464 (N_1464,N_818,N_1080);
xnor U1465 (N_1465,N_1405,In_369);
nand U1466 (N_1466,N_738,N_1224);
nand U1467 (N_1467,In_1333,N_745);
and U1468 (N_1468,N_1332,N_1403);
or U1469 (N_1469,N_783,In_1595);
and U1470 (N_1470,In_421,N_622);
and U1471 (N_1471,N_1094,N_1250);
xnor U1472 (N_1472,N_1432,N_1306);
nand U1473 (N_1473,N_1047,N_977);
or U1474 (N_1474,N_1315,N_1363);
nor U1475 (N_1475,N_421,N_992);
and U1476 (N_1476,In_93,In_1288);
or U1477 (N_1477,In_1934,N_702);
and U1478 (N_1478,N_994,N_1283);
xnor U1479 (N_1479,N_1012,N_1354);
nand U1480 (N_1480,N_1435,N_1352);
nor U1481 (N_1481,N_975,N_1142);
and U1482 (N_1482,N_1314,In_1888);
xor U1483 (N_1483,N_887,N_926);
nand U1484 (N_1484,In_221,N_1322);
and U1485 (N_1485,In_264,N_1347);
and U1486 (N_1486,N_1334,N_1183);
nor U1487 (N_1487,N_993,N_1327);
xor U1488 (N_1488,N_1439,N_672);
or U1489 (N_1489,N_1300,In_1285);
and U1490 (N_1490,In_636,N_1159);
and U1491 (N_1491,In_1572,N_1061);
and U1492 (N_1492,In_1892,N_730);
and U1493 (N_1493,N_1043,N_1134);
nand U1494 (N_1494,N_1009,In_15);
or U1495 (N_1495,N_621,N_1393);
xnor U1496 (N_1496,N_1213,N_1148);
xnor U1497 (N_1497,In_1399,N_1324);
nor U1498 (N_1498,N_1395,N_1077);
nand U1499 (N_1499,N_435,In_1498);
or U1500 (N_1500,N_379,N_376);
nand U1501 (N_1501,In_243,N_1049);
xnor U1502 (N_1502,In_801,N_1368);
nor U1503 (N_1503,N_1399,N_1285);
xor U1504 (N_1504,N_972,N_1343);
nor U1505 (N_1505,N_1112,N_1400);
xor U1506 (N_1506,N_1404,N_272);
and U1507 (N_1507,In_42,N_1365);
nor U1508 (N_1508,N_539,N_1381);
nor U1509 (N_1509,N_1397,N_1036);
xor U1510 (N_1510,N_1388,N_1135);
or U1511 (N_1511,N_952,N_1131);
xnor U1512 (N_1512,N_141,N_1264);
nor U1513 (N_1513,N_1350,N_489);
nor U1514 (N_1514,N_1075,N_1437);
nor U1515 (N_1515,In_1202,N_1402);
and U1516 (N_1516,N_1188,N_75);
or U1517 (N_1517,N_1024,N_1356);
or U1518 (N_1518,In_1548,N_834);
or U1519 (N_1519,N_1114,N_351);
nor U1520 (N_1520,N_1010,In_200);
nor U1521 (N_1521,N_1038,N_1280);
nor U1522 (N_1522,N_1419,In_1062);
and U1523 (N_1523,In_1075,N_861);
xnor U1524 (N_1524,N_1342,N_828);
nor U1525 (N_1525,In_362,N_1302);
or U1526 (N_1526,In_1149,N_618);
xor U1527 (N_1527,In_484,In_1633);
and U1528 (N_1528,N_1323,N_357);
nand U1529 (N_1529,N_915,N_554);
and U1530 (N_1530,N_1040,N_592);
or U1531 (N_1531,N_814,N_1317);
nand U1532 (N_1532,N_1281,N_1175);
xor U1533 (N_1533,N_723,N_1165);
xnor U1534 (N_1534,In_1642,N_1223);
xor U1535 (N_1535,N_1358,N_1233);
nand U1536 (N_1536,N_1290,N_826);
or U1537 (N_1537,N_1424,N_1228);
or U1538 (N_1538,N_1293,N_1409);
and U1539 (N_1539,N_1187,N_1387);
or U1540 (N_1540,N_744,N_1231);
and U1541 (N_1541,N_696,N_1398);
nand U1542 (N_1542,N_1240,N_218);
or U1543 (N_1543,In_417,In_1596);
nor U1544 (N_1544,N_1177,N_1335);
or U1545 (N_1545,N_331,N_1418);
nand U1546 (N_1546,N_865,N_1304);
or U1547 (N_1547,In_1265,N_1386);
nand U1548 (N_1548,N_1058,In_1114);
xor U1549 (N_1549,N_1340,N_1372);
nor U1550 (N_1550,N_1168,N_1429);
or U1551 (N_1551,N_1319,In_1512);
and U1552 (N_1552,N_670,N_681);
or U1553 (N_1553,In_1846,N_1167);
xor U1554 (N_1554,N_1069,N_1086);
xor U1555 (N_1555,N_153,N_1057);
nor U1556 (N_1556,N_749,In_1144);
or U1557 (N_1557,N_1034,In_1229);
nor U1558 (N_1558,N_1308,N_920);
nor U1559 (N_1559,N_1170,N_1211);
or U1560 (N_1560,In_289,In_94);
and U1561 (N_1561,In_33,N_1218);
or U1562 (N_1562,In_1124,N_633);
xor U1563 (N_1563,N_998,N_1318);
nand U1564 (N_1564,In_1963,In_1370);
nor U1565 (N_1565,In_108,N_1380);
and U1566 (N_1566,N_1146,N_1230);
nor U1567 (N_1567,N_1247,N_1421);
nand U1568 (N_1568,N_1195,N_905);
and U1569 (N_1569,N_1312,N_1305);
xnor U1570 (N_1570,In_201,N_1413);
xnor U1571 (N_1571,In_888,N_1174);
or U1572 (N_1572,N_1180,N_686);
or U1573 (N_1573,N_1366,N_1065);
xnor U1574 (N_1574,In_1978,In_796);
or U1575 (N_1575,In_869,N_1383);
or U1576 (N_1576,In_1959,In_155);
and U1577 (N_1577,N_1396,N_1196);
nand U1578 (N_1578,N_334,N_1359);
nor U1579 (N_1579,In_1728,In_719);
nand U1580 (N_1580,N_1426,N_1153);
and U1581 (N_1581,In_962,N_1151);
xnor U1582 (N_1582,N_1361,In_368);
nand U1583 (N_1583,In_1518,N_1325);
nand U1584 (N_1584,N_1391,In_294);
nor U1585 (N_1585,N_1122,In_1481);
nand U1586 (N_1586,In_556,N_1212);
and U1587 (N_1587,N_709,In_704);
xor U1588 (N_1588,In_337,N_1269);
nor U1589 (N_1589,N_782,N_1333);
nor U1590 (N_1590,In_1908,N_775);
or U1591 (N_1591,N_629,N_835);
or U1592 (N_1592,N_1060,N_1433);
and U1593 (N_1593,N_1423,N_1276);
nand U1594 (N_1594,N_658,N_1371);
and U1595 (N_1595,N_1416,N_1227);
or U1596 (N_1596,In_1778,N_1436);
nand U1597 (N_1597,N_251,N_1367);
nor U1598 (N_1598,N_1221,N_1310);
xor U1599 (N_1599,N_1329,In_1715);
and U1600 (N_1600,N_1595,N_1337);
nand U1601 (N_1601,N_963,N_1488);
nor U1602 (N_1602,N_1016,N_1533);
nand U1603 (N_1603,In_699,N_1417);
and U1604 (N_1604,N_1379,N_1483);
xor U1605 (N_1605,In_1862,N_1508);
or U1606 (N_1606,In_680,N_1422);
xor U1607 (N_1607,N_1147,N_1064);
or U1608 (N_1608,N_1524,N_1470);
nand U1609 (N_1609,N_827,N_1385);
or U1610 (N_1610,N_756,N_1512);
nand U1611 (N_1611,N_699,N_1184);
and U1612 (N_1612,N_852,N_1594);
or U1613 (N_1613,N_1563,N_1472);
xnor U1614 (N_1614,N_1525,In_884);
or U1615 (N_1615,N_1507,N_1096);
or U1616 (N_1616,In_9,N_1570);
nand U1617 (N_1617,N_1258,N_1186);
or U1618 (N_1618,N_1456,N_1450);
and U1619 (N_1619,N_1394,N_1464);
nand U1620 (N_1620,In_1102,N_1558);
nand U1621 (N_1621,In_1040,N_1540);
nand U1622 (N_1622,N_294,N_1505);
or U1623 (N_1623,N_970,N_1547);
nor U1624 (N_1624,N_1535,N_1289);
nand U1625 (N_1625,N_1369,N_573);
xor U1626 (N_1626,N_662,N_1268);
or U1627 (N_1627,N_1521,N_1130);
xnor U1628 (N_1628,N_1330,N_1542);
and U1629 (N_1629,N_1355,N_1494);
and U1630 (N_1630,N_1480,In_1515);
nor U1631 (N_1631,In_1925,N_1585);
nand U1632 (N_1632,In_692,In_1858);
or U1633 (N_1633,N_1033,In_1476);
nor U1634 (N_1634,N_902,N_1215);
or U1635 (N_1635,N_838,N_1573);
nor U1636 (N_1636,N_1297,N_1475);
and U1637 (N_1637,N_1107,N_1090);
xor U1638 (N_1638,N_1501,In_1334);
xnor U1639 (N_1639,N_1062,N_1462);
xnor U1640 (N_1640,N_1572,N_1097);
or U1641 (N_1641,N_1441,N_1362);
xnor U1642 (N_1642,N_1382,N_1497);
xnor U1643 (N_1643,N_1449,N_1376);
or U1644 (N_1644,N_1554,N_973);
xnor U1645 (N_1645,N_1448,N_1357);
nand U1646 (N_1646,N_604,In_1761);
xnor U1647 (N_1647,N_470,N_873);
or U1648 (N_1648,N_1556,N_1452);
xor U1649 (N_1649,N_1243,N_1444);
nand U1650 (N_1650,N_1270,N_1331);
xor U1651 (N_1651,N_1539,N_1581);
nand U1652 (N_1652,N_1538,N_1478);
nand U1653 (N_1653,In_1067,N_1537);
xnor U1654 (N_1654,N_377,N_1427);
nand U1655 (N_1655,N_1408,N_1063);
nor U1656 (N_1656,In_954,N_787);
and U1657 (N_1657,In_1057,N_1552);
nand U1658 (N_1658,In_324,N_1261);
or U1659 (N_1659,N_1575,N_1442);
nand U1660 (N_1660,N_1516,N_1313);
xor U1661 (N_1661,N_1353,N_1295);
and U1662 (N_1662,N_1469,N_1320);
or U1663 (N_1663,N_1377,N_1447);
and U1664 (N_1664,N_1345,N_1364);
nand U1665 (N_1665,N_1294,N_1232);
or U1666 (N_1666,N_529,In_1129);
or U1667 (N_1667,In_68,In_349);
or U1668 (N_1668,N_1198,N_1181);
nand U1669 (N_1669,N_1291,N_593);
nand U1670 (N_1670,In_1218,N_1415);
or U1671 (N_1671,N_1443,In_35);
nor U1672 (N_1672,N_1529,In_1649);
nand U1673 (N_1673,N_1067,N_989);
nand U1674 (N_1674,N_1035,N_483);
xnor U1675 (N_1675,N_1490,N_1336);
and U1676 (N_1676,N_297,N_1495);
nand U1677 (N_1677,N_1102,N_1392);
nor U1678 (N_1678,N_610,N_1500);
nor U1679 (N_1679,N_751,N_1136);
xnor U1680 (N_1680,N_1510,In_325);
and U1681 (N_1681,N_1477,N_1229);
and U1682 (N_1682,N_1502,N_1143);
or U1683 (N_1683,N_1513,N_1303);
nand U1684 (N_1684,N_415,N_1496);
nand U1685 (N_1685,In_1592,N_1517);
or U1686 (N_1686,N_1059,In_787);
xor U1687 (N_1687,N_1584,N_1316);
nand U1688 (N_1688,N_535,N_1428);
xor U1689 (N_1689,N_1209,N_1473);
xor U1690 (N_1690,N_1282,N_1526);
xnor U1691 (N_1691,N_683,N_897);
or U1692 (N_1692,N_1589,N_1546);
nor U1693 (N_1693,N_1561,N_1503);
nor U1694 (N_1694,N_1048,N_1286);
nor U1695 (N_1695,N_1438,N_1425);
nor U1696 (N_1696,N_1468,N_1590);
or U1697 (N_1697,N_1555,N_980);
nand U1698 (N_1698,N_772,N_1346);
nand U1699 (N_1699,N_1586,N_1037);
nor U1700 (N_1700,N_1531,N_1566);
or U1701 (N_1701,In_935,N_1466);
or U1702 (N_1702,N_1152,N_1520);
nand U1703 (N_1703,N_1522,In_1354);
nor U1704 (N_1704,N_1491,N_1266);
and U1705 (N_1705,N_1138,N_191);
nor U1706 (N_1706,N_1471,N_1574);
or U1707 (N_1707,N_1192,N_1592);
nor U1708 (N_1708,N_1476,N_1598);
nor U1709 (N_1709,N_1583,N_1249);
or U1710 (N_1710,N_1005,N_1527);
nor U1711 (N_1711,In_274,N_895);
xor U1712 (N_1712,N_1292,N_1541);
or U1713 (N_1713,N_1349,In_1777);
or U1714 (N_1714,N_1545,N_1401);
xnor U1715 (N_1715,In_1876,N_1489);
or U1716 (N_1716,N_1599,N_1588);
nor U1717 (N_1717,In_1484,N_166);
or U1718 (N_1718,N_1518,N_1197);
xnor U1719 (N_1719,N_1596,N_1499);
and U1720 (N_1720,N_1509,N_1562);
nor U1721 (N_1721,N_904,N_1420);
or U1722 (N_1722,N_1560,In_639);
nor U1723 (N_1723,N_1463,N_1474);
xor U1724 (N_1724,N_1523,N_1298);
or U1725 (N_1725,N_1498,N_1559);
nand U1726 (N_1726,N_1458,N_1479);
nor U1727 (N_1727,In_1579,N_801);
xor U1728 (N_1728,N_1536,N_1412);
or U1729 (N_1729,N_82,N_1564);
or U1730 (N_1730,N_1373,N_1571);
or U1731 (N_1731,N_881,N_1576);
xnor U1732 (N_1732,N_1532,N_1236);
nand U1733 (N_1733,N_1550,N_1485);
nand U1734 (N_1734,N_689,N_1321);
nand U1735 (N_1735,In_1047,N_1284);
and U1736 (N_1736,N_1021,N_1275);
nand U1737 (N_1737,N_1073,N_705);
nand U1738 (N_1738,N_1484,N_1482);
nand U1739 (N_1739,N_1549,N_1193);
nand U1740 (N_1740,N_1341,N_1378);
xor U1741 (N_1741,N_876,N_1465);
xor U1742 (N_1742,N_1453,N_1191);
and U1743 (N_1743,In_1551,N_1591);
nor U1744 (N_1744,N_1567,N_1351);
nand U1745 (N_1745,N_758,N_706);
and U1746 (N_1746,N_1519,In_1983);
xnor U1747 (N_1747,In_366,N_1460);
and U1748 (N_1748,N_1092,N_1457);
xnor U1749 (N_1749,N_1565,N_1580);
nand U1750 (N_1750,N_1182,N_1461);
nand U1751 (N_1751,N_1577,N_308);
and U1752 (N_1752,N_111,N_1551);
and U1753 (N_1753,N_1455,N_1145);
xor U1754 (N_1754,N_1451,N_1578);
and U1755 (N_1755,N_1257,N_223);
or U1756 (N_1756,N_1579,N_1534);
nor U1757 (N_1757,N_1434,N_1504);
xor U1758 (N_1758,N_1548,N_1311);
nor U1759 (N_1759,N_864,N_1486);
or U1760 (N_1760,N_1696,N_1655);
or U1761 (N_1761,N_1120,N_1657);
and U1762 (N_1762,N_1742,N_1117);
nor U1763 (N_1763,N_1756,N_1467);
or U1764 (N_1764,In_166,N_1597);
nor U1765 (N_1765,N_1242,N_1659);
and U1766 (N_1766,N_1296,N_1757);
nand U1767 (N_1767,N_1680,In_654);
nor U1768 (N_1768,N_1301,N_682);
and U1769 (N_1769,N_1239,N_1039);
and U1770 (N_1770,N_1741,N_1709);
or U1771 (N_1771,N_1620,N_927);
and U1772 (N_1772,N_1644,N_1672);
nor U1773 (N_1773,N_1671,N_1514);
and U1774 (N_1774,N_1661,N_1748);
nor U1775 (N_1775,N_1743,N_1481);
or U1776 (N_1776,N_1624,N_1528);
or U1777 (N_1777,N_1669,N_396);
and U1778 (N_1778,N_1716,N_1692);
xor U1779 (N_1779,N_1654,N_1370);
xnor U1780 (N_1780,N_1019,N_822);
nand U1781 (N_1781,N_1721,N_1326);
nor U1782 (N_1782,N_1616,N_731);
xor U1783 (N_1783,N_1446,N_1271);
or U1784 (N_1784,N_1758,N_1374);
nand U1785 (N_1785,N_1726,N_1717);
or U1786 (N_1786,N_1205,N_1600);
nor U1787 (N_1787,N_1493,N_1611);
nand U1788 (N_1788,N_1652,N_1687);
nor U1789 (N_1789,N_1623,In_865);
xor U1790 (N_1790,N_1593,N_1662);
xor U1791 (N_1791,N_1587,N_1744);
nand U1792 (N_1792,N_1750,N_1630);
and U1793 (N_1793,N_1627,N_1738);
xor U1794 (N_1794,N_1653,N_1689);
or U1795 (N_1795,N_1607,N_1664);
nand U1796 (N_1796,N_1723,In_1184);
or U1797 (N_1797,N_1082,In_804);
or U1798 (N_1798,In_150,In_1847);
or U1799 (N_1799,N_1734,N_1701);
and U1800 (N_1800,N_1622,N_1718);
xnor U1801 (N_1801,N_1632,N_1730);
and U1802 (N_1802,N_1700,N_1606);
or U1803 (N_1803,N_1732,N_727);
nor U1804 (N_1804,N_1633,N_1642);
nand U1805 (N_1805,N_1629,In_388);
or U1806 (N_1806,N_1407,N_1641);
nor U1807 (N_1807,N_1678,N_661);
xnor U1808 (N_1808,N_1088,N_1656);
xor U1809 (N_1809,N_1712,N_1706);
xnor U1810 (N_1810,N_1698,N_1645);
xnor U1811 (N_1811,N_1759,N_1582);
or U1812 (N_1812,N_1615,N_1515);
nor U1813 (N_1813,N_358,N_1660);
nand U1814 (N_1814,N_1618,N_1544);
xnor U1815 (N_1815,N_1747,N_1328);
nand U1816 (N_1816,N_1699,N_1634);
nand U1817 (N_1817,N_1635,N_1702);
and U1818 (N_1818,N_1650,N_1714);
nor U1819 (N_1819,N_1668,N_1704);
xnor U1820 (N_1820,N_1603,N_1608);
xnor U1821 (N_1821,N_1569,N_1601);
or U1822 (N_1822,N_1728,In_474);
nand U1823 (N_1823,N_1612,In_939);
and U1824 (N_1824,N_1454,N_1686);
and U1825 (N_1825,N_595,N_1663);
or U1826 (N_1826,N_1339,N_1729);
and U1827 (N_1827,N_1736,N_1722);
xnor U1828 (N_1828,N_1649,N_1719);
and U1829 (N_1829,N_1673,N_1628);
nand U1830 (N_1830,N_1626,N_1749);
and U1831 (N_1831,N_1648,N_1530);
xnor U1832 (N_1832,N_1681,N_1506);
or U1833 (N_1833,N_1713,N_1431);
or U1834 (N_1834,N_1711,N_1487);
nor U1835 (N_1835,N_1705,N_1674);
nand U1836 (N_1836,In_1527,N_1752);
nand U1837 (N_1837,N_1707,N_1724);
nor U1838 (N_1838,N_1658,In_158);
or U1839 (N_1839,N_1619,N_1625);
xor U1840 (N_1840,N_1693,N_1440);
nor U1841 (N_1841,N_1735,N_1676);
and U1842 (N_1842,N_1631,N_1703);
nor U1843 (N_1843,N_1127,N_1651);
or U1844 (N_1844,N_1076,N_1751);
or U1845 (N_1845,N_1727,N_1708);
nor U1846 (N_1846,N_1665,N_1754);
xnor U1847 (N_1847,N_1695,N_1604);
nor U1848 (N_1848,N_1685,N_1639);
or U1849 (N_1849,In_1622,N_1492);
xnor U1850 (N_1850,N_1740,N_1638);
nand U1851 (N_1851,N_1725,N_1666);
or U1852 (N_1852,N_341,N_1670);
and U1853 (N_1853,N_1690,N_1675);
xnor U1854 (N_1854,N_1610,N_1609);
or U1855 (N_1855,N_1746,N_1287);
nor U1856 (N_1856,N_1206,N_1720);
or U1857 (N_1857,N_1677,N_1613);
or U1858 (N_1858,N_1688,N_708);
and U1859 (N_1859,N_1445,N_1646);
nor U1860 (N_1860,N_1511,N_1683);
xor U1861 (N_1861,N_1715,N_1733);
nand U1862 (N_1862,N_1737,N_1647);
or U1863 (N_1863,N_1411,N_1274);
or U1864 (N_1864,N_1753,N_1710);
and U1865 (N_1865,N_1636,N_1682);
nand U1866 (N_1866,N_1621,N_1731);
and U1867 (N_1867,In_1554,N_1617);
and U1868 (N_1868,N_1667,N_1755);
xnor U1869 (N_1869,N_1684,N_1553);
and U1870 (N_1870,N_1543,N_1459);
or U1871 (N_1871,N_1694,N_1614);
nor U1872 (N_1872,N_1691,N_1679);
xor U1873 (N_1873,N_1338,N_1640);
or U1874 (N_1874,N_1176,N_1267);
or U1875 (N_1875,N_1643,N_1745);
nor U1876 (N_1876,N_1637,N_1602);
nand U1877 (N_1877,N_1697,N_1299);
nand U1878 (N_1878,N_1739,N_1605);
xor U1879 (N_1879,N_1568,N_1557);
nor U1880 (N_1880,N_1445,N_1706);
and U1881 (N_1881,N_1602,N_822);
nand U1882 (N_1882,N_1679,N_1683);
and U1883 (N_1883,N_1759,N_1735);
nand U1884 (N_1884,N_1607,N_1690);
and U1885 (N_1885,N_1659,N_1711);
xor U1886 (N_1886,N_1446,N_1612);
nor U1887 (N_1887,N_1681,In_158);
and U1888 (N_1888,N_708,N_1679);
nor U1889 (N_1889,N_1511,In_1184);
and U1890 (N_1890,N_1710,N_1659);
and U1891 (N_1891,N_1608,In_474);
nor U1892 (N_1892,In_166,N_1647);
nor U1893 (N_1893,N_1636,N_1722);
or U1894 (N_1894,N_1705,N_1267);
and U1895 (N_1895,N_1757,N_1729);
nor U1896 (N_1896,N_1674,N_1271);
xor U1897 (N_1897,N_1326,N_1752);
nor U1898 (N_1898,In_1184,In_150);
and U1899 (N_1899,In_474,N_1082);
or U1900 (N_1900,N_1411,N_1487);
nor U1901 (N_1901,N_1626,N_1467);
nand U1902 (N_1902,N_661,N_396);
xor U1903 (N_1903,In_1527,N_1687);
xor U1904 (N_1904,N_1744,N_1127);
nor U1905 (N_1905,N_1737,N_1699);
nand U1906 (N_1906,N_727,N_1593);
nor U1907 (N_1907,N_1720,N_1618);
and U1908 (N_1908,N_1301,N_1338);
and U1909 (N_1909,N_1609,N_1481);
and U1910 (N_1910,N_1039,N_1714);
or U1911 (N_1911,N_727,N_1657);
and U1912 (N_1912,N_1753,N_1715);
nor U1913 (N_1913,N_1544,N_1697);
nand U1914 (N_1914,N_1370,N_1431);
nor U1915 (N_1915,N_1735,N_1662);
xor U1916 (N_1916,N_1693,N_1608);
nor U1917 (N_1917,In_804,In_158);
xnor U1918 (N_1918,N_1672,N_1709);
nand U1919 (N_1919,N_1626,N_1663);
or U1920 (N_1920,N_1805,N_1840);
xnor U1921 (N_1921,N_1830,N_1896);
and U1922 (N_1922,N_1795,N_1774);
nor U1923 (N_1923,N_1890,N_1845);
or U1924 (N_1924,N_1772,N_1867);
nand U1925 (N_1925,N_1898,N_1823);
or U1926 (N_1926,N_1869,N_1891);
nand U1927 (N_1927,N_1858,N_1872);
nand U1928 (N_1928,N_1894,N_1905);
and U1929 (N_1929,N_1783,N_1770);
nor U1930 (N_1930,N_1849,N_1822);
and U1931 (N_1931,N_1819,N_1800);
nor U1932 (N_1932,N_1818,N_1862);
xor U1933 (N_1933,N_1804,N_1900);
xnor U1934 (N_1934,N_1850,N_1885);
nand U1935 (N_1935,N_1766,N_1827);
nor U1936 (N_1936,N_1812,N_1919);
and U1937 (N_1937,N_1832,N_1851);
nand U1938 (N_1938,N_1767,N_1917);
nor U1939 (N_1939,N_1776,N_1874);
and U1940 (N_1940,N_1848,N_1870);
nand U1941 (N_1941,N_1771,N_1881);
nor U1942 (N_1942,N_1834,N_1857);
and U1943 (N_1943,N_1781,N_1798);
nor U1944 (N_1944,N_1908,N_1789);
or U1945 (N_1945,N_1793,N_1824);
and U1946 (N_1946,N_1906,N_1790);
nand U1947 (N_1947,N_1765,N_1763);
nor U1948 (N_1948,N_1846,N_1784);
xnor U1949 (N_1949,N_1762,N_1809);
nor U1950 (N_1950,N_1817,N_1909);
or U1951 (N_1951,N_1859,N_1841);
nand U1952 (N_1952,N_1785,N_1887);
nand U1953 (N_1953,N_1799,N_1807);
nand U1954 (N_1954,N_1813,N_1820);
or U1955 (N_1955,N_1892,N_1842);
nand U1956 (N_1956,N_1777,N_1878);
or U1957 (N_1957,N_1801,N_1907);
or U1958 (N_1958,N_1914,N_1915);
nand U1959 (N_1959,N_1902,N_1828);
nor U1960 (N_1960,N_1833,N_1856);
xor U1961 (N_1961,N_1837,N_1911);
nand U1962 (N_1962,N_1791,N_1860);
and U1963 (N_1963,N_1883,N_1855);
nor U1964 (N_1964,N_1916,N_1844);
nand U1965 (N_1965,N_1853,N_1880);
nor U1966 (N_1966,N_1904,N_1780);
nor U1967 (N_1967,N_1864,N_1810);
nor U1968 (N_1968,N_1893,N_1821);
or U1969 (N_1969,N_1792,N_1873);
xnor U1970 (N_1970,N_1879,N_1788);
or U1971 (N_1971,N_1760,N_1811);
or U1972 (N_1972,N_1768,N_1838);
xnor U1973 (N_1973,N_1847,N_1852);
nand U1974 (N_1974,N_1871,N_1786);
xor U1975 (N_1975,N_1787,N_1836);
and U1976 (N_1976,N_1861,N_1875);
nor U1977 (N_1977,N_1884,N_1897);
nor U1978 (N_1978,N_1796,N_1773);
nand U1979 (N_1979,N_1865,N_1816);
nand U1980 (N_1980,N_1808,N_1901);
xnor U1981 (N_1981,N_1829,N_1854);
nand U1982 (N_1982,N_1888,N_1782);
or U1983 (N_1983,N_1903,N_1803);
nand U1984 (N_1984,N_1868,N_1826);
and U1985 (N_1985,N_1882,N_1912);
and U1986 (N_1986,N_1876,N_1797);
nand U1987 (N_1987,N_1910,N_1831);
and U1988 (N_1988,N_1825,N_1835);
and U1989 (N_1989,N_1761,N_1764);
and U1990 (N_1990,N_1806,N_1899);
nand U1991 (N_1991,N_1886,N_1913);
xor U1992 (N_1992,N_1839,N_1863);
xor U1993 (N_1993,N_1779,N_1775);
xor U1994 (N_1994,N_1889,N_1802);
xor U1995 (N_1995,N_1769,N_1814);
xnor U1996 (N_1996,N_1918,N_1877);
nor U1997 (N_1997,N_1895,N_1866);
nand U1998 (N_1998,N_1843,N_1778);
nor U1999 (N_1999,N_1815,N_1794);
or U2000 (N_2000,N_1863,N_1780);
xor U2001 (N_2001,N_1850,N_1884);
nor U2002 (N_2002,N_1815,N_1801);
nand U2003 (N_2003,N_1914,N_1846);
nand U2004 (N_2004,N_1820,N_1889);
nand U2005 (N_2005,N_1806,N_1767);
nor U2006 (N_2006,N_1855,N_1811);
and U2007 (N_2007,N_1877,N_1777);
or U2008 (N_2008,N_1881,N_1764);
xnor U2009 (N_2009,N_1784,N_1794);
nor U2010 (N_2010,N_1829,N_1883);
or U2011 (N_2011,N_1802,N_1820);
nand U2012 (N_2012,N_1840,N_1789);
or U2013 (N_2013,N_1820,N_1862);
and U2014 (N_2014,N_1911,N_1782);
or U2015 (N_2015,N_1814,N_1810);
and U2016 (N_2016,N_1791,N_1802);
nor U2017 (N_2017,N_1872,N_1822);
nor U2018 (N_2018,N_1896,N_1762);
nor U2019 (N_2019,N_1836,N_1764);
and U2020 (N_2020,N_1763,N_1841);
nor U2021 (N_2021,N_1860,N_1767);
or U2022 (N_2022,N_1844,N_1771);
and U2023 (N_2023,N_1814,N_1870);
nor U2024 (N_2024,N_1780,N_1828);
nor U2025 (N_2025,N_1837,N_1891);
nand U2026 (N_2026,N_1903,N_1831);
or U2027 (N_2027,N_1883,N_1881);
and U2028 (N_2028,N_1908,N_1775);
nor U2029 (N_2029,N_1874,N_1908);
and U2030 (N_2030,N_1786,N_1826);
or U2031 (N_2031,N_1794,N_1839);
nand U2032 (N_2032,N_1889,N_1902);
and U2033 (N_2033,N_1811,N_1875);
xnor U2034 (N_2034,N_1828,N_1896);
nand U2035 (N_2035,N_1902,N_1904);
nand U2036 (N_2036,N_1855,N_1911);
and U2037 (N_2037,N_1907,N_1850);
and U2038 (N_2038,N_1763,N_1857);
nor U2039 (N_2039,N_1867,N_1836);
nor U2040 (N_2040,N_1853,N_1865);
or U2041 (N_2041,N_1914,N_1810);
nor U2042 (N_2042,N_1833,N_1869);
or U2043 (N_2043,N_1899,N_1761);
or U2044 (N_2044,N_1839,N_1792);
and U2045 (N_2045,N_1906,N_1771);
nor U2046 (N_2046,N_1805,N_1783);
and U2047 (N_2047,N_1908,N_1814);
or U2048 (N_2048,N_1883,N_1813);
nor U2049 (N_2049,N_1905,N_1811);
nand U2050 (N_2050,N_1894,N_1791);
or U2051 (N_2051,N_1764,N_1827);
or U2052 (N_2052,N_1785,N_1899);
and U2053 (N_2053,N_1861,N_1766);
nand U2054 (N_2054,N_1860,N_1867);
xor U2055 (N_2055,N_1877,N_1917);
xor U2056 (N_2056,N_1762,N_1777);
xnor U2057 (N_2057,N_1871,N_1909);
xor U2058 (N_2058,N_1880,N_1918);
nor U2059 (N_2059,N_1880,N_1899);
or U2060 (N_2060,N_1819,N_1804);
nand U2061 (N_2061,N_1890,N_1833);
xor U2062 (N_2062,N_1905,N_1804);
nand U2063 (N_2063,N_1842,N_1835);
or U2064 (N_2064,N_1868,N_1885);
or U2065 (N_2065,N_1822,N_1893);
and U2066 (N_2066,N_1903,N_1867);
nand U2067 (N_2067,N_1844,N_1762);
nand U2068 (N_2068,N_1893,N_1827);
nor U2069 (N_2069,N_1906,N_1853);
nand U2070 (N_2070,N_1824,N_1787);
xnor U2071 (N_2071,N_1872,N_1806);
or U2072 (N_2072,N_1831,N_1851);
xor U2073 (N_2073,N_1792,N_1774);
or U2074 (N_2074,N_1853,N_1881);
nor U2075 (N_2075,N_1833,N_1787);
xnor U2076 (N_2076,N_1815,N_1882);
or U2077 (N_2077,N_1781,N_1822);
and U2078 (N_2078,N_1862,N_1873);
xor U2079 (N_2079,N_1838,N_1852);
or U2080 (N_2080,N_1938,N_1993);
nand U2081 (N_2081,N_1975,N_2012);
nor U2082 (N_2082,N_1948,N_1969);
xnor U2083 (N_2083,N_2010,N_2040);
xnor U2084 (N_2084,N_2032,N_1956);
nor U2085 (N_2085,N_1924,N_1953);
or U2086 (N_2086,N_2076,N_1958);
and U2087 (N_2087,N_1921,N_2042);
xor U2088 (N_2088,N_1964,N_1951);
and U2089 (N_2089,N_1941,N_2072);
nor U2090 (N_2090,N_2051,N_2035);
or U2091 (N_2091,N_2023,N_1926);
or U2092 (N_2092,N_1957,N_2068);
or U2093 (N_2093,N_1949,N_1954);
nand U2094 (N_2094,N_2027,N_1986);
and U2095 (N_2095,N_1991,N_2052);
or U2096 (N_2096,N_1945,N_2043);
nor U2097 (N_2097,N_2011,N_2046);
nand U2098 (N_2098,N_1947,N_2029);
nand U2099 (N_2099,N_2015,N_1929);
nand U2100 (N_2100,N_1989,N_2039);
xnor U2101 (N_2101,N_1960,N_1950);
xnor U2102 (N_2102,N_2031,N_2008);
nand U2103 (N_2103,N_2077,N_2013);
and U2104 (N_2104,N_1979,N_2048);
or U2105 (N_2105,N_1976,N_1928);
xor U2106 (N_2106,N_2073,N_1982);
or U2107 (N_2107,N_2007,N_2054);
or U2108 (N_2108,N_2030,N_2071);
and U2109 (N_2109,N_2066,N_2003);
or U2110 (N_2110,N_2049,N_1981);
nor U2111 (N_2111,N_2026,N_2056);
and U2112 (N_2112,N_2070,N_2033);
nor U2113 (N_2113,N_1971,N_1999);
or U2114 (N_2114,N_2079,N_2057);
nor U2115 (N_2115,N_1978,N_2037);
nand U2116 (N_2116,N_2050,N_1946);
nor U2117 (N_2117,N_2047,N_2059);
nand U2118 (N_2118,N_1988,N_1931);
xor U2119 (N_2119,N_2038,N_2065);
or U2120 (N_2120,N_1955,N_1968);
xor U2121 (N_2121,N_1962,N_1992);
nand U2122 (N_2122,N_1972,N_2062);
or U2123 (N_2123,N_2014,N_1977);
nor U2124 (N_2124,N_1923,N_1998);
or U2125 (N_2125,N_2074,N_2058);
and U2126 (N_2126,N_1997,N_1967);
nand U2127 (N_2127,N_1922,N_1996);
or U2128 (N_2128,N_1980,N_1987);
nand U2129 (N_2129,N_2067,N_2020);
or U2130 (N_2130,N_2028,N_2024);
xor U2131 (N_2131,N_1952,N_1934);
or U2132 (N_2132,N_1974,N_2069);
nand U2133 (N_2133,N_2016,N_1963);
nand U2134 (N_2134,N_2022,N_1984);
and U2135 (N_2135,N_2002,N_1942);
or U2136 (N_2136,N_2044,N_2006);
xnor U2137 (N_2137,N_1995,N_1920);
xor U2138 (N_2138,N_2078,N_2018);
and U2139 (N_2139,N_1965,N_2053);
and U2140 (N_2140,N_1994,N_1940);
nor U2141 (N_2141,N_2055,N_2000);
xor U2142 (N_2142,N_1927,N_1930);
and U2143 (N_2143,N_2021,N_1936);
nor U2144 (N_2144,N_2041,N_2001);
or U2145 (N_2145,N_2075,N_1935);
nand U2146 (N_2146,N_1933,N_2017);
nand U2147 (N_2147,N_1966,N_1944);
or U2148 (N_2148,N_2009,N_2045);
nor U2149 (N_2149,N_1970,N_1939);
and U2150 (N_2150,N_2060,N_1943);
nor U2151 (N_2151,N_1925,N_1961);
and U2152 (N_2152,N_1937,N_1932);
and U2153 (N_2153,N_1983,N_2025);
and U2154 (N_2154,N_2004,N_2019);
nand U2155 (N_2155,N_2036,N_2061);
xnor U2156 (N_2156,N_2005,N_1990);
xnor U2157 (N_2157,N_2063,N_1973);
nor U2158 (N_2158,N_2064,N_1985);
nor U2159 (N_2159,N_1959,N_2034);
or U2160 (N_2160,N_2007,N_2050);
or U2161 (N_2161,N_1979,N_2020);
xor U2162 (N_2162,N_1986,N_1920);
or U2163 (N_2163,N_1971,N_2026);
or U2164 (N_2164,N_1953,N_2019);
and U2165 (N_2165,N_1978,N_2049);
or U2166 (N_2166,N_2025,N_2076);
xnor U2167 (N_2167,N_2026,N_2006);
nor U2168 (N_2168,N_1990,N_1978);
nor U2169 (N_2169,N_1995,N_2076);
or U2170 (N_2170,N_1979,N_2044);
and U2171 (N_2171,N_2070,N_1928);
or U2172 (N_2172,N_2016,N_2002);
or U2173 (N_2173,N_2035,N_2031);
xor U2174 (N_2174,N_2079,N_1947);
nor U2175 (N_2175,N_2016,N_1972);
and U2176 (N_2176,N_1991,N_2013);
nor U2177 (N_2177,N_1940,N_1935);
nand U2178 (N_2178,N_2033,N_1965);
or U2179 (N_2179,N_2072,N_1943);
and U2180 (N_2180,N_2068,N_1942);
nand U2181 (N_2181,N_1960,N_2032);
and U2182 (N_2182,N_2009,N_2031);
nand U2183 (N_2183,N_2022,N_1987);
xor U2184 (N_2184,N_1957,N_1929);
nor U2185 (N_2185,N_2039,N_2073);
or U2186 (N_2186,N_2034,N_2079);
nand U2187 (N_2187,N_2025,N_1958);
nand U2188 (N_2188,N_2022,N_2015);
and U2189 (N_2189,N_2063,N_1978);
or U2190 (N_2190,N_2073,N_2076);
xnor U2191 (N_2191,N_2064,N_2003);
or U2192 (N_2192,N_2079,N_2002);
xnor U2193 (N_2193,N_1954,N_2009);
and U2194 (N_2194,N_2000,N_1954);
xnor U2195 (N_2195,N_1935,N_1963);
and U2196 (N_2196,N_1930,N_2034);
nor U2197 (N_2197,N_1984,N_2008);
nand U2198 (N_2198,N_1943,N_1925);
nor U2199 (N_2199,N_1957,N_2011);
and U2200 (N_2200,N_2055,N_1937);
nand U2201 (N_2201,N_1966,N_1931);
xnor U2202 (N_2202,N_2077,N_1974);
and U2203 (N_2203,N_1961,N_1996);
or U2204 (N_2204,N_1939,N_1988);
nand U2205 (N_2205,N_1972,N_1933);
and U2206 (N_2206,N_2026,N_2052);
and U2207 (N_2207,N_2059,N_1928);
nand U2208 (N_2208,N_2059,N_2036);
and U2209 (N_2209,N_1998,N_2012);
or U2210 (N_2210,N_2010,N_1929);
nand U2211 (N_2211,N_2017,N_1939);
and U2212 (N_2212,N_1990,N_1979);
xor U2213 (N_2213,N_2056,N_1954);
nand U2214 (N_2214,N_2076,N_2034);
and U2215 (N_2215,N_2046,N_1936);
nand U2216 (N_2216,N_2069,N_2074);
nor U2217 (N_2217,N_1978,N_2042);
xor U2218 (N_2218,N_1931,N_2037);
xor U2219 (N_2219,N_1922,N_2052);
or U2220 (N_2220,N_2051,N_2014);
nor U2221 (N_2221,N_2034,N_1943);
or U2222 (N_2222,N_2044,N_1953);
and U2223 (N_2223,N_1960,N_2028);
nor U2224 (N_2224,N_1947,N_2028);
nor U2225 (N_2225,N_1984,N_2031);
xor U2226 (N_2226,N_1921,N_1949);
and U2227 (N_2227,N_2007,N_2016);
or U2228 (N_2228,N_2004,N_1933);
nand U2229 (N_2229,N_2044,N_2070);
xor U2230 (N_2230,N_1939,N_2035);
xnor U2231 (N_2231,N_1935,N_2052);
xor U2232 (N_2232,N_2050,N_2018);
and U2233 (N_2233,N_1968,N_1941);
nor U2234 (N_2234,N_2067,N_2056);
nor U2235 (N_2235,N_2058,N_2046);
xor U2236 (N_2236,N_1920,N_2054);
or U2237 (N_2237,N_2016,N_2049);
or U2238 (N_2238,N_2025,N_2001);
nor U2239 (N_2239,N_2011,N_1944);
xor U2240 (N_2240,N_2191,N_2234);
xor U2241 (N_2241,N_2207,N_2202);
or U2242 (N_2242,N_2120,N_2105);
xor U2243 (N_2243,N_2224,N_2166);
xor U2244 (N_2244,N_2170,N_2082);
xor U2245 (N_2245,N_2216,N_2171);
xor U2246 (N_2246,N_2092,N_2194);
nor U2247 (N_2247,N_2142,N_2238);
nor U2248 (N_2248,N_2156,N_2165);
nor U2249 (N_2249,N_2237,N_2198);
nor U2250 (N_2250,N_2160,N_2192);
nor U2251 (N_2251,N_2154,N_2175);
nor U2252 (N_2252,N_2152,N_2102);
or U2253 (N_2253,N_2219,N_2090);
nand U2254 (N_2254,N_2086,N_2201);
or U2255 (N_2255,N_2123,N_2239);
nand U2256 (N_2256,N_2195,N_2108);
nor U2257 (N_2257,N_2188,N_2163);
nand U2258 (N_2258,N_2081,N_2126);
or U2259 (N_2259,N_2098,N_2227);
and U2260 (N_2260,N_2214,N_2184);
or U2261 (N_2261,N_2099,N_2114);
nor U2262 (N_2262,N_2230,N_2159);
and U2263 (N_2263,N_2233,N_2168);
and U2264 (N_2264,N_2180,N_2228);
xnor U2265 (N_2265,N_2130,N_2220);
nand U2266 (N_2266,N_2183,N_2193);
nor U2267 (N_2267,N_2179,N_2203);
or U2268 (N_2268,N_2136,N_2093);
nor U2269 (N_2269,N_2147,N_2174);
xor U2270 (N_2270,N_2199,N_2218);
xor U2271 (N_2271,N_2118,N_2209);
xor U2272 (N_2272,N_2104,N_2155);
xnor U2273 (N_2273,N_2149,N_2217);
and U2274 (N_2274,N_2181,N_2131);
nand U2275 (N_2275,N_2101,N_2221);
nand U2276 (N_2276,N_2117,N_2119);
or U2277 (N_2277,N_2177,N_2084);
xnor U2278 (N_2278,N_2088,N_2097);
nor U2279 (N_2279,N_2129,N_2185);
nand U2280 (N_2280,N_2158,N_2124);
xor U2281 (N_2281,N_2127,N_2205);
or U2282 (N_2282,N_2215,N_2137);
nand U2283 (N_2283,N_2167,N_2115);
nand U2284 (N_2284,N_2135,N_2206);
xor U2285 (N_2285,N_2133,N_2080);
nand U2286 (N_2286,N_2157,N_2189);
or U2287 (N_2287,N_2107,N_2197);
or U2288 (N_2288,N_2094,N_2146);
nor U2289 (N_2289,N_2103,N_2116);
or U2290 (N_2290,N_2161,N_2208);
xor U2291 (N_2291,N_2132,N_2169);
and U2292 (N_2292,N_2210,N_2083);
or U2293 (N_2293,N_2187,N_2196);
xor U2294 (N_2294,N_2148,N_2178);
nor U2295 (N_2295,N_2091,N_2113);
or U2296 (N_2296,N_2225,N_2134);
nand U2297 (N_2297,N_2235,N_2204);
nand U2298 (N_2298,N_2222,N_2186);
and U2299 (N_2299,N_2150,N_2176);
or U2300 (N_2300,N_2138,N_2164);
nand U2301 (N_2301,N_2125,N_2121);
nor U2302 (N_2302,N_2085,N_2139);
or U2303 (N_2303,N_2212,N_2190);
nand U2304 (N_2304,N_2106,N_2096);
and U2305 (N_2305,N_2109,N_2143);
nand U2306 (N_2306,N_2144,N_2110);
xor U2307 (N_2307,N_2236,N_2100);
and U2308 (N_2308,N_2229,N_2153);
and U2309 (N_2309,N_2122,N_2226);
or U2310 (N_2310,N_2182,N_2213);
xnor U2311 (N_2311,N_2145,N_2128);
xor U2312 (N_2312,N_2232,N_2162);
xor U2313 (N_2313,N_2172,N_2231);
nand U2314 (N_2314,N_2200,N_2140);
and U2315 (N_2315,N_2173,N_2112);
nand U2316 (N_2316,N_2151,N_2089);
and U2317 (N_2317,N_2211,N_2223);
nor U2318 (N_2318,N_2141,N_2087);
and U2319 (N_2319,N_2095,N_2111);
and U2320 (N_2320,N_2138,N_2154);
and U2321 (N_2321,N_2103,N_2223);
and U2322 (N_2322,N_2148,N_2231);
xor U2323 (N_2323,N_2207,N_2080);
nor U2324 (N_2324,N_2117,N_2128);
nor U2325 (N_2325,N_2226,N_2157);
nand U2326 (N_2326,N_2217,N_2092);
xor U2327 (N_2327,N_2233,N_2087);
nor U2328 (N_2328,N_2087,N_2132);
and U2329 (N_2329,N_2093,N_2159);
nor U2330 (N_2330,N_2199,N_2150);
xor U2331 (N_2331,N_2100,N_2082);
nand U2332 (N_2332,N_2183,N_2167);
nor U2333 (N_2333,N_2232,N_2196);
nand U2334 (N_2334,N_2147,N_2127);
nand U2335 (N_2335,N_2217,N_2126);
xor U2336 (N_2336,N_2110,N_2098);
and U2337 (N_2337,N_2150,N_2204);
or U2338 (N_2338,N_2186,N_2144);
and U2339 (N_2339,N_2191,N_2107);
or U2340 (N_2340,N_2179,N_2222);
xnor U2341 (N_2341,N_2188,N_2191);
or U2342 (N_2342,N_2083,N_2121);
and U2343 (N_2343,N_2163,N_2210);
nand U2344 (N_2344,N_2100,N_2163);
xnor U2345 (N_2345,N_2201,N_2175);
nor U2346 (N_2346,N_2117,N_2228);
and U2347 (N_2347,N_2097,N_2149);
or U2348 (N_2348,N_2185,N_2237);
xor U2349 (N_2349,N_2197,N_2201);
nand U2350 (N_2350,N_2210,N_2167);
and U2351 (N_2351,N_2213,N_2107);
nand U2352 (N_2352,N_2182,N_2143);
nor U2353 (N_2353,N_2158,N_2104);
and U2354 (N_2354,N_2217,N_2165);
nor U2355 (N_2355,N_2144,N_2131);
nor U2356 (N_2356,N_2202,N_2217);
xor U2357 (N_2357,N_2084,N_2183);
and U2358 (N_2358,N_2211,N_2109);
nor U2359 (N_2359,N_2110,N_2196);
xnor U2360 (N_2360,N_2148,N_2144);
nor U2361 (N_2361,N_2151,N_2138);
and U2362 (N_2362,N_2219,N_2230);
xnor U2363 (N_2363,N_2147,N_2149);
nand U2364 (N_2364,N_2219,N_2234);
nor U2365 (N_2365,N_2119,N_2125);
nand U2366 (N_2366,N_2125,N_2185);
nor U2367 (N_2367,N_2083,N_2128);
and U2368 (N_2368,N_2137,N_2181);
and U2369 (N_2369,N_2133,N_2094);
or U2370 (N_2370,N_2152,N_2162);
or U2371 (N_2371,N_2141,N_2232);
and U2372 (N_2372,N_2160,N_2150);
nand U2373 (N_2373,N_2141,N_2215);
xor U2374 (N_2374,N_2189,N_2160);
and U2375 (N_2375,N_2126,N_2183);
xnor U2376 (N_2376,N_2087,N_2101);
nor U2377 (N_2377,N_2100,N_2147);
xor U2378 (N_2378,N_2191,N_2200);
nand U2379 (N_2379,N_2119,N_2239);
nand U2380 (N_2380,N_2200,N_2206);
xnor U2381 (N_2381,N_2127,N_2237);
and U2382 (N_2382,N_2222,N_2100);
nor U2383 (N_2383,N_2145,N_2224);
nor U2384 (N_2384,N_2232,N_2139);
nor U2385 (N_2385,N_2133,N_2157);
nand U2386 (N_2386,N_2091,N_2126);
xnor U2387 (N_2387,N_2218,N_2189);
and U2388 (N_2388,N_2162,N_2225);
nand U2389 (N_2389,N_2091,N_2120);
and U2390 (N_2390,N_2215,N_2090);
and U2391 (N_2391,N_2097,N_2209);
nand U2392 (N_2392,N_2212,N_2218);
and U2393 (N_2393,N_2146,N_2117);
nor U2394 (N_2394,N_2084,N_2152);
xor U2395 (N_2395,N_2119,N_2122);
nor U2396 (N_2396,N_2233,N_2085);
xor U2397 (N_2397,N_2108,N_2161);
or U2398 (N_2398,N_2236,N_2090);
nor U2399 (N_2399,N_2186,N_2130);
or U2400 (N_2400,N_2318,N_2240);
nand U2401 (N_2401,N_2287,N_2372);
nand U2402 (N_2402,N_2357,N_2360);
and U2403 (N_2403,N_2380,N_2307);
nand U2404 (N_2404,N_2362,N_2366);
or U2405 (N_2405,N_2286,N_2387);
nand U2406 (N_2406,N_2273,N_2323);
nor U2407 (N_2407,N_2399,N_2359);
or U2408 (N_2408,N_2330,N_2292);
nand U2409 (N_2409,N_2276,N_2332);
and U2410 (N_2410,N_2396,N_2316);
and U2411 (N_2411,N_2314,N_2383);
nor U2412 (N_2412,N_2294,N_2302);
nor U2413 (N_2413,N_2335,N_2310);
and U2414 (N_2414,N_2348,N_2271);
and U2415 (N_2415,N_2326,N_2261);
nor U2416 (N_2416,N_2245,N_2241);
or U2417 (N_2417,N_2319,N_2244);
nor U2418 (N_2418,N_2279,N_2277);
and U2419 (N_2419,N_2263,N_2290);
xnor U2420 (N_2420,N_2243,N_2392);
xor U2421 (N_2421,N_2376,N_2375);
nand U2422 (N_2422,N_2338,N_2252);
or U2423 (N_2423,N_2378,N_2353);
nor U2424 (N_2424,N_2299,N_2272);
or U2425 (N_2425,N_2345,N_2343);
xnor U2426 (N_2426,N_2363,N_2374);
nand U2427 (N_2427,N_2305,N_2367);
xnor U2428 (N_2428,N_2331,N_2295);
nand U2429 (N_2429,N_2262,N_2265);
or U2430 (N_2430,N_2312,N_2341);
and U2431 (N_2431,N_2301,N_2354);
or U2432 (N_2432,N_2300,N_2311);
nor U2433 (N_2433,N_2266,N_2355);
or U2434 (N_2434,N_2267,N_2282);
or U2435 (N_2435,N_2368,N_2306);
nor U2436 (N_2436,N_2291,N_2296);
or U2437 (N_2437,N_2303,N_2391);
nor U2438 (N_2438,N_2395,N_2248);
or U2439 (N_2439,N_2242,N_2346);
nor U2440 (N_2440,N_2397,N_2336);
nand U2441 (N_2441,N_2344,N_2390);
or U2442 (N_2442,N_2264,N_2351);
xor U2443 (N_2443,N_2246,N_2322);
and U2444 (N_2444,N_2356,N_2280);
and U2445 (N_2445,N_2373,N_2254);
or U2446 (N_2446,N_2347,N_2281);
xor U2447 (N_2447,N_2274,N_2329);
or U2448 (N_2448,N_2289,N_2389);
or U2449 (N_2449,N_2258,N_2257);
nor U2450 (N_2450,N_2337,N_2384);
or U2451 (N_2451,N_2255,N_2269);
nand U2452 (N_2452,N_2385,N_2249);
nor U2453 (N_2453,N_2358,N_2365);
nor U2454 (N_2454,N_2253,N_2361);
or U2455 (N_2455,N_2352,N_2304);
nor U2456 (N_2456,N_2340,N_2381);
nor U2457 (N_2457,N_2283,N_2315);
nand U2458 (N_2458,N_2298,N_2278);
nand U2459 (N_2459,N_2328,N_2275);
or U2460 (N_2460,N_2398,N_2270);
and U2461 (N_2461,N_2250,N_2268);
nor U2462 (N_2462,N_2386,N_2317);
nor U2463 (N_2463,N_2325,N_2393);
nor U2464 (N_2464,N_2260,N_2288);
nor U2465 (N_2465,N_2327,N_2364);
xnor U2466 (N_2466,N_2394,N_2382);
xor U2467 (N_2467,N_2321,N_2350);
nand U2468 (N_2468,N_2339,N_2247);
and U2469 (N_2469,N_2334,N_2333);
or U2470 (N_2470,N_2284,N_2308);
or U2471 (N_2471,N_2297,N_2256);
nand U2472 (N_2472,N_2251,N_2349);
or U2473 (N_2473,N_2377,N_2371);
or U2474 (N_2474,N_2259,N_2379);
and U2475 (N_2475,N_2313,N_2309);
nor U2476 (N_2476,N_2370,N_2388);
and U2477 (N_2477,N_2320,N_2342);
nor U2478 (N_2478,N_2285,N_2324);
nor U2479 (N_2479,N_2369,N_2293);
or U2480 (N_2480,N_2325,N_2293);
or U2481 (N_2481,N_2284,N_2292);
xor U2482 (N_2482,N_2394,N_2333);
or U2483 (N_2483,N_2269,N_2348);
xnor U2484 (N_2484,N_2264,N_2337);
or U2485 (N_2485,N_2263,N_2387);
nand U2486 (N_2486,N_2357,N_2327);
or U2487 (N_2487,N_2265,N_2345);
or U2488 (N_2488,N_2281,N_2360);
and U2489 (N_2489,N_2373,N_2243);
nand U2490 (N_2490,N_2317,N_2240);
or U2491 (N_2491,N_2343,N_2257);
nor U2492 (N_2492,N_2318,N_2331);
nand U2493 (N_2493,N_2353,N_2340);
nand U2494 (N_2494,N_2288,N_2302);
nor U2495 (N_2495,N_2338,N_2279);
and U2496 (N_2496,N_2344,N_2284);
nand U2497 (N_2497,N_2293,N_2305);
nand U2498 (N_2498,N_2250,N_2351);
and U2499 (N_2499,N_2282,N_2342);
and U2500 (N_2500,N_2353,N_2386);
nand U2501 (N_2501,N_2264,N_2389);
xor U2502 (N_2502,N_2329,N_2316);
and U2503 (N_2503,N_2275,N_2374);
or U2504 (N_2504,N_2280,N_2315);
xor U2505 (N_2505,N_2394,N_2395);
nand U2506 (N_2506,N_2320,N_2385);
xor U2507 (N_2507,N_2260,N_2289);
nor U2508 (N_2508,N_2377,N_2290);
nor U2509 (N_2509,N_2270,N_2347);
nor U2510 (N_2510,N_2255,N_2355);
nand U2511 (N_2511,N_2254,N_2379);
nor U2512 (N_2512,N_2284,N_2319);
or U2513 (N_2513,N_2326,N_2387);
xor U2514 (N_2514,N_2271,N_2296);
or U2515 (N_2515,N_2288,N_2305);
and U2516 (N_2516,N_2325,N_2352);
xnor U2517 (N_2517,N_2310,N_2249);
and U2518 (N_2518,N_2359,N_2281);
and U2519 (N_2519,N_2373,N_2316);
or U2520 (N_2520,N_2249,N_2351);
xnor U2521 (N_2521,N_2280,N_2363);
and U2522 (N_2522,N_2297,N_2352);
xnor U2523 (N_2523,N_2309,N_2360);
nand U2524 (N_2524,N_2294,N_2245);
xnor U2525 (N_2525,N_2383,N_2265);
xnor U2526 (N_2526,N_2242,N_2345);
or U2527 (N_2527,N_2300,N_2266);
xor U2528 (N_2528,N_2335,N_2306);
nand U2529 (N_2529,N_2293,N_2254);
nand U2530 (N_2530,N_2382,N_2315);
and U2531 (N_2531,N_2304,N_2351);
and U2532 (N_2532,N_2345,N_2279);
nor U2533 (N_2533,N_2277,N_2312);
nand U2534 (N_2534,N_2275,N_2304);
nor U2535 (N_2535,N_2277,N_2287);
nand U2536 (N_2536,N_2380,N_2324);
nor U2537 (N_2537,N_2347,N_2272);
nor U2538 (N_2538,N_2302,N_2390);
nor U2539 (N_2539,N_2286,N_2278);
and U2540 (N_2540,N_2396,N_2362);
and U2541 (N_2541,N_2315,N_2250);
or U2542 (N_2542,N_2256,N_2282);
or U2543 (N_2543,N_2256,N_2271);
nor U2544 (N_2544,N_2291,N_2277);
nand U2545 (N_2545,N_2302,N_2306);
nand U2546 (N_2546,N_2271,N_2311);
nor U2547 (N_2547,N_2336,N_2367);
nand U2548 (N_2548,N_2397,N_2276);
or U2549 (N_2549,N_2256,N_2390);
nand U2550 (N_2550,N_2396,N_2337);
nand U2551 (N_2551,N_2248,N_2351);
nor U2552 (N_2552,N_2255,N_2396);
xor U2553 (N_2553,N_2391,N_2380);
and U2554 (N_2554,N_2307,N_2376);
nand U2555 (N_2555,N_2348,N_2278);
xnor U2556 (N_2556,N_2321,N_2314);
xor U2557 (N_2557,N_2253,N_2265);
and U2558 (N_2558,N_2381,N_2241);
xor U2559 (N_2559,N_2268,N_2356);
nor U2560 (N_2560,N_2548,N_2464);
or U2561 (N_2561,N_2502,N_2527);
or U2562 (N_2562,N_2495,N_2516);
nand U2563 (N_2563,N_2526,N_2411);
xnor U2564 (N_2564,N_2423,N_2428);
and U2565 (N_2565,N_2446,N_2543);
nand U2566 (N_2566,N_2538,N_2505);
nor U2567 (N_2567,N_2454,N_2449);
xnor U2568 (N_2568,N_2465,N_2555);
xnor U2569 (N_2569,N_2523,N_2457);
and U2570 (N_2570,N_2473,N_2540);
or U2571 (N_2571,N_2458,N_2522);
xor U2572 (N_2572,N_2414,N_2463);
nor U2573 (N_2573,N_2497,N_2453);
and U2574 (N_2574,N_2422,N_2450);
nor U2575 (N_2575,N_2407,N_2421);
nand U2576 (N_2576,N_2503,N_2461);
nor U2577 (N_2577,N_2435,N_2507);
and U2578 (N_2578,N_2438,N_2429);
or U2579 (N_2579,N_2445,N_2460);
nor U2580 (N_2580,N_2425,N_2432);
or U2581 (N_2581,N_2418,N_2529);
nor U2582 (N_2582,N_2536,N_2549);
nor U2583 (N_2583,N_2492,N_2470);
nor U2584 (N_2584,N_2410,N_2535);
or U2585 (N_2585,N_2406,N_2439);
xor U2586 (N_2586,N_2520,N_2525);
or U2587 (N_2587,N_2510,N_2517);
nor U2588 (N_2588,N_2452,N_2403);
nor U2589 (N_2589,N_2466,N_2482);
xnor U2590 (N_2590,N_2559,N_2402);
nand U2591 (N_2591,N_2542,N_2509);
or U2592 (N_2592,N_2534,N_2486);
xnor U2593 (N_2593,N_2551,N_2431);
or U2594 (N_2594,N_2469,N_2400);
nand U2595 (N_2595,N_2413,N_2412);
or U2596 (N_2596,N_2488,N_2485);
xnor U2597 (N_2597,N_2513,N_2480);
and U2598 (N_2598,N_2448,N_2436);
nand U2599 (N_2599,N_2401,N_2496);
and U2600 (N_2600,N_2530,N_2443);
xor U2601 (N_2601,N_2440,N_2408);
nand U2602 (N_2602,N_2471,N_2532);
or U2603 (N_2603,N_2541,N_2478);
xor U2604 (N_2604,N_2444,N_2491);
nand U2605 (N_2605,N_2437,N_2511);
nand U2606 (N_2606,N_2506,N_2524);
or U2607 (N_2607,N_2494,N_2528);
xor U2608 (N_2608,N_2467,N_2420);
and U2609 (N_2609,N_2547,N_2493);
xnor U2610 (N_2610,N_2557,N_2462);
or U2611 (N_2611,N_2531,N_2515);
and U2612 (N_2612,N_2476,N_2424);
nor U2613 (N_2613,N_2427,N_2415);
xnor U2614 (N_2614,N_2405,N_2442);
xnor U2615 (N_2615,N_2416,N_2550);
xnor U2616 (N_2616,N_2498,N_2499);
xnor U2617 (N_2617,N_2426,N_2447);
and U2618 (N_2618,N_2419,N_2459);
or U2619 (N_2619,N_2479,N_2500);
nand U2620 (N_2620,N_2477,N_2451);
xor U2621 (N_2621,N_2556,N_2504);
nor U2622 (N_2622,N_2481,N_2456);
xnor U2623 (N_2623,N_2521,N_2519);
or U2624 (N_2624,N_2518,N_2409);
nand U2625 (N_2625,N_2489,N_2474);
nand U2626 (N_2626,N_2533,N_2558);
and U2627 (N_2627,N_2441,N_2545);
nand U2628 (N_2628,N_2472,N_2514);
and U2629 (N_2629,N_2553,N_2487);
nand U2630 (N_2630,N_2501,N_2554);
nor U2631 (N_2631,N_2552,N_2484);
nand U2632 (N_2632,N_2434,N_2483);
and U2633 (N_2633,N_2468,N_2455);
and U2634 (N_2634,N_2508,N_2544);
xnor U2635 (N_2635,N_2539,N_2512);
or U2636 (N_2636,N_2417,N_2475);
nand U2637 (N_2637,N_2546,N_2537);
nand U2638 (N_2638,N_2490,N_2404);
xnor U2639 (N_2639,N_2430,N_2433);
and U2640 (N_2640,N_2470,N_2435);
xnor U2641 (N_2641,N_2444,N_2471);
and U2642 (N_2642,N_2469,N_2526);
and U2643 (N_2643,N_2467,N_2409);
xor U2644 (N_2644,N_2538,N_2410);
and U2645 (N_2645,N_2505,N_2524);
or U2646 (N_2646,N_2455,N_2555);
and U2647 (N_2647,N_2497,N_2416);
and U2648 (N_2648,N_2417,N_2422);
xor U2649 (N_2649,N_2547,N_2427);
nand U2650 (N_2650,N_2459,N_2514);
nand U2651 (N_2651,N_2450,N_2548);
and U2652 (N_2652,N_2470,N_2432);
and U2653 (N_2653,N_2455,N_2432);
nor U2654 (N_2654,N_2469,N_2454);
and U2655 (N_2655,N_2510,N_2542);
or U2656 (N_2656,N_2434,N_2455);
or U2657 (N_2657,N_2401,N_2457);
nand U2658 (N_2658,N_2450,N_2424);
or U2659 (N_2659,N_2425,N_2405);
or U2660 (N_2660,N_2444,N_2541);
nand U2661 (N_2661,N_2525,N_2433);
nor U2662 (N_2662,N_2447,N_2521);
or U2663 (N_2663,N_2472,N_2441);
nor U2664 (N_2664,N_2450,N_2447);
and U2665 (N_2665,N_2552,N_2519);
nor U2666 (N_2666,N_2405,N_2512);
xnor U2667 (N_2667,N_2415,N_2554);
nor U2668 (N_2668,N_2530,N_2453);
and U2669 (N_2669,N_2491,N_2548);
xor U2670 (N_2670,N_2514,N_2449);
nand U2671 (N_2671,N_2494,N_2400);
and U2672 (N_2672,N_2539,N_2559);
nand U2673 (N_2673,N_2526,N_2437);
or U2674 (N_2674,N_2502,N_2425);
nor U2675 (N_2675,N_2434,N_2482);
xnor U2676 (N_2676,N_2514,N_2465);
or U2677 (N_2677,N_2503,N_2511);
nor U2678 (N_2678,N_2471,N_2473);
or U2679 (N_2679,N_2519,N_2400);
and U2680 (N_2680,N_2408,N_2447);
nand U2681 (N_2681,N_2518,N_2441);
nand U2682 (N_2682,N_2440,N_2452);
nand U2683 (N_2683,N_2422,N_2553);
and U2684 (N_2684,N_2486,N_2449);
nand U2685 (N_2685,N_2410,N_2501);
and U2686 (N_2686,N_2511,N_2509);
nand U2687 (N_2687,N_2464,N_2545);
and U2688 (N_2688,N_2478,N_2414);
nor U2689 (N_2689,N_2418,N_2557);
nor U2690 (N_2690,N_2539,N_2537);
and U2691 (N_2691,N_2487,N_2518);
nor U2692 (N_2692,N_2501,N_2459);
and U2693 (N_2693,N_2508,N_2491);
xor U2694 (N_2694,N_2442,N_2524);
nor U2695 (N_2695,N_2439,N_2506);
nor U2696 (N_2696,N_2412,N_2527);
nand U2697 (N_2697,N_2400,N_2551);
xor U2698 (N_2698,N_2463,N_2443);
nand U2699 (N_2699,N_2502,N_2536);
xnor U2700 (N_2700,N_2482,N_2544);
nand U2701 (N_2701,N_2496,N_2405);
nor U2702 (N_2702,N_2419,N_2557);
nand U2703 (N_2703,N_2439,N_2423);
or U2704 (N_2704,N_2554,N_2506);
nor U2705 (N_2705,N_2509,N_2504);
and U2706 (N_2706,N_2530,N_2415);
xor U2707 (N_2707,N_2508,N_2528);
nand U2708 (N_2708,N_2431,N_2439);
xnor U2709 (N_2709,N_2439,N_2480);
nor U2710 (N_2710,N_2438,N_2410);
xor U2711 (N_2711,N_2413,N_2496);
and U2712 (N_2712,N_2520,N_2439);
and U2713 (N_2713,N_2424,N_2429);
xnor U2714 (N_2714,N_2512,N_2422);
or U2715 (N_2715,N_2433,N_2467);
nor U2716 (N_2716,N_2520,N_2544);
nor U2717 (N_2717,N_2557,N_2440);
xor U2718 (N_2718,N_2409,N_2522);
xor U2719 (N_2719,N_2403,N_2542);
or U2720 (N_2720,N_2592,N_2671);
and U2721 (N_2721,N_2681,N_2589);
nor U2722 (N_2722,N_2673,N_2651);
and U2723 (N_2723,N_2713,N_2698);
or U2724 (N_2724,N_2603,N_2571);
and U2725 (N_2725,N_2628,N_2659);
nor U2726 (N_2726,N_2689,N_2683);
xor U2727 (N_2727,N_2636,N_2601);
and U2728 (N_2728,N_2575,N_2648);
and U2729 (N_2729,N_2703,N_2595);
and U2730 (N_2730,N_2699,N_2570);
nor U2731 (N_2731,N_2604,N_2608);
and U2732 (N_2732,N_2702,N_2690);
nand U2733 (N_2733,N_2582,N_2580);
nor U2734 (N_2734,N_2662,N_2563);
nor U2735 (N_2735,N_2645,N_2630);
xor U2736 (N_2736,N_2694,N_2562);
and U2737 (N_2737,N_2599,N_2632);
nand U2738 (N_2738,N_2717,N_2611);
and U2739 (N_2739,N_2578,N_2586);
xor U2740 (N_2740,N_2684,N_2661);
or U2741 (N_2741,N_2652,N_2682);
nand U2742 (N_2742,N_2711,N_2621);
nand U2743 (N_2743,N_2638,N_2590);
and U2744 (N_2744,N_2685,N_2709);
nor U2745 (N_2745,N_2649,N_2688);
and U2746 (N_2746,N_2719,N_2610);
nor U2747 (N_2747,N_2627,N_2677);
nand U2748 (N_2748,N_2576,N_2680);
and U2749 (N_2749,N_2633,N_2705);
and U2750 (N_2750,N_2697,N_2602);
nor U2751 (N_2751,N_2672,N_2606);
xor U2752 (N_2752,N_2605,N_2568);
and U2753 (N_2753,N_2584,N_2618);
xnor U2754 (N_2754,N_2670,N_2676);
xor U2755 (N_2755,N_2666,N_2566);
xor U2756 (N_2756,N_2612,N_2567);
or U2757 (N_2757,N_2695,N_2643);
nand U2758 (N_2758,N_2667,N_2646);
nor U2759 (N_2759,N_2701,N_2663);
and U2760 (N_2760,N_2565,N_2615);
or U2761 (N_2761,N_2708,N_2686);
or U2762 (N_2762,N_2658,N_2613);
and U2763 (N_2763,N_2640,N_2718);
or U2764 (N_2764,N_2572,N_2642);
or U2765 (N_2765,N_2660,N_2573);
nand U2766 (N_2766,N_2675,N_2707);
nor U2767 (N_2767,N_2692,N_2623);
xor U2768 (N_2768,N_2593,N_2583);
or U2769 (N_2769,N_2609,N_2691);
and U2770 (N_2770,N_2647,N_2664);
nand U2771 (N_2771,N_2594,N_2607);
or U2772 (N_2772,N_2581,N_2600);
xor U2773 (N_2773,N_2579,N_2668);
and U2774 (N_2774,N_2624,N_2631);
nor U2775 (N_2775,N_2696,N_2650);
and U2776 (N_2776,N_2569,N_2588);
nand U2777 (N_2777,N_2679,N_2669);
or U2778 (N_2778,N_2712,N_2641);
or U2779 (N_2779,N_2693,N_2674);
and U2780 (N_2780,N_2564,N_2587);
and U2781 (N_2781,N_2591,N_2619);
and U2782 (N_2782,N_2598,N_2620);
xor U2783 (N_2783,N_2706,N_2596);
and U2784 (N_2784,N_2710,N_2616);
nand U2785 (N_2785,N_2617,N_2629);
nand U2786 (N_2786,N_2635,N_2560);
and U2787 (N_2787,N_2656,N_2655);
or U2788 (N_2788,N_2715,N_2614);
and U2789 (N_2789,N_2678,N_2639);
nand U2790 (N_2790,N_2716,N_2704);
xor U2791 (N_2791,N_2574,N_2687);
nor U2792 (N_2792,N_2597,N_2714);
nand U2793 (N_2793,N_2577,N_2625);
xnor U2794 (N_2794,N_2626,N_2654);
nand U2795 (N_2795,N_2622,N_2637);
xnor U2796 (N_2796,N_2585,N_2644);
and U2797 (N_2797,N_2561,N_2634);
and U2798 (N_2798,N_2700,N_2665);
xor U2799 (N_2799,N_2657,N_2653);
nor U2800 (N_2800,N_2718,N_2666);
xnor U2801 (N_2801,N_2710,N_2591);
xnor U2802 (N_2802,N_2683,N_2595);
and U2803 (N_2803,N_2637,N_2679);
or U2804 (N_2804,N_2645,N_2582);
nor U2805 (N_2805,N_2716,N_2586);
nor U2806 (N_2806,N_2575,N_2645);
and U2807 (N_2807,N_2614,N_2708);
or U2808 (N_2808,N_2601,N_2595);
or U2809 (N_2809,N_2652,N_2591);
or U2810 (N_2810,N_2711,N_2598);
nor U2811 (N_2811,N_2629,N_2646);
or U2812 (N_2812,N_2662,N_2713);
and U2813 (N_2813,N_2594,N_2696);
or U2814 (N_2814,N_2663,N_2649);
or U2815 (N_2815,N_2605,N_2619);
and U2816 (N_2816,N_2651,N_2677);
xor U2817 (N_2817,N_2717,N_2686);
or U2818 (N_2818,N_2627,N_2575);
xor U2819 (N_2819,N_2675,N_2655);
nand U2820 (N_2820,N_2718,N_2698);
or U2821 (N_2821,N_2581,N_2680);
or U2822 (N_2822,N_2674,N_2623);
nand U2823 (N_2823,N_2656,N_2624);
and U2824 (N_2824,N_2638,N_2691);
xor U2825 (N_2825,N_2618,N_2578);
nor U2826 (N_2826,N_2619,N_2696);
and U2827 (N_2827,N_2600,N_2619);
nand U2828 (N_2828,N_2687,N_2588);
or U2829 (N_2829,N_2591,N_2686);
nand U2830 (N_2830,N_2625,N_2693);
and U2831 (N_2831,N_2626,N_2636);
xnor U2832 (N_2832,N_2593,N_2627);
or U2833 (N_2833,N_2576,N_2636);
nor U2834 (N_2834,N_2593,N_2575);
and U2835 (N_2835,N_2650,N_2700);
nand U2836 (N_2836,N_2613,N_2625);
xor U2837 (N_2837,N_2574,N_2701);
nor U2838 (N_2838,N_2568,N_2611);
nand U2839 (N_2839,N_2640,N_2620);
nand U2840 (N_2840,N_2717,N_2624);
nand U2841 (N_2841,N_2642,N_2595);
and U2842 (N_2842,N_2668,N_2652);
and U2843 (N_2843,N_2679,N_2702);
or U2844 (N_2844,N_2680,N_2644);
nand U2845 (N_2845,N_2591,N_2608);
xnor U2846 (N_2846,N_2682,N_2672);
or U2847 (N_2847,N_2692,N_2592);
and U2848 (N_2848,N_2606,N_2653);
or U2849 (N_2849,N_2705,N_2707);
or U2850 (N_2850,N_2594,N_2715);
nand U2851 (N_2851,N_2690,N_2719);
nor U2852 (N_2852,N_2620,N_2623);
or U2853 (N_2853,N_2712,N_2706);
nand U2854 (N_2854,N_2689,N_2567);
nand U2855 (N_2855,N_2586,N_2664);
or U2856 (N_2856,N_2618,N_2600);
xor U2857 (N_2857,N_2602,N_2627);
or U2858 (N_2858,N_2570,N_2644);
xor U2859 (N_2859,N_2687,N_2618);
nor U2860 (N_2860,N_2654,N_2686);
and U2861 (N_2861,N_2593,N_2708);
xnor U2862 (N_2862,N_2695,N_2647);
and U2863 (N_2863,N_2574,N_2696);
xor U2864 (N_2864,N_2644,N_2687);
or U2865 (N_2865,N_2633,N_2635);
xnor U2866 (N_2866,N_2622,N_2676);
xor U2867 (N_2867,N_2622,N_2609);
and U2868 (N_2868,N_2707,N_2579);
nand U2869 (N_2869,N_2689,N_2617);
nor U2870 (N_2870,N_2624,N_2618);
and U2871 (N_2871,N_2571,N_2598);
and U2872 (N_2872,N_2668,N_2592);
nand U2873 (N_2873,N_2625,N_2705);
xnor U2874 (N_2874,N_2689,N_2595);
or U2875 (N_2875,N_2653,N_2596);
nand U2876 (N_2876,N_2681,N_2656);
xnor U2877 (N_2877,N_2623,N_2682);
and U2878 (N_2878,N_2621,N_2667);
nor U2879 (N_2879,N_2677,N_2626);
xor U2880 (N_2880,N_2782,N_2844);
nand U2881 (N_2881,N_2738,N_2728);
nand U2882 (N_2882,N_2752,N_2839);
nand U2883 (N_2883,N_2760,N_2867);
or U2884 (N_2884,N_2737,N_2869);
nor U2885 (N_2885,N_2855,N_2789);
and U2886 (N_2886,N_2746,N_2857);
nor U2887 (N_2887,N_2836,N_2872);
xor U2888 (N_2888,N_2847,N_2819);
nand U2889 (N_2889,N_2798,N_2775);
or U2890 (N_2890,N_2854,N_2841);
or U2891 (N_2891,N_2758,N_2723);
nand U2892 (N_2892,N_2809,N_2829);
nor U2893 (N_2893,N_2779,N_2795);
and U2894 (N_2894,N_2826,N_2731);
nand U2895 (N_2895,N_2761,N_2832);
or U2896 (N_2896,N_2864,N_2755);
and U2897 (N_2897,N_2787,N_2858);
xor U2898 (N_2898,N_2743,N_2754);
nor U2899 (N_2899,N_2863,N_2773);
nand U2900 (N_2900,N_2767,N_2830);
and U2901 (N_2901,N_2786,N_2763);
nor U2902 (N_2902,N_2720,N_2772);
nand U2903 (N_2903,N_2784,N_2876);
or U2904 (N_2904,N_2785,N_2843);
and U2905 (N_2905,N_2825,N_2821);
xnor U2906 (N_2906,N_2769,N_2842);
and U2907 (N_2907,N_2848,N_2736);
nand U2908 (N_2908,N_2845,N_2726);
xor U2909 (N_2909,N_2794,N_2878);
or U2910 (N_2910,N_2788,N_2822);
and U2911 (N_2911,N_2730,N_2727);
nand U2912 (N_2912,N_2808,N_2824);
nand U2913 (N_2913,N_2729,N_2862);
nor U2914 (N_2914,N_2765,N_2770);
or U2915 (N_2915,N_2846,N_2879);
nand U2916 (N_2916,N_2766,N_2762);
xor U2917 (N_2917,N_2865,N_2817);
and U2918 (N_2918,N_2820,N_2732);
nand U2919 (N_2919,N_2800,N_2834);
nand U2920 (N_2920,N_2813,N_2733);
or U2921 (N_2921,N_2793,N_2870);
xor U2922 (N_2922,N_2757,N_2764);
nor U2923 (N_2923,N_2840,N_2810);
or U2924 (N_2924,N_2749,N_2837);
and U2925 (N_2925,N_2747,N_2814);
xnor U2926 (N_2926,N_2853,N_2861);
xnor U2927 (N_2927,N_2828,N_2807);
and U2928 (N_2928,N_2748,N_2792);
nor U2929 (N_2929,N_2734,N_2801);
or U2930 (N_2930,N_2774,N_2781);
xor U2931 (N_2931,N_2850,N_2722);
xnor U2932 (N_2932,N_2753,N_2735);
nand U2933 (N_2933,N_2750,N_2739);
and U2934 (N_2934,N_2740,N_2803);
or U2935 (N_2935,N_2721,N_2851);
nand U2936 (N_2936,N_2768,N_2790);
nor U2937 (N_2937,N_2776,N_2804);
xor U2938 (N_2938,N_2783,N_2812);
xor U2939 (N_2939,N_2744,N_2833);
nand U2940 (N_2940,N_2875,N_2823);
nor U2941 (N_2941,N_2802,N_2791);
and U2942 (N_2942,N_2741,N_2860);
nand U2943 (N_2943,N_2871,N_2759);
xor U2944 (N_2944,N_2745,N_2797);
and U2945 (N_2945,N_2796,N_2856);
nor U2946 (N_2946,N_2877,N_2806);
nor U2947 (N_2947,N_2778,N_2874);
xor U2948 (N_2948,N_2756,N_2835);
nor U2949 (N_2949,N_2777,N_2815);
and U2950 (N_2950,N_2742,N_2816);
xnor U2951 (N_2951,N_2780,N_2831);
or U2952 (N_2952,N_2811,N_2868);
xnor U2953 (N_2953,N_2838,N_2818);
or U2954 (N_2954,N_2852,N_2859);
or U2955 (N_2955,N_2751,N_2873);
xor U2956 (N_2956,N_2827,N_2799);
nor U2957 (N_2957,N_2771,N_2849);
nand U2958 (N_2958,N_2724,N_2725);
nand U2959 (N_2959,N_2805,N_2866);
nor U2960 (N_2960,N_2795,N_2735);
or U2961 (N_2961,N_2783,N_2837);
nor U2962 (N_2962,N_2813,N_2849);
or U2963 (N_2963,N_2814,N_2800);
nor U2964 (N_2964,N_2869,N_2850);
xor U2965 (N_2965,N_2822,N_2781);
xnor U2966 (N_2966,N_2771,N_2752);
or U2967 (N_2967,N_2871,N_2842);
and U2968 (N_2968,N_2877,N_2829);
nand U2969 (N_2969,N_2724,N_2752);
and U2970 (N_2970,N_2729,N_2741);
xnor U2971 (N_2971,N_2745,N_2856);
nor U2972 (N_2972,N_2850,N_2822);
xnor U2973 (N_2973,N_2801,N_2759);
or U2974 (N_2974,N_2724,N_2860);
nand U2975 (N_2975,N_2752,N_2783);
xnor U2976 (N_2976,N_2810,N_2782);
or U2977 (N_2977,N_2815,N_2825);
nor U2978 (N_2978,N_2844,N_2725);
or U2979 (N_2979,N_2736,N_2785);
or U2980 (N_2980,N_2779,N_2832);
nor U2981 (N_2981,N_2841,N_2745);
xnor U2982 (N_2982,N_2733,N_2794);
nand U2983 (N_2983,N_2788,N_2728);
nand U2984 (N_2984,N_2761,N_2848);
nor U2985 (N_2985,N_2859,N_2764);
nand U2986 (N_2986,N_2783,N_2797);
nor U2987 (N_2987,N_2723,N_2875);
nand U2988 (N_2988,N_2773,N_2741);
and U2989 (N_2989,N_2791,N_2770);
or U2990 (N_2990,N_2725,N_2803);
nor U2991 (N_2991,N_2743,N_2807);
nor U2992 (N_2992,N_2779,N_2787);
nor U2993 (N_2993,N_2770,N_2783);
nand U2994 (N_2994,N_2759,N_2857);
nor U2995 (N_2995,N_2734,N_2768);
nand U2996 (N_2996,N_2802,N_2850);
nand U2997 (N_2997,N_2813,N_2727);
nor U2998 (N_2998,N_2774,N_2828);
and U2999 (N_2999,N_2832,N_2855);
and U3000 (N_3000,N_2841,N_2869);
xor U3001 (N_3001,N_2736,N_2876);
nor U3002 (N_3002,N_2865,N_2868);
nor U3003 (N_3003,N_2746,N_2833);
or U3004 (N_3004,N_2831,N_2806);
nand U3005 (N_3005,N_2787,N_2781);
nand U3006 (N_3006,N_2832,N_2738);
nand U3007 (N_3007,N_2807,N_2774);
nand U3008 (N_3008,N_2822,N_2759);
xnor U3009 (N_3009,N_2799,N_2731);
or U3010 (N_3010,N_2754,N_2878);
nor U3011 (N_3011,N_2726,N_2741);
xor U3012 (N_3012,N_2815,N_2748);
and U3013 (N_3013,N_2755,N_2784);
nor U3014 (N_3014,N_2743,N_2767);
nor U3015 (N_3015,N_2819,N_2724);
nand U3016 (N_3016,N_2840,N_2867);
nor U3017 (N_3017,N_2837,N_2728);
nor U3018 (N_3018,N_2845,N_2830);
and U3019 (N_3019,N_2774,N_2870);
and U3020 (N_3020,N_2852,N_2725);
xnor U3021 (N_3021,N_2855,N_2733);
xor U3022 (N_3022,N_2746,N_2876);
and U3023 (N_3023,N_2809,N_2738);
xor U3024 (N_3024,N_2868,N_2801);
or U3025 (N_3025,N_2738,N_2769);
nor U3026 (N_3026,N_2832,N_2782);
nor U3027 (N_3027,N_2825,N_2856);
xnor U3028 (N_3028,N_2847,N_2828);
or U3029 (N_3029,N_2875,N_2788);
and U3030 (N_3030,N_2724,N_2849);
nand U3031 (N_3031,N_2874,N_2817);
or U3032 (N_3032,N_2845,N_2727);
or U3033 (N_3033,N_2832,N_2844);
nor U3034 (N_3034,N_2797,N_2860);
nand U3035 (N_3035,N_2753,N_2782);
xor U3036 (N_3036,N_2749,N_2787);
or U3037 (N_3037,N_2758,N_2872);
and U3038 (N_3038,N_2734,N_2859);
or U3039 (N_3039,N_2862,N_2818);
or U3040 (N_3040,N_2969,N_3002);
or U3041 (N_3041,N_3035,N_2923);
xnor U3042 (N_3042,N_3025,N_2973);
or U3043 (N_3043,N_3017,N_2920);
nor U3044 (N_3044,N_2949,N_2884);
nor U3045 (N_3045,N_2895,N_2885);
and U3046 (N_3046,N_2937,N_2948);
nand U3047 (N_3047,N_2927,N_2914);
nand U3048 (N_3048,N_3030,N_2989);
nor U3049 (N_3049,N_3027,N_2993);
xor U3050 (N_3050,N_2947,N_2894);
or U3051 (N_3051,N_3019,N_2881);
and U3052 (N_3052,N_2925,N_2886);
nand U3053 (N_3053,N_2913,N_2896);
xnor U3054 (N_3054,N_2965,N_2901);
xor U3055 (N_3055,N_3022,N_2990);
nand U3056 (N_3056,N_2982,N_2961);
nor U3057 (N_3057,N_2916,N_2955);
and U3058 (N_3058,N_2981,N_3010);
nand U3059 (N_3059,N_2977,N_2960);
and U3060 (N_3060,N_2984,N_2908);
nor U3061 (N_3061,N_2883,N_2942);
or U3062 (N_3062,N_2946,N_3023);
nand U3063 (N_3063,N_3012,N_2970);
or U3064 (N_3064,N_2903,N_3016);
or U3065 (N_3065,N_3028,N_2939);
nor U3066 (N_3066,N_2902,N_2924);
or U3067 (N_3067,N_3018,N_3033);
or U3068 (N_3068,N_2882,N_2880);
xor U3069 (N_3069,N_2985,N_3007);
or U3070 (N_3070,N_2935,N_2958);
xnor U3071 (N_3071,N_2918,N_2889);
nor U3072 (N_3072,N_2929,N_3034);
or U3073 (N_3073,N_2968,N_2988);
nor U3074 (N_3074,N_2967,N_2928);
or U3075 (N_3075,N_2892,N_2907);
nor U3076 (N_3076,N_2911,N_2997);
nand U3077 (N_3077,N_2963,N_2953);
or U3078 (N_3078,N_3005,N_2945);
xor U3079 (N_3079,N_3036,N_2943);
or U3080 (N_3080,N_3037,N_2976);
xnor U3081 (N_3081,N_2995,N_3026);
xnor U3082 (N_3082,N_2932,N_2952);
xor U3083 (N_3083,N_2917,N_2954);
nor U3084 (N_3084,N_3003,N_2986);
or U3085 (N_3085,N_2926,N_3006);
nor U3086 (N_3086,N_2922,N_3014);
and U3087 (N_3087,N_2890,N_2910);
or U3088 (N_3088,N_3004,N_2998);
or U3089 (N_3089,N_2944,N_2893);
nor U3090 (N_3090,N_2888,N_2950);
nor U3091 (N_3091,N_2938,N_2956);
or U3092 (N_3092,N_3013,N_2992);
or U3093 (N_3093,N_2900,N_2962);
and U3094 (N_3094,N_2983,N_2940);
nand U3095 (N_3095,N_2999,N_2897);
nor U3096 (N_3096,N_2975,N_3001);
nand U3097 (N_3097,N_3039,N_2957);
and U3098 (N_3098,N_3000,N_3024);
nor U3099 (N_3099,N_2933,N_2904);
nand U3100 (N_3100,N_3029,N_2915);
and U3101 (N_3101,N_2966,N_2971);
or U3102 (N_3102,N_2951,N_2898);
or U3103 (N_3103,N_3021,N_2887);
xnor U3104 (N_3104,N_2934,N_2978);
nor U3105 (N_3105,N_2994,N_2919);
nor U3106 (N_3106,N_2936,N_2987);
nor U3107 (N_3107,N_3008,N_2899);
xor U3108 (N_3108,N_2921,N_2972);
and U3109 (N_3109,N_2906,N_2905);
or U3110 (N_3110,N_2964,N_2979);
nand U3111 (N_3111,N_2980,N_3011);
and U3112 (N_3112,N_3015,N_2912);
or U3113 (N_3113,N_2891,N_3032);
nand U3114 (N_3114,N_2959,N_2974);
or U3115 (N_3115,N_3038,N_2930);
nor U3116 (N_3116,N_2996,N_3009);
nand U3117 (N_3117,N_2931,N_2909);
xor U3118 (N_3118,N_3031,N_2941);
or U3119 (N_3119,N_3020,N_2991);
and U3120 (N_3120,N_2880,N_2919);
nand U3121 (N_3121,N_2894,N_2935);
nor U3122 (N_3122,N_3035,N_2895);
nor U3123 (N_3123,N_3032,N_2881);
and U3124 (N_3124,N_2914,N_2967);
and U3125 (N_3125,N_2953,N_2946);
nor U3126 (N_3126,N_2948,N_2992);
nor U3127 (N_3127,N_3014,N_2976);
nor U3128 (N_3128,N_2995,N_2982);
nor U3129 (N_3129,N_3030,N_2956);
xor U3130 (N_3130,N_2976,N_2932);
and U3131 (N_3131,N_2881,N_3015);
nand U3132 (N_3132,N_3030,N_3000);
or U3133 (N_3133,N_2920,N_2999);
nand U3134 (N_3134,N_3011,N_3038);
nand U3135 (N_3135,N_3038,N_3017);
nor U3136 (N_3136,N_2973,N_2958);
or U3137 (N_3137,N_3019,N_2936);
xnor U3138 (N_3138,N_2946,N_2881);
or U3139 (N_3139,N_2952,N_2968);
nor U3140 (N_3140,N_2897,N_2942);
and U3141 (N_3141,N_2949,N_3038);
xnor U3142 (N_3142,N_2889,N_2969);
and U3143 (N_3143,N_2887,N_2988);
xor U3144 (N_3144,N_2889,N_2921);
nor U3145 (N_3145,N_2887,N_2972);
nand U3146 (N_3146,N_3028,N_2891);
nand U3147 (N_3147,N_2885,N_2897);
and U3148 (N_3148,N_2939,N_2987);
xnor U3149 (N_3149,N_2937,N_3018);
and U3150 (N_3150,N_3038,N_3014);
nor U3151 (N_3151,N_2955,N_2940);
nor U3152 (N_3152,N_3014,N_2918);
and U3153 (N_3153,N_2968,N_2886);
nor U3154 (N_3154,N_3001,N_2942);
or U3155 (N_3155,N_2881,N_3008);
or U3156 (N_3156,N_2930,N_2962);
and U3157 (N_3157,N_2997,N_2976);
nand U3158 (N_3158,N_2958,N_3008);
nor U3159 (N_3159,N_2957,N_2961);
nand U3160 (N_3160,N_3011,N_2948);
nor U3161 (N_3161,N_2981,N_2921);
nor U3162 (N_3162,N_2918,N_3022);
nand U3163 (N_3163,N_2897,N_2970);
and U3164 (N_3164,N_2933,N_3032);
nand U3165 (N_3165,N_2913,N_2914);
xor U3166 (N_3166,N_2960,N_2962);
nand U3167 (N_3167,N_2882,N_2906);
nor U3168 (N_3168,N_2941,N_3018);
or U3169 (N_3169,N_2976,N_2894);
or U3170 (N_3170,N_2981,N_2996);
or U3171 (N_3171,N_2991,N_2948);
nor U3172 (N_3172,N_2947,N_2963);
nand U3173 (N_3173,N_2912,N_2967);
or U3174 (N_3174,N_2985,N_2897);
xnor U3175 (N_3175,N_2966,N_3004);
xor U3176 (N_3176,N_2956,N_2880);
nand U3177 (N_3177,N_2969,N_2940);
or U3178 (N_3178,N_2939,N_3014);
and U3179 (N_3179,N_2983,N_2956);
and U3180 (N_3180,N_2894,N_2980);
xnor U3181 (N_3181,N_2953,N_3028);
nand U3182 (N_3182,N_2969,N_2891);
xnor U3183 (N_3183,N_3037,N_2993);
nand U3184 (N_3184,N_3018,N_2901);
or U3185 (N_3185,N_3033,N_2954);
nand U3186 (N_3186,N_2948,N_2975);
nor U3187 (N_3187,N_2898,N_3026);
or U3188 (N_3188,N_2984,N_2930);
or U3189 (N_3189,N_2897,N_3032);
xnor U3190 (N_3190,N_3027,N_3022);
and U3191 (N_3191,N_2974,N_2969);
and U3192 (N_3192,N_2894,N_2997);
xnor U3193 (N_3193,N_2996,N_2916);
nor U3194 (N_3194,N_3031,N_2943);
nor U3195 (N_3195,N_2985,N_2969);
and U3196 (N_3196,N_3014,N_3031);
nand U3197 (N_3197,N_2938,N_3007);
or U3198 (N_3198,N_2906,N_2966);
nand U3199 (N_3199,N_3000,N_2939);
or U3200 (N_3200,N_3081,N_3063);
or U3201 (N_3201,N_3187,N_3055);
nand U3202 (N_3202,N_3110,N_3159);
nand U3203 (N_3203,N_3146,N_3067);
nor U3204 (N_3204,N_3073,N_3065);
and U3205 (N_3205,N_3164,N_3145);
xnor U3206 (N_3206,N_3050,N_3053);
nor U3207 (N_3207,N_3101,N_3113);
or U3208 (N_3208,N_3041,N_3044);
or U3209 (N_3209,N_3096,N_3132);
nand U3210 (N_3210,N_3177,N_3047);
xnor U3211 (N_3211,N_3066,N_3048);
or U3212 (N_3212,N_3056,N_3153);
nor U3213 (N_3213,N_3119,N_3160);
or U3214 (N_3214,N_3173,N_3071);
and U3215 (N_3215,N_3049,N_3078);
xnor U3216 (N_3216,N_3165,N_3123);
nand U3217 (N_3217,N_3114,N_3057);
nand U3218 (N_3218,N_3128,N_3196);
xnor U3219 (N_3219,N_3106,N_3095);
or U3220 (N_3220,N_3180,N_3094);
and U3221 (N_3221,N_3140,N_3188);
or U3222 (N_3222,N_3148,N_3116);
nand U3223 (N_3223,N_3150,N_3062);
nand U3224 (N_3224,N_3195,N_3058);
nor U3225 (N_3225,N_3069,N_3137);
or U3226 (N_3226,N_3126,N_3133);
and U3227 (N_3227,N_3109,N_3163);
and U3228 (N_3228,N_3117,N_3098);
or U3229 (N_3229,N_3134,N_3147);
xnor U3230 (N_3230,N_3197,N_3168);
nand U3231 (N_3231,N_3099,N_3089);
nand U3232 (N_3232,N_3182,N_3157);
and U3233 (N_3233,N_3179,N_3108);
and U3234 (N_3234,N_3152,N_3174);
nand U3235 (N_3235,N_3190,N_3072);
xnor U3236 (N_3236,N_3161,N_3143);
xnor U3237 (N_3237,N_3064,N_3111);
nor U3238 (N_3238,N_3046,N_3189);
and U3239 (N_3239,N_3130,N_3199);
nand U3240 (N_3240,N_3070,N_3198);
and U3241 (N_3241,N_3043,N_3155);
nor U3242 (N_3242,N_3084,N_3135);
nand U3243 (N_3243,N_3091,N_3139);
and U3244 (N_3244,N_3131,N_3076);
or U3245 (N_3245,N_3127,N_3104);
nand U3246 (N_3246,N_3086,N_3136);
or U3247 (N_3247,N_3051,N_3083);
or U3248 (N_3248,N_3054,N_3112);
xor U3249 (N_3249,N_3079,N_3176);
or U3250 (N_3250,N_3080,N_3171);
nor U3251 (N_3251,N_3097,N_3118);
and U3252 (N_3252,N_3040,N_3120);
or U3253 (N_3253,N_3059,N_3138);
xnor U3254 (N_3254,N_3186,N_3162);
nor U3255 (N_3255,N_3122,N_3103);
and U3256 (N_3256,N_3100,N_3181);
and U3257 (N_3257,N_3105,N_3107);
nand U3258 (N_3258,N_3169,N_3102);
or U3259 (N_3259,N_3172,N_3074);
nand U3260 (N_3260,N_3125,N_3121);
nand U3261 (N_3261,N_3052,N_3194);
and U3262 (N_3262,N_3124,N_3061);
and U3263 (N_3263,N_3185,N_3085);
or U3264 (N_3264,N_3142,N_3144);
nand U3265 (N_3265,N_3166,N_3088);
nand U3266 (N_3266,N_3156,N_3082);
and U3267 (N_3267,N_3167,N_3193);
nand U3268 (N_3268,N_3154,N_3060);
nor U3269 (N_3269,N_3191,N_3075);
and U3270 (N_3270,N_3129,N_3045);
nand U3271 (N_3271,N_3093,N_3141);
nand U3272 (N_3272,N_3170,N_3184);
nor U3273 (N_3273,N_3183,N_3158);
nand U3274 (N_3274,N_3178,N_3192);
nand U3275 (N_3275,N_3087,N_3149);
and U3276 (N_3276,N_3068,N_3090);
nand U3277 (N_3277,N_3092,N_3175);
or U3278 (N_3278,N_3151,N_3077);
nand U3279 (N_3279,N_3115,N_3042);
nor U3280 (N_3280,N_3099,N_3127);
nor U3281 (N_3281,N_3157,N_3065);
nor U3282 (N_3282,N_3195,N_3199);
xnor U3283 (N_3283,N_3116,N_3181);
nor U3284 (N_3284,N_3048,N_3082);
nand U3285 (N_3285,N_3173,N_3088);
and U3286 (N_3286,N_3041,N_3070);
nand U3287 (N_3287,N_3132,N_3194);
xnor U3288 (N_3288,N_3139,N_3056);
nand U3289 (N_3289,N_3180,N_3159);
xor U3290 (N_3290,N_3144,N_3150);
or U3291 (N_3291,N_3073,N_3137);
nor U3292 (N_3292,N_3165,N_3156);
nor U3293 (N_3293,N_3124,N_3052);
nand U3294 (N_3294,N_3087,N_3080);
xnor U3295 (N_3295,N_3045,N_3169);
or U3296 (N_3296,N_3170,N_3089);
nand U3297 (N_3297,N_3061,N_3105);
and U3298 (N_3298,N_3163,N_3179);
and U3299 (N_3299,N_3178,N_3184);
or U3300 (N_3300,N_3047,N_3082);
xor U3301 (N_3301,N_3076,N_3062);
nor U3302 (N_3302,N_3142,N_3099);
and U3303 (N_3303,N_3173,N_3171);
xor U3304 (N_3304,N_3123,N_3180);
and U3305 (N_3305,N_3180,N_3040);
nand U3306 (N_3306,N_3198,N_3179);
or U3307 (N_3307,N_3074,N_3044);
or U3308 (N_3308,N_3059,N_3168);
nand U3309 (N_3309,N_3124,N_3060);
xnor U3310 (N_3310,N_3128,N_3050);
xnor U3311 (N_3311,N_3145,N_3193);
nor U3312 (N_3312,N_3071,N_3171);
nand U3313 (N_3313,N_3130,N_3044);
xor U3314 (N_3314,N_3184,N_3120);
nand U3315 (N_3315,N_3072,N_3070);
nand U3316 (N_3316,N_3171,N_3166);
nor U3317 (N_3317,N_3059,N_3114);
or U3318 (N_3318,N_3080,N_3151);
nand U3319 (N_3319,N_3128,N_3146);
xnor U3320 (N_3320,N_3113,N_3091);
nand U3321 (N_3321,N_3053,N_3079);
or U3322 (N_3322,N_3148,N_3086);
xnor U3323 (N_3323,N_3084,N_3044);
and U3324 (N_3324,N_3149,N_3133);
nand U3325 (N_3325,N_3080,N_3195);
nand U3326 (N_3326,N_3090,N_3046);
nand U3327 (N_3327,N_3111,N_3114);
or U3328 (N_3328,N_3191,N_3082);
or U3329 (N_3329,N_3198,N_3048);
or U3330 (N_3330,N_3172,N_3176);
nand U3331 (N_3331,N_3177,N_3168);
xor U3332 (N_3332,N_3100,N_3180);
nor U3333 (N_3333,N_3103,N_3092);
nand U3334 (N_3334,N_3178,N_3152);
xnor U3335 (N_3335,N_3126,N_3152);
nand U3336 (N_3336,N_3191,N_3185);
nand U3337 (N_3337,N_3101,N_3120);
and U3338 (N_3338,N_3165,N_3076);
xnor U3339 (N_3339,N_3073,N_3119);
xor U3340 (N_3340,N_3052,N_3184);
and U3341 (N_3341,N_3162,N_3173);
nand U3342 (N_3342,N_3177,N_3053);
or U3343 (N_3343,N_3064,N_3107);
or U3344 (N_3344,N_3102,N_3135);
or U3345 (N_3345,N_3063,N_3097);
nor U3346 (N_3346,N_3089,N_3058);
xnor U3347 (N_3347,N_3096,N_3122);
nand U3348 (N_3348,N_3186,N_3170);
nor U3349 (N_3349,N_3153,N_3101);
nor U3350 (N_3350,N_3052,N_3130);
or U3351 (N_3351,N_3091,N_3120);
nor U3352 (N_3352,N_3195,N_3057);
nand U3353 (N_3353,N_3114,N_3116);
xor U3354 (N_3354,N_3054,N_3168);
or U3355 (N_3355,N_3060,N_3164);
and U3356 (N_3356,N_3084,N_3181);
nor U3357 (N_3357,N_3170,N_3046);
nor U3358 (N_3358,N_3165,N_3174);
xor U3359 (N_3359,N_3177,N_3130);
or U3360 (N_3360,N_3245,N_3257);
nand U3361 (N_3361,N_3327,N_3213);
xor U3362 (N_3362,N_3214,N_3232);
nand U3363 (N_3363,N_3247,N_3292);
nor U3364 (N_3364,N_3201,N_3342);
or U3365 (N_3365,N_3304,N_3288);
xnor U3366 (N_3366,N_3268,N_3223);
nor U3367 (N_3367,N_3348,N_3266);
or U3368 (N_3368,N_3273,N_3321);
nor U3369 (N_3369,N_3295,N_3280);
nor U3370 (N_3370,N_3258,N_3317);
nand U3371 (N_3371,N_3315,N_3303);
xnor U3372 (N_3372,N_3281,N_3320);
nand U3373 (N_3373,N_3328,N_3322);
and U3374 (N_3374,N_3284,N_3262);
and U3375 (N_3375,N_3345,N_3259);
nor U3376 (N_3376,N_3243,N_3310);
nand U3377 (N_3377,N_3233,N_3236);
or U3378 (N_3378,N_3336,N_3324);
and U3379 (N_3379,N_3301,N_3294);
nor U3380 (N_3380,N_3282,N_3216);
nor U3381 (N_3381,N_3253,N_3238);
xor U3382 (N_3382,N_3334,N_3285);
xnor U3383 (N_3383,N_3225,N_3209);
nand U3384 (N_3384,N_3237,N_3202);
nor U3385 (N_3385,N_3274,N_3332);
or U3386 (N_3386,N_3219,N_3260);
xnor U3387 (N_3387,N_3265,N_3251);
xor U3388 (N_3388,N_3299,N_3316);
and U3389 (N_3389,N_3211,N_3312);
or U3390 (N_3390,N_3212,N_3226);
nor U3391 (N_3391,N_3318,N_3341);
nand U3392 (N_3392,N_3290,N_3256);
and U3393 (N_3393,N_3337,N_3331);
nand U3394 (N_3394,N_3264,N_3261);
xor U3395 (N_3395,N_3286,N_3297);
or U3396 (N_3396,N_3291,N_3335);
nor U3397 (N_3397,N_3340,N_3267);
nor U3398 (N_3398,N_3287,N_3306);
nand U3399 (N_3399,N_3222,N_3203);
or U3400 (N_3400,N_3204,N_3235);
and U3401 (N_3401,N_3206,N_3283);
xor U3402 (N_3402,N_3263,N_3242);
or U3403 (N_3403,N_3240,N_3200);
and U3404 (N_3404,N_3329,N_3246);
nand U3405 (N_3405,N_3230,N_3305);
and U3406 (N_3406,N_3356,N_3215);
xor U3407 (N_3407,N_3248,N_3349);
xnor U3408 (N_3408,N_3325,N_3227);
nand U3409 (N_3409,N_3269,N_3293);
or U3410 (N_3410,N_3277,N_3224);
nor U3411 (N_3411,N_3307,N_3338);
or U3412 (N_3412,N_3358,N_3276);
xnor U3413 (N_3413,N_3359,N_3229);
nand U3414 (N_3414,N_3221,N_3234);
or U3415 (N_3415,N_3309,N_3355);
and U3416 (N_3416,N_3323,N_3339);
and U3417 (N_3417,N_3250,N_3220);
and U3418 (N_3418,N_3352,N_3344);
and U3419 (N_3419,N_3228,N_3354);
xnor U3420 (N_3420,N_3353,N_3231);
xor U3421 (N_3421,N_3289,N_3208);
nand U3422 (N_3422,N_3296,N_3271);
or U3423 (N_3423,N_3218,N_3350);
xnor U3424 (N_3424,N_3272,N_3249);
xnor U3425 (N_3425,N_3330,N_3351);
and U3426 (N_3426,N_3314,N_3205);
nor U3427 (N_3427,N_3298,N_3279);
nand U3428 (N_3428,N_3239,N_3254);
nand U3429 (N_3429,N_3270,N_3313);
xnor U3430 (N_3430,N_3207,N_3346);
xor U3431 (N_3431,N_3210,N_3311);
or U3432 (N_3432,N_3326,N_3255);
xnor U3433 (N_3433,N_3347,N_3300);
xnor U3434 (N_3434,N_3217,N_3252);
or U3435 (N_3435,N_3302,N_3319);
or U3436 (N_3436,N_3357,N_3343);
or U3437 (N_3437,N_3241,N_3308);
or U3438 (N_3438,N_3244,N_3278);
nor U3439 (N_3439,N_3275,N_3333);
xnor U3440 (N_3440,N_3211,N_3313);
xnor U3441 (N_3441,N_3347,N_3330);
xnor U3442 (N_3442,N_3301,N_3310);
and U3443 (N_3443,N_3325,N_3296);
and U3444 (N_3444,N_3278,N_3314);
xnor U3445 (N_3445,N_3334,N_3341);
nand U3446 (N_3446,N_3258,N_3293);
or U3447 (N_3447,N_3325,N_3306);
nor U3448 (N_3448,N_3303,N_3222);
nor U3449 (N_3449,N_3253,N_3250);
nand U3450 (N_3450,N_3329,N_3233);
nor U3451 (N_3451,N_3263,N_3326);
and U3452 (N_3452,N_3213,N_3230);
and U3453 (N_3453,N_3211,N_3297);
nand U3454 (N_3454,N_3250,N_3216);
nor U3455 (N_3455,N_3323,N_3206);
xnor U3456 (N_3456,N_3293,N_3235);
or U3457 (N_3457,N_3314,N_3257);
or U3458 (N_3458,N_3313,N_3323);
xor U3459 (N_3459,N_3311,N_3355);
and U3460 (N_3460,N_3267,N_3304);
and U3461 (N_3461,N_3258,N_3328);
nor U3462 (N_3462,N_3333,N_3256);
xnor U3463 (N_3463,N_3202,N_3288);
nor U3464 (N_3464,N_3262,N_3293);
or U3465 (N_3465,N_3358,N_3210);
nand U3466 (N_3466,N_3213,N_3305);
or U3467 (N_3467,N_3281,N_3277);
nor U3468 (N_3468,N_3208,N_3272);
xor U3469 (N_3469,N_3223,N_3272);
nor U3470 (N_3470,N_3223,N_3274);
nand U3471 (N_3471,N_3217,N_3210);
or U3472 (N_3472,N_3235,N_3280);
and U3473 (N_3473,N_3284,N_3345);
and U3474 (N_3474,N_3315,N_3301);
nor U3475 (N_3475,N_3286,N_3322);
xor U3476 (N_3476,N_3233,N_3311);
or U3477 (N_3477,N_3349,N_3325);
xnor U3478 (N_3478,N_3206,N_3277);
nand U3479 (N_3479,N_3258,N_3311);
nand U3480 (N_3480,N_3314,N_3358);
xnor U3481 (N_3481,N_3255,N_3202);
or U3482 (N_3482,N_3356,N_3206);
nor U3483 (N_3483,N_3309,N_3352);
xor U3484 (N_3484,N_3358,N_3232);
xor U3485 (N_3485,N_3347,N_3325);
xor U3486 (N_3486,N_3237,N_3236);
xor U3487 (N_3487,N_3240,N_3324);
or U3488 (N_3488,N_3326,N_3315);
and U3489 (N_3489,N_3267,N_3291);
nand U3490 (N_3490,N_3228,N_3322);
and U3491 (N_3491,N_3285,N_3291);
or U3492 (N_3492,N_3304,N_3309);
or U3493 (N_3493,N_3234,N_3257);
xor U3494 (N_3494,N_3228,N_3221);
and U3495 (N_3495,N_3348,N_3216);
nand U3496 (N_3496,N_3214,N_3262);
nor U3497 (N_3497,N_3250,N_3255);
and U3498 (N_3498,N_3261,N_3269);
nor U3499 (N_3499,N_3240,N_3234);
xor U3500 (N_3500,N_3296,N_3254);
xnor U3501 (N_3501,N_3355,N_3274);
nor U3502 (N_3502,N_3329,N_3212);
and U3503 (N_3503,N_3215,N_3232);
nand U3504 (N_3504,N_3314,N_3268);
or U3505 (N_3505,N_3278,N_3335);
nand U3506 (N_3506,N_3327,N_3287);
nand U3507 (N_3507,N_3213,N_3290);
xnor U3508 (N_3508,N_3273,N_3303);
nand U3509 (N_3509,N_3298,N_3226);
or U3510 (N_3510,N_3280,N_3344);
nand U3511 (N_3511,N_3317,N_3346);
and U3512 (N_3512,N_3286,N_3216);
nand U3513 (N_3513,N_3281,N_3279);
and U3514 (N_3514,N_3320,N_3279);
or U3515 (N_3515,N_3354,N_3280);
nor U3516 (N_3516,N_3356,N_3247);
nand U3517 (N_3517,N_3307,N_3333);
xnor U3518 (N_3518,N_3282,N_3296);
or U3519 (N_3519,N_3203,N_3224);
and U3520 (N_3520,N_3502,N_3463);
nand U3521 (N_3521,N_3441,N_3489);
or U3522 (N_3522,N_3454,N_3388);
or U3523 (N_3523,N_3488,N_3370);
xor U3524 (N_3524,N_3421,N_3496);
nand U3525 (N_3525,N_3472,N_3400);
xnor U3526 (N_3526,N_3425,N_3360);
nor U3527 (N_3527,N_3437,N_3452);
or U3528 (N_3528,N_3442,N_3427);
nand U3529 (N_3529,N_3398,N_3467);
xor U3530 (N_3530,N_3436,N_3375);
nand U3531 (N_3531,N_3422,N_3376);
nand U3532 (N_3532,N_3405,N_3382);
and U3533 (N_3533,N_3414,N_3482);
or U3534 (N_3534,N_3429,N_3368);
or U3535 (N_3535,N_3387,N_3444);
nor U3536 (N_3536,N_3448,N_3395);
or U3537 (N_3537,N_3457,N_3426);
and U3538 (N_3538,N_3424,N_3413);
and U3539 (N_3539,N_3419,N_3417);
and U3540 (N_3540,N_3471,N_3487);
and U3541 (N_3541,N_3476,N_3386);
and U3542 (N_3542,N_3495,N_3434);
and U3543 (N_3543,N_3506,N_3420);
or U3544 (N_3544,N_3513,N_3407);
nand U3545 (N_3545,N_3456,N_3464);
or U3546 (N_3546,N_3381,N_3443);
nand U3547 (N_3547,N_3483,N_3469);
nor U3548 (N_3548,N_3449,N_3401);
nor U3549 (N_3549,N_3412,N_3518);
nor U3550 (N_3550,N_3432,N_3475);
nor U3551 (N_3551,N_3460,N_3404);
xnor U3552 (N_3552,N_3519,N_3508);
and U3553 (N_3553,N_3498,N_3435);
nor U3554 (N_3554,N_3372,N_3497);
nand U3555 (N_3555,N_3415,N_3416);
nor U3556 (N_3556,N_3408,N_3394);
or U3557 (N_3557,N_3481,N_3411);
nor U3558 (N_3558,N_3410,N_3465);
xor U3559 (N_3559,N_3371,N_3430);
nor U3560 (N_3560,N_3440,N_3458);
nor U3561 (N_3561,N_3491,N_3493);
xnor U3562 (N_3562,N_3505,N_3445);
xnor U3563 (N_3563,N_3369,N_3361);
xor U3564 (N_3564,N_3365,N_3478);
nor U3565 (N_3565,N_3367,N_3499);
nand U3566 (N_3566,N_3378,N_3377);
nor U3567 (N_3567,N_3516,N_3366);
nor U3568 (N_3568,N_3439,N_3406);
xnor U3569 (N_3569,N_3392,N_3517);
xnor U3570 (N_3570,N_3501,N_3450);
nor U3571 (N_3571,N_3477,N_3461);
xor U3572 (N_3572,N_3409,N_3390);
and U3573 (N_3573,N_3403,N_3374);
nand U3574 (N_3574,N_3399,N_3385);
and U3575 (N_3575,N_3364,N_3391);
nor U3576 (N_3576,N_3468,N_3466);
nand U3577 (N_3577,N_3509,N_3511);
nor U3578 (N_3578,N_3363,N_3433);
or U3579 (N_3579,N_3447,N_3494);
and U3580 (N_3580,N_3384,N_3453);
nor U3581 (N_3581,N_3362,N_3393);
xor U3582 (N_3582,N_3484,N_3490);
nand U3583 (N_3583,N_3512,N_3383);
nor U3584 (N_3584,N_3451,N_3510);
and U3585 (N_3585,N_3380,N_3485);
xnor U3586 (N_3586,N_3402,N_3470);
nor U3587 (N_3587,N_3423,N_3507);
xnor U3588 (N_3588,N_3504,N_3438);
xor U3589 (N_3589,N_3462,N_3389);
xnor U3590 (N_3590,N_3397,N_3480);
and U3591 (N_3591,N_3503,N_3492);
or U3592 (N_3592,N_3486,N_3418);
or U3593 (N_3593,N_3515,N_3514);
xnor U3594 (N_3594,N_3474,N_3473);
nand U3595 (N_3595,N_3428,N_3459);
or U3596 (N_3596,N_3431,N_3479);
nand U3597 (N_3597,N_3373,N_3396);
xor U3598 (N_3598,N_3446,N_3379);
nor U3599 (N_3599,N_3500,N_3455);
nand U3600 (N_3600,N_3362,N_3446);
nor U3601 (N_3601,N_3415,N_3519);
and U3602 (N_3602,N_3365,N_3387);
nor U3603 (N_3603,N_3498,N_3464);
or U3604 (N_3604,N_3489,N_3399);
or U3605 (N_3605,N_3426,N_3423);
xor U3606 (N_3606,N_3490,N_3499);
nand U3607 (N_3607,N_3417,N_3460);
and U3608 (N_3608,N_3395,N_3405);
nand U3609 (N_3609,N_3493,N_3463);
and U3610 (N_3610,N_3462,N_3436);
xnor U3611 (N_3611,N_3478,N_3489);
and U3612 (N_3612,N_3417,N_3372);
xor U3613 (N_3613,N_3419,N_3431);
xor U3614 (N_3614,N_3379,N_3494);
nor U3615 (N_3615,N_3362,N_3361);
nand U3616 (N_3616,N_3464,N_3516);
nor U3617 (N_3617,N_3444,N_3371);
or U3618 (N_3618,N_3380,N_3396);
nor U3619 (N_3619,N_3469,N_3363);
xor U3620 (N_3620,N_3457,N_3389);
nand U3621 (N_3621,N_3392,N_3486);
nand U3622 (N_3622,N_3466,N_3422);
xnor U3623 (N_3623,N_3471,N_3401);
nor U3624 (N_3624,N_3377,N_3463);
xnor U3625 (N_3625,N_3452,N_3376);
or U3626 (N_3626,N_3456,N_3430);
nand U3627 (N_3627,N_3456,N_3424);
nor U3628 (N_3628,N_3360,N_3473);
nand U3629 (N_3629,N_3460,N_3416);
and U3630 (N_3630,N_3380,N_3459);
xor U3631 (N_3631,N_3499,N_3493);
or U3632 (N_3632,N_3427,N_3517);
nand U3633 (N_3633,N_3508,N_3377);
or U3634 (N_3634,N_3505,N_3454);
xnor U3635 (N_3635,N_3414,N_3441);
nor U3636 (N_3636,N_3434,N_3411);
xnor U3637 (N_3637,N_3487,N_3504);
and U3638 (N_3638,N_3491,N_3450);
xnor U3639 (N_3639,N_3368,N_3391);
and U3640 (N_3640,N_3385,N_3433);
nand U3641 (N_3641,N_3490,N_3380);
and U3642 (N_3642,N_3491,N_3419);
nor U3643 (N_3643,N_3395,N_3420);
nor U3644 (N_3644,N_3469,N_3410);
nand U3645 (N_3645,N_3492,N_3413);
and U3646 (N_3646,N_3373,N_3452);
nand U3647 (N_3647,N_3434,N_3413);
and U3648 (N_3648,N_3364,N_3481);
and U3649 (N_3649,N_3430,N_3490);
or U3650 (N_3650,N_3463,N_3422);
or U3651 (N_3651,N_3437,N_3389);
xor U3652 (N_3652,N_3451,N_3511);
nor U3653 (N_3653,N_3418,N_3434);
and U3654 (N_3654,N_3513,N_3451);
and U3655 (N_3655,N_3492,N_3474);
nand U3656 (N_3656,N_3504,N_3453);
or U3657 (N_3657,N_3381,N_3498);
xnor U3658 (N_3658,N_3462,N_3480);
and U3659 (N_3659,N_3453,N_3459);
nand U3660 (N_3660,N_3374,N_3409);
nor U3661 (N_3661,N_3491,N_3425);
nand U3662 (N_3662,N_3494,N_3404);
or U3663 (N_3663,N_3403,N_3463);
xor U3664 (N_3664,N_3441,N_3514);
or U3665 (N_3665,N_3381,N_3482);
nand U3666 (N_3666,N_3470,N_3377);
nor U3667 (N_3667,N_3444,N_3436);
nor U3668 (N_3668,N_3510,N_3363);
or U3669 (N_3669,N_3490,N_3437);
or U3670 (N_3670,N_3497,N_3473);
and U3671 (N_3671,N_3417,N_3462);
or U3672 (N_3672,N_3372,N_3489);
nor U3673 (N_3673,N_3403,N_3506);
and U3674 (N_3674,N_3514,N_3453);
and U3675 (N_3675,N_3519,N_3484);
xnor U3676 (N_3676,N_3420,N_3419);
or U3677 (N_3677,N_3476,N_3460);
xnor U3678 (N_3678,N_3387,N_3482);
nand U3679 (N_3679,N_3382,N_3371);
and U3680 (N_3680,N_3542,N_3650);
or U3681 (N_3681,N_3548,N_3579);
and U3682 (N_3682,N_3522,N_3604);
and U3683 (N_3683,N_3552,N_3611);
and U3684 (N_3684,N_3607,N_3633);
nor U3685 (N_3685,N_3667,N_3544);
or U3686 (N_3686,N_3655,N_3556);
and U3687 (N_3687,N_3644,N_3618);
nand U3688 (N_3688,N_3576,N_3614);
nor U3689 (N_3689,N_3674,N_3539);
nor U3690 (N_3690,N_3570,N_3608);
or U3691 (N_3691,N_3567,N_3565);
nor U3692 (N_3692,N_3589,N_3596);
or U3693 (N_3693,N_3609,N_3669);
nand U3694 (N_3694,N_3605,N_3640);
and U3695 (N_3695,N_3617,N_3591);
or U3696 (N_3696,N_3584,N_3677);
xnor U3697 (N_3697,N_3534,N_3612);
or U3698 (N_3698,N_3602,N_3530);
nand U3699 (N_3699,N_3631,N_3659);
and U3700 (N_3700,N_3594,N_3625);
xnor U3701 (N_3701,N_3676,N_3597);
or U3702 (N_3702,N_3661,N_3581);
xor U3703 (N_3703,N_3603,N_3638);
nand U3704 (N_3704,N_3538,N_3559);
or U3705 (N_3705,N_3563,N_3657);
xor U3706 (N_3706,N_3598,N_3653);
nand U3707 (N_3707,N_3529,N_3645);
and U3708 (N_3708,N_3652,N_3547);
or U3709 (N_3709,N_3610,N_3558);
nand U3710 (N_3710,N_3524,N_3540);
xnor U3711 (N_3711,N_3639,N_3564);
and U3712 (N_3712,N_3566,N_3553);
nand U3713 (N_3713,N_3649,N_3623);
nor U3714 (N_3714,N_3543,N_3660);
nand U3715 (N_3715,N_3600,N_3629);
xor U3716 (N_3716,N_3574,N_3537);
nor U3717 (N_3717,N_3678,N_3672);
nor U3718 (N_3718,N_3626,N_3580);
and U3719 (N_3719,N_3533,N_3572);
nand U3720 (N_3720,N_3521,N_3654);
and U3721 (N_3721,N_3630,N_3583);
nor U3722 (N_3722,N_3624,N_3599);
nand U3723 (N_3723,N_3595,N_3627);
nand U3724 (N_3724,N_3545,N_3535);
or U3725 (N_3725,N_3635,N_3658);
nand U3726 (N_3726,N_3585,N_3647);
xnor U3727 (N_3727,N_3641,N_3541);
or U3728 (N_3728,N_3670,N_3648);
nor U3729 (N_3729,N_3621,N_3668);
and U3730 (N_3730,N_3527,N_3665);
nor U3731 (N_3731,N_3646,N_3628);
and U3732 (N_3732,N_3622,N_3666);
xnor U3733 (N_3733,N_3577,N_3588);
nor U3734 (N_3734,N_3528,N_3642);
and U3735 (N_3735,N_3673,N_3531);
or U3736 (N_3736,N_3571,N_3663);
and U3737 (N_3737,N_3651,N_3606);
nor U3738 (N_3738,N_3590,N_3554);
nor U3739 (N_3739,N_3560,N_3578);
and U3740 (N_3740,N_3526,N_3619);
and U3741 (N_3741,N_3557,N_3549);
or U3742 (N_3742,N_3634,N_3555);
or U3743 (N_3743,N_3636,N_3620);
xor U3744 (N_3744,N_3601,N_3546);
or U3745 (N_3745,N_3675,N_3593);
and U3746 (N_3746,N_3550,N_3587);
nand U3747 (N_3747,N_3569,N_3568);
or U3748 (N_3748,N_3586,N_3532);
nand U3749 (N_3749,N_3523,N_3615);
or U3750 (N_3750,N_3613,N_3671);
nor U3751 (N_3751,N_3536,N_3520);
xor U3752 (N_3752,N_3575,N_3562);
nand U3753 (N_3753,N_3632,N_3643);
nor U3754 (N_3754,N_3679,N_3561);
or U3755 (N_3755,N_3664,N_3592);
nor U3756 (N_3756,N_3637,N_3582);
xor U3757 (N_3757,N_3551,N_3573);
or U3758 (N_3758,N_3616,N_3656);
and U3759 (N_3759,N_3662,N_3525);
nand U3760 (N_3760,N_3578,N_3582);
and U3761 (N_3761,N_3563,N_3585);
nor U3762 (N_3762,N_3640,N_3576);
xnor U3763 (N_3763,N_3653,N_3664);
and U3764 (N_3764,N_3679,N_3594);
nor U3765 (N_3765,N_3643,N_3591);
xnor U3766 (N_3766,N_3566,N_3576);
and U3767 (N_3767,N_3627,N_3620);
xnor U3768 (N_3768,N_3576,N_3554);
and U3769 (N_3769,N_3541,N_3562);
and U3770 (N_3770,N_3602,N_3525);
nor U3771 (N_3771,N_3620,N_3584);
xnor U3772 (N_3772,N_3618,N_3541);
nand U3773 (N_3773,N_3651,N_3603);
and U3774 (N_3774,N_3657,N_3678);
nor U3775 (N_3775,N_3655,N_3646);
and U3776 (N_3776,N_3567,N_3595);
nand U3777 (N_3777,N_3662,N_3635);
and U3778 (N_3778,N_3615,N_3600);
xor U3779 (N_3779,N_3520,N_3610);
xor U3780 (N_3780,N_3521,N_3568);
nor U3781 (N_3781,N_3604,N_3664);
and U3782 (N_3782,N_3606,N_3641);
nor U3783 (N_3783,N_3528,N_3656);
and U3784 (N_3784,N_3548,N_3522);
and U3785 (N_3785,N_3595,N_3562);
or U3786 (N_3786,N_3561,N_3672);
xnor U3787 (N_3787,N_3667,N_3679);
xor U3788 (N_3788,N_3547,N_3561);
nand U3789 (N_3789,N_3613,N_3646);
nor U3790 (N_3790,N_3541,N_3649);
and U3791 (N_3791,N_3634,N_3522);
and U3792 (N_3792,N_3570,N_3548);
and U3793 (N_3793,N_3673,N_3551);
or U3794 (N_3794,N_3578,N_3622);
nor U3795 (N_3795,N_3643,N_3614);
and U3796 (N_3796,N_3580,N_3651);
xor U3797 (N_3797,N_3637,N_3551);
xor U3798 (N_3798,N_3601,N_3588);
nand U3799 (N_3799,N_3522,N_3626);
nor U3800 (N_3800,N_3609,N_3662);
nor U3801 (N_3801,N_3544,N_3604);
nand U3802 (N_3802,N_3523,N_3643);
or U3803 (N_3803,N_3558,N_3573);
xor U3804 (N_3804,N_3638,N_3590);
and U3805 (N_3805,N_3589,N_3581);
nand U3806 (N_3806,N_3528,N_3610);
nand U3807 (N_3807,N_3583,N_3671);
xor U3808 (N_3808,N_3665,N_3609);
and U3809 (N_3809,N_3655,N_3650);
xor U3810 (N_3810,N_3645,N_3606);
and U3811 (N_3811,N_3547,N_3658);
and U3812 (N_3812,N_3550,N_3597);
nand U3813 (N_3813,N_3599,N_3627);
or U3814 (N_3814,N_3552,N_3646);
xor U3815 (N_3815,N_3556,N_3634);
and U3816 (N_3816,N_3542,N_3533);
or U3817 (N_3817,N_3659,N_3525);
nand U3818 (N_3818,N_3591,N_3578);
and U3819 (N_3819,N_3540,N_3621);
or U3820 (N_3820,N_3601,N_3557);
or U3821 (N_3821,N_3615,N_3640);
or U3822 (N_3822,N_3534,N_3582);
nand U3823 (N_3823,N_3630,N_3671);
nand U3824 (N_3824,N_3659,N_3620);
xor U3825 (N_3825,N_3638,N_3596);
xnor U3826 (N_3826,N_3577,N_3610);
nand U3827 (N_3827,N_3531,N_3616);
nand U3828 (N_3828,N_3545,N_3663);
xnor U3829 (N_3829,N_3578,N_3606);
xor U3830 (N_3830,N_3674,N_3587);
or U3831 (N_3831,N_3598,N_3640);
nand U3832 (N_3832,N_3533,N_3650);
xnor U3833 (N_3833,N_3638,N_3672);
and U3834 (N_3834,N_3572,N_3652);
nand U3835 (N_3835,N_3676,N_3577);
nor U3836 (N_3836,N_3616,N_3639);
xor U3837 (N_3837,N_3654,N_3665);
or U3838 (N_3838,N_3573,N_3566);
xor U3839 (N_3839,N_3599,N_3559);
nor U3840 (N_3840,N_3703,N_3724);
xnor U3841 (N_3841,N_3803,N_3762);
nand U3842 (N_3842,N_3777,N_3827);
and U3843 (N_3843,N_3701,N_3711);
and U3844 (N_3844,N_3794,N_3831);
nand U3845 (N_3845,N_3826,N_3782);
and U3846 (N_3846,N_3742,N_3771);
xor U3847 (N_3847,N_3744,N_3765);
nand U3848 (N_3848,N_3773,N_3787);
xnor U3849 (N_3849,N_3730,N_3761);
xnor U3850 (N_3850,N_3792,N_3752);
nor U3851 (N_3851,N_3784,N_3796);
nand U3852 (N_3852,N_3722,N_3797);
xnor U3853 (N_3853,N_3770,N_3790);
xnor U3854 (N_3854,N_3731,N_3769);
or U3855 (N_3855,N_3830,N_3834);
and U3856 (N_3856,N_3682,N_3727);
and U3857 (N_3857,N_3779,N_3763);
nand U3858 (N_3858,N_3718,N_3819);
nand U3859 (N_3859,N_3814,N_3753);
or U3860 (N_3860,N_3680,N_3820);
xnor U3861 (N_3861,N_3683,N_3800);
or U3862 (N_3862,N_3810,N_3729);
nand U3863 (N_3863,N_3723,N_3710);
and U3864 (N_3864,N_3740,N_3786);
nand U3865 (N_3865,N_3749,N_3738);
nor U3866 (N_3866,N_3766,N_3696);
xor U3867 (N_3867,N_3818,N_3805);
nor U3868 (N_3868,N_3745,N_3747);
and U3869 (N_3869,N_3739,N_3821);
nand U3870 (N_3870,N_3709,N_3833);
or U3871 (N_3871,N_3807,N_3832);
nand U3872 (N_3872,N_3788,N_3695);
nand U3873 (N_3873,N_3697,N_3726);
or U3874 (N_3874,N_3716,N_3717);
nor U3875 (N_3875,N_3715,N_3780);
and U3876 (N_3876,N_3774,N_3746);
nand U3877 (N_3877,N_3760,N_3789);
nor U3878 (N_3878,N_3829,N_3793);
and U3879 (N_3879,N_3692,N_3781);
and U3880 (N_3880,N_3741,N_3836);
or U3881 (N_3881,N_3720,N_3775);
nand U3882 (N_3882,N_3751,N_3733);
or U3883 (N_3883,N_3798,N_3705);
xnor U3884 (N_3884,N_3783,N_3702);
and U3885 (N_3885,N_3725,N_3755);
nand U3886 (N_3886,N_3758,N_3808);
or U3887 (N_3887,N_3838,N_3748);
nor U3888 (N_3888,N_3813,N_3691);
xnor U3889 (N_3889,N_3815,N_3734);
or U3890 (N_3890,N_3809,N_3822);
and U3891 (N_3891,N_3735,N_3700);
nand U3892 (N_3892,N_3686,N_3721);
nor U3893 (N_3893,N_3759,N_3806);
nor U3894 (N_3894,N_3764,N_3736);
or U3895 (N_3895,N_3685,N_3698);
xor U3896 (N_3896,N_3681,N_3835);
nand U3897 (N_3897,N_3699,N_3714);
nand U3898 (N_3898,N_3785,N_3684);
nand U3899 (N_3899,N_3791,N_3778);
nand U3900 (N_3900,N_3706,N_3743);
xnor U3901 (N_3901,N_3690,N_3795);
xnor U3902 (N_3902,N_3776,N_3694);
xor U3903 (N_3903,N_3719,N_3689);
or U3904 (N_3904,N_3767,N_3811);
nor U3905 (N_3905,N_3824,N_3828);
xor U3906 (N_3906,N_3687,N_3802);
or U3907 (N_3907,N_3768,N_3693);
and U3908 (N_3908,N_3707,N_3737);
and U3909 (N_3909,N_3757,N_3728);
and U3910 (N_3910,N_3816,N_3704);
nor U3911 (N_3911,N_3708,N_3837);
or U3912 (N_3912,N_3772,N_3712);
and U3913 (N_3913,N_3750,N_3823);
nor U3914 (N_3914,N_3839,N_3812);
xor U3915 (N_3915,N_3804,N_3688);
and U3916 (N_3916,N_3825,N_3754);
and U3917 (N_3917,N_3756,N_3732);
nor U3918 (N_3918,N_3713,N_3817);
and U3919 (N_3919,N_3799,N_3801);
and U3920 (N_3920,N_3729,N_3803);
xnor U3921 (N_3921,N_3802,N_3810);
or U3922 (N_3922,N_3800,N_3713);
or U3923 (N_3923,N_3780,N_3762);
nand U3924 (N_3924,N_3780,N_3708);
and U3925 (N_3925,N_3694,N_3828);
and U3926 (N_3926,N_3837,N_3759);
or U3927 (N_3927,N_3826,N_3753);
nor U3928 (N_3928,N_3823,N_3729);
and U3929 (N_3929,N_3788,N_3819);
nand U3930 (N_3930,N_3824,N_3776);
nand U3931 (N_3931,N_3693,N_3706);
nand U3932 (N_3932,N_3715,N_3820);
or U3933 (N_3933,N_3835,N_3787);
nand U3934 (N_3934,N_3727,N_3755);
and U3935 (N_3935,N_3752,N_3703);
nor U3936 (N_3936,N_3839,N_3814);
nor U3937 (N_3937,N_3729,N_3757);
or U3938 (N_3938,N_3693,N_3720);
nor U3939 (N_3939,N_3753,N_3817);
xor U3940 (N_3940,N_3681,N_3763);
xnor U3941 (N_3941,N_3688,N_3767);
nand U3942 (N_3942,N_3684,N_3801);
or U3943 (N_3943,N_3762,N_3820);
nor U3944 (N_3944,N_3798,N_3769);
and U3945 (N_3945,N_3794,N_3730);
xor U3946 (N_3946,N_3788,N_3826);
nor U3947 (N_3947,N_3738,N_3789);
or U3948 (N_3948,N_3706,N_3801);
xnor U3949 (N_3949,N_3755,N_3736);
xor U3950 (N_3950,N_3826,N_3762);
or U3951 (N_3951,N_3723,N_3805);
nor U3952 (N_3952,N_3807,N_3751);
nand U3953 (N_3953,N_3791,N_3739);
xnor U3954 (N_3954,N_3727,N_3700);
nand U3955 (N_3955,N_3693,N_3718);
or U3956 (N_3956,N_3772,N_3681);
or U3957 (N_3957,N_3779,N_3724);
nand U3958 (N_3958,N_3836,N_3686);
xnor U3959 (N_3959,N_3680,N_3770);
and U3960 (N_3960,N_3739,N_3755);
and U3961 (N_3961,N_3825,N_3820);
nor U3962 (N_3962,N_3699,N_3726);
nor U3963 (N_3963,N_3695,N_3801);
or U3964 (N_3964,N_3687,N_3735);
and U3965 (N_3965,N_3687,N_3708);
nand U3966 (N_3966,N_3744,N_3824);
nor U3967 (N_3967,N_3774,N_3736);
nor U3968 (N_3968,N_3797,N_3832);
nor U3969 (N_3969,N_3715,N_3799);
nor U3970 (N_3970,N_3837,N_3817);
or U3971 (N_3971,N_3709,N_3752);
nor U3972 (N_3972,N_3755,N_3693);
or U3973 (N_3973,N_3777,N_3821);
xnor U3974 (N_3974,N_3814,N_3816);
or U3975 (N_3975,N_3804,N_3702);
nand U3976 (N_3976,N_3723,N_3739);
nand U3977 (N_3977,N_3732,N_3801);
and U3978 (N_3978,N_3716,N_3815);
and U3979 (N_3979,N_3726,N_3808);
and U3980 (N_3980,N_3793,N_3763);
and U3981 (N_3981,N_3753,N_3787);
and U3982 (N_3982,N_3777,N_3730);
xor U3983 (N_3983,N_3768,N_3802);
nand U3984 (N_3984,N_3697,N_3827);
and U3985 (N_3985,N_3721,N_3734);
xor U3986 (N_3986,N_3700,N_3787);
or U3987 (N_3987,N_3818,N_3727);
or U3988 (N_3988,N_3806,N_3738);
nor U3989 (N_3989,N_3828,N_3685);
and U3990 (N_3990,N_3754,N_3691);
nand U3991 (N_3991,N_3713,N_3693);
nor U3992 (N_3992,N_3835,N_3796);
nand U3993 (N_3993,N_3746,N_3789);
xnor U3994 (N_3994,N_3745,N_3752);
and U3995 (N_3995,N_3830,N_3730);
nand U3996 (N_3996,N_3735,N_3818);
nand U3997 (N_3997,N_3821,N_3747);
or U3998 (N_3998,N_3820,N_3807);
xnor U3999 (N_3999,N_3789,N_3778);
xnor U4000 (N_4000,N_3842,N_3848);
or U4001 (N_4001,N_3973,N_3902);
or U4002 (N_4002,N_3905,N_3878);
and U4003 (N_4003,N_3939,N_3976);
or U4004 (N_4004,N_3850,N_3966);
and U4005 (N_4005,N_3984,N_3950);
nand U4006 (N_4006,N_3868,N_3870);
xnor U4007 (N_4007,N_3864,N_3912);
nor U4008 (N_4008,N_3956,N_3860);
nor U4009 (N_4009,N_3986,N_3847);
and U4010 (N_4010,N_3840,N_3849);
or U4011 (N_4011,N_3994,N_3867);
nand U4012 (N_4012,N_3885,N_3882);
or U4013 (N_4013,N_3856,N_3853);
and U4014 (N_4014,N_3843,N_3858);
xor U4015 (N_4015,N_3958,N_3917);
xnor U4016 (N_4016,N_3933,N_3880);
xor U4017 (N_4017,N_3972,N_3918);
nor U4018 (N_4018,N_3938,N_3895);
nor U4019 (N_4019,N_3996,N_3985);
xnor U4020 (N_4020,N_3990,N_3999);
nand U4021 (N_4021,N_3946,N_3910);
nand U4022 (N_4022,N_3998,N_3906);
xor U4023 (N_4023,N_3965,N_3937);
xor U4024 (N_4024,N_3931,N_3940);
xor U4025 (N_4025,N_3925,N_3873);
nor U4026 (N_4026,N_3963,N_3943);
nor U4027 (N_4027,N_3876,N_3967);
nor U4028 (N_4028,N_3897,N_3989);
and U4029 (N_4029,N_3975,N_3911);
nand U4030 (N_4030,N_3941,N_3899);
and U4031 (N_4031,N_3852,N_3892);
nor U4032 (N_4032,N_3949,N_3907);
or U4033 (N_4033,N_3859,N_3888);
xnor U4034 (N_4034,N_3982,N_3960);
or U4035 (N_4035,N_3898,N_3954);
and U4036 (N_4036,N_3934,N_3924);
and U4037 (N_4037,N_3957,N_3970);
or U4038 (N_4038,N_3865,N_3900);
nor U4039 (N_4039,N_3955,N_3977);
nand U4040 (N_4040,N_3932,N_3862);
or U4041 (N_4041,N_3961,N_3871);
nand U4042 (N_4042,N_3874,N_3971);
nand U4043 (N_4043,N_3863,N_3944);
and U4044 (N_4044,N_3929,N_3968);
nor U4045 (N_4045,N_3980,N_3959);
nand U4046 (N_4046,N_3926,N_3915);
nand U4047 (N_4047,N_3974,N_3869);
xnor U4048 (N_4048,N_3936,N_3845);
xnor U4049 (N_4049,N_3997,N_3904);
or U4050 (N_4050,N_3935,N_3993);
and U4051 (N_4051,N_3881,N_3914);
and U4052 (N_4052,N_3861,N_3893);
or U4053 (N_4053,N_3964,N_3969);
nand U4054 (N_4054,N_3953,N_3992);
or U4055 (N_4055,N_3908,N_3981);
nor U4056 (N_4056,N_3922,N_3841);
nand U4057 (N_4057,N_3879,N_3896);
or U4058 (N_4058,N_3883,N_3890);
nand U4059 (N_4059,N_3979,N_3903);
xnor U4060 (N_4060,N_3952,N_3916);
xor U4061 (N_4061,N_3945,N_3844);
and U4062 (N_4062,N_3991,N_3987);
xor U4063 (N_4063,N_3942,N_3962);
and U4064 (N_4064,N_3919,N_3875);
xnor U4065 (N_4065,N_3983,N_3846);
xnor U4066 (N_4066,N_3889,N_3978);
and U4067 (N_4067,N_3901,N_3886);
nor U4068 (N_4068,N_3872,N_3923);
or U4069 (N_4069,N_3851,N_3928);
and U4070 (N_4070,N_3891,N_3866);
and U4071 (N_4071,N_3947,N_3988);
or U4072 (N_4072,N_3855,N_3920);
and U4073 (N_4073,N_3948,N_3894);
and U4074 (N_4074,N_3921,N_3913);
nand U4075 (N_4075,N_3877,N_3857);
and U4076 (N_4076,N_3951,N_3854);
nor U4077 (N_4077,N_3995,N_3884);
nand U4078 (N_4078,N_3887,N_3927);
and U4079 (N_4079,N_3909,N_3930);
nand U4080 (N_4080,N_3948,N_3951);
xnor U4081 (N_4081,N_3942,N_3913);
nand U4082 (N_4082,N_3916,N_3844);
xnor U4083 (N_4083,N_3840,N_3977);
and U4084 (N_4084,N_3891,N_3886);
and U4085 (N_4085,N_3963,N_3960);
xor U4086 (N_4086,N_3856,N_3963);
or U4087 (N_4087,N_3929,N_3875);
xor U4088 (N_4088,N_3914,N_3843);
nor U4089 (N_4089,N_3981,N_3944);
nand U4090 (N_4090,N_3880,N_3942);
or U4091 (N_4091,N_3875,N_3991);
or U4092 (N_4092,N_3891,N_3880);
and U4093 (N_4093,N_3890,N_3942);
nor U4094 (N_4094,N_3865,N_3976);
xnor U4095 (N_4095,N_3924,N_3893);
nand U4096 (N_4096,N_3928,N_3916);
nor U4097 (N_4097,N_3963,N_3904);
nand U4098 (N_4098,N_3859,N_3889);
nand U4099 (N_4099,N_3981,N_3851);
xor U4100 (N_4100,N_3871,N_3875);
and U4101 (N_4101,N_3883,N_3847);
xnor U4102 (N_4102,N_3985,N_3971);
nand U4103 (N_4103,N_3874,N_3997);
and U4104 (N_4104,N_3990,N_3907);
or U4105 (N_4105,N_3995,N_3906);
and U4106 (N_4106,N_3998,N_3971);
xnor U4107 (N_4107,N_3875,N_3855);
nor U4108 (N_4108,N_3932,N_3867);
nor U4109 (N_4109,N_3943,N_3899);
nor U4110 (N_4110,N_3940,N_3906);
nor U4111 (N_4111,N_3884,N_3989);
or U4112 (N_4112,N_3899,N_3935);
or U4113 (N_4113,N_3898,N_3999);
xor U4114 (N_4114,N_3909,N_3929);
or U4115 (N_4115,N_3913,N_3967);
nor U4116 (N_4116,N_3950,N_3907);
nand U4117 (N_4117,N_3863,N_3854);
nand U4118 (N_4118,N_3905,N_3953);
nor U4119 (N_4119,N_3921,N_3975);
xor U4120 (N_4120,N_3983,N_3947);
nand U4121 (N_4121,N_3972,N_3958);
and U4122 (N_4122,N_3892,N_3929);
nor U4123 (N_4123,N_3879,N_3950);
xnor U4124 (N_4124,N_3986,N_3859);
nand U4125 (N_4125,N_3856,N_3948);
nor U4126 (N_4126,N_3981,N_3998);
and U4127 (N_4127,N_3877,N_3912);
and U4128 (N_4128,N_3964,N_3909);
and U4129 (N_4129,N_3948,N_3891);
nand U4130 (N_4130,N_3953,N_3955);
xor U4131 (N_4131,N_3854,N_3927);
and U4132 (N_4132,N_3970,N_3924);
and U4133 (N_4133,N_3906,N_3922);
nor U4134 (N_4134,N_3882,N_3970);
nand U4135 (N_4135,N_3882,N_3869);
and U4136 (N_4136,N_3995,N_3957);
xnor U4137 (N_4137,N_3944,N_3898);
xor U4138 (N_4138,N_3979,N_3897);
xor U4139 (N_4139,N_3849,N_3889);
and U4140 (N_4140,N_3884,N_3844);
xnor U4141 (N_4141,N_3861,N_3916);
xor U4142 (N_4142,N_3949,N_3987);
nand U4143 (N_4143,N_3997,N_3980);
nand U4144 (N_4144,N_3929,N_3925);
nand U4145 (N_4145,N_3980,N_3961);
nor U4146 (N_4146,N_3938,N_3857);
nand U4147 (N_4147,N_3869,N_3862);
nand U4148 (N_4148,N_3844,N_3876);
nor U4149 (N_4149,N_3963,N_3897);
and U4150 (N_4150,N_3906,N_3858);
nor U4151 (N_4151,N_3868,N_3952);
nor U4152 (N_4152,N_3898,N_3855);
or U4153 (N_4153,N_3881,N_3989);
or U4154 (N_4154,N_3906,N_3956);
nand U4155 (N_4155,N_3928,N_3880);
xnor U4156 (N_4156,N_3994,N_3937);
nand U4157 (N_4157,N_3890,N_3979);
xor U4158 (N_4158,N_3911,N_3866);
or U4159 (N_4159,N_3847,N_3952);
xnor U4160 (N_4160,N_4025,N_4063);
or U4161 (N_4161,N_4080,N_4075);
xnor U4162 (N_4162,N_4147,N_4021);
nand U4163 (N_4163,N_4148,N_4159);
xnor U4164 (N_4164,N_4132,N_4048);
and U4165 (N_4165,N_4098,N_4001);
and U4166 (N_4166,N_4000,N_4109);
nor U4167 (N_4167,N_4122,N_4118);
nand U4168 (N_4168,N_4018,N_4117);
and U4169 (N_4169,N_4125,N_4066);
nand U4170 (N_4170,N_4022,N_4143);
and U4171 (N_4171,N_4090,N_4041);
xor U4172 (N_4172,N_4124,N_4015);
xor U4173 (N_4173,N_4129,N_4131);
and U4174 (N_4174,N_4058,N_4141);
xnor U4175 (N_4175,N_4043,N_4068);
nand U4176 (N_4176,N_4037,N_4042);
or U4177 (N_4177,N_4091,N_4156);
and U4178 (N_4178,N_4086,N_4049);
xnor U4179 (N_4179,N_4111,N_4099);
xor U4180 (N_4180,N_4070,N_4083);
xor U4181 (N_4181,N_4146,N_4060);
nor U4182 (N_4182,N_4084,N_4158);
nor U4183 (N_4183,N_4007,N_4027);
or U4184 (N_4184,N_4039,N_4026);
nor U4185 (N_4185,N_4008,N_4123);
xnor U4186 (N_4186,N_4016,N_4036);
nor U4187 (N_4187,N_4040,N_4020);
nand U4188 (N_4188,N_4009,N_4051);
nand U4189 (N_4189,N_4057,N_4054);
nand U4190 (N_4190,N_4013,N_4137);
nand U4191 (N_4191,N_4116,N_4134);
xor U4192 (N_4192,N_4076,N_4155);
or U4193 (N_4193,N_4050,N_4088);
and U4194 (N_4194,N_4120,N_4014);
nand U4195 (N_4195,N_4130,N_4074);
nand U4196 (N_4196,N_4073,N_4071);
nor U4197 (N_4197,N_4126,N_4085);
nand U4198 (N_4198,N_4062,N_4149);
nand U4199 (N_4199,N_4096,N_4104);
nor U4200 (N_4200,N_4067,N_4002);
or U4201 (N_4201,N_4005,N_4065);
nand U4202 (N_4202,N_4038,N_4028);
nand U4203 (N_4203,N_4072,N_4059);
nand U4204 (N_4204,N_4079,N_4004);
nor U4205 (N_4205,N_4114,N_4077);
xor U4206 (N_4206,N_4144,N_4097);
and U4207 (N_4207,N_4121,N_4105);
nand U4208 (N_4208,N_4157,N_4113);
xnor U4209 (N_4209,N_4064,N_4138);
nor U4210 (N_4210,N_4133,N_4069);
xnor U4211 (N_4211,N_4107,N_4047);
nand U4212 (N_4212,N_4019,N_4082);
and U4213 (N_4213,N_4110,N_4017);
or U4214 (N_4214,N_4151,N_4095);
or U4215 (N_4215,N_4046,N_4093);
or U4216 (N_4216,N_4052,N_4119);
nand U4217 (N_4217,N_4128,N_4100);
nand U4218 (N_4218,N_4103,N_4150);
nand U4219 (N_4219,N_4029,N_4145);
xor U4220 (N_4220,N_4034,N_4035);
and U4221 (N_4221,N_4044,N_4092);
nor U4222 (N_4222,N_4112,N_4106);
or U4223 (N_4223,N_4024,N_4032);
nor U4224 (N_4224,N_4006,N_4089);
or U4225 (N_4225,N_4031,N_4056);
or U4226 (N_4226,N_4135,N_4108);
and U4227 (N_4227,N_4102,N_4053);
xor U4228 (N_4228,N_4139,N_4078);
xor U4229 (N_4229,N_4011,N_4153);
nand U4230 (N_4230,N_4140,N_4152);
nor U4231 (N_4231,N_4045,N_4030);
nand U4232 (N_4232,N_4127,N_4101);
and U4233 (N_4233,N_4012,N_4033);
nand U4234 (N_4234,N_4094,N_4003);
and U4235 (N_4235,N_4136,N_4061);
or U4236 (N_4236,N_4010,N_4055);
xor U4237 (N_4237,N_4023,N_4142);
or U4238 (N_4238,N_4087,N_4154);
nand U4239 (N_4239,N_4081,N_4115);
or U4240 (N_4240,N_4085,N_4036);
nand U4241 (N_4241,N_4142,N_4017);
or U4242 (N_4242,N_4058,N_4112);
and U4243 (N_4243,N_4156,N_4113);
and U4244 (N_4244,N_4065,N_4018);
and U4245 (N_4245,N_4052,N_4090);
or U4246 (N_4246,N_4035,N_4116);
and U4247 (N_4247,N_4007,N_4093);
nand U4248 (N_4248,N_4050,N_4002);
and U4249 (N_4249,N_4096,N_4023);
and U4250 (N_4250,N_4112,N_4097);
nand U4251 (N_4251,N_4142,N_4000);
nand U4252 (N_4252,N_4023,N_4061);
and U4253 (N_4253,N_4133,N_4061);
and U4254 (N_4254,N_4065,N_4030);
xor U4255 (N_4255,N_4071,N_4078);
xnor U4256 (N_4256,N_4094,N_4020);
nor U4257 (N_4257,N_4001,N_4096);
nand U4258 (N_4258,N_4051,N_4159);
or U4259 (N_4259,N_4103,N_4116);
nor U4260 (N_4260,N_4066,N_4111);
nand U4261 (N_4261,N_4148,N_4095);
and U4262 (N_4262,N_4148,N_4003);
xnor U4263 (N_4263,N_4077,N_4001);
xnor U4264 (N_4264,N_4050,N_4043);
or U4265 (N_4265,N_4122,N_4119);
or U4266 (N_4266,N_4044,N_4084);
xor U4267 (N_4267,N_4018,N_4032);
nand U4268 (N_4268,N_4050,N_4107);
or U4269 (N_4269,N_4150,N_4082);
xnor U4270 (N_4270,N_4103,N_4024);
nor U4271 (N_4271,N_4060,N_4108);
nand U4272 (N_4272,N_4063,N_4067);
nand U4273 (N_4273,N_4010,N_4150);
xnor U4274 (N_4274,N_4085,N_4131);
nand U4275 (N_4275,N_4084,N_4140);
xnor U4276 (N_4276,N_4131,N_4143);
nor U4277 (N_4277,N_4021,N_4070);
xnor U4278 (N_4278,N_4030,N_4105);
nand U4279 (N_4279,N_4053,N_4157);
or U4280 (N_4280,N_4024,N_4010);
nor U4281 (N_4281,N_4052,N_4154);
and U4282 (N_4282,N_4154,N_4078);
nor U4283 (N_4283,N_4043,N_4012);
or U4284 (N_4284,N_4081,N_4145);
or U4285 (N_4285,N_4087,N_4116);
or U4286 (N_4286,N_4105,N_4097);
xnor U4287 (N_4287,N_4059,N_4086);
and U4288 (N_4288,N_4084,N_4109);
nor U4289 (N_4289,N_4102,N_4082);
or U4290 (N_4290,N_4042,N_4125);
and U4291 (N_4291,N_4043,N_4128);
xnor U4292 (N_4292,N_4009,N_4091);
nand U4293 (N_4293,N_4010,N_4067);
nor U4294 (N_4294,N_4057,N_4115);
and U4295 (N_4295,N_4034,N_4127);
nand U4296 (N_4296,N_4070,N_4144);
or U4297 (N_4297,N_4013,N_4142);
and U4298 (N_4298,N_4101,N_4106);
or U4299 (N_4299,N_4038,N_4108);
nand U4300 (N_4300,N_4080,N_4014);
or U4301 (N_4301,N_4000,N_4046);
nor U4302 (N_4302,N_4134,N_4051);
nand U4303 (N_4303,N_4021,N_4051);
nand U4304 (N_4304,N_4024,N_4082);
nand U4305 (N_4305,N_4131,N_4119);
nand U4306 (N_4306,N_4132,N_4091);
or U4307 (N_4307,N_4081,N_4156);
and U4308 (N_4308,N_4112,N_4055);
xor U4309 (N_4309,N_4111,N_4058);
nor U4310 (N_4310,N_4010,N_4120);
nor U4311 (N_4311,N_4098,N_4021);
or U4312 (N_4312,N_4119,N_4009);
nand U4313 (N_4313,N_4006,N_4050);
xnor U4314 (N_4314,N_4026,N_4128);
xnor U4315 (N_4315,N_4046,N_4026);
or U4316 (N_4316,N_4075,N_4088);
nand U4317 (N_4317,N_4151,N_4038);
nand U4318 (N_4318,N_4154,N_4152);
and U4319 (N_4319,N_4020,N_4129);
or U4320 (N_4320,N_4311,N_4223);
and U4321 (N_4321,N_4283,N_4255);
or U4322 (N_4322,N_4197,N_4249);
or U4323 (N_4323,N_4240,N_4258);
nand U4324 (N_4324,N_4307,N_4179);
nor U4325 (N_4325,N_4243,N_4186);
xnor U4326 (N_4326,N_4187,N_4199);
and U4327 (N_4327,N_4289,N_4174);
nor U4328 (N_4328,N_4276,N_4294);
nor U4329 (N_4329,N_4252,N_4266);
or U4330 (N_4330,N_4189,N_4182);
nand U4331 (N_4331,N_4278,N_4163);
xor U4332 (N_4332,N_4306,N_4277);
nand U4333 (N_4333,N_4198,N_4268);
nand U4334 (N_4334,N_4195,N_4280);
nor U4335 (N_4335,N_4305,N_4295);
nand U4336 (N_4336,N_4309,N_4260);
nand U4337 (N_4337,N_4253,N_4271);
and U4338 (N_4338,N_4300,N_4217);
nor U4339 (N_4339,N_4211,N_4219);
and U4340 (N_4340,N_4239,N_4287);
nand U4341 (N_4341,N_4191,N_4184);
nor U4342 (N_4342,N_4263,N_4190);
or U4343 (N_4343,N_4227,N_4297);
and U4344 (N_4344,N_4226,N_4284);
nor U4345 (N_4345,N_4233,N_4248);
or U4346 (N_4346,N_4235,N_4232);
or U4347 (N_4347,N_4177,N_4317);
nor U4348 (N_4348,N_4301,N_4230);
or U4349 (N_4349,N_4238,N_4312);
or U4350 (N_4350,N_4242,N_4279);
and U4351 (N_4351,N_4264,N_4194);
or U4352 (N_4352,N_4208,N_4168);
nand U4353 (N_4353,N_4293,N_4218);
nand U4354 (N_4354,N_4161,N_4267);
and U4355 (N_4355,N_4180,N_4178);
and U4356 (N_4356,N_4285,N_4291);
or U4357 (N_4357,N_4196,N_4234);
nand U4358 (N_4358,N_4192,N_4173);
or U4359 (N_4359,N_4273,N_4250);
nor U4360 (N_4360,N_4315,N_4172);
xor U4361 (N_4361,N_4205,N_4310);
nor U4362 (N_4362,N_4188,N_4319);
or U4363 (N_4363,N_4286,N_4222);
or U4364 (N_4364,N_4202,N_4270);
or U4365 (N_4365,N_4251,N_4200);
and U4366 (N_4366,N_4169,N_4170);
or U4367 (N_4367,N_4212,N_4206);
or U4368 (N_4368,N_4210,N_4171);
xor U4369 (N_4369,N_4216,N_4313);
nor U4370 (N_4370,N_4167,N_4245);
xnor U4371 (N_4371,N_4304,N_4308);
xor U4372 (N_4372,N_4176,N_4231);
or U4373 (N_4373,N_4257,N_4274);
xor U4374 (N_4374,N_4213,N_4298);
nor U4375 (N_4375,N_4256,N_4290);
nor U4376 (N_4376,N_4225,N_4224);
nand U4377 (N_4377,N_4201,N_4207);
nor U4378 (N_4378,N_4236,N_4220);
nand U4379 (N_4379,N_4237,N_4316);
nor U4380 (N_4380,N_4275,N_4183);
or U4381 (N_4381,N_4296,N_4318);
nand U4382 (N_4382,N_4303,N_4164);
nand U4383 (N_4383,N_4244,N_4281);
xor U4384 (N_4384,N_4269,N_4292);
or U4385 (N_4385,N_4214,N_4229);
nand U4386 (N_4386,N_4272,N_4162);
and U4387 (N_4387,N_4204,N_4175);
or U4388 (N_4388,N_4209,N_4261);
or U4389 (N_4389,N_4165,N_4160);
and U4390 (N_4390,N_4166,N_4181);
nand U4391 (N_4391,N_4288,N_4185);
or U4392 (N_4392,N_4265,N_4314);
and U4393 (N_4393,N_4282,N_4299);
and U4394 (N_4394,N_4246,N_4193);
nand U4395 (N_4395,N_4228,N_4241);
or U4396 (N_4396,N_4215,N_4254);
nand U4397 (N_4397,N_4221,N_4247);
xor U4398 (N_4398,N_4203,N_4262);
xor U4399 (N_4399,N_4259,N_4302);
nand U4400 (N_4400,N_4289,N_4286);
or U4401 (N_4401,N_4233,N_4179);
nor U4402 (N_4402,N_4249,N_4252);
or U4403 (N_4403,N_4219,N_4272);
and U4404 (N_4404,N_4300,N_4238);
and U4405 (N_4405,N_4272,N_4278);
nand U4406 (N_4406,N_4250,N_4257);
nor U4407 (N_4407,N_4284,N_4270);
nor U4408 (N_4408,N_4266,N_4306);
nor U4409 (N_4409,N_4234,N_4204);
xnor U4410 (N_4410,N_4187,N_4217);
and U4411 (N_4411,N_4164,N_4230);
or U4412 (N_4412,N_4225,N_4189);
xnor U4413 (N_4413,N_4188,N_4256);
or U4414 (N_4414,N_4315,N_4216);
nor U4415 (N_4415,N_4234,N_4165);
or U4416 (N_4416,N_4305,N_4186);
xor U4417 (N_4417,N_4311,N_4274);
nand U4418 (N_4418,N_4245,N_4220);
and U4419 (N_4419,N_4168,N_4224);
or U4420 (N_4420,N_4286,N_4177);
or U4421 (N_4421,N_4288,N_4257);
xnor U4422 (N_4422,N_4310,N_4222);
nor U4423 (N_4423,N_4188,N_4312);
xor U4424 (N_4424,N_4200,N_4301);
xnor U4425 (N_4425,N_4204,N_4178);
nor U4426 (N_4426,N_4237,N_4201);
or U4427 (N_4427,N_4292,N_4239);
nand U4428 (N_4428,N_4216,N_4235);
xor U4429 (N_4429,N_4272,N_4249);
xor U4430 (N_4430,N_4300,N_4185);
and U4431 (N_4431,N_4215,N_4286);
and U4432 (N_4432,N_4247,N_4287);
or U4433 (N_4433,N_4173,N_4221);
xor U4434 (N_4434,N_4283,N_4196);
and U4435 (N_4435,N_4301,N_4222);
or U4436 (N_4436,N_4190,N_4225);
nand U4437 (N_4437,N_4219,N_4278);
xor U4438 (N_4438,N_4193,N_4214);
nor U4439 (N_4439,N_4230,N_4171);
or U4440 (N_4440,N_4169,N_4282);
or U4441 (N_4441,N_4302,N_4253);
or U4442 (N_4442,N_4271,N_4190);
xor U4443 (N_4443,N_4295,N_4262);
nor U4444 (N_4444,N_4163,N_4288);
nand U4445 (N_4445,N_4170,N_4262);
and U4446 (N_4446,N_4199,N_4185);
xor U4447 (N_4447,N_4254,N_4201);
nor U4448 (N_4448,N_4251,N_4196);
nor U4449 (N_4449,N_4287,N_4194);
or U4450 (N_4450,N_4282,N_4291);
xor U4451 (N_4451,N_4208,N_4185);
and U4452 (N_4452,N_4273,N_4297);
or U4453 (N_4453,N_4226,N_4250);
nand U4454 (N_4454,N_4236,N_4244);
xnor U4455 (N_4455,N_4162,N_4274);
nor U4456 (N_4456,N_4316,N_4165);
or U4457 (N_4457,N_4285,N_4179);
or U4458 (N_4458,N_4295,N_4270);
xor U4459 (N_4459,N_4160,N_4249);
or U4460 (N_4460,N_4234,N_4242);
nand U4461 (N_4461,N_4233,N_4267);
nand U4462 (N_4462,N_4187,N_4296);
nor U4463 (N_4463,N_4231,N_4298);
nand U4464 (N_4464,N_4201,N_4302);
and U4465 (N_4465,N_4192,N_4281);
xnor U4466 (N_4466,N_4283,N_4306);
nor U4467 (N_4467,N_4193,N_4231);
xnor U4468 (N_4468,N_4169,N_4209);
and U4469 (N_4469,N_4278,N_4297);
xnor U4470 (N_4470,N_4248,N_4171);
or U4471 (N_4471,N_4201,N_4306);
nor U4472 (N_4472,N_4275,N_4176);
nand U4473 (N_4473,N_4296,N_4181);
xor U4474 (N_4474,N_4237,N_4214);
or U4475 (N_4475,N_4220,N_4223);
or U4476 (N_4476,N_4236,N_4227);
nor U4477 (N_4477,N_4205,N_4210);
and U4478 (N_4478,N_4253,N_4229);
nand U4479 (N_4479,N_4172,N_4199);
nor U4480 (N_4480,N_4388,N_4322);
xnor U4481 (N_4481,N_4363,N_4421);
nand U4482 (N_4482,N_4477,N_4468);
xnor U4483 (N_4483,N_4361,N_4370);
and U4484 (N_4484,N_4359,N_4323);
and U4485 (N_4485,N_4402,N_4331);
xnor U4486 (N_4486,N_4367,N_4466);
or U4487 (N_4487,N_4464,N_4434);
and U4488 (N_4488,N_4471,N_4354);
or U4489 (N_4489,N_4392,N_4460);
nand U4490 (N_4490,N_4357,N_4385);
nor U4491 (N_4491,N_4320,N_4475);
and U4492 (N_4492,N_4458,N_4479);
nor U4493 (N_4493,N_4472,N_4436);
and U4494 (N_4494,N_4336,N_4447);
and U4495 (N_4495,N_4337,N_4412);
nor U4496 (N_4496,N_4400,N_4365);
xor U4497 (N_4497,N_4444,N_4343);
or U4498 (N_4498,N_4457,N_4426);
and U4499 (N_4499,N_4425,N_4362);
or U4500 (N_4500,N_4403,N_4478);
nor U4501 (N_4501,N_4369,N_4470);
or U4502 (N_4502,N_4358,N_4356);
xor U4503 (N_4503,N_4414,N_4465);
or U4504 (N_4504,N_4416,N_4341);
nor U4505 (N_4505,N_4391,N_4374);
nand U4506 (N_4506,N_4404,N_4342);
xnor U4507 (N_4507,N_4340,N_4422);
xnor U4508 (N_4508,N_4372,N_4351);
nor U4509 (N_4509,N_4439,N_4427);
nor U4510 (N_4510,N_4364,N_4383);
and U4511 (N_4511,N_4330,N_4469);
nor U4512 (N_4512,N_4352,N_4454);
and U4513 (N_4513,N_4419,N_4459);
nand U4514 (N_4514,N_4446,N_4455);
xnor U4515 (N_4515,N_4409,N_4355);
and U4516 (N_4516,N_4467,N_4395);
xor U4517 (N_4517,N_4393,N_4329);
or U4518 (N_4518,N_4435,N_4335);
xor U4519 (N_4519,N_4389,N_4324);
or U4520 (N_4520,N_4452,N_4376);
xor U4521 (N_4521,N_4373,N_4417);
nor U4522 (N_4522,N_4440,N_4347);
xnor U4523 (N_4523,N_4390,N_4381);
nand U4524 (N_4524,N_4325,N_4420);
xnor U4525 (N_4525,N_4476,N_4378);
or U4526 (N_4526,N_4406,N_4375);
and U4527 (N_4527,N_4360,N_4451);
xor U4528 (N_4528,N_4349,N_4368);
and U4529 (N_4529,N_4462,N_4411);
xnor U4530 (N_4530,N_4344,N_4430);
and U4531 (N_4531,N_4449,N_4461);
or U4532 (N_4532,N_4334,N_4433);
nand U4533 (N_4533,N_4380,N_4431);
xor U4534 (N_4534,N_4401,N_4410);
nand U4535 (N_4535,N_4398,N_4443);
xnor U4536 (N_4536,N_4438,N_4405);
or U4537 (N_4537,N_4339,N_4327);
nand U4538 (N_4538,N_4453,N_4321);
xor U4539 (N_4539,N_4366,N_4345);
and U4540 (N_4540,N_4397,N_4332);
nand U4541 (N_4541,N_4338,N_4415);
nor U4542 (N_4542,N_4326,N_4386);
or U4543 (N_4543,N_4371,N_4429);
or U4544 (N_4544,N_4445,N_4346);
nand U4545 (N_4545,N_4450,N_4413);
and U4546 (N_4546,N_4387,N_4408);
and U4547 (N_4547,N_4394,N_4353);
nand U4548 (N_4548,N_4456,N_4350);
nor U4549 (N_4549,N_4424,N_4379);
xnor U4550 (N_4550,N_4407,N_4473);
nor U4551 (N_4551,N_4399,N_4442);
and U4552 (N_4552,N_4382,N_4328);
and U4553 (N_4553,N_4384,N_4432);
nand U4554 (N_4554,N_4333,N_4448);
xor U4555 (N_4555,N_4463,N_4348);
xnor U4556 (N_4556,N_4396,N_4423);
or U4557 (N_4557,N_4437,N_4428);
xor U4558 (N_4558,N_4418,N_4377);
or U4559 (N_4559,N_4474,N_4441);
nor U4560 (N_4560,N_4351,N_4428);
nor U4561 (N_4561,N_4461,N_4433);
or U4562 (N_4562,N_4373,N_4478);
or U4563 (N_4563,N_4447,N_4360);
xor U4564 (N_4564,N_4365,N_4402);
xnor U4565 (N_4565,N_4385,N_4457);
and U4566 (N_4566,N_4412,N_4403);
or U4567 (N_4567,N_4448,N_4393);
or U4568 (N_4568,N_4451,N_4478);
nor U4569 (N_4569,N_4363,N_4344);
or U4570 (N_4570,N_4400,N_4359);
or U4571 (N_4571,N_4344,N_4427);
and U4572 (N_4572,N_4469,N_4327);
nand U4573 (N_4573,N_4329,N_4398);
or U4574 (N_4574,N_4362,N_4400);
nor U4575 (N_4575,N_4378,N_4452);
xor U4576 (N_4576,N_4439,N_4422);
or U4577 (N_4577,N_4358,N_4458);
nand U4578 (N_4578,N_4359,N_4325);
nor U4579 (N_4579,N_4412,N_4342);
nor U4580 (N_4580,N_4418,N_4360);
xnor U4581 (N_4581,N_4457,N_4458);
xor U4582 (N_4582,N_4467,N_4331);
nor U4583 (N_4583,N_4444,N_4451);
nand U4584 (N_4584,N_4321,N_4438);
and U4585 (N_4585,N_4363,N_4414);
or U4586 (N_4586,N_4374,N_4443);
or U4587 (N_4587,N_4368,N_4467);
nand U4588 (N_4588,N_4367,N_4462);
nor U4589 (N_4589,N_4374,N_4369);
or U4590 (N_4590,N_4419,N_4386);
and U4591 (N_4591,N_4434,N_4468);
nor U4592 (N_4592,N_4373,N_4370);
and U4593 (N_4593,N_4354,N_4394);
nor U4594 (N_4594,N_4373,N_4466);
nand U4595 (N_4595,N_4362,N_4422);
and U4596 (N_4596,N_4335,N_4427);
nand U4597 (N_4597,N_4425,N_4466);
nand U4598 (N_4598,N_4325,N_4407);
or U4599 (N_4599,N_4456,N_4328);
xnor U4600 (N_4600,N_4336,N_4467);
nor U4601 (N_4601,N_4433,N_4402);
and U4602 (N_4602,N_4365,N_4374);
xor U4603 (N_4603,N_4332,N_4370);
or U4604 (N_4604,N_4341,N_4322);
xor U4605 (N_4605,N_4471,N_4477);
or U4606 (N_4606,N_4442,N_4349);
and U4607 (N_4607,N_4473,N_4390);
xnor U4608 (N_4608,N_4452,N_4338);
nor U4609 (N_4609,N_4350,N_4344);
xor U4610 (N_4610,N_4408,N_4432);
nor U4611 (N_4611,N_4470,N_4438);
nand U4612 (N_4612,N_4351,N_4420);
nor U4613 (N_4613,N_4409,N_4471);
nand U4614 (N_4614,N_4401,N_4408);
xnor U4615 (N_4615,N_4444,N_4438);
nor U4616 (N_4616,N_4464,N_4323);
xor U4617 (N_4617,N_4430,N_4391);
xor U4618 (N_4618,N_4458,N_4456);
and U4619 (N_4619,N_4452,N_4331);
nor U4620 (N_4620,N_4341,N_4373);
nand U4621 (N_4621,N_4410,N_4360);
nand U4622 (N_4622,N_4479,N_4332);
nand U4623 (N_4623,N_4408,N_4366);
nor U4624 (N_4624,N_4365,N_4367);
nand U4625 (N_4625,N_4423,N_4361);
nor U4626 (N_4626,N_4448,N_4412);
nand U4627 (N_4627,N_4330,N_4419);
and U4628 (N_4628,N_4475,N_4344);
and U4629 (N_4629,N_4475,N_4342);
or U4630 (N_4630,N_4321,N_4417);
and U4631 (N_4631,N_4455,N_4458);
or U4632 (N_4632,N_4382,N_4420);
and U4633 (N_4633,N_4391,N_4437);
xnor U4634 (N_4634,N_4455,N_4361);
xor U4635 (N_4635,N_4442,N_4354);
and U4636 (N_4636,N_4363,N_4327);
and U4637 (N_4637,N_4338,N_4368);
nor U4638 (N_4638,N_4403,N_4433);
nand U4639 (N_4639,N_4460,N_4422);
nor U4640 (N_4640,N_4544,N_4541);
nor U4641 (N_4641,N_4561,N_4483);
nand U4642 (N_4642,N_4484,N_4564);
nand U4643 (N_4643,N_4591,N_4542);
and U4644 (N_4644,N_4572,N_4594);
or U4645 (N_4645,N_4620,N_4536);
xor U4646 (N_4646,N_4508,N_4548);
nor U4647 (N_4647,N_4516,N_4543);
nand U4648 (N_4648,N_4610,N_4527);
nor U4649 (N_4649,N_4575,N_4525);
or U4650 (N_4650,N_4517,N_4623);
and U4651 (N_4651,N_4639,N_4530);
nor U4652 (N_4652,N_4574,N_4554);
nor U4653 (N_4653,N_4491,N_4628);
nand U4654 (N_4654,N_4488,N_4563);
xor U4655 (N_4655,N_4606,N_4532);
nor U4656 (N_4656,N_4493,N_4570);
or U4657 (N_4657,N_4630,N_4545);
nor U4658 (N_4658,N_4569,N_4593);
and U4659 (N_4659,N_4513,N_4546);
or U4660 (N_4660,N_4553,N_4596);
or U4661 (N_4661,N_4582,N_4534);
nand U4662 (N_4662,N_4556,N_4528);
xnor U4663 (N_4663,N_4494,N_4565);
or U4664 (N_4664,N_4578,N_4571);
nor U4665 (N_4665,N_4537,N_4637);
nand U4666 (N_4666,N_4634,N_4624);
nand U4667 (N_4667,N_4573,N_4585);
or U4668 (N_4668,N_4502,N_4560);
nor U4669 (N_4669,N_4609,N_4605);
nand U4670 (N_4670,N_4557,N_4566);
and U4671 (N_4671,N_4567,N_4602);
nor U4672 (N_4672,N_4498,N_4601);
nand U4673 (N_4673,N_4616,N_4568);
nor U4674 (N_4674,N_4580,N_4559);
or U4675 (N_4675,N_4581,N_4617);
xnor U4676 (N_4676,N_4501,N_4608);
xor U4677 (N_4677,N_4549,N_4509);
or U4678 (N_4678,N_4495,N_4550);
and U4679 (N_4679,N_4539,N_4551);
nor U4680 (N_4680,N_4636,N_4562);
xnor U4681 (N_4681,N_4535,N_4552);
or U4682 (N_4682,N_4592,N_4506);
nand U4683 (N_4683,N_4529,N_4489);
nor U4684 (N_4684,N_4518,N_4587);
nand U4685 (N_4685,N_4604,N_4597);
xnor U4686 (N_4686,N_4635,N_4621);
or U4687 (N_4687,N_4599,N_4555);
and U4688 (N_4688,N_4531,N_4490);
nor U4689 (N_4689,N_4638,N_4611);
xor U4690 (N_4690,N_4590,N_4607);
xor U4691 (N_4691,N_4503,N_4523);
nor U4692 (N_4692,N_4510,N_4512);
nand U4693 (N_4693,N_4505,N_4586);
or U4694 (N_4694,N_4576,N_4482);
and U4695 (N_4695,N_4507,N_4589);
xor U4696 (N_4696,N_4558,N_4603);
or U4697 (N_4697,N_4492,N_4497);
nand U4698 (N_4698,N_4533,N_4538);
or U4699 (N_4699,N_4579,N_4519);
nor U4700 (N_4700,N_4515,N_4577);
or U4701 (N_4701,N_4588,N_4629);
xnor U4702 (N_4702,N_4522,N_4481);
xor U4703 (N_4703,N_4524,N_4547);
or U4704 (N_4704,N_4584,N_4500);
xor U4705 (N_4705,N_4632,N_4600);
xnor U4706 (N_4706,N_4487,N_4622);
and U4707 (N_4707,N_4499,N_4486);
nor U4708 (N_4708,N_4540,N_4625);
nor U4709 (N_4709,N_4631,N_4598);
nand U4710 (N_4710,N_4514,N_4614);
or U4711 (N_4711,N_4595,N_4619);
xnor U4712 (N_4712,N_4520,N_4521);
xor U4713 (N_4713,N_4511,N_4626);
nand U4714 (N_4714,N_4627,N_4583);
nand U4715 (N_4715,N_4613,N_4633);
xnor U4716 (N_4716,N_4485,N_4615);
and U4717 (N_4717,N_4480,N_4612);
xor U4718 (N_4718,N_4526,N_4504);
nand U4719 (N_4719,N_4496,N_4618);
or U4720 (N_4720,N_4628,N_4518);
nand U4721 (N_4721,N_4543,N_4618);
or U4722 (N_4722,N_4635,N_4634);
xor U4723 (N_4723,N_4631,N_4596);
and U4724 (N_4724,N_4609,N_4491);
or U4725 (N_4725,N_4484,N_4636);
xor U4726 (N_4726,N_4560,N_4606);
or U4727 (N_4727,N_4602,N_4543);
xor U4728 (N_4728,N_4566,N_4545);
and U4729 (N_4729,N_4483,N_4564);
or U4730 (N_4730,N_4550,N_4584);
nand U4731 (N_4731,N_4604,N_4621);
nand U4732 (N_4732,N_4524,N_4560);
nor U4733 (N_4733,N_4597,N_4511);
nand U4734 (N_4734,N_4535,N_4548);
or U4735 (N_4735,N_4493,N_4574);
or U4736 (N_4736,N_4571,N_4495);
nor U4737 (N_4737,N_4489,N_4542);
nand U4738 (N_4738,N_4504,N_4580);
xnor U4739 (N_4739,N_4591,N_4566);
xnor U4740 (N_4740,N_4560,N_4638);
xnor U4741 (N_4741,N_4576,N_4616);
and U4742 (N_4742,N_4485,N_4576);
nand U4743 (N_4743,N_4514,N_4618);
or U4744 (N_4744,N_4593,N_4518);
and U4745 (N_4745,N_4636,N_4584);
and U4746 (N_4746,N_4625,N_4598);
and U4747 (N_4747,N_4600,N_4527);
or U4748 (N_4748,N_4634,N_4516);
or U4749 (N_4749,N_4578,N_4506);
nor U4750 (N_4750,N_4573,N_4513);
or U4751 (N_4751,N_4591,N_4541);
or U4752 (N_4752,N_4562,N_4595);
nand U4753 (N_4753,N_4567,N_4633);
or U4754 (N_4754,N_4484,N_4510);
or U4755 (N_4755,N_4609,N_4511);
xor U4756 (N_4756,N_4563,N_4572);
xnor U4757 (N_4757,N_4523,N_4489);
nor U4758 (N_4758,N_4602,N_4568);
nand U4759 (N_4759,N_4610,N_4544);
xnor U4760 (N_4760,N_4524,N_4624);
and U4761 (N_4761,N_4534,N_4543);
xnor U4762 (N_4762,N_4496,N_4552);
and U4763 (N_4763,N_4623,N_4533);
or U4764 (N_4764,N_4572,N_4622);
or U4765 (N_4765,N_4489,N_4582);
nand U4766 (N_4766,N_4545,N_4539);
nand U4767 (N_4767,N_4522,N_4615);
and U4768 (N_4768,N_4575,N_4522);
nor U4769 (N_4769,N_4529,N_4509);
nor U4770 (N_4770,N_4606,N_4618);
nor U4771 (N_4771,N_4587,N_4548);
nor U4772 (N_4772,N_4532,N_4497);
xor U4773 (N_4773,N_4491,N_4570);
and U4774 (N_4774,N_4569,N_4574);
or U4775 (N_4775,N_4606,N_4520);
xnor U4776 (N_4776,N_4541,N_4518);
and U4777 (N_4777,N_4628,N_4555);
xnor U4778 (N_4778,N_4487,N_4620);
or U4779 (N_4779,N_4623,N_4522);
and U4780 (N_4780,N_4625,N_4525);
nand U4781 (N_4781,N_4626,N_4560);
and U4782 (N_4782,N_4621,N_4583);
or U4783 (N_4783,N_4498,N_4585);
nand U4784 (N_4784,N_4586,N_4610);
nor U4785 (N_4785,N_4580,N_4585);
nand U4786 (N_4786,N_4626,N_4517);
nor U4787 (N_4787,N_4481,N_4552);
or U4788 (N_4788,N_4639,N_4606);
or U4789 (N_4789,N_4634,N_4629);
nand U4790 (N_4790,N_4584,N_4484);
nor U4791 (N_4791,N_4516,N_4605);
or U4792 (N_4792,N_4596,N_4637);
nand U4793 (N_4793,N_4564,N_4560);
xnor U4794 (N_4794,N_4536,N_4590);
nand U4795 (N_4795,N_4591,N_4519);
and U4796 (N_4796,N_4580,N_4634);
and U4797 (N_4797,N_4524,N_4485);
and U4798 (N_4798,N_4574,N_4502);
or U4799 (N_4799,N_4612,N_4598);
and U4800 (N_4800,N_4767,N_4729);
xor U4801 (N_4801,N_4662,N_4770);
nor U4802 (N_4802,N_4739,N_4671);
nand U4803 (N_4803,N_4711,N_4656);
nor U4804 (N_4804,N_4670,N_4666);
and U4805 (N_4805,N_4645,N_4728);
nand U4806 (N_4806,N_4693,N_4796);
nor U4807 (N_4807,N_4753,N_4771);
and U4808 (N_4808,N_4741,N_4734);
nand U4809 (N_4809,N_4648,N_4651);
or U4810 (N_4810,N_4777,N_4669);
nand U4811 (N_4811,N_4680,N_4794);
or U4812 (N_4812,N_4756,N_4791);
nor U4813 (N_4813,N_4712,N_4726);
or U4814 (N_4814,N_4682,N_4787);
nor U4815 (N_4815,N_4719,N_4774);
xnor U4816 (N_4816,N_4642,N_4709);
xor U4817 (N_4817,N_4676,N_4701);
nor U4818 (N_4818,N_4768,N_4754);
xor U4819 (N_4819,N_4647,N_4673);
xnor U4820 (N_4820,N_4749,N_4686);
and U4821 (N_4821,N_4762,N_4688);
nand U4822 (N_4822,N_4748,N_4699);
xnor U4823 (N_4823,N_4653,N_4740);
nor U4824 (N_4824,N_4786,N_4717);
nor U4825 (N_4825,N_4720,N_4722);
or U4826 (N_4826,N_4759,N_4750);
xor U4827 (N_4827,N_4696,N_4674);
or U4828 (N_4828,N_4657,N_4658);
or U4829 (N_4829,N_4714,N_4725);
and U4830 (N_4830,N_4691,N_4751);
nor U4831 (N_4831,N_4705,N_4763);
or U4832 (N_4832,N_4778,N_4640);
and U4833 (N_4833,N_4667,N_4732);
and U4834 (N_4834,N_4795,N_4681);
and U4835 (N_4835,N_4797,N_4746);
xor U4836 (N_4836,N_4735,N_4769);
nand U4837 (N_4837,N_4702,N_4718);
and U4838 (N_4838,N_4788,N_4672);
nor U4839 (N_4839,N_4742,N_4697);
nand U4840 (N_4840,N_4689,N_4773);
xor U4841 (N_4841,N_4747,N_4780);
xnor U4842 (N_4842,N_4687,N_4781);
xor U4843 (N_4843,N_4761,N_4721);
xor U4844 (N_4844,N_4695,N_4752);
and U4845 (N_4845,N_4760,N_4664);
nor U4846 (N_4846,N_4785,N_4736);
nor U4847 (N_4847,N_4779,N_4799);
nand U4848 (N_4848,N_4743,N_4793);
and U4849 (N_4849,N_4663,N_4744);
or U4850 (N_4850,N_4703,N_4641);
xor U4851 (N_4851,N_4652,N_4792);
nor U4852 (N_4852,N_4710,N_4668);
nand U4853 (N_4853,N_4650,N_4757);
nor U4854 (N_4854,N_4683,N_4655);
xor U4855 (N_4855,N_4776,N_4772);
xnor U4856 (N_4856,N_4775,N_4708);
nand U4857 (N_4857,N_4755,N_4764);
and U4858 (N_4858,N_4692,N_4716);
and U4859 (N_4859,N_4738,N_4707);
nand U4860 (N_4860,N_4789,N_4727);
and U4861 (N_4861,N_4715,N_4706);
and U4862 (N_4862,N_4731,N_4790);
xnor U4863 (N_4863,N_4733,N_4643);
xnor U4864 (N_4864,N_4737,N_4690);
and U4865 (N_4865,N_4685,N_4649);
and U4866 (N_4866,N_4758,N_4660);
nand U4867 (N_4867,N_4675,N_4766);
and U4868 (N_4868,N_4783,N_4782);
nand U4869 (N_4869,N_4724,N_4698);
or U4870 (N_4870,N_4704,N_4677);
nand U4871 (N_4871,N_4659,N_4694);
xor U4872 (N_4872,N_4713,N_4654);
nand U4873 (N_4873,N_4784,N_4665);
or U4874 (N_4874,N_4730,N_4745);
nor U4875 (N_4875,N_4679,N_4684);
or U4876 (N_4876,N_4661,N_4644);
xor U4877 (N_4877,N_4646,N_4700);
nor U4878 (N_4878,N_4765,N_4798);
or U4879 (N_4879,N_4678,N_4723);
nand U4880 (N_4880,N_4763,N_4663);
nand U4881 (N_4881,N_4786,N_4759);
nand U4882 (N_4882,N_4703,N_4640);
xnor U4883 (N_4883,N_4642,N_4734);
or U4884 (N_4884,N_4777,N_4704);
xor U4885 (N_4885,N_4701,N_4719);
nand U4886 (N_4886,N_4799,N_4734);
nor U4887 (N_4887,N_4713,N_4645);
and U4888 (N_4888,N_4767,N_4697);
or U4889 (N_4889,N_4789,N_4772);
nand U4890 (N_4890,N_4696,N_4772);
nor U4891 (N_4891,N_4643,N_4783);
nor U4892 (N_4892,N_4740,N_4696);
nand U4893 (N_4893,N_4713,N_4738);
nand U4894 (N_4894,N_4745,N_4687);
nor U4895 (N_4895,N_4708,N_4787);
xnor U4896 (N_4896,N_4723,N_4798);
nor U4897 (N_4897,N_4703,N_4654);
xor U4898 (N_4898,N_4653,N_4794);
and U4899 (N_4899,N_4765,N_4744);
xnor U4900 (N_4900,N_4649,N_4713);
nor U4901 (N_4901,N_4690,N_4675);
and U4902 (N_4902,N_4754,N_4707);
or U4903 (N_4903,N_4696,N_4687);
xnor U4904 (N_4904,N_4658,N_4691);
and U4905 (N_4905,N_4760,N_4653);
nand U4906 (N_4906,N_4766,N_4746);
and U4907 (N_4907,N_4717,N_4646);
xor U4908 (N_4908,N_4647,N_4728);
nand U4909 (N_4909,N_4741,N_4671);
xor U4910 (N_4910,N_4679,N_4759);
nand U4911 (N_4911,N_4783,N_4745);
xnor U4912 (N_4912,N_4764,N_4773);
nand U4913 (N_4913,N_4766,N_4733);
xor U4914 (N_4914,N_4782,N_4781);
nor U4915 (N_4915,N_4738,N_4690);
and U4916 (N_4916,N_4783,N_4784);
nand U4917 (N_4917,N_4660,N_4654);
nand U4918 (N_4918,N_4793,N_4765);
and U4919 (N_4919,N_4653,N_4727);
and U4920 (N_4920,N_4784,N_4777);
or U4921 (N_4921,N_4686,N_4741);
nor U4922 (N_4922,N_4702,N_4671);
nor U4923 (N_4923,N_4692,N_4739);
and U4924 (N_4924,N_4757,N_4794);
or U4925 (N_4925,N_4644,N_4649);
or U4926 (N_4926,N_4733,N_4767);
and U4927 (N_4927,N_4723,N_4704);
nand U4928 (N_4928,N_4796,N_4797);
nor U4929 (N_4929,N_4714,N_4731);
and U4930 (N_4930,N_4781,N_4739);
or U4931 (N_4931,N_4772,N_4785);
xnor U4932 (N_4932,N_4649,N_4737);
nand U4933 (N_4933,N_4667,N_4727);
and U4934 (N_4934,N_4672,N_4722);
or U4935 (N_4935,N_4676,N_4753);
xor U4936 (N_4936,N_4764,N_4784);
and U4937 (N_4937,N_4665,N_4723);
nor U4938 (N_4938,N_4757,N_4735);
nor U4939 (N_4939,N_4776,N_4774);
nor U4940 (N_4940,N_4754,N_4735);
xnor U4941 (N_4941,N_4702,N_4649);
nand U4942 (N_4942,N_4761,N_4765);
nand U4943 (N_4943,N_4756,N_4766);
or U4944 (N_4944,N_4645,N_4792);
xnor U4945 (N_4945,N_4677,N_4681);
and U4946 (N_4946,N_4716,N_4651);
nand U4947 (N_4947,N_4673,N_4740);
nor U4948 (N_4948,N_4678,N_4688);
or U4949 (N_4949,N_4717,N_4647);
nand U4950 (N_4950,N_4743,N_4668);
and U4951 (N_4951,N_4797,N_4686);
nand U4952 (N_4952,N_4751,N_4776);
nand U4953 (N_4953,N_4697,N_4669);
and U4954 (N_4954,N_4774,N_4769);
xor U4955 (N_4955,N_4696,N_4735);
nor U4956 (N_4956,N_4788,N_4658);
xnor U4957 (N_4957,N_4679,N_4694);
nor U4958 (N_4958,N_4714,N_4656);
xnor U4959 (N_4959,N_4765,N_4737);
and U4960 (N_4960,N_4907,N_4944);
nor U4961 (N_4961,N_4841,N_4810);
and U4962 (N_4962,N_4865,N_4846);
and U4963 (N_4963,N_4870,N_4850);
nor U4964 (N_4964,N_4940,N_4834);
or U4965 (N_4965,N_4819,N_4913);
or U4966 (N_4966,N_4882,N_4879);
and U4967 (N_4967,N_4847,N_4875);
or U4968 (N_4968,N_4895,N_4933);
nand U4969 (N_4969,N_4936,N_4904);
nor U4970 (N_4970,N_4874,N_4830);
nor U4971 (N_4971,N_4941,N_4843);
xor U4972 (N_4972,N_4837,N_4833);
nor U4973 (N_4973,N_4923,N_4884);
nand U4974 (N_4974,N_4948,N_4937);
and U4975 (N_4975,N_4854,N_4823);
xnor U4976 (N_4976,N_4954,N_4851);
and U4977 (N_4977,N_4886,N_4832);
nand U4978 (N_4978,N_4950,N_4845);
and U4979 (N_4979,N_4826,N_4909);
nor U4980 (N_4980,N_4932,N_4888);
xnor U4981 (N_4981,N_4828,N_4947);
nor U4982 (N_4982,N_4929,N_4956);
and U4983 (N_4983,N_4926,N_4800);
or U4984 (N_4984,N_4928,N_4910);
nor U4985 (N_4985,N_4939,N_4957);
nor U4986 (N_4986,N_4822,N_4942);
nor U4987 (N_4987,N_4927,N_4838);
and U4988 (N_4988,N_4938,N_4801);
nand U4989 (N_4989,N_4859,N_4813);
and U4990 (N_4990,N_4815,N_4809);
nand U4991 (N_4991,N_4821,N_4849);
xor U4992 (N_4992,N_4871,N_4931);
nor U4993 (N_4993,N_4864,N_4958);
and U4994 (N_4994,N_4839,N_4860);
xnor U4995 (N_4995,N_4921,N_4869);
xnor U4996 (N_4996,N_4827,N_4959);
xnor U4997 (N_4997,N_4872,N_4807);
nor U4998 (N_4998,N_4912,N_4906);
or U4999 (N_4999,N_4891,N_4855);
nand U5000 (N_5000,N_4914,N_4862);
or U5001 (N_5001,N_4935,N_4951);
and U5002 (N_5002,N_4863,N_4840);
nor U5003 (N_5003,N_4892,N_4848);
or U5004 (N_5004,N_4812,N_4878);
or U5005 (N_5005,N_4901,N_4803);
or U5006 (N_5006,N_4861,N_4804);
or U5007 (N_5007,N_4818,N_4955);
or U5008 (N_5008,N_4805,N_4814);
nand U5009 (N_5009,N_4946,N_4896);
nand U5010 (N_5010,N_4816,N_4877);
nor U5011 (N_5011,N_4842,N_4918);
and U5012 (N_5012,N_4873,N_4857);
xor U5013 (N_5013,N_4922,N_4953);
or U5014 (N_5014,N_4903,N_4916);
xnor U5015 (N_5015,N_4889,N_4945);
xor U5016 (N_5016,N_4852,N_4887);
xor U5017 (N_5017,N_4808,N_4915);
xor U5018 (N_5018,N_4917,N_4911);
and U5019 (N_5019,N_4924,N_4893);
nand U5020 (N_5020,N_4806,N_4876);
and U5021 (N_5021,N_4949,N_4899);
or U5022 (N_5022,N_4898,N_4824);
or U5023 (N_5023,N_4890,N_4934);
nand U5024 (N_5024,N_4925,N_4902);
and U5025 (N_5025,N_4908,N_4868);
nor U5026 (N_5026,N_4858,N_4866);
or U5027 (N_5027,N_4829,N_4880);
nand U5028 (N_5028,N_4811,N_4920);
and U5029 (N_5029,N_4952,N_4856);
or U5030 (N_5030,N_4897,N_4943);
nor U5031 (N_5031,N_4825,N_4817);
and U5032 (N_5032,N_4844,N_4867);
nor U5033 (N_5033,N_4883,N_4885);
nor U5034 (N_5034,N_4836,N_4881);
nor U5035 (N_5035,N_4820,N_4835);
xnor U5036 (N_5036,N_4853,N_4802);
nand U5037 (N_5037,N_4919,N_4894);
xnor U5038 (N_5038,N_4905,N_4831);
nand U5039 (N_5039,N_4930,N_4900);
nor U5040 (N_5040,N_4808,N_4860);
nand U5041 (N_5041,N_4936,N_4875);
nand U5042 (N_5042,N_4873,N_4904);
xor U5043 (N_5043,N_4850,N_4843);
and U5044 (N_5044,N_4874,N_4952);
and U5045 (N_5045,N_4940,N_4888);
or U5046 (N_5046,N_4881,N_4928);
and U5047 (N_5047,N_4897,N_4861);
xor U5048 (N_5048,N_4888,N_4824);
nor U5049 (N_5049,N_4803,N_4940);
and U5050 (N_5050,N_4935,N_4810);
nand U5051 (N_5051,N_4894,N_4926);
or U5052 (N_5052,N_4828,N_4821);
and U5053 (N_5053,N_4953,N_4897);
nand U5054 (N_5054,N_4803,N_4855);
or U5055 (N_5055,N_4871,N_4807);
and U5056 (N_5056,N_4830,N_4951);
xor U5057 (N_5057,N_4949,N_4826);
or U5058 (N_5058,N_4875,N_4873);
xnor U5059 (N_5059,N_4860,N_4813);
or U5060 (N_5060,N_4929,N_4897);
or U5061 (N_5061,N_4822,N_4828);
or U5062 (N_5062,N_4912,N_4930);
nand U5063 (N_5063,N_4870,N_4908);
xor U5064 (N_5064,N_4874,N_4939);
or U5065 (N_5065,N_4926,N_4802);
or U5066 (N_5066,N_4907,N_4874);
nor U5067 (N_5067,N_4868,N_4830);
nand U5068 (N_5068,N_4922,N_4950);
and U5069 (N_5069,N_4941,N_4926);
and U5070 (N_5070,N_4844,N_4933);
nor U5071 (N_5071,N_4840,N_4934);
xnor U5072 (N_5072,N_4929,N_4825);
nor U5073 (N_5073,N_4951,N_4810);
nand U5074 (N_5074,N_4935,N_4928);
and U5075 (N_5075,N_4936,N_4924);
or U5076 (N_5076,N_4814,N_4889);
xnor U5077 (N_5077,N_4870,N_4884);
nand U5078 (N_5078,N_4884,N_4803);
xor U5079 (N_5079,N_4891,N_4801);
nand U5080 (N_5080,N_4932,N_4841);
nand U5081 (N_5081,N_4935,N_4896);
and U5082 (N_5082,N_4916,N_4862);
nor U5083 (N_5083,N_4812,N_4957);
nor U5084 (N_5084,N_4899,N_4861);
xor U5085 (N_5085,N_4851,N_4870);
xor U5086 (N_5086,N_4882,N_4908);
and U5087 (N_5087,N_4893,N_4816);
and U5088 (N_5088,N_4851,N_4829);
xnor U5089 (N_5089,N_4914,N_4887);
nand U5090 (N_5090,N_4911,N_4820);
xnor U5091 (N_5091,N_4897,N_4915);
nor U5092 (N_5092,N_4880,N_4921);
xor U5093 (N_5093,N_4825,N_4839);
and U5094 (N_5094,N_4923,N_4912);
xor U5095 (N_5095,N_4885,N_4889);
or U5096 (N_5096,N_4901,N_4826);
nand U5097 (N_5097,N_4921,N_4933);
or U5098 (N_5098,N_4847,N_4811);
or U5099 (N_5099,N_4880,N_4841);
nand U5100 (N_5100,N_4943,N_4827);
and U5101 (N_5101,N_4813,N_4955);
nand U5102 (N_5102,N_4910,N_4924);
xnor U5103 (N_5103,N_4909,N_4800);
nand U5104 (N_5104,N_4952,N_4899);
nor U5105 (N_5105,N_4924,N_4917);
and U5106 (N_5106,N_4901,N_4917);
nor U5107 (N_5107,N_4871,N_4914);
nor U5108 (N_5108,N_4805,N_4920);
nor U5109 (N_5109,N_4874,N_4892);
xor U5110 (N_5110,N_4887,N_4922);
nand U5111 (N_5111,N_4909,N_4832);
nor U5112 (N_5112,N_4830,N_4870);
or U5113 (N_5113,N_4882,N_4922);
nor U5114 (N_5114,N_4959,N_4958);
nand U5115 (N_5115,N_4821,N_4953);
and U5116 (N_5116,N_4945,N_4878);
and U5117 (N_5117,N_4828,N_4944);
xnor U5118 (N_5118,N_4877,N_4909);
nor U5119 (N_5119,N_4801,N_4824);
nor U5120 (N_5120,N_4990,N_5070);
or U5121 (N_5121,N_5004,N_5097);
xor U5122 (N_5122,N_5071,N_5093);
nor U5123 (N_5123,N_5040,N_5056);
nor U5124 (N_5124,N_4976,N_4968);
nand U5125 (N_5125,N_5008,N_5047);
and U5126 (N_5126,N_5058,N_5082);
and U5127 (N_5127,N_5061,N_5030);
and U5128 (N_5128,N_4973,N_4988);
and U5129 (N_5129,N_5081,N_5089);
or U5130 (N_5130,N_4978,N_5118);
and U5131 (N_5131,N_5038,N_5067);
and U5132 (N_5132,N_5087,N_5112);
or U5133 (N_5133,N_5031,N_5104);
or U5134 (N_5134,N_5057,N_5079);
and U5135 (N_5135,N_5003,N_5105);
nor U5136 (N_5136,N_5043,N_5010);
and U5137 (N_5137,N_5012,N_4992);
or U5138 (N_5138,N_4977,N_4974);
nor U5139 (N_5139,N_4981,N_5090);
or U5140 (N_5140,N_5014,N_4994);
nor U5141 (N_5141,N_5078,N_5054);
or U5142 (N_5142,N_4960,N_5013);
or U5143 (N_5143,N_5033,N_5052);
nand U5144 (N_5144,N_4969,N_5044);
nand U5145 (N_5145,N_4983,N_5002);
nor U5146 (N_5146,N_5066,N_5034);
nor U5147 (N_5147,N_4961,N_5045);
nand U5148 (N_5148,N_5111,N_4999);
and U5149 (N_5149,N_5072,N_5108);
and U5150 (N_5150,N_5059,N_5060);
and U5151 (N_5151,N_4998,N_5019);
xnor U5152 (N_5152,N_5009,N_5102);
and U5153 (N_5153,N_5063,N_4984);
nand U5154 (N_5154,N_5021,N_4964);
and U5155 (N_5155,N_5015,N_5035);
and U5156 (N_5156,N_5088,N_5098);
nor U5157 (N_5157,N_4971,N_5049);
xnor U5158 (N_5158,N_5101,N_5023);
nand U5159 (N_5159,N_5116,N_5017);
nor U5160 (N_5160,N_5053,N_5022);
nand U5161 (N_5161,N_4975,N_4967);
and U5162 (N_5162,N_5007,N_4962);
and U5163 (N_5163,N_5115,N_4995);
and U5164 (N_5164,N_5074,N_5037);
xor U5165 (N_5165,N_5099,N_5027);
xor U5166 (N_5166,N_4993,N_5064);
and U5167 (N_5167,N_5011,N_5086);
xor U5168 (N_5168,N_5041,N_5000);
nand U5169 (N_5169,N_5069,N_5096);
xnor U5170 (N_5170,N_4965,N_5028);
and U5171 (N_5171,N_5032,N_5062);
or U5172 (N_5172,N_5110,N_5076);
nand U5173 (N_5173,N_5048,N_5085);
nand U5174 (N_5174,N_5001,N_4982);
nor U5175 (N_5175,N_5077,N_5106);
and U5176 (N_5176,N_5113,N_4997);
or U5177 (N_5177,N_5018,N_5091);
nor U5178 (N_5178,N_5095,N_4963);
xnor U5179 (N_5179,N_5094,N_4980);
and U5180 (N_5180,N_4972,N_5065);
nor U5181 (N_5181,N_4991,N_5046);
nor U5182 (N_5182,N_5107,N_5075);
and U5183 (N_5183,N_4986,N_5092);
nand U5184 (N_5184,N_5114,N_5100);
and U5185 (N_5185,N_4979,N_5024);
nor U5186 (N_5186,N_5036,N_5025);
xnor U5187 (N_5187,N_5039,N_5026);
xor U5188 (N_5188,N_5103,N_5084);
or U5189 (N_5189,N_5016,N_4989);
nand U5190 (N_5190,N_5083,N_5109);
and U5191 (N_5191,N_5042,N_5073);
or U5192 (N_5192,N_4996,N_4987);
and U5193 (N_5193,N_5051,N_4966);
nand U5194 (N_5194,N_5005,N_5006);
and U5195 (N_5195,N_5050,N_5068);
nor U5196 (N_5196,N_5117,N_5029);
or U5197 (N_5197,N_5119,N_5055);
xor U5198 (N_5198,N_5080,N_5020);
xnor U5199 (N_5199,N_4985,N_4970);
nand U5200 (N_5200,N_5097,N_5038);
and U5201 (N_5201,N_5080,N_5102);
or U5202 (N_5202,N_5063,N_5051);
nor U5203 (N_5203,N_5059,N_5015);
nor U5204 (N_5204,N_5050,N_5038);
xnor U5205 (N_5205,N_4972,N_5115);
nor U5206 (N_5206,N_4969,N_5023);
or U5207 (N_5207,N_5092,N_5016);
and U5208 (N_5208,N_5078,N_5020);
or U5209 (N_5209,N_5003,N_5040);
or U5210 (N_5210,N_4985,N_5005);
nor U5211 (N_5211,N_5029,N_4961);
or U5212 (N_5212,N_5091,N_5102);
nand U5213 (N_5213,N_5052,N_4996);
or U5214 (N_5214,N_5005,N_5064);
nor U5215 (N_5215,N_5006,N_4970);
nor U5216 (N_5216,N_4988,N_5108);
nor U5217 (N_5217,N_5051,N_5058);
nand U5218 (N_5218,N_5046,N_5052);
or U5219 (N_5219,N_4978,N_5097);
and U5220 (N_5220,N_5024,N_5038);
and U5221 (N_5221,N_5093,N_5108);
nor U5222 (N_5222,N_4975,N_5114);
nor U5223 (N_5223,N_5107,N_4991);
nand U5224 (N_5224,N_5107,N_5002);
nand U5225 (N_5225,N_5093,N_5041);
or U5226 (N_5226,N_5023,N_4989);
xnor U5227 (N_5227,N_4961,N_4972);
xor U5228 (N_5228,N_5028,N_4966);
xor U5229 (N_5229,N_4997,N_5014);
or U5230 (N_5230,N_5015,N_5088);
and U5231 (N_5231,N_5078,N_5071);
and U5232 (N_5232,N_5097,N_5040);
or U5233 (N_5233,N_5056,N_5037);
or U5234 (N_5234,N_5027,N_5040);
nand U5235 (N_5235,N_4995,N_5021);
nor U5236 (N_5236,N_5070,N_4993);
nand U5237 (N_5237,N_5100,N_4968);
xor U5238 (N_5238,N_5083,N_5047);
or U5239 (N_5239,N_5003,N_5089);
or U5240 (N_5240,N_5012,N_4966);
or U5241 (N_5241,N_4972,N_5029);
nor U5242 (N_5242,N_4986,N_4973);
nand U5243 (N_5243,N_5061,N_5100);
nand U5244 (N_5244,N_4984,N_4969);
and U5245 (N_5245,N_5008,N_5107);
nand U5246 (N_5246,N_5038,N_5074);
xor U5247 (N_5247,N_5012,N_5103);
nor U5248 (N_5248,N_5065,N_5108);
xnor U5249 (N_5249,N_4995,N_5069);
and U5250 (N_5250,N_5004,N_5052);
xor U5251 (N_5251,N_5060,N_5040);
xor U5252 (N_5252,N_4976,N_5009);
nor U5253 (N_5253,N_5055,N_5047);
nand U5254 (N_5254,N_4979,N_5018);
nor U5255 (N_5255,N_5115,N_4985);
nand U5256 (N_5256,N_5047,N_4960);
or U5257 (N_5257,N_5096,N_5003);
nand U5258 (N_5258,N_5093,N_4994);
or U5259 (N_5259,N_5091,N_4977);
nand U5260 (N_5260,N_4974,N_5059);
and U5261 (N_5261,N_4968,N_5065);
nor U5262 (N_5262,N_5025,N_5102);
and U5263 (N_5263,N_5058,N_5048);
nor U5264 (N_5264,N_5097,N_5051);
nand U5265 (N_5265,N_5025,N_5013);
and U5266 (N_5266,N_5101,N_5091);
or U5267 (N_5267,N_5039,N_4969);
or U5268 (N_5268,N_5118,N_5067);
xnor U5269 (N_5269,N_4967,N_4989);
nand U5270 (N_5270,N_5095,N_5092);
nor U5271 (N_5271,N_4995,N_5074);
nor U5272 (N_5272,N_5069,N_5008);
or U5273 (N_5273,N_5105,N_5103);
and U5274 (N_5274,N_5110,N_5055);
or U5275 (N_5275,N_4973,N_5104);
nor U5276 (N_5276,N_5042,N_5049);
or U5277 (N_5277,N_5022,N_5020);
and U5278 (N_5278,N_5005,N_5033);
nand U5279 (N_5279,N_5052,N_5067);
or U5280 (N_5280,N_5218,N_5272);
and U5281 (N_5281,N_5246,N_5128);
xor U5282 (N_5282,N_5160,N_5194);
or U5283 (N_5283,N_5209,N_5240);
xnor U5284 (N_5284,N_5261,N_5135);
xnor U5285 (N_5285,N_5239,N_5174);
xnor U5286 (N_5286,N_5200,N_5179);
xnor U5287 (N_5287,N_5274,N_5185);
xnor U5288 (N_5288,N_5196,N_5172);
nor U5289 (N_5289,N_5173,N_5182);
or U5290 (N_5290,N_5247,N_5217);
nor U5291 (N_5291,N_5277,N_5276);
xor U5292 (N_5292,N_5273,N_5165);
and U5293 (N_5293,N_5213,N_5251);
and U5294 (N_5294,N_5186,N_5188);
and U5295 (N_5295,N_5171,N_5221);
xnor U5296 (N_5296,N_5145,N_5159);
nor U5297 (N_5297,N_5219,N_5190);
nand U5298 (N_5298,N_5270,N_5214);
nor U5299 (N_5299,N_5131,N_5252);
or U5300 (N_5300,N_5170,N_5279);
nor U5301 (N_5301,N_5138,N_5268);
nand U5302 (N_5302,N_5226,N_5258);
nand U5303 (N_5303,N_5167,N_5208);
and U5304 (N_5304,N_5123,N_5233);
or U5305 (N_5305,N_5275,N_5205);
xnor U5306 (N_5306,N_5125,N_5155);
xnor U5307 (N_5307,N_5147,N_5154);
nor U5308 (N_5308,N_5262,N_5121);
or U5309 (N_5309,N_5151,N_5265);
and U5310 (N_5310,N_5169,N_5212);
and U5311 (N_5311,N_5161,N_5242);
nand U5312 (N_5312,N_5253,N_5143);
xor U5313 (N_5313,N_5207,N_5178);
and U5314 (N_5314,N_5193,N_5223);
nor U5315 (N_5315,N_5263,N_5140);
nor U5316 (N_5316,N_5231,N_5235);
or U5317 (N_5317,N_5199,N_5237);
or U5318 (N_5318,N_5177,N_5228);
or U5319 (N_5319,N_5148,N_5243);
nand U5320 (N_5320,N_5198,N_5126);
xnor U5321 (N_5321,N_5271,N_5144);
and U5322 (N_5322,N_5176,N_5163);
and U5323 (N_5323,N_5156,N_5211);
or U5324 (N_5324,N_5254,N_5189);
nand U5325 (N_5325,N_5249,N_5229);
nor U5326 (N_5326,N_5181,N_5215);
and U5327 (N_5327,N_5238,N_5130);
nand U5328 (N_5328,N_5162,N_5142);
or U5329 (N_5329,N_5267,N_5203);
nand U5330 (N_5330,N_5256,N_5187);
and U5331 (N_5331,N_5132,N_5134);
nand U5332 (N_5332,N_5250,N_5278);
or U5333 (N_5333,N_5192,N_5216);
xor U5334 (N_5334,N_5139,N_5195);
nor U5335 (N_5335,N_5120,N_5168);
nand U5336 (N_5336,N_5153,N_5206);
xnor U5337 (N_5337,N_5197,N_5164);
or U5338 (N_5338,N_5224,N_5129);
nand U5339 (N_5339,N_5136,N_5204);
nand U5340 (N_5340,N_5269,N_5241);
nor U5341 (N_5341,N_5230,N_5137);
xnor U5342 (N_5342,N_5244,N_5266);
xnor U5343 (N_5343,N_5260,N_5124);
and U5344 (N_5344,N_5158,N_5175);
and U5345 (N_5345,N_5191,N_5166);
nor U5346 (N_5346,N_5245,N_5127);
nor U5347 (N_5347,N_5222,N_5227);
nand U5348 (N_5348,N_5210,N_5152);
nand U5349 (N_5349,N_5234,N_5236);
or U5350 (N_5350,N_5259,N_5150);
or U5351 (N_5351,N_5133,N_5184);
and U5352 (N_5352,N_5220,N_5202);
nand U5353 (N_5353,N_5180,N_5225);
or U5354 (N_5354,N_5255,N_5122);
nor U5355 (N_5355,N_5248,N_5257);
and U5356 (N_5356,N_5264,N_5183);
nand U5357 (N_5357,N_5149,N_5157);
and U5358 (N_5358,N_5201,N_5232);
or U5359 (N_5359,N_5146,N_5141);
nor U5360 (N_5360,N_5154,N_5125);
nand U5361 (N_5361,N_5175,N_5156);
nand U5362 (N_5362,N_5205,N_5184);
nand U5363 (N_5363,N_5193,N_5256);
and U5364 (N_5364,N_5255,N_5177);
or U5365 (N_5365,N_5228,N_5264);
nand U5366 (N_5366,N_5229,N_5250);
nor U5367 (N_5367,N_5222,N_5145);
and U5368 (N_5368,N_5212,N_5237);
nor U5369 (N_5369,N_5126,N_5240);
nor U5370 (N_5370,N_5172,N_5186);
xnor U5371 (N_5371,N_5166,N_5123);
and U5372 (N_5372,N_5247,N_5189);
xnor U5373 (N_5373,N_5137,N_5167);
xnor U5374 (N_5374,N_5124,N_5156);
or U5375 (N_5375,N_5249,N_5211);
xnor U5376 (N_5376,N_5190,N_5124);
xor U5377 (N_5377,N_5133,N_5181);
and U5378 (N_5378,N_5170,N_5246);
nand U5379 (N_5379,N_5198,N_5240);
xor U5380 (N_5380,N_5192,N_5239);
or U5381 (N_5381,N_5127,N_5209);
nand U5382 (N_5382,N_5238,N_5260);
nand U5383 (N_5383,N_5131,N_5130);
xor U5384 (N_5384,N_5186,N_5251);
nand U5385 (N_5385,N_5124,N_5141);
or U5386 (N_5386,N_5268,N_5154);
nor U5387 (N_5387,N_5239,N_5218);
or U5388 (N_5388,N_5243,N_5231);
nand U5389 (N_5389,N_5170,N_5176);
nor U5390 (N_5390,N_5141,N_5209);
nand U5391 (N_5391,N_5168,N_5205);
or U5392 (N_5392,N_5148,N_5175);
and U5393 (N_5393,N_5133,N_5256);
or U5394 (N_5394,N_5137,N_5272);
or U5395 (N_5395,N_5190,N_5185);
or U5396 (N_5396,N_5217,N_5206);
xnor U5397 (N_5397,N_5253,N_5241);
and U5398 (N_5398,N_5196,N_5165);
and U5399 (N_5399,N_5124,N_5200);
nand U5400 (N_5400,N_5158,N_5267);
nor U5401 (N_5401,N_5169,N_5241);
nand U5402 (N_5402,N_5142,N_5159);
and U5403 (N_5403,N_5248,N_5261);
or U5404 (N_5404,N_5151,N_5226);
or U5405 (N_5405,N_5191,N_5136);
xnor U5406 (N_5406,N_5256,N_5222);
nand U5407 (N_5407,N_5207,N_5193);
or U5408 (N_5408,N_5207,N_5145);
and U5409 (N_5409,N_5210,N_5178);
nor U5410 (N_5410,N_5178,N_5144);
xor U5411 (N_5411,N_5197,N_5193);
xnor U5412 (N_5412,N_5252,N_5254);
or U5413 (N_5413,N_5216,N_5193);
nor U5414 (N_5414,N_5191,N_5243);
nand U5415 (N_5415,N_5123,N_5178);
or U5416 (N_5416,N_5121,N_5266);
xor U5417 (N_5417,N_5147,N_5254);
nand U5418 (N_5418,N_5122,N_5171);
xor U5419 (N_5419,N_5142,N_5136);
nand U5420 (N_5420,N_5261,N_5184);
nand U5421 (N_5421,N_5263,N_5251);
and U5422 (N_5422,N_5152,N_5183);
or U5423 (N_5423,N_5159,N_5205);
and U5424 (N_5424,N_5190,N_5255);
or U5425 (N_5425,N_5129,N_5263);
nor U5426 (N_5426,N_5255,N_5246);
nand U5427 (N_5427,N_5153,N_5226);
nor U5428 (N_5428,N_5197,N_5175);
and U5429 (N_5429,N_5218,N_5237);
or U5430 (N_5430,N_5278,N_5170);
and U5431 (N_5431,N_5168,N_5196);
and U5432 (N_5432,N_5271,N_5132);
xnor U5433 (N_5433,N_5131,N_5186);
xor U5434 (N_5434,N_5217,N_5199);
nand U5435 (N_5435,N_5269,N_5225);
nand U5436 (N_5436,N_5232,N_5167);
nand U5437 (N_5437,N_5235,N_5196);
nand U5438 (N_5438,N_5248,N_5181);
and U5439 (N_5439,N_5219,N_5126);
xor U5440 (N_5440,N_5395,N_5432);
and U5441 (N_5441,N_5341,N_5426);
nor U5442 (N_5442,N_5321,N_5373);
nand U5443 (N_5443,N_5309,N_5387);
xnor U5444 (N_5444,N_5382,N_5376);
or U5445 (N_5445,N_5351,N_5427);
nand U5446 (N_5446,N_5331,N_5339);
xnor U5447 (N_5447,N_5295,N_5299);
or U5448 (N_5448,N_5413,N_5396);
xor U5449 (N_5449,N_5398,N_5345);
nand U5450 (N_5450,N_5320,N_5438);
and U5451 (N_5451,N_5423,N_5288);
nor U5452 (N_5452,N_5401,N_5359);
or U5453 (N_5453,N_5352,N_5412);
or U5454 (N_5454,N_5439,N_5374);
or U5455 (N_5455,N_5294,N_5364);
xor U5456 (N_5456,N_5346,N_5297);
nor U5457 (N_5457,N_5305,N_5362);
xor U5458 (N_5458,N_5325,N_5327);
nand U5459 (N_5459,N_5317,N_5322);
or U5460 (N_5460,N_5293,N_5306);
xor U5461 (N_5461,N_5409,N_5381);
nor U5462 (N_5462,N_5436,N_5290);
nand U5463 (N_5463,N_5348,N_5433);
nor U5464 (N_5464,N_5425,N_5302);
xor U5465 (N_5465,N_5361,N_5437);
and U5466 (N_5466,N_5282,N_5386);
nor U5467 (N_5467,N_5407,N_5329);
nor U5468 (N_5468,N_5336,N_5343);
nand U5469 (N_5469,N_5404,N_5307);
nor U5470 (N_5470,N_5405,N_5399);
xor U5471 (N_5471,N_5372,N_5408);
or U5472 (N_5472,N_5291,N_5333);
and U5473 (N_5473,N_5323,N_5349);
nand U5474 (N_5474,N_5410,N_5357);
nand U5475 (N_5475,N_5337,N_5281);
or U5476 (N_5476,N_5344,N_5356);
xnor U5477 (N_5477,N_5324,N_5429);
xnor U5478 (N_5478,N_5384,N_5388);
nor U5479 (N_5479,N_5316,N_5390);
or U5480 (N_5480,N_5280,N_5419);
nor U5481 (N_5481,N_5416,N_5363);
and U5482 (N_5482,N_5338,N_5421);
nor U5483 (N_5483,N_5431,N_5313);
nand U5484 (N_5484,N_5355,N_5418);
and U5485 (N_5485,N_5370,N_5296);
and U5486 (N_5486,N_5292,N_5430);
nor U5487 (N_5487,N_5285,N_5286);
and U5488 (N_5488,N_5332,N_5415);
xor U5489 (N_5489,N_5330,N_5365);
nor U5490 (N_5490,N_5434,N_5342);
nor U5491 (N_5491,N_5301,N_5367);
nor U5492 (N_5492,N_5389,N_5368);
nand U5493 (N_5493,N_5334,N_5284);
nand U5494 (N_5494,N_5397,N_5353);
nand U5495 (N_5495,N_5377,N_5300);
and U5496 (N_5496,N_5420,N_5318);
xnor U5497 (N_5497,N_5304,N_5414);
xnor U5498 (N_5498,N_5383,N_5394);
nand U5499 (N_5499,N_5310,N_5375);
xnor U5500 (N_5500,N_5287,N_5392);
or U5501 (N_5501,N_5385,N_5350);
or U5502 (N_5502,N_5380,N_5358);
or U5503 (N_5503,N_5314,N_5366);
nand U5504 (N_5504,N_5347,N_5315);
xor U5505 (N_5505,N_5406,N_5311);
and U5506 (N_5506,N_5435,N_5403);
or U5507 (N_5507,N_5422,N_5283);
nor U5508 (N_5508,N_5411,N_5308);
or U5509 (N_5509,N_5312,N_5417);
xnor U5510 (N_5510,N_5400,N_5360);
and U5511 (N_5511,N_5328,N_5428);
or U5512 (N_5512,N_5371,N_5424);
nor U5513 (N_5513,N_5289,N_5326);
xor U5514 (N_5514,N_5402,N_5319);
or U5515 (N_5515,N_5393,N_5340);
nand U5516 (N_5516,N_5369,N_5379);
and U5517 (N_5517,N_5298,N_5303);
or U5518 (N_5518,N_5335,N_5391);
nor U5519 (N_5519,N_5378,N_5354);
nand U5520 (N_5520,N_5371,N_5425);
xnor U5521 (N_5521,N_5344,N_5411);
nand U5522 (N_5522,N_5434,N_5341);
nor U5523 (N_5523,N_5316,N_5310);
or U5524 (N_5524,N_5406,N_5404);
xnor U5525 (N_5525,N_5299,N_5311);
or U5526 (N_5526,N_5431,N_5294);
and U5527 (N_5527,N_5309,N_5357);
xor U5528 (N_5528,N_5285,N_5297);
nand U5529 (N_5529,N_5416,N_5399);
nor U5530 (N_5530,N_5361,N_5395);
xor U5531 (N_5531,N_5438,N_5395);
nand U5532 (N_5532,N_5351,N_5375);
xnor U5533 (N_5533,N_5353,N_5326);
xor U5534 (N_5534,N_5433,N_5349);
and U5535 (N_5535,N_5416,N_5350);
nor U5536 (N_5536,N_5390,N_5328);
or U5537 (N_5537,N_5384,N_5310);
xor U5538 (N_5538,N_5337,N_5405);
nor U5539 (N_5539,N_5366,N_5436);
xnor U5540 (N_5540,N_5328,N_5304);
or U5541 (N_5541,N_5303,N_5330);
xnor U5542 (N_5542,N_5385,N_5344);
or U5543 (N_5543,N_5369,N_5417);
xnor U5544 (N_5544,N_5411,N_5402);
xor U5545 (N_5545,N_5432,N_5425);
xnor U5546 (N_5546,N_5317,N_5354);
nand U5547 (N_5547,N_5380,N_5381);
or U5548 (N_5548,N_5318,N_5385);
and U5549 (N_5549,N_5327,N_5411);
xor U5550 (N_5550,N_5316,N_5395);
and U5551 (N_5551,N_5306,N_5429);
or U5552 (N_5552,N_5283,N_5282);
and U5553 (N_5553,N_5346,N_5356);
nor U5554 (N_5554,N_5350,N_5312);
and U5555 (N_5555,N_5437,N_5313);
nand U5556 (N_5556,N_5340,N_5287);
nor U5557 (N_5557,N_5342,N_5339);
nand U5558 (N_5558,N_5415,N_5325);
or U5559 (N_5559,N_5332,N_5311);
xnor U5560 (N_5560,N_5334,N_5424);
and U5561 (N_5561,N_5328,N_5376);
nand U5562 (N_5562,N_5423,N_5305);
and U5563 (N_5563,N_5318,N_5316);
nand U5564 (N_5564,N_5391,N_5352);
nand U5565 (N_5565,N_5378,N_5397);
nand U5566 (N_5566,N_5344,N_5287);
nand U5567 (N_5567,N_5430,N_5406);
nand U5568 (N_5568,N_5381,N_5332);
nand U5569 (N_5569,N_5292,N_5357);
or U5570 (N_5570,N_5297,N_5388);
xor U5571 (N_5571,N_5329,N_5321);
or U5572 (N_5572,N_5424,N_5340);
xor U5573 (N_5573,N_5399,N_5313);
nand U5574 (N_5574,N_5323,N_5342);
nand U5575 (N_5575,N_5373,N_5374);
or U5576 (N_5576,N_5380,N_5312);
nor U5577 (N_5577,N_5314,N_5415);
nand U5578 (N_5578,N_5375,N_5392);
xor U5579 (N_5579,N_5335,N_5312);
xor U5580 (N_5580,N_5310,N_5342);
nor U5581 (N_5581,N_5317,N_5409);
or U5582 (N_5582,N_5281,N_5371);
or U5583 (N_5583,N_5315,N_5437);
xnor U5584 (N_5584,N_5285,N_5348);
and U5585 (N_5585,N_5336,N_5340);
and U5586 (N_5586,N_5349,N_5322);
or U5587 (N_5587,N_5319,N_5361);
xnor U5588 (N_5588,N_5294,N_5324);
xnor U5589 (N_5589,N_5382,N_5361);
xor U5590 (N_5590,N_5399,N_5412);
and U5591 (N_5591,N_5313,N_5319);
or U5592 (N_5592,N_5370,N_5306);
nand U5593 (N_5593,N_5312,N_5373);
and U5594 (N_5594,N_5433,N_5374);
or U5595 (N_5595,N_5363,N_5361);
or U5596 (N_5596,N_5330,N_5416);
xnor U5597 (N_5597,N_5307,N_5309);
xor U5598 (N_5598,N_5345,N_5370);
and U5599 (N_5599,N_5434,N_5414);
xnor U5600 (N_5600,N_5494,N_5559);
or U5601 (N_5601,N_5512,N_5567);
and U5602 (N_5602,N_5446,N_5493);
nand U5603 (N_5603,N_5485,N_5482);
xnor U5604 (N_5604,N_5538,N_5531);
and U5605 (N_5605,N_5560,N_5481);
nor U5606 (N_5606,N_5546,N_5581);
xor U5607 (N_5607,N_5444,N_5585);
nand U5608 (N_5608,N_5599,N_5584);
nor U5609 (N_5609,N_5460,N_5596);
nand U5610 (N_5610,N_5586,N_5449);
and U5611 (N_5611,N_5479,N_5452);
nand U5612 (N_5612,N_5540,N_5443);
nor U5613 (N_5613,N_5467,N_5490);
xnor U5614 (N_5614,N_5447,N_5553);
nor U5615 (N_5615,N_5568,N_5530);
nor U5616 (N_5616,N_5549,N_5453);
nand U5617 (N_5617,N_5473,N_5489);
nor U5618 (N_5618,N_5552,N_5517);
nand U5619 (N_5619,N_5442,N_5574);
or U5620 (N_5620,N_5528,N_5470);
and U5621 (N_5621,N_5544,N_5569);
or U5622 (N_5622,N_5510,N_5504);
xnor U5623 (N_5623,N_5562,N_5537);
nor U5624 (N_5624,N_5580,N_5514);
nand U5625 (N_5625,N_5573,N_5595);
nor U5626 (N_5626,N_5505,N_5476);
and U5627 (N_5627,N_5561,N_5448);
xor U5628 (N_5628,N_5457,N_5475);
or U5629 (N_5629,N_5550,N_5486);
xnor U5630 (N_5630,N_5471,N_5511);
or U5631 (N_5631,N_5454,N_5542);
nor U5632 (N_5632,N_5590,N_5513);
nand U5633 (N_5633,N_5507,N_5480);
nand U5634 (N_5634,N_5536,N_5483);
nand U5635 (N_5635,N_5527,N_5594);
and U5636 (N_5636,N_5566,N_5492);
and U5637 (N_5637,N_5455,N_5456);
xnor U5638 (N_5638,N_5466,N_5541);
xor U5639 (N_5639,N_5491,N_5555);
or U5640 (N_5640,N_5548,N_5441);
and U5641 (N_5641,N_5522,N_5521);
nand U5642 (N_5642,N_5589,N_5462);
nor U5643 (N_5643,N_5488,N_5524);
or U5644 (N_5644,N_5529,N_5571);
xnor U5645 (N_5645,N_5583,N_5472);
nand U5646 (N_5646,N_5469,N_5445);
xnor U5647 (N_5647,N_5478,N_5463);
and U5648 (N_5648,N_5558,N_5464);
and U5649 (N_5649,N_5496,N_5565);
xor U5650 (N_5650,N_5556,N_5503);
nor U5651 (N_5651,N_5465,N_5534);
and U5652 (N_5652,N_5579,N_5539);
or U5653 (N_5653,N_5557,N_5500);
and U5654 (N_5654,N_5547,N_5508);
xor U5655 (N_5655,N_5591,N_5575);
xnor U5656 (N_5656,N_5461,N_5487);
nand U5657 (N_5657,N_5577,N_5515);
nand U5658 (N_5658,N_5459,N_5495);
xnor U5659 (N_5659,N_5597,N_5578);
and U5660 (N_5660,N_5576,N_5451);
xnor U5661 (N_5661,N_5532,N_5572);
nor U5662 (N_5662,N_5598,N_5554);
nor U5663 (N_5663,N_5523,N_5502);
or U5664 (N_5664,N_5477,N_5440);
nor U5665 (N_5665,N_5450,N_5592);
and U5666 (N_5666,N_5499,N_5468);
nor U5667 (N_5667,N_5543,N_5533);
nand U5668 (N_5668,N_5474,N_5551);
and U5669 (N_5669,N_5582,N_5526);
or U5670 (N_5670,N_5516,N_5535);
nand U5671 (N_5671,N_5564,N_5588);
and U5672 (N_5672,N_5587,N_5506);
or U5673 (N_5673,N_5497,N_5484);
or U5674 (N_5674,N_5525,N_5570);
and U5675 (N_5675,N_5545,N_5593);
xor U5676 (N_5676,N_5498,N_5520);
xor U5677 (N_5677,N_5518,N_5458);
xor U5678 (N_5678,N_5501,N_5509);
or U5679 (N_5679,N_5519,N_5563);
nor U5680 (N_5680,N_5576,N_5597);
nand U5681 (N_5681,N_5514,N_5596);
xor U5682 (N_5682,N_5486,N_5481);
nand U5683 (N_5683,N_5545,N_5529);
or U5684 (N_5684,N_5454,N_5506);
nor U5685 (N_5685,N_5480,N_5472);
and U5686 (N_5686,N_5503,N_5552);
nand U5687 (N_5687,N_5595,N_5507);
nand U5688 (N_5688,N_5560,N_5532);
and U5689 (N_5689,N_5594,N_5519);
nor U5690 (N_5690,N_5461,N_5445);
nand U5691 (N_5691,N_5506,N_5446);
xor U5692 (N_5692,N_5440,N_5492);
nor U5693 (N_5693,N_5507,N_5567);
nand U5694 (N_5694,N_5581,N_5572);
and U5695 (N_5695,N_5598,N_5517);
nor U5696 (N_5696,N_5472,N_5459);
xnor U5697 (N_5697,N_5449,N_5597);
nand U5698 (N_5698,N_5568,N_5469);
nor U5699 (N_5699,N_5510,N_5518);
xor U5700 (N_5700,N_5533,N_5464);
nor U5701 (N_5701,N_5572,N_5590);
or U5702 (N_5702,N_5451,N_5531);
nand U5703 (N_5703,N_5480,N_5596);
or U5704 (N_5704,N_5583,N_5579);
and U5705 (N_5705,N_5578,N_5454);
or U5706 (N_5706,N_5583,N_5452);
nand U5707 (N_5707,N_5577,N_5481);
nand U5708 (N_5708,N_5598,N_5521);
xor U5709 (N_5709,N_5453,N_5555);
and U5710 (N_5710,N_5528,N_5486);
or U5711 (N_5711,N_5588,N_5512);
or U5712 (N_5712,N_5457,N_5459);
nand U5713 (N_5713,N_5522,N_5584);
xor U5714 (N_5714,N_5546,N_5563);
nor U5715 (N_5715,N_5588,N_5511);
and U5716 (N_5716,N_5546,N_5542);
nor U5717 (N_5717,N_5560,N_5554);
and U5718 (N_5718,N_5499,N_5581);
and U5719 (N_5719,N_5508,N_5581);
or U5720 (N_5720,N_5463,N_5499);
xnor U5721 (N_5721,N_5539,N_5506);
nor U5722 (N_5722,N_5457,N_5542);
nand U5723 (N_5723,N_5555,N_5539);
xor U5724 (N_5724,N_5459,N_5467);
xor U5725 (N_5725,N_5486,N_5500);
nand U5726 (N_5726,N_5501,N_5572);
nor U5727 (N_5727,N_5455,N_5457);
and U5728 (N_5728,N_5510,N_5508);
xnor U5729 (N_5729,N_5465,N_5571);
nor U5730 (N_5730,N_5488,N_5547);
nand U5731 (N_5731,N_5493,N_5445);
nor U5732 (N_5732,N_5561,N_5476);
xnor U5733 (N_5733,N_5579,N_5505);
xnor U5734 (N_5734,N_5472,N_5477);
nand U5735 (N_5735,N_5491,N_5574);
or U5736 (N_5736,N_5461,N_5492);
xor U5737 (N_5737,N_5545,N_5557);
or U5738 (N_5738,N_5563,N_5450);
nand U5739 (N_5739,N_5448,N_5525);
nand U5740 (N_5740,N_5562,N_5532);
and U5741 (N_5741,N_5447,N_5578);
or U5742 (N_5742,N_5521,N_5563);
xnor U5743 (N_5743,N_5548,N_5505);
nor U5744 (N_5744,N_5542,N_5554);
nand U5745 (N_5745,N_5461,N_5448);
nor U5746 (N_5746,N_5506,N_5597);
or U5747 (N_5747,N_5463,N_5457);
nand U5748 (N_5748,N_5488,N_5546);
nor U5749 (N_5749,N_5468,N_5464);
xnor U5750 (N_5750,N_5443,N_5584);
nor U5751 (N_5751,N_5478,N_5508);
nor U5752 (N_5752,N_5586,N_5555);
or U5753 (N_5753,N_5481,N_5499);
nand U5754 (N_5754,N_5527,N_5463);
nor U5755 (N_5755,N_5482,N_5590);
nand U5756 (N_5756,N_5445,N_5540);
xnor U5757 (N_5757,N_5532,N_5479);
or U5758 (N_5758,N_5447,N_5465);
nor U5759 (N_5759,N_5484,N_5546);
xor U5760 (N_5760,N_5620,N_5704);
or U5761 (N_5761,N_5710,N_5701);
xor U5762 (N_5762,N_5652,N_5744);
nand U5763 (N_5763,N_5617,N_5644);
or U5764 (N_5764,N_5612,N_5705);
nand U5765 (N_5765,N_5694,N_5697);
or U5766 (N_5766,N_5624,N_5610);
and U5767 (N_5767,N_5750,N_5604);
and U5768 (N_5768,N_5731,N_5737);
xnor U5769 (N_5769,N_5732,N_5699);
or U5770 (N_5770,N_5692,N_5665);
nor U5771 (N_5771,N_5717,N_5713);
or U5772 (N_5772,N_5660,N_5729);
nand U5773 (N_5773,N_5600,N_5675);
and U5774 (N_5774,N_5645,N_5679);
nand U5775 (N_5775,N_5639,N_5643);
nand U5776 (N_5776,N_5661,N_5629);
nand U5777 (N_5777,N_5642,N_5685);
nor U5778 (N_5778,N_5608,N_5693);
nor U5779 (N_5779,N_5637,N_5700);
nand U5780 (N_5780,N_5736,N_5621);
nand U5781 (N_5781,N_5616,N_5690);
nor U5782 (N_5782,N_5618,N_5681);
or U5783 (N_5783,N_5635,N_5672);
xor U5784 (N_5784,N_5633,N_5686);
and U5785 (N_5785,N_5657,N_5676);
xnor U5786 (N_5786,N_5726,N_5725);
or U5787 (N_5787,N_5655,N_5709);
or U5788 (N_5788,N_5683,N_5647);
nor U5789 (N_5789,N_5626,N_5735);
xnor U5790 (N_5790,N_5748,N_5730);
or U5791 (N_5791,N_5670,N_5752);
nand U5792 (N_5792,N_5611,N_5663);
or U5793 (N_5793,N_5684,N_5739);
and U5794 (N_5794,N_5678,N_5677);
nor U5795 (N_5795,N_5651,N_5747);
nor U5796 (N_5796,N_5720,N_5641);
nand U5797 (N_5797,N_5619,N_5664);
or U5798 (N_5798,N_5671,N_5719);
nand U5799 (N_5799,N_5646,N_5627);
nor U5800 (N_5800,N_5716,N_5602);
and U5801 (N_5801,N_5613,N_5636);
and U5802 (N_5802,N_5696,N_5695);
or U5803 (N_5803,N_5754,N_5656);
nand U5804 (N_5804,N_5625,N_5756);
or U5805 (N_5805,N_5640,N_5740);
nor U5806 (N_5806,N_5638,N_5698);
or U5807 (N_5807,N_5666,N_5674);
or U5808 (N_5808,N_5615,N_5673);
nor U5809 (N_5809,N_5734,N_5614);
or U5810 (N_5810,N_5605,N_5668);
or U5811 (N_5811,N_5711,N_5741);
xnor U5812 (N_5812,N_5733,N_5745);
and U5813 (N_5813,N_5703,N_5723);
nor U5814 (N_5814,N_5749,N_5667);
xnor U5815 (N_5815,N_5758,N_5682);
and U5816 (N_5816,N_5738,N_5722);
nor U5817 (N_5817,N_5728,N_5628);
or U5818 (N_5818,N_5757,N_5632);
or U5819 (N_5819,N_5688,N_5727);
or U5820 (N_5820,N_5707,N_5708);
or U5821 (N_5821,N_5622,N_5631);
nand U5822 (N_5822,N_5746,N_5751);
or U5823 (N_5823,N_5653,N_5654);
xor U5824 (N_5824,N_5650,N_5680);
nand U5825 (N_5825,N_5609,N_5759);
nand U5826 (N_5826,N_5662,N_5715);
and U5827 (N_5827,N_5649,N_5702);
or U5828 (N_5828,N_5607,N_5658);
and U5829 (N_5829,N_5659,N_5648);
nand U5830 (N_5830,N_5691,N_5601);
nor U5831 (N_5831,N_5743,N_5689);
nand U5832 (N_5832,N_5606,N_5634);
and U5833 (N_5833,N_5712,N_5718);
or U5834 (N_5834,N_5742,N_5706);
xor U5835 (N_5835,N_5603,N_5630);
nand U5836 (N_5836,N_5721,N_5687);
or U5837 (N_5837,N_5753,N_5669);
xnor U5838 (N_5838,N_5714,N_5623);
or U5839 (N_5839,N_5755,N_5724);
xnor U5840 (N_5840,N_5759,N_5686);
nand U5841 (N_5841,N_5729,N_5656);
xor U5842 (N_5842,N_5617,N_5698);
or U5843 (N_5843,N_5756,N_5667);
and U5844 (N_5844,N_5703,N_5634);
or U5845 (N_5845,N_5740,N_5728);
nand U5846 (N_5846,N_5631,N_5670);
nor U5847 (N_5847,N_5744,N_5600);
nor U5848 (N_5848,N_5727,N_5720);
nand U5849 (N_5849,N_5624,N_5677);
and U5850 (N_5850,N_5665,N_5614);
or U5851 (N_5851,N_5618,N_5669);
and U5852 (N_5852,N_5721,N_5659);
or U5853 (N_5853,N_5668,N_5611);
and U5854 (N_5854,N_5693,N_5741);
nor U5855 (N_5855,N_5715,N_5702);
or U5856 (N_5856,N_5636,N_5737);
or U5857 (N_5857,N_5667,N_5629);
nor U5858 (N_5858,N_5756,N_5653);
and U5859 (N_5859,N_5625,N_5671);
nor U5860 (N_5860,N_5712,N_5623);
or U5861 (N_5861,N_5634,N_5750);
nand U5862 (N_5862,N_5626,N_5664);
or U5863 (N_5863,N_5742,N_5680);
or U5864 (N_5864,N_5689,N_5729);
nor U5865 (N_5865,N_5655,N_5713);
or U5866 (N_5866,N_5611,N_5636);
xnor U5867 (N_5867,N_5753,N_5759);
nand U5868 (N_5868,N_5727,N_5748);
nor U5869 (N_5869,N_5718,N_5659);
nor U5870 (N_5870,N_5698,N_5702);
nor U5871 (N_5871,N_5708,N_5629);
and U5872 (N_5872,N_5650,N_5695);
and U5873 (N_5873,N_5743,N_5614);
nand U5874 (N_5874,N_5724,N_5632);
xor U5875 (N_5875,N_5601,N_5703);
and U5876 (N_5876,N_5752,N_5676);
nor U5877 (N_5877,N_5649,N_5708);
nor U5878 (N_5878,N_5630,N_5699);
and U5879 (N_5879,N_5753,N_5639);
nor U5880 (N_5880,N_5744,N_5601);
xnor U5881 (N_5881,N_5660,N_5677);
nor U5882 (N_5882,N_5647,N_5686);
nand U5883 (N_5883,N_5709,N_5719);
xnor U5884 (N_5884,N_5653,N_5608);
xor U5885 (N_5885,N_5732,N_5627);
nand U5886 (N_5886,N_5662,N_5680);
nor U5887 (N_5887,N_5708,N_5700);
and U5888 (N_5888,N_5672,N_5734);
or U5889 (N_5889,N_5670,N_5714);
nand U5890 (N_5890,N_5734,N_5661);
nand U5891 (N_5891,N_5656,N_5660);
nor U5892 (N_5892,N_5610,N_5739);
or U5893 (N_5893,N_5721,N_5608);
and U5894 (N_5894,N_5661,N_5644);
nand U5895 (N_5895,N_5638,N_5657);
nor U5896 (N_5896,N_5724,N_5751);
nor U5897 (N_5897,N_5716,N_5689);
nand U5898 (N_5898,N_5701,N_5706);
and U5899 (N_5899,N_5687,N_5632);
or U5900 (N_5900,N_5605,N_5757);
nor U5901 (N_5901,N_5710,N_5637);
or U5902 (N_5902,N_5741,N_5615);
nor U5903 (N_5903,N_5718,N_5685);
nand U5904 (N_5904,N_5673,N_5756);
xor U5905 (N_5905,N_5632,N_5600);
and U5906 (N_5906,N_5666,N_5717);
nor U5907 (N_5907,N_5724,N_5662);
nand U5908 (N_5908,N_5651,N_5707);
xor U5909 (N_5909,N_5614,N_5723);
xnor U5910 (N_5910,N_5659,N_5711);
nand U5911 (N_5911,N_5671,N_5608);
nor U5912 (N_5912,N_5695,N_5745);
or U5913 (N_5913,N_5660,N_5606);
or U5914 (N_5914,N_5717,N_5687);
and U5915 (N_5915,N_5719,N_5629);
nand U5916 (N_5916,N_5696,N_5711);
or U5917 (N_5917,N_5694,N_5638);
nor U5918 (N_5918,N_5625,N_5647);
nor U5919 (N_5919,N_5646,N_5620);
xnor U5920 (N_5920,N_5862,N_5875);
and U5921 (N_5921,N_5852,N_5816);
or U5922 (N_5922,N_5801,N_5840);
nand U5923 (N_5923,N_5910,N_5828);
nand U5924 (N_5924,N_5807,N_5774);
nand U5925 (N_5925,N_5825,N_5768);
nor U5926 (N_5926,N_5834,N_5863);
nand U5927 (N_5927,N_5765,N_5841);
nand U5928 (N_5928,N_5900,N_5796);
nand U5929 (N_5929,N_5790,N_5906);
xnor U5930 (N_5930,N_5783,N_5874);
and U5931 (N_5931,N_5919,N_5847);
or U5932 (N_5932,N_5800,N_5916);
and U5933 (N_5933,N_5907,N_5788);
nor U5934 (N_5934,N_5785,N_5819);
or U5935 (N_5935,N_5802,N_5791);
or U5936 (N_5936,N_5867,N_5818);
or U5937 (N_5937,N_5808,N_5879);
nor U5938 (N_5938,N_5858,N_5870);
nand U5939 (N_5939,N_5918,N_5766);
nand U5940 (N_5940,N_5781,N_5780);
nor U5941 (N_5941,N_5833,N_5821);
xor U5942 (N_5942,N_5865,N_5849);
nand U5943 (N_5943,N_5776,N_5813);
and U5944 (N_5944,N_5851,N_5794);
xor U5945 (N_5945,N_5835,N_5837);
and U5946 (N_5946,N_5886,N_5798);
nor U5947 (N_5947,N_5857,N_5823);
and U5948 (N_5948,N_5839,N_5806);
nor U5949 (N_5949,N_5889,N_5830);
xor U5950 (N_5950,N_5903,N_5860);
or U5951 (N_5951,N_5804,N_5898);
and U5952 (N_5952,N_5799,N_5905);
nand U5953 (N_5953,N_5812,N_5913);
nor U5954 (N_5954,N_5911,N_5760);
nand U5955 (N_5955,N_5909,N_5885);
nor U5956 (N_5956,N_5769,N_5854);
or U5957 (N_5957,N_5787,N_5881);
or U5958 (N_5958,N_5864,N_5843);
nand U5959 (N_5959,N_5868,N_5891);
and U5960 (N_5960,N_5767,N_5883);
nand U5961 (N_5961,N_5772,N_5856);
nor U5962 (N_5962,N_5827,N_5888);
or U5963 (N_5963,N_5895,N_5904);
and U5964 (N_5964,N_5782,N_5887);
xor U5965 (N_5965,N_5764,N_5873);
or U5966 (N_5966,N_5882,N_5773);
and U5967 (N_5967,N_5771,N_5917);
and U5968 (N_5968,N_5853,N_5899);
or U5969 (N_5969,N_5784,N_5877);
or U5970 (N_5970,N_5792,N_5778);
xnor U5971 (N_5971,N_5815,N_5878);
nand U5972 (N_5972,N_5844,N_5829);
nor U5973 (N_5973,N_5859,N_5901);
nand U5974 (N_5974,N_5850,N_5848);
nand U5975 (N_5975,N_5762,N_5914);
xnor U5976 (N_5976,N_5793,N_5822);
or U5977 (N_5977,N_5820,N_5894);
xor U5978 (N_5978,N_5779,N_5795);
nand U5979 (N_5979,N_5805,N_5869);
nand U5980 (N_5980,N_5876,N_5797);
nor U5981 (N_5981,N_5810,N_5880);
or U5982 (N_5982,N_5831,N_5838);
xnor U5983 (N_5983,N_5893,N_5912);
and U5984 (N_5984,N_5884,N_5763);
nor U5985 (N_5985,N_5872,N_5842);
nor U5986 (N_5986,N_5786,N_5908);
and U5987 (N_5987,N_5892,N_5896);
and U5988 (N_5988,N_5789,N_5824);
and U5989 (N_5989,N_5761,N_5855);
nand U5990 (N_5990,N_5890,N_5777);
xor U5991 (N_5991,N_5826,N_5770);
or U5992 (N_5992,N_5871,N_5814);
nor U5993 (N_5993,N_5845,N_5803);
and U5994 (N_5994,N_5915,N_5866);
nand U5995 (N_5995,N_5775,N_5811);
xnor U5996 (N_5996,N_5861,N_5846);
and U5997 (N_5997,N_5817,N_5897);
xor U5998 (N_5998,N_5809,N_5836);
or U5999 (N_5999,N_5902,N_5832);
and U6000 (N_6000,N_5786,N_5819);
and U6001 (N_6001,N_5912,N_5775);
xnor U6002 (N_6002,N_5805,N_5873);
or U6003 (N_6003,N_5762,N_5792);
and U6004 (N_6004,N_5859,N_5789);
nand U6005 (N_6005,N_5900,N_5912);
and U6006 (N_6006,N_5832,N_5888);
or U6007 (N_6007,N_5830,N_5846);
or U6008 (N_6008,N_5764,N_5841);
and U6009 (N_6009,N_5820,N_5842);
nor U6010 (N_6010,N_5889,N_5907);
or U6011 (N_6011,N_5897,N_5834);
nor U6012 (N_6012,N_5826,N_5842);
and U6013 (N_6013,N_5898,N_5846);
nand U6014 (N_6014,N_5835,N_5906);
xnor U6015 (N_6015,N_5882,N_5803);
or U6016 (N_6016,N_5905,N_5834);
or U6017 (N_6017,N_5766,N_5789);
nor U6018 (N_6018,N_5793,N_5878);
nand U6019 (N_6019,N_5770,N_5885);
nand U6020 (N_6020,N_5805,N_5902);
xnor U6021 (N_6021,N_5805,N_5858);
xor U6022 (N_6022,N_5821,N_5765);
nand U6023 (N_6023,N_5878,N_5900);
xnor U6024 (N_6024,N_5760,N_5850);
and U6025 (N_6025,N_5857,N_5892);
xor U6026 (N_6026,N_5907,N_5770);
and U6027 (N_6027,N_5864,N_5868);
xor U6028 (N_6028,N_5855,N_5816);
nor U6029 (N_6029,N_5904,N_5877);
nand U6030 (N_6030,N_5902,N_5873);
or U6031 (N_6031,N_5836,N_5878);
nand U6032 (N_6032,N_5761,N_5817);
nor U6033 (N_6033,N_5761,N_5852);
nand U6034 (N_6034,N_5859,N_5762);
nand U6035 (N_6035,N_5830,N_5810);
nand U6036 (N_6036,N_5826,N_5794);
or U6037 (N_6037,N_5807,N_5884);
or U6038 (N_6038,N_5873,N_5867);
nor U6039 (N_6039,N_5810,N_5771);
or U6040 (N_6040,N_5773,N_5823);
nor U6041 (N_6041,N_5855,N_5910);
nand U6042 (N_6042,N_5884,N_5864);
and U6043 (N_6043,N_5788,N_5867);
and U6044 (N_6044,N_5882,N_5909);
xnor U6045 (N_6045,N_5908,N_5917);
and U6046 (N_6046,N_5871,N_5791);
xnor U6047 (N_6047,N_5854,N_5908);
and U6048 (N_6048,N_5862,N_5823);
nor U6049 (N_6049,N_5880,N_5919);
nand U6050 (N_6050,N_5770,N_5801);
xor U6051 (N_6051,N_5862,N_5883);
or U6052 (N_6052,N_5855,N_5860);
or U6053 (N_6053,N_5782,N_5767);
nand U6054 (N_6054,N_5769,N_5805);
and U6055 (N_6055,N_5805,N_5859);
nor U6056 (N_6056,N_5807,N_5782);
nor U6057 (N_6057,N_5895,N_5859);
nor U6058 (N_6058,N_5845,N_5854);
and U6059 (N_6059,N_5832,N_5841);
or U6060 (N_6060,N_5892,N_5887);
and U6061 (N_6061,N_5773,N_5816);
or U6062 (N_6062,N_5775,N_5852);
nor U6063 (N_6063,N_5859,N_5770);
and U6064 (N_6064,N_5846,N_5777);
nor U6065 (N_6065,N_5821,N_5842);
and U6066 (N_6066,N_5763,N_5807);
nand U6067 (N_6067,N_5833,N_5857);
nor U6068 (N_6068,N_5798,N_5896);
nand U6069 (N_6069,N_5828,N_5885);
or U6070 (N_6070,N_5810,N_5809);
nand U6071 (N_6071,N_5803,N_5848);
or U6072 (N_6072,N_5907,N_5851);
xnor U6073 (N_6073,N_5913,N_5916);
nand U6074 (N_6074,N_5778,N_5834);
or U6075 (N_6075,N_5836,N_5867);
xor U6076 (N_6076,N_5893,N_5823);
and U6077 (N_6077,N_5789,N_5876);
xor U6078 (N_6078,N_5790,N_5890);
nand U6079 (N_6079,N_5854,N_5852);
nor U6080 (N_6080,N_5974,N_5998);
and U6081 (N_6081,N_5962,N_6004);
nand U6082 (N_6082,N_5956,N_5921);
or U6083 (N_6083,N_6024,N_5990);
xor U6084 (N_6084,N_6007,N_5950);
nand U6085 (N_6085,N_6069,N_6011);
xnor U6086 (N_6086,N_5922,N_5984);
and U6087 (N_6087,N_6067,N_5959);
nor U6088 (N_6088,N_6030,N_5960);
nand U6089 (N_6089,N_6040,N_5971);
nand U6090 (N_6090,N_6012,N_6073);
or U6091 (N_6091,N_6025,N_5924);
xnor U6092 (N_6092,N_5938,N_5980);
nor U6093 (N_6093,N_5951,N_6066);
nand U6094 (N_6094,N_5929,N_6054);
nand U6095 (N_6095,N_6039,N_6049);
and U6096 (N_6096,N_5995,N_6014);
nand U6097 (N_6097,N_6060,N_5994);
nand U6098 (N_6098,N_6070,N_5927);
nand U6099 (N_6099,N_6061,N_5997);
nand U6100 (N_6100,N_6074,N_6010);
nor U6101 (N_6101,N_5957,N_6063);
or U6102 (N_6102,N_6037,N_6003);
or U6103 (N_6103,N_5958,N_6051);
or U6104 (N_6104,N_5977,N_5996);
or U6105 (N_6105,N_6034,N_5967);
xnor U6106 (N_6106,N_5948,N_6057);
or U6107 (N_6107,N_6026,N_6045);
or U6108 (N_6108,N_5949,N_5985);
xor U6109 (N_6109,N_6016,N_6027);
xor U6110 (N_6110,N_5981,N_5932);
xnor U6111 (N_6111,N_6006,N_6005);
or U6112 (N_6112,N_5968,N_5972);
or U6113 (N_6113,N_6013,N_5931);
nor U6114 (N_6114,N_5930,N_5934);
nand U6115 (N_6115,N_6023,N_5925);
or U6116 (N_6116,N_6009,N_5976);
nor U6117 (N_6117,N_5953,N_6062);
or U6118 (N_6118,N_6031,N_5952);
xnor U6119 (N_6119,N_6015,N_5975);
nand U6120 (N_6120,N_6002,N_5923);
xnor U6121 (N_6121,N_5983,N_6068);
or U6122 (N_6122,N_5966,N_6017);
or U6123 (N_6123,N_6021,N_5947);
nand U6124 (N_6124,N_6071,N_5939);
nand U6125 (N_6125,N_6036,N_6075);
and U6126 (N_6126,N_5978,N_6048);
nor U6127 (N_6127,N_6050,N_6079);
nor U6128 (N_6128,N_5946,N_6022);
and U6129 (N_6129,N_5945,N_6020);
or U6130 (N_6130,N_5954,N_6059);
or U6131 (N_6131,N_5935,N_6028);
and U6132 (N_6132,N_6000,N_6038);
nor U6133 (N_6133,N_5989,N_6047);
nor U6134 (N_6134,N_6029,N_6042);
nand U6135 (N_6135,N_6035,N_5993);
nor U6136 (N_6136,N_5926,N_5999);
or U6137 (N_6137,N_5965,N_6008);
xnor U6138 (N_6138,N_6033,N_5942);
nand U6139 (N_6139,N_6052,N_6041);
xnor U6140 (N_6140,N_5955,N_6032);
nand U6141 (N_6141,N_5944,N_5964);
xnor U6142 (N_6142,N_6046,N_5963);
nand U6143 (N_6143,N_5988,N_6064);
nor U6144 (N_6144,N_5920,N_5961);
nand U6145 (N_6145,N_5937,N_5986);
nand U6146 (N_6146,N_6001,N_6018);
nor U6147 (N_6147,N_5992,N_5973);
nand U6148 (N_6148,N_5928,N_6072);
or U6149 (N_6149,N_6065,N_5982);
nand U6150 (N_6150,N_5936,N_5987);
nor U6151 (N_6151,N_5969,N_6019);
nand U6152 (N_6152,N_5940,N_6044);
and U6153 (N_6153,N_5991,N_6077);
nand U6154 (N_6154,N_6056,N_6053);
nor U6155 (N_6155,N_5941,N_5943);
xor U6156 (N_6156,N_6076,N_5970);
xnor U6157 (N_6157,N_6078,N_6043);
and U6158 (N_6158,N_5933,N_6058);
or U6159 (N_6159,N_6055,N_5979);
and U6160 (N_6160,N_5971,N_6033);
nand U6161 (N_6161,N_6009,N_6074);
or U6162 (N_6162,N_5923,N_5964);
nor U6163 (N_6163,N_5982,N_6037);
nand U6164 (N_6164,N_6012,N_6074);
and U6165 (N_6165,N_6076,N_6056);
or U6166 (N_6166,N_6042,N_5934);
nor U6167 (N_6167,N_5981,N_6030);
xor U6168 (N_6168,N_6028,N_6059);
nand U6169 (N_6169,N_5982,N_5986);
nand U6170 (N_6170,N_6068,N_6044);
or U6171 (N_6171,N_6062,N_5955);
and U6172 (N_6172,N_5941,N_5961);
xor U6173 (N_6173,N_6065,N_6047);
nor U6174 (N_6174,N_6003,N_5988);
nor U6175 (N_6175,N_6019,N_6068);
nor U6176 (N_6176,N_5975,N_6077);
nand U6177 (N_6177,N_5927,N_5984);
and U6178 (N_6178,N_5925,N_5995);
nor U6179 (N_6179,N_5928,N_6046);
nor U6180 (N_6180,N_5967,N_5921);
or U6181 (N_6181,N_5988,N_5960);
nand U6182 (N_6182,N_5930,N_6059);
and U6183 (N_6183,N_5941,N_6036);
xnor U6184 (N_6184,N_5953,N_6014);
or U6185 (N_6185,N_6079,N_6064);
and U6186 (N_6186,N_5973,N_6025);
nor U6187 (N_6187,N_6063,N_5967);
xor U6188 (N_6188,N_6041,N_6056);
or U6189 (N_6189,N_5978,N_6037);
nor U6190 (N_6190,N_6027,N_6062);
nor U6191 (N_6191,N_6053,N_6044);
and U6192 (N_6192,N_6066,N_6008);
and U6193 (N_6193,N_6049,N_5984);
nor U6194 (N_6194,N_6011,N_6001);
xor U6195 (N_6195,N_5962,N_5971);
or U6196 (N_6196,N_5950,N_5983);
xnor U6197 (N_6197,N_5959,N_5982);
xor U6198 (N_6198,N_6033,N_5985);
xnor U6199 (N_6199,N_5999,N_6012);
nand U6200 (N_6200,N_6032,N_5979);
or U6201 (N_6201,N_6073,N_5921);
or U6202 (N_6202,N_6046,N_6026);
nor U6203 (N_6203,N_6073,N_5974);
or U6204 (N_6204,N_5934,N_6078);
or U6205 (N_6205,N_5936,N_5958);
nand U6206 (N_6206,N_5940,N_6000);
or U6207 (N_6207,N_5946,N_6002);
and U6208 (N_6208,N_5954,N_5952);
nand U6209 (N_6209,N_5949,N_6001);
or U6210 (N_6210,N_5980,N_6046);
and U6211 (N_6211,N_6018,N_6021);
or U6212 (N_6212,N_6014,N_5984);
or U6213 (N_6213,N_5953,N_6068);
nor U6214 (N_6214,N_5973,N_5938);
xor U6215 (N_6215,N_5966,N_6012);
and U6216 (N_6216,N_6006,N_5981);
nor U6217 (N_6217,N_5931,N_6051);
or U6218 (N_6218,N_5942,N_5944);
or U6219 (N_6219,N_5951,N_6020);
or U6220 (N_6220,N_5972,N_5946);
nand U6221 (N_6221,N_6076,N_5979);
and U6222 (N_6222,N_5973,N_6048);
or U6223 (N_6223,N_5961,N_5951);
and U6224 (N_6224,N_6026,N_6040);
xor U6225 (N_6225,N_5995,N_6071);
nand U6226 (N_6226,N_6001,N_6021);
or U6227 (N_6227,N_6053,N_5955);
or U6228 (N_6228,N_5937,N_6034);
nor U6229 (N_6229,N_6024,N_6074);
nand U6230 (N_6230,N_6068,N_5970);
xor U6231 (N_6231,N_6049,N_6046);
or U6232 (N_6232,N_6053,N_6047);
xor U6233 (N_6233,N_5960,N_5926);
nand U6234 (N_6234,N_6050,N_6073);
nor U6235 (N_6235,N_6048,N_5964);
and U6236 (N_6236,N_6045,N_5940);
nor U6237 (N_6237,N_5961,N_6039);
nor U6238 (N_6238,N_6014,N_6013);
xor U6239 (N_6239,N_5938,N_6007);
or U6240 (N_6240,N_6141,N_6229);
xor U6241 (N_6241,N_6101,N_6150);
and U6242 (N_6242,N_6225,N_6140);
or U6243 (N_6243,N_6085,N_6171);
and U6244 (N_6244,N_6181,N_6220);
xor U6245 (N_6245,N_6131,N_6134);
and U6246 (N_6246,N_6228,N_6168);
or U6247 (N_6247,N_6207,N_6180);
xor U6248 (N_6248,N_6139,N_6158);
nand U6249 (N_6249,N_6217,N_6223);
nor U6250 (N_6250,N_6184,N_6126);
and U6251 (N_6251,N_6209,N_6200);
xnor U6252 (N_6252,N_6179,N_6084);
or U6253 (N_6253,N_6176,N_6191);
or U6254 (N_6254,N_6195,N_6110);
nand U6255 (N_6255,N_6104,N_6095);
nand U6256 (N_6256,N_6128,N_6203);
and U6257 (N_6257,N_6182,N_6196);
xnor U6258 (N_6258,N_6144,N_6118);
nor U6259 (N_6259,N_6113,N_6163);
nand U6260 (N_6260,N_6233,N_6100);
nor U6261 (N_6261,N_6216,N_6197);
nor U6262 (N_6262,N_6164,N_6167);
and U6263 (N_6263,N_6129,N_6230);
nand U6264 (N_6264,N_6156,N_6108);
or U6265 (N_6265,N_6124,N_6114);
nor U6266 (N_6266,N_6119,N_6091);
or U6267 (N_6267,N_6115,N_6210);
nor U6268 (N_6268,N_6090,N_6080);
or U6269 (N_6269,N_6143,N_6178);
nor U6270 (N_6270,N_6147,N_6165);
xor U6271 (N_6271,N_6125,N_6121);
nor U6272 (N_6272,N_6183,N_6112);
nand U6273 (N_6273,N_6224,N_6227);
xnor U6274 (N_6274,N_6219,N_6117);
and U6275 (N_6275,N_6087,N_6206);
nand U6276 (N_6276,N_6116,N_6086);
nand U6277 (N_6277,N_6106,N_6082);
nor U6278 (N_6278,N_6161,N_6093);
xor U6279 (N_6279,N_6089,N_6149);
nand U6280 (N_6280,N_6205,N_6226);
or U6281 (N_6281,N_6187,N_6154);
and U6282 (N_6282,N_6218,N_6155);
nor U6283 (N_6283,N_6169,N_6120);
xor U6284 (N_6284,N_6103,N_6092);
xor U6285 (N_6285,N_6174,N_6185);
xor U6286 (N_6286,N_6214,N_6152);
and U6287 (N_6287,N_6109,N_6202);
nand U6288 (N_6288,N_6098,N_6221);
xnor U6289 (N_6289,N_6142,N_6212);
or U6290 (N_6290,N_6083,N_6081);
nand U6291 (N_6291,N_6138,N_6135);
nand U6292 (N_6292,N_6193,N_6105);
and U6293 (N_6293,N_6127,N_6190);
and U6294 (N_6294,N_6173,N_6204);
xor U6295 (N_6295,N_6136,N_6222);
and U6296 (N_6296,N_6215,N_6213);
nor U6297 (N_6297,N_6122,N_6111);
or U6298 (N_6298,N_6236,N_6102);
xnor U6299 (N_6299,N_6198,N_6189);
xor U6300 (N_6300,N_6130,N_6172);
or U6301 (N_6301,N_6153,N_6235);
nor U6302 (N_6302,N_6160,N_6162);
and U6303 (N_6303,N_6170,N_6133);
xnor U6304 (N_6304,N_6192,N_6199);
and U6305 (N_6305,N_6132,N_6099);
and U6306 (N_6306,N_6177,N_6094);
xor U6307 (N_6307,N_6201,N_6232);
or U6308 (N_6308,N_6175,N_6237);
or U6309 (N_6309,N_6146,N_6188);
and U6310 (N_6310,N_6159,N_6208);
or U6311 (N_6311,N_6123,N_6186);
nand U6312 (N_6312,N_6107,N_6194);
xor U6313 (N_6313,N_6231,N_6088);
or U6314 (N_6314,N_6239,N_6137);
xor U6315 (N_6315,N_6151,N_6145);
or U6316 (N_6316,N_6148,N_6234);
nand U6317 (N_6317,N_6166,N_6211);
xnor U6318 (N_6318,N_6096,N_6097);
or U6319 (N_6319,N_6238,N_6157);
nor U6320 (N_6320,N_6155,N_6150);
xor U6321 (N_6321,N_6127,N_6097);
xor U6322 (N_6322,N_6188,N_6120);
or U6323 (N_6323,N_6136,N_6133);
nand U6324 (N_6324,N_6136,N_6169);
xor U6325 (N_6325,N_6232,N_6181);
and U6326 (N_6326,N_6201,N_6156);
or U6327 (N_6327,N_6153,N_6133);
and U6328 (N_6328,N_6197,N_6164);
and U6329 (N_6329,N_6159,N_6211);
nor U6330 (N_6330,N_6160,N_6081);
xor U6331 (N_6331,N_6208,N_6118);
nand U6332 (N_6332,N_6160,N_6166);
nand U6333 (N_6333,N_6141,N_6225);
nand U6334 (N_6334,N_6204,N_6124);
xor U6335 (N_6335,N_6088,N_6155);
xor U6336 (N_6336,N_6099,N_6157);
or U6337 (N_6337,N_6224,N_6203);
and U6338 (N_6338,N_6133,N_6206);
nor U6339 (N_6339,N_6135,N_6123);
or U6340 (N_6340,N_6144,N_6237);
xnor U6341 (N_6341,N_6239,N_6133);
nor U6342 (N_6342,N_6153,N_6111);
nand U6343 (N_6343,N_6156,N_6163);
xnor U6344 (N_6344,N_6143,N_6161);
and U6345 (N_6345,N_6153,N_6114);
xor U6346 (N_6346,N_6134,N_6209);
or U6347 (N_6347,N_6188,N_6142);
or U6348 (N_6348,N_6214,N_6210);
nand U6349 (N_6349,N_6170,N_6171);
or U6350 (N_6350,N_6111,N_6181);
and U6351 (N_6351,N_6139,N_6196);
nor U6352 (N_6352,N_6207,N_6214);
or U6353 (N_6353,N_6110,N_6182);
nand U6354 (N_6354,N_6146,N_6170);
or U6355 (N_6355,N_6208,N_6199);
nor U6356 (N_6356,N_6091,N_6152);
or U6357 (N_6357,N_6120,N_6143);
nor U6358 (N_6358,N_6180,N_6219);
nand U6359 (N_6359,N_6229,N_6158);
xnor U6360 (N_6360,N_6199,N_6180);
and U6361 (N_6361,N_6083,N_6162);
or U6362 (N_6362,N_6114,N_6202);
and U6363 (N_6363,N_6178,N_6235);
or U6364 (N_6364,N_6191,N_6080);
and U6365 (N_6365,N_6209,N_6123);
nor U6366 (N_6366,N_6142,N_6183);
or U6367 (N_6367,N_6147,N_6101);
xor U6368 (N_6368,N_6151,N_6165);
or U6369 (N_6369,N_6119,N_6155);
or U6370 (N_6370,N_6215,N_6227);
nor U6371 (N_6371,N_6120,N_6108);
nor U6372 (N_6372,N_6194,N_6222);
or U6373 (N_6373,N_6188,N_6144);
xnor U6374 (N_6374,N_6226,N_6124);
nand U6375 (N_6375,N_6191,N_6091);
nor U6376 (N_6376,N_6143,N_6233);
and U6377 (N_6377,N_6174,N_6167);
nand U6378 (N_6378,N_6209,N_6118);
or U6379 (N_6379,N_6184,N_6206);
nor U6380 (N_6380,N_6233,N_6191);
xnor U6381 (N_6381,N_6145,N_6212);
nand U6382 (N_6382,N_6149,N_6222);
xor U6383 (N_6383,N_6215,N_6120);
or U6384 (N_6384,N_6201,N_6110);
xor U6385 (N_6385,N_6082,N_6096);
xnor U6386 (N_6386,N_6158,N_6108);
or U6387 (N_6387,N_6105,N_6210);
nor U6388 (N_6388,N_6171,N_6182);
or U6389 (N_6389,N_6238,N_6132);
xnor U6390 (N_6390,N_6128,N_6206);
nor U6391 (N_6391,N_6203,N_6137);
or U6392 (N_6392,N_6126,N_6200);
nand U6393 (N_6393,N_6135,N_6176);
nor U6394 (N_6394,N_6183,N_6159);
and U6395 (N_6395,N_6186,N_6135);
or U6396 (N_6396,N_6185,N_6109);
xor U6397 (N_6397,N_6194,N_6167);
xnor U6398 (N_6398,N_6113,N_6114);
nor U6399 (N_6399,N_6179,N_6122);
nand U6400 (N_6400,N_6347,N_6296);
nor U6401 (N_6401,N_6244,N_6270);
or U6402 (N_6402,N_6254,N_6286);
nand U6403 (N_6403,N_6341,N_6325);
nor U6404 (N_6404,N_6354,N_6276);
and U6405 (N_6405,N_6336,N_6307);
nor U6406 (N_6406,N_6317,N_6299);
xnor U6407 (N_6407,N_6258,N_6368);
nor U6408 (N_6408,N_6346,N_6326);
nand U6409 (N_6409,N_6337,N_6288);
nand U6410 (N_6410,N_6315,N_6331);
and U6411 (N_6411,N_6324,N_6261);
xnor U6412 (N_6412,N_6320,N_6396);
nand U6413 (N_6413,N_6333,N_6362);
xor U6414 (N_6414,N_6295,N_6260);
and U6415 (N_6415,N_6314,N_6287);
nor U6416 (N_6416,N_6308,N_6273);
or U6417 (N_6417,N_6392,N_6340);
nand U6418 (N_6418,N_6247,N_6257);
nand U6419 (N_6419,N_6343,N_6387);
nor U6420 (N_6420,N_6266,N_6309);
and U6421 (N_6421,N_6366,N_6361);
and U6422 (N_6422,N_6353,N_6311);
or U6423 (N_6423,N_6253,N_6291);
nor U6424 (N_6424,N_6375,N_6256);
xnor U6425 (N_6425,N_6269,N_6395);
nor U6426 (N_6426,N_6355,N_6328);
nand U6427 (N_6427,N_6268,N_6312);
xor U6428 (N_6428,N_6391,N_6240);
xor U6429 (N_6429,N_6359,N_6356);
and U6430 (N_6430,N_6252,N_6304);
and U6431 (N_6431,N_6388,N_6245);
nor U6432 (N_6432,N_6390,N_6372);
nand U6433 (N_6433,N_6381,N_6250);
nand U6434 (N_6434,N_6259,N_6351);
nand U6435 (N_6435,N_6301,N_6345);
nor U6436 (N_6436,N_6383,N_6321);
nand U6437 (N_6437,N_6335,N_6318);
or U6438 (N_6438,N_6322,N_6279);
nand U6439 (N_6439,N_6248,N_6349);
or U6440 (N_6440,N_6389,N_6364);
nand U6441 (N_6441,N_6365,N_6305);
nor U6442 (N_6442,N_6399,N_6243);
and U6443 (N_6443,N_6274,N_6313);
xor U6444 (N_6444,N_6344,N_6264);
or U6445 (N_6445,N_6246,N_6371);
nand U6446 (N_6446,N_6369,N_6262);
nand U6447 (N_6447,N_6306,N_6384);
or U6448 (N_6448,N_6310,N_6398);
nor U6449 (N_6449,N_6293,N_6339);
xnor U6450 (N_6450,N_6377,N_6378);
nor U6451 (N_6451,N_6373,N_6316);
xnor U6452 (N_6452,N_6255,N_6298);
or U6453 (N_6453,N_6358,N_6397);
nand U6454 (N_6454,N_6319,N_6360);
or U6455 (N_6455,N_6342,N_6267);
or U6456 (N_6456,N_6278,N_6242);
and U6457 (N_6457,N_6334,N_6282);
nand U6458 (N_6458,N_6329,N_6393);
and U6459 (N_6459,N_6327,N_6376);
and U6460 (N_6460,N_6241,N_6303);
nand U6461 (N_6461,N_6263,N_6272);
xnor U6462 (N_6462,N_6350,N_6265);
xnor U6463 (N_6463,N_6363,N_6374);
xor U6464 (N_6464,N_6297,N_6271);
nor U6465 (N_6465,N_6284,N_6394);
and U6466 (N_6466,N_6249,N_6332);
and U6467 (N_6467,N_6281,N_6251);
and U6468 (N_6468,N_6289,N_6348);
nand U6469 (N_6469,N_6338,N_6292);
or U6470 (N_6470,N_6386,N_6323);
nand U6471 (N_6471,N_6357,N_6285);
and U6472 (N_6472,N_6277,N_6370);
xnor U6473 (N_6473,N_6380,N_6283);
nor U6474 (N_6474,N_6352,N_6330);
nand U6475 (N_6475,N_6302,N_6280);
nand U6476 (N_6476,N_6275,N_6382);
and U6477 (N_6477,N_6294,N_6379);
nor U6478 (N_6478,N_6300,N_6367);
nand U6479 (N_6479,N_6290,N_6385);
nor U6480 (N_6480,N_6308,N_6266);
or U6481 (N_6481,N_6320,N_6327);
and U6482 (N_6482,N_6248,N_6345);
nor U6483 (N_6483,N_6272,N_6275);
xnor U6484 (N_6484,N_6361,N_6390);
and U6485 (N_6485,N_6351,N_6306);
nor U6486 (N_6486,N_6369,N_6340);
nand U6487 (N_6487,N_6243,N_6267);
and U6488 (N_6488,N_6284,N_6371);
xor U6489 (N_6489,N_6314,N_6364);
and U6490 (N_6490,N_6349,N_6393);
or U6491 (N_6491,N_6378,N_6392);
nor U6492 (N_6492,N_6323,N_6350);
or U6493 (N_6493,N_6314,N_6293);
nor U6494 (N_6494,N_6385,N_6252);
xor U6495 (N_6495,N_6315,N_6258);
nand U6496 (N_6496,N_6267,N_6380);
xnor U6497 (N_6497,N_6306,N_6338);
nand U6498 (N_6498,N_6321,N_6396);
nand U6499 (N_6499,N_6369,N_6258);
or U6500 (N_6500,N_6337,N_6365);
and U6501 (N_6501,N_6272,N_6367);
and U6502 (N_6502,N_6264,N_6357);
nor U6503 (N_6503,N_6374,N_6330);
and U6504 (N_6504,N_6354,N_6271);
xnor U6505 (N_6505,N_6326,N_6319);
xor U6506 (N_6506,N_6297,N_6390);
nand U6507 (N_6507,N_6328,N_6277);
or U6508 (N_6508,N_6379,N_6240);
nor U6509 (N_6509,N_6311,N_6276);
nor U6510 (N_6510,N_6377,N_6254);
nand U6511 (N_6511,N_6278,N_6318);
xor U6512 (N_6512,N_6380,N_6372);
xnor U6513 (N_6513,N_6297,N_6340);
nor U6514 (N_6514,N_6356,N_6254);
nand U6515 (N_6515,N_6316,N_6244);
and U6516 (N_6516,N_6336,N_6311);
nor U6517 (N_6517,N_6350,N_6250);
xor U6518 (N_6518,N_6304,N_6359);
and U6519 (N_6519,N_6352,N_6341);
or U6520 (N_6520,N_6345,N_6284);
and U6521 (N_6521,N_6384,N_6369);
nand U6522 (N_6522,N_6296,N_6380);
nor U6523 (N_6523,N_6340,N_6338);
nor U6524 (N_6524,N_6314,N_6296);
or U6525 (N_6525,N_6252,N_6311);
or U6526 (N_6526,N_6292,N_6362);
or U6527 (N_6527,N_6335,N_6278);
and U6528 (N_6528,N_6283,N_6243);
nor U6529 (N_6529,N_6360,N_6395);
and U6530 (N_6530,N_6281,N_6341);
and U6531 (N_6531,N_6299,N_6249);
and U6532 (N_6532,N_6256,N_6329);
and U6533 (N_6533,N_6266,N_6348);
or U6534 (N_6534,N_6247,N_6302);
and U6535 (N_6535,N_6382,N_6295);
or U6536 (N_6536,N_6300,N_6359);
or U6537 (N_6537,N_6343,N_6353);
or U6538 (N_6538,N_6351,N_6398);
xor U6539 (N_6539,N_6253,N_6390);
nor U6540 (N_6540,N_6351,N_6243);
and U6541 (N_6541,N_6323,N_6302);
or U6542 (N_6542,N_6317,N_6264);
xor U6543 (N_6543,N_6296,N_6307);
xor U6544 (N_6544,N_6383,N_6398);
xor U6545 (N_6545,N_6275,N_6248);
nand U6546 (N_6546,N_6348,N_6304);
nor U6547 (N_6547,N_6304,N_6336);
or U6548 (N_6548,N_6261,N_6249);
or U6549 (N_6549,N_6277,N_6292);
or U6550 (N_6550,N_6322,N_6328);
nand U6551 (N_6551,N_6287,N_6297);
or U6552 (N_6552,N_6378,N_6330);
and U6553 (N_6553,N_6347,N_6396);
and U6554 (N_6554,N_6264,N_6289);
xnor U6555 (N_6555,N_6371,N_6336);
and U6556 (N_6556,N_6366,N_6339);
nor U6557 (N_6557,N_6277,N_6335);
nand U6558 (N_6558,N_6249,N_6369);
nor U6559 (N_6559,N_6246,N_6256);
or U6560 (N_6560,N_6413,N_6494);
nor U6561 (N_6561,N_6498,N_6453);
and U6562 (N_6562,N_6501,N_6465);
xor U6563 (N_6563,N_6410,N_6428);
nand U6564 (N_6564,N_6401,N_6499);
xor U6565 (N_6565,N_6478,N_6531);
nor U6566 (N_6566,N_6526,N_6475);
and U6567 (N_6567,N_6437,N_6402);
or U6568 (N_6568,N_6549,N_6540);
and U6569 (N_6569,N_6552,N_6408);
xnor U6570 (N_6570,N_6455,N_6488);
nor U6571 (N_6571,N_6415,N_6514);
nand U6572 (N_6572,N_6405,N_6556);
nor U6573 (N_6573,N_6462,N_6440);
nand U6574 (N_6574,N_6544,N_6481);
and U6575 (N_6575,N_6536,N_6541);
or U6576 (N_6576,N_6513,N_6418);
and U6577 (N_6577,N_6557,N_6445);
and U6578 (N_6578,N_6473,N_6400);
nand U6579 (N_6579,N_6442,N_6438);
and U6580 (N_6580,N_6502,N_6407);
nor U6581 (N_6581,N_6450,N_6510);
nor U6582 (N_6582,N_6483,N_6467);
xnor U6583 (N_6583,N_6530,N_6482);
or U6584 (N_6584,N_6468,N_6419);
and U6585 (N_6585,N_6446,N_6421);
nand U6586 (N_6586,N_6411,N_6529);
or U6587 (N_6587,N_6550,N_6451);
xor U6588 (N_6588,N_6527,N_6495);
and U6589 (N_6589,N_6409,N_6534);
and U6590 (N_6590,N_6430,N_6535);
nor U6591 (N_6591,N_6471,N_6470);
xor U6592 (N_6592,N_6447,N_6558);
nor U6593 (N_6593,N_6448,N_6537);
xor U6594 (N_6594,N_6511,N_6479);
and U6595 (N_6595,N_6507,N_6457);
or U6596 (N_6596,N_6476,N_6449);
and U6597 (N_6597,N_6554,N_6420);
and U6598 (N_6598,N_6458,N_6406);
nor U6599 (N_6599,N_6493,N_6486);
xnor U6600 (N_6600,N_6484,N_6439);
or U6601 (N_6601,N_6508,N_6553);
nand U6602 (N_6602,N_6515,N_6469);
nand U6603 (N_6603,N_6443,N_6456);
nand U6604 (N_6604,N_6461,N_6506);
xnor U6605 (N_6605,N_6533,N_6539);
nand U6606 (N_6606,N_6485,N_6417);
nand U6607 (N_6607,N_6546,N_6525);
nor U6608 (N_6608,N_6489,N_6512);
nor U6609 (N_6609,N_6496,N_6505);
nor U6610 (N_6610,N_6490,N_6542);
and U6611 (N_6611,N_6441,N_6538);
xor U6612 (N_6612,N_6414,N_6422);
or U6613 (N_6613,N_6491,N_6466);
xor U6614 (N_6614,N_6412,N_6545);
or U6615 (N_6615,N_6423,N_6472);
xor U6616 (N_6616,N_6524,N_6436);
nor U6617 (N_6617,N_6500,N_6403);
and U6618 (N_6618,N_6521,N_6474);
nand U6619 (N_6619,N_6532,N_6523);
or U6620 (N_6620,N_6424,N_6463);
or U6621 (N_6621,N_6492,N_6480);
xor U6622 (N_6622,N_6559,N_6519);
and U6623 (N_6623,N_6497,N_6555);
nor U6624 (N_6624,N_6551,N_6547);
nor U6625 (N_6625,N_6404,N_6548);
xor U6626 (N_6626,N_6509,N_6477);
nand U6627 (N_6627,N_6433,N_6487);
xnor U6628 (N_6628,N_6432,N_6464);
nand U6629 (N_6629,N_6522,N_6426);
nand U6630 (N_6630,N_6427,N_6504);
and U6631 (N_6631,N_6520,N_6516);
nor U6632 (N_6632,N_6517,N_6431);
xnor U6633 (N_6633,N_6425,N_6460);
or U6634 (N_6634,N_6528,N_6518);
nor U6635 (N_6635,N_6452,N_6416);
or U6636 (N_6636,N_6435,N_6459);
or U6637 (N_6637,N_6503,N_6429);
xnor U6638 (N_6638,N_6434,N_6454);
and U6639 (N_6639,N_6444,N_6543);
nand U6640 (N_6640,N_6519,N_6475);
nor U6641 (N_6641,N_6461,N_6512);
xor U6642 (N_6642,N_6422,N_6439);
and U6643 (N_6643,N_6431,N_6445);
and U6644 (N_6644,N_6456,N_6528);
xor U6645 (N_6645,N_6512,N_6452);
and U6646 (N_6646,N_6439,N_6418);
and U6647 (N_6647,N_6461,N_6548);
xnor U6648 (N_6648,N_6557,N_6502);
xnor U6649 (N_6649,N_6547,N_6512);
nand U6650 (N_6650,N_6473,N_6511);
or U6651 (N_6651,N_6435,N_6537);
xor U6652 (N_6652,N_6530,N_6473);
and U6653 (N_6653,N_6522,N_6554);
and U6654 (N_6654,N_6473,N_6487);
xnor U6655 (N_6655,N_6551,N_6441);
nand U6656 (N_6656,N_6551,N_6554);
and U6657 (N_6657,N_6400,N_6552);
xnor U6658 (N_6658,N_6536,N_6530);
or U6659 (N_6659,N_6478,N_6557);
or U6660 (N_6660,N_6446,N_6492);
xor U6661 (N_6661,N_6482,N_6529);
xnor U6662 (N_6662,N_6487,N_6537);
xnor U6663 (N_6663,N_6554,N_6542);
nor U6664 (N_6664,N_6557,N_6490);
and U6665 (N_6665,N_6420,N_6431);
and U6666 (N_6666,N_6442,N_6411);
or U6667 (N_6667,N_6483,N_6457);
xor U6668 (N_6668,N_6535,N_6548);
and U6669 (N_6669,N_6558,N_6400);
and U6670 (N_6670,N_6423,N_6539);
nand U6671 (N_6671,N_6536,N_6531);
xnor U6672 (N_6672,N_6493,N_6475);
nor U6673 (N_6673,N_6535,N_6550);
xnor U6674 (N_6674,N_6484,N_6558);
nor U6675 (N_6675,N_6493,N_6522);
xor U6676 (N_6676,N_6531,N_6462);
xnor U6677 (N_6677,N_6511,N_6523);
and U6678 (N_6678,N_6549,N_6413);
nor U6679 (N_6679,N_6412,N_6421);
xor U6680 (N_6680,N_6547,N_6533);
nand U6681 (N_6681,N_6545,N_6415);
and U6682 (N_6682,N_6522,N_6420);
or U6683 (N_6683,N_6553,N_6503);
xor U6684 (N_6684,N_6415,N_6458);
xor U6685 (N_6685,N_6474,N_6479);
or U6686 (N_6686,N_6404,N_6454);
nand U6687 (N_6687,N_6556,N_6559);
or U6688 (N_6688,N_6518,N_6509);
xor U6689 (N_6689,N_6556,N_6413);
and U6690 (N_6690,N_6433,N_6555);
nand U6691 (N_6691,N_6437,N_6550);
xor U6692 (N_6692,N_6407,N_6525);
nand U6693 (N_6693,N_6485,N_6429);
nor U6694 (N_6694,N_6550,N_6543);
and U6695 (N_6695,N_6528,N_6500);
nand U6696 (N_6696,N_6446,N_6414);
nand U6697 (N_6697,N_6408,N_6445);
nand U6698 (N_6698,N_6432,N_6545);
and U6699 (N_6699,N_6416,N_6431);
and U6700 (N_6700,N_6554,N_6461);
xor U6701 (N_6701,N_6505,N_6462);
nand U6702 (N_6702,N_6521,N_6548);
nor U6703 (N_6703,N_6430,N_6529);
nor U6704 (N_6704,N_6492,N_6469);
nand U6705 (N_6705,N_6504,N_6524);
xor U6706 (N_6706,N_6427,N_6407);
nor U6707 (N_6707,N_6544,N_6530);
or U6708 (N_6708,N_6545,N_6431);
nand U6709 (N_6709,N_6511,N_6488);
nand U6710 (N_6710,N_6539,N_6537);
and U6711 (N_6711,N_6490,N_6441);
or U6712 (N_6712,N_6545,N_6420);
nand U6713 (N_6713,N_6476,N_6408);
or U6714 (N_6714,N_6496,N_6410);
or U6715 (N_6715,N_6536,N_6475);
xnor U6716 (N_6716,N_6549,N_6435);
and U6717 (N_6717,N_6448,N_6518);
nor U6718 (N_6718,N_6495,N_6420);
and U6719 (N_6719,N_6546,N_6496);
nor U6720 (N_6720,N_6682,N_6716);
nand U6721 (N_6721,N_6674,N_6715);
or U6722 (N_6722,N_6713,N_6608);
xnor U6723 (N_6723,N_6574,N_6630);
or U6724 (N_6724,N_6647,N_6579);
or U6725 (N_6725,N_6623,N_6650);
nand U6726 (N_6726,N_6569,N_6649);
nand U6727 (N_6727,N_6576,N_6658);
and U6728 (N_6728,N_6560,N_6690);
and U6729 (N_6729,N_6667,N_6693);
nand U6730 (N_6730,N_6592,N_6669);
or U6731 (N_6731,N_6666,N_6645);
nand U6732 (N_6732,N_6708,N_6718);
and U6733 (N_6733,N_6598,N_6611);
and U6734 (N_6734,N_6678,N_6565);
xor U6735 (N_6735,N_6656,N_6607);
nor U6736 (N_6736,N_6651,N_6627);
or U6737 (N_6737,N_6590,N_6687);
nand U6738 (N_6738,N_6573,N_6706);
nand U6739 (N_6739,N_6683,N_6717);
or U6740 (N_6740,N_6566,N_6616);
xnor U6741 (N_6741,N_6695,N_6652);
xor U6742 (N_6742,N_6660,N_6614);
xnor U6743 (N_6743,N_6628,N_6671);
or U6744 (N_6744,N_6668,N_6578);
nor U6745 (N_6745,N_6691,N_6584);
nor U6746 (N_6746,N_6620,N_6684);
xor U6747 (N_6747,N_6585,N_6700);
nor U6748 (N_6748,N_6696,N_6698);
and U6749 (N_6749,N_6679,N_6634);
nor U6750 (N_6750,N_6655,N_6665);
nand U6751 (N_6751,N_6653,N_6638);
and U6752 (N_6752,N_6694,N_6680);
nor U6753 (N_6753,N_6632,N_6625);
nor U6754 (N_6754,N_6677,N_6676);
nor U6755 (N_6755,N_6577,N_6613);
nand U6756 (N_6756,N_6575,N_6563);
or U6757 (N_6757,N_6685,N_6709);
xnor U6758 (N_6758,N_6640,N_6600);
or U6759 (N_6759,N_6712,N_6639);
or U6760 (N_6760,N_6597,N_6701);
or U6761 (N_6761,N_6692,N_6587);
nor U6762 (N_6762,N_6681,N_6619);
xor U6763 (N_6763,N_6703,N_6641);
nor U6764 (N_6764,N_6621,N_6675);
nor U6765 (N_6765,N_6705,N_6561);
or U6766 (N_6766,N_6648,N_6661);
nor U6767 (N_6767,N_6711,N_6606);
nor U6768 (N_6768,N_6672,N_6605);
nor U6769 (N_6769,N_6688,N_6588);
nand U6770 (N_6770,N_6626,N_6670);
nor U6771 (N_6771,N_6654,N_6644);
nor U6772 (N_6772,N_6591,N_6699);
nor U6773 (N_6773,N_6593,N_6702);
nor U6774 (N_6774,N_6599,N_6646);
nand U6775 (N_6775,N_6637,N_6689);
nand U6776 (N_6776,N_6562,N_6617);
and U6777 (N_6777,N_6615,N_6572);
xor U6778 (N_6778,N_6612,N_6707);
or U6779 (N_6779,N_6697,N_6582);
or U6780 (N_6780,N_6642,N_6581);
or U6781 (N_6781,N_6609,N_6571);
nand U6782 (N_6782,N_6568,N_6586);
xor U6783 (N_6783,N_6657,N_6610);
and U6784 (N_6784,N_6622,N_6714);
and U6785 (N_6785,N_6580,N_6564);
or U6786 (N_6786,N_6629,N_6618);
nor U6787 (N_6787,N_6570,N_6643);
xnor U6788 (N_6788,N_6604,N_6601);
xor U6789 (N_6789,N_6589,N_6686);
nor U6790 (N_6790,N_6633,N_6673);
nand U6791 (N_6791,N_6631,N_6659);
nand U6792 (N_6792,N_6595,N_6662);
or U6793 (N_6793,N_6602,N_6704);
nor U6794 (N_6794,N_6719,N_6594);
nand U6795 (N_6795,N_6636,N_6596);
nand U6796 (N_6796,N_6583,N_6624);
and U6797 (N_6797,N_6635,N_6710);
xor U6798 (N_6798,N_6567,N_6664);
xor U6799 (N_6799,N_6603,N_6663);
and U6800 (N_6800,N_6644,N_6603);
or U6801 (N_6801,N_6593,N_6711);
or U6802 (N_6802,N_6652,N_6604);
nor U6803 (N_6803,N_6657,N_6679);
or U6804 (N_6804,N_6580,N_6660);
nor U6805 (N_6805,N_6600,N_6562);
nor U6806 (N_6806,N_6676,N_6623);
xnor U6807 (N_6807,N_6653,N_6655);
and U6808 (N_6808,N_6638,N_6687);
nor U6809 (N_6809,N_6624,N_6597);
and U6810 (N_6810,N_6685,N_6651);
and U6811 (N_6811,N_6624,N_6587);
and U6812 (N_6812,N_6684,N_6562);
nor U6813 (N_6813,N_6683,N_6675);
nor U6814 (N_6814,N_6573,N_6569);
xnor U6815 (N_6815,N_6645,N_6617);
and U6816 (N_6816,N_6563,N_6706);
nor U6817 (N_6817,N_6588,N_6563);
xor U6818 (N_6818,N_6604,N_6571);
and U6819 (N_6819,N_6573,N_6604);
xnor U6820 (N_6820,N_6621,N_6637);
and U6821 (N_6821,N_6690,N_6635);
or U6822 (N_6822,N_6692,N_6603);
nand U6823 (N_6823,N_6718,N_6565);
or U6824 (N_6824,N_6677,N_6589);
nor U6825 (N_6825,N_6581,N_6579);
or U6826 (N_6826,N_6569,N_6653);
or U6827 (N_6827,N_6667,N_6607);
nor U6828 (N_6828,N_6621,N_6660);
and U6829 (N_6829,N_6564,N_6574);
nand U6830 (N_6830,N_6663,N_6626);
xnor U6831 (N_6831,N_6650,N_6686);
or U6832 (N_6832,N_6560,N_6593);
nor U6833 (N_6833,N_6714,N_6630);
xor U6834 (N_6834,N_6578,N_6628);
xnor U6835 (N_6835,N_6615,N_6707);
or U6836 (N_6836,N_6716,N_6705);
xor U6837 (N_6837,N_6566,N_6600);
and U6838 (N_6838,N_6645,N_6688);
or U6839 (N_6839,N_6617,N_6568);
xor U6840 (N_6840,N_6572,N_6625);
or U6841 (N_6841,N_6569,N_6670);
and U6842 (N_6842,N_6678,N_6643);
nand U6843 (N_6843,N_6670,N_6655);
or U6844 (N_6844,N_6677,N_6661);
nor U6845 (N_6845,N_6599,N_6705);
and U6846 (N_6846,N_6648,N_6707);
or U6847 (N_6847,N_6623,N_6593);
xnor U6848 (N_6848,N_6621,N_6685);
nand U6849 (N_6849,N_6566,N_6620);
nand U6850 (N_6850,N_6656,N_6680);
or U6851 (N_6851,N_6620,N_6605);
xnor U6852 (N_6852,N_6712,N_6619);
nor U6853 (N_6853,N_6590,N_6622);
nand U6854 (N_6854,N_6642,N_6706);
or U6855 (N_6855,N_6689,N_6714);
nor U6856 (N_6856,N_6621,N_6707);
or U6857 (N_6857,N_6703,N_6645);
nor U6858 (N_6858,N_6629,N_6561);
or U6859 (N_6859,N_6610,N_6700);
xor U6860 (N_6860,N_6705,N_6631);
or U6861 (N_6861,N_6683,N_6645);
nand U6862 (N_6862,N_6666,N_6606);
nand U6863 (N_6863,N_6687,N_6677);
nand U6864 (N_6864,N_6669,N_6597);
or U6865 (N_6865,N_6707,N_6664);
and U6866 (N_6866,N_6636,N_6639);
xnor U6867 (N_6867,N_6665,N_6634);
nor U6868 (N_6868,N_6682,N_6615);
or U6869 (N_6869,N_6668,N_6681);
and U6870 (N_6870,N_6660,N_6690);
xor U6871 (N_6871,N_6596,N_6681);
nor U6872 (N_6872,N_6619,N_6580);
and U6873 (N_6873,N_6567,N_6569);
xnor U6874 (N_6874,N_6602,N_6665);
or U6875 (N_6875,N_6704,N_6638);
nand U6876 (N_6876,N_6674,N_6701);
and U6877 (N_6877,N_6600,N_6667);
nand U6878 (N_6878,N_6640,N_6696);
and U6879 (N_6879,N_6678,N_6637);
nor U6880 (N_6880,N_6753,N_6786);
xor U6881 (N_6881,N_6818,N_6754);
nand U6882 (N_6882,N_6758,N_6853);
xnor U6883 (N_6883,N_6774,N_6802);
nand U6884 (N_6884,N_6816,N_6827);
or U6885 (N_6885,N_6746,N_6830);
and U6886 (N_6886,N_6727,N_6834);
nor U6887 (N_6887,N_6809,N_6726);
and U6888 (N_6888,N_6879,N_6783);
nor U6889 (N_6889,N_6843,N_6878);
nor U6890 (N_6890,N_6870,N_6750);
or U6891 (N_6891,N_6864,N_6781);
nor U6892 (N_6892,N_6771,N_6728);
or U6893 (N_6893,N_6779,N_6875);
nand U6894 (N_6894,N_6787,N_6757);
or U6895 (N_6895,N_6840,N_6838);
xor U6896 (N_6896,N_6831,N_6729);
nor U6897 (N_6897,N_6814,N_6862);
and U6898 (N_6898,N_6720,N_6723);
nand U6899 (N_6899,N_6833,N_6795);
nor U6900 (N_6900,N_6798,N_6822);
xor U6901 (N_6901,N_6744,N_6734);
and U6902 (N_6902,N_6841,N_6839);
and U6903 (N_6903,N_6749,N_6866);
and U6904 (N_6904,N_6731,N_6776);
nand U6905 (N_6905,N_6836,N_6860);
or U6906 (N_6906,N_6855,N_6764);
nand U6907 (N_6907,N_6785,N_6821);
and U6908 (N_6908,N_6807,N_6765);
nand U6909 (N_6909,N_6782,N_6763);
or U6910 (N_6910,N_6722,N_6861);
xor U6911 (N_6911,N_6872,N_6767);
nor U6912 (N_6912,N_6778,N_6773);
nor U6913 (N_6913,N_6751,N_6733);
or U6914 (N_6914,N_6837,N_6748);
nor U6915 (N_6915,N_6825,N_6777);
nand U6916 (N_6916,N_6817,N_6747);
or U6917 (N_6917,N_6819,N_6732);
or U6918 (N_6918,N_6775,N_6806);
xor U6919 (N_6919,N_6868,N_6770);
nor U6920 (N_6920,N_6730,N_6796);
or U6921 (N_6921,N_6736,N_6735);
and U6922 (N_6922,N_6865,N_6812);
or U6923 (N_6923,N_6784,N_6808);
and U6924 (N_6924,N_6755,N_6801);
nor U6925 (N_6925,N_6725,N_6856);
and U6926 (N_6926,N_6863,N_6762);
nand U6927 (N_6927,N_6799,N_6846);
and U6928 (N_6928,N_6791,N_6845);
xnor U6929 (N_6929,N_6790,N_6738);
xnor U6930 (N_6930,N_6828,N_6760);
xor U6931 (N_6931,N_6852,N_6829);
xnor U6932 (N_6932,N_6874,N_6844);
and U6933 (N_6933,N_6857,N_6854);
xnor U6934 (N_6934,N_6850,N_6737);
and U6935 (N_6935,N_6849,N_6803);
xnor U6936 (N_6936,N_6724,N_6823);
and U6937 (N_6937,N_6805,N_6813);
xor U6938 (N_6938,N_6780,N_6804);
and U6939 (N_6939,N_6769,N_6811);
nand U6940 (N_6940,N_6794,N_6873);
or U6941 (N_6941,N_6797,N_6826);
nor U6942 (N_6942,N_6789,N_6788);
xor U6943 (N_6943,N_6792,N_6721);
nand U6944 (N_6944,N_6876,N_6772);
or U6945 (N_6945,N_6745,N_6851);
nand U6946 (N_6946,N_6756,N_6871);
nand U6947 (N_6947,N_6742,N_6869);
or U6948 (N_6948,N_6761,N_6824);
and U6949 (N_6949,N_6858,N_6842);
or U6950 (N_6950,N_6768,N_6741);
nand U6951 (N_6951,N_6848,N_6793);
or U6952 (N_6952,N_6835,N_6810);
nor U6953 (N_6953,N_6877,N_6740);
xor U6954 (N_6954,N_6815,N_6847);
xor U6955 (N_6955,N_6832,N_6752);
and U6956 (N_6956,N_6859,N_6820);
xnor U6957 (N_6957,N_6739,N_6867);
and U6958 (N_6958,N_6766,N_6800);
xnor U6959 (N_6959,N_6759,N_6743);
or U6960 (N_6960,N_6828,N_6845);
nor U6961 (N_6961,N_6810,N_6752);
and U6962 (N_6962,N_6776,N_6850);
nor U6963 (N_6963,N_6732,N_6860);
or U6964 (N_6964,N_6794,N_6830);
nor U6965 (N_6965,N_6843,N_6799);
and U6966 (N_6966,N_6745,N_6870);
xnor U6967 (N_6967,N_6787,N_6802);
and U6968 (N_6968,N_6750,N_6741);
and U6969 (N_6969,N_6789,N_6855);
and U6970 (N_6970,N_6730,N_6803);
and U6971 (N_6971,N_6763,N_6858);
xor U6972 (N_6972,N_6747,N_6821);
and U6973 (N_6973,N_6734,N_6732);
nand U6974 (N_6974,N_6740,N_6777);
nor U6975 (N_6975,N_6865,N_6788);
or U6976 (N_6976,N_6760,N_6819);
and U6977 (N_6977,N_6783,N_6771);
nand U6978 (N_6978,N_6784,N_6845);
and U6979 (N_6979,N_6780,N_6865);
or U6980 (N_6980,N_6859,N_6865);
or U6981 (N_6981,N_6745,N_6733);
and U6982 (N_6982,N_6822,N_6858);
xor U6983 (N_6983,N_6862,N_6753);
nor U6984 (N_6984,N_6842,N_6821);
and U6985 (N_6985,N_6811,N_6752);
and U6986 (N_6986,N_6754,N_6838);
nand U6987 (N_6987,N_6729,N_6862);
nand U6988 (N_6988,N_6750,N_6789);
or U6989 (N_6989,N_6830,N_6873);
nand U6990 (N_6990,N_6776,N_6827);
or U6991 (N_6991,N_6767,N_6727);
nand U6992 (N_6992,N_6754,N_6738);
xnor U6993 (N_6993,N_6820,N_6752);
and U6994 (N_6994,N_6837,N_6740);
and U6995 (N_6995,N_6813,N_6751);
xor U6996 (N_6996,N_6774,N_6793);
or U6997 (N_6997,N_6767,N_6756);
nand U6998 (N_6998,N_6851,N_6750);
xnor U6999 (N_6999,N_6857,N_6845);
and U7000 (N_7000,N_6838,N_6774);
xor U7001 (N_7001,N_6765,N_6784);
or U7002 (N_7002,N_6745,N_6803);
or U7003 (N_7003,N_6748,N_6735);
or U7004 (N_7004,N_6733,N_6858);
xnor U7005 (N_7005,N_6767,N_6742);
nand U7006 (N_7006,N_6878,N_6819);
nor U7007 (N_7007,N_6727,N_6749);
nand U7008 (N_7008,N_6749,N_6821);
nor U7009 (N_7009,N_6747,N_6858);
xor U7010 (N_7010,N_6873,N_6771);
or U7011 (N_7011,N_6744,N_6829);
and U7012 (N_7012,N_6804,N_6731);
and U7013 (N_7013,N_6875,N_6831);
or U7014 (N_7014,N_6735,N_6839);
nand U7015 (N_7015,N_6861,N_6790);
xnor U7016 (N_7016,N_6760,N_6876);
and U7017 (N_7017,N_6791,N_6782);
nand U7018 (N_7018,N_6745,N_6749);
or U7019 (N_7019,N_6845,N_6811);
and U7020 (N_7020,N_6794,N_6785);
xnor U7021 (N_7021,N_6762,N_6764);
or U7022 (N_7022,N_6733,N_6801);
or U7023 (N_7023,N_6794,N_6759);
nand U7024 (N_7024,N_6834,N_6748);
or U7025 (N_7025,N_6804,N_6825);
nor U7026 (N_7026,N_6729,N_6849);
xor U7027 (N_7027,N_6860,N_6768);
nand U7028 (N_7028,N_6787,N_6828);
nand U7029 (N_7029,N_6762,N_6876);
nand U7030 (N_7030,N_6743,N_6831);
and U7031 (N_7031,N_6860,N_6721);
nand U7032 (N_7032,N_6859,N_6796);
nand U7033 (N_7033,N_6776,N_6785);
nor U7034 (N_7034,N_6841,N_6788);
nor U7035 (N_7035,N_6785,N_6759);
xnor U7036 (N_7036,N_6759,N_6767);
and U7037 (N_7037,N_6865,N_6782);
nor U7038 (N_7038,N_6854,N_6852);
nand U7039 (N_7039,N_6852,N_6822);
xnor U7040 (N_7040,N_6938,N_6992);
and U7041 (N_7041,N_6960,N_6946);
nor U7042 (N_7042,N_6950,N_6895);
nand U7043 (N_7043,N_6997,N_6922);
xnor U7044 (N_7044,N_6903,N_7001);
or U7045 (N_7045,N_7000,N_6885);
xnor U7046 (N_7046,N_6906,N_6988);
xor U7047 (N_7047,N_6959,N_7031);
and U7048 (N_7048,N_6970,N_6886);
and U7049 (N_7049,N_6991,N_6894);
nand U7050 (N_7050,N_6899,N_7002);
nor U7051 (N_7051,N_6928,N_6985);
or U7052 (N_7052,N_6882,N_6890);
nor U7053 (N_7053,N_6986,N_6915);
and U7054 (N_7054,N_6980,N_6943);
xor U7055 (N_7055,N_7029,N_6995);
xor U7056 (N_7056,N_6926,N_7005);
xnor U7057 (N_7057,N_6956,N_6896);
or U7058 (N_7058,N_6919,N_7035);
and U7059 (N_7059,N_7004,N_7026);
xnor U7060 (N_7060,N_6936,N_6880);
nor U7061 (N_7061,N_6898,N_6884);
nand U7062 (N_7062,N_6908,N_7010);
and U7063 (N_7063,N_7023,N_6920);
and U7064 (N_7064,N_7017,N_6923);
nand U7065 (N_7065,N_6994,N_7030);
or U7066 (N_7066,N_6955,N_6989);
xnor U7067 (N_7067,N_6982,N_6953);
or U7068 (N_7068,N_6999,N_7009);
xnor U7069 (N_7069,N_6973,N_7037);
xor U7070 (N_7070,N_6891,N_6993);
or U7071 (N_7071,N_6947,N_6962);
nand U7072 (N_7072,N_6921,N_6961);
or U7073 (N_7073,N_6957,N_6912);
and U7074 (N_7074,N_6935,N_7014);
nor U7075 (N_7075,N_7018,N_6978);
xor U7076 (N_7076,N_7008,N_6889);
nor U7077 (N_7077,N_6881,N_6941);
and U7078 (N_7078,N_6925,N_6937);
or U7079 (N_7079,N_6969,N_6887);
or U7080 (N_7080,N_6954,N_6967);
or U7081 (N_7081,N_7016,N_6944);
and U7082 (N_7082,N_6975,N_6902);
or U7083 (N_7083,N_6974,N_6966);
xnor U7084 (N_7084,N_6952,N_6996);
nand U7085 (N_7085,N_6927,N_6984);
xnor U7086 (N_7086,N_6901,N_6892);
nor U7087 (N_7087,N_6958,N_7038);
nand U7088 (N_7088,N_7007,N_6940);
and U7089 (N_7089,N_6917,N_6964);
nor U7090 (N_7090,N_6945,N_6951);
nand U7091 (N_7091,N_6971,N_6911);
xnor U7092 (N_7092,N_6968,N_6897);
nor U7093 (N_7093,N_6931,N_6888);
nand U7094 (N_7094,N_6998,N_6990);
or U7095 (N_7095,N_7021,N_7032);
and U7096 (N_7096,N_6900,N_6907);
xor U7097 (N_7097,N_6942,N_7028);
or U7098 (N_7098,N_7020,N_7013);
nand U7099 (N_7099,N_6913,N_6983);
nor U7100 (N_7100,N_7015,N_6930);
nor U7101 (N_7101,N_6976,N_6972);
and U7102 (N_7102,N_6910,N_6883);
nor U7103 (N_7103,N_6909,N_7011);
xor U7104 (N_7104,N_7019,N_6939);
or U7105 (N_7105,N_6914,N_7034);
and U7106 (N_7106,N_7006,N_6949);
nor U7107 (N_7107,N_6924,N_7027);
xnor U7108 (N_7108,N_6918,N_7024);
xnor U7109 (N_7109,N_7025,N_6916);
nand U7110 (N_7110,N_6981,N_6929);
nor U7111 (N_7111,N_7033,N_6934);
or U7112 (N_7112,N_7022,N_6904);
or U7113 (N_7113,N_7039,N_7003);
nand U7114 (N_7114,N_6948,N_6905);
or U7115 (N_7115,N_6987,N_6963);
or U7116 (N_7116,N_7012,N_6893);
and U7117 (N_7117,N_6979,N_7036);
or U7118 (N_7118,N_6933,N_6965);
xor U7119 (N_7119,N_6977,N_6932);
xnor U7120 (N_7120,N_6884,N_7019);
xnor U7121 (N_7121,N_6956,N_6910);
nor U7122 (N_7122,N_6919,N_6946);
nor U7123 (N_7123,N_6884,N_6961);
or U7124 (N_7124,N_6897,N_7034);
xor U7125 (N_7125,N_6940,N_6966);
or U7126 (N_7126,N_6886,N_6930);
or U7127 (N_7127,N_6926,N_6980);
and U7128 (N_7128,N_7017,N_7010);
and U7129 (N_7129,N_6909,N_6914);
nand U7130 (N_7130,N_6892,N_6904);
or U7131 (N_7131,N_7006,N_6936);
xor U7132 (N_7132,N_6986,N_6958);
nand U7133 (N_7133,N_6989,N_6957);
xnor U7134 (N_7134,N_7033,N_6979);
and U7135 (N_7135,N_6947,N_6885);
and U7136 (N_7136,N_7015,N_6948);
xnor U7137 (N_7137,N_7006,N_6946);
or U7138 (N_7138,N_6890,N_6885);
or U7139 (N_7139,N_7012,N_6964);
or U7140 (N_7140,N_6884,N_6922);
and U7141 (N_7141,N_6918,N_6943);
and U7142 (N_7142,N_6962,N_7019);
and U7143 (N_7143,N_7018,N_6883);
or U7144 (N_7144,N_6940,N_6994);
nor U7145 (N_7145,N_6986,N_6886);
nor U7146 (N_7146,N_6931,N_6986);
nand U7147 (N_7147,N_6948,N_6986);
nor U7148 (N_7148,N_6955,N_6892);
or U7149 (N_7149,N_7031,N_6932);
nor U7150 (N_7150,N_6995,N_6907);
and U7151 (N_7151,N_6948,N_7016);
xnor U7152 (N_7152,N_7002,N_6906);
and U7153 (N_7153,N_6953,N_6940);
nand U7154 (N_7154,N_6957,N_7020);
nand U7155 (N_7155,N_7011,N_6951);
and U7156 (N_7156,N_6930,N_6943);
xnor U7157 (N_7157,N_6923,N_6917);
and U7158 (N_7158,N_7005,N_6948);
xor U7159 (N_7159,N_6910,N_6969);
nor U7160 (N_7160,N_6918,N_6881);
xnor U7161 (N_7161,N_7003,N_6965);
and U7162 (N_7162,N_6939,N_6932);
nand U7163 (N_7163,N_6933,N_6938);
nor U7164 (N_7164,N_7020,N_6903);
nor U7165 (N_7165,N_6991,N_6885);
xnor U7166 (N_7166,N_7013,N_6944);
or U7167 (N_7167,N_6916,N_7024);
and U7168 (N_7168,N_6942,N_7032);
and U7169 (N_7169,N_7029,N_7022);
and U7170 (N_7170,N_6953,N_6931);
nand U7171 (N_7171,N_6972,N_6990);
nor U7172 (N_7172,N_6966,N_6883);
xor U7173 (N_7173,N_6960,N_7022);
nand U7174 (N_7174,N_6990,N_6942);
or U7175 (N_7175,N_6900,N_6946);
or U7176 (N_7176,N_6885,N_6895);
or U7177 (N_7177,N_6997,N_6987);
or U7178 (N_7178,N_6935,N_6895);
nor U7179 (N_7179,N_6954,N_7037);
nand U7180 (N_7180,N_6977,N_6897);
xor U7181 (N_7181,N_6911,N_6882);
nor U7182 (N_7182,N_7032,N_6972);
and U7183 (N_7183,N_6897,N_6957);
and U7184 (N_7184,N_6887,N_6956);
xor U7185 (N_7185,N_7036,N_6931);
nor U7186 (N_7186,N_7011,N_6993);
xor U7187 (N_7187,N_6982,N_6957);
xor U7188 (N_7188,N_7036,N_6954);
nand U7189 (N_7189,N_6985,N_6977);
or U7190 (N_7190,N_7020,N_7010);
xor U7191 (N_7191,N_6911,N_6986);
xor U7192 (N_7192,N_6981,N_6942);
nor U7193 (N_7193,N_6936,N_6989);
and U7194 (N_7194,N_6913,N_7031);
nor U7195 (N_7195,N_7027,N_6890);
nand U7196 (N_7196,N_6956,N_6961);
nor U7197 (N_7197,N_6937,N_7035);
and U7198 (N_7198,N_6975,N_7002);
or U7199 (N_7199,N_6995,N_6978);
xnor U7200 (N_7200,N_7072,N_7145);
or U7201 (N_7201,N_7050,N_7067);
or U7202 (N_7202,N_7074,N_7129);
or U7203 (N_7203,N_7149,N_7070);
or U7204 (N_7204,N_7097,N_7046);
or U7205 (N_7205,N_7068,N_7196);
nand U7206 (N_7206,N_7141,N_7102);
nor U7207 (N_7207,N_7194,N_7139);
and U7208 (N_7208,N_7047,N_7041);
xnor U7209 (N_7209,N_7126,N_7083);
nand U7210 (N_7210,N_7190,N_7091);
nand U7211 (N_7211,N_7100,N_7099);
nand U7212 (N_7212,N_7175,N_7191);
and U7213 (N_7213,N_7110,N_7171);
and U7214 (N_7214,N_7106,N_7147);
or U7215 (N_7215,N_7179,N_7162);
nor U7216 (N_7216,N_7136,N_7119);
xor U7217 (N_7217,N_7157,N_7195);
nand U7218 (N_7218,N_7154,N_7057);
nor U7219 (N_7219,N_7174,N_7095);
nand U7220 (N_7220,N_7111,N_7121);
and U7221 (N_7221,N_7082,N_7058);
and U7222 (N_7222,N_7170,N_7138);
xor U7223 (N_7223,N_7090,N_7164);
xnor U7224 (N_7224,N_7186,N_7115);
nand U7225 (N_7225,N_7081,N_7167);
nor U7226 (N_7226,N_7084,N_7131);
and U7227 (N_7227,N_7188,N_7159);
nor U7228 (N_7228,N_7108,N_7112);
and U7229 (N_7229,N_7080,N_7069);
and U7230 (N_7230,N_7150,N_7061);
nand U7231 (N_7231,N_7189,N_7182);
nor U7232 (N_7232,N_7042,N_7076);
or U7233 (N_7233,N_7176,N_7053);
and U7234 (N_7234,N_7087,N_7144);
nor U7235 (N_7235,N_7140,N_7142);
and U7236 (N_7236,N_7060,N_7079);
or U7237 (N_7237,N_7077,N_7094);
xor U7238 (N_7238,N_7064,N_7107);
nand U7239 (N_7239,N_7166,N_7146);
and U7240 (N_7240,N_7173,N_7089);
nor U7241 (N_7241,N_7130,N_7105);
and U7242 (N_7242,N_7104,N_7052);
and U7243 (N_7243,N_7184,N_7181);
or U7244 (N_7244,N_7093,N_7177);
or U7245 (N_7245,N_7043,N_7143);
xor U7246 (N_7246,N_7169,N_7075);
nand U7247 (N_7247,N_7096,N_7122);
xnor U7248 (N_7248,N_7168,N_7065);
xnor U7249 (N_7249,N_7133,N_7045);
xnor U7250 (N_7250,N_7180,N_7098);
and U7251 (N_7251,N_7199,N_7055);
nor U7252 (N_7252,N_7160,N_7148);
and U7253 (N_7253,N_7063,N_7135);
nor U7254 (N_7254,N_7156,N_7128);
and U7255 (N_7255,N_7086,N_7187);
nand U7256 (N_7256,N_7103,N_7153);
or U7257 (N_7257,N_7051,N_7049);
nor U7258 (N_7258,N_7123,N_7165);
or U7259 (N_7259,N_7092,N_7101);
and U7260 (N_7260,N_7193,N_7132);
nor U7261 (N_7261,N_7134,N_7071);
nand U7262 (N_7262,N_7198,N_7172);
nor U7263 (N_7263,N_7116,N_7088);
nand U7264 (N_7264,N_7127,N_7183);
and U7265 (N_7265,N_7161,N_7073);
nand U7266 (N_7266,N_7155,N_7185);
or U7267 (N_7267,N_7124,N_7109);
nor U7268 (N_7268,N_7085,N_7125);
nor U7269 (N_7269,N_7117,N_7192);
nand U7270 (N_7270,N_7056,N_7113);
xor U7271 (N_7271,N_7066,N_7152);
nor U7272 (N_7272,N_7078,N_7114);
nand U7273 (N_7273,N_7197,N_7118);
or U7274 (N_7274,N_7163,N_7054);
and U7275 (N_7275,N_7120,N_7040);
xnor U7276 (N_7276,N_7151,N_7158);
or U7277 (N_7277,N_7178,N_7044);
nor U7278 (N_7278,N_7059,N_7137);
xnor U7279 (N_7279,N_7048,N_7062);
and U7280 (N_7280,N_7147,N_7174);
xnor U7281 (N_7281,N_7045,N_7102);
nor U7282 (N_7282,N_7101,N_7087);
and U7283 (N_7283,N_7168,N_7109);
nor U7284 (N_7284,N_7121,N_7182);
or U7285 (N_7285,N_7103,N_7082);
xnor U7286 (N_7286,N_7052,N_7071);
and U7287 (N_7287,N_7166,N_7076);
nand U7288 (N_7288,N_7072,N_7058);
and U7289 (N_7289,N_7148,N_7117);
nor U7290 (N_7290,N_7083,N_7138);
nor U7291 (N_7291,N_7086,N_7064);
or U7292 (N_7292,N_7095,N_7085);
nand U7293 (N_7293,N_7043,N_7150);
xor U7294 (N_7294,N_7151,N_7119);
nand U7295 (N_7295,N_7062,N_7154);
xnor U7296 (N_7296,N_7167,N_7115);
xor U7297 (N_7297,N_7077,N_7166);
nand U7298 (N_7298,N_7158,N_7055);
nand U7299 (N_7299,N_7171,N_7122);
xor U7300 (N_7300,N_7184,N_7165);
nor U7301 (N_7301,N_7173,N_7157);
xnor U7302 (N_7302,N_7130,N_7107);
nor U7303 (N_7303,N_7113,N_7177);
and U7304 (N_7304,N_7071,N_7131);
and U7305 (N_7305,N_7141,N_7066);
nand U7306 (N_7306,N_7179,N_7195);
nand U7307 (N_7307,N_7161,N_7192);
and U7308 (N_7308,N_7104,N_7078);
and U7309 (N_7309,N_7154,N_7163);
and U7310 (N_7310,N_7095,N_7082);
nand U7311 (N_7311,N_7152,N_7072);
xnor U7312 (N_7312,N_7093,N_7155);
and U7313 (N_7313,N_7083,N_7048);
nor U7314 (N_7314,N_7040,N_7045);
or U7315 (N_7315,N_7169,N_7175);
xnor U7316 (N_7316,N_7085,N_7124);
and U7317 (N_7317,N_7171,N_7191);
or U7318 (N_7318,N_7169,N_7144);
xor U7319 (N_7319,N_7117,N_7057);
and U7320 (N_7320,N_7053,N_7052);
and U7321 (N_7321,N_7183,N_7078);
and U7322 (N_7322,N_7041,N_7119);
nor U7323 (N_7323,N_7129,N_7068);
nand U7324 (N_7324,N_7068,N_7078);
xnor U7325 (N_7325,N_7146,N_7101);
or U7326 (N_7326,N_7144,N_7051);
nand U7327 (N_7327,N_7112,N_7174);
xnor U7328 (N_7328,N_7121,N_7095);
xnor U7329 (N_7329,N_7191,N_7071);
xnor U7330 (N_7330,N_7046,N_7168);
xnor U7331 (N_7331,N_7140,N_7104);
xnor U7332 (N_7332,N_7161,N_7080);
nor U7333 (N_7333,N_7070,N_7170);
or U7334 (N_7334,N_7091,N_7082);
nor U7335 (N_7335,N_7147,N_7187);
or U7336 (N_7336,N_7044,N_7063);
nor U7337 (N_7337,N_7073,N_7189);
or U7338 (N_7338,N_7080,N_7197);
or U7339 (N_7339,N_7150,N_7079);
and U7340 (N_7340,N_7119,N_7130);
nor U7341 (N_7341,N_7125,N_7093);
xor U7342 (N_7342,N_7095,N_7193);
nand U7343 (N_7343,N_7067,N_7082);
or U7344 (N_7344,N_7096,N_7158);
nor U7345 (N_7345,N_7115,N_7087);
and U7346 (N_7346,N_7112,N_7131);
nor U7347 (N_7347,N_7040,N_7100);
or U7348 (N_7348,N_7057,N_7084);
and U7349 (N_7349,N_7181,N_7088);
or U7350 (N_7350,N_7122,N_7078);
and U7351 (N_7351,N_7118,N_7051);
or U7352 (N_7352,N_7148,N_7171);
xnor U7353 (N_7353,N_7095,N_7184);
nor U7354 (N_7354,N_7110,N_7130);
and U7355 (N_7355,N_7118,N_7094);
nand U7356 (N_7356,N_7090,N_7067);
and U7357 (N_7357,N_7180,N_7102);
nand U7358 (N_7358,N_7045,N_7164);
xor U7359 (N_7359,N_7192,N_7188);
or U7360 (N_7360,N_7277,N_7275);
xnor U7361 (N_7361,N_7305,N_7206);
or U7362 (N_7362,N_7251,N_7297);
nor U7363 (N_7363,N_7327,N_7213);
nor U7364 (N_7364,N_7293,N_7210);
nand U7365 (N_7365,N_7328,N_7320);
nand U7366 (N_7366,N_7258,N_7336);
and U7367 (N_7367,N_7240,N_7232);
nand U7368 (N_7368,N_7235,N_7302);
xnor U7369 (N_7369,N_7299,N_7237);
or U7370 (N_7370,N_7223,N_7215);
or U7371 (N_7371,N_7264,N_7250);
or U7372 (N_7372,N_7344,N_7311);
nand U7373 (N_7373,N_7312,N_7291);
and U7374 (N_7374,N_7342,N_7244);
and U7375 (N_7375,N_7321,N_7225);
and U7376 (N_7376,N_7339,N_7203);
and U7377 (N_7377,N_7289,N_7332);
xor U7378 (N_7378,N_7292,N_7241);
and U7379 (N_7379,N_7238,N_7316);
nand U7380 (N_7380,N_7356,N_7208);
and U7381 (N_7381,N_7260,N_7246);
nand U7382 (N_7382,N_7353,N_7284);
nor U7383 (N_7383,N_7247,N_7278);
nor U7384 (N_7384,N_7288,N_7233);
and U7385 (N_7385,N_7211,N_7267);
xnor U7386 (N_7386,N_7347,N_7317);
nor U7387 (N_7387,N_7285,N_7354);
or U7388 (N_7388,N_7352,N_7337);
or U7389 (N_7389,N_7358,N_7214);
or U7390 (N_7390,N_7303,N_7341);
nand U7391 (N_7391,N_7252,N_7338);
or U7392 (N_7392,N_7209,N_7282);
nand U7393 (N_7393,N_7300,N_7221);
or U7394 (N_7394,N_7229,N_7350);
nand U7395 (N_7395,N_7329,N_7242);
nor U7396 (N_7396,N_7217,N_7220);
xor U7397 (N_7397,N_7255,N_7248);
nand U7398 (N_7398,N_7205,N_7330);
or U7399 (N_7399,N_7273,N_7228);
xnor U7400 (N_7400,N_7226,N_7343);
nand U7401 (N_7401,N_7348,N_7243);
or U7402 (N_7402,N_7314,N_7274);
and U7403 (N_7403,N_7310,N_7323);
xnor U7404 (N_7404,N_7334,N_7286);
and U7405 (N_7405,N_7218,N_7201);
nor U7406 (N_7406,N_7234,N_7280);
xnor U7407 (N_7407,N_7325,N_7259);
xor U7408 (N_7408,N_7268,N_7290);
or U7409 (N_7409,N_7324,N_7270);
nand U7410 (N_7410,N_7322,N_7313);
nor U7411 (N_7411,N_7212,N_7295);
or U7412 (N_7412,N_7256,N_7272);
or U7413 (N_7413,N_7222,N_7253);
nand U7414 (N_7414,N_7296,N_7266);
nor U7415 (N_7415,N_7254,N_7331);
xnor U7416 (N_7416,N_7257,N_7304);
nor U7417 (N_7417,N_7281,N_7261);
nor U7418 (N_7418,N_7306,N_7359);
or U7419 (N_7419,N_7351,N_7294);
nand U7420 (N_7420,N_7202,N_7276);
nand U7421 (N_7421,N_7283,N_7224);
and U7422 (N_7422,N_7262,N_7236);
and U7423 (N_7423,N_7219,N_7307);
or U7424 (N_7424,N_7271,N_7357);
and U7425 (N_7425,N_7315,N_7301);
or U7426 (N_7426,N_7279,N_7263);
nand U7427 (N_7427,N_7204,N_7239);
xnor U7428 (N_7428,N_7326,N_7345);
and U7429 (N_7429,N_7340,N_7265);
nor U7430 (N_7430,N_7287,N_7216);
or U7431 (N_7431,N_7319,N_7346);
nand U7432 (N_7432,N_7355,N_7231);
nor U7433 (N_7433,N_7227,N_7318);
nand U7434 (N_7434,N_7298,N_7349);
and U7435 (N_7435,N_7333,N_7335);
or U7436 (N_7436,N_7249,N_7200);
and U7437 (N_7437,N_7245,N_7230);
or U7438 (N_7438,N_7309,N_7207);
nor U7439 (N_7439,N_7308,N_7269);
nor U7440 (N_7440,N_7284,N_7301);
and U7441 (N_7441,N_7300,N_7206);
xnor U7442 (N_7442,N_7214,N_7325);
nand U7443 (N_7443,N_7215,N_7337);
or U7444 (N_7444,N_7320,N_7265);
or U7445 (N_7445,N_7309,N_7266);
or U7446 (N_7446,N_7315,N_7343);
xnor U7447 (N_7447,N_7317,N_7353);
nor U7448 (N_7448,N_7318,N_7283);
or U7449 (N_7449,N_7264,N_7356);
and U7450 (N_7450,N_7319,N_7356);
nor U7451 (N_7451,N_7276,N_7346);
or U7452 (N_7452,N_7252,N_7258);
and U7453 (N_7453,N_7338,N_7261);
xnor U7454 (N_7454,N_7257,N_7256);
xnor U7455 (N_7455,N_7305,N_7200);
or U7456 (N_7456,N_7218,N_7306);
nor U7457 (N_7457,N_7236,N_7295);
and U7458 (N_7458,N_7232,N_7293);
or U7459 (N_7459,N_7238,N_7349);
and U7460 (N_7460,N_7330,N_7337);
or U7461 (N_7461,N_7224,N_7223);
or U7462 (N_7462,N_7306,N_7333);
nor U7463 (N_7463,N_7224,N_7313);
nor U7464 (N_7464,N_7243,N_7250);
nand U7465 (N_7465,N_7302,N_7266);
and U7466 (N_7466,N_7297,N_7282);
xor U7467 (N_7467,N_7341,N_7261);
and U7468 (N_7468,N_7316,N_7322);
nand U7469 (N_7469,N_7337,N_7260);
nand U7470 (N_7470,N_7342,N_7298);
and U7471 (N_7471,N_7268,N_7265);
and U7472 (N_7472,N_7297,N_7295);
or U7473 (N_7473,N_7341,N_7306);
and U7474 (N_7474,N_7276,N_7355);
xor U7475 (N_7475,N_7305,N_7207);
nor U7476 (N_7476,N_7354,N_7260);
or U7477 (N_7477,N_7354,N_7290);
and U7478 (N_7478,N_7237,N_7356);
nand U7479 (N_7479,N_7201,N_7286);
nor U7480 (N_7480,N_7227,N_7210);
xor U7481 (N_7481,N_7203,N_7238);
or U7482 (N_7482,N_7325,N_7251);
and U7483 (N_7483,N_7267,N_7315);
and U7484 (N_7484,N_7333,N_7255);
nand U7485 (N_7485,N_7200,N_7324);
or U7486 (N_7486,N_7292,N_7204);
and U7487 (N_7487,N_7207,N_7312);
or U7488 (N_7488,N_7338,N_7309);
nor U7489 (N_7489,N_7256,N_7355);
or U7490 (N_7490,N_7248,N_7267);
nand U7491 (N_7491,N_7274,N_7275);
xor U7492 (N_7492,N_7329,N_7289);
nor U7493 (N_7493,N_7248,N_7238);
nor U7494 (N_7494,N_7269,N_7234);
nor U7495 (N_7495,N_7346,N_7218);
nand U7496 (N_7496,N_7208,N_7219);
nand U7497 (N_7497,N_7341,N_7221);
or U7498 (N_7498,N_7350,N_7323);
and U7499 (N_7499,N_7295,N_7335);
nand U7500 (N_7500,N_7253,N_7241);
and U7501 (N_7501,N_7200,N_7261);
nand U7502 (N_7502,N_7234,N_7232);
and U7503 (N_7503,N_7346,N_7245);
or U7504 (N_7504,N_7349,N_7267);
and U7505 (N_7505,N_7250,N_7341);
nand U7506 (N_7506,N_7237,N_7232);
nand U7507 (N_7507,N_7239,N_7229);
nand U7508 (N_7508,N_7347,N_7312);
and U7509 (N_7509,N_7305,N_7347);
nand U7510 (N_7510,N_7219,N_7205);
or U7511 (N_7511,N_7269,N_7213);
nor U7512 (N_7512,N_7355,N_7320);
and U7513 (N_7513,N_7255,N_7261);
and U7514 (N_7514,N_7282,N_7279);
or U7515 (N_7515,N_7236,N_7302);
xnor U7516 (N_7516,N_7204,N_7290);
nand U7517 (N_7517,N_7214,N_7281);
and U7518 (N_7518,N_7317,N_7283);
xor U7519 (N_7519,N_7296,N_7313);
or U7520 (N_7520,N_7469,N_7442);
xor U7521 (N_7521,N_7451,N_7386);
nand U7522 (N_7522,N_7473,N_7516);
or U7523 (N_7523,N_7375,N_7455);
nand U7524 (N_7524,N_7437,N_7502);
xor U7525 (N_7525,N_7500,N_7420);
nor U7526 (N_7526,N_7454,N_7394);
nand U7527 (N_7527,N_7362,N_7441);
nand U7528 (N_7528,N_7507,N_7392);
xnor U7529 (N_7529,N_7389,N_7448);
and U7530 (N_7530,N_7511,N_7404);
nor U7531 (N_7531,N_7503,N_7400);
nand U7532 (N_7532,N_7518,N_7369);
nand U7533 (N_7533,N_7373,N_7402);
xnor U7534 (N_7534,N_7427,N_7505);
xnor U7535 (N_7535,N_7364,N_7464);
and U7536 (N_7536,N_7489,N_7498);
xnor U7537 (N_7537,N_7499,N_7467);
and U7538 (N_7538,N_7422,N_7496);
nand U7539 (N_7539,N_7483,N_7478);
or U7540 (N_7540,N_7462,N_7378);
or U7541 (N_7541,N_7419,N_7415);
nor U7542 (N_7542,N_7474,N_7361);
xnor U7543 (N_7543,N_7497,N_7501);
and U7544 (N_7544,N_7433,N_7468);
nand U7545 (N_7545,N_7488,N_7424);
xnor U7546 (N_7546,N_7508,N_7475);
or U7547 (N_7547,N_7363,N_7492);
and U7548 (N_7548,N_7381,N_7396);
xnor U7549 (N_7549,N_7519,N_7494);
and U7550 (N_7550,N_7432,N_7490);
nor U7551 (N_7551,N_7374,N_7379);
xor U7552 (N_7552,N_7382,N_7365);
or U7553 (N_7553,N_7418,N_7436);
xnor U7554 (N_7554,N_7383,N_7449);
or U7555 (N_7555,N_7506,N_7514);
nor U7556 (N_7556,N_7480,N_7510);
or U7557 (N_7557,N_7457,N_7385);
or U7558 (N_7558,N_7367,N_7443);
xor U7559 (N_7559,N_7460,N_7406);
xor U7560 (N_7560,N_7368,N_7513);
and U7561 (N_7561,N_7405,N_7435);
nand U7562 (N_7562,N_7479,N_7459);
or U7563 (N_7563,N_7430,N_7487);
or U7564 (N_7564,N_7412,N_7517);
or U7565 (N_7565,N_7452,N_7472);
or U7566 (N_7566,N_7429,N_7399);
nor U7567 (N_7567,N_7413,N_7384);
and U7568 (N_7568,N_7393,N_7463);
nand U7569 (N_7569,N_7438,N_7376);
nand U7570 (N_7570,N_7471,N_7388);
and U7571 (N_7571,N_7504,N_7421);
or U7572 (N_7572,N_7366,N_7425);
nor U7573 (N_7573,N_7515,N_7447);
nor U7574 (N_7574,N_7409,N_7493);
xnor U7575 (N_7575,N_7445,N_7398);
nor U7576 (N_7576,N_7417,N_7416);
or U7577 (N_7577,N_7484,N_7476);
nor U7578 (N_7578,N_7370,N_7391);
and U7579 (N_7579,N_7509,N_7414);
xor U7580 (N_7580,N_7495,N_7380);
and U7581 (N_7581,N_7360,N_7408);
xor U7582 (N_7582,N_7485,N_7411);
nor U7583 (N_7583,N_7450,N_7423);
or U7584 (N_7584,N_7371,N_7456);
xnor U7585 (N_7585,N_7486,N_7470);
or U7586 (N_7586,N_7395,N_7461);
nand U7587 (N_7587,N_7397,N_7465);
xor U7588 (N_7588,N_7446,N_7512);
and U7589 (N_7589,N_7403,N_7440);
nor U7590 (N_7590,N_7410,N_7482);
or U7591 (N_7591,N_7434,N_7477);
and U7592 (N_7592,N_7401,N_7372);
and U7593 (N_7593,N_7407,N_7439);
xnor U7594 (N_7594,N_7387,N_7453);
nor U7595 (N_7595,N_7481,N_7428);
nand U7596 (N_7596,N_7426,N_7491);
or U7597 (N_7597,N_7377,N_7431);
or U7598 (N_7598,N_7444,N_7390);
or U7599 (N_7599,N_7466,N_7458);
and U7600 (N_7600,N_7409,N_7387);
or U7601 (N_7601,N_7469,N_7420);
xor U7602 (N_7602,N_7393,N_7387);
nor U7603 (N_7603,N_7450,N_7433);
or U7604 (N_7604,N_7518,N_7414);
and U7605 (N_7605,N_7381,N_7464);
or U7606 (N_7606,N_7375,N_7390);
xnor U7607 (N_7607,N_7473,N_7421);
and U7608 (N_7608,N_7454,N_7364);
and U7609 (N_7609,N_7372,N_7378);
and U7610 (N_7610,N_7489,N_7443);
xor U7611 (N_7611,N_7432,N_7455);
xnor U7612 (N_7612,N_7365,N_7478);
xor U7613 (N_7613,N_7481,N_7442);
or U7614 (N_7614,N_7427,N_7499);
and U7615 (N_7615,N_7514,N_7365);
and U7616 (N_7616,N_7466,N_7505);
or U7617 (N_7617,N_7507,N_7470);
nand U7618 (N_7618,N_7362,N_7403);
xnor U7619 (N_7619,N_7431,N_7514);
nor U7620 (N_7620,N_7507,N_7366);
and U7621 (N_7621,N_7517,N_7400);
xnor U7622 (N_7622,N_7480,N_7378);
or U7623 (N_7623,N_7379,N_7365);
xnor U7624 (N_7624,N_7413,N_7406);
nor U7625 (N_7625,N_7498,N_7429);
nand U7626 (N_7626,N_7382,N_7385);
nand U7627 (N_7627,N_7490,N_7386);
nor U7628 (N_7628,N_7411,N_7392);
or U7629 (N_7629,N_7515,N_7384);
or U7630 (N_7630,N_7457,N_7426);
or U7631 (N_7631,N_7471,N_7411);
or U7632 (N_7632,N_7432,N_7368);
nand U7633 (N_7633,N_7368,N_7434);
nand U7634 (N_7634,N_7399,N_7410);
nor U7635 (N_7635,N_7367,N_7438);
nand U7636 (N_7636,N_7384,N_7464);
xnor U7637 (N_7637,N_7417,N_7443);
nand U7638 (N_7638,N_7467,N_7489);
xnor U7639 (N_7639,N_7370,N_7397);
nor U7640 (N_7640,N_7494,N_7424);
xor U7641 (N_7641,N_7488,N_7478);
and U7642 (N_7642,N_7417,N_7380);
nand U7643 (N_7643,N_7493,N_7460);
nor U7644 (N_7644,N_7433,N_7421);
or U7645 (N_7645,N_7478,N_7464);
and U7646 (N_7646,N_7428,N_7375);
and U7647 (N_7647,N_7438,N_7380);
or U7648 (N_7648,N_7467,N_7497);
xor U7649 (N_7649,N_7465,N_7429);
and U7650 (N_7650,N_7458,N_7408);
and U7651 (N_7651,N_7392,N_7406);
nor U7652 (N_7652,N_7444,N_7374);
and U7653 (N_7653,N_7447,N_7362);
or U7654 (N_7654,N_7400,N_7496);
and U7655 (N_7655,N_7462,N_7396);
or U7656 (N_7656,N_7464,N_7411);
nor U7657 (N_7657,N_7469,N_7472);
nand U7658 (N_7658,N_7479,N_7464);
xnor U7659 (N_7659,N_7416,N_7510);
nor U7660 (N_7660,N_7362,N_7468);
xor U7661 (N_7661,N_7380,N_7508);
nand U7662 (N_7662,N_7484,N_7373);
nor U7663 (N_7663,N_7410,N_7404);
and U7664 (N_7664,N_7509,N_7502);
or U7665 (N_7665,N_7439,N_7384);
or U7666 (N_7666,N_7451,N_7491);
nor U7667 (N_7667,N_7503,N_7481);
or U7668 (N_7668,N_7451,N_7382);
and U7669 (N_7669,N_7367,N_7496);
nand U7670 (N_7670,N_7432,N_7404);
and U7671 (N_7671,N_7494,N_7497);
or U7672 (N_7672,N_7426,N_7508);
or U7673 (N_7673,N_7381,N_7514);
nand U7674 (N_7674,N_7426,N_7410);
xnor U7675 (N_7675,N_7424,N_7480);
and U7676 (N_7676,N_7424,N_7475);
xnor U7677 (N_7677,N_7476,N_7383);
nor U7678 (N_7678,N_7369,N_7426);
nand U7679 (N_7679,N_7445,N_7463);
xor U7680 (N_7680,N_7621,N_7664);
nor U7681 (N_7681,N_7678,N_7541);
or U7682 (N_7682,N_7628,N_7554);
nand U7683 (N_7683,N_7633,N_7656);
and U7684 (N_7684,N_7632,N_7679);
nand U7685 (N_7685,N_7596,N_7649);
or U7686 (N_7686,N_7615,N_7545);
xnor U7687 (N_7687,N_7599,N_7673);
nand U7688 (N_7688,N_7666,N_7587);
nand U7689 (N_7689,N_7579,N_7555);
nor U7690 (N_7690,N_7601,N_7524);
nor U7691 (N_7691,N_7648,N_7660);
or U7692 (N_7692,N_7622,N_7607);
or U7693 (N_7693,N_7550,N_7667);
nor U7694 (N_7694,N_7618,N_7677);
nor U7695 (N_7695,N_7563,N_7573);
nor U7696 (N_7696,N_7652,N_7610);
nand U7697 (N_7697,N_7543,N_7551);
xnor U7698 (N_7698,N_7674,N_7576);
xor U7699 (N_7699,N_7523,N_7529);
nor U7700 (N_7700,N_7577,N_7564);
nand U7701 (N_7701,N_7569,N_7591);
nand U7702 (N_7702,N_7560,N_7672);
nor U7703 (N_7703,N_7568,N_7557);
nand U7704 (N_7704,N_7640,N_7631);
nor U7705 (N_7705,N_7534,N_7532);
and U7706 (N_7706,N_7589,N_7556);
xnor U7707 (N_7707,N_7655,N_7586);
nand U7708 (N_7708,N_7604,N_7608);
or U7709 (N_7709,N_7613,N_7606);
nor U7710 (N_7710,N_7583,N_7575);
xor U7711 (N_7711,N_7572,N_7567);
nor U7712 (N_7712,N_7661,N_7566);
xor U7713 (N_7713,N_7641,N_7571);
or U7714 (N_7714,N_7623,N_7647);
nand U7715 (N_7715,N_7605,N_7558);
or U7716 (N_7716,N_7578,N_7539);
nor U7717 (N_7717,N_7562,N_7644);
nand U7718 (N_7718,N_7609,N_7553);
xor U7719 (N_7719,N_7552,N_7593);
and U7720 (N_7720,N_7528,N_7602);
and U7721 (N_7721,N_7559,N_7665);
nor U7722 (N_7722,N_7625,N_7636);
nor U7723 (N_7723,N_7547,N_7630);
or U7724 (N_7724,N_7663,N_7643);
nand U7725 (N_7725,N_7634,N_7581);
nor U7726 (N_7726,N_7670,N_7595);
nor U7727 (N_7727,N_7530,N_7574);
xnor U7728 (N_7728,N_7635,N_7544);
and U7729 (N_7729,N_7637,N_7525);
xor U7730 (N_7730,N_7662,N_7600);
nand U7731 (N_7731,N_7520,N_7542);
or U7732 (N_7732,N_7584,N_7582);
nand U7733 (N_7733,N_7639,N_7597);
xor U7734 (N_7734,N_7646,N_7671);
xor U7735 (N_7735,N_7522,N_7676);
xor U7736 (N_7736,N_7533,N_7540);
nor U7737 (N_7737,N_7653,N_7675);
xnor U7738 (N_7738,N_7620,N_7526);
xor U7739 (N_7739,N_7546,N_7614);
nor U7740 (N_7740,N_7537,N_7626);
nor U7741 (N_7741,N_7651,N_7590);
or U7742 (N_7742,N_7594,N_7531);
nand U7743 (N_7743,N_7603,N_7536);
nor U7744 (N_7744,N_7669,N_7617);
or U7745 (N_7745,N_7592,N_7619);
or U7746 (N_7746,N_7548,N_7521);
or U7747 (N_7747,N_7645,N_7629);
and U7748 (N_7748,N_7585,N_7616);
nor U7749 (N_7749,N_7561,N_7527);
nand U7750 (N_7750,N_7598,N_7588);
or U7751 (N_7751,N_7612,N_7624);
nor U7752 (N_7752,N_7642,N_7654);
nand U7753 (N_7753,N_7549,N_7535);
nor U7754 (N_7754,N_7638,N_7570);
nor U7755 (N_7755,N_7650,N_7565);
nor U7756 (N_7756,N_7611,N_7659);
and U7757 (N_7757,N_7580,N_7657);
xnor U7758 (N_7758,N_7627,N_7658);
nand U7759 (N_7759,N_7538,N_7668);
nor U7760 (N_7760,N_7666,N_7577);
nand U7761 (N_7761,N_7555,N_7529);
xnor U7762 (N_7762,N_7663,N_7600);
xor U7763 (N_7763,N_7678,N_7538);
nor U7764 (N_7764,N_7656,N_7551);
and U7765 (N_7765,N_7551,N_7542);
xnor U7766 (N_7766,N_7653,N_7534);
xor U7767 (N_7767,N_7639,N_7532);
nand U7768 (N_7768,N_7551,N_7534);
nand U7769 (N_7769,N_7592,N_7568);
or U7770 (N_7770,N_7591,N_7557);
or U7771 (N_7771,N_7608,N_7620);
xnor U7772 (N_7772,N_7625,N_7556);
xor U7773 (N_7773,N_7621,N_7606);
xnor U7774 (N_7774,N_7608,N_7649);
or U7775 (N_7775,N_7534,N_7584);
nor U7776 (N_7776,N_7531,N_7579);
nand U7777 (N_7777,N_7640,N_7555);
nand U7778 (N_7778,N_7530,N_7678);
xor U7779 (N_7779,N_7623,N_7541);
nand U7780 (N_7780,N_7571,N_7597);
nand U7781 (N_7781,N_7593,N_7637);
or U7782 (N_7782,N_7569,N_7677);
nand U7783 (N_7783,N_7668,N_7583);
nand U7784 (N_7784,N_7676,N_7575);
nand U7785 (N_7785,N_7590,N_7640);
or U7786 (N_7786,N_7655,N_7601);
nor U7787 (N_7787,N_7643,N_7671);
and U7788 (N_7788,N_7544,N_7600);
nand U7789 (N_7789,N_7638,N_7558);
nor U7790 (N_7790,N_7671,N_7547);
nand U7791 (N_7791,N_7679,N_7669);
nand U7792 (N_7792,N_7661,N_7643);
or U7793 (N_7793,N_7669,N_7533);
or U7794 (N_7794,N_7669,N_7543);
xnor U7795 (N_7795,N_7631,N_7522);
or U7796 (N_7796,N_7607,N_7659);
and U7797 (N_7797,N_7584,N_7661);
nand U7798 (N_7798,N_7584,N_7553);
or U7799 (N_7799,N_7562,N_7525);
xnor U7800 (N_7800,N_7666,N_7664);
or U7801 (N_7801,N_7663,N_7674);
nand U7802 (N_7802,N_7627,N_7609);
or U7803 (N_7803,N_7613,N_7678);
nand U7804 (N_7804,N_7634,N_7537);
or U7805 (N_7805,N_7608,N_7537);
nand U7806 (N_7806,N_7657,N_7643);
or U7807 (N_7807,N_7584,N_7644);
nand U7808 (N_7808,N_7587,N_7637);
nor U7809 (N_7809,N_7625,N_7615);
xor U7810 (N_7810,N_7527,N_7591);
nand U7811 (N_7811,N_7606,N_7641);
or U7812 (N_7812,N_7540,N_7671);
xnor U7813 (N_7813,N_7583,N_7620);
or U7814 (N_7814,N_7530,N_7552);
nor U7815 (N_7815,N_7637,N_7575);
and U7816 (N_7816,N_7633,N_7617);
nand U7817 (N_7817,N_7596,N_7650);
and U7818 (N_7818,N_7534,N_7531);
nand U7819 (N_7819,N_7573,N_7634);
or U7820 (N_7820,N_7642,N_7671);
or U7821 (N_7821,N_7672,N_7546);
xnor U7822 (N_7822,N_7541,N_7591);
and U7823 (N_7823,N_7576,N_7527);
or U7824 (N_7824,N_7585,N_7623);
nand U7825 (N_7825,N_7630,N_7553);
or U7826 (N_7826,N_7597,N_7577);
nand U7827 (N_7827,N_7651,N_7530);
or U7828 (N_7828,N_7536,N_7668);
xnor U7829 (N_7829,N_7570,N_7550);
or U7830 (N_7830,N_7638,N_7553);
and U7831 (N_7831,N_7678,N_7587);
and U7832 (N_7832,N_7592,N_7638);
nand U7833 (N_7833,N_7621,N_7598);
or U7834 (N_7834,N_7649,N_7556);
or U7835 (N_7835,N_7630,N_7585);
or U7836 (N_7836,N_7571,N_7545);
nor U7837 (N_7837,N_7578,N_7573);
xor U7838 (N_7838,N_7531,N_7591);
nor U7839 (N_7839,N_7658,N_7645);
or U7840 (N_7840,N_7792,N_7685);
xnor U7841 (N_7841,N_7717,N_7791);
xnor U7842 (N_7842,N_7813,N_7732);
and U7843 (N_7843,N_7838,N_7693);
xor U7844 (N_7844,N_7686,N_7727);
or U7845 (N_7845,N_7746,N_7698);
nor U7846 (N_7846,N_7702,N_7822);
nor U7847 (N_7847,N_7767,N_7747);
nor U7848 (N_7848,N_7709,N_7785);
and U7849 (N_7849,N_7832,N_7711);
and U7850 (N_7850,N_7815,N_7793);
or U7851 (N_7851,N_7798,N_7824);
or U7852 (N_7852,N_7758,N_7777);
and U7853 (N_7853,N_7722,N_7703);
and U7854 (N_7854,N_7690,N_7837);
or U7855 (N_7855,N_7802,N_7789);
nor U7856 (N_7856,N_7683,N_7765);
nand U7857 (N_7857,N_7740,N_7821);
nor U7858 (N_7858,N_7807,N_7707);
and U7859 (N_7859,N_7819,N_7796);
nand U7860 (N_7860,N_7826,N_7755);
xor U7861 (N_7861,N_7804,N_7719);
and U7862 (N_7862,N_7816,N_7737);
nor U7863 (N_7863,N_7823,N_7766);
nor U7864 (N_7864,N_7771,N_7801);
and U7865 (N_7865,N_7752,N_7811);
and U7866 (N_7866,N_7708,N_7778);
or U7867 (N_7867,N_7809,N_7695);
nand U7868 (N_7868,N_7741,N_7772);
or U7869 (N_7869,N_7699,N_7739);
and U7870 (N_7870,N_7805,N_7720);
xnor U7871 (N_7871,N_7724,N_7692);
and U7872 (N_7872,N_7762,N_7748);
nor U7873 (N_7873,N_7743,N_7757);
nand U7874 (N_7874,N_7728,N_7730);
nand U7875 (N_7875,N_7721,N_7688);
and U7876 (N_7876,N_7713,N_7790);
nor U7877 (N_7877,N_7770,N_7705);
nand U7878 (N_7878,N_7835,N_7803);
nand U7879 (N_7879,N_7818,N_7726);
and U7880 (N_7880,N_7806,N_7782);
or U7881 (N_7881,N_7714,N_7750);
nand U7882 (N_7882,N_7756,N_7774);
xor U7883 (N_7883,N_7723,N_7833);
nand U7884 (N_7884,N_7817,N_7810);
xnor U7885 (N_7885,N_7700,N_7694);
or U7886 (N_7886,N_7754,N_7829);
nor U7887 (N_7887,N_7780,N_7800);
xor U7888 (N_7888,N_7799,N_7718);
xor U7889 (N_7889,N_7689,N_7775);
xor U7890 (N_7890,N_7706,N_7751);
xor U7891 (N_7891,N_7773,N_7787);
nor U7892 (N_7892,N_7836,N_7701);
nor U7893 (N_7893,N_7795,N_7786);
and U7894 (N_7894,N_7749,N_7715);
nor U7895 (N_7895,N_7729,N_7761);
xor U7896 (N_7896,N_7776,N_7682);
or U7897 (N_7897,N_7753,N_7696);
and U7898 (N_7898,N_7704,N_7764);
nand U7899 (N_7899,N_7794,N_7760);
nor U7900 (N_7900,N_7759,N_7684);
and U7901 (N_7901,N_7783,N_7839);
nor U7902 (N_7902,N_7788,N_7834);
nand U7903 (N_7903,N_7731,N_7687);
nand U7904 (N_7904,N_7710,N_7763);
nor U7905 (N_7905,N_7742,N_7745);
xnor U7906 (N_7906,N_7716,N_7734);
or U7907 (N_7907,N_7744,N_7735);
or U7908 (N_7908,N_7733,N_7736);
nand U7909 (N_7909,N_7814,N_7831);
or U7910 (N_7910,N_7769,N_7820);
and U7911 (N_7911,N_7808,N_7812);
xnor U7912 (N_7912,N_7797,N_7697);
and U7913 (N_7913,N_7828,N_7784);
and U7914 (N_7914,N_7681,N_7691);
and U7915 (N_7915,N_7827,N_7779);
nand U7916 (N_7916,N_7712,N_7738);
and U7917 (N_7917,N_7725,N_7781);
nor U7918 (N_7918,N_7680,N_7768);
or U7919 (N_7919,N_7830,N_7825);
or U7920 (N_7920,N_7684,N_7740);
nand U7921 (N_7921,N_7783,N_7724);
and U7922 (N_7922,N_7681,N_7806);
and U7923 (N_7923,N_7765,N_7759);
nand U7924 (N_7924,N_7736,N_7790);
xnor U7925 (N_7925,N_7811,N_7818);
nand U7926 (N_7926,N_7692,N_7812);
nor U7927 (N_7927,N_7705,N_7831);
nand U7928 (N_7928,N_7684,N_7741);
or U7929 (N_7929,N_7758,N_7747);
nor U7930 (N_7930,N_7744,N_7701);
nand U7931 (N_7931,N_7815,N_7759);
nor U7932 (N_7932,N_7817,N_7783);
nand U7933 (N_7933,N_7806,N_7838);
and U7934 (N_7934,N_7798,N_7749);
nor U7935 (N_7935,N_7681,N_7832);
nor U7936 (N_7936,N_7816,N_7793);
nand U7937 (N_7937,N_7786,N_7723);
nand U7938 (N_7938,N_7690,N_7830);
or U7939 (N_7939,N_7816,N_7763);
xor U7940 (N_7940,N_7715,N_7698);
nor U7941 (N_7941,N_7777,N_7736);
xnor U7942 (N_7942,N_7766,N_7741);
or U7943 (N_7943,N_7763,N_7687);
xnor U7944 (N_7944,N_7698,N_7748);
xor U7945 (N_7945,N_7732,N_7710);
or U7946 (N_7946,N_7698,N_7839);
xor U7947 (N_7947,N_7790,N_7766);
and U7948 (N_7948,N_7729,N_7823);
nand U7949 (N_7949,N_7796,N_7760);
and U7950 (N_7950,N_7836,N_7694);
xor U7951 (N_7951,N_7820,N_7703);
or U7952 (N_7952,N_7787,N_7836);
xor U7953 (N_7953,N_7741,N_7694);
and U7954 (N_7954,N_7732,N_7786);
and U7955 (N_7955,N_7715,N_7707);
and U7956 (N_7956,N_7740,N_7694);
and U7957 (N_7957,N_7767,N_7757);
nand U7958 (N_7958,N_7729,N_7741);
xnor U7959 (N_7959,N_7689,N_7821);
nor U7960 (N_7960,N_7795,N_7812);
nand U7961 (N_7961,N_7707,N_7788);
xnor U7962 (N_7962,N_7771,N_7825);
nand U7963 (N_7963,N_7706,N_7818);
xor U7964 (N_7964,N_7717,N_7684);
nor U7965 (N_7965,N_7729,N_7827);
or U7966 (N_7966,N_7770,N_7709);
nand U7967 (N_7967,N_7769,N_7826);
xnor U7968 (N_7968,N_7818,N_7805);
nor U7969 (N_7969,N_7704,N_7723);
or U7970 (N_7970,N_7783,N_7747);
nor U7971 (N_7971,N_7762,N_7801);
xnor U7972 (N_7972,N_7795,N_7690);
xnor U7973 (N_7973,N_7686,N_7718);
nand U7974 (N_7974,N_7811,N_7801);
or U7975 (N_7975,N_7799,N_7750);
nand U7976 (N_7976,N_7726,N_7766);
or U7977 (N_7977,N_7693,N_7833);
and U7978 (N_7978,N_7831,N_7683);
nand U7979 (N_7979,N_7709,N_7682);
xnor U7980 (N_7980,N_7753,N_7765);
xor U7981 (N_7981,N_7832,N_7773);
nor U7982 (N_7982,N_7776,N_7766);
xnor U7983 (N_7983,N_7799,N_7815);
and U7984 (N_7984,N_7715,N_7768);
and U7985 (N_7985,N_7771,N_7737);
and U7986 (N_7986,N_7680,N_7836);
nor U7987 (N_7987,N_7692,N_7767);
xor U7988 (N_7988,N_7728,N_7735);
or U7989 (N_7989,N_7682,N_7765);
nor U7990 (N_7990,N_7802,N_7738);
or U7991 (N_7991,N_7754,N_7795);
xor U7992 (N_7992,N_7784,N_7802);
nand U7993 (N_7993,N_7697,N_7831);
and U7994 (N_7994,N_7725,N_7827);
nand U7995 (N_7995,N_7815,N_7722);
nor U7996 (N_7996,N_7693,N_7689);
or U7997 (N_7997,N_7823,N_7812);
xor U7998 (N_7998,N_7750,N_7822);
xnor U7999 (N_7999,N_7703,N_7737);
nand U8000 (N_8000,N_7854,N_7849);
and U8001 (N_8001,N_7949,N_7893);
nand U8002 (N_8002,N_7875,N_7887);
nor U8003 (N_8003,N_7963,N_7894);
nor U8004 (N_8004,N_7948,N_7972);
nor U8005 (N_8005,N_7888,N_7996);
or U8006 (N_8006,N_7879,N_7883);
xor U8007 (N_8007,N_7993,N_7873);
nor U8008 (N_8008,N_7923,N_7850);
and U8009 (N_8009,N_7907,N_7899);
nand U8010 (N_8010,N_7847,N_7848);
nand U8011 (N_8011,N_7960,N_7930);
xor U8012 (N_8012,N_7917,N_7976);
nand U8013 (N_8013,N_7920,N_7941);
xor U8014 (N_8014,N_7871,N_7898);
and U8015 (N_8015,N_7856,N_7981);
xnor U8016 (N_8016,N_7989,N_7927);
or U8017 (N_8017,N_7896,N_7924);
xor U8018 (N_8018,N_7866,N_7890);
xor U8019 (N_8019,N_7971,N_7946);
nand U8020 (N_8020,N_7918,N_7880);
or U8021 (N_8021,N_7964,N_7953);
or U8022 (N_8022,N_7882,N_7936);
nand U8023 (N_8023,N_7852,N_7841);
or U8024 (N_8024,N_7878,N_7952);
nor U8025 (N_8025,N_7905,N_7954);
xor U8026 (N_8026,N_7915,N_7886);
nor U8027 (N_8027,N_7877,N_7855);
or U8028 (N_8028,N_7922,N_7900);
xnor U8029 (N_8029,N_7947,N_7874);
nor U8030 (N_8030,N_7925,N_7932);
xor U8031 (N_8031,N_7926,N_7982);
nor U8032 (N_8032,N_7944,N_7913);
or U8033 (N_8033,N_7974,N_7869);
and U8034 (N_8034,N_7906,N_7979);
or U8035 (N_8035,N_7966,N_7951);
and U8036 (N_8036,N_7889,N_7937);
and U8037 (N_8037,N_7994,N_7990);
and U8038 (N_8038,N_7921,N_7903);
nand U8039 (N_8039,N_7844,N_7911);
xnor U8040 (N_8040,N_7934,N_7929);
xnor U8041 (N_8041,N_7998,N_7985);
xor U8042 (N_8042,N_7851,N_7916);
xnor U8043 (N_8043,N_7965,N_7992);
xor U8044 (N_8044,N_7955,N_7864);
and U8045 (N_8045,N_7958,N_7959);
or U8046 (N_8046,N_7872,N_7909);
and U8047 (N_8047,N_7912,N_7988);
xor U8048 (N_8048,N_7862,N_7970);
xor U8049 (N_8049,N_7861,N_7858);
nor U8050 (N_8050,N_7931,N_7868);
xor U8051 (N_8051,N_7968,N_7956);
nor U8052 (N_8052,N_7940,N_7863);
xor U8053 (N_8053,N_7857,N_7902);
nor U8054 (N_8054,N_7867,N_7939);
and U8055 (N_8055,N_7840,N_7876);
nand U8056 (N_8056,N_7870,N_7980);
nand U8057 (N_8057,N_7919,N_7950);
nor U8058 (N_8058,N_7859,N_7991);
nand U8059 (N_8059,N_7975,N_7967);
xor U8060 (N_8060,N_7978,N_7997);
or U8061 (N_8061,N_7995,N_7933);
and U8062 (N_8062,N_7938,N_7910);
nand U8063 (N_8063,N_7908,N_7842);
and U8064 (N_8064,N_7891,N_7860);
xnor U8065 (N_8065,N_7904,N_7986);
and U8066 (N_8066,N_7892,N_7957);
and U8067 (N_8067,N_7942,N_7987);
nand U8068 (N_8068,N_7984,N_7914);
and U8069 (N_8069,N_7961,N_7881);
nand U8070 (N_8070,N_7853,N_7865);
xnor U8071 (N_8071,N_7846,N_7977);
or U8072 (N_8072,N_7973,N_7884);
nor U8073 (N_8073,N_7983,N_7945);
and U8074 (N_8074,N_7843,N_7895);
xnor U8075 (N_8075,N_7935,N_7943);
or U8076 (N_8076,N_7845,N_7969);
and U8077 (N_8077,N_7999,N_7901);
nor U8078 (N_8078,N_7962,N_7885);
or U8079 (N_8079,N_7928,N_7897);
or U8080 (N_8080,N_7865,N_7926);
nor U8081 (N_8081,N_7925,N_7943);
nor U8082 (N_8082,N_7860,N_7843);
nand U8083 (N_8083,N_7932,N_7965);
xor U8084 (N_8084,N_7883,N_7843);
xnor U8085 (N_8085,N_7896,N_7953);
or U8086 (N_8086,N_7846,N_7990);
or U8087 (N_8087,N_7905,N_7961);
and U8088 (N_8088,N_7964,N_7844);
nand U8089 (N_8089,N_7974,N_7886);
nand U8090 (N_8090,N_7919,N_7974);
nor U8091 (N_8091,N_7873,N_7991);
nand U8092 (N_8092,N_7878,N_7886);
xor U8093 (N_8093,N_7930,N_7967);
and U8094 (N_8094,N_7842,N_7864);
nand U8095 (N_8095,N_7978,N_7856);
nand U8096 (N_8096,N_7883,N_7953);
or U8097 (N_8097,N_7992,N_7949);
xnor U8098 (N_8098,N_7882,N_7875);
and U8099 (N_8099,N_7969,N_7943);
and U8100 (N_8100,N_7842,N_7954);
and U8101 (N_8101,N_7912,N_7946);
nor U8102 (N_8102,N_7991,N_7922);
nand U8103 (N_8103,N_7897,N_7912);
or U8104 (N_8104,N_7959,N_7907);
and U8105 (N_8105,N_7938,N_7922);
nor U8106 (N_8106,N_7953,N_7975);
xor U8107 (N_8107,N_7847,N_7922);
and U8108 (N_8108,N_7909,N_7869);
nor U8109 (N_8109,N_7860,N_7991);
nor U8110 (N_8110,N_7982,N_7865);
and U8111 (N_8111,N_7886,N_7981);
nand U8112 (N_8112,N_7860,N_7911);
and U8113 (N_8113,N_7966,N_7948);
nor U8114 (N_8114,N_7912,N_7879);
nand U8115 (N_8115,N_7976,N_7922);
nand U8116 (N_8116,N_7919,N_7866);
nand U8117 (N_8117,N_7928,N_7841);
and U8118 (N_8118,N_7897,N_7923);
and U8119 (N_8119,N_7998,N_7886);
or U8120 (N_8120,N_7978,N_7910);
or U8121 (N_8121,N_7935,N_7870);
nand U8122 (N_8122,N_7985,N_7886);
and U8123 (N_8123,N_7850,N_7981);
xnor U8124 (N_8124,N_7890,N_7984);
nor U8125 (N_8125,N_7917,N_7857);
xor U8126 (N_8126,N_7980,N_7967);
nand U8127 (N_8127,N_7866,N_7885);
nand U8128 (N_8128,N_7849,N_7907);
and U8129 (N_8129,N_7975,N_7922);
and U8130 (N_8130,N_7935,N_7876);
nor U8131 (N_8131,N_7899,N_7900);
or U8132 (N_8132,N_7889,N_7945);
nand U8133 (N_8133,N_7924,N_7855);
nor U8134 (N_8134,N_7960,N_7997);
xor U8135 (N_8135,N_7860,N_7888);
or U8136 (N_8136,N_7870,N_7982);
nand U8137 (N_8137,N_7978,N_7952);
nand U8138 (N_8138,N_7884,N_7980);
nor U8139 (N_8139,N_7984,N_7952);
xor U8140 (N_8140,N_7954,N_7894);
nand U8141 (N_8141,N_7929,N_7895);
nor U8142 (N_8142,N_7977,N_7998);
and U8143 (N_8143,N_7935,N_7844);
or U8144 (N_8144,N_7930,N_7918);
nor U8145 (N_8145,N_7888,N_7862);
or U8146 (N_8146,N_7942,N_7885);
or U8147 (N_8147,N_7960,N_7968);
or U8148 (N_8148,N_7918,N_7999);
or U8149 (N_8149,N_7964,N_7960);
xnor U8150 (N_8150,N_7974,N_7962);
xor U8151 (N_8151,N_7934,N_7943);
nor U8152 (N_8152,N_7850,N_7993);
and U8153 (N_8153,N_7940,N_7948);
or U8154 (N_8154,N_7856,N_7947);
nor U8155 (N_8155,N_7964,N_7993);
nor U8156 (N_8156,N_7944,N_7981);
xnor U8157 (N_8157,N_7858,N_7857);
xnor U8158 (N_8158,N_7877,N_7996);
or U8159 (N_8159,N_7870,N_7948);
nor U8160 (N_8160,N_8069,N_8043);
nor U8161 (N_8161,N_8130,N_8106);
xor U8162 (N_8162,N_8143,N_8035);
nand U8163 (N_8163,N_8118,N_8009);
nor U8164 (N_8164,N_8025,N_8121);
or U8165 (N_8165,N_8045,N_8087);
xnor U8166 (N_8166,N_8018,N_8100);
or U8167 (N_8167,N_8063,N_8010);
and U8168 (N_8168,N_8111,N_8086);
nor U8169 (N_8169,N_8078,N_8131);
xnor U8170 (N_8170,N_8117,N_8090);
nor U8171 (N_8171,N_8155,N_8052);
and U8172 (N_8172,N_8079,N_8049);
or U8173 (N_8173,N_8039,N_8098);
nand U8174 (N_8174,N_8076,N_8151);
xnor U8175 (N_8175,N_8119,N_8051);
xnor U8176 (N_8176,N_8032,N_8073);
xor U8177 (N_8177,N_8031,N_8152);
xor U8178 (N_8178,N_8089,N_8081);
nor U8179 (N_8179,N_8096,N_8147);
and U8180 (N_8180,N_8088,N_8122);
and U8181 (N_8181,N_8065,N_8114);
nand U8182 (N_8182,N_8099,N_8072);
xor U8183 (N_8183,N_8110,N_8084);
nand U8184 (N_8184,N_8091,N_8128);
and U8185 (N_8185,N_8064,N_8029);
and U8186 (N_8186,N_8056,N_8034);
or U8187 (N_8187,N_8095,N_8006);
and U8188 (N_8188,N_8129,N_8156);
and U8189 (N_8189,N_8127,N_8037);
nor U8190 (N_8190,N_8120,N_8158);
xnor U8191 (N_8191,N_8001,N_8014);
nand U8192 (N_8192,N_8057,N_8137);
and U8193 (N_8193,N_8139,N_8093);
nor U8194 (N_8194,N_8007,N_8062);
and U8195 (N_8195,N_8135,N_8005);
nor U8196 (N_8196,N_8144,N_8027);
or U8197 (N_8197,N_8003,N_8134);
nor U8198 (N_8198,N_8109,N_8150);
nor U8199 (N_8199,N_8132,N_8146);
nor U8200 (N_8200,N_8097,N_8116);
or U8201 (N_8201,N_8080,N_8000);
nand U8202 (N_8202,N_8055,N_8105);
nand U8203 (N_8203,N_8040,N_8094);
nor U8204 (N_8204,N_8024,N_8054);
xnor U8205 (N_8205,N_8153,N_8145);
nor U8206 (N_8206,N_8019,N_8041);
and U8207 (N_8207,N_8157,N_8103);
and U8208 (N_8208,N_8036,N_8101);
or U8209 (N_8209,N_8112,N_8070);
nand U8210 (N_8210,N_8044,N_8074);
xnor U8211 (N_8211,N_8108,N_8060);
or U8212 (N_8212,N_8021,N_8004);
xor U8213 (N_8213,N_8113,N_8059);
nor U8214 (N_8214,N_8008,N_8015);
and U8215 (N_8215,N_8107,N_8142);
nand U8216 (N_8216,N_8083,N_8159);
or U8217 (N_8217,N_8071,N_8038);
and U8218 (N_8218,N_8066,N_8077);
nor U8219 (N_8219,N_8046,N_8012);
or U8220 (N_8220,N_8141,N_8033);
or U8221 (N_8221,N_8082,N_8154);
or U8222 (N_8222,N_8042,N_8017);
xnor U8223 (N_8223,N_8067,N_8020);
xor U8224 (N_8224,N_8148,N_8126);
nand U8225 (N_8225,N_8092,N_8016);
xnor U8226 (N_8226,N_8068,N_8053);
or U8227 (N_8227,N_8133,N_8022);
or U8228 (N_8228,N_8104,N_8123);
nor U8229 (N_8229,N_8026,N_8047);
or U8230 (N_8230,N_8050,N_8136);
nor U8231 (N_8231,N_8058,N_8028);
or U8232 (N_8232,N_8140,N_8013);
nand U8233 (N_8233,N_8125,N_8030);
nand U8234 (N_8234,N_8002,N_8023);
nor U8235 (N_8235,N_8048,N_8124);
nor U8236 (N_8236,N_8102,N_8075);
nand U8237 (N_8237,N_8085,N_8061);
or U8238 (N_8238,N_8138,N_8011);
nand U8239 (N_8239,N_8149,N_8115);
nor U8240 (N_8240,N_8079,N_8035);
xnor U8241 (N_8241,N_8004,N_8090);
nand U8242 (N_8242,N_8013,N_8149);
or U8243 (N_8243,N_8082,N_8030);
nor U8244 (N_8244,N_8140,N_8088);
nand U8245 (N_8245,N_8126,N_8089);
xnor U8246 (N_8246,N_8034,N_8032);
xnor U8247 (N_8247,N_8008,N_8148);
xor U8248 (N_8248,N_8059,N_8130);
or U8249 (N_8249,N_8064,N_8105);
xnor U8250 (N_8250,N_8095,N_8003);
and U8251 (N_8251,N_8023,N_8105);
xor U8252 (N_8252,N_8072,N_8103);
xnor U8253 (N_8253,N_8128,N_8013);
nand U8254 (N_8254,N_8114,N_8030);
and U8255 (N_8255,N_8057,N_8131);
xnor U8256 (N_8256,N_8141,N_8120);
and U8257 (N_8257,N_8012,N_8060);
or U8258 (N_8258,N_8114,N_8100);
and U8259 (N_8259,N_8100,N_8103);
and U8260 (N_8260,N_8022,N_8156);
xor U8261 (N_8261,N_8061,N_8092);
nor U8262 (N_8262,N_8125,N_8041);
xnor U8263 (N_8263,N_8003,N_8060);
nand U8264 (N_8264,N_8139,N_8077);
nor U8265 (N_8265,N_8128,N_8014);
and U8266 (N_8266,N_8025,N_8141);
nand U8267 (N_8267,N_8131,N_8128);
and U8268 (N_8268,N_8019,N_8070);
and U8269 (N_8269,N_8059,N_8088);
nor U8270 (N_8270,N_8090,N_8099);
nor U8271 (N_8271,N_8016,N_8063);
nand U8272 (N_8272,N_8023,N_8016);
xor U8273 (N_8273,N_8076,N_8018);
and U8274 (N_8274,N_8090,N_8096);
nor U8275 (N_8275,N_8007,N_8001);
xnor U8276 (N_8276,N_8129,N_8013);
nand U8277 (N_8277,N_8136,N_8065);
nor U8278 (N_8278,N_8096,N_8119);
xor U8279 (N_8279,N_8049,N_8085);
nor U8280 (N_8280,N_8033,N_8022);
and U8281 (N_8281,N_8017,N_8143);
nor U8282 (N_8282,N_8153,N_8022);
and U8283 (N_8283,N_8156,N_8079);
xor U8284 (N_8284,N_8007,N_8125);
xor U8285 (N_8285,N_8117,N_8029);
nand U8286 (N_8286,N_8012,N_8015);
nor U8287 (N_8287,N_8049,N_8117);
nand U8288 (N_8288,N_8021,N_8055);
nor U8289 (N_8289,N_8079,N_8102);
nor U8290 (N_8290,N_8112,N_8097);
nand U8291 (N_8291,N_8076,N_8108);
and U8292 (N_8292,N_8014,N_8022);
nand U8293 (N_8293,N_8159,N_8071);
and U8294 (N_8294,N_8035,N_8109);
xor U8295 (N_8295,N_8154,N_8002);
and U8296 (N_8296,N_8010,N_8050);
and U8297 (N_8297,N_8137,N_8116);
nor U8298 (N_8298,N_8093,N_8081);
or U8299 (N_8299,N_8148,N_8100);
xnor U8300 (N_8300,N_8123,N_8074);
or U8301 (N_8301,N_8144,N_8152);
xnor U8302 (N_8302,N_8072,N_8081);
nor U8303 (N_8303,N_8152,N_8018);
and U8304 (N_8304,N_8088,N_8023);
nor U8305 (N_8305,N_8057,N_8000);
nand U8306 (N_8306,N_8142,N_8058);
and U8307 (N_8307,N_8028,N_8130);
and U8308 (N_8308,N_8069,N_8026);
nor U8309 (N_8309,N_8068,N_8049);
nor U8310 (N_8310,N_8111,N_8031);
or U8311 (N_8311,N_8038,N_8023);
nor U8312 (N_8312,N_8136,N_8080);
nand U8313 (N_8313,N_8034,N_8053);
xnor U8314 (N_8314,N_8001,N_8000);
xnor U8315 (N_8315,N_8003,N_8051);
and U8316 (N_8316,N_8125,N_8029);
and U8317 (N_8317,N_8058,N_8104);
nor U8318 (N_8318,N_8155,N_8094);
nand U8319 (N_8319,N_8128,N_8079);
or U8320 (N_8320,N_8318,N_8262);
or U8321 (N_8321,N_8298,N_8223);
nor U8322 (N_8322,N_8186,N_8273);
xor U8323 (N_8323,N_8279,N_8270);
or U8324 (N_8324,N_8231,N_8218);
or U8325 (N_8325,N_8203,N_8288);
nand U8326 (N_8326,N_8167,N_8233);
nand U8327 (N_8327,N_8302,N_8198);
nand U8328 (N_8328,N_8282,N_8224);
and U8329 (N_8329,N_8217,N_8205);
and U8330 (N_8330,N_8236,N_8283);
xor U8331 (N_8331,N_8240,N_8162);
or U8332 (N_8332,N_8238,N_8177);
or U8333 (N_8333,N_8163,N_8164);
nand U8334 (N_8334,N_8274,N_8160);
nand U8335 (N_8335,N_8253,N_8241);
xnor U8336 (N_8336,N_8250,N_8249);
and U8337 (N_8337,N_8245,N_8277);
nor U8338 (N_8338,N_8263,N_8285);
nand U8339 (N_8339,N_8174,N_8182);
nand U8340 (N_8340,N_8294,N_8210);
or U8341 (N_8341,N_8313,N_8222);
or U8342 (N_8342,N_8161,N_8275);
and U8343 (N_8343,N_8171,N_8190);
and U8344 (N_8344,N_8196,N_8309);
xnor U8345 (N_8345,N_8312,N_8214);
nor U8346 (N_8346,N_8310,N_8227);
and U8347 (N_8347,N_8244,N_8185);
or U8348 (N_8348,N_8281,N_8200);
xor U8349 (N_8349,N_8254,N_8181);
nand U8350 (N_8350,N_8195,N_8306);
xor U8351 (N_8351,N_8170,N_8204);
nand U8352 (N_8352,N_8258,N_8246);
or U8353 (N_8353,N_8303,N_8284);
xnor U8354 (N_8354,N_8219,N_8266);
nor U8355 (N_8355,N_8191,N_8278);
nand U8356 (N_8356,N_8307,N_8280);
nand U8357 (N_8357,N_8319,N_8269);
or U8358 (N_8358,N_8296,N_8297);
xor U8359 (N_8359,N_8315,N_8248);
xor U8360 (N_8360,N_8252,N_8187);
or U8361 (N_8361,N_8168,N_8234);
nor U8362 (N_8362,N_8211,N_8251);
and U8363 (N_8363,N_8301,N_8220);
nand U8364 (N_8364,N_8267,N_8208);
and U8365 (N_8365,N_8299,N_8265);
xor U8366 (N_8366,N_8256,N_8188);
or U8367 (N_8367,N_8264,N_8165);
xor U8368 (N_8368,N_8289,N_8247);
or U8369 (N_8369,N_8268,N_8286);
xor U8370 (N_8370,N_8260,N_8276);
nand U8371 (N_8371,N_8175,N_8178);
and U8372 (N_8372,N_8225,N_8295);
xor U8373 (N_8373,N_8189,N_8308);
and U8374 (N_8374,N_8184,N_8305);
or U8375 (N_8375,N_8237,N_8176);
and U8376 (N_8376,N_8179,N_8215);
nor U8377 (N_8377,N_8207,N_8293);
nand U8378 (N_8378,N_8194,N_8173);
xor U8379 (N_8379,N_8202,N_8199);
nor U8380 (N_8380,N_8197,N_8201);
nand U8381 (N_8381,N_8180,N_8257);
nor U8382 (N_8382,N_8316,N_8213);
and U8383 (N_8383,N_8287,N_8261);
or U8384 (N_8384,N_8239,N_8235);
xnor U8385 (N_8385,N_8272,N_8216);
xnor U8386 (N_8386,N_8311,N_8172);
or U8387 (N_8387,N_8300,N_8291);
and U8388 (N_8388,N_8314,N_8221);
nand U8389 (N_8389,N_8209,N_8259);
nor U8390 (N_8390,N_8193,N_8229);
nand U8391 (N_8391,N_8242,N_8255);
and U8392 (N_8392,N_8292,N_8232);
xor U8393 (N_8393,N_8226,N_8228);
or U8394 (N_8394,N_8212,N_8243);
nand U8395 (N_8395,N_8290,N_8183);
and U8396 (N_8396,N_8304,N_8206);
nor U8397 (N_8397,N_8271,N_8169);
nand U8398 (N_8398,N_8166,N_8230);
nand U8399 (N_8399,N_8317,N_8192);
nor U8400 (N_8400,N_8288,N_8275);
nor U8401 (N_8401,N_8298,N_8266);
nand U8402 (N_8402,N_8231,N_8316);
nand U8403 (N_8403,N_8300,N_8268);
xor U8404 (N_8404,N_8260,N_8169);
and U8405 (N_8405,N_8256,N_8282);
or U8406 (N_8406,N_8174,N_8178);
or U8407 (N_8407,N_8226,N_8208);
nor U8408 (N_8408,N_8230,N_8265);
or U8409 (N_8409,N_8255,N_8297);
and U8410 (N_8410,N_8211,N_8169);
nand U8411 (N_8411,N_8265,N_8164);
nor U8412 (N_8412,N_8222,N_8293);
nand U8413 (N_8413,N_8309,N_8264);
or U8414 (N_8414,N_8175,N_8308);
nand U8415 (N_8415,N_8187,N_8306);
nand U8416 (N_8416,N_8184,N_8317);
and U8417 (N_8417,N_8222,N_8289);
nor U8418 (N_8418,N_8289,N_8298);
xnor U8419 (N_8419,N_8314,N_8168);
and U8420 (N_8420,N_8252,N_8295);
and U8421 (N_8421,N_8167,N_8246);
nor U8422 (N_8422,N_8223,N_8273);
xor U8423 (N_8423,N_8240,N_8288);
xnor U8424 (N_8424,N_8205,N_8194);
xnor U8425 (N_8425,N_8222,N_8290);
or U8426 (N_8426,N_8206,N_8199);
nand U8427 (N_8427,N_8172,N_8211);
and U8428 (N_8428,N_8191,N_8215);
xor U8429 (N_8429,N_8170,N_8199);
or U8430 (N_8430,N_8238,N_8292);
xnor U8431 (N_8431,N_8256,N_8248);
xnor U8432 (N_8432,N_8314,N_8258);
and U8433 (N_8433,N_8237,N_8296);
nor U8434 (N_8434,N_8263,N_8316);
nand U8435 (N_8435,N_8272,N_8230);
xnor U8436 (N_8436,N_8317,N_8298);
and U8437 (N_8437,N_8203,N_8307);
or U8438 (N_8438,N_8255,N_8268);
nand U8439 (N_8439,N_8231,N_8264);
or U8440 (N_8440,N_8264,N_8294);
or U8441 (N_8441,N_8305,N_8234);
nor U8442 (N_8442,N_8297,N_8286);
nand U8443 (N_8443,N_8262,N_8230);
xnor U8444 (N_8444,N_8262,N_8261);
and U8445 (N_8445,N_8301,N_8212);
xnor U8446 (N_8446,N_8257,N_8297);
and U8447 (N_8447,N_8304,N_8248);
or U8448 (N_8448,N_8191,N_8295);
or U8449 (N_8449,N_8255,N_8276);
or U8450 (N_8450,N_8313,N_8294);
and U8451 (N_8451,N_8206,N_8314);
nand U8452 (N_8452,N_8245,N_8247);
nor U8453 (N_8453,N_8289,N_8295);
and U8454 (N_8454,N_8184,N_8306);
xor U8455 (N_8455,N_8290,N_8200);
and U8456 (N_8456,N_8250,N_8184);
nand U8457 (N_8457,N_8261,N_8296);
xnor U8458 (N_8458,N_8190,N_8270);
nand U8459 (N_8459,N_8164,N_8230);
nor U8460 (N_8460,N_8227,N_8251);
nand U8461 (N_8461,N_8194,N_8247);
nor U8462 (N_8462,N_8170,N_8300);
xor U8463 (N_8463,N_8259,N_8216);
or U8464 (N_8464,N_8167,N_8211);
xor U8465 (N_8465,N_8257,N_8193);
nand U8466 (N_8466,N_8167,N_8316);
nand U8467 (N_8467,N_8235,N_8165);
and U8468 (N_8468,N_8307,N_8231);
or U8469 (N_8469,N_8293,N_8221);
xor U8470 (N_8470,N_8204,N_8193);
and U8471 (N_8471,N_8271,N_8243);
or U8472 (N_8472,N_8220,N_8298);
nor U8473 (N_8473,N_8279,N_8278);
xor U8474 (N_8474,N_8222,N_8311);
and U8475 (N_8475,N_8255,N_8265);
or U8476 (N_8476,N_8245,N_8313);
and U8477 (N_8477,N_8210,N_8232);
nand U8478 (N_8478,N_8311,N_8264);
nor U8479 (N_8479,N_8278,N_8262);
nor U8480 (N_8480,N_8426,N_8478);
xor U8481 (N_8481,N_8385,N_8394);
or U8482 (N_8482,N_8373,N_8463);
and U8483 (N_8483,N_8379,N_8449);
nand U8484 (N_8484,N_8432,N_8436);
nor U8485 (N_8485,N_8351,N_8349);
xor U8486 (N_8486,N_8337,N_8418);
and U8487 (N_8487,N_8381,N_8365);
nor U8488 (N_8488,N_8361,N_8444);
xnor U8489 (N_8489,N_8479,N_8459);
nor U8490 (N_8490,N_8421,N_8399);
nand U8491 (N_8491,N_8362,N_8442);
nand U8492 (N_8492,N_8414,N_8419);
nand U8493 (N_8493,N_8453,N_8359);
xor U8494 (N_8494,N_8409,N_8375);
or U8495 (N_8495,N_8398,N_8346);
nand U8496 (N_8496,N_8456,N_8323);
or U8497 (N_8497,N_8383,N_8446);
xor U8498 (N_8498,N_8338,N_8401);
or U8499 (N_8499,N_8376,N_8367);
nand U8500 (N_8500,N_8455,N_8356);
or U8501 (N_8501,N_8405,N_8335);
nand U8502 (N_8502,N_8352,N_8371);
and U8503 (N_8503,N_8331,N_8425);
xnor U8504 (N_8504,N_8332,N_8407);
xnor U8505 (N_8505,N_8474,N_8420);
nand U8506 (N_8506,N_8438,N_8393);
nor U8507 (N_8507,N_8475,N_8465);
nand U8508 (N_8508,N_8357,N_8358);
and U8509 (N_8509,N_8450,N_8427);
xor U8510 (N_8510,N_8325,N_8443);
xor U8511 (N_8511,N_8400,N_8368);
xnor U8512 (N_8512,N_8329,N_8433);
and U8513 (N_8513,N_8363,N_8350);
and U8514 (N_8514,N_8452,N_8347);
nand U8515 (N_8515,N_8328,N_8431);
nand U8516 (N_8516,N_8406,N_8374);
or U8517 (N_8517,N_8339,N_8461);
nand U8518 (N_8518,N_8330,N_8320);
nor U8519 (N_8519,N_8360,N_8334);
nor U8520 (N_8520,N_8324,N_8454);
and U8521 (N_8521,N_8377,N_8370);
and U8522 (N_8522,N_8355,N_8429);
nor U8523 (N_8523,N_8457,N_8411);
or U8524 (N_8524,N_8413,N_8340);
and U8525 (N_8525,N_8326,N_8447);
xnor U8526 (N_8526,N_8392,N_8471);
or U8527 (N_8527,N_8412,N_8386);
and U8528 (N_8528,N_8364,N_8333);
nor U8529 (N_8529,N_8458,N_8430);
nor U8530 (N_8530,N_8353,N_8342);
xor U8531 (N_8531,N_8397,N_8372);
nor U8532 (N_8532,N_8391,N_8462);
nor U8533 (N_8533,N_8466,N_8387);
xor U8534 (N_8534,N_8434,N_8423);
or U8535 (N_8535,N_8467,N_8344);
nor U8536 (N_8536,N_8380,N_8468);
xnor U8537 (N_8537,N_8476,N_8404);
xor U8538 (N_8538,N_8396,N_8470);
nor U8539 (N_8539,N_8321,N_8322);
xnor U8540 (N_8540,N_8451,N_8384);
nor U8541 (N_8541,N_8435,N_8415);
and U8542 (N_8542,N_8382,N_8390);
or U8543 (N_8543,N_8440,N_8477);
xnor U8544 (N_8544,N_8408,N_8460);
nand U8545 (N_8545,N_8327,N_8366);
or U8546 (N_8546,N_8341,N_8369);
nand U8547 (N_8547,N_8437,N_8410);
nor U8548 (N_8548,N_8416,N_8417);
or U8549 (N_8549,N_8336,N_8469);
nor U8550 (N_8550,N_8428,N_8424);
xnor U8551 (N_8551,N_8348,N_8395);
xor U8552 (N_8552,N_8448,N_8345);
nand U8553 (N_8553,N_8389,N_8388);
and U8554 (N_8554,N_8464,N_8343);
nor U8555 (N_8555,N_8402,N_8472);
nor U8556 (N_8556,N_8378,N_8441);
or U8557 (N_8557,N_8403,N_8439);
nand U8558 (N_8558,N_8445,N_8473);
nor U8559 (N_8559,N_8354,N_8422);
nand U8560 (N_8560,N_8364,N_8346);
nor U8561 (N_8561,N_8322,N_8479);
xor U8562 (N_8562,N_8472,N_8380);
and U8563 (N_8563,N_8358,N_8413);
nand U8564 (N_8564,N_8468,N_8473);
xnor U8565 (N_8565,N_8387,N_8392);
nand U8566 (N_8566,N_8333,N_8471);
or U8567 (N_8567,N_8460,N_8396);
xnor U8568 (N_8568,N_8451,N_8449);
nor U8569 (N_8569,N_8422,N_8449);
nand U8570 (N_8570,N_8344,N_8359);
nand U8571 (N_8571,N_8384,N_8403);
and U8572 (N_8572,N_8337,N_8399);
xnor U8573 (N_8573,N_8418,N_8363);
nor U8574 (N_8574,N_8392,N_8391);
or U8575 (N_8575,N_8379,N_8368);
nand U8576 (N_8576,N_8456,N_8362);
nor U8577 (N_8577,N_8375,N_8425);
nand U8578 (N_8578,N_8420,N_8458);
nor U8579 (N_8579,N_8451,N_8358);
and U8580 (N_8580,N_8412,N_8402);
or U8581 (N_8581,N_8465,N_8321);
and U8582 (N_8582,N_8330,N_8416);
nor U8583 (N_8583,N_8407,N_8426);
or U8584 (N_8584,N_8325,N_8338);
and U8585 (N_8585,N_8402,N_8466);
or U8586 (N_8586,N_8393,N_8435);
xor U8587 (N_8587,N_8461,N_8383);
nor U8588 (N_8588,N_8410,N_8374);
nor U8589 (N_8589,N_8338,N_8425);
or U8590 (N_8590,N_8475,N_8374);
or U8591 (N_8591,N_8385,N_8456);
xor U8592 (N_8592,N_8463,N_8358);
and U8593 (N_8593,N_8362,N_8469);
nor U8594 (N_8594,N_8436,N_8440);
or U8595 (N_8595,N_8425,N_8359);
nand U8596 (N_8596,N_8356,N_8342);
nor U8597 (N_8597,N_8465,N_8356);
nand U8598 (N_8598,N_8452,N_8376);
nand U8599 (N_8599,N_8471,N_8475);
xor U8600 (N_8600,N_8477,N_8429);
and U8601 (N_8601,N_8467,N_8331);
or U8602 (N_8602,N_8368,N_8377);
or U8603 (N_8603,N_8412,N_8329);
or U8604 (N_8604,N_8349,N_8411);
nor U8605 (N_8605,N_8332,N_8360);
nor U8606 (N_8606,N_8382,N_8328);
or U8607 (N_8607,N_8451,N_8416);
or U8608 (N_8608,N_8428,N_8347);
and U8609 (N_8609,N_8417,N_8414);
xnor U8610 (N_8610,N_8396,N_8419);
nand U8611 (N_8611,N_8448,N_8412);
and U8612 (N_8612,N_8424,N_8453);
xor U8613 (N_8613,N_8402,N_8403);
xor U8614 (N_8614,N_8456,N_8359);
xnor U8615 (N_8615,N_8471,N_8468);
nor U8616 (N_8616,N_8411,N_8470);
and U8617 (N_8617,N_8439,N_8436);
and U8618 (N_8618,N_8397,N_8362);
xnor U8619 (N_8619,N_8385,N_8340);
nor U8620 (N_8620,N_8383,N_8439);
nor U8621 (N_8621,N_8398,N_8450);
xnor U8622 (N_8622,N_8361,N_8363);
nand U8623 (N_8623,N_8451,N_8459);
or U8624 (N_8624,N_8390,N_8369);
or U8625 (N_8625,N_8418,N_8476);
or U8626 (N_8626,N_8453,N_8348);
xnor U8627 (N_8627,N_8326,N_8400);
nand U8628 (N_8628,N_8365,N_8415);
and U8629 (N_8629,N_8458,N_8393);
nor U8630 (N_8630,N_8444,N_8457);
or U8631 (N_8631,N_8330,N_8406);
or U8632 (N_8632,N_8426,N_8368);
and U8633 (N_8633,N_8355,N_8333);
xnor U8634 (N_8634,N_8459,N_8377);
nor U8635 (N_8635,N_8350,N_8418);
nand U8636 (N_8636,N_8448,N_8464);
or U8637 (N_8637,N_8413,N_8371);
nand U8638 (N_8638,N_8322,N_8382);
and U8639 (N_8639,N_8384,N_8396);
or U8640 (N_8640,N_8590,N_8625);
nand U8641 (N_8641,N_8579,N_8636);
nand U8642 (N_8642,N_8598,N_8480);
nand U8643 (N_8643,N_8549,N_8530);
or U8644 (N_8644,N_8639,N_8504);
nor U8645 (N_8645,N_8554,N_8518);
or U8646 (N_8646,N_8584,N_8546);
xor U8647 (N_8647,N_8575,N_8487);
nand U8648 (N_8648,N_8519,N_8565);
nand U8649 (N_8649,N_8553,N_8631);
xor U8650 (N_8650,N_8500,N_8588);
xnor U8651 (N_8651,N_8482,N_8545);
and U8652 (N_8652,N_8562,N_8527);
nor U8653 (N_8653,N_8503,N_8592);
nor U8654 (N_8654,N_8566,N_8568);
nand U8655 (N_8655,N_8548,N_8542);
nand U8656 (N_8656,N_8596,N_8629);
or U8657 (N_8657,N_8624,N_8564);
and U8658 (N_8658,N_8623,N_8573);
nor U8659 (N_8659,N_8593,N_8638);
or U8660 (N_8660,N_8589,N_8616);
and U8661 (N_8661,N_8614,N_8569);
xnor U8662 (N_8662,N_8601,N_8594);
and U8663 (N_8663,N_8507,N_8634);
nor U8664 (N_8664,N_8541,N_8617);
and U8665 (N_8665,N_8502,N_8612);
or U8666 (N_8666,N_8574,N_8558);
nand U8667 (N_8667,N_8511,N_8633);
and U8668 (N_8668,N_8556,N_8497);
nor U8669 (N_8669,N_8505,N_8595);
nand U8670 (N_8670,N_8615,N_8628);
and U8671 (N_8671,N_8627,N_8637);
nor U8672 (N_8672,N_8534,N_8524);
nand U8673 (N_8673,N_8525,N_8585);
xnor U8674 (N_8674,N_8533,N_8635);
nand U8675 (N_8675,N_8512,N_8516);
xnor U8676 (N_8676,N_8608,N_8611);
xor U8677 (N_8677,N_8539,N_8528);
nor U8678 (N_8678,N_8515,N_8621);
xnor U8679 (N_8679,N_8485,N_8506);
xor U8680 (N_8680,N_8537,N_8560);
or U8681 (N_8681,N_8600,N_8520);
and U8682 (N_8682,N_8561,N_8559);
nor U8683 (N_8683,N_8572,N_8510);
nor U8684 (N_8684,N_8587,N_8578);
nor U8685 (N_8685,N_8547,N_8603);
nand U8686 (N_8686,N_8540,N_8495);
and U8687 (N_8687,N_8609,N_8514);
xnor U8688 (N_8688,N_8491,N_8498);
xor U8689 (N_8689,N_8552,N_8490);
nand U8690 (N_8690,N_8576,N_8481);
or U8691 (N_8691,N_8582,N_8496);
xnor U8692 (N_8692,N_8632,N_8580);
xor U8693 (N_8693,N_8622,N_8494);
and U8694 (N_8694,N_8581,N_8529);
xnor U8695 (N_8695,N_8499,N_8610);
xor U8696 (N_8696,N_8523,N_8489);
nor U8697 (N_8697,N_8535,N_8488);
nand U8698 (N_8698,N_8483,N_8618);
xnor U8699 (N_8699,N_8538,N_8619);
and U8700 (N_8700,N_8521,N_8630);
nand U8701 (N_8701,N_8571,N_8577);
and U8702 (N_8702,N_8551,N_8620);
and U8703 (N_8703,N_8509,N_8599);
and U8704 (N_8704,N_8567,N_8602);
nand U8705 (N_8705,N_8626,N_8604);
nand U8706 (N_8706,N_8517,N_8606);
and U8707 (N_8707,N_8597,N_8563);
or U8708 (N_8708,N_8532,N_8531);
nand U8709 (N_8709,N_8508,N_8484);
xnor U8710 (N_8710,N_8513,N_8522);
xnor U8711 (N_8711,N_8526,N_8555);
or U8712 (N_8712,N_8501,N_8543);
xor U8713 (N_8713,N_8550,N_8605);
xor U8714 (N_8714,N_8536,N_8486);
or U8715 (N_8715,N_8607,N_8591);
or U8716 (N_8716,N_8492,N_8570);
and U8717 (N_8717,N_8586,N_8613);
nand U8718 (N_8718,N_8544,N_8583);
nand U8719 (N_8719,N_8493,N_8557);
and U8720 (N_8720,N_8597,N_8535);
xnor U8721 (N_8721,N_8491,N_8561);
nor U8722 (N_8722,N_8567,N_8565);
nor U8723 (N_8723,N_8620,N_8593);
or U8724 (N_8724,N_8523,N_8619);
and U8725 (N_8725,N_8492,N_8556);
or U8726 (N_8726,N_8632,N_8606);
and U8727 (N_8727,N_8628,N_8484);
nor U8728 (N_8728,N_8621,N_8601);
nand U8729 (N_8729,N_8505,N_8600);
xnor U8730 (N_8730,N_8540,N_8581);
nand U8731 (N_8731,N_8586,N_8638);
and U8732 (N_8732,N_8528,N_8525);
nor U8733 (N_8733,N_8581,N_8632);
or U8734 (N_8734,N_8619,N_8543);
or U8735 (N_8735,N_8607,N_8559);
and U8736 (N_8736,N_8628,N_8498);
and U8737 (N_8737,N_8571,N_8562);
or U8738 (N_8738,N_8581,N_8607);
or U8739 (N_8739,N_8627,N_8631);
xor U8740 (N_8740,N_8581,N_8624);
nor U8741 (N_8741,N_8617,N_8628);
xnor U8742 (N_8742,N_8597,N_8607);
or U8743 (N_8743,N_8522,N_8510);
nand U8744 (N_8744,N_8531,N_8587);
or U8745 (N_8745,N_8546,N_8626);
nor U8746 (N_8746,N_8551,N_8549);
nand U8747 (N_8747,N_8516,N_8633);
nand U8748 (N_8748,N_8524,N_8502);
nor U8749 (N_8749,N_8572,N_8535);
or U8750 (N_8750,N_8525,N_8568);
and U8751 (N_8751,N_8556,N_8571);
nand U8752 (N_8752,N_8538,N_8631);
and U8753 (N_8753,N_8608,N_8527);
nor U8754 (N_8754,N_8514,N_8570);
xnor U8755 (N_8755,N_8547,N_8638);
nand U8756 (N_8756,N_8495,N_8571);
nor U8757 (N_8757,N_8497,N_8638);
xor U8758 (N_8758,N_8553,N_8590);
xor U8759 (N_8759,N_8517,N_8584);
and U8760 (N_8760,N_8635,N_8634);
or U8761 (N_8761,N_8501,N_8504);
xnor U8762 (N_8762,N_8531,N_8571);
nor U8763 (N_8763,N_8543,N_8596);
xor U8764 (N_8764,N_8605,N_8509);
and U8765 (N_8765,N_8528,N_8638);
xnor U8766 (N_8766,N_8621,N_8497);
xnor U8767 (N_8767,N_8597,N_8637);
nor U8768 (N_8768,N_8597,N_8525);
nand U8769 (N_8769,N_8492,N_8531);
xor U8770 (N_8770,N_8603,N_8513);
nand U8771 (N_8771,N_8568,N_8489);
and U8772 (N_8772,N_8523,N_8515);
xor U8773 (N_8773,N_8490,N_8512);
or U8774 (N_8774,N_8562,N_8605);
or U8775 (N_8775,N_8597,N_8537);
and U8776 (N_8776,N_8626,N_8529);
xor U8777 (N_8777,N_8596,N_8634);
nor U8778 (N_8778,N_8488,N_8555);
and U8779 (N_8779,N_8609,N_8489);
or U8780 (N_8780,N_8507,N_8517);
or U8781 (N_8781,N_8513,N_8548);
nand U8782 (N_8782,N_8504,N_8519);
nand U8783 (N_8783,N_8549,N_8555);
nand U8784 (N_8784,N_8616,N_8568);
and U8785 (N_8785,N_8543,N_8512);
xor U8786 (N_8786,N_8576,N_8564);
or U8787 (N_8787,N_8517,N_8619);
or U8788 (N_8788,N_8508,N_8560);
or U8789 (N_8789,N_8582,N_8508);
xnor U8790 (N_8790,N_8624,N_8520);
nor U8791 (N_8791,N_8609,N_8492);
nand U8792 (N_8792,N_8591,N_8572);
nand U8793 (N_8793,N_8482,N_8546);
nor U8794 (N_8794,N_8519,N_8482);
nor U8795 (N_8795,N_8585,N_8545);
nand U8796 (N_8796,N_8497,N_8504);
nand U8797 (N_8797,N_8548,N_8495);
or U8798 (N_8798,N_8518,N_8488);
xor U8799 (N_8799,N_8596,N_8611);
and U8800 (N_8800,N_8773,N_8752);
and U8801 (N_8801,N_8686,N_8774);
nor U8802 (N_8802,N_8798,N_8654);
nand U8803 (N_8803,N_8720,N_8709);
xor U8804 (N_8804,N_8664,N_8663);
nor U8805 (N_8805,N_8667,N_8756);
xor U8806 (N_8806,N_8685,N_8697);
or U8807 (N_8807,N_8710,N_8688);
xnor U8808 (N_8808,N_8699,N_8706);
xnor U8809 (N_8809,N_8791,N_8769);
or U8810 (N_8810,N_8708,N_8764);
xnor U8811 (N_8811,N_8722,N_8660);
nand U8812 (N_8812,N_8726,N_8658);
and U8813 (N_8813,N_8747,N_8781);
nor U8814 (N_8814,N_8641,N_8775);
xor U8815 (N_8815,N_8653,N_8787);
xnor U8816 (N_8816,N_8724,N_8647);
nand U8817 (N_8817,N_8717,N_8770);
nand U8818 (N_8818,N_8691,N_8668);
xor U8819 (N_8819,N_8694,N_8777);
nor U8820 (N_8820,N_8753,N_8671);
nor U8821 (N_8821,N_8767,N_8799);
nor U8822 (N_8822,N_8744,N_8696);
xor U8823 (N_8823,N_8736,N_8716);
and U8824 (N_8824,N_8788,N_8760);
nand U8825 (N_8825,N_8795,N_8678);
or U8826 (N_8826,N_8758,N_8739);
or U8827 (N_8827,N_8683,N_8714);
and U8828 (N_8828,N_8754,N_8711);
or U8829 (N_8829,N_8785,N_8677);
and U8830 (N_8830,N_8784,N_8674);
xnor U8831 (N_8831,N_8790,N_8650);
or U8832 (N_8832,N_8651,N_8682);
and U8833 (N_8833,N_8649,N_8745);
or U8834 (N_8834,N_8733,N_8762);
nor U8835 (N_8835,N_8780,N_8797);
nor U8836 (N_8836,N_8771,N_8734);
xnor U8837 (N_8837,N_8675,N_8738);
xor U8838 (N_8838,N_8778,N_8643);
nor U8839 (N_8839,N_8721,N_8676);
nor U8840 (N_8840,N_8761,N_8765);
nor U8841 (N_8841,N_8692,N_8743);
xor U8842 (N_8842,N_8687,N_8693);
and U8843 (N_8843,N_8792,N_8703);
or U8844 (N_8844,N_8700,N_8695);
or U8845 (N_8845,N_8672,N_8742);
and U8846 (N_8846,N_8698,N_8645);
nand U8847 (N_8847,N_8679,N_8746);
nor U8848 (N_8848,N_8719,N_8732);
and U8849 (N_8849,N_8656,N_8757);
nand U8850 (N_8850,N_8665,N_8766);
and U8851 (N_8851,N_8735,N_8646);
or U8852 (N_8852,N_8670,N_8680);
xor U8853 (N_8853,N_8759,N_8715);
nor U8854 (N_8854,N_8748,N_8728);
nor U8855 (N_8855,N_8684,N_8750);
xnor U8856 (N_8856,N_8713,N_8776);
or U8857 (N_8857,N_8657,N_8718);
nand U8858 (N_8858,N_8749,N_8755);
nand U8859 (N_8859,N_8690,N_8707);
or U8860 (N_8860,N_8725,N_8669);
nand U8861 (N_8861,N_8723,N_8730);
nand U8862 (N_8862,N_8727,N_8768);
and U8863 (N_8863,N_8794,N_8779);
and U8864 (N_8864,N_8659,N_8789);
nor U8865 (N_8865,N_8729,N_8763);
or U8866 (N_8866,N_8796,N_8740);
nor U8867 (N_8867,N_8648,N_8655);
nor U8868 (N_8868,N_8741,N_8712);
and U8869 (N_8869,N_8731,N_8642);
or U8870 (N_8870,N_8681,N_8704);
and U8871 (N_8871,N_8652,N_8783);
and U8872 (N_8872,N_8737,N_8702);
nand U8873 (N_8873,N_8772,N_8666);
or U8874 (N_8874,N_8786,N_8689);
or U8875 (N_8875,N_8640,N_8644);
nand U8876 (N_8876,N_8782,N_8751);
nor U8877 (N_8877,N_8793,N_8701);
or U8878 (N_8878,N_8673,N_8705);
nor U8879 (N_8879,N_8661,N_8662);
or U8880 (N_8880,N_8643,N_8683);
and U8881 (N_8881,N_8670,N_8767);
nand U8882 (N_8882,N_8747,N_8691);
nor U8883 (N_8883,N_8674,N_8683);
and U8884 (N_8884,N_8793,N_8777);
xnor U8885 (N_8885,N_8775,N_8657);
xnor U8886 (N_8886,N_8662,N_8799);
nand U8887 (N_8887,N_8655,N_8684);
or U8888 (N_8888,N_8745,N_8797);
or U8889 (N_8889,N_8747,N_8740);
and U8890 (N_8890,N_8738,N_8768);
nand U8891 (N_8891,N_8705,N_8641);
xor U8892 (N_8892,N_8669,N_8674);
or U8893 (N_8893,N_8655,N_8650);
and U8894 (N_8894,N_8700,N_8665);
nor U8895 (N_8895,N_8728,N_8796);
or U8896 (N_8896,N_8763,N_8688);
nor U8897 (N_8897,N_8730,N_8681);
and U8898 (N_8898,N_8782,N_8645);
nand U8899 (N_8899,N_8659,N_8739);
xnor U8900 (N_8900,N_8751,N_8729);
xor U8901 (N_8901,N_8747,N_8765);
and U8902 (N_8902,N_8654,N_8786);
or U8903 (N_8903,N_8746,N_8780);
nand U8904 (N_8904,N_8681,N_8794);
or U8905 (N_8905,N_8724,N_8731);
and U8906 (N_8906,N_8771,N_8691);
nor U8907 (N_8907,N_8783,N_8716);
nor U8908 (N_8908,N_8718,N_8698);
nand U8909 (N_8909,N_8665,N_8788);
xor U8910 (N_8910,N_8724,N_8728);
xor U8911 (N_8911,N_8644,N_8657);
or U8912 (N_8912,N_8712,N_8761);
nand U8913 (N_8913,N_8708,N_8766);
xnor U8914 (N_8914,N_8792,N_8791);
nor U8915 (N_8915,N_8742,N_8733);
nand U8916 (N_8916,N_8753,N_8780);
xnor U8917 (N_8917,N_8727,N_8767);
or U8918 (N_8918,N_8761,N_8724);
and U8919 (N_8919,N_8755,N_8675);
or U8920 (N_8920,N_8732,N_8751);
xor U8921 (N_8921,N_8657,N_8723);
and U8922 (N_8922,N_8760,N_8754);
and U8923 (N_8923,N_8699,N_8748);
and U8924 (N_8924,N_8666,N_8709);
and U8925 (N_8925,N_8688,N_8693);
or U8926 (N_8926,N_8656,N_8779);
xor U8927 (N_8927,N_8732,N_8660);
or U8928 (N_8928,N_8725,N_8744);
nand U8929 (N_8929,N_8743,N_8677);
xnor U8930 (N_8930,N_8690,N_8784);
and U8931 (N_8931,N_8699,N_8653);
nand U8932 (N_8932,N_8679,N_8762);
and U8933 (N_8933,N_8756,N_8693);
xor U8934 (N_8934,N_8745,N_8655);
nor U8935 (N_8935,N_8761,N_8748);
or U8936 (N_8936,N_8766,N_8705);
nand U8937 (N_8937,N_8707,N_8742);
xnor U8938 (N_8938,N_8704,N_8713);
and U8939 (N_8939,N_8689,N_8729);
xor U8940 (N_8940,N_8705,N_8644);
nand U8941 (N_8941,N_8754,N_8793);
xnor U8942 (N_8942,N_8735,N_8757);
xor U8943 (N_8943,N_8730,N_8769);
or U8944 (N_8944,N_8709,N_8724);
nand U8945 (N_8945,N_8764,N_8723);
or U8946 (N_8946,N_8706,N_8755);
nor U8947 (N_8947,N_8709,N_8656);
or U8948 (N_8948,N_8777,N_8698);
and U8949 (N_8949,N_8721,N_8771);
nand U8950 (N_8950,N_8769,N_8650);
nor U8951 (N_8951,N_8728,N_8749);
xor U8952 (N_8952,N_8700,N_8710);
or U8953 (N_8953,N_8732,N_8668);
nand U8954 (N_8954,N_8688,N_8716);
or U8955 (N_8955,N_8719,N_8658);
xor U8956 (N_8956,N_8772,N_8787);
nor U8957 (N_8957,N_8653,N_8794);
xor U8958 (N_8958,N_8711,N_8728);
and U8959 (N_8959,N_8661,N_8669);
xnor U8960 (N_8960,N_8948,N_8943);
xnor U8961 (N_8961,N_8811,N_8851);
xor U8962 (N_8962,N_8847,N_8933);
and U8963 (N_8963,N_8925,N_8853);
xor U8964 (N_8964,N_8821,N_8806);
or U8965 (N_8965,N_8843,N_8824);
xor U8966 (N_8966,N_8862,N_8803);
xor U8967 (N_8967,N_8873,N_8952);
and U8968 (N_8968,N_8841,N_8831);
nor U8969 (N_8969,N_8856,N_8860);
or U8970 (N_8970,N_8867,N_8926);
nor U8971 (N_8971,N_8953,N_8822);
or U8972 (N_8972,N_8904,N_8813);
nand U8973 (N_8973,N_8839,N_8917);
nand U8974 (N_8974,N_8914,N_8954);
or U8975 (N_8975,N_8950,N_8901);
xor U8976 (N_8976,N_8840,N_8956);
and U8977 (N_8977,N_8949,N_8946);
or U8978 (N_8978,N_8820,N_8842);
nor U8979 (N_8979,N_8834,N_8898);
and U8980 (N_8980,N_8912,N_8855);
nor U8981 (N_8981,N_8823,N_8832);
nor U8982 (N_8982,N_8909,N_8878);
nand U8983 (N_8983,N_8868,N_8886);
or U8984 (N_8984,N_8807,N_8902);
nand U8985 (N_8985,N_8939,N_8876);
nor U8986 (N_8986,N_8830,N_8893);
nor U8987 (N_8987,N_8866,N_8857);
and U8988 (N_8988,N_8828,N_8864);
nand U8989 (N_8989,N_8833,N_8815);
or U8990 (N_8990,N_8908,N_8883);
nand U8991 (N_8991,N_8836,N_8848);
nor U8992 (N_8992,N_8881,N_8935);
nor U8993 (N_8993,N_8920,N_8919);
xnor U8994 (N_8994,N_8882,N_8812);
or U8995 (N_8995,N_8814,N_8896);
xnor U8996 (N_8996,N_8889,N_8869);
and U8997 (N_8997,N_8931,N_8850);
and U8998 (N_8998,N_8861,N_8957);
nand U8999 (N_8999,N_8955,N_8958);
nor U9000 (N_9000,N_8825,N_8819);
nor U9001 (N_9001,N_8880,N_8802);
or U9002 (N_9002,N_8945,N_8906);
xor U9003 (N_9003,N_8877,N_8849);
or U9004 (N_9004,N_8863,N_8959);
xor U9005 (N_9005,N_8894,N_8846);
nand U9006 (N_9006,N_8907,N_8818);
nor U9007 (N_9007,N_8899,N_8944);
nor U9008 (N_9008,N_8844,N_8929);
or U9009 (N_9009,N_8942,N_8936);
nor U9010 (N_9010,N_8941,N_8891);
nor U9011 (N_9011,N_8927,N_8951);
xnor U9012 (N_9012,N_8879,N_8816);
or U9013 (N_9013,N_8910,N_8801);
nor U9014 (N_9014,N_8872,N_8921);
nor U9015 (N_9015,N_8810,N_8918);
or U9016 (N_9016,N_8911,N_8903);
or U9017 (N_9017,N_8940,N_8829);
nand U9018 (N_9018,N_8938,N_8838);
and U9019 (N_9019,N_8808,N_8865);
nor U9020 (N_9020,N_8887,N_8905);
nand U9021 (N_9021,N_8930,N_8817);
and U9022 (N_9022,N_8892,N_8845);
nand U9023 (N_9023,N_8934,N_8897);
or U9024 (N_9024,N_8900,N_8895);
and U9025 (N_9025,N_8884,N_8859);
or U9026 (N_9026,N_8852,N_8854);
or U9027 (N_9027,N_8947,N_8924);
or U9028 (N_9028,N_8837,N_8858);
nor U9029 (N_9029,N_8915,N_8835);
nor U9030 (N_9030,N_8916,N_8804);
nor U9031 (N_9031,N_8870,N_8871);
nand U9032 (N_9032,N_8809,N_8805);
or U9033 (N_9033,N_8932,N_8923);
xnor U9034 (N_9034,N_8827,N_8875);
nor U9035 (N_9035,N_8800,N_8913);
and U9036 (N_9036,N_8937,N_8890);
xnor U9037 (N_9037,N_8826,N_8888);
nor U9038 (N_9038,N_8885,N_8928);
nand U9039 (N_9039,N_8922,N_8874);
or U9040 (N_9040,N_8921,N_8846);
and U9041 (N_9041,N_8843,N_8860);
or U9042 (N_9042,N_8922,N_8862);
nor U9043 (N_9043,N_8930,N_8831);
or U9044 (N_9044,N_8860,N_8897);
xor U9045 (N_9045,N_8845,N_8809);
and U9046 (N_9046,N_8928,N_8846);
nand U9047 (N_9047,N_8956,N_8948);
xor U9048 (N_9048,N_8956,N_8863);
or U9049 (N_9049,N_8888,N_8812);
xor U9050 (N_9050,N_8926,N_8871);
or U9051 (N_9051,N_8801,N_8905);
xor U9052 (N_9052,N_8880,N_8935);
or U9053 (N_9053,N_8888,N_8836);
nand U9054 (N_9054,N_8946,N_8957);
nor U9055 (N_9055,N_8866,N_8949);
nor U9056 (N_9056,N_8918,N_8950);
or U9057 (N_9057,N_8814,N_8875);
nor U9058 (N_9058,N_8943,N_8910);
or U9059 (N_9059,N_8852,N_8904);
xnor U9060 (N_9060,N_8894,N_8888);
and U9061 (N_9061,N_8940,N_8895);
xor U9062 (N_9062,N_8889,N_8899);
nand U9063 (N_9063,N_8878,N_8856);
nor U9064 (N_9064,N_8943,N_8949);
nand U9065 (N_9065,N_8818,N_8823);
nand U9066 (N_9066,N_8950,N_8920);
or U9067 (N_9067,N_8903,N_8841);
or U9068 (N_9068,N_8862,N_8816);
and U9069 (N_9069,N_8895,N_8816);
xnor U9070 (N_9070,N_8959,N_8846);
nor U9071 (N_9071,N_8824,N_8882);
xnor U9072 (N_9072,N_8824,N_8953);
and U9073 (N_9073,N_8861,N_8923);
nor U9074 (N_9074,N_8827,N_8857);
nor U9075 (N_9075,N_8818,N_8812);
and U9076 (N_9076,N_8842,N_8893);
or U9077 (N_9077,N_8911,N_8829);
or U9078 (N_9078,N_8836,N_8949);
and U9079 (N_9079,N_8813,N_8802);
nor U9080 (N_9080,N_8871,N_8822);
or U9081 (N_9081,N_8923,N_8845);
or U9082 (N_9082,N_8824,N_8881);
nand U9083 (N_9083,N_8855,N_8926);
nor U9084 (N_9084,N_8916,N_8938);
and U9085 (N_9085,N_8953,N_8894);
xnor U9086 (N_9086,N_8908,N_8862);
nor U9087 (N_9087,N_8945,N_8855);
xor U9088 (N_9088,N_8925,N_8807);
or U9089 (N_9089,N_8946,N_8803);
nand U9090 (N_9090,N_8887,N_8942);
and U9091 (N_9091,N_8943,N_8824);
xor U9092 (N_9092,N_8813,N_8896);
nor U9093 (N_9093,N_8926,N_8891);
nor U9094 (N_9094,N_8916,N_8870);
and U9095 (N_9095,N_8827,N_8899);
and U9096 (N_9096,N_8819,N_8923);
and U9097 (N_9097,N_8884,N_8800);
xnor U9098 (N_9098,N_8800,N_8807);
or U9099 (N_9099,N_8937,N_8938);
xnor U9100 (N_9100,N_8936,N_8908);
and U9101 (N_9101,N_8931,N_8851);
nand U9102 (N_9102,N_8861,N_8927);
and U9103 (N_9103,N_8860,N_8937);
nand U9104 (N_9104,N_8820,N_8945);
and U9105 (N_9105,N_8805,N_8909);
xor U9106 (N_9106,N_8845,N_8806);
nand U9107 (N_9107,N_8826,N_8844);
xor U9108 (N_9108,N_8829,N_8855);
or U9109 (N_9109,N_8816,N_8882);
xnor U9110 (N_9110,N_8904,N_8888);
nand U9111 (N_9111,N_8839,N_8910);
nand U9112 (N_9112,N_8838,N_8830);
xor U9113 (N_9113,N_8815,N_8865);
and U9114 (N_9114,N_8820,N_8904);
and U9115 (N_9115,N_8951,N_8875);
nor U9116 (N_9116,N_8935,N_8827);
and U9117 (N_9117,N_8914,N_8812);
or U9118 (N_9118,N_8853,N_8899);
nand U9119 (N_9119,N_8959,N_8938);
nor U9120 (N_9120,N_9047,N_8970);
nand U9121 (N_9121,N_9023,N_8991);
nand U9122 (N_9122,N_9113,N_9119);
or U9123 (N_9123,N_8990,N_9079);
nand U9124 (N_9124,N_9044,N_9108);
xor U9125 (N_9125,N_8987,N_9078);
xnor U9126 (N_9126,N_9006,N_9067);
or U9127 (N_9127,N_9036,N_9109);
and U9128 (N_9128,N_9086,N_9014);
and U9129 (N_9129,N_9083,N_9071);
xor U9130 (N_9130,N_9062,N_9076);
nand U9131 (N_9131,N_9055,N_9016);
nand U9132 (N_9132,N_9033,N_9097);
nand U9133 (N_9133,N_9061,N_9038);
xor U9134 (N_9134,N_8982,N_8960);
and U9135 (N_9135,N_9018,N_9104);
nor U9136 (N_9136,N_8974,N_9030);
nand U9137 (N_9137,N_9054,N_8975);
xor U9138 (N_9138,N_9080,N_9089);
and U9139 (N_9139,N_9019,N_8979);
and U9140 (N_9140,N_9117,N_9042);
or U9141 (N_9141,N_8973,N_8967);
or U9142 (N_9142,N_9091,N_9077);
nor U9143 (N_9143,N_9082,N_9060);
nand U9144 (N_9144,N_8962,N_9065);
nand U9145 (N_9145,N_8972,N_8968);
or U9146 (N_9146,N_8983,N_9081);
xor U9147 (N_9147,N_9028,N_9029);
xnor U9148 (N_9148,N_8996,N_9051);
or U9149 (N_9149,N_8997,N_8961);
xor U9150 (N_9150,N_9064,N_9010);
and U9151 (N_9151,N_8984,N_9073);
nand U9152 (N_9152,N_9003,N_9072);
xnor U9153 (N_9153,N_9090,N_8966);
nor U9154 (N_9154,N_9074,N_9068);
nand U9155 (N_9155,N_8969,N_9093);
and U9156 (N_9156,N_9106,N_9008);
nand U9157 (N_9157,N_9011,N_9114);
and U9158 (N_9158,N_8977,N_9001);
or U9159 (N_9159,N_8988,N_9024);
or U9160 (N_9160,N_9118,N_9115);
and U9161 (N_9161,N_9020,N_9111);
xnor U9162 (N_9162,N_9009,N_8976);
and U9163 (N_9163,N_9000,N_9092);
or U9164 (N_9164,N_9039,N_9035);
xor U9165 (N_9165,N_9085,N_9049);
nor U9166 (N_9166,N_9059,N_9063);
xnor U9167 (N_9167,N_9057,N_9084);
nor U9168 (N_9168,N_8986,N_8994);
nand U9169 (N_9169,N_9070,N_9099);
nand U9170 (N_9170,N_8981,N_8993);
or U9171 (N_9171,N_9100,N_9046);
or U9172 (N_9172,N_9052,N_9058);
nand U9173 (N_9173,N_9017,N_9107);
nand U9174 (N_9174,N_9015,N_8995);
and U9175 (N_9175,N_9053,N_9094);
or U9176 (N_9176,N_9087,N_9102);
and U9177 (N_9177,N_9007,N_9095);
xnor U9178 (N_9178,N_9096,N_9037);
or U9179 (N_9179,N_9013,N_9021);
or U9180 (N_9180,N_8992,N_9027);
xor U9181 (N_9181,N_9031,N_8964);
and U9182 (N_9182,N_9101,N_9050);
nand U9183 (N_9183,N_9026,N_9005);
nand U9184 (N_9184,N_8965,N_9098);
xnor U9185 (N_9185,N_9103,N_9112);
or U9186 (N_9186,N_9075,N_8971);
nor U9187 (N_9187,N_9110,N_8978);
and U9188 (N_9188,N_9048,N_9032);
or U9189 (N_9189,N_9045,N_9116);
or U9190 (N_9190,N_9043,N_8963);
or U9191 (N_9191,N_9066,N_9056);
nand U9192 (N_9192,N_8980,N_8985);
and U9193 (N_9193,N_8999,N_8998);
or U9194 (N_9194,N_9002,N_9004);
or U9195 (N_9195,N_9088,N_9012);
xor U9196 (N_9196,N_8989,N_9022);
xor U9197 (N_9197,N_9040,N_9025);
nor U9198 (N_9198,N_9069,N_9041);
and U9199 (N_9199,N_9034,N_9105);
xnor U9200 (N_9200,N_9097,N_9053);
nor U9201 (N_9201,N_9042,N_8996);
and U9202 (N_9202,N_9067,N_8977);
or U9203 (N_9203,N_9031,N_9081);
or U9204 (N_9204,N_9067,N_8981);
nand U9205 (N_9205,N_9067,N_9016);
nor U9206 (N_9206,N_8988,N_9010);
or U9207 (N_9207,N_9092,N_9067);
and U9208 (N_9208,N_9117,N_9066);
nand U9209 (N_9209,N_8960,N_9100);
or U9210 (N_9210,N_9016,N_9026);
nor U9211 (N_9211,N_8997,N_9105);
nor U9212 (N_9212,N_8978,N_9002);
or U9213 (N_9213,N_9098,N_8998);
xnor U9214 (N_9214,N_9090,N_9054);
or U9215 (N_9215,N_9118,N_9015);
or U9216 (N_9216,N_9112,N_9077);
nand U9217 (N_9217,N_9076,N_9043);
xnor U9218 (N_9218,N_9085,N_9003);
nor U9219 (N_9219,N_9075,N_8995);
and U9220 (N_9220,N_9079,N_8976);
xnor U9221 (N_9221,N_9084,N_9097);
and U9222 (N_9222,N_9036,N_9011);
nand U9223 (N_9223,N_9074,N_9032);
and U9224 (N_9224,N_9066,N_9104);
nand U9225 (N_9225,N_8979,N_9028);
nor U9226 (N_9226,N_8967,N_9066);
nor U9227 (N_9227,N_9071,N_8998);
nand U9228 (N_9228,N_9064,N_9036);
nand U9229 (N_9229,N_8963,N_9057);
or U9230 (N_9230,N_9107,N_9092);
and U9231 (N_9231,N_9095,N_8967);
or U9232 (N_9232,N_9093,N_9054);
nor U9233 (N_9233,N_9035,N_9030);
xor U9234 (N_9234,N_9062,N_9060);
nor U9235 (N_9235,N_9029,N_9068);
and U9236 (N_9236,N_8994,N_9058);
xnor U9237 (N_9237,N_8963,N_9096);
or U9238 (N_9238,N_9016,N_9011);
and U9239 (N_9239,N_9030,N_8997);
xor U9240 (N_9240,N_9111,N_8969);
nor U9241 (N_9241,N_9038,N_9073);
nor U9242 (N_9242,N_9050,N_9075);
xor U9243 (N_9243,N_9043,N_9014);
or U9244 (N_9244,N_9077,N_9055);
xnor U9245 (N_9245,N_8999,N_9071);
nand U9246 (N_9246,N_9112,N_9007);
xor U9247 (N_9247,N_9061,N_9055);
or U9248 (N_9248,N_9002,N_9046);
or U9249 (N_9249,N_9098,N_8968);
or U9250 (N_9250,N_9000,N_8987);
nand U9251 (N_9251,N_9107,N_9023);
nor U9252 (N_9252,N_9093,N_8988);
nor U9253 (N_9253,N_9009,N_9119);
nand U9254 (N_9254,N_9116,N_9065);
or U9255 (N_9255,N_9099,N_9055);
nor U9256 (N_9256,N_9042,N_8976);
nand U9257 (N_9257,N_9087,N_9043);
or U9258 (N_9258,N_9075,N_8968);
xor U9259 (N_9259,N_8997,N_9013);
xor U9260 (N_9260,N_9074,N_9052);
or U9261 (N_9261,N_8995,N_9097);
nand U9262 (N_9262,N_9098,N_8960);
xnor U9263 (N_9263,N_9083,N_9062);
nand U9264 (N_9264,N_9024,N_9044);
nor U9265 (N_9265,N_8964,N_9073);
or U9266 (N_9266,N_9078,N_8980);
nand U9267 (N_9267,N_9052,N_8961);
or U9268 (N_9268,N_9040,N_8994);
xnor U9269 (N_9269,N_9047,N_9070);
nor U9270 (N_9270,N_9119,N_9099);
xor U9271 (N_9271,N_8981,N_9019);
nor U9272 (N_9272,N_8992,N_9060);
and U9273 (N_9273,N_9093,N_9024);
nor U9274 (N_9274,N_9070,N_9056);
nor U9275 (N_9275,N_8994,N_9073);
or U9276 (N_9276,N_9110,N_8969);
or U9277 (N_9277,N_9112,N_9109);
and U9278 (N_9278,N_9025,N_8967);
nand U9279 (N_9279,N_8962,N_8982);
nand U9280 (N_9280,N_9238,N_9187);
xnor U9281 (N_9281,N_9135,N_9189);
or U9282 (N_9282,N_9169,N_9124);
or U9283 (N_9283,N_9200,N_9165);
nand U9284 (N_9284,N_9232,N_9196);
or U9285 (N_9285,N_9137,N_9258);
xor U9286 (N_9286,N_9166,N_9184);
xnor U9287 (N_9287,N_9193,N_9229);
xor U9288 (N_9288,N_9235,N_9242);
nor U9289 (N_9289,N_9228,N_9253);
or U9290 (N_9290,N_9263,N_9239);
and U9291 (N_9291,N_9222,N_9148);
nor U9292 (N_9292,N_9233,N_9139);
nand U9293 (N_9293,N_9218,N_9248);
nand U9294 (N_9294,N_9131,N_9206);
and U9295 (N_9295,N_9154,N_9252);
nand U9296 (N_9296,N_9278,N_9132);
nor U9297 (N_9297,N_9126,N_9171);
xnor U9298 (N_9298,N_9257,N_9237);
nand U9299 (N_9299,N_9246,N_9264);
nor U9300 (N_9300,N_9152,N_9244);
or U9301 (N_9301,N_9217,N_9256);
xor U9302 (N_9302,N_9142,N_9122);
nor U9303 (N_9303,N_9213,N_9129);
nand U9304 (N_9304,N_9134,N_9143);
and U9305 (N_9305,N_9163,N_9262);
xnor U9306 (N_9306,N_9153,N_9150);
nor U9307 (N_9307,N_9121,N_9260);
nand U9308 (N_9308,N_9130,N_9211);
nand U9309 (N_9309,N_9199,N_9234);
and U9310 (N_9310,N_9266,N_9145);
or U9311 (N_9311,N_9147,N_9174);
xor U9312 (N_9312,N_9128,N_9191);
nand U9313 (N_9313,N_9255,N_9172);
nand U9314 (N_9314,N_9197,N_9123);
nand U9315 (N_9315,N_9159,N_9269);
or U9316 (N_9316,N_9270,N_9219);
and U9317 (N_9317,N_9204,N_9138);
or U9318 (N_9318,N_9195,N_9168);
xor U9319 (N_9319,N_9220,N_9251);
xnor U9320 (N_9320,N_9136,N_9203);
nand U9321 (N_9321,N_9144,N_9167);
xnor U9322 (N_9322,N_9201,N_9223);
xnor U9323 (N_9323,N_9198,N_9180);
and U9324 (N_9324,N_9276,N_9140);
or U9325 (N_9325,N_9271,N_9164);
xnor U9326 (N_9326,N_9208,N_9236);
nand U9327 (N_9327,N_9190,N_9162);
or U9328 (N_9328,N_9182,N_9151);
nand U9329 (N_9329,N_9177,N_9254);
or U9330 (N_9330,N_9157,N_9212);
xor U9331 (N_9331,N_9240,N_9181);
or U9332 (N_9332,N_9230,N_9158);
nor U9333 (N_9333,N_9202,N_9149);
or U9334 (N_9334,N_9216,N_9249);
and U9335 (N_9335,N_9178,N_9170);
nand U9336 (N_9336,N_9250,N_9194);
and U9337 (N_9337,N_9267,N_9245);
nand U9338 (N_9338,N_9155,N_9225);
nor U9339 (N_9339,N_9175,N_9259);
nor U9340 (N_9340,N_9146,N_9179);
nand U9341 (N_9341,N_9183,N_9141);
or U9342 (N_9342,N_9272,N_9277);
and U9343 (N_9343,N_9161,N_9268);
or U9344 (N_9344,N_9215,N_9127);
or U9345 (N_9345,N_9185,N_9173);
nand U9346 (N_9346,N_9209,N_9241);
and U9347 (N_9347,N_9231,N_9188);
xnor U9348 (N_9348,N_9275,N_9221);
or U9349 (N_9349,N_9176,N_9133);
and U9350 (N_9350,N_9226,N_9265);
or U9351 (N_9351,N_9120,N_9186);
and U9352 (N_9352,N_9192,N_9224);
and U9353 (N_9353,N_9210,N_9160);
or U9354 (N_9354,N_9227,N_9273);
or U9355 (N_9355,N_9243,N_9261);
or U9356 (N_9356,N_9205,N_9207);
nor U9357 (N_9357,N_9274,N_9156);
nor U9358 (N_9358,N_9247,N_9125);
nand U9359 (N_9359,N_9279,N_9214);
and U9360 (N_9360,N_9245,N_9139);
xnor U9361 (N_9361,N_9201,N_9199);
nand U9362 (N_9362,N_9127,N_9120);
or U9363 (N_9363,N_9267,N_9158);
xor U9364 (N_9364,N_9272,N_9198);
xor U9365 (N_9365,N_9127,N_9130);
nor U9366 (N_9366,N_9151,N_9191);
xnor U9367 (N_9367,N_9163,N_9208);
nand U9368 (N_9368,N_9130,N_9244);
or U9369 (N_9369,N_9127,N_9277);
xor U9370 (N_9370,N_9261,N_9257);
nor U9371 (N_9371,N_9246,N_9228);
nor U9372 (N_9372,N_9142,N_9193);
xnor U9373 (N_9373,N_9214,N_9208);
xor U9374 (N_9374,N_9254,N_9246);
and U9375 (N_9375,N_9120,N_9258);
or U9376 (N_9376,N_9193,N_9153);
or U9377 (N_9377,N_9197,N_9226);
or U9378 (N_9378,N_9160,N_9213);
and U9379 (N_9379,N_9275,N_9141);
nand U9380 (N_9380,N_9127,N_9275);
nand U9381 (N_9381,N_9142,N_9187);
nand U9382 (N_9382,N_9123,N_9215);
nand U9383 (N_9383,N_9234,N_9173);
or U9384 (N_9384,N_9199,N_9181);
nand U9385 (N_9385,N_9139,N_9261);
nand U9386 (N_9386,N_9206,N_9164);
xor U9387 (N_9387,N_9159,N_9256);
or U9388 (N_9388,N_9200,N_9235);
and U9389 (N_9389,N_9136,N_9274);
xor U9390 (N_9390,N_9243,N_9212);
or U9391 (N_9391,N_9228,N_9125);
and U9392 (N_9392,N_9238,N_9258);
or U9393 (N_9393,N_9217,N_9178);
nand U9394 (N_9394,N_9134,N_9168);
and U9395 (N_9395,N_9146,N_9163);
or U9396 (N_9396,N_9144,N_9148);
and U9397 (N_9397,N_9172,N_9169);
nor U9398 (N_9398,N_9206,N_9178);
nor U9399 (N_9399,N_9157,N_9235);
nor U9400 (N_9400,N_9140,N_9189);
or U9401 (N_9401,N_9192,N_9202);
xnor U9402 (N_9402,N_9272,N_9132);
xor U9403 (N_9403,N_9133,N_9225);
xor U9404 (N_9404,N_9272,N_9190);
nand U9405 (N_9405,N_9253,N_9245);
or U9406 (N_9406,N_9167,N_9259);
nor U9407 (N_9407,N_9258,N_9268);
nor U9408 (N_9408,N_9164,N_9124);
nand U9409 (N_9409,N_9236,N_9226);
nor U9410 (N_9410,N_9211,N_9220);
nand U9411 (N_9411,N_9234,N_9244);
nor U9412 (N_9412,N_9238,N_9233);
nand U9413 (N_9413,N_9139,N_9141);
and U9414 (N_9414,N_9169,N_9229);
nor U9415 (N_9415,N_9226,N_9199);
nor U9416 (N_9416,N_9270,N_9182);
xnor U9417 (N_9417,N_9224,N_9168);
xnor U9418 (N_9418,N_9256,N_9144);
or U9419 (N_9419,N_9225,N_9153);
or U9420 (N_9420,N_9244,N_9228);
nor U9421 (N_9421,N_9121,N_9199);
nand U9422 (N_9422,N_9255,N_9227);
or U9423 (N_9423,N_9179,N_9245);
nor U9424 (N_9424,N_9139,N_9240);
or U9425 (N_9425,N_9223,N_9168);
and U9426 (N_9426,N_9182,N_9245);
or U9427 (N_9427,N_9251,N_9244);
nand U9428 (N_9428,N_9200,N_9125);
or U9429 (N_9429,N_9203,N_9155);
nor U9430 (N_9430,N_9157,N_9276);
xor U9431 (N_9431,N_9138,N_9253);
or U9432 (N_9432,N_9247,N_9143);
nor U9433 (N_9433,N_9226,N_9121);
nand U9434 (N_9434,N_9140,N_9193);
nand U9435 (N_9435,N_9181,N_9247);
nor U9436 (N_9436,N_9178,N_9143);
nand U9437 (N_9437,N_9145,N_9226);
xor U9438 (N_9438,N_9274,N_9273);
nor U9439 (N_9439,N_9143,N_9199);
nor U9440 (N_9440,N_9397,N_9371);
and U9441 (N_9441,N_9384,N_9387);
nand U9442 (N_9442,N_9435,N_9294);
or U9443 (N_9443,N_9300,N_9299);
nor U9444 (N_9444,N_9433,N_9365);
nand U9445 (N_9445,N_9291,N_9415);
nor U9446 (N_9446,N_9438,N_9336);
or U9447 (N_9447,N_9292,N_9411);
and U9448 (N_9448,N_9305,N_9417);
and U9449 (N_9449,N_9400,N_9301);
or U9450 (N_9450,N_9376,N_9385);
and U9451 (N_9451,N_9333,N_9367);
nand U9452 (N_9452,N_9394,N_9364);
or U9453 (N_9453,N_9287,N_9398);
xnor U9454 (N_9454,N_9401,N_9338);
and U9455 (N_9455,N_9379,N_9372);
and U9456 (N_9456,N_9361,N_9374);
nand U9457 (N_9457,N_9410,N_9334);
nand U9458 (N_9458,N_9363,N_9422);
or U9459 (N_9459,N_9418,N_9399);
nor U9460 (N_9460,N_9329,N_9310);
nor U9461 (N_9461,N_9437,N_9284);
and U9462 (N_9462,N_9351,N_9402);
and U9463 (N_9463,N_9405,N_9344);
nand U9464 (N_9464,N_9290,N_9357);
xnor U9465 (N_9465,N_9431,N_9308);
nor U9466 (N_9466,N_9359,N_9386);
nor U9467 (N_9467,N_9335,N_9315);
nand U9468 (N_9468,N_9413,N_9281);
and U9469 (N_9469,N_9286,N_9377);
nand U9470 (N_9470,N_9346,N_9375);
or U9471 (N_9471,N_9289,N_9341);
or U9472 (N_9472,N_9391,N_9436);
or U9473 (N_9473,N_9288,N_9404);
or U9474 (N_9474,N_9347,N_9409);
and U9475 (N_9475,N_9423,N_9358);
nor U9476 (N_9476,N_9362,N_9407);
xor U9477 (N_9477,N_9432,N_9370);
or U9478 (N_9478,N_9312,N_9378);
or U9479 (N_9479,N_9406,N_9350);
nand U9480 (N_9480,N_9317,N_9314);
nand U9481 (N_9481,N_9421,N_9313);
nor U9482 (N_9482,N_9393,N_9352);
nand U9483 (N_9483,N_9381,N_9320);
nand U9484 (N_9484,N_9354,N_9439);
nor U9485 (N_9485,N_9368,N_9337);
and U9486 (N_9486,N_9340,N_9343);
xor U9487 (N_9487,N_9285,N_9403);
or U9488 (N_9488,N_9321,N_9280);
and U9489 (N_9489,N_9296,N_9424);
nor U9490 (N_9490,N_9318,N_9353);
xnor U9491 (N_9491,N_9425,N_9295);
or U9492 (N_9492,N_9382,N_9360);
or U9493 (N_9493,N_9390,N_9328);
and U9494 (N_9494,N_9327,N_9369);
xnor U9495 (N_9495,N_9396,N_9389);
nor U9496 (N_9496,N_9380,N_9395);
xor U9497 (N_9497,N_9388,N_9306);
and U9498 (N_9498,N_9416,N_9373);
and U9499 (N_9499,N_9383,N_9419);
or U9500 (N_9500,N_9330,N_9326);
xnor U9501 (N_9501,N_9331,N_9430);
nor U9502 (N_9502,N_9304,N_9332);
or U9503 (N_9503,N_9302,N_9426);
nor U9504 (N_9504,N_9307,N_9309);
and U9505 (N_9505,N_9319,N_9392);
xnor U9506 (N_9506,N_9428,N_9322);
xnor U9507 (N_9507,N_9408,N_9412);
and U9508 (N_9508,N_9345,N_9356);
nor U9509 (N_9509,N_9293,N_9282);
nor U9510 (N_9510,N_9355,N_9342);
nor U9511 (N_9511,N_9366,N_9348);
nor U9512 (N_9512,N_9303,N_9420);
and U9513 (N_9513,N_9297,N_9298);
nor U9514 (N_9514,N_9324,N_9311);
and U9515 (N_9515,N_9339,N_9323);
or U9516 (N_9516,N_9434,N_9349);
nor U9517 (N_9517,N_9325,N_9283);
xnor U9518 (N_9518,N_9429,N_9414);
and U9519 (N_9519,N_9316,N_9427);
and U9520 (N_9520,N_9389,N_9338);
or U9521 (N_9521,N_9421,N_9434);
and U9522 (N_9522,N_9304,N_9363);
nand U9523 (N_9523,N_9406,N_9343);
nand U9524 (N_9524,N_9333,N_9287);
nand U9525 (N_9525,N_9394,N_9339);
nand U9526 (N_9526,N_9400,N_9382);
or U9527 (N_9527,N_9394,N_9326);
nand U9528 (N_9528,N_9380,N_9295);
nand U9529 (N_9529,N_9344,N_9280);
and U9530 (N_9530,N_9305,N_9304);
nor U9531 (N_9531,N_9401,N_9428);
xor U9532 (N_9532,N_9289,N_9362);
nor U9533 (N_9533,N_9301,N_9355);
nand U9534 (N_9534,N_9405,N_9428);
nor U9535 (N_9535,N_9313,N_9327);
nand U9536 (N_9536,N_9374,N_9396);
or U9537 (N_9537,N_9310,N_9382);
xor U9538 (N_9538,N_9360,N_9313);
or U9539 (N_9539,N_9317,N_9432);
nor U9540 (N_9540,N_9340,N_9366);
xor U9541 (N_9541,N_9423,N_9357);
xor U9542 (N_9542,N_9350,N_9402);
xor U9543 (N_9543,N_9389,N_9291);
nor U9544 (N_9544,N_9306,N_9333);
nand U9545 (N_9545,N_9295,N_9407);
or U9546 (N_9546,N_9368,N_9353);
or U9547 (N_9547,N_9280,N_9419);
xor U9548 (N_9548,N_9385,N_9349);
nand U9549 (N_9549,N_9337,N_9376);
and U9550 (N_9550,N_9428,N_9285);
nor U9551 (N_9551,N_9380,N_9283);
nor U9552 (N_9552,N_9357,N_9318);
and U9553 (N_9553,N_9366,N_9317);
and U9554 (N_9554,N_9433,N_9358);
or U9555 (N_9555,N_9359,N_9346);
xnor U9556 (N_9556,N_9380,N_9421);
nor U9557 (N_9557,N_9399,N_9412);
nor U9558 (N_9558,N_9329,N_9322);
or U9559 (N_9559,N_9310,N_9421);
and U9560 (N_9560,N_9395,N_9399);
or U9561 (N_9561,N_9419,N_9339);
xor U9562 (N_9562,N_9285,N_9418);
and U9563 (N_9563,N_9360,N_9372);
or U9564 (N_9564,N_9364,N_9436);
xnor U9565 (N_9565,N_9433,N_9438);
and U9566 (N_9566,N_9300,N_9328);
nor U9567 (N_9567,N_9377,N_9322);
xor U9568 (N_9568,N_9292,N_9314);
nor U9569 (N_9569,N_9320,N_9349);
or U9570 (N_9570,N_9286,N_9285);
nor U9571 (N_9571,N_9373,N_9312);
and U9572 (N_9572,N_9359,N_9352);
xnor U9573 (N_9573,N_9332,N_9396);
or U9574 (N_9574,N_9339,N_9329);
nand U9575 (N_9575,N_9295,N_9286);
or U9576 (N_9576,N_9361,N_9291);
nor U9577 (N_9577,N_9402,N_9403);
nand U9578 (N_9578,N_9336,N_9314);
or U9579 (N_9579,N_9355,N_9328);
nor U9580 (N_9580,N_9409,N_9289);
or U9581 (N_9581,N_9344,N_9336);
and U9582 (N_9582,N_9436,N_9341);
xnor U9583 (N_9583,N_9318,N_9338);
or U9584 (N_9584,N_9424,N_9338);
nand U9585 (N_9585,N_9308,N_9367);
or U9586 (N_9586,N_9432,N_9412);
and U9587 (N_9587,N_9419,N_9347);
and U9588 (N_9588,N_9289,N_9311);
nor U9589 (N_9589,N_9337,N_9321);
xor U9590 (N_9590,N_9337,N_9309);
and U9591 (N_9591,N_9305,N_9376);
or U9592 (N_9592,N_9388,N_9287);
or U9593 (N_9593,N_9294,N_9346);
xor U9594 (N_9594,N_9381,N_9411);
or U9595 (N_9595,N_9284,N_9418);
and U9596 (N_9596,N_9290,N_9373);
xor U9597 (N_9597,N_9364,N_9379);
xor U9598 (N_9598,N_9388,N_9319);
and U9599 (N_9599,N_9334,N_9307);
nor U9600 (N_9600,N_9555,N_9448);
nand U9601 (N_9601,N_9597,N_9532);
and U9602 (N_9602,N_9477,N_9514);
nand U9603 (N_9603,N_9599,N_9454);
nand U9604 (N_9604,N_9483,N_9465);
nand U9605 (N_9605,N_9549,N_9573);
nand U9606 (N_9606,N_9474,N_9510);
nor U9607 (N_9607,N_9476,N_9547);
xnor U9608 (N_9608,N_9468,N_9533);
and U9609 (N_9609,N_9472,N_9498);
or U9610 (N_9610,N_9564,N_9522);
nand U9611 (N_9611,N_9579,N_9525);
or U9612 (N_9612,N_9517,N_9445);
and U9613 (N_9613,N_9459,N_9570);
and U9614 (N_9614,N_9528,N_9586);
nor U9615 (N_9615,N_9482,N_9469);
nand U9616 (N_9616,N_9464,N_9512);
or U9617 (N_9617,N_9507,N_9557);
or U9618 (N_9618,N_9450,N_9592);
or U9619 (N_9619,N_9521,N_9538);
nor U9620 (N_9620,N_9488,N_9506);
and U9621 (N_9621,N_9572,N_9508);
nor U9622 (N_9622,N_9527,N_9475);
or U9623 (N_9623,N_9560,N_9554);
and U9624 (N_9624,N_9567,N_9545);
xor U9625 (N_9625,N_9568,N_9504);
or U9626 (N_9626,N_9453,N_9496);
nand U9627 (N_9627,N_9487,N_9451);
and U9628 (N_9628,N_9523,N_9544);
xnor U9629 (N_9629,N_9542,N_9509);
nor U9630 (N_9630,N_9582,N_9561);
and U9631 (N_9631,N_9574,N_9580);
nand U9632 (N_9632,N_9553,N_9478);
nor U9633 (N_9633,N_9558,N_9490);
nor U9634 (N_9634,N_9484,N_9443);
and U9635 (N_9635,N_9563,N_9565);
nor U9636 (N_9636,N_9536,N_9587);
nor U9637 (N_9637,N_9576,N_9534);
nand U9638 (N_9638,N_9497,N_9492);
nand U9639 (N_9639,N_9452,N_9460);
and U9640 (N_9640,N_9591,N_9589);
or U9641 (N_9641,N_9455,N_9585);
or U9642 (N_9642,N_9458,N_9505);
nor U9643 (N_9643,N_9539,N_9531);
xor U9644 (N_9644,N_9526,N_9449);
or U9645 (N_9645,N_9594,N_9493);
and U9646 (N_9646,N_9494,N_9513);
xnor U9647 (N_9647,N_9593,N_9556);
or U9648 (N_9648,N_9516,N_9479);
nor U9649 (N_9649,N_9596,N_9456);
and U9650 (N_9650,N_9446,N_9501);
xnor U9651 (N_9651,N_9444,N_9535);
or U9652 (N_9652,N_9486,N_9502);
nor U9653 (N_9653,N_9515,N_9569);
nor U9654 (N_9654,N_9584,N_9598);
xnor U9655 (N_9655,N_9485,N_9473);
or U9656 (N_9656,N_9511,N_9577);
nand U9657 (N_9657,N_9489,N_9480);
and U9658 (N_9658,N_9590,N_9546);
or U9659 (N_9659,N_9467,N_9550);
xnor U9660 (N_9660,N_9440,N_9495);
nand U9661 (N_9661,N_9552,N_9551);
nor U9662 (N_9662,N_9559,N_9441);
or U9663 (N_9663,N_9537,N_9524);
nor U9664 (N_9664,N_9530,N_9500);
nor U9665 (N_9665,N_9529,N_9583);
nor U9666 (N_9666,N_9470,N_9466);
nor U9667 (N_9667,N_9519,N_9471);
xor U9668 (N_9668,N_9457,N_9481);
or U9669 (N_9669,N_9566,N_9578);
xor U9670 (N_9670,N_9543,N_9575);
xnor U9671 (N_9671,N_9571,N_9548);
nand U9672 (N_9672,N_9588,N_9503);
or U9673 (N_9673,N_9518,N_9595);
or U9674 (N_9674,N_9520,N_9462);
xnor U9675 (N_9675,N_9541,N_9562);
xor U9676 (N_9676,N_9499,N_9491);
xnor U9677 (N_9677,N_9447,N_9581);
and U9678 (N_9678,N_9461,N_9540);
nand U9679 (N_9679,N_9463,N_9442);
xnor U9680 (N_9680,N_9585,N_9447);
and U9681 (N_9681,N_9445,N_9456);
and U9682 (N_9682,N_9574,N_9595);
nor U9683 (N_9683,N_9591,N_9530);
or U9684 (N_9684,N_9552,N_9485);
nor U9685 (N_9685,N_9582,N_9599);
xor U9686 (N_9686,N_9572,N_9560);
nand U9687 (N_9687,N_9458,N_9498);
or U9688 (N_9688,N_9476,N_9533);
and U9689 (N_9689,N_9550,N_9553);
nor U9690 (N_9690,N_9574,N_9498);
nand U9691 (N_9691,N_9564,N_9511);
nand U9692 (N_9692,N_9500,N_9540);
nor U9693 (N_9693,N_9516,N_9470);
or U9694 (N_9694,N_9558,N_9526);
nor U9695 (N_9695,N_9459,N_9576);
nand U9696 (N_9696,N_9520,N_9505);
nand U9697 (N_9697,N_9459,N_9527);
nand U9698 (N_9698,N_9466,N_9514);
and U9699 (N_9699,N_9464,N_9597);
nand U9700 (N_9700,N_9576,N_9524);
xnor U9701 (N_9701,N_9495,N_9508);
and U9702 (N_9702,N_9567,N_9490);
and U9703 (N_9703,N_9532,N_9477);
and U9704 (N_9704,N_9510,N_9487);
and U9705 (N_9705,N_9587,N_9502);
nor U9706 (N_9706,N_9490,N_9579);
nor U9707 (N_9707,N_9446,N_9492);
nand U9708 (N_9708,N_9562,N_9509);
xnor U9709 (N_9709,N_9523,N_9479);
or U9710 (N_9710,N_9544,N_9573);
nand U9711 (N_9711,N_9556,N_9596);
nand U9712 (N_9712,N_9513,N_9575);
nor U9713 (N_9713,N_9597,N_9456);
and U9714 (N_9714,N_9555,N_9516);
xnor U9715 (N_9715,N_9481,N_9492);
or U9716 (N_9716,N_9474,N_9483);
nor U9717 (N_9717,N_9531,N_9468);
xor U9718 (N_9718,N_9592,N_9468);
or U9719 (N_9719,N_9451,N_9526);
or U9720 (N_9720,N_9469,N_9513);
xnor U9721 (N_9721,N_9481,N_9511);
or U9722 (N_9722,N_9495,N_9507);
xnor U9723 (N_9723,N_9599,N_9587);
or U9724 (N_9724,N_9445,N_9523);
nand U9725 (N_9725,N_9473,N_9540);
or U9726 (N_9726,N_9591,N_9570);
xnor U9727 (N_9727,N_9478,N_9568);
or U9728 (N_9728,N_9532,N_9471);
nor U9729 (N_9729,N_9521,N_9522);
xor U9730 (N_9730,N_9463,N_9524);
or U9731 (N_9731,N_9579,N_9538);
nor U9732 (N_9732,N_9589,N_9488);
nand U9733 (N_9733,N_9491,N_9478);
or U9734 (N_9734,N_9515,N_9579);
nand U9735 (N_9735,N_9481,N_9515);
xor U9736 (N_9736,N_9586,N_9577);
xnor U9737 (N_9737,N_9588,N_9477);
nor U9738 (N_9738,N_9523,N_9484);
nand U9739 (N_9739,N_9590,N_9511);
nor U9740 (N_9740,N_9553,N_9447);
or U9741 (N_9741,N_9558,N_9447);
xnor U9742 (N_9742,N_9472,N_9552);
nor U9743 (N_9743,N_9448,N_9501);
nand U9744 (N_9744,N_9484,N_9469);
nand U9745 (N_9745,N_9507,N_9501);
nand U9746 (N_9746,N_9549,N_9536);
xor U9747 (N_9747,N_9522,N_9445);
nor U9748 (N_9748,N_9557,N_9553);
or U9749 (N_9749,N_9553,N_9455);
xor U9750 (N_9750,N_9504,N_9581);
xor U9751 (N_9751,N_9457,N_9551);
and U9752 (N_9752,N_9533,N_9450);
nand U9753 (N_9753,N_9462,N_9442);
or U9754 (N_9754,N_9456,N_9552);
or U9755 (N_9755,N_9469,N_9563);
nand U9756 (N_9756,N_9553,N_9507);
nand U9757 (N_9757,N_9553,N_9466);
and U9758 (N_9758,N_9473,N_9445);
and U9759 (N_9759,N_9596,N_9520);
nand U9760 (N_9760,N_9604,N_9627);
xor U9761 (N_9761,N_9730,N_9742);
and U9762 (N_9762,N_9620,N_9677);
nand U9763 (N_9763,N_9651,N_9618);
or U9764 (N_9764,N_9608,N_9704);
or U9765 (N_9765,N_9713,N_9706);
xor U9766 (N_9766,N_9645,N_9639);
and U9767 (N_9767,N_9626,N_9664);
and U9768 (N_9768,N_9747,N_9603);
nand U9769 (N_9769,N_9656,N_9633);
nand U9770 (N_9770,N_9754,N_9734);
or U9771 (N_9771,N_9668,N_9721);
xnor U9772 (N_9772,N_9748,N_9700);
nand U9773 (N_9773,N_9631,N_9741);
or U9774 (N_9774,N_9657,N_9684);
nand U9775 (N_9775,N_9649,N_9724);
nand U9776 (N_9776,N_9710,N_9723);
nor U9777 (N_9777,N_9628,N_9670);
nor U9778 (N_9778,N_9673,N_9735);
or U9779 (N_9779,N_9712,N_9680);
xnor U9780 (N_9780,N_9757,N_9634);
xor U9781 (N_9781,N_9717,N_9669);
nor U9782 (N_9782,N_9652,N_9701);
and U9783 (N_9783,N_9660,N_9722);
nand U9784 (N_9784,N_9600,N_9705);
xnor U9785 (N_9785,N_9688,N_9637);
nand U9786 (N_9786,N_9689,N_9648);
or U9787 (N_9787,N_9699,N_9753);
nor U9788 (N_9788,N_9672,N_9729);
nand U9789 (N_9789,N_9733,N_9725);
nand U9790 (N_9790,N_9715,N_9659);
and U9791 (N_9791,N_9638,N_9625);
nor U9792 (N_9792,N_9666,N_9610);
nand U9793 (N_9793,N_9607,N_9663);
or U9794 (N_9794,N_9644,N_9693);
xnor U9795 (N_9795,N_9726,N_9737);
or U9796 (N_9796,N_9685,N_9629);
xnor U9797 (N_9797,N_9690,N_9750);
xnor U9798 (N_9798,N_9630,N_9661);
nand U9799 (N_9799,N_9703,N_9727);
nand U9800 (N_9800,N_9681,N_9686);
or U9801 (N_9801,N_9653,N_9731);
nor U9802 (N_9802,N_9702,N_9635);
xnor U9803 (N_9803,N_9611,N_9697);
xnor U9804 (N_9804,N_9622,N_9759);
nand U9805 (N_9805,N_9636,N_9751);
and U9806 (N_9806,N_9728,N_9738);
and U9807 (N_9807,N_9758,N_9665);
and U9808 (N_9808,N_9691,N_9732);
xnor U9809 (N_9809,N_9740,N_9711);
and U9810 (N_9810,N_9707,N_9716);
and U9811 (N_9811,N_9667,N_9709);
nor U9812 (N_9812,N_9679,N_9617);
and U9813 (N_9813,N_9675,N_9708);
xnor U9814 (N_9814,N_9683,N_9719);
xor U9815 (N_9815,N_9739,N_9624);
xnor U9816 (N_9816,N_9743,N_9640);
xnor U9817 (N_9817,N_9605,N_9641);
and U9818 (N_9818,N_9650,N_9615);
or U9819 (N_9819,N_9692,N_9696);
nand U9820 (N_9820,N_9749,N_9642);
nor U9821 (N_9821,N_9643,N_9720);
and U9822 (N_9822,N_9674,N_9744);
and U9823 (N_9823,N_9745,N_9647);
nor U9824 (N_9824,N_9613,N_9718);
or U9825 (N_9825,N_9678,N_9682);
and U9826 (N_9826,N_9746,N_9655);
nand U9827 (N_9827,N_9714,N_9646);
nor U9828 (N_9828,N_9695,N_9601);
xnor U9829 (N_9829,N_9687,N_9756);
xor U9830 (N_9830,N_9694,N_9671);
or U9831 (N_9831,N_9621,N_9612);
xnor U9832 (N_9832,N_9755,N_9654);
or U9833 (N_9833,N_9632,N_9602);
xnor U9834 (N_9834,N_9614,N_9619);
and U9835 (N_9835,N_9623,N_9609);
and U9836 (N_9836,N_9658,N_9662);
xor U9837 (N_9837,N_9736,N_9616);
or U9838 (N_9838,N_9752,N_9676);
or U9839 (N_9839,N_9606,N_9698);
and U9840 (N_9840,N_9614,N_9740);
and U9841 (N_9841,N_9735,N_9705);
or U9842 (N_9842,N_9605,N_9642);
or U9843 (N_9843,N_9617,N_9683);
nand U9844 (N_9844,N_9736,N_9697);
and U9845 (N_9845,N_9613,N_9636);
and U9846 (N_9846,N_9746,N_9652);
nand U9847 (N_9847,N_9705,N_9633);
nand U9848 (N_9848,N_9647,N_9744);
and U9849 (N_9849,N_9720,N_9667);
nor U9850 (N_9850,N_9711,N_9668);
and U9851 (N_9851,N_9650,N_9754);
nand U9852 (N_9852,N_9721,N_9611);
nand U9853 (N_9853,N_9724,N_9672);
nand U9854 (N_9854,N_9658,N_9618);
xor U9855 (N_9855,N_9671,N_9652);
and U9856 (N_9856,N_9675,N_9700);
or U9857 (N_9857,N_9755,N_9677);
xor U9858 (N_9858,N_9673,N_9629);
xor U9859 (N_9859,N_9678,N_9647);
nand U9860 (N_9860,N_9735,N_9674);
nor U9861 (N_9861,N_9751,N_9725);
nand U9862 (N_9862,N_9738,N_9657);
xnor U9863 (N_9863,N_9726,N_9747);
or U9864 (N_9864,N_9736,N_9713);
or U9865 (N_9865,N_9721,N_9739);
and U9866 (N_9866,N_9623,N_9630);
and U9867 (N_9867,N_9637,N_9708);
nand U9868 (N_9868,N_9700,N_9721);
nand U9869 (N_9869,N_9604,N_9656);
xor U9870 (N_9870,N_9612,N_9715);
or U9871 (N_9871,N_9648,N_9712);
or U9872 (N_9872,N_9642,N_9705);
nand U9873 (N_9873,N_9674,N_9652);
nor U9874 (N_9874,N_9672,N_9677);
nand U9875 (N_9875,N_9705,N_9707);
nor U9876 (N_9876,N_9621,N_9689);
or U9877 (N_9877,N_9650,N_9729);
or U9878 (N_9878,N_9739,N_9748);
or U9879 (N_9879,N_9716,N_9626);
nor U9880 (N_9880,N_9699,N_9651);
xnor U9881 (N_9881,N_9607,N_9694);
xor U9882 (N_9882,N_9637,N_9654);
xor U9883 (N_9883,N_9726,N_9697);
nor U9884 (N_9884,N_9740,N_9695);
and U9885 (N_9885,N_9628,N_9734);
or U9886 (N_9886,N_9739,N_9710);
xnor U9887 (N_9887,N_9759,N_9670);
xnor U9888 (N_9888,N_9734,N_9616);
and U9889 (N_9889,N_9613,N_9729);
and U9890 (N_9890,N_9718,N_9697);
xor U9891 (N_9891,N_9665,N_9756);
nor U9892 (N_9892,N_9743,N_9705);
xnor U9893 (N_9893,N_9711,N_9738);
xnor U9894 (N_9894,N_9609,N_9757);
xnor U9895 (N_9895,N_9648,N_9609);
or U9896 (N_9896,N_9704,N_9727);
and U9897 (N_9897,N_9728,N_9614);
or U9898 (N_9898,N_9663,N_9660);
and U9899 (N_9899,N_9756,N_9711);
nand U9900 (N_9900,N_9673,N_9712);
nand U9901 (N_9901,N_9678,N_9676);
xnor U9902 (N_9902,N_9705,N_9627);
or U9903 (N_9903,N_9627,N_9702);
nor U9904 (N_9904,N_9699,N_9625);
nor U9905 (N_9905,N_9755,N_9730);
and U9906 (N_9906,N_9702,N_9738);
nor U9907 (N_9907,N_9732,N_9615);
nor U9908 (N_9908,N_9718,N_9682);
xor U9909 (N_9909,N_9748,N_9632);
nor U9910 (N_9910,N_9654,N_9649);
and U9911 (N_9911,N_9714,N_9696);
xor U9912 (N_9912,N_9721,N_9670);
or U9913 (N_9913,N_9726,N_9661);
nor U9914 (N_9914,N_9718,N_9629);
or U9915 (N_9915,N_9634,N_9643);
and U9916 (N_9916,N_9708,N_9679);
nor U9917 (N_9917,N_9680,N_9655);
and U9918 (N_9918,N_9717,N_9656);
nor U9919 (N_9919,N_9634,N_9691);
nand U9920 (N_9920,N_9885,N_9896);
or U9921 (N_9921,N_9897,N_9882);
or U9922 (N_9922,N_9784,N_9856);
or U9923 (N_9923,N_9809,N_9862);
nor U9924 (N_9924,N_9762,N_9813);
nor U9925 (N_9925,N_9889,N_9798);
or U9926 (N_9926,N_9841,N_9913);
or U9927 (N_9927,N_9845,N_9837);
xnor U9928 (N_9928,N_9779,N_9760);
xor U9929 (N_9929,N_9789,N_9768);
or U9930 (N_9930,N_9817,N_9905);
xnor U9931 (N_9931,N_9843,N_9761);
and U9932 (N_9932,N_9892,N_9820);
xor U9933 (N_9933,N_9829,N_9911);
nor U9934 (N_9934,N_9824,N_9791);
xnor U9935 (N_9935,N_9812,N_9888);
or U9936 (N_9936,N_9803,N_9800);
and U9937 (N_9937,N_9898,N_9873);
xnor U9938 (N_9938,N_9855,N_9783);
nand U9939 (N_9939,N_9894,N_9836);
nand U9940 (N_9940,N_9854,N_9786);
and U9941 (N_9941,N_9805,N_9793);
xnor U9942 (N_9942,N_9859,N_9877);
xor U9943 (N_9943,N_9828,N_9878);
xnor U9944 (N_9944,N_9775,N_9814);
and U9945 (N_9945,N_9808,N_9876);
xor U9946 (N_9946,N_9777,N_9880);
nand U9947 (N_9947,N_9868,N_9794);
or U9948 (N_9948,N_9899,N_9839);
nand U9949 (N_9949,N_9861,N_9884);
and U9950 (N_9950,N_9869,N_9860);
xor U9951 (N_9951,N_9858,N_9915);
and U9952 (N_9952,N_9830,N_9870);
nand U9953 (N_9953,N_9810,N_9823);
or U9954 (N_9954,N_9790,N_9827);
and U9955 (N_9955,N_9907,N_9846);
xnor U9956 (N_9956,N_9792,N_9785);
and U9957 (N_9957,N_9819,N_9893);
and U9958 (N_9958,N_9916,N_9776);
xnor U9959 (N_9959,N_9866,N_9788);
nor U9960 (N_9960,N_9804,N_9795);
nand U9961 (N_9961,N_9909,N_9879);
and U9962 (N_9962,N_9887,N_9796);
nor U9963 (N_9963,N_9815,N_9811);
nor U9964 (N_9964,N_9857,N_9891);
and U9965 (N_9965,N_9765,N_9881);
nand U9966 (N_9966,N_9833,N_9801);
and U9967 (N_9967,N_9764,N_9781);
and U9968 (N_9968,N_9919,N_9852);
and U9969 (N_9969,N_9842,N_9902);
nor U9970 (N_9970,N_9863,N_9770);
nor U9971 (N_9971,N_9825,N_9780);
or U9972 (N_9972,N_9797,N_9912);
and U9973 (N_9973,N_9838,N_9848);
nand U9974 (N_9974,N_9872,N_9900);
nor U9975 (N_9975,N_9883,N_9840);
or U9976 (N_9976,N_9903,N_9895);
nor U9977 (N_9977,N_9763,N_9864);
xor U9978 (N_9978,N_9910,N_9871);
xnor U9979 (N_9979,N_9832,N_9782);
and U9980 (N_9980,N_9914,N_9875);
nand U9981 (N_9981,N_9807,N_9917);
and U9982 (N_9982,N_9799,N_9806);
nor U9983 (N_9983,N_9865,N_9906);
xor U9984 (N_9984,N_9835,N_9834);
nand U9985 (N_9985,N_9847,N_9904);
or U9986 (N_9986,N_9908,N_9767);
xnor U9987 (N_9987,N_9774,N_9851);
xnor U9988 (N_9988,N_9918,N_9874);
nor U9989 (N_9989,N_9853,N_9849);
xor U9990 (N_9990,N_9850,N_9773);
nor U9991 (N_9991,N_9890,N_9831);
xnor U9992 (N_9992,N_9802,N_9769);
nor U9993 (N_9993,N_9816,N_9766);
nand U9994 (N_9994,N_9778,N_9787);
nand U9995 (N_9995,N_9867,N_9772);
or U9996 (N_9996,N_9822,N_9818);
nor U9997 (N_9997,N_9886,N_9821);
or U9998 (N_9998,N_9826,N_9844);
xor U9999 (N_9999,N_9901,N_9771);
and U10000 (N_10000,N_9905,N_9814);
nand U10001 (N_10001,N_9916,N_9785);
nand U10002 (N_10002,N_9793,N_9780);
nand U10003 (N_10003,N_9881,N_9913);
xnor U10004 (N_10004,N_9898,N_9833);
nor U10005 (N_10005,N_9770,N_9913);
xor U10006 (N_10006,N_9801,N_9823);
and U10007 (N_10007,N_9849,N_9761);
nand U10008 (N_10008,N_9819,N_9888);
nand U10009 (N_10009,N_9868,N_9774);
nand U10010 (N_10010,N_9915,N_9825);
or U10011 (N_10011,N_9905,N_9804);
nor U10012 (N_10012,N_9828,N_9900);
xnor U10013 (N_10013,N_9796,N_9914);
or U10014 (N_10014,N_9767,N_9816);
nor U10015 (N_10015,N_9843,N_9917);
xor U10016 (N_10016,N_9876,N_9864);
nand U10017 (N_10017,N_9895,N_9850);
nand U10018 (N_10018,N_9906,N_9795);
xnor U10019 (N_10019,N_9915,N_9822);
nor U10020 (N_10020,N_9844,N_9764);
nand U10021 (N_10021,N_9846,N_9838);
nand U10022 (N_10022,N_9789,N_9868);
or U10023 (N_10023,N_9873,N_9852);
nand U10024 (N_10024,N_9914,N_9806);
nor U10025 (N_10025,N_9858,N_9776);
nor U10026 (N_10026,N_9838,N_9888);
xor U10027 (N_10027,N_9807,N_9883);
or U10028 (N_10028,N_9785,N_9910);
nor U10029 (N_10029,N_9798,N_9918);
nor U10030 (N_10030,N_9873,N_9811);
nand U10031 (N_10031,N_9772,N_9836);
nor U10032 (N_10032,N_9916,N_9900);
nand U10033 (N_10033,N_9915,N_9889);
and U10034 (N_10034,N_9783,N_9836);
nand U10035 (N_10035,N_9762,N_9877);
and U10036 (N_10036,N_9863,N_9825);
nand U10037 (N_10037,N_9820,N_9809);
and U10038 (N_10038,N_9797,N_9878);
nand U10039 (N_10039,N_9810,N_9892);
xnor U10040 (N_10040,N_9831,N_9909);
nor U10041 (N_10041,N_9883,N_9882);
or U10042 (N_10042,N_9852,N_9846);
xnor U10043 (N_10043,N_9873,N_9772);
nand U10044 (N_10044,N_9833,N_9774);
xnor U10045 (N_10045,N_9763,N_9848);
and U10046 (N_10046,N_9825,N_9794);
and U10047 (N_10047,N_9823,N_9776);
nand U10048 (N_10048,N_9800,N_9787);
or U10049 (N_10049,N_9833,N_9857);
or U10050 (N_10050,N_9776,N_9784);
and U10051 (N_10051,N_9792,N_9859);
or U10052 (N_10052,N_9894,N_9893);
or U10053 (N_10053,N_9817,N_9846);
nand U10054 (N_10054,N_9876,N_9891);
and U10055 (N_10055,N_9845,N_9839);
nand U10056 (N_10056,N_9918,N_9845);
xor U10057 (N_10057,N_9858,N_9762);
nor U10058 (N_10058,N_9915,N_9783);
nor U10059 (N_10059,N_9781,N_9847);
or U10060 (N_10060,N_9909,N_9888);
and U10061 (N_10061,N_9918,N_9776);
nand U10062 (N_10062,N_9904,N_9864);
nand U10063 (N_10063,N_9903,N_9918);
nor U10064 (N_10064,N_9847,N_9878);
xor U10065 (N_10065,N_9832,N_9763);
and U10066 (N_10066,N_9786,N_9767);
or U10067 (N_10067,N_9894,N_9834);
nor U10068 (N_10068,N_9830,N_9856);
and U10069 (N_10069,N_9849,N_9769);
or U10070 (N_10070,N_9910,N_9781);
and U10071 (N_10071,N_9906,N_9855);
or U10072 (N_10072,N_9799,N_9855);
or U10073 (N_10073,N_9866,N_9865);
or U10074 (N_10074,N_9835,N_9827);
nand U10075 (N_10075,N_9842,N_9870);
and U10076 (N_10076,N_9913,N_9789);
and U10077 (N_10077,N_9845,N_9768);
xnor U10078 (N_10078,N_9793,N_9862);
and U10079 (N_10079,N_9812,N_9826);
and U10080 (N_10080,N_9960,N_10013);
xnor U10081 (N_10081,N_10030,N_10019);
nor U10082 (N_10082,N_10023,N_9986);
and U10083 (N_10083,N_9938,N_10018);
or U10084 (N_10084,N_10020,N_10050);
nand U10085 (N_10085,N_10028,N_10016);
or U10086 (N_10086,N_10044,N_9925);
xor U10087 (N_10087,N_9988,N_9963);
and U10088 (N_10088,N_9921,N_9980);
nor U10089 (N_10089,N_10055,N_10042);
nand U10090 (N_10090,N_9977,N_10054);
nor U10091 (N_10091,N_10072,N_9924);
or U10092 (N_10092,N_10032,N_9984);
nand U10093 (N_10093,N_9927,N_9949);
or U10094 (N_10094,N_10043,N_10068);
nand U10095 (N_10095,N_9941,N_10078);
or U10096 (N_10096,N_10006,N_9934);
or U10097 (N_10097,N_9944,N_9976);
nand U10098 (N_10098,N_9951,N_9936);
nand U10099 (N_10099,N_10041,N_9952);
nand U10100 (N_10100,N_10004,N_10024);
nor U10101 (N_10101,N_10035,N_9994);
nand U10102 (N_10102,N_9970,N_9968);
or U10103 (N_10103,N_9945,N_10056);
and U10104 (N_10104,N_9962,N_10046);
xnor U10105 (N_10105,N_9943,N_9932);
or U10106 (N_10106,N_9981,N_10075);
or U10107 (N_10107,N_9955,N_10001);
nor U10108 (N_10108,N_9990,N_10034);
and U10109 (N_10109,N_10037,N_9978);
and U10110 (N_10110,N_9957,N_9935);
nor U10111 (N_10111,N_10015,N_9964);
or U10112 (N_10112,N_10059,N_9965);
nor U10113 (N_10113,N_9923,N_9939);
nor U10114 (N_10114,N_10073,N_9983);
xor U10115 (N_10115,N_9928,N_9999);
or U10116 (N_10116,N_9953,N_9996);
or U10117 (N_10117,N_9940,N_10045);
and U10118 (N_10118,N_10011,N_10036);
nor U10119 (N_10119,N_9974,N_10014);
xor U10120 (N_10120,N_10077,N_9997);
nand U10121 (N_10121,N_9979,N_10010);
nand U10122 (N_10122,N_9971,N_9966);
xnor U10123 (N_10123,N_9989,N_10038);
or U10124 (N_10124,N_10065,N_10017);
nand U10125 (N_10125,N_9975,N_9958);
xor U10126 (N_10126,N_9937,N_10025);
nand U10127 (N_10127,N_9929,N_9992);
and U10128 (N_10128,N_10058,N_9982);
or U10129 (N_10129,N_10079,N_10039);
nor U10130 (N_10130,N_10052,N_10005);
or U10131 (N_10131,N_10029,N_10064);
xor U10132 (N_10132,N_10026,N_9922);
xor U10133 (N_10133,N_10000,N_10067);
or U10134 (N_10134,N_10048,N_9930);
and U10135 (N_10135,N_9998,N_9956);
xor U10136 (N_10136,N_9946,N_9947);
nor U10137 (N_10137,N_9920,N_9926);
nor U10138 (N_10138,N_9972,N_10053);
nand U10139 (N_10139,N_10040,N_10033);
xnor U10140 (N_10140,N_10069,N_10071);
nor U10141 (N_10141,N_9959,N_10008);
xor U10142 (N_10142,N_9987,N_10007);
xor U10143 (N_10143,N_10051,N_10070);
and U10144 (N_10144,N_10002,N_9931);
xor U10145 (N_10145,N_10009,N_10031);
xnor U10146 (N_10146,N_10062,N_10049);
or U10147 (N_10147,N_9933,N_10021);
nor U10148 (N_10148,N_9954,N_9942);
or U10149 (N_10149,N_10022,N_10047);
nand U10150 (N_10150,N_10066,N_9985);
nor U10151 (N_10151,N_10061,N_10060);
and U10152 (N_10152,N_9995,N_9950);
and U10153 (N_10153,N_9967,N_10074);
and U10154 (N_10154,N_10003,N_10012);
nand U10155 (N_10155,N_10027,N_10057);
and U10156 (N_10156,N_9991,N_9973);
or U10157 (N_10157,N_9961,N_10076);
xnor U10158 (N_10158,N_9948,N_9993);
nand U10159 (N_10159,N_10063,N_9969);
or U10160 (N_10160,N_10006,N_10054);
nand U10161 (N_10161,N_9959,N_10057);
and U10162 (N_10162,N_10079,N_10040);
xor U10163 (N_10163,N_10022,N_10042);
and U10164 (N_10164,N_9988,N_9927);
and U10165 (N_10165,N_9945,N_9949);
nand U10166 (N_10166,N_9990,N_9955);
or U10167 (N_10167,N_10056,N_10037);
nand U10168 (N_10168,N_9926,N_9976);
nand U10169 (N_10169,N_9990,N_10039);
or U10170 (N_10170,N_10004,N_9983);
or U10171 (N_10171,N_10041,N_10065);
or U10172 (N_10172,N_10000,N_10041);
nor U10173 (N_10173,N_10004,N_10076);
nand U10174 (N_10174,N_10017,N_10026);
or U10175 (N_10175,N_10047,N_10006);
xnor U10176 (N_10176,N_10069,N_10032);
xnor U10177 (N_10177,N_10008,N_10024);
or U10178 (N_10178,N_9942,N_9989);
nand U10179 (N_10179,N_9936,N_9962);
nand U10180 (N_10180,N_9954,N_10052);
xnor U10181 (N_10181,N_9960,N_9975);
xnor U10182 (N_10182,N_9975,N_9970);
nand U10183 (N_10183,N_10028,N_10056);
or U10184 (N_10184,N_9967,N_9969);
xnor U10185 (N_10185,N_10005,N_10064);
nand U10186 (N_10186,N_9967,N_9930);
nor U10187 (N_10187,N_9990,N_10073);
nor U10188 (N_10188,N_10023,N_9944);
nand U10189 (N_10189,N_10076,N_9947);
xnor U10190 (N_10190,N_10057,N_9950);
nor U10191 (N_10191,N_10029,N_9939);
and U10192 (N_10192,N_9934,N_9925);
xor U10193 (N_10193,N_9992,N_10007);
nor U10194 (N_10194,N_9936,N_9943);
xnor U10195 (N_10195,N_9966,N_9926);
xor U10196 (N_10196,N_10069,N_9960);
or U10197 (N_10197,N_10036,N_10030);
or U10198 (N_10198,N_9989,N_10053);
nor U10199 (N_10199,N_9923,N_10035);
nand U10200 (N_10200,N_9986,N_10076);
nand U10201 (N_10201,N_10012,N_9948);
nor U10202 (N_10202,N_10074,N_9939);
nand U10203 (N_10203,N_9953,N_9940);
and U10204 (N_10204,N_9989,N_10058);
nand U10205 (N_10205,N_9952,N_9942);
nand U10206 (N_10206,N_9935,N_10053);
nand U10207 (N_10207,N_9974,N_9977);
xnor U10208 (N_10208,N_10062,N_10066);
xor U10209 (N_10209,N_9930,N_9925);
nor U10210 (N_10210,N_9978,N_9981);
or U10211 (N_10211,N_9998,N_9933);
or U10212 (N_10212,N_9958,N_10015);
nand U10213 (N_10213,N_9925,N_9973);
or U10214 (N_10214,N_9935,N_10042);
nand U10215 (N_10215,N_10058,N_10036);
nor U10216 (N_10216,N_9925,N_10074);
and U10217 (N_10217,N_9945,N_9985);
nand U10218 (N_10218,N_9964,N_10020);
xnor U10219 (N_10219,N_9984,N_9954);
or U10220 (N_10220,N_9997,N_9974);
xor U10221 (N_10221,N_10033,N_10029);
nand U10222 (N_10222,N_10021,N_9956);
and U10223 (N_10223,N_10023,N_10010);
xor U10224 (N_10224,N_10026,N_10037);
nor U10225 (N_10225,N_9935,N_9960);
and U10226 (N_10226,N_9949,N_9960);
xnor U10227 (N_10227,N_10065,N_10011);
xnor U10228 (N_10228,N_9972,N_9955);
or U10229 (N_10229,N_9960,N_10022);
and U10230 (N_10230,N_10024,N_10018);
and U10231 (N_10231,N_9966,N_10019);
nand U10232 (N_10232,N_9992,N_9998);
xor U10233 (N_10233,N_10047,N_10018);
nand U10234 (N_10234,N_9936,N_10052);
xnor U10235 (N_10235,N_10007,N_10026);
and U10236 (N_10236,N_9962,N_10055);
and U10237 (N_10237,N_10009,N_9956);
xnor U10238 (N_10238,N_9968,N_9946);
xnor U10239 (N_10239,N_9952,N_9947);
or U10240 (N_10240,N_10126,N_10142);
or U10241 (N_10241,N_10085,N_10103);
nand U10242 (N_10242,N_10211,N_10117);
nand U10243 (N_10243,N_10159,N_10167);
or U10244 (N_10244,N_10146,N_10200);
nand U10245 (N_10245,N_10172,N_10083);
and U10246 (N_10246,N_10107,N_10082);
nand U10247 (N_10247,N_10180,N_10130);
nor U10248 (N_10248,N_10101,N_10080);
nor U10249 (N_10249,N_10204,N_10164);
and U10250 (N_10250,N_10136,N_10230);
nor U10251 (N_10251,N_10148,N_10187);
or U10252 (N_10252,N_10210,N_10218);
xor U10253 (N_10253,N_10095,N_10150);
nand U10254 (N_10254,N_10115,N_10223);
or U10255 (N_10255,N_10125,N_10176);
and U10256 (N_10256,N_10089,N_10081);
nor U10257 (N_10257,N_10151,N_10161);
xnor U10258 (N_10258,N_10197,N_10145);
or U10259 (N_10259,N_10198,N_10179);
nand U10260 (N_10260,N_10238,N_10157);
or U10261 (N_10261,N_10122,N_10124);
nor U10262 (N_10262,N_10165,N_10141);
nand U10263 (N_10263,N_10096,N_10154);
xor U10264 (N_10264,N_10129,N_10111);
nor U10265 (N_10265,N_10227,N_10114);
xor U10266 (N_10266,N_10087,N_10175);
nand U10267 (N_10267,N_10160,N_10086);
or U10268 (N_10268,N_10168,N_10118);
and U10269 (N_10269,N_10215,N_10216);
and U10270 (N_10270,N_10104,N_10193);
nor U10271 (N_10271,N_10110,N_10162);
or U10272 (N_10272,N_10237,N_10133);
or U10273 (N_10273,N_10173,N_10090);
and U10274 (N_10274,N_10236,N_10171);
nor U10275 (N_10275,N_10220,N_10178);
xor U10276 (N_10276,N_10144,N_10093);
xor U10277 (N_10277,N_10135,N_10099);
nor U10278 (N_10278,N_10208,N_10155);
nor U10279 (N_10279,N_10232,N_10112);
nor U10280 (N_10280,N_10094,N_10152);
nor U10281 (N_10281,N_10098,N_10108);
and U10282 (N_10282,N_10105,N_10182);
nor U10283 (N_10283,N_10209,N_10132);
nor U10284 (N_10284,N_10183,N_10192);
xnor U10285 (N_10285,N_10234,N_10127);
xor U10286 (N_10286,N_10194,N_10225);
nand U10287 (N_10287,N_10185,N_10239);
nand U10288 (N_10288,N_10226,N_10158);
nor U10289 (N_10289,N_10143,N_10088);
and U10290 (N_10290,N_10131,N_10134);
and U10291 (N_10291,N_10100,N_10106);
nor U10292 (N_10292,N_10181,N_10217);
nor U10293 (N_10293,N_10221,N_10189);
or U10294 (N_10294,N_10229,N_10137);
nor U10295 (N_10295,N_10196,N_10199);
xnor U10296 (N_10296,N_10119,N_10233);
and U10297 (N_10297,N_10166,N_10205);
and U10298 (N_10298,N_10121,N_10203);
xnor U10299 (N_10299,N_10228,N_10156);
or U10300 (N_10300,N_10092,N_10091);
xor U10301 (N_10301,N_10214,N_10202);
or U10302 (N_10302,N_10174,N_10097);
or U10303 (N_10303,N_10170,N_10120);
nand U10304 (N_10304,N_10149,N_10184);
or U10305 (N_10305,N_10102,N_10109);
nor U10306 (N_10306,N_10219,N_10222);
or U10307 (N_10307,N_10169,N_10224);
nor U10308 (N_10308,N_10138,N_10186);
nor U10309 (N_10309,N_10147,N_10212);
nand U10310 (N_10310,N_10191,N_10188);
and U10311 (N_10311,N_10206,N_10213);
or U10312 (N_10312,N_10207,N_10201);
and U10313 (N_10313,N_10235,N_10113);
nand U10314 (N_10314,N_10163,N_10195);
nor U10315 (N_10315,N_10140,N_10177);
nand U10316 (N_10316,N_10139,N_10190);
nand U10317 (N_10317,N_10123,N_10116);
xor U10318 (N_10318,N_10153,N_10231);
nand U10319 (N_10319,N_10084,N_10128);
and U10320 (N_10320,N_10126,N_10160);
nand U10321 (N_10321,N_10090,N_10127);
nor U10322 (N_10322,N_10082,N_10225);
xnor U10323 (N_10323,N_10175,N_10095);
nor U10324 (N_10324,N_10145,N_10090);
nand U10325 (N_10325,N_10146,N_10214);
xor U10326 (N_10326,N_10193,N_10091);
or U10327 (N_10327,N_10163,N_10150);
or U10328 (N_10328,N_10222,N_10239);
nand U10329 (N_10329,N_10113,N_10142);
xor U10330 (N_10330,N_10224,N_10125);
and U10331 (N_10331,N_10216,N_10158);
xnor U10332 (N_10332,N_10106,N_10090);
nand U10333 (N_10333,N_10218,N_10123);
and U10334 (N_10334,N_10145,N_10114);
nand U10335 (N_10335,N_10104,N_10100);
and U10336 (N_10336,N_10119,N_10103);
or U10337 (N_10337,N_10194,N_10199);
nand U10338 (N_10338,N_10221,N_10137);
and U10339 (N_10339,N_10129,N_10151);
nand U10340 (N_10340,N_10232,N_10083);
xor U10341 (N_10341,N_10157,N_10142);
nand U10342 (N_10342,N_10201,N_10187);
and U10343 (N_10343,N_10197,N_10122);
or U10344 (N_10344,N_10211,N_10122);
nand U10345 (N_10345,N_10189,N_10131);
or U10346 (N_10346,N_10109,N_10235);
or U10347 (N_10347,N_10106,N_10168);
nand U10348 (N_10348,N_10103,N_10186);
or U10349 (N_10349,N_10228,N_10163);
or U10350 (N_10350,N_10229,N_10207);
and U10351 (N_10351,N_10099,N_10211);
nor U10352 (N_10352,N_10185,N_10224);
or U10353 (N_10353,N_10104,N_10230);
and U10354 (N_10354,N_10104,N_10099);
xor U10355 (N_10355,N_10080,N_10095);
xor U10356 (N_10356,N_10190,N_10083);
and U10357 (N_10357,N_10081,N_10156);
nor U10358 (N_10358,N_10224,N_10154);
or U10359 (N_10359,N_10167,N_10215);
or U10360 (N_10360,N_10148,N_10095);
xor U10361 (N_10361,N_10099,N_10144);
nand U10362 (N_10362,N_10094,N_10111);
xor U10363 (N_10363,N_10168,N_10115);
or U10364 (N_10364,N_10134,N_10184);
xnor U10365 (N_10365,N_10113,N_10093);
nand U10366 (N_10366,N_10197,N_10220);
or U10367 (N_10367,N_10108,N_10228);
and U10368 (N_10368,N_10128,N_10098);
nand U10369 (N_10369,N_10203,N_10198);
and U10370 (N_10370,N_10161,N_10228);
or U10371 (N_10371,N_10166,N_10096);
nand U10372 (N_10372,N_10189,N_10178);
or U10373 (N_10373,N_10172,N_10190);
or U10374 (N_10374,N_10118,N_10159);
or U10375 (N_10375,N_10134,N_10188);
and U10376 (N_10376,N_10233,N_10206);
and U10377 (N_10377,N_10237,N_10160);
nand U10378 (N_10378,N_10117,N_10090);
nand U10379 (N_10379,N_10121,N_10149);
or U10380 (N_10380,N_10183,N_10165);
and U10381 (N_10381,N_10196,N_10225);
xnor U10382 (N_10382,N_10095,N_10170);
xor U10383 (N_10383,N_10199,N_10083);
nor U10384 (N_10384,N_10239,N_10157);
nand U10385 (N_10385,N_10112,N_10149);
nor U10386 (N_10386,N_10108,N_10209);
xnor U10387 (N_10387,N_10084,N_10232);
xnor U10388 (N_10388,N_10226,N_10149);
and U10389 (N_10389,N_10145,N_10122);
and U10390 (N_10390,N_10165,N_10081);
and U10391 (N_10391,N_10196,N_10137);
xnor U10392 (N_10392,N_10204,N_10219);
xor U10393 (N_10393,N_10207,N_10105);
xnor U10394 (N_10394,N_10139,N_10230);
xnor U10395 (N_10395,N_10085,N_10235);
and U10396 (N_10396,N_10176,N_10181);
xnor U10397 (N_10397,N_10090,N_10186);
and U10398 (N_10398,N_10103,N_10107);
nor U10399 (N_10399,N_10197,N_10091);
and U10400 (N_10400,N_10395,N_10249);
nand U10401 (N_10401,N_10348,N_10336);
nand U10402 (N_10402,N_10298,N_10359);
nand U10403 (N_10403,N_10372,N_10253);
or U10404 (N_10404,N_10251,N_10399);
and U10405 (N_10405,N_10296,N_10278);
and U10406 (N_10406,N_10271,N_10355);
and U10407 (N_10407,N_10288,N_10293);
and U10408 (N_10408,N_10259,N_10285);
nor U10409 (N_10409,N_10264,N_10313);
nand U10410 (N_10410,N_10290,N_10316);
nor U10411 (N_10411,N_10341,N_10283);
xnor U10412 (N_10412,N_10242,N_10369);
nand U10413 (N_10413,N_10273,N_10319);
and U10414 (N_10414,N_10324,N_10277);
nand U10415 (N_10415,N_10361,N_10310);
nand U10416 (N_10416,N_10276,N_10292);
nand U10417 (N_10417,N_10279,N_10309);
xnor U10418 (N_10418,N_10389,N_10246);
xnor U10419 (N_10419,N_10392,N_10267);
or U10420 (N_10420,N_10280,N_10304);
nand U10421 (N_10421,N_10344,N_10388);
nor U10422 (N_10422,N_10254,N_10243);
or U10423 (N_10423,N_10294,N_10373);
or U10424 (N_10424,N_10262,N_10332);
and U10425 (N_10425,N_10323,N_10260);
and U10426 (N_10426,N_10358,N_10295);
nor U10427 (N_10427,N_10274,N_10393);
xnor U10428 (N_10428,N_10345,N_10378);
and U10429 (N_10429,N_10370,N_10318);
xnor U10430 (N_10430,N_10360,N_10391);
nand U10431 (N_10431,N_10380,N_10287);
nand U10432 (N_10432,N_10347,N_10351);
nor U10433 (N_10433,N_10275,N_10320);
nor U10434 (N_10434,N_10303,N_10301);
or U10435 (N_10435,N_10248,N_10329);
nor U10436 (N_10436,N_10289,N_10334);
nand U10437 (N_10437,N_10371,N_10382);
nor U10438 (N_10438,N_10256,N_10314);
nor U10439 (N_10439,N_10317,N_10270);
xnor U10440 (N_10440,N_10349,N_10321);
nand U10441 (N_10441,N_10250,N_10308);
xor U10442 (N_10442,N_10241,N_10396);
nor U10443 (N_10443,N_10247,N_10357);
xnor U10444 (N_10444,N_10255,N_10365);
and U10445 (N_10445,N_10268,N_10387);
nand U10446 (N_10446,N_10331,N_10311);
nand U10447 (N_10447,N_10266,N_10379);
xnor U10448 (N_10448,N_10328,N_10252);
and U10449 (N_10449,N_10272,N_10281);
nand U10450 (N_10450,N_10383,N_10269);
nor U10451 (N_10451,N_10377,N_10245);
nor U10452 (N_10452,N_10265,N_10297);
nor U10453 (N_10453,N_10305,N_10300);
or U10454 (N_10454,N_10327,N_10325);
xor U10455 (N_10455,N_10367,N_10335);
or U10456 (N_10456,N_10330,N_10362);
nor U10457 (N_10457,N_10354,N_10315);
nand U10458 (N_10458,N_10394,N_10390);
nand U10459 (N_10459,N_10397,N_10261);
and U10460 (N_10460,N_10384,N_10291);
or U10461 (N_10461,N_10374,N_10333);
and U10462 (N_10462,N_10381,N_10263);
nand U10463 (N_10463,N_10352,N_10353);
xor U10464 (N_10464,N_10340,N_10363);
or U10465 (N_10465,N_10385,N_10299);
or U10466 (N_10466,N_10343,N_10375);
and U10467 (N_10467,N_10244,N_10398);
and U10468 (N_10468,N_10306,N_10326);
nand U10469 (N_10469,N_10282,N_10346);
and U10470 (N_10470,N_10322,N_10240);
xnor U10471 (N_10471,N_10302,N_10350);
nor U10472 (N_10472,N_10258,N_10368);
nand U10473 (N_10473,N_10386,N_10338);
xor U10474 (N_10474,N_10312,N_10339);
nor U10475 (N_10475,N_10286,N_10307);
and U10476 (N_10476,N_10364,N_10342);
xor U10477 (N_10477,N_10376,N_10257);
nor U10478 (N_10478,N_10284,N_10356);
nand U10479 (N_10479,N_10337,N_10366);
and U10480 (N_10480,N_10394,N_10352);
or U10481 (N_10481,N_10359,N_10338);
xor U10482 (N_10482,N_10314,N_10281);
nand U10483 (N_10483,N_10298,N_10290);
and U10484 (N_10484,N_10328,N_10347);
or U10485 (N_10485,N_10356,N_10288);
or U10486 (N_10486,N_10253,N_10319);
nor U10487 (N_10487,N_10294,N_10320);
xnor U10488 (N_10488,N_10360,N_10387);
nand U10489 (N_10489,N_10352,N_10317);
nor U10490 (N_10490,N_10245,N_10383);
and U10491 (N_10491,N_10354,N_10382);
or U10492 (N_10492,N_10359,N_10345);
and U10493 (N_10493,N_10317,N_10280);
and U10494 (N_10494,N_10255,N_10359);
xnor U10495 (N_10495,N_10247,N_10375);
nor U10496 (N_10496,N_10322,N_10376);
nor U10497 (N_10497,N_10366,N_10368);
or U10498 (N_10498,N_10316,N_10327);
nand U10499 (N_10499,N_10246,N_10299);
xnor U10500 (N_10500,N_10282,N_10270);
nor U10501 (N_10501,N_10274,N_10290);
and U10502 (N_10502,N_10266,N_10324);
nand U10503 (N_10503,N_10361,N_10259);
xnor U10504 (N_10504,N_10259,N_10255);
and U10505 (N_10505,N_10263,N_10294);
nand U10506 (N_10506,N_10274,N_10253);
nand U10507 (N_10507,N_10337,N_10274);
or U10508 (N_10508,N_10399,N_10290);
and U10509 (N_10509,N_10268,N_10254);
xnor U10510 (N_10510,N_10256,N_10371);
xnor U10511 (N_10511,N_10253,N_10366);
or U10512 (N_10512,N_10254,N_10318);
or U10513 (N_10513,N_10377,N_10298);
nand U10514 (N_10514,N_10346,N_10392);
nand U10515 (N_10515,N_10356,N_10334);
nor U10516 (N_10516,N_10243,N_10339);
and U10517 (N_10517,N_10359,N_10377);
or U10518 (N_10518,N_10326,N_10321);
nor U10519 (N_10519,N_10342,N_10247);
xnor U10520 (N_10520,N_10385,N_10283);
nand U10521 (N_10521,N_10341,N_10285);
xnor U10522 (N_10522,N_10254,N_10341);
and U10523 (N_10523,N_10344,N_10263);
or U10524 (N_10524,N_10318,N_10292);
nor U10525 (N_10525,N_10387,N_10330);
or U10526 (N_10526,N_10356,N_10279);
or U10527 (N_10527,N_10355,N_10391);
xnor U10528 (N_10528,N_10341,N_10314);
xnor U10529 (N_10529,N_10317,N_10243);
nor U10530 (N_10530,N_10290,N_10269);
xnor U10531 (N_10531,N_10360,N_10363);
nand U10532 (N_10532,N_10262,N_10320);
nand U10533 (N_10533,N_10371,N_10307);
or U10534 (N_10534,N_10357,N_10334);
nand U10535 (N_10535,N_10335,N_10388);
nand U10536 (N_10536,N_10314,N_10299);
and U10537 (N_10537,N_10267,N_10370);
and U10538 (N_10538,N_10345,N_10287);
or U10539 (N_10539,N_10269,N_10393);
nand U10540 (N_10540,N_10248,N_10295);
or U10541 (N_10541,N_10338,N_10364);
xnor U10542 (N_10542,N_10346,N_10286);
xnor U10543 (N_10543,N_10261,N_10270);
and U10544 (N_10544,N_10367,N_10257);
nor U10545 (N_10545,N_10307,N_10301);
nand U10546 (N_10546,N_10389,N_10384);
or U10547 (N_10547,N_10290,N_10321);
or U10548 (N_10548,N_10388,N_10346);
xor U10549 (N_10549,N_10307,N_10380);
nand U10550 (N_10550,N_10290,N_10360);
nor U10551 (N_10551,N_10352,N_10290);
nand U10552 (N_10552,N_10347,N_10242);
and U10553 (N_10553,N_10382,N_10284);
nand U10554 (N_10554,N_10256,N_10398);
nor U10555 (N_10555,N_10350,N_10328);
or U10556 (N_10556,N_10338,N_10293);
nand U10557 (N_10557,N_10272,N_10378);
xor U10558 (N_10558,N_10349,N_10267);
or U10559 (N_10559,N_10277,N_10290);
and U10560 (N_10560,N_10518,N_10421);
and U10561 (N_10561,N_10532,N_10435);
nand U10562 (N_10562,N_10449,N_10539);
xnor U10563 (N_10563,N_10450,N_10445);
nand U10564 (N_10564,N_10550,N_10515);
nor U10565 (N_10565,N_10436,N_10499);
and U10566 (N_10566,N_10426,N_10545);
or U10567 (N_10567,N_10433,N_10519);
and U10568 (N_10568,N_10520,N_10521);
and U10569 (N_10569,N_10488,N_10505);
nor U10570 (N_10570,N_10552,N_10412);
nand U10571 (N_10571,N_10479,N_10454);
and U10572 (N_10572,N_10418,N_10405);
nor U10573 (N_10573,N_10459,N_10487);
and U10574 (N_10574,N_10528,N_10540);
xor U10575 (N_10575,N_10489,N_10456);
and U10576 (N_10576,N_10547,N_10525);
xor U10577 (N_10577,N_10441,N_10512);
xnor U10578 (N_10578,N_10478,N_10482);
xor U10579 (N_10579,N_10473,N_10500);
xnor U10580 (N_10580,N_10542,N_10442);
xor U10581 (N_10581,N_10472,N_10413);
nor U10582 (N_10582,N_10486,N_10533);
nor U10583 (N_10583,N_10553,N_10534);
and U10584 (N_10584,N_10530,N_10496);
and U10585 (N_10585,N_10529,N_10419);
nand U10586 (N_10586,N_10506,N_10440);
nor U10587 (N_10587,N_10497,N_10546);
or U10588 (N_10588,N_10493,N_10471);
xnor U10589 (N_10589,N_10531,N_10402);
and U10590 (N_10590,N_10463,N_10406);
and U10591 (N_10591,N_10424,N_10514);
nand U10592 (N_10592,N_10536,N_10523);
xnor U10593 (N_10593,N_10467,N_10522);
or U10594 (N_10594,N_10470,N_10510);
or U10595 (N_10595,N_10416,N_10404);
nor U10596 (N_10596,N_10554,N_10485);
and U10597 (N_10597,N_10508,N_10556);
xor U10598 (N_10598,N_10446,N_10495);
nor U10599 (N_10599,N_10464,N_10502);
xnor U10600 (N_10600,N_10503,N_10403);
or U10601 (N_10601,N_10535,N_10455);
nand U10602 (N_10602,N_10409,N_10551);
or U10603 (N_10603,N_10559,N_10453);
nor U10604 (N_10604,N_10461,N_10490);
nand U10605 (N_10605,N_10468,N_10526);
or U10606 (N_10606,N_10483,N_10538);
and U10607 (N_10607,N_10549,N_10558);
nor U10608 (N_10608,N_10415,N_10475);
or U10609 (N_10609,N_10462,N_10410);
and U10610 (N_10610,N_10432,N_10491);
nand U10611 (N_10611,N_10474,N_10524);
or U10612 (N_10612,N_10427,N_10411);
nor U10613 (N_10613,N_10481,N_10452);
nand U10614 (N_10614,N_10548,N_10430);
xnor U10615 (N_10615,N_10507,N_10543);
nand U10616 (N_10616,N_10460,N_10555);
xor U10617 (N_10617,N_10428,N_10420);
or U10618 (N_10618,N_10465,N_10458);
and U10619 (N_10619,N_10476,N_10466);
nand U10620 (N_10620,N_10451,N_10448);
nand U10621 (N_10621,N_10513,N_10517);
nor U10622 (N_10622,N_10422,N_10431);
or U10623 (N_10623,N_10511,N_10504);
or U10624 (N_10624,N_10541,N_10469);
and U10625 (N_10625,N_10480,N_10438);
xnor U10626 (N_10626,N_10429,N_10501);
and U10627 (N_10627,N_10477,N_10443);
nor U10628 (N_10628,N_10423,N_10407);
and U10629 (N_10629,N_10457,N_10417);
or U10630 (N_10630,N_10557,N_10498);
or U10631 (N_10631,N_10447,N_10494);
nand U10632 (N_10632,N_10444,N_10527);
nand U10633 (N_10633,N_10434,N_10492);
or U10634 (N_10634,N_10408,N_10484);
nand U10635 (N_10635,N_10544,N_10437);
nor U10636 (N_10636,N_10439,N_10516);
xnor U10637 (N_10637,N_10537,N_10425);
xnor U10638 (N_10638,N_10401,N_10400);
nor U10639 (N_10639,N_10414,N_10509);
and U10640 (N_10640,N_10416,N_10533);
and U10641 (N_10641,N_10440,N_10520);
and U10642 (N_10642,N_10428,N_10439);
nor U10643 (N_10643,N_10527,N_10520);
and U10644 (N_10644,N_10408,N_10433);
nor U10645 (N_10645,N_10491,N_10512);
or U10646 (N_10646,N_10406,N_10543);
xor U10647 (N_10647,N_10532,N_10534);
xnor U10648 (N_10648,N_10456,N_10553);
nand U10649 (N_10649,N_10417,N_10474);
nor U10650 (N_10650,N_10445,N_10430);
nor U10651 (N_10651,N_10423,N_10430);
or U10652 (N_10652,N_10485,N_10488);
nor U10653 (N_10653,N_10401,N_10520);
nor U10654 (N_10654,N_10524,N_10547);
nor U10655 (N_10655,N_10420,N_10429);
xnor U10656 (N_10656,N_10527,N_10552);
or U10657 (N_10657,N_10473,N_10549);
xnor U10658 (N_10658,N_10411,N_10546);
xor U10659 (N_10659,N_10541,N_10457);
and U10660 (N_10660,N_10453,N_10526);
xnor U10661 (N_10661,N_10522,N_10444);
xnor U10662 (N_10662,N_10541,N_10440);
nand U10663 (N_10663,N_10534,N_10424);
xnor U10664 (N_10664,N_10554,N_10559);
nand U10665 (N_10665,N_10534,N_10559);
nand U10666 (N_10666,N_10421,N_10475);
nand U10667 (N_10667,N_10422,N_10496);
nand U10668 (N_10668,N_10417,N_10480);
xor U10669 (N_10669,N_10522,N_10488);
or U10670 (N_10670,N_10453,N_10443);
xnor U10671 (N_10671,N_10442,N_10437);
nand U10672 (N_10672,N_10479,N_10435);
nor U10673 (N_10673,N_10501,N_10505);
or U10674 (N_10674,N_10459,N_10433);
and U10675 (N_10675,N_10555,N_10501);
nand U10676 (N_10676,N_10465,N_10482);
xnor U10677 (N_10677,N_10420,N_10457);
nand U10678 (N_10678,N_10413,N_10534);
nand U10679 (N_10679,N_10427,N_10533);
nand U10680 (N_10680,N_10425,N_10475);
xor U10681 (N_10681,N_10472,N_10490);
and U10682 (N_10682,N_10555,N_10458);
or U10683 (N_10683,N_10536,N_10538);
nand U10684 (N_10684,N_10423,N_10479);
and U10685 (N_10685,N_10477,N_10544);
nand U10686 (N_10686,N_10400,N_10424);
nand U10687 (N_10687,N_10547,N_10533);
and U10688 (N_10688,N_10504,N_10412);
and U10689 (N_10689,N_10528,N_10426);
xor U10690 (N_10690,N_10509,N_10491);
or U10691 (N_10691,N_10444,N_10537);
and U10692 (N_10692,N_10403,N_10486);
nor U10693 (N_10693,N_10422,N_10462);
and U10694 (N_10694,N_10448,N_10547);
xnor U10695 (N_10695,N_10511,N_10491);
xnor U10696 (N_10696,N_10450,N_10444);
nor U10697 (N_10697,N_10448,N_10407);
or U10698 (N_10698,N_10490,N_10475);
nand U10699 (N_10699,N_10495,N_10420);
xnor U10700 (N_10700,N_10446,N_10491);
and U10701 (N_10701,N_10492,N_10471);
nand U10702 (N_10702,N_10553,N_10558);
xor U10703 (N_10703,N_10473,N_10537);
nand U10704 (N_10704,N_10449,N_10533);
nor U10705 (N_10705,N_10550,N_10433);
xor U10706 (N_10706,N_10422,N_10513);
nand U10707 (N_10707,N_10420,N_10492);
nand U10708 (N_10708,N_10409,N_10536);
nand U10709 (N_10709,N_10498,N_10469);
xor U10710 (N_10710,N_10482,N_10544);
and U10711 (N_10711,N_10537,N_10426);
nand U10712 (N_10712,N_10431,N_10545);
nor U10713 (N_10713,N_10542,N_10412);
and U10714 (N_10714,N_10495,N_10435);
nand U10715 (N_10715,N_10412,N_10401);
xor U10716 (N_10716,N_10548,N_10407);
or U10717 (N_10717,N_10468,N_10407);
and U10718 (N_10718,N_10453,N_10462);
nor U10719 (N_10719,N_10418,N_10509);
nand U10720 (N_10720,N_10625,N_10644);
nand U10721 (N_10721,N_10626,N_10699);
xnor U10722 (N_10722,N_10616,N_10700);
and U10723 (N_10723,N_10610,N_10632);
xnor U10724 (N_10724,N_10595,N_10584);
xor U10725 (N_10725,N_10707,N_10660);
nand U10726 (N_10726,N_10648,N_10578);
and U10727 (N_10727,N_10577,N_10679);
nor U10728 (N_10728,N_10667,N_10689);
nand U10729 (N_10729,N_10654,N_10688);
nor U10730 (N_10730,N_10593,N_10596);
xor U10731 (N_10731,N_10709,N_10647);
or U10732 (N_10732,N_10718,N_10617);
xnor U10733 (N_10733,N_10708,N_10560);
xor U10734 (N_10734,N_10716,N_10687);
nand U10735 (N_10735,N_10640,N_10587);
and U10736 (N_10736,N_10698,N_10591);
and U10737 (N_10737,N_10603,N_10572);
or U10738 (N_10738,N_10583,N_10562);
nand U10739 (N_10739,N_10636,N_10717);
and U10740 (N_10740,N_10592,N_10713);
nor U10741 (N_10741,N_10702,N_10658);
nor U10742 (N_10742,N_10678,N_10590);
nor U10743 (N_10743,N_10613,N_10705);
or U10744 (N_10744,N_10564,N_10696);
nand U10745 (N_10745,N_10670,N_10657);
nand U10746 (N_10746,N_10711,N_10597);
and U10747 (N_10747,N_10686,N_10609);
or U10748 (N_10748,N_10715,N_10682);
xor U10749 (N_10749,N_10568,N_10674);
xnor U10750 (N_10750,N_10575,N_10661);
nor U10751 (N_10751,N_10604,N_10579);
xor U10752 (N_10752,N_10651,N_10684);
nand U10753 (N_10753,N_10628,N_10642);
xor U10754 (N_10754,N_10668,N_10599);
nand U10755 (N_10755,N_10662,N_10574);
nor U10756 (N_10756,N_10618,N_10563);
and U10757 (N_10757,N_10681,N_10677);
xor U10758 (N_10758,N_10680,N_10652);
nor U10759 (N_10759,N_10580,N_10582);
and U10760 (N_10760,N_10685,N_10573);
and U10761 (N_10761,N_10676,N_10581);
or U10762 (N_10762,N_10695,N_10589);
nor U10763 (N_10763,N_10630,N_10602);
and U10764 (N_10764,N_10719,N_10619);
nand U10765 (N_10765,N_10653,N_10561);
or U10766 (N_10766,N_10671,N_10566);
nand U10767 (N_10767,N_10620,N_10569);
xnor U10768 (N_10768,N_10665,N_10675);
xnor U10769 (N_10769,N_10594,N_10643);
and U10770 (N_10770,N_10627,N_10570);
nor U10771 (N_10771,N_10614,N_10683);
nand U10772 (N_10772,N_10611,N_10649);
xnor U10773 (N_10773,N_10714,N_10664);
xnor U10774 (N_10774,N_10704,N_10706);
nand U10775 (N_10775,N_10598,N_10633);
or U10776 (N_10776,N_10607,N_10703);
nand U10777 (N_10777,N_10585,N_10701);
xor U10778 (N_10778,N_10588,N_10571);
and U10779 (N_10779,N_10576,N_10622);
or U10780 (N_10780,N_10565,N_10656);
or U10781 (N_10781,N_10623,N_10669);
or U10782 (N_10782,N_10673,N_10672);
and U10783 (N_10783,N_10637,N_10600);
xnor U10784 (N_10784,N_10641,N_10567);
nor U10785 (N_10785,N_10586,N_10693);
xor U10786 (N_10786,N_10615,N_10601);
nor U10787 (N_10787,N_10631,N_10697);
or U10788 (N_10788,N_10650,N_10638);
xnor U10789 (N_10789,N_10666,N_10634);
or U10790 (N_10790,N_10606,N_10639);
nand U10791 (N_10791,N_10629,N_10691);
xnor U10792 (N_10792,N_10605,N_10694);
xor U10793 (N_10793,N_10612,N_10635);
nor U10794 (N_10794,N_10659,N_10621);
nor U10795 (N_10795,N_10608,N_10663);
xor U10796 (N_10796,N_10690,N_10645);
and U10797 (N_10797,N_10692,N_10624);
nand U10798 (N_10798,N_10712,N_10710);
nor U10799 (N_10799,N_10646,N_10655);
or U10800 (N_10800,N_10651,N_10603);
nor U10801 (N_10801,N_10574,N_10616);
xor U10802 (N_10802,N_10704,N_10711);
nand U10803 (N_10803,N_10570,N_10644);
xor U10804 (N_10804,N_10659,N_10670);
nand U10805 (N_10805,N_10710,N_10602);
xnor U10806 (N_10806,N_10659,N_10564);
nor U10807 (N_10807,N_10562,N_10623);
or U10808 (N_10808,N_10697,N_10699);
and U10809 (N_10809,N_10587,N_10637);
and U10810 (N_10810,N_10572,N_10644);
nor U10811 (N_10811,N_10627,N_10613);
nand U10812 (N_10812,N_10573,N_10643);
xor U10813 (N_10813,N_10672,N_10616);
nand U10814 (N_10814,N_10571,N_10657);
xnor U10815 (N_10815,N_10598,N_10663);
nor U10816 (N_10816,N_10678,N_10589);
xnor U10817 (N_10817,N_10572,N_10589);
nand U10818 (N_10818,N_10561,N_10641);
and U10819 (N_10819,N_10601,N_10666);
xor U10820 (N_10820,N_10693,N_10648);
nand U10821 (N_10821,N_10602,N_10681);
and U10822 (N_10822,N_10641,N_10638);
and U10823 (N_10823,N_10648,N_10602);
or U10824 (N_10824,N_10629,N_10708);
nand U10825 (N_10825,N_10681,N_10578);
nand U10826 (N_10826,N_10626,N_10714);
nand U10827 (N_10827,N_10674,N_10623);
nor U10828 (N_10828,N_10675,N_10572);
nor U10829 (N_10829,N_10716,N_10711);
xnor U10830 (N_10830,N_10694,N_10703);
and U10831 (N_10831,N_10628,N_10657);
nor U10832 (N_10832,N_10635,N_10631);
and U10833 (N_10833,N_10564,N_10604);
nor U10834 (N_10834,N_10579,N_10634);
nand U10835 (N_10835,N_10709,N_10652);
nor U10836 (N_10836,N_10560,N_10685);
nand U10837 (N_10837,N_10648,N_10601);
and U10838 (N_10838,N_10653,N_10654);
nand U10839 (N_10839,N_10568,N_10663);
and U10840 (N_10840,N_10678,N_10571);
or U10841 (N_10841,N_10638,N_10665);
or U10842 (N_10842,N_10619,N_10663);
or U10843 (N_10843,N_10707,N_10615);
nand U10844 (N_10844,N_10598,N_10688);
nor U10845 (N_10845,N_10710,N_10653);
and U10846 (N_10846,N_10696,N_10598);
nor U10847 (N_10847,N_10583,N_10675);
nand U10848 (N_10848,N_10665,N_10693);
xor U10849 (N_10849,N_10632,N_10624);
or U10850 (N_10850,N_10649,N_10640);
nor U10851 (N_10851,N_10641,N_10564);
xor U10852 (N_10852,N_10718,N_10639);
nor U10853 (N_10853,N_10658,N_10587);
xnor U10854 (N_10854,N_10642,N_10586);
nor U10855 (N_10855,N_10619,N_10639);
and U10856 (N_10856,N_10665,N_10581);
nor U10857 (N_10857,N_10706,N_10703);
nor U10858 (N_10858,N_10632,N_10666);
xor U10859 (N_10859,N_10666,N_10647);
nand U10860 (N_10860,N_10648,N_10675);
or U10861 (N_10861,N_10662,N_10584);
or U10862 (N_10862,N_10664,N_10599);
and U10863 (N_10863,N_10713,N_10655);
and U10864 (N_10864,N_10641,N_10706);
nor U10865 (N_10865,N_10705,N_10666);
xnor U10866 (N_10866,N_10588,N_10662);
and U10867 (N_10867,N_10718,N_10641);
or U10868 (N_10868,N_10626,N_10614);
nand U10869 (N_10869,N_10696,N_10560);
and U10870 (N_10870,N_10575,N_10643);
and U10871 (N_10871,N_10707,N_10620);
and U10872 (N_10872,N_10693,N_10603);
nand U10873 (N_10873,N_10581,N_10620);
and U10874 (N_10874,N_10706,N_10694);
and U10875 (N_10875,N_10655,N_10630);
and U10876 (N_10876,N_10707,N_10648);
xnor U10877 (N_10877,N_10639,N_10644);
xnor U10878 (N_10878,N_10682,N_10708);
nand U10879 (N_10879,N_10634,N_10643);
or U10880 (N_10880,N_10753,N_10866);
nand U10881 (N_10881,N_10790,N_10774);
or U10882 (N_10882,N_10860,N_10841);
or U10883 (N_10883,N_10822,N_10721);
or U10884 (N_10884,N_10874,N_10806);
nand U10885 (N_10885,N_10749,N_10724);
nand U10886 (N_10886,N_10793,N_10761);
or U10887 (N_10887,N_10819,N_10772);
nand U10888 (N_10888,N_10789,N_10856);
nand U10889 (N_10889,N_10843,N_10823);
nor U10890 (N_10890,N_10754,N_10800);
or U10891 (N_10891,N_10760,N_10871);
and U10892 (N_10892,N_10723,N_10763);
nand U10893 (N_10893,N_10861,N_10862);
nand U10894 (N_10894,N_10788,N_10814);
xnor U10895 (N_10895,N_10835,N_10870);
nor U10896 (N_10896,N_10836,N_10734);
nand U10897 (N_10897,N_10869,N_10816);
or U10898 (N_10898,N_10801,N_10787);
xor U10899 (N_10899,N_10757,N_10762);
xor U10900 (N_10900,N_10837,N_10865);
nor U10901 (N_10901,N_10833,N_10778);
nand U10902 (N_10902,N_10838,N_10737);
or U10903 (N_10903,N_10847,N_10868);
nand U10904 (N_10904,N_10776,N_10805);
or U10905 (N_10905,N_10840,N_10767);
nand U10906 (N_10906,N_10794,N_10829);
nand U10907 (N_10907,N_10875,N_10784);
or U10908 (N_10908,N_10852,N_10810);
or U10909 (N_10909,N_10849,N_10797);
and U10910 (N_10910,N_10732,N_10850);
xor U10911 (N_10911,N_10781,N_10831);
nor U10912 (N_10912,N_10786,N_10742);
and U10913 (N_10913,N_10809,N_10820);
nor U10914 (N_10914,N_10857,N_10878);
nor U10915 (N_10915,N_10755,N_10791);
and U10916 (N_10916,N_10792,N_10879);
xnor U10917 (N_10917,N_10745,N_10783);
nor U10918 (N_10918,N_10825,N_10863);
or U10919 (N_10919,N_10785,N_10813);
and U10920 (N_10920,N_10733,N_10779);
or U10921 (N_10921,N_10811,N_10771);
or U10922 (N_10922,N_10777,N_10746);
nand U10923 (N_10923,N_10769,N_10817);
xnor U10924 (N_10924,N_10802,N_10750);
nand U10925 (N_10925,N_10877,N_10738);
and U10926 (N_10926,N_10828,N_10842);
nor U10927 (N_10927,N_10747,N_10764);
nor U10928 (N_10928,N_10832,N_10848);
xnor U10929 (N_10929,N_10798,N_10720);
nand U10930 (N_10930,N_10859,N_10864);
xnor U10931 (N_10931,N_10751,N_10766);
xnor U10932 (N_10932,N_10728,N_10815);
or U10933 (N_10933,N_10872,N_10743);
and U10934 (N_10934,N_10729,N_10854);
xor U10935 (N_10935,N_10808,N_10827);
xor U10936 (N_10936,N_10727,N_10844);
xor U10937 (N_10937,N_10873,N_10758);
xnor U10938 (N_10938,N_10830,N_10834);
nor U10939 (N_10939,N_10818,N_10765);
nor U10940 (N_10940,N_10735,N_10775);
nand U10941 (N_10941,N_10744,N_10722);
or U10942 (N_10942,N_10799,N_10812);
xnor U10943 (N_10943,N_10851,N_10773);
xnor U10944 (N_10944,N_10845,N_10853);
xor U10945 (N_10945,N_10770,N_10780);
or U10946 (N_10946,N_10795,N_10756);
or U10947 (N_10947,N_10807,N_10736);
nand U10948 (N_10948,N_10748,N_10826);
nor U10949 (N_10949,N_10730,N_10739);
xnor U10950 (N_10950,N_10846,N_10867);
or U10951 (N_10951,N_10803,N_10725);
or U10952 (N_10952,N_10824,N_10821);
nand U10953 (N_10953,N_10876,N_10782);
or U10954 (N_10954,N_10804,N_10752);
nor U10955 (N_10955,N_10796,N_10741);
xor U10956 (N_10956,N_10858,N_10768);
and U10957 (N_10957,N_10731,N_10855);
nand U10958 (N_10958,N_10726,N_10839);
xnor U10959 (N_10959,N_10740,N_10759);
or U10960 (N_10960,N_10864,N_10764);
or U10961 (N_10961,N_10751,N_10840);
or U10962 (N_10962,N_10769,N_10863);
and U10963 (N_10963,N_10742,N_10782);
and U10964 (N_10964,N_10774,N_10848);
nor U10965 (N_10965,N_10813,N_10864);
or U10966 (N_10966,N_10807,N_10869);
nor U10967 (N_10967,N_10816,N_10862);
xor U10968 (N_10968,N_10788,N_10819);
xnor U10969 (N_10969,N_10738,N_10759);
nor U10970 (N_10970,N_10853,N_10765);
nor U10971 (N_10971,N_10833,N_10775);
or U10972 (N_10972,N_10802,N_10741);
nand U10973 (N_10973,N_10737,N_10795);
xor U10974 (N_10974,N_10729,N_10802);
or U10975 (N_10975,N_10786,N_10723);
nand U10976 (N_10976,N_10815,N_10758);
or U10977 (N_10977,N_10829,N_10772);
xor U10978 (N_10978,N_10819,N_10802);
or U10979 (N_10979,N_10865,N_10738);
nor U10980 (N_10980,N_10772,N_10799);
xnor U10981 (N_10981,N_10732,N_10781);
or U10982 (N_10982,N_10846,N_10829);
or U10983 (N_10983,N_10815,N_10801);
xor U10984 (N_10984,N_10866,N_10876);
and U10985 (N_10985,N_10721,N_10829);
nor U10986 (N_10986,N_10733,N_10720);
nand U10987 (N_10987,N_10747,N_10756);
nand U10988 (N_10988,N_10776,N_10819);
nor U10989 (N_10989,N_10854,N_10769);
xor U10990 (N_10990,N_10878,N_10839);
nor U10991 (N_10991,N_10725,N_10833);
xnor U10992 (N_10992,N_10726,N_10815);
nand U10993 (N_10993,N_10843,N_10820);
and U10994 (N_10994,N_10752,N_10748);
and U10995 (N_10995,N_10866,N_10747);
and U10996 (N_10996,N_10820,N_10754);
nor U10997 (N_10997,N_10876,N_10721);
and U10998 (N_10998,N_10781,N_10761);
xor U10999 (N_10999,N_10727,N_10734);
nor U11000 (N_11000,N_10817,N_10836);
nor U11001 (N_11001,N_10817,N_10767);
nand U11002 (N_11002,N_10771,N_10785);
nor U11003 (N_11003,N_10770,N_10831);
nand U11004 (N_11004,N_10821,N_10733);
and U11005 (N_11005,N_10806,N_10840);
nand U11006 (N_11006,N_10769,N_10841);
nand U11007 (N_11007,N_10797,N_10726);
xor U11008 (N_11008,N_10767,N_10850);
and U11009 (N_11009,N_10772,N_10861);
nand U11010 (N_11010,N_10766,N_10786);
nor U11011 (N_11011,N_10766,N_10875);
or U11012 (N_11012,N_10775,N_10802);
nand U11013 (N_11013,N_10767,N_10819);
and U11014 (N_11014,N_10802,N_10724);
and U11015 (N_11015,N_10746,N_10876);
nand U11016 (N_11016,N_10756,N_10772);
nor U11017 (N_11017,N_10753,N_10855);
nand U11018 (N_11018,N_10870,N_10731);
xor U11019 (N_11019,N_10813,N_10814);
nand U11020 (N_11020,N_10729,N_10750);
or U11021 (N_11021,N_10878,N_10773);
and U11022 (N_11022,N_10754,N_10848);
nor U11023 (N_11023,N_10760,N_10774);
xnor U11024 (N_11024,N_10725,N_10850);
nor U11025 (N_11025,N_10772,N_10846);
nand U11026 (N_11026,N_10768,N_10722);
xor U11027 (N_11027,N_10830,N_10791);
or U11028 (N_11028,N_10840,N_10720);
nor U11029 (N_11029,N_10834,N_10859);
or U11030 (N_11030,N_10807,N_10835);
xor U11031 (N_11031,N_10739,N_10835);
or U11032 (N_11032,N_10857,N_10753);
and U11033 (N_11033,N_10810,N_10809);
and U11034 (N_11034,N_10850,N_10722);
and U11035 (N_11035,N_10870,N_10792);
nor U11036 (N_11036,N_10729,N_10773);
and U11037 (N_11037,N_10872,N_10788);
and U11038 (N_11038,N_10722,N_10811);
nor U11039 (N_11039,N_10878,N_10796);
or U11040 (N_11040,N_10941,N_10886);
xor U11041 (N_11041,N_10921,N_11035);
nor U11042 (N_11042,N_10949,N_10978);
and U11043 (N_11043,N_10983,N_10982);
xnor U11044 (N_11044,N_10912,N_10891);
xnor U11045 (N_11045,N_11000,N_10996);
xnor U11046 (N_11046,N_10954,N_11029);
nand U11047 (N_11047,N_10992,N_10976);
xnor U11048 (N_11048,N_10936,N_10993);
nor U11049 (N_11049,N_11023,N_11024);
and U11050 (N_11050,N_10947,N_10920);
or U11051 (N_11051,N_11003,N_10986);
xnor U11052 (N_11052,N_10940,N_10990);
nand U11053 (N_11053,N_10881,N_10950);
nor U11054 (N_11054,N_11014,N_10952);
xnor U11055 (N_11055,N_10926,N_10893);
or U11056 (N_11056,N_10977,N_10973);
xnor U11057 (N_11057,N_10960,N_10905);
nor U11058 (N_11058,N_10894,N_10904);
xnor U11059 (N_11059,N_11012,N_10907);
and U11060 (N_11060,N_10919,N_11020);
xnor U11061 (N_11061,N_11028,N_10901);
nor U11062 (N_11062,N_11039,N_10974);
nand U11063 (N_11063,N_11038,N_11002);
nand U11064 (N_11064,N_10968,N_10911);
and U11065 (N_11065,N_10975,N_10943);
xnor U11066 (N_11066,N_10909,N_11027);
xnor U11067 (N_11067,N_11011,N_10998);
nor U11068 (N_11068,N_10979,N_10938);
xor U11069 (N_11069,N_10903,N_10981);
nand U11070 (N_11070,N_10970,N_11026);
nor U11071 (N_11071,N_10971,N_10924);
and U11072 (N_11072,N_11034,N_10980);
xor U11073 (N_11073,N_11030,N_10929);
xnor U11074 (N_11074,N_10908,N_11009);
nand U11075 (N_11075,N_10999,N_10984);
xnor U11076 (N_11076,N_10895,N_11005);
nor U11077 (N_11077,N_11031,N_10923);
nand U11078 (N_11078,N_10932,N_10964);
xnor U11079 (N_11079,N_10946,N_10906);
xnor U11080 (N_11080,N_10898,N_10933);
or U11081 (N_11081,N_10955,N_11018);
xnor U11082 (N_11082,N_11008,N_10945);
or U11083 (N_11083,N_10918,N_10953);
or U11084 (N_11084,N_10888,N_10887);
or U11085 (N_11085,N_10997,N_10957);
xnor U11086 (N_11086,N_10958,N_11010);
xor U11087 (N_11087,N_10956,N_11036);
xnor U11088 (N_11088,N_10899,N_10935);
nor U11089 (N_11089,N_11016,N_10966);
or U11090 (N_11090,N_10927,N_10934);
and U11091 (N_11091,N_11004,N_10959);
or U11092 (N_11092,N_10922,N_10914);
or U11093 (N_11093,N_10944,N_11019);
nor U11094 (N_11094,N_10967,N_10937);
xor U11095 (N_11095,N_10913,N_10931);
or U11096 (N_11096,N_10987,N_11006);
nand U11097 (N_11097,N_11021,N_10961);
and U11098 (N_11098,N_11037,N_11032);
and U11099 (N_11099,N_10902,N_10951);
or U11100 (N_11100,N_10916,N_10889);
nand U11101 (N_11101,N_10884,N_11017);
nor U11102 (N_11102,N_10942,N_10896);
nor U11103 (N_11103,N_11007,N_10885);
nand U11104 (N_11104,N_11025,N_10910);
or U11105 (N_11105,N_10962,N_10948);
and U11106 (N_11106,N_11013,N_10989);
or U11107 (N_11107,N_10880,N_10882);
nand U11108 (N_11108,N_11033,N_10883);
and U11109 (N_11109,N_10988,N_11022);
or U11110 (N_11110,N_10965,N_10928);
or U11111 (N_11111,N_10925,N_11001);
nor U11112 (N_11112,N_10963,N_10994);
nor U11113 (N_11113,N_10939,N_10985);
and U11114 (N_11114,N_10995,N_10890);
xnor U11115 (N_11115,N_10917,N_10915);
xor U11116 (N_11116,N_10892,N_10900);
and U11117 (N_11117,N_11015,N_10897);
and U11118 (N_11118,N_10972,N_10969);
nor U11119 (N_11119,N_10930,N_10991);
nor U11120 (N_11120,N_10926,N_10979);
and U11121 (N_11121,N_10904,N_10999);
or U11122 (N_11122,N_11027,N_10934);
xnor U11123 (N_11123,N_11036,N_10931);
xnor U11124 (N_11124,N_10925,N_10970);
nand U11125 (N_11125,N_10940,N_10978);
xnor U11126 (N_11126,N_10984,N_10966);
nand U11127 (N_11127,N_10978,N_10882);
nor U11128 (N_11128,N_10918,N_10982);
or U11129 (N_11129,N_10908,N_10920);
nor U11130 (N_11130,N_10944,N_10893);
or U11131 (N_11131,N_11003,N_10988);
or U11132 (N_11132,N_10915,N_10921);
or U11133 (N_11133,N_10992,N_10986);
nand U11134 (N_11134,N_10909,N_10992);
or U11135 (N_11135,N_10937,N_10964);
xnor U11136 (N_11136,N_10957,N_10906);
and U11137 (N_11137,N_10971,N_10983);
nand U11138 (N_11138,N_10990,N_10982);
and U11139 (N_11139,N_10906,N_11012);
nand U11140 (N_11140,N_11016,N_11032);
nor U11141 (N_11141,N_11015,N_10971);
nor U11142 (N_11142,N_10972,N_11027);
and U11143 (N_11143,N_10978,N_10963);
and U11144 (N_11144,N_10984,N_10949);
xor U11145 (N_11145,N_10884,N_10993);
nor U11146 (N_11146,N_11007,N_10923);
or U11147 (N_11147,N_10897,N_10987);
and U11148 (N_11148,N_11000,N_10938);
nand U11149 (N_11149,N_10961,N_11011);
nor U11150 (N_11150,N_10979,N_10959);
and U11151 (N_11151,N_10923,N_10883);
xor U11152 (N_11152,N_11016,N_10911);
and U11153 (N_11153,N_10979,N_10963);
nor U11154 (N_11154,N_10997,N_10929);
or U11155 (N_11155,N_11001,N_10904);
nor U11156 (N_11156,N_10956,N_10992);
xor U11157 (N_11157,N_11033,N_10990);
nand U11158 (N_11158,N_10931,N_10996);
nor U11159 (N_11159,N_10925,N_11030);
or U11160 (N_11160,N_10995,N_10952);
xnor U11161 (N_11161,N_10963,N_11039);
xnor U11162 (N_11162,N_10935,N_10965);
nor U11163 (N_11163,N_10950,N_11003);
or U11164 (N_11164,N_10992,N_11036);
and U11165 (N_11165,N_11032,N_10947);
and U11166 (N_11166,N_10918,N_10955);
or U11167 (N_11167,N_10971,N_10968);
or U11168 (N_11168,N_10931,N_10950);
nor U11169 (N_11169,N_10922,N_10885);
xnor U11170 (N_11170,N_10975,N_10917);
nand U11171 (N_11171,N_10895,N_10948);
and U11172 (N_11172,N_10967,N_11023);
and U11173 (N_11173,N_10970,N_10914);
nor U11174 (N_11174,N_10902,N_10979);
and U11175 (N_11175,N_11009,N_11005);
and U11176 (N_11176,N_10998,N_11000);
or U11177 (N_11177,N_10921,N_10975);
xnor U11178 (N_11178,N_10979,N_11039);
xnor U11179 (N_11179,N_10994,N_10945);
or U11180 (N_11180,N_10968,N_10983);
nand U11181 (N_11181,N_10912,N_10959);
and U11182 (N_11182,N_10954,N_11007);
nand U11183 (N_11183,N_11003,N_10897);
xnor U11184 (N_11184,N_10925,N_10894);
nand U11185 (N_11185,N_10949,N_10891);
nor U11186 (N_11186,N_10976,N_10926);
nor U11187 (N_11187,N_10931,N_11011);
or U11188 (N_11188,N_10911,N_10919);
nand U11189 (N_11189,N_10988,N_11034);
xor U11190 (N_11190,N_10887,N_11031);
nand U11191 (N_11191,N_10908,N_11035);
and U11192 (N_11192,N_11026,N_10932);
nand U11193 (N_11193,N_10927,N_10890);
nand U11194 (N_11194,N_11015,N_10894);
xnor U11195 (N_11195,N_10896,N_10919);
or U11196 (N_11196,N_11006,N_11020);
nor U11197 (N_11197,N_10892,N_10996);
nand U11198 (N_11198,N_11036,N_10918);
and U11199 (N_11199,N_10957,N_10890);
xnor U11200 (N_11200,N_11115,N_11117);
or U11201 (N_11201,N_11064,N_11065);
xor U11202 (N_11202,N_11073,N_11173);
or U11203 (N_11203,N_11103,N_11070);
xnor U11204 (N_11204,N_11194,N_11084);
nor U11205 (N_11205,N_11056,N_11133);
xnor U11206 (N_11206,N_11152,N_11192);
xnor U11207 (N_11207,N_11150,N_11040);
nor U11208 (N_11208,N_11042,N_11162);
nand U11209 (N_11209,N_11161,N_11090);
and U11210 (N_11210,N_11100,N_11049);
nor U11211 (N_11211,N_11186,N_11195);
or U11212 (N_11212,N_11104,N_11156);
or U11213 (N_11213,N_11149,N_11093);
nor U11214 (N_11214,N_11168,N_11105);
xor U11215 (N_11215,N_11191,N_11153);
or U11216 (N_11216,N_11116,N_11190);
nand U11217 (N_11217,N_11126,N_11158);
xor U11218 (N_11218,N_11148,N_11199);
nor U11219 (N_11219,N_11159,N_11166);
or U11220 (N_11220,N_11139,N_11167);
nor U11221 (N_11221,N_11055,N_11170);
and U11222 (N_11222,N_11118,N_11050);
nor U11223 (N_11223,N_11079,N_11089);
nor U11224 (N_11224,N_11151,N_11130);
xor U11225 (N_11225,N_11075,N_11163);
or U11226 (N_11226,N_11086,N_11185);
xnor U11227 (N_11227,N_11140,N_11196);
nor U11228 (N_11228,N_11189,N_11077);
xor U11229 (N_11229,N_11107,N_11085);
xnor U11230 (N_11230,N_11069,N_11178);
nor U11231 (N_11231,N_11063,N_11045);
and U11232 (N_11232,N_11059,N_11113);
nor U11233 (N_11233,N_11138,N_11147);
nor U11234 (N_11234,N_11124,N_11154);
nand U11235 (N_11235,N_11076,N_11082);
nand U11236 (N_11236,N_11088,N_11143);
nand U11237 (N_11237,N_11125,N_11068);
nor U11238 (N_11238,N_11146,N_11127);
nand U11239 (N_11239,N_11081,N_11180);
nand U11240 (N_11240,N_11046,N_11112);
nor U11241 (N_11241,N_11181,N_11187);
nand U11242 (N_11242,N_11054,N_11182);
xor U11243 (N_11243,N_11141,N_11179);
nor U11244 (N_11244,N_11135,N_11109);
nand U11245 (N_11245,N_11155,N_11106);
nand U11246 (N_11246,N_11131,N_11053);
nor U11247 (N_11247,N_11080,N_11071);
nor U11248 (N_11248,N_11043,N_11165);
or U11249 (N_11249,N_11169,N_11094);
or U11250 (N_11250,N_11122,N_11099);
nand U11251 (N_11251,N_11066,N_11092);
or U11252 (N_11252,N_11123,N_11128);
and U11253 (N_11253,N_11176,N_11078);
and U11254 (N_11254,N_11072,N_11041);
or U11255 (N_11255,N_11157,N_11160);
or U11256 (N_11256,N_11096,N_11102);
nor U11257 (N_11257,N_11174,N_11175);
xor U11258 (N_11258,N_11184,N_11058);
and U11259 (N_11259,N_11047,N_11120);
and U11260 (N_11260,N_11091,N_11101);
nand U11261 (N_11261,N_11132,N_11098);
and U11262 (N_11262,N_11145,N_11121);
nor U11263 (N_11263,N_11044,N_11060);
xnor U11264 (N_11264,N_11083,N_11188);
nor U11265 (N_11265,N_11142,N_11134);
or U11266 (N_11266,N_11061,N_11111);
nor U11267 (N_11267,N_11108,N_11137);
xnor U11268 (N_11268,N_11129,N_11057);
nand U11269 (N_11269,N_11067,N_11087);
or U11270 (N_11270,N_11097,N_11177);
xor U11271 (N_11271,N_11183,N_11052);
or U11272 (N_11272,N_11198,N_11119);
xor U11273 (N_11273,N_11062,N_11144);
nor U11274 (N_11274,N_11095,N_11074);
and U11275 (N_11275,N_11114,N_11136);
nand U11276 (N_11276,N_11051,N_11193);
xor U11277 (N_11277,N_11172,N_11171);
or U11278 (N_11278,N_11197,N_11110);
nand U11279 (N_11279,N_11164,N_11048);
nor U11280 (N_11280,N_11120,N_11055);
xor U11281 (N_11281,N_11114,N_11175);
or U11282 (N_11282,N_11080,N_11163);
xnor U11283 (N_11283,N_11136,N_11066);
and U11284 (N_11284,N_11138,N_11063);
nand U11285 (N_11285,N_11150,N_11095);
nand U11286 (N_11286,N_11102,N_11167);
nand U11287 (N_11287,N_11092,N_11161);
nand U11288 (N_11288,N_11180,N_11083);
or U11289 (N_11289,N_11129,N_11070);
or U11290 (N_11290,N_11139,N_11096);
nand U11291 (N_11291,N_11190,N_11098);
xnor U11292 (N_11292,N_11167,N_11040);
nor U11293 (N_11293,N_11159,N_11164);
and U11294 (N_11294,N_11123,N_11080);
xnor U11295 (N_11295,N_11140,N_11103);
and U11296 (N_11296,N_11148,N_11143);
or U11297 (N_11297,N_11135,N_11149);
and U11298 (N_11298,N_11179,N_11149);
or U11299 (N_11299,N_11079,N_11184);
or U11300 (N_11300,N_11198,N_11155);
xnor U11301 (N_11301,N_11062,N_11041);
or U11302 (N_11302,N_11050,N_11180);
nand U11303 (N_11303,N_11162,N_11180);
nand U11304 (N_11304,N_11195,N_11135);
xor U11305 (N_11305,N_11061,N_11073);
or U11306 (N_11306,N_11170,N_11131);
nor U11307 (N_11307,N_11141,N_11108);
or U11308 (N_11308,N_11069,N_11133);
xor U11309 (N_11309,N_11109,N_11091);
nor U11310 (N_11310,N_11168,N_11093);
or U11311 (N_11311,N_11148,N_11128);
and U11312 (N_11312,N_11124,N_11108);
xor U11313 (N_11313,N_11093,N_11138);
or U11314 (N_11314,N_11048,N_11127);
or U11315 (N_11315,N_11051,N_11123);
or U11316 (N_11316,N_11162,N_11046);
xnor U11317 (N_11317,N_11171,N_11041);
or U11318 (N_11318,N_11055,N_11183);
xnor U11319 (N_11319,N_11055,N_11122);
nand U11320 (N_11320,N_11116,N_11065);
xor U11321 (N_11321,N_11125,N_11194);
nand U11322 (N_11322,N_11054,N_11173);
or U11323 (N_11323,N_11197,N_11103);
xnor U11324 (N_11324,N_11112,N_11145);
xnor U11325 (N_11325,N_11156,N_11132);
or U11326 (N_11326,N_11168,N_11138);
nand U11327 (N_11327,N_11059,N_11086);
nand U11328 (N_11328,N_11096,N_11066);
or U11329 (N_11329,N_11049,N_11144);
nor U11330 (N_11330,N_11189,N_11051);
xnor U11331 (N_11331,N_11086,N_11107);
nand U11332 (N_11332,N_11114,N_11097);
and U11333 (N_11333,N_11159,N_11157);
and U11334 (N_11334,N_11199,N_11081);
nand U11335 (N_11335,N_11177,N_11163);
nand U11336 (N_11336,N_11114,N_11106);
nor U11337 (N_11337,N_11188,N_11194);
nand U11338 (N_11338,N_11163,N_11198);
nand U11339 (N_11339,N_11194,N_11070);
nand U11340 (N_11340,N_11198,N_11189);
nor U11341 (N_11341,N_11042,N_11120);
or U11342 (N_11342,N_11143,N_11195);
xnor U11343 (N_11343,N_11167,N_11180);
xor U11344 (N_11344,N_11162,N_11161);
nand U11345 (N_11345,N_11069,N_11177);
nor U11346 (N_11346,N_11146,N_11089);
xor U11347 (N_11347,N_11061,N_11134);
nor U11348 (N_11348,N_11132,N_11148);
and U11349 (N_11349,N_11068,N_11089);
xnor U11350 (N_11350,N_11132,N_11166);
or U11351 (N_11351,N_11156,N_11099);
and U11352 (N_11352,N_11165,N_11156);
nand U11353 (N_11353,N_11162,N_11072);
or U11354 (N_11354,N_11098,N_11075);
nand U11355 (N_11355,N_11056,N_11186);
xor U11356 (N_11356,N_11055,N_11040);
xnor U11357 (N_11357,N_11186,N_11100);
xnor U11358 (N_11358,N_11120,N_11044);
and U11359 (N_11359,N_11142,N_11157);
or U11360 (N_11360,N_11303,N_11277);
and U11361 (N_11361,N_11245,N_11330);
and U11362 (N_11362,N_11235,N_11205);
nor U11363 (N_11363,N_11229,N_11333);
xnor U11364 (N_11364,N_11358,N_11304);
and U11365 (N_11365,N_11266,N_11272);
nor U11366 (N_11366,N_11265,N_11209);
and U11367 (N_11367,N_11359,N_11356);
nand U11368 (N_11368,N_11280,N_11217);
and U11369 (N_11369,N_11345,N_11253);
xnor U11370 (N_11370,N_11309,N_11326);
nor U11371 (N_11371,N_11224,N_11262);
or U11372 (N_11372,N_11246,N_11307);
nor U11373 (N_11373,N_11222,N_11216);
or U11374 (N_11374,N_11221,N_11301);
nor U11375 (N_11375,N_11236,N_11278);
and U11376 (N_11376,N_11276,N_11249);
nand U11377 (N_11377,N_11287,N_11200);
nand U11378 (N_11378,N_11352,N_11263);
nand U11379 (N_11379,N_11256,N_11315);
or U11380 (N_11380,N_11243,N_11284);
and U11381 (N_11381,N_11259,N_11232);
nor U11382 (N_11382,N_11294,N_11312);
or U11383 (N_11383,N_11241,N_11317);
or U11384 (N_11384,N_11225,N_11231);
and U11385 (N_11385,N_11215,N_11282);
xnor U11386 (N_11386,N_11201,N_11336);
or U11387 (N_11387,N_11291,N_11223);
xor U11388 (N_11388,N_11230,N_11323);
and U11389 (N_11389,N_11227,N_11237);
nor U11390 (N_11390,N_11239,N_11350);
xnor U11391 (N_11391,N_11335,N_11268);
xnor U11392 (N_11392,N_11273,N_11305);
nor U11393 (N_11393,N_11210,N_11327);
nand U11394 (N_11394,N_11238,N_11355);
or U11395 (N_11395,N_11347,N_11218);
xnor U11396 (N_11396,N_11343,N_11319);
nor U11397 (N_11397,N_11339,N_11270);
nand U11398 (N_11398,N_11214,N_11290);
nor U11399 (N_11399,N_11255,N_11334);
and U11400 (N_11400,N_11204,N_11310);
nand U11401 (N_11401,N_11283,N_11340);
xor U11402 (N_11402,N_11267,N_11254);
and U11403 (N_11403,N_11331,N_11341);
and U11404 (N_11404,N_11332,N_11349);
or U11405 (N_11405,N_11322,N_11329);
nor U11406 (N_11406,N_11279,N_11342);
nor U11407 (N_11407,N_11348,N_11328);
and U11408 (N_11408,N_11296,N_11308);
or U11409 (N_11409,N_11306,N_11299);
nor U11410 (N_11410,N_11258,N_11269);
xnor U11411 (N_11411,N_11321,N_11257);
or U11412 (N_11412,N_11320,N_11213);
or U11413 (N_11413,N_11357,N_11233);
xor U11414 (N_11414,N_11260,N_11289);
nand U11415 (N_11415,N_11298,N_11264);
nor U11416 (N_11416,N_11344,N_11300);
nor U11417 (N_11417,N_11261,N_11314);
or U11418 (N_11418,N_11228,N_11297);
xor U11419 (N_11419,N_11313,N_11234);
nand U11420 (N_11420,N_11286,N_11351);
xnor U11421 (N_11421,N_11324,N_11353);
or U11422 (N_11422,N_11202,N_11295);
nand U11423 (N_11423,N_11244,N_11354);
and U11424 (N_11424,N_11281,N_11302);
xor U11425 (N_11425,N_11285,N_11240);
nor U11426 (N_11426,N_11212,N_11219);
nor U11427 (N_11427,N_11207,N_11220);
and U11428 (N_11428,N_11293,N_11203);
or U11429 (N_11429,N_11226,N_11242);
nor U11430 (N_11430,N_11292,N_11252);
nand U11431 (N_11431,N_11250,N_11247);
nand U11432 (N_11432,N_11338,N_11311);
nor U11433 (N_11433,N_11211,N_11325);
and U11434 (N_11434,N_11318,N_11206);
or U11435 (N_11435,N_11271,N_11275);
and U11436 (N_11436,N_11251,N_11316);
xor U11437 (N_11437,N_11337,N_11346);
nand U11438 (N_11438,N_11288,N_11274);
nor U11439 (N_11439,N_11248,N_11208);
nor U11440 (N_11440,N_11240,N_11343);
nand U11441 (N_11441,N_11208,N_11298);
nand U11442 (N_11442,N_11273,N_11324);
nor U11443 (N_11443,N_11307,N_11238);
and U11444 (N_11444,N_11295,N_11229);
xor U11445 (N_11445,N_11232,N_11300);
nor U11446 (N_11446,N_11346,N_11248);
xnor U11447 (N_11447,N_11286,N_11293);
nor U11448 (N_11448,N_11276,N_11232);
nand U11449 (N_11449,N_11304,N_11328);
nand U11450 (N_11450,N_11288,N_11245);
and U11451 (N_11451,N_11207,N_11234);
and U11452 (N_11452,N_11275,N_11200);
xor U11453 (N_11453,N_11233,N_11336);
and U11454 (N_11454,N_11288,N_11265);
or U11455 (N_11455,N_11320,N_11257);
nand U11456 (N_11456,N_11231,N_11222);
nor U11457 (N_11457,N_11323,N_11314);
xor U11458 (N_11458,N_11269,N_11203);
or U11459 (N_11459,N_11237,N_11304);
xnor U11460 (N_11460,N_11310,N_11237);
xor U11461 (N_11461,N_11299,N_11285);
nor U11462 (N_11462,N_11205,N_11229);
nor U11463 (N_11463,N_11240,N_11337);
or U11464 (N_11464,N_11216,N_11308);
nand U11465 (N_11465,N_11295,N_11315);
nor U11466 (N_11466,N_11334,N_11262);
or U11467 (N_11467,N_11315,N_11345);
and U11468 (N_11468,N_11226,N_11246);
xnor U11469 (N_11469,N_11320,N_11300);
and U11470 (N_11470,N_11217,N_11323);
or U11471 (N_11471,N_11342,N_11314);
or U11472 (N_11472,N_11302,N_11209);
or U11473 (N_11473,N_11351,N_11316);
nor U11474 (N_11474,N_11231,N_11212);
nor U11475 (N_11475,N_11319,N_11358);
nor U11476 (N_11476,N_11305,N_11339);
nor U11477 (N_11477,N_11356,N_11276);
or U11478 (N_11478,N_11304,N_11329);
nand U11479 (N_11479,N_11215,N_11343);
nor U11480 (N_11480,N_11313,N_11258);
and U11481 (N_11481,N_11278,N_11300);
nor U11482 (N_11482,N_11335,N_11224);
or U11483 (N_11483,N_11251,N_11268);
or U11484 (N_11484,N_11217,N_11352);
or U11485 (N_11485,N_11344,N_11294);
nand U11486 (N_11486,N_11325,N_11225);
nor U11487 (N_11487,N_11334,N_11329);
nand U11488 (N_11488,N_11245,N_11243);
or U11489 (N_11489,N_11274,N_11310);
nor U11490 (N_11490,N_11332,N_11257);
or U11491 (N_11491,N_11309,N_11214);
nand U11492 (N_11492,N_11249,N_11209);
nand U11493 (N_11493,N_11234,N_11346);
xnor U11494 (N_11494,N_11263,N_11307);
or U11495 (N_11495,N_11264,N_11253);
and U11496 (N_11496,N_11202,N_11205);
xor U11497 (N_11497,N_11216,N_11334);
and U11498 (N_11498,N_11228,N_11282);
or U11499 (N_11499,N_11218,N_11311);
xnor U11500 (N_11500,N_11205,N_11281);
xor U11501 (N_11501,N_11288,N_11306);
and U11502 (N_11502,N_11244,N_11311);
nor U11503 (N_11503,N_11255,N_11288);
nand U11504 (N_11504,N_11314,N_11294);
nor U11505 (N_11505,N_11255,N_11312);
xnor U11506 (N_11506,N_11244,N_11279);
nor U11507 (N_11507,N_11315,N_11348);
or U11508 (N_11508,N_11325,N_11237);
and U11509 (N_11509,N_11271,N_11227);
and U11510 (N_11510,N_11288,N_11309);
xnor U11511 (N_11511,N_11230,N_11310);
nor U11512 (N_11512,N_11221,N_11291);
nor U11513 (N_11513,N_11257,N_11276);
or U11514 (N_11514,N_11250,N_11210);
nand U11515 (N_11515,N_11250,N_11290);
or U11516 (N_11516,N_11281,N_11319);
nor U11517 (N_11517,N_11255,N_11308);
nor U11518 (N_11518,N_11246,N_11244);
xor U11519 (N_11519,N_11275,N_11205);
nor U11520 (N_11520,N_11518,N_11491);
nand U11521 (N_11521,N_11402,N_11427);
nand U11522 (N_11522,N_11511,N_11488);
or U11523 (N_11523,N_11418,N_11423);
or U11524 (N_11524,N_11469,N_11376);
and U11525 (N_11525,N_11366,N_11519);
nand U11526 (N_11526,N_11407,N_11479);
or U11527 (N_11527,N_11365,N_11362);
xnor U11528 (N_11528,N_11450,N_11506);
nor U11529 (N_11529,N_11382,N_11425);
nand U11530 (N_11530,N_11367,N_11493);
or U11531 (N_11531,N_11455,N_11411);
and U11532 (N_11532,N_11426,N_11422);
xor U11533 (N_11533,N_11448,N_11489);
and U11534 (N_11534,N_11442,N_11464);
or U11535 (N_11535,N_11398,N_11463);
and U11536 (N_11536,N_11377,N_11412);
nand U11537 (N_11537,N_11393,N_11458);
nor U11538 (N_11538,N_11410,N_11401);
nor U11539 (N_11539,N_11421,N_11431);
nand U11540 (N_11540,N_11485,N_11372);
nor U11541 (N_11541,N_11378,N_11394);
and U11542 (N_11542,N_11510,N_11496);
xnor U11543 (N_11543,N_11483,N_11409);
nor U11544 (N_11544,N_11446,N_11397);
xor U11545 (N_11545,N_11507,N_11375);
nand U11546 (N_11546,N_11404,N_11486);
nor U11547 (N_11547,N_11403,N_11452);
nor U11548 (N_11548,N_11443,N_11381);
or U11549 (N_11549,N_11392,N_11439);
and U11550 (N_11550,N_11508,N_11445);
nand U11551 (N_11551,N_11494,N_11460);
and U11552 (N_11552,N_11435,N_11476);
nand U11553 (N_11553,N_11472,N_11454);
nor U11554 (N_11554,N_11468,N_11373);
xnor U11555 (N_11555,N_11500,N_11395);
nand U11556 (N_11556,N_11363,N_11505);
nor U11557 (N_11557,N_11461,N_11503);
nand U11558 (N_11558,N_11499,N_11437);
or U11559 (N_11559,N_11504,N_11492);
or U11560 (N_11560,N_11419,N_11441);
nor U11561 (N_11561,N_11424,N_11498);
nand U11562 (N_11562,N_11416,N_11368);
xnor U11563 (N_11563,N_11387,N_11432);
nor U11564 (N_11564,N_11447,N_11462);
nor U11565 (N_11565,N_11513,N_11433);
or U11566 (N_11566,N_11434,N_11475);
nand U11567 (N_11567,N_11390,N_11474);
and U11568 (N_11568,N_11371,N_11495);
xnor U11569 (N_11569,N_11514,N_11497);
and U11570 (N_11570,N_11396,N_11369);
and U11571 (N_11571,N_11457,N_11490);
nand U11572 (N_11572,N_11440,N_11484);
or U11573 (N_11573,N_11444,N_11406);
or U11574 (N_11574,N_11471,N_11517);
nand U11575 (N_11575,N_11413,N_11470);
nor U11576 (N_11576,N_11438,N_11430);
xor U11577 (N_11577,N_11399,N_11515);
xnor U11578 (N_11578,N_11459,N_11512);
nor U11579 (N_11579,N_11436,N_11391);
or U11580 (N_11580,N_11516,N_11415);
or U11581 (N_11581,N_11487,N_11502);
xnor U11582 (N_11582,N_11501,N_11385);
or U11583 (N_11583,N_11453,N_11364);
nor U11584 (N_11584,N_11389,N_11456);
or U11585 (N_11585,N_11400,N_11509);
nor U11586 (N_11586,N_11386,N_11405);
or U11587 (N_11587,N_11360,N_11383);
or U11588 (N_11588,N_11465,N_11408);
and U11589 (N_11589,N_11361,N_11370);
xnor U11590 (N_11590,N_11481,N_11467);
and U11591 (N_11591,N_11379,N_11429);
and U11592 (N_11592,N_11480,N_11374);
nand U11593 (N_11593,N_11414,N_11451);
nand U11594 (N_11594,N_11384,N_11417);
and U11595 (N_11595,N_11478,N_11482);
and U11596 (N_11596,N_11388,N_11449);
nand U11597 (N_11597,N_11380,N_11477);
nor U11598 (N_11598,N_11428,N_11420);
nor U11599 (N_11599,N_11473,N_11466);
nand U11600 (N_11600,N_11482,N_11451);
or U11601 (N_11601,N_11459,N_11502);
nor U11602 (N_11602,N_11480,N_11496);
and U11603 (N_11603,N_11467,N_11504);
or U11604 (N_11604,N_11399,N_11398);
or U11605 (N_11605,N_11443,N_11395);
and U11606 (N_11606,N_11456,N_11421);
nand U11607 (N_11607,N_11363,N_11368);
nand U11608 (N_11608,N_11369,N_11409);
nand U11609 (N_11609,N_11476,N_11364);
xnor U11610 (N_11610,N_11438,N_11513);
or U11611 (N_11611,N_11479,N_11514);
nor U11612 (N_11612,N_11502,N_11414);
nor U11613 (N_11613,N_11504,N_11493);
and U11614 (N_11614,N_11453,N_11394);
or U11615 (N_11615,N_11434,N_11423);
or U11616 (N_11616,N_11519,N_11415);
and U11617 (N_11617,N_11503,N_11452);
and U11618 (N_11618,N_11419,N_11442);
nand U11619 (N_11619,N_11501,N_11454);
xnor U11620 (N_11620,N_11428,N_11412);
nor U11621 (N_11621,N_11478,N_11372);
nand U11622 (N_11622,N_11485,N_11381);
nand U11623 (N_11623,N_11492,N_11500);
and U11624 (N_11624,N_11426,N_11419);
and U11625 (N_11625,N_11494,N_11451);
xor U11626 (N_11626,N_11381,N_11421);
xnor U11627 (N_11627,N_11502,N_11496);
or U11628 (N_11628,N_11441,N_11469);
nand U11629 (N_11629,N_11406,N_11440);
or U11630 (N_11630,N_11517,N_11509);
nand U11631 (N_11631,N_11480,N_11366);
nor U11632 (N_11632,N_11398,N_11447);
and U11633 (N_11633,N_11519,N_11399);
nand U11634 (N_11634,N_11434,N_11393);
or U11635 (N_11635,N_11511,N_11502);
nand U11636 (N_11636,N_11390,N_11444);
xnor U11637 (N_11637,N_11386,N_11460);
xor U11638 (N_11638,N_11514,N_11400);
or U11639 (N_11639,N_11409,N_11467);
nor U11640 (N_11640,N_11454,N_11391);
nand U11641 (N_11641,N_11402,N_11463);
or U11642 (N_11642,N_11370,N_11385);
xnor U11643 (N_11643,N_11498,N_11486);
and U11644 (N_11644,N_11457,N_11433);
and U11645 (N_11645,N_11401,N_11459);
nor U11646 (N_11646,N_11447,N_11482);
and U11647 (N_11647,N_11377,N_11390);
and U11648 (N_11648,N_11484,N_11514);
and U11649 (N_11649,N_11381,N_11503);
xnor U11650 (N_11650,N_11479,N_11461);
nand U11651 (N_11651,N_11503,N_11422);
xor U11652 (N_11652,N_11445,N_11381);
or U11653 (N_11653,N_11422,N_11466);
xor U11654 (N_11654,N_11475,N_11439);
nand U11655 (N_11655,N_11449,N_11378);
or U11656 (N_11656,N_11477,N_11377);
nor U11657 (N_11657,N_11367,N_11360);
nand U11658 (N_11658,N_11406,N_11464);
or U11659 (N_11659,N_11432,N_11363);
nand U11660 (N_11660,N_11477,N_11379);
nor U11661 (N_11661,N_11367,N_11497);
and U11662 (N_11662,N_11446,N_11421);
or U11663 (N_11663,N_11405,N_11451);
and U11664 (N_11664,N_11493,N_11508);
nor U11665 (N_11665,N_11363,N_11471);
nor U11666 (N_11666,N_11388,N_11509);
and U11667 (N_11667,N_11495,N_11461);
and U11668 (N_11668,N_11451,N_11372);
or U11669 (N_11669,N_11437,N_11484);
nor U11670 (N_11670,N_11445,N_11412);
nand U11671 (N_11671,N_11417,N_11431);
nor U11672 (N_11672,N_11488,N_11417);
or U11673 (N_11673,N_11468,N_11405);
xnor U11674 (N_11674,N_11455,N_11486);
nand U11675 (N_11675,N_11414,N_11469);
and U11676 (N_11676,N_11436,N_11457);
xor U11677 (N_11677,N_11463,N_11481);
xor U11678 (N_11678,N_11361,N_11410);
xor U11679 (N_11679,N_11444,N_11481);
and U11680 (N_11680,N_11611,N_11583);
nor U11681 (N_11681,N_11528,N_11633);
xor U11682 (N_11682,N_11672,N_11588);
and U11683 (N_11683,N_11658,N_11553);
nor U11684 (N_11684,N_11679,N_11634);
nand U11685 (N_11685,N_11655,N_11545);
and U11686 (N_11686,N_11638,N_11676);
xnor U11687 (N_11687,N_11582,N_11656);
nand U11688 (N_11688,N_11620,N_11570);
nand U11689 (N_11689,N_11636,N_11657);
xor U11690 (N_11690,N_11563,N_11617);
nand U11691 (N_11691,N_11542,N_11642);
nor U11692 (N_11692,N_11590,N_11576);
xnor U11693 (N_11693,N_11623,N_11541);
xnor U11694 (N_11694,N_11674,N_11532);
or U11695 (N_11695,N_11549,N_11527);
nor U11696 (N_11696,N_11520,N_11529);
or U11697 (N_11697,N_11653,N_11561);
and U11698 (N_11698,N_11600,N_11578);
and U11699 (N_11699,N_11615,N_11643);
nand U11700 (N_11700,N_11585,N_11637);
nand U11701 (N_11701,N_11586,N_11622);
nand U11702 (N_11702,N_11651,N_11677);
xor U11703 (N_11703,N_11665,N_11612);
and U11704 (N_11704,N_11605,N_11571);
or U11705 (N_11705,N_11530,N_11670);
nand U11706 (N_11706,N_11628,N_11531);
nand U11707 (N_11707,N_11551,N_11543);
nand U11708 (N_11708,N_11522,N_11630);
and U11709 (N_11709,N_11648,N_11647);
and U11710 (N_11710,N_11629,N_11610);
and U11711 (N_11711,N_11552,N_11639);
or U11712 (N_11712,N_11624,N_11601);
or U11713 (N_11713,N_11604,N_11635);
xnor U11714 (N_11714,N_11618,N_11626);
nand U11715 (N_11715,N_11525,N_11556);
nor U11716 (N_11716,N_11593,N_11607);
nor U11717 (N_11717,N_11587,N_11538);
nor U11718 (N_11718,N_11641,N_11592);
nor U11719 (N_11719,N_11640,N_11540);
and U11720 (N_11720,N_11614,N_11663);
xor U11721 (N_11721,N_11631,N_11539);
xor U11722 (N_11722,N_11566,N_11535);
or U11723 (N_11723,N_11557,N_11548);
and U11724 (N_11724,N_11537,N_11565);
nor U11725 (N_11725,N_11569,N_11603);
xnor U11726 (N_11726,N_11568,N_11577);
or U11727 (N_11727,N_11567,N_11621);
and U11728 (N_11728,N_11564,N_11596);
and U11729 (N_11729,N_11533,N_11599);
and U11730 (N_11730,N_11609,N_11616);
or U11731 (N_11731,N_11597,N_11667);
and U11732 (N_11732,N_11544,N_11625);
nor U11733 (N_11733,N_11521,N_11524);
or U11734 (N_11734,N_11591,N_11652);
xnor U11735 (N_11735,N_11666,N_11560);
or U11736 (N_11736,N_11550,N_11606);
and U11737 (N_11737,N_11668,N_11673);
xnor U11738 (N_11738,N_11650,N_11574);
and U11739 (N_11739,N_11572,N_11660);
xor U11740 (N_11740,N_11654,N_11594);
nor U11741 (N_11741,N_11536,N_11547);
or U11742 (N_11742,N_11581,N_11555);
and U11743 (N_11743,N_11661,N_11598);
xor U11744 (N_11744,N_11575,N_11649);
xnor U11745 (N_11745,N_11627,N_11619);
or U11746 (N_11746,N_11526,N_11669);
nand U11747 (N_11747,N_11662,N_11678);
nor U11748 (N_11748,N_11613,N_11589);
xnor U11749 (N_11749,N_11645,N_11580);
or U11750 (N_11750,N_11595,N_11675);
nand U11751 (N_11751,N_11546,N_11671);
or U11752 (N_11752,N_11602,N_11659);
and U11753 (N_11753,N_11584,N_11646);
and U11754 (N_11754,N_11558,N_11523);
nand U11755 (N_11755,N_11534,N_11573);
or U11756 (N_11756,N_11664,N_11644);
nor U11757 (N_11757,N_11579,N_11632);
or U11758 (N_11758,N_11554,N_11559);
or U11759 (N_11759,N_11562,N_11608);
and U11760 (N_11760,N_11523,N_11632);
xor U11761 (N_11761,N_11601,N_11610);
nand U11762 (N_11762,N_11651,N_11593);
nand U11763 (N_11763,N_11664,N_11633);
nor U11764 (N_11764,N_11574,N_11625);
xnor U11765 (N_11765,N_11542,N_11677);
and U11766 (N_11766,N_11544,N_11570);
or U11767 (N_11767,N_11583,N_11607);
xnor U11768 (N_11768,N_11594,N_11604);
nand U11769 (N_11769,N_11609,N_11638);
or U11770 (N_11770,N_11555,N_11575);
and U11771 (N_11771,N_11552,N_11641);
nor U11772 (N_11772,N_11597,N_11578);
and U11773 (N_11773,N_11607,N_11544);
nor U11774 (N_11774,N_11636,N_11616);
or U11775 (N_11775,N_11522,N_11641);
and U11776 (N_11776,N_11585,N_11564);
nor U11777 (N_11777,N_11556,N_11577);
nand U11778 (N_11778,N_11602,N_11583);
xnor U11779 (N_11779,N_11657,N_11598);
nand U11780 (N_11780,N_11545,N_11530);
or U11781 (N_11781,N_11559,N_11522);
or U11782 (N_11782,N_11607,N_11674);
nand U11783 (N_11783,N_11524,N_11578);
or U11784 (N_11784,N_11551,N_11677);
and U11785 (N_11785,N_11549,N_11662);
nand U11786 (N_11786,N_11646,N_11671);
nor U11787 (N_11787,N_11640,N_11538);
or U11788 (N_11788,N_11545,N_11570);
xor U11789 (N_11789,N_11614,N_11669);
xor U11790 (N_11790,N_11633,N_11639);
or U11791 (N_11791,N_11648,N_11560);
xor U11792 (N_11792,N_11560,N_11612);
and U11793 (N_11793,N_11595,N_11616);
or U11794 (N_11794,N_11606,N_11540);
and U11795 (N_11795,N_11583,N_11633);
nand U11796 (N_11796,N_11534,N_11546);
or U11797 (N_11797,N_11576,N_11581);
nor U11798 (N_11798,N_11572,N_11523);
or U11799 (N_11799,N_11624,N_11610);
xnor U11800 (N_11800,N_11656,N_11625);
or U11801 (N_11801,N_11619,N_11636);
and U11802 (N_11802,N_11527,N_11671);
nand U11803 (N_11803,N_11579,N_11555);
nor U11804 (N_11804,N_11678,N_11644);
nor U11805 (N_11805,N_11556,N_11542);
nor U11806 (N_11806,N_11636,N_11679);
nor U11807 (N_11807,N_11532,N_11637);
or U11808 (N_11808,N_11543,N_11675);
nor U11809 (N_11809,N_11582,N_11611);
or U11810 (N_11810,N_11616,N_11637);
and U11811 (N_11811,N_11646,N_11649);
nand U11812 (N_11812,N_11653,N_11581);
and U11813 (N_11813,N_11642,N_11631);
or U11814 (N_11814,N_11570,N_11618);
nor U11815 (N_11815,N_11594,N_11535);
or U11816 (N_11816,N_11584,N_11590);
and U11817 (N_11817,N_11567,N_11589);
xor U11818 (N_11818,N_11616,N_11599);
nor U11819 (N_11819,N_11549,N_11587);
nand U11820 (N_11820,N_11582,N_11657);
or U11821 (N_11821,N_11532,N_11570);
nand U11822 (N_11822,N_11574,N_11669);
and U11823 (N_11823,N_11674,N_11675);
or U11824 (N_11824,N_11524,N_11540);
nor U11825 (N_11825,N_11589,N_11543);
xnor U11826 (N_11826,N_11539,N_11543);
and U11827 (N_11827,N_11552,N_11588);
and U11828 (N_11828,N_11535,N_11603);
nor U11829 (N_11829,N_11617,N_11627);
and U11830 (N_11830,N_11578,N_11567);
or U11831 (N_11831,N_11597,N_11674);
nand U11832 (N_11832,N_11641,N_11622);
nor U11833 (N_11833,N_11672,N_11619);
or U11834 (N_11834,N_11582,N_11647);
or U11835 (N_11835,N_11634,N_11631);
nor U11836 (N_11836,N_11568,N_11527);
nand U11837 (N_11837,N_11656,N_11673);
nand U11838 (N_11838,N_11562,N_11581);
nand U11839 (N_11839,N_11643,N_11555);
and U11840 (N_11840,N_11784,N_11744);
xor U11841 (N_11841,N_11776,N_11725);
xor U11842 (N_11842,N_11729,N_11785);
nor U11843 (N_11843,N_11794,N_11796);
nor U11844 (N_11844,N_11745,N_11734);
or U11845 (N_11845,N_11823,N_11737);
and U11846 (N_11846,N_11838,N_11686);
nand U11847 (N_11847,N_11791,N_11719);
nand U11848 (N_11848,N_11777,N_11773);
nor U11849 (N_11849,N_11748,N_11781);
and U11850 (N_11850,N_11795,N_11722);
xor U11851 (N_11851,N_11807,N_11752);
nor U11852 (N_11852,N_11782,N_11819);
and U11853 (N_11853,N_11695,N_11802);
nand U11854 (N_11854,N_11754,N_11790);
and U11855 (N_11855,N_11780,N_11835);
or U11856 (N_11856,N_11788,N_11820);
nor U11857 (N_11857,N_11713,N_11809);
and U11858 (N_11858,N_11724,N_11770);
nor U11859 (N_11859,N_11803,N_11825);
and U11860 (N_11860,N_11683,N_11694);
and U11861 (N_11861,N_11816,N_11743);
or U11862 (N_11862,N_11704,N_11710);
and U11863 (N_11863,N_11698,N_11757);
xnor U11864 (N_11864,N_11783,N_11834);
nand U11865 (N_11865,N_11800,N_11739);
xor U11866 (N_11866,N_11708,N_11736);
and U11867 (N_11867,N_11789,N_11700);
or U11868 (N_11868,N_11762,N_11755);
xnor U11869 (N_11869,N_11793,N_11684);
nor U11870 (N_11870,N_11830,N_11717);
and U11871 (N_11871,N_11828,N_11798);
nand U11872 (N_11872,N_11697,N_11772);
nor U11873 (N_11873,N_11814,N_11797);
xor U11874 (N_11874,N_11718,N_11693);
or U11875 (N_11875,N_11808,N_11758);
nand U11876 (N_11876,N_11681,N_11806);
xnor U11877 (N_11877,N_11760,N_11692);
nor U11878 (N_11878,N_11733,N_11716);
or U11879 (N_11879,N_11715,N_11742);
and U11880 (N_11880,N_11727,N_11741);
nand U11881 (N_11881,N_11767,N_11761);
or U11882 (N_11882,N_11766,N_11839);
or U11883 (N_11883,N_11735,N_11836);
nor U11884 (N_11884,N_11696,N_11801);
or U11885 (N_11885,N_11821,N_11827);
nand U11886 (N_11886,N_11706,N_11682);
nand U11887 (N_11887,N_11810,N_11813);
or U11888 (N_11888,N_11826,N_11711);
nand U11889 (N_11889,N_11832,N_11690);
nor U11890 (N_11890,N_11759,N_11732);
and U11891 (N_11891,N_11817,N_11756);
xor U11892 (N_11892,N_11799,N_11753);
and U11893 (N_11893,N_11815,N_11751);
or U11894 (N_11894,N_11764,N_11685);
nor U11895 (N_11895,N_11822,N_11831);
or U11896 (N_11896,N_11701,N_11699);
or U11897 (N_11897,N_11774,N_11786);
or U11898 (N_11898,N_11829,N_11721);
nor U11899 (N_11899,N_11689,N_11720);
and U11900 (N_11900,N_11728,N_11726);
and U11901 (N_11901,N_11804,N_11749);
nor U11902 (N_11902,N_11812,N_11723);
xnor U11903 (N_11903,N_11805,N_11771);
or U11904 (N_11904,N_11750,N_11818);
nor U11905 (N_11905,N_11769,N_11792);
nor U11906 (N_11906,N_11775,N_11768);
and U11907 (N_11907,N_11833,N_11779);
nor U11908 (N_11908,N_11731,N_11778);
or U11909 (N_11909,N_11687,N_11824);
nand U11910 (N_11910,N_11747,N_11746);
nand U11911 (N_11911,N_11705,N_11707);
xnor U11912 (N_11912,N_11738,N_11765);
and U11913 (N_11913,N_11703,N_11680);
nand U11914 (N_11914,N_11740,N_11709);
nor U11915 (N_11915,N_11702,N_11811);
or U11916 (N_11916,N_11763,N_11714);
xor U11917 (N_11917,N_11837,N_11712);
nand U11918 (N_11918,N_11730,N_11691);
xor U11919 (N_11919,N_11688,N_11787);
nand U11920 (N_11920,N_11727,N_11811);
or U11921 (N_11921,N_11757,N_11822);
xor U11922 (N_11922,N_11692,N_11748);
nor U11923 (N_11923,N_11801,N_11757);
nor U11924 (N_11924,N_11754,N_11786);
and U11925 (N_11925,N_11816,N_11723);
and U11926 (N_11926,N_11805,N_11765);
xor U11927 (N_11927,N_11813,N_11726);
or U11928 (N_11928,N_11817,N_11716);
and U11929 (N_11929,N_11746,N_11764);
nand U11930 (N_11930,N_11752,N_11715);
nor U11931 (N_11931,N_11691,N_11748);
nand U11932 (N_11932,N_11820,N_11838);
xor U11933 (N_11933,N_11799,N_11820);
nand U11934 (N_11934,N_11775,N_11745);
xnor U11935 (N_11935,N_11705,N_11808);
nor U11936 (N_11936,N_11682,N_11688);
nand U11937 (N_11937,N_11698,N_11706);
or U11938 (N_11938,N_11742,N_11806);
and U11939 (N_11939,N_11723,N_11684);
xor U11940 (N_11940,N_11751,N_11828);
and U11941 (N_11941,N_11749,N_11752);
or U11942 (N_11942,N_11712,N_11723);
and U11943 (N_11943,N_11790,N_11796);
or U11944 (N_11944,N_11714,N_11815);
or U11945 (N_11945,N_11729,N_11758);
or U11946 (N_11946,N_11723,N_11728);
and U11947 (N_11947,N_11751,N_11757);
nor U11948 (N_11948,N_11765,N_11767);
nand U11949 (N_11949,N_11817,N_11738);
xor U11950 (N_11950,N_11725,N_11728);
or U11951 (N_11951,N_11784,N_11758);
or U11952 (N_11952,N_11717,N_11829);
or U11953 (N_11953,N_11716,N_11685);
or U11954 (N_11954,N_11790,N_11708);
and U11955 (N_11955,N_11778,N_11746);
nor U11956 (N_11956,N_11810,N_11799);
xnor U11957 (N_11957,N_11723,N_11706);
xnor U11958 (N_11958,N_11724,N_11741);
xnor U11959 (N_11959,N_11774,N_11789);
nand U11960 (N_11960,N_11764,N_11769);
or U11961 (N_11961,N_11777,N_11774);
and U11962 (N_11962,N_11701,N_11724);
nand U11963 (N_11963,N_11821,N_11706);
nand U11964 (N_11964,N_11820,N_11680);
nor U11965 (N_11965,N_11732,N_11834);
xnor U11966 (N_11966,N_11693,N_11703);
xnor U11967 (N_11967,N_11749,N_11694);
xnor U11968 (N_11968,N_11816,N_11768);
and U11969 (N_11969,N_11764,N_11763);
or U11970 (N_11970,N_11712,N_11788);
xor U11971 (N_11971,N_11719,N_11706);
nand U11972 (N_11972,N_11821,N_11778);
and U11973 (N_11973,N_11699,N_11782);
and U11974 (N_11974,N_11683,N_11736);
or U11975 (N_11975,N_11825,N_11729);
nor U11976 (N_11976,N_11813,N_11738);
and U11977 (N_11977,N_11832,N_11719);
nand U11978 (N_11978,N_11797,N_11818);
or U11979 (N_11979,N_11838,N_11819);
xor U11980 (N_11980,N_11745,N_11710);
or U11981 (N_11981,N_11797,N_11713);
or U11982 (N_11982,N_11779,N_11685);
or U11983 (N_11983,N_11806,N_11724);
and U11984 (N_11984,N_11757,N_11780);
nor U11985 (N_11985,N_11811,N_11770);
nor U11986 (N_11986,N_11682,N_11808);
xor U11987 (N_11987,N_11768,N_11764);
or U11988 (N_11988,N_11715,N_11793);
nor U11989 (N_11989,N_11771,N_11756);
nand U11990 (N_11990,N_11823,N_11747);
and U11991 (N_11991,N_11717,N_11706);
xor U11992 (N_11992,N_11823,N_11782);
nand U11993 (N_11993,N_11735,N_11822);
or U11994 (N_11994,N_11810,N_11831);
and U11995 (N_11995,N_11822,N_11702);
xnor U11996 (N_11996,N_11783,N_11774);
nor U11997 (N_11997,N_11789,N_11733);
or U11998 (N_11998,N_11792,N_11830);
nor U11999 (N_11999,N_11710,N_11753);
nand U12000 (N_12000,N_11882,N_11851);
nor U12001 (N_12001,N_11894,N_11883);
xor U12002 (N_12002,N_11867,N_11937);
xnor U12003 (N_12003,N_11887,N_11999);
or U12004 (N_12004,N_11860,N_11929);
nand U12005 (N_12005,N_11903,N_11840);
or U12006 (N_12006,N_11971,N_11873);
nor U12007 (N_12007,N_11977,N_11944);
nor U12008 (N_12008,N_11920,N_11962);
or U12009 (N_12009,N_11906,N_11921);
or U12010 (N_12010,N_11852,N_11913);
xor U12011 (N_12011,N_11948,N_11998);
and U12012 (N_12012,N_11924,N_11980);
nor U12013 (N_12013,N_11861,N_11933);
and U12014 (N_12014,N_11985,N_11952);
xor U12015 (N_12015,N_11848,N_11915);
and U12016 (N_12016,N_11969,N_11931);
and U12017 (N_12017,N_11947,N_11982);
or U12018 (N_12018,N_11935,N_11918);
nor U12019 (N_12019,N_11951,N_11890);
and U12020 (N_12020,N_11871,N_11965);
and U12021 (N_12021,N_11925,N_11934);
or U12022 (N_12022,N_11919,N_11912);
nand U12023 (N_12023,N_11922,N_11870);
nand U12024 (N_12024,N_11943,N_11939);
and U12025 (N_12025,N_11895,N_11996);
xnor U12026 (N_12026,N_11897,N_11972);
xnor U12027 (N_12027,N_11955,N_11850);
nand U12028 (N_12028,N_11917,N_11988);
nor U12029 (N_12029,N_11875,N_11844);
nand U12030 (N_12030,N_11868,N_11940);
nand U12031 (N_12031,N_11841,N_11849);
nand U12032 (N_12032,N_11909,N_11884);
and U12033 (N_12033,N_11879,N_11872);
nand U12034 (N_12034,N_11994,N_11888);
nand U12035 (N_12035,N_11869,N_11910);
or U12036 (N_12036,N_11855,N_11974);
nor U12037 (N_12037,N_11953,N_11949);
xor U12038 (N_12038,N_11853,N_11865);
and U12039 (N_12039,N_11958,N_11970);
nor U12040 (N_12040,N_11968,N_11950);
and U12041 (N_12041,N_11960,N_11959);
or U12042 (N_12042,N_11901,N_11984);
xor U12043 (N_12043,N_11862,N_11889);
and U12044 (N_12044,N_11843,N_11926);
xor U12045 (N_12045,N_11956,N_11886);
or U12046 (N_12046,N_11945,N_11957);
xnor U12047 (N_12047,N_11993,N_11863);
nand U12048 (N_12048,N_11990,N_11846);
and U12049 (N_12049,N_11928,N_11842);
nor U12050 (N_12050,N_11991,N_11847);
nand U12051 (N_12051,N_11859,N_11881);
or U12052 (N_12052,N_11967,N_11992);
nor U12053 (N_12053,N_11979,N_11927);
nand U12054 (N_12054,N_11885,N_11942);
nor U12055 (N_12055,N_11973,N_11857);
xor U12056 (N_12056,N_11892,N_11966);
xor U12057 (N_12057,N_11954,N_11975);
and U12058 (N_12058,N_11900,N_11878);
xnor U12059 (N_12059,N_11854,N_11946);
nand U12060 (N_12060,N_11858,N_11941);
and U12061 (N_12061,N_11864,N_11930);
or U12062 (N_12062,N_11914,N_11891);
or U12063 (N_12063,N_11981,N_11963);
or U12064 (N_12064,N_11983,N_11902);
nor U12065 (N_12065,N_11899,N_11898);
or U12066 (N_12066,N_11876,N_11893);
or U12067 (N_12067,N_11916,N_11907);
nand U12068 (N_12068,N_11908,N_11932);
and U12069 (N_12069,N_11911,N_11997);
nor U12070 (N_12070,N_11905,N_11856);
xnor U12071 (N_12071,N_11936,N_11874);
and U12072 (N_12072,N_11877,N_11923);
nor U12073 (N_12073,N_11986,N_11978);
and U12074 (N_12074,N_11989,N_11866);
xor U12075 (N_12075,N_11964,N_11938);
nand U12076 (N_12076,N_11987,N_11845);
and U12077 (N_12077,N_11896,N_11961);
nand U12078 (N_12078,N_11904,N_11976);
nand U12079 (N_12079,N_11880,N_11995);
nand U12080 (N_12080,N_11959,N_11860);
or U12081 (N_12081,N_11912,N_11849);
and U12082 (N_12082,N_11995,N_11869);
xnor U12083 (N_12083,N_11963,N_11978);
and U12084 (N_12084,N_11977,N_11971);
nor U12085 (N_12085,N_11920,N_11929);
nor U12086 (N_12086,N_11987,N_11885);
xnor U12087 (N_12087,N_11937,N_11896);
nor U12088 (N_12088,N_11898,N_11903);
nor U12089 (N_12089,N_11933,N_11975);
xnor U12090 (N_12090,N_11969,N_11876);
nand U12091 (N_12091,N_11871,N_11901);
or U12092 (N_12092,N_11859,N_11907);
nor U12093 (N_12093,N_11883,N_11853);
nand U12094 (N_12094,N_11953,N_11911);
nor U12095 (N_12095,N_11854,N_11993);
nand U12096 (N_12096,N_11858,N_11848);
nand U12097 (N_12097,N_11961,N_11998);
or U12098 (N_12098,N_11847,N_11870);
nand U12099 (N_12099,N_11885,N_11995);
xor U12100 (N_12100,N_11887,N_11961);
and U12101 (N_12101,N_11940,N_11962);
xor U12102 (N_12102,N_11872,N_11873);
nor U12103 (N_12103,N_11943,N_11973);
nor U12104 (N_12104,N_11923,N_11908);
xnor U12105 (N_12105,N_11897,N_11892);
nand U12106 (N_12106,N_11916,N_11941);
nor U12107 (N_12107,N_11895,N_11985);
nor U12108 (N_12108,N_11850,N_11975);
or U12109 (N_12109,N_11933,N_11884);
nor U12110 (N_12110,N_11916,N_11936);
nor U12111 (N_12111,N_11953,N_11882);
or U12112 (N_12112,N_11951,N_11978);
xor U12113 (N_12113,N_11968,N_11873);
xnor U12114 (N_12114,N_11931,N_11985);
nand U12115 (N_12115,N_11906,N_11939);
or U12116 (N_12116,N_11906,N_11902);
or U12117 (N_12117,N_11985,N_11937);
and U12118 (N_12118,N_11966,N_11996);
and U12119 (N_12119,N_11851,N_11915);
and U12120 (N_12120,N_11939,N_11995);
and U12121 (N_12121,N_11985,N_11907);
and U12122 (N_12122,N_11873,N_11944);
and U12123 (N_12123,N_11883,N_11972);
or U12124 (N_12124,N_11954,N_11956);
or U12125 (N_12125,N_11974,N_11960);
or U12126 (N_12126,N_11909,N_11841);
nor U12127 (N_12127,N_11905,N_11974);
nor U12128 (N_12128,N_11980,N_11904);
nand U12129 (N_12129,N_11981,N_11890);
nor U12130 (N_12130,N_11844,N_11897);
or U12131 (N_12131,N_11977,N_11848);
xor U12132 (N_12132,N_11926,N_11991);
nor U12133 (N_12133,N_11883,N_11934);
nand U12134 (N_12134,N_11849,N_11885);
nand U12135 (N_12135,N_11997,N_11980);
and U12136 (N_12136,N_11906,N_11917);
nor U12137 (N_12137,N_11935,N_11968);
nor U12138 (N_12138,N_11882,N_11990);
nand U12139 (N_12139,N_11894,N_11906);
or U12140 (N_12140,N_11872,N_11840);
nor U12141 (N_12141,N_11988,N_11975);
nand U12142 (N_12142,N_11972,N_11997);
nand U12143 (N_12143,N_11907,N_11972);
nand U12144 (N_12144,N_11866,N_11952);
or U12145 (N_12145,N_11986,N_11846);
and U12146 (N_12146,N_11864,N_11842);
nand U12147 (N_12147,N_11928,N_11884);
or U12148 (N_12148,N_11934,N_11990);
or U12149 (N_12149,N_11864,N_11855);
nor U12150 (N_12150,N_11880,N_11958);
nand U12151 (N_12151,N_11931,N_11842);
nor U12152 (N_12152,N_11920,N_11901);
nand U12153 (N_12153,N_11948,N_11841);
xnor U12154 (N_12154,N_11851,N_11840);
xor U12155 (N_12155,N_11951,N_11864);
xor U12156 (N_12156,N_11928,N_11861);
nor U12157 (N_12157,N_11860,N_11843);
nand U12158 (N_12158,N_11885,N_11947);
nor U12159 (N_12159,N_11876,N_11859);
and U12160 (N_12160,N_12102,N_12031);
nand U12161 (N_12161,N_12079,N_12120);
and U12162 (N_12162,N_12116,N_12097);
and U12163 (N_12163,N_12080,N_12125);
and U12164 (N_12164,N_12137,N_12052);
and U12165 (N_12165,N_12155,N_12115);
nor U12166 (N_12166,N_12094,N_12127);
nand U12167 (N_12167,N_12009,N_12103);
nand U12168 (N_12168,N_12023,N_12071);
nand U12169 (N_12169,N_12068,N_12096);
xor U12170 (N_12170,N_12018,N_12133);
xnor U12171 (N_12171,N_12148,N_12064);
or U12172 (N_12172,N_12082,N_12063);
and U12173 (N_12173,N_12140,N_12123);
or U12174 (N_12174,N_12003,N_12026);
nand U12175 (N_12175,N_12114,N_12067);
nor U12176 (N_12176,N_12001,N_12065);
nand U12177 (N_12177,N_12154,N_12143);
and U12178 (N_12178,N_12016,N_12099);
xnor U12179 (N_12179,N_12104,N_12066);
or U12180 (N_12180,N_12044,N_12084);
nand U12181 (N_12181,N_12090,N_12083);
nor U12182 (N_12182,N_12017,N_12054);
xnor U12183 (N_12183,N_12135,N_12002);
or U12184 (N_12184,N_12076,N_12077);
nor U12185 (N_12185,N_12153,N_12110);
and U12186 (N_12186,N_12086,N_12000);
and U12187 (N_12187,N_12129,N_12046);
or U12188 (N_12188,N_12081,N_12058);
xnor U12189 (N_12189,N_12033,N_12147);
xnor U12190 (N_12190,N_12151,N_12139);
or U12191 (N_12191,N_12108,N_12075);
and U12192 (N_12192,N_12029,N_12078);
nand U12193 (N_12193,N_12109,N_12021);
xor U12194 (N_12194,N_12050,N_12022);
and U12195 (N_12195,N_12149,N_12034);
nand U12196 (N_12196,N_12117,N_12124);
xor U12197 (N_12197,N_12131,N_12118);
xnor U12198 (N_12198,N_12038,N_12025);
nand U12199 (N_12199,N_12037,N_12128);
and U12200 (N_12200,N_12056,N_12111);
nor U12201 (N_12201,N_12013,N_12152);
nand U12202 (N_12202,N_12014,N_12057);
xor U12203 (N_12203,N_12005,N_12091);
and U12204 (N_12204,N_12088,N_12010);
xnor U12205 (N_12205,N_12074,N_12055);
xor U12206 (N_12206,N_12136,N_12141);
xor U12207 (N_12207,N_12073,N_12012);
nor U12208 (N_12208,N_12007,N_12100);
nand U12209 (N_12209,N_12020,N_12011);
xnor U12210 (N_12210,N_12105,N_12047);
or U12211 (N_12211,N_12146,N_12035);
nand U12212 (N_12212,N_12028,N_12041);
nor U12213 (N_12213,N_12107,N_12145);
or U12214 (N_12214,N_12051,N_12126);
xor U12215 (N_12215,N_12142,N_12061);
xor U12216 (N_12216,N_12089,N_12039);
and U12217 (N_12217,N_12036,N_12015);
or U12218 (N_12218,N_12112,N_12159);
or U12219 (N_12219,N_12030,N_12042);
xnor U12220 (N_12220,N_12150,N_12092);
nand U12221 (N_12221,N_12119,N_12070);
xor U12222 (N_12222,N_12134,N_12062);
and U12223 (N_12223,N_12045,N_12132);
nor U12224 (N_12224,N_12072,N_12101);
nand U12225 (N_12225,N_12060,N_12156);
and U12226 (N_12226,N_12106,N_12144);
nor U12227 (N_12227,N_12157,N_12053);
and U12228 (N_12228,N_12043,N_12085);
nand U12229 (N_12229,N_12024,N_12113);
nor U12230 (N_12230,N_12008,N_12087);
xnor U12231 (N_12231,N_12006,N_12048);
or U12232 (N_12232,N_12098,N_12093);
xnor U12233 (N_12233,N_12049,N_12122);
xnor U12234 (N_12234,N_12040,N_12019);
or U12235 (N_12235,N_12004,N_12095);
nor U12236 (N_12236,N_12069,N_12032);
nand U12237 (N_12237,N_12121,N_12158);
nor U12238 (N_12238,N_12027,N_12130);
nor U12239 (N_12239,N_12138,N_12059);
nor U12240 (N_12240,N_12021,N_12033);
nand U12241 (N_12241,N_12027,N_12055);
or U12242 (N_12242,N_12028,N_12157);
nand U12243 (N_12243,N_12046,N_12130);
nand U12244 (N_12244,N_12055,N_12013);
nor U12245 (N_12245,N_12049,N_12025);
xor U12246 (N_12246,N_12052,N_12116);
nand U12247 (N_12247,N_12123,N_12085);
nor U12248 (N_12248,N_12055,N_12052);
xor U12249 (N_12249,N_12155,N_12013);
nor U12250 (N_12250,N_12017,N_12040);
nor U12251 (N_12251,N_12011,N_12082);
or U12252 (N_12252,N_12084,N_12104);
xnor U12253 (N_12253,N_12059,N_12078);
and U12254 (N_12254,N_12117,N_12029);
nor U12255 (N_12255,N_12091,N_12094);
nor U12256 (N_12256,N_12062,N_12034);
xor U12257 (N_12257,N_12021,N_12038);
nand U12258 (N_12258,N_12025,N_12096);
or U12259 (N_12259,N_12063,N_12133);
nand U12260 (N_12260,N_12005,N_12053);
nand U12261 (N_12261,N_12002,N_12043);
or U12262 (N_12262,N_12013,N_12068);
and U12263 (N_12263,N_12090,N_12117);
or U12264 (N_12264,N_12140,N_12103);
nand U12265 (N_12265,N_12085,N_12090);
nor U12266 (N_12266,N_12087,N_12153);
xor U12267 (N_12267,N_12059,N_12070);
or U12268 (N_12268,N_12010,N_12036);
or U12269 (N_12269,N_12155,N_12083);
nand U12270 (N_12270,N_12022,N_12035);
xnor U12271 (N_12271,N_12011,N_12148);
or U12272 (N_12272,N_12123,N_12105);
or U12273 (N_12273,N_12091,N_12117);
nand U12274 (N_12274,N_12046,N_12029);
xnor U12275 (N_12275,N_12005,N_12120);
or U12276 (N_12276,N_12024,N_12063);
nor U12277 (N_12277,N_12048,N_12149);
or U12278 (N_12278,N_12129,N_12154);
nand U12279 (N_12279,N_12131,N_12055);
or U12280 (N_12280,N_12147,N_12097);
nor U12281 (N_12281,N_12082,N_12049);
xor U12282 (N_12282,N_12095,N_12064);
nor U12283 (N_12283,N_12084,N_12148);
or U12284 (N_12284,N_12038,N_12045);
or U12285 (N_12285,N_12001,N_12130);
and U12286 (N_12286,N_12074,N_12148);
nor U12287 (N_12287,N_12128,N_12062);
or U12288 (N_12288,N_12150,N_12027);
nand U12289 (N_12289,N_12005,N_12121);
xor U12290 (N_12290,N_12159,N_12091);
and U12291 (N_12291,N_12116,N_12084);
or U12292 (N_12292,N_12127,N_12158);
xor U12293 (N_12293,N_12022,N_12021);
xor U12294 (N_12294,N_12043,N_12159);
or U12295 (N_12295,N_12088,N_12050);
or U12296 (N_12296,N_12021,N_12123);
or U12297 (N_12297,N_12096,N_12129);
and U12298 (N_12298,N_12032,N_12046);
or U12299 (N_12299,N_12157,N_12073);
or U12300 (N_12300,N_12122,N_12100);
and U12301 (N_12301,N_12027,N_12067);
xnor U12302 (N_12302,N_12155,N_12124);
and U12303 (N_12303,N_12052,N_12048);
nand U12304 (N_12304,N_12126,N_12145);
nand U12305 (N_12305,N_12037,N_12028);
nand U12306 (N_12306,N_12031,N_12044);
nor U12307 (N_12307,N_12152,N_12091);
and U12308 (N_12308,N_12046,N_12149);
xnor U12309 (N_12309,N_12059,N_12131);
or U12310 (N_12310,N_12072,N_12125);
nand U12311 (N_12311,N_12025,N_12155);
nor U12312 (N_12312,N_12147,N_12053);
nor U12313 (N_12313,N_12059,N_12093);
nand U12314 (N_12314,N_12032,N_12041);
or U12315 (N_12315,N_12089,N_12117);
or U12316 (N_12316,N_12081,N_12126);
nand U12317 (N_12317,N_12044,N_12119);
and U12318 (N_12318,N_12064,N_12017);
and U12319 (N_12319,N_12151,N_12100);
and U12320 (N_12320,N_12201,N_12303);
nand U12321 (N_12321,N_12206,N_12188);
and U12322 (N_12322,N_12179,N_12254);
xor U12323 (N_12323,N_12308,N_12287);
and U12324 (N_12324,N_12272,N_12279);
and U12325 (N_12325,N_12196,N_12277);
nor U12326 (N_12326,N_12205,N_12311);
or U12327 (N_12327,N_12191,N_12202);
and U12328 (N_12328,N_12235,N_12265);
and U12329 (N_12329,N_12247,N_12283);
and U12330 (N_12330,N_12227,N_12195);
or U12331 (N_12331,N_12302,N_12172);
nor U12332 (N_12332,N_12203,N_12298);
and U12333 (N_12333,N_12255,N_12305);
nand U12334 (N_12334,N_12192,N_12163);
xor U12335 (N_12335,N_12278,N_12187);
nand U12336 (N_12336,N_12160,N_12269);
xor U12337 (N_12337,N_12245,N_12292);
or U12338 (N_12338,N_12310,N_12171);
or U12339 (N_12339,N_12166,N_12319);
nor U12340 (N_12340,N_12197,N_12209);
nor U12341 (N_12341,N_12316,N_12271);
or U12342 (N_12342,N_12309,N_12304);
nor U12343 (N_12343,N_12264,N_12226);
or U12344 (N_12344,N_12299,N_12266);
and U12345 (N_12345,N_12216,N_12220);
or U12346 (N_12346,N_12244,N_12274);
xor U12347 (N_12347,N_12284,N_12248);
nor U12348 (N_12348,N_12260,N_12225);
nor U12349 (N_12349,N_12208,N_12259);
and U12350 (N_12350,N_12175,N_12290);
xor U12351 (N_12351,N_12210,N_12193);
xnor U12352 (N_12352,N_12189,N_12261);
or U12353 (N_12353,N_12176,N_12306);
xnor U12354 (N_12354,N_12240,N_12246);
nor U12355 (N_12355,N_12204,N_12293);
and U12356 (N_12356,N_12230,N_12281);
or U12357 (N_12357,N_12314,N_12317);
nor U12358 (N_12358,N_12174,N_12273);
or U12359 (N_12359,N_12252,N_12262);
nand U12360 (N_12360,N_12224,N_12291);
nor U12361 (N_12361,N_12180,N_12285);
nor U12362 (N_12362,N_12256,N_12268);
xnor U12363 (N_12363,N_12307,N_12250);
and U12364 (N_12364,N_12267,N_12286);
or U12365 (N_12365,N_12295,N_12270);
or U12366 (N_12366,N_12276,N_12289);
nand U12367 (N_12367,N_12184,N_12190);
xor U12368 (N_12368,N_12243,N_12238);
and U12369 (N_12369,N_12164,N_12239);
nor U12370 (N_12370,N_12237,N_12167);
or U12371 (N_12371,N_12258,N_12231);
xnor U12372 (N_12372,N_12182,N_12257);
xnor U12373 (N_12373,N_12318,N_12212);
or U12374 (N_12374,N_12242,N_12253);
and U12375 (N_12375,N_12297,N_12300);
or U12376 (N_12376,N_12301,N_12200);
xnor U12377 (N_12377,N_12282,N_12222);
and U12378 (N_12378,N_12236,N_12168);
nand U12379 (N_12379,N_12296,N_12161);
nand U12380 (N_12380,N_12207,N_12263);
and U12381 (N_12381,N_12186,N_12183);
and U12382 (N_12382,N_12165,N_12280);
xnor U12383 (N_12383,N_12223,N_12234);
nor U12384 (N_12384,N_12313,N_12173);
nand U12385 (N_12385,N_12198,N_12178);
and U12386 (N_12386,N_12169,N_12233);
or U12387 (N_12387,N_12221,N_12217);
nor U12388 (N_12388,N_12211,N_12194);
or U12389 (N_12389,N_12312,N_12275);
nand U12390 (N_12390,N_12232,N_12241);
xnor U12391 (N_12391,N_12218,N_12162);
or U12392 (N_12392,N_12213,N_12249);
xor U12393 (N_12393,N_12177,N_12219);
or U12394 (N_12394,N_12228,N_12229);
nor U12395 (N_12395,N_12294,N_12170);
or U12396 (N_12396,N_12214,N_12288);
or U12397 (N_12397,N_12185,N_12315);
nand U12398 (N_12398,N_12215,N_12251);
xor U12399 (N_12399,N_12181,N_12199);
xor U12400 (N_12400,N_12221,N_12271);
or U12401 (N_12401,N_12201,N_12176);
nand U12402 (N_12402,N_12301,N_12300);
nor U12403 (N_12403,N_12194,N_12301);
nor U12404 (N_12404,N_12305,N_12190);
nor U12405 (N_12405,N_12197,N_12193);
nand U12406 (N_12406,N_12312,N_12314);
xor U12407 (N_12407,N_12259,N_12183);
nor U12408 (N_12408,N_12318,N_12265);
or U12409 (N_12409,N_12203,N_12274);
or U12410 (N_12410,N_12313,N_12300);
nor U12411 (N_12411,N_12288,N_12304);
nand U12412 (N_12412,N_12234,N_12236);
or U12413 (N_12413,N_12313,N_12175);
nand U12414 (N_12414,N_12169,N_12163);
or U12415 (N_12415,N_12260,N_12235);
xor U12416 (N_12416,N_12170,N_12191);
nor U12417 (N_12417,N_12233,N_12184);
xnor U12418 (N_12418,N_12228,N_12266);
or U12419 (N_12419,N_12206,N_12258);
xor U12420 (N_12420,N_12266,N_12257);
nand U12421 (N_12421,N_12188,N_12180);
or U12422 (N_12422,N_12223,N_12240);
nand U12423 (N_12423,N_12253,N_12310);
nand U12424 (N_12424,N_12197,N_12295);
nand U12425 (N_12425,N_12208,N_12196);
or U12426 (N_12426,N_12283,N_12242);
xnor U12427 (N_12427,N_12298,N_12218);
and U12428 (N_12428,N_12247,N_12271);
or U12429 (N_12429,N_12182,N_12212);
nor U12430 (N_12430,N_12223,N_12262);
and U12431 (N_12431,N_12220,N_12192);
xnor U12432 (N_12432,N_12293,N_12249);
nand U12433 (N_12433,N_12306,N_12285);
nand U12434 (N_12434,N_12214,N_12271);
nand U12435 (N_12435,N_12229,N_12169);
nand U12436 (N_12436,N_12160,N_12255);
nor U12437 (N_12437,N_12172,N_12232);
or U12438 (N_12438,N_12290,N_12171);
and U12439 (N_12439,N_12194,N_12248);
and U12440 (N_12440,N_12209,N_12285);
nor U12441 (N_12441,N_12308,N_12254);
nor U12442 (N_12442,N_12177,N_12307);
xnor U12443 (N_12443,N_12313,N_12166);
and U12444 (N_12444,N_12202,N_12285);
xnor U12445 (N_12445,N_12199,N_12269);
and U12446 (N_12446,N_12231,N_12276);
or U12447 (N_12447,N_12308,N_12188);
nor U12448 (N_12448,N_12245,N_12168);
nor U12449 (N_12449,N_12241,N_12216);
xnor U12450 (N_12450,N_12211,N_12272);
nor U12451 (N_12451,N_12313,N_12253);
xor U12452 (N_12452,N_12163,N_12291);
and U12453 (N_12453,N_12312,N_12192);
nand U12454 (N_12454,N_12276,N_12303);
nand U12455 (N_12455,N_12291,N_12217);
and U12456 (N_12456,N_12270,N_12298);
and U12457 (N_12457,N_12309,N_12250);
nor U12458 (N_12458,N_12225,N_12161);
nor U12459 (N_12459,N_12226,N_12166);
nor U12460 (N_12460,N_12213,N_12209);
nand U12461 (N_12461,N_12283,N_12224);
xnor U12462 (N_12462,N_12272,N_12182);
nor U12463 (N_12463,N_12226,N_12185);
and U12464 (N_12464,N_12209,N_12201);
nand U12465 (N_12465,N_12191,N_12291);
nand U12466 (N_12466,N_12198,N_12253);
and U12467 (N_12467,N_12307,N_12314);
xor U12468 (N_12468,N_12217,N_12302);
or U12469 (N_12469,N_12298,N_12236);
xnor U12470 (N_12470,N_12208,N_12308);
nor U12471 (N_12471,N_12240,N_12198);
or U12472 (N_12472,N_12255,N_12207);
and U12473 (N_12473,N_12167,N_12199);
nand U12474 (N_12474,N_12315,N_12236);
and U12475 (N_12475,N_12165,N_12302);
and U12476 (N_12476,N_12166,N_12244);
or U12477 (N_12477,N_12185,N_12316);
nor U12478 (N_12478,N_12198,N_12173);
nand U12479 (N_12479,N_12229,N_12289);
nor U12480 (N_12480,N_12473,N_12400);
or U12481 (N_12481,N_12438,N_12381);
nand U12482 (N_12482,N_12460,N_12322);
nand U12483 (N_12483,N_12335,N_12339);
nor U12484 (N_12484,N_12340,N_12467);
nor U12485 (N_12485,N_12437,N_12362);
xor U12486 (N_12486,N_12457,N_12398);
nor U12487 (N_12487,N_12336,N_12409);
nor U12488 (N_12488,N_12374,N_12359);
nor U12489 (N_12489,N_12380,N_12356);
or U12490 (N_12490,N_12401,N_12393);
nand U12491 (N_12491,N_12446,N_12430);
nand U12492 (N_12492,N_12447,N_12432);
nor U12493 (N_12493,N_12370,N_12453);
xnor U12494 (N_12494,N_12429,N_12358);
nand U12495 (N_12495,N_12441,N_12476);
or U12496 (N_12496,N_12406,N_12452);
and U12497 (N_12497,N_12385,N_12458);
and U12498 (N_12498,N_12348,N_12331);
and U12499 (N_12499,N_12355,N_12433);
and U12500 (N_12500,N_12407,N_12346);
nand U12501 (N_12501,N_12404,N_12361);
or U12502 (N_12502,N_12451,N_12450);
nor U12503 (N_12503,N_12320,N_12466);
nor U12504 (N_12504,N_12440,N_12412);
or U12505 (N_12505,N_12354,N_12352);
nand U12506 (N_12506,N_12428,N_12449);
xor U12507 (N_12507,N_12366,N_12454);
nand U12508 (N_12508,N_12479,N_12341);
xnor U12509 (N_12509,N_12367,N_12371);
nor U12510 (N_12510,N_12464,N_12329);
nor U12511 (N_12511,N_12465,N_12389);
xnor U12512 (N_12512,N_12388,N_12342);
xnor U12513 (N_12513,N_12394,N_12382);
nor U12514 (N_12514,N_12413,N_12363);
nor U12515 (N_12515,N_12416,N_12372);
or U12516 (N_12516,N_12425,N_12326);
and U12517 (N_12517,N_12375,N_12418);
and U12518 (N_12518,N_12330,N_12477);
xor U12519 (N_12519,N_12327,N_12419);
and U12520 (N_12520,N_12436,N_12334);
or U12521 (N_12521,N_12369,N_12420);
and U12522 (N_12522,N_12349,N_12325);
or U12523 (N_12523,N_12445,N_12468);
nand U12524 (N_12524,N_12396,N_12414);
and U12525 (N_12525,N_12455,N_12444);
and U12526 (N_12526,N_12377,N_12392);
xnor U12527 (N_12527,N_12360,N_12442);
xor U12528 (N_12528,N_12475,N_12390);
and U12529 (N_12529,N_12474,N_12345);
nor U12530 (N_12530,N_12422,N_12344);
and U12531 (N_12531,N_12373,N_12402);
nand U12532 (N_12532,N_12347,N_12383);
nand U12533 (N_12533,N_12386,N_12459);
nand U12534 (N_12534,N_12463,N_12461);
nand U12535 (N_12535,N_12368,N_12353);
nand U12536 (N_12536,N_12434,N_12378);
or U12537 (N_12537,N_12423,N_12338);
xor U12538 (N_12538,N_12376,N_12426);
nand U12539 (N_12539,N_12469,N_12343);
nand U12540 (N_12540,N_12328,N_12435);
xnor U12541 (N_12541,N_12364,N_12324);
xor U12542 (N_12542,N_12478,N_12421);
or U12543 (N_12543,N_12337,N_12456);
xnor U12544 (N_12544,N_12424,N_12365);
or U12545 (N_12545,N_12462,N_12391);
xor U12546 (N_12546,N_12411,N_12399);
xnor U12547 (N_12547,N_12332,N_12448);
nor U12548 (N_12548,N_12471,N_12351);
nor U12549 (N_12549,N_12403,N_12415);
nor U12550 (N_12550,N_12417,N_12410);
and U12551 (N_12551,N_12395,N_12397);
xor U12552 (N_12552,N_12379,N_12439);
and U12553 (N_12553,N_12333,N_12431);
or U12554 (N_12554,N_12408,N_12405);
and U12555 (N_12555,N_12470,N_12357);
xnor U12556 (N_12556,N_12427,N_12323);
xnor U12557 (N_12557,N_12387,N_12472);
and U12558 (N_12558,N_12321,N_12443);
nor U12559 (N_12559,N_12384,N_12350);
and U12560 (N_12560,N_12462,N_12386);
nor U12561 (N_12561,N_12335,N_12326);
nand U12562 (N_12562,N_12375,N_12427);
or U12563 (N_12563,N_12391,N_12351);
or U12564 (N_12564,N_12394,N_12396);
and U12565 (N_12565,N_12353,N_12474);
nand U12566 (N_12566,N_12469,N_12393);
and U12567 (N_12567,N_12321,N_12458);
xor U12568 (N_12568,N_12390,N_12479);
xor U12569 (N_12569,N_12439,N_12468);
nor U12570 (N_12570,N_12443,N_12447);
xnor U12571 (N_12571,N_12411,N_12356);
nor U12572 (N_12572,N_12451,N_12340);
xor U12573 (N_12573,N_12361,N_12369);
xor U12574 (N_12574,N_12460,N_12408);
and U12575 (N_12575,N_12412,N_12476);
nor U12576 (N_12576,N_12362,N_12363);
xor U12577 (N_12577,N_12393,N_12429);
nor U12578 (N_12578,N_12404,N_12427);
and U12579 (N_12579,N_12335,N_12410);
nand U12580 (N_12580,N_12409,N_12386);
nor U12581 (N_12581,N_12451,N_12390);
nand U12582 (N_12582,N_12372,N_12395);
nand U12583 (N_12583,N_12476,N_12370);
and U12584 (N_12584,N_12437,N_12431);
xnor U12585 (N_12585,N_12448,N_12328);
nand U12586 (N_12586,N_12448,N_12456);
and U12587 (N_12587,N_12364,N_12455);
and U12588 (N_12588,N_12456,N_12357);
or U12589 (N_12589,N_12425,N_12455);
or U12590 (N_12590,N_12385,N_12400);
or U12591 (N_12591,N_12367,N_12473);
nand U12592 (N_12592,N_12425,N_12468);
or U12593 (N_12593,N_12420,N_12323);
or U12594 (N_12594,N_12331,N_12472);
and U12595 (N_12595,N_12375,N_12430);
or U12596 (N_12596,N_12366,N_12411);
xnor U12597 (N_12597,N_12476,N_12329);
nand U12598 (N_12598,N_12473,N_12453);
or U12599 (N_12599,N_12340,N_12408);
nand U12600 (N_12600,N_12474,N_12375);
or U12601 (N_12601,N_12363,N_12378);
and U12602 (N_12602,N_12424,N_12370);
or U12603 (N_12603,N_12342,N_12345);
xnor U12604 (N_12604,N_12341,N_12347);
xor U12605 (N_12605,N_12327,N_12379);
and U12606 (N_12606,N_12478,N_12401);
nand U12607 (N_12607,N_12361,N_12336);
xnor U12608 (N_12608,N_12413,N_12343);
and U12609 (N_12609,N_12407,N_12413);
and U12610 (N_12610,N_12338,N_12346);
nor U12611 (N_12611,N_12402,N_12423);
and U12612 (N_12612,N_12467,N_12426);
or U12613 (N_12613,N_12347,N_12435);
and U12614 (N_12614,N_12449,N_12466);
nor U12615 (N_12615,N_12346,N_12402);
nor U12616 (N_12616,N_12434,N_12350);
nand U12617 (N_12617,N_12378,N_12447);
nand U12618 (N_12618,N_12446,N_12339);
xnor U12619 (N_12619,N_12412,N_12432);
nand U12620 (N_12620,N_12321,N_12423);
or U12621 (N_12621,N_12332,N_12343);
or U12622 (N_12622,N_12463,N_12367);
nand U12623 (N_12623,N_12368,N_12440);
and U12624 (N_12624,N_12405,N_12476);
xor U12625 (N_12625,N_12458,N_12405);
nor U12626 (N_12626,N_12410,N_12356);
nor U12627 (N_12627,N_12472,N_12360);
or U12628 (N_12628,N_12397,N_12430);
nand U12629 (N_12629,N_12377,N_12334);
or U12630 (N_12630,N_12356,N_12379);
xnor U12631 (N_12631,N_12373,N_12426);
nand U12632 (N_12632,N_12391,N_12375);
and U12633 (N_12633,N_12411,N_12409);
nor U12634 (N_12634,N_12390,N_12420);
xor U12635 (N_12635,N_12444,N_12380);
nor U12636 (N_12636,N_12349,N_12423);
and U12637 (N_12637,N_12375,N_12324);
xnor U12638 (N_12638,N_12457,N_12382);
nand U12639 (N_12639,N_12408,N_12339);
nand U12640 (N_12640,N_12608,N_12558);
and U12641 (N_12641,N_12520,N_12539);
xor U12642 (N_12642,N_12535,N_12487);
and U12643 (N_12643,N_12616,N_12540);
xor U12644 (N_12644,N_12497,N_12560);
nor U12645 (N_12645,N_12615,N_12514);
xor U12646 (N_12646,N_12585,N_12627);
nor U12647 (N_12647,N_12529,N_12511);
nor U12648 (N_12648,N_12552,N_12480);
xnor U12649 (N_12649,N_12619,N_12607);
nand U12650 (N_12650,N_12524,N_12574);
nand U12651 (N_12651,N_12617,N_12588);
nor U12652 (N_12652,N_12532,N_12629);
nand U12653 (N_12653,N_12569,N_12525);
nor U12654 (N_12654,N_12572,N_12559);
xnor U12655 (N_12655,N_12515,N_12519);
and U12656 (N_12656,N_12577,N_12634);
or U12657 (N_12657,N_12481,N_12489);
nor U12658 (N_12658,N_12562,N_12604);
nor U12659 (N_12659,N_12530,N_12492);
xnor U12660 (N_12660,N_12485,N_12486);
and U12661 (N_12661,N_12541,N_12606);
nand U12662 (N_12662,N_12533,N_12504);
and U12663 (N_12663,N_12591,N_12551);
and U12664 (N_12664,N_12547,N_12639);
or U12665 (N_12665,N_12488,N_12637);
and U12666 (N_12666,N_12605,N_12484);
and U12667 (N_12667,N_12502,N_12496);
or U12668 (N_12668,N_12596,N_12542);
and U12669 (N_12669,N_12581,N_12590);
nand U12670 (N_12670,N_12493,N_12509);
xor U12671 (N_12671,N_12550,N_12506);
nor U12672 (N_12672,N_12531,N_12490);
nand U12673 (N_12673,N_12614,N_12561);
or U12674 (N_12674,N_12512,N_12571);
or U12675 (N_12675,N_12554,N_12568);
xnor U12676 (N_12676,N_12587,N_12521);
nand U12677 (N_12677,N_12631,N_12618);
nand U12678 (N_12678,N_12513,N_12538);
nand U12679 (N_12679,N_12517,N_12602);
and U12680 (N_12680,N_12597,N_12621);
or U12681 (N_12681,N_12623,N_12546);
nor U12682 (N_12682,N_12491,N_12576);
or U12683 (N_12683,N_12545,N_12522);
nor U12684 (N_12684,N_12593,N_12635);
nor U12685 (N_12685,N_12483,N_12501);
or U12686 (N_12686,N_12638,N_12589);
nand U12687 (N_12687,N_12595,N_12573);
or U12688 (N_12688,N_12537,N_12570);
or U12689 (N_12689,N_12556,N_12523);
and U12690 (N_12690,N_12603,N_12527);
or U12691 (N_12691,N_12609,N_12613);
xnor U12692 (N_12692,N_12633,N_12536);
and U12693 (N_12693,N_12544,N_12620);
xor U12694 (N_12694,N_12636,N_12575);
or U12695 (N_12695,N_12630,N_12494);
and U12696 (N_12696,N_12495,N_12579);
nor U12697 (N_12697,N_12600,N_12586);
xor U12698 (N_12698,N_12516,N_12594);
and U12699 (N_12699,N_12625,N_12632);
nand U12700 (N_12700,N_12592,N_12528);
nor U12701 (N_12701,N_12611,N_12510);
and U12702 (N_12702,N_12564,N_12548);
nor U12703 (N_12703,N_12557,N_12505);
xor U12704 (N_12704,N_12555,N_12580);
nor U12705 (N_12705,N_12601,N_12518);
and U12706 (N_12706,N_12612,N_12622);
and U12707 (N_12707,N_12543,N_12628);
and U12708 (N_12708,N_12500,N_12507);
nand U12709 (N_12709,N_12499,N_12563);
and U12710 (N_12710,N_12503,N_12582);
xnor U12711 (N_12711,N_12626,N_12553);
xor U12712 (N_12712,N_12508,N_12610);
or U12713 (N_12713,N_12565,N_12598);
nand U12714 (N_12714,N_12584,N_12583);
nand U12715 (N_12715,N_12534,N_12624);
xnor U12716 (N_12716,N_12482,N_12549);
or U12717 (N_12717,N_12526,N_12498);
nor U12718 (N_12718,N_12578,N_12567);
nor U12719 (N_12719,N_12599,N_12566);
or U12720 (N_12720,N_12510,N_12589);
nand U12721 (N_12721,N_12631,N_12512);
or U12722 (N_12722,N_12484,N_12487);
nand U12723 (N_12723,N_12560,N_12572);
xor U12724 (N_12724,N_12579,N_12520);
nand U12725 (N_12725,N_12524,N_12493);
nand U12726 (N_12726,N_12485,N_12519);
or U12727 (N_12727,N_12499,N_12491);
xor U12728 (N_12728,N_12561,N_12618);
and U12729 (N_12729,N_12511,N_12492);
and U12730 (N_12730,N_12516,N_12499);
xnor U12731 (N_12731,N_12633,N_12558);
nand U12732 (N_12732,N_12570,N_12484);
nand U12733 (N_12733,N_12481,N_12534);
or U12734 (N_12734,N_12551,N_12509);
and U12735 (N_12735,N_12631,N_12508);
xnor U12736 (N_12736,N_12617,N_12601);
nand U12737 (N_12737,N_12531,N_12547);
xor U12738 (N_12738,N_12576,N_12488);
xnor U12739 (N_12739,N_12605,N_12616);
nand U12740 (N_12740,N_12631,N_12497);
nand U12741 (N_12741,N_12605,N_12573);
and U12742 (N_12742,N_12605,N_12539);
or U12743 (N_12743,N_12534,N_12510);
or U12744 (N_12744,N_12618,N_12592);
and U12745 (N_12745,N_12597,N_12589);
or U12746 (N_12746,N_12543,N_12490);
nor U12747 (N_12747,N_12548,N_12483);
and U12748 (N_12748,N_12626,N_12614);
or U12749 (N_12749,N_12501,N_12517);
and U12750 (N_12750,N_12598,N_12619);
nor U12751 (N_12751,N_12632,N_12557);
nor U12752 (N_12752,N_12614,N_12551);
nand U12753 (N_12753,N_12506,N_12623);
and U12754 (N_12754,N_12579,N_12636);
nor U12755 (N_12755,N_12636,N_12550);
or U12756 (N_12756,N_12521,N_12487);
and U12757 (N_12757,N_12512,N_12602);
nand U12758 (N_12758,N_12516,N_12591);
nand U12759 (N_12759,N_12587,N_12619);
xnor U12760 (N_12760,N_12595,N_12537);
xor U12761 (N_12761,N_12484,N_12556);
nor U12762 (N_12762,N_12546,N_12552);
xor U12763 (N_12763,N_12606,N_12561);
xnor U12764 (N_12764,N_12538,N_12620);
xnor U12765 (N_12765,N_12595,N_12605);
xor U12766 (N_12766,N_12480,N_12530);
nand U12767 (N_12767,N_12525,N_12496);
or U12768 (N_12768,N_12634,N_12636);
nor U12769 (N_12769,N_12631,N_12627);
nand U12770 (N_12770,N_12592,N_12632);
nand U12771 (N_12771,N_12520,N_12573);
nor U12772 (N_12772,N_12527,N_12534);
nor U12773 (N_12773,N_12489,N_12486);
nand U12774 (N_12774,N_12536,N_12565);
and U12775 (N_12775,N_12613,N_12501);
xnor U12776 (N_12776,N_12528,N_12566);
xor U12777 (N_12777,N_12485,N_12503);
xor U12778 (N_12778,N_12615,N_12535);
xor U12779 (N_12779,N_12492,N_12634);
nor U12780 (N_12780,N_12627,N_12536);
xor U12781 (N_12781,N_12516,N_12605);
nand U12782 (N_12782,N_12540,N_12613);
and U12783 (N_12783,N_12534,N_12603);
nor U12784 (N_12784,N_12498,N_12537);
nor U12785 (N_12785,N_12595,N_12623);
or U12786 (N_12786,N_12520,N_12612);
nand U12787 (N_12787,N_12623,N_12534);
or U12788 (N_12788,N_12636,N_12582);
xnor U12789 (N_12789,N_12516,N_12502);
nor U12790 (N_12790,N_12488,N_12554);
and U12791 (N_12791,N_12612,N_12511);
xor U12792 (N_12792,N_12611,N_12582);
or U12793 (N_12793,N_12596,N_12574);
nand U12794 (N_12794,N_12586,N_12574);
nor U12795 (N_12795,N_12481,N_12576);
nand U12796 (N_12796,N_12542,N_12605);
nand U12797 (N_12797,N_12574,N_12566);
xnor U12798 (N_12798,N_12595,N_12486);
xor U12799 (N_12799,N_12508,N_12637);
and U12800 (N_12800,N_12797,N_12759);
or U12801 (N_12801,N_12660,N_12670);
nand U12802 (N_12802,N_12745,N_12724);
xor U12803 (N_12803,N_12756,N_12699);
nand U12804 (N_12804,N_12694,N_12776);
or U12805 (N_12805,N_12781,N_12738);
xor U12806 (N_12806,N_12767,N_12741);
xor U12807 (N_12807,N_12731,N_12791);
xnor U12808 (N_12808,N_12760,N_12779);
and U12809 (N_12809,N_12720,N_12763);
and U12810 (N_12810,N_12689,N_12790);
nor U12811 (N_12811,N_12798,N_12751);
nand U12812 (N_12812,N_12769,N_12764);
and U12813 (N_12813,N_12685,N_12642);
nor U12814 (N_12814,N_12799,N_12795);
nor U12815 (N_12815,N_12677,N_12789);
xor U12816 (N_12816,N_12770,N_12723);
or U12817 (N_12817,N_12754,N_12659);
nand U12818 (N_12818,N_12717,N_12655);
nand U12819 (N_12819,N_12713,N_12698);
nand U12820 (N_12820,N_12705,N_12788);
or U12821 (N_12821,N_12703,N_12786);
xnor U12822 (N_12822,N_12712,N_12704);
nand U12823 (N_12823,N_12701,N_12708);
nand U12824 (N_12824,N_12785,N_12796);
nand U12825 (N_12825,N_12772,N_12755);
or U12826 (N_12826,N_12707,N_12729);
and U12827 (N_12827,N_12671,N_12710);
xor U12828 (N_12828,N_12647,N_12657);
and U12829 (N_12829,N_12641,N_12679);
and U12830 (N_12830,N_12654,N_12652);
xnor U12831 (N_12831,N_12664,N_12761);
or U12832 (N_12832,N_12743,N_12750);
nor U12833 (N_12833,N_12669,N_12658);
nand U12834 (N_12834,N_12780,N_12668);
and U12835 (N_12835,N_12653,N_12722);
or U12836 (N_12836,N_12691,N_12680);
xnor U12837 (N_12837,N_12687,N_12681);
nand U12838 (N_12838,N_12700,N_12739);
nand U12839 (N_12839,N_12673,N_12674);
and U12840 (N_12840,N_12640,N_12648);
nand U12841 (N_12841,N_12771,N_12778);
xnor U12842 (N_12842,N_12676,N_12725);
nor U12843 (N_12843,N_12646,N_12715);
and U12844 (N_12844,N_12783,N_12742);
or U12845 (N_12845,N_12716,N_12721);
nor U12846 (N_12846,N_12645,N_12726);
nand U12847 (N_12847,N_12749,N_12667);
nor U12848 (N_12848,N_12686,N_12736);
nand U12849 (N_12849,N_12782,N_12768);
nor U12850 (N_12850,N_12794,N_12651);
or U12851 (N_12851,N_12650,N_12682);
nor U12852 (N_12852,N_12662,N_12683);
xor U12853 (N_12853,N_12695,N_12727);
nand U12854 (N_12854,N_12643,N_12787);
and U12855 (N_12855,N_12784,N_12661);
xnor U12856 (N_12856,N_12684,N_12762);
and U12857 (N_12857,N_12649,N_12714);
or U12858 (N_12858,N_12777,N_12678);
and U12859 (N_12859,N_12792,N_12752);
and U12860 (N_12860,N_12663,N_12697);
xnor U12861 (N_12861,N_12735,N_12711);
and U12862 (N_12862,N_12718,N_12737);
nor U12863 (N_12863,N_12719,N_12734);
nand U12864 (N_12864,N_12692,N_12656);
and U12865 (N_12865,N_12665,N_12696);
or U12866 (N_12866,N_12765,N_12644);
nand U12867 (N_12867,N_12774,N_12746);
nand U12868 (N_12868,N_12730,N_12666);
xor U12869 (N_12869,N_12693,N_12675);
nand U12870 (N_12870,N_12753,N_12728);
nor U12871 (N_12871,N_12793,N_12706);
nor U12872 (N_12872,N_12744,N_12747);
and U12873 (N_12873,N_12766,N_12758);
and U12874 (N_12874,N_12757,N_12775);
and U12875 (N_12875,N_12688,N_12672);
nor U12876 (N_12876,N_12748,N_12733);
nor U12877 (N_12877,N_12740,N_12690);
and U12878 (N_12878,N_12773,N_12732);
or U12879 (N_12879,N_12709,N_12702);
nand U12880 (N_12880,N_12680,N_12714);
or U12881 (N_12881,N_12774,N_12669);
xor U12882 (N_12882,N_12640,N_12795);
nand U12883 (N_12883,N_12723,N_12690);
or U12884 (N_12884,N_12673,N_12659);
or U12885 (N_12885,N_12779,N_12689);
nor U12886 (N_12886,N_12659,N_12787);
and U12887 (N_12887,N_12689,N_12774);
nand U12888 (N_12888,N_12678,N_12699);
xor U12889 (N_12889,N_12747,N_12756);
xnor U12890 (N_12890,N_12798,N_12688);
nand U12891 (N_12891,N_12677,N_12791);
nor U12892 (N_12892,N_12755,N_12751);
nor U12893 (N_12893,N_12795,N_12721);
or U12894 (N_12894,N_12687,N_12790);
nor U12895 (N_12895,N_12760,N_12753);
xnor U12896 (N_12896,N_12659,N_12735);
nor U12897 (N_12897,N_12746,N_12748);
nor U12898 (N_12898,N_12660,N_12788);
nor U12899 (N_12899,N_12727,N_12744);
nand U12900 (N_12900,N_12689,N_12752);
nand U12901 (N_12901,N_12710,N_12694);
nor U12902 (N_12902,N_12651,N_12714);
nand U12903 (N_12903,N_12797,N_12642);
nor U12904 (N_12904,N_12777,N_12650);
nand U12905 (N_12905,N_12731,N_12740);
and U12906 (N_12906,N_12694,N_12745);
nand U12907 (N_12907,N_12670,N_12715);
nor U12908 (N_12908,N_12686,N_12646);
nor U12909 (N_12909,N_12691,N_12756);
nand U12910 (N_12910,N_12709,N_12725);
xor U12911 (N_12911,N_12764,N_12691);
or U12912 (N_12912,N_12736,N_12717);
xnor U12913 (N_12913,N_12770,N_12685);
nand U12914 (N_12914,N_12795,N_12745);
or U12915 (N_12915,N_12759,N_12662);
nand U12916 (N_12916,N_12730,N_12739);
xor U12917 (N_12917,N_12673,N_12757);
nand U12918 (N_12918,N_12660,N_12725);
nand U12919 (N_12919,N_12791,N_12669);
nand U12920 (N_12920,N_12767,N_12745);
and U12921 (N_12921,N_12690,N_12677);
nand U12922 (N_12922,N_12784,N_12702);
or U12923 (N_12923,N_12654,N_12750);
nand U12924 (N_12924,N_12773,N_12721);
nor U12925 (N_12925,N_12767,N_12655);
and U12926 (N_12926,N_12730,N_12770);
nor U12927 (N_12927,N_12690,N_12729);
xnor U12928 (N_12928,N_12784,N_12699);
or U12929 (N_12929,N_12661,N_12684);
nand U12930 (N_12930,N_12787,N_12711);
nand U12931 (N_12931,N_12778,N_12713);
and U12932 (N_12932,N_12751,N_12773);
xnor U12933 (N_12933,N_12768,N_12755);
and U12934 (N_12934,N_12763,N_12673);
nand U12935 (N_12935,N_12778,N_12649);
and U12936 (N_12936,N_12748,N_12677);
and U12937 (N_12937,N_12747,N_12738);
nor U12938 (N_12938,N_12727,N_12767);
nand U12939 (N_12939,N_12698,N_12787);
or U12940 (N_12940,N_12759,N_12656);
nor U12941 (N_12941,N_12649,N_12780);
or U12942 (N_12942,N_12712,N_12725);
and U12943 (N_12943,N_12661,N_12746);
and U12944 (N_12944,N_12788,N_12791);
nor U12945 (N_12945,N_12650,N_12739);
nand U12946 (N_12946,N_12762,N_12782);
or U12947 (N_12947,N_12716,N_12742);
and U12948 (N_12948,N_12784,N_12692);
nor U12949 (N_12949,N_12785,N_12709);
nor U12950 (N_12950,N_12655,N_12761);
xor U12951 (N_12951,N_12699,N_12783);
and U12952 (N_12952,N_12712,N_12663);
nor U12953 (N_12953,N_12681,N_12780);
or U12954 (N_12954,N_12732,N_12786);
or U12955 (N_12955,N_12680,N_12681);
nand U12956 (N_12956,N_12736,N_12791);
nand U12957 (N_12957,N_12711,N_12766);
and U12958 (N_12958,N_12768,N_12772);
or U12959 (N_12959,N_12662,N_12654);
and U12960 (N_12960,N_12889,N_12878);
nand U12961 (N_12961,N_12944,N_12868);
nor U12962 (N_12962,N_12920,N_12946);
nand U12963 (N_12963,N_12871,N_12882);
or U12964 (N_12964,N_12805,N_12851);
xor U12965 (N_12965,N_12822,N_12865);
xnor U12966 (N_12966,N_12834,N_12823);
or U12967 (N_12967,N_12890,N_12840);
nand U12968 (N_12968,N_12828,N_12810);
nor U12969 (N_12969,N_12912,N_12895);
nor U12970 (N_12970,N_12813,N_12854);
nor U12971 (N_12971,N_12869,N_12837);
nor U12972 (N_12972,N_12941,N_12943);
nor U12973 (N_12973,N_12959,N_12860);
nor U12974 (N_12974,N_12926,N_12815);
and U12975 (N_12975,N_12826,N_12929);
nand U12976 (N_12976,N_12887,N_12803);
and U12977 (N_12977,N_12931,N_12948);
xor U12978 (N_12978,N_12885,N_12924);
nand U12979 (N_12979,N_12855,N_12893);
nor U12980 (N_12980,N_12872,N_12807);
nor U12981 (N_12981,N_12870,N_12888);
xor U12982 (N_12982,N_12945,N_12915);
or U12983 (N_12983,N_12841,N_12910);
nand U12984 (N_12984,N_12932,N_12938);
nand U12985 (N_12985,N_12809,N_12853);
xor U12986 (N_12986,N_12858,N_12862);
and U12987 (N_12987,N_12914,N_12825);
and U12988 (N_12988,N_12843,N_12874);
nand U12989 (N_12989,N_12952,N_12824);
or U12990 (N_12990,N_12867,N_12933);
nand U12991 (N_12991,N_12886,N_12901);
xor U12992 (N_12992,N_12935,N_12896);
and U12993 (N_12993,N_12849,N_12930);
and U12994 (N_12994,N_12908,N_12831);
and U12995 (N_12995,N_12922,N_12953);
or U12996 (N_12996,N_12898,N_12857);
nand U12997 (N_12997,N_12835,N_12934);
nand U12998 (N_12998,N_12808,N_12917);
xor U12999 (N_12999,N_12838,N_12847);
and U13000 (N_13000,N_12942,N_12883);
nor U13001 (N_13001,N_12906,N_12864);
or U13002 (N_13002,N_12909,N_12891);
xnor U13003 (N_13003,N_12881,N_12859);
nor U13004 (N_13004,N_12925,N_12830);
nand U13005 (N_13005,N_12844,N_12816);
or U13006 (N_13006,N_12812,N_12875);
xor U13007 (N_13007,N_12877,N_12905);
xnor U13008 (N_13008,N_12897,N_12928);
nor U13009 (N_13009,N_12842,N_12940);
xnor U13010 (N_13010,N_12818,N_12845);
xnor U13011 (N_13011,N_12800,N_12956);
nor U13012 (N_13012,N_12879,N_12923);
or U13013 (N_13013,N_12902,N_12957);
xnor U13014 (N_13014,N_12900,N_12866);
xor U13015 (N_13015,N_12819,N_12904);
xnor U13016 (N_13016,N_12829,N_12846);
and U13017 (N_13017,N_12958,N_12913);
nand U13018 (N_13018,N_12947,N_12833);
nor U13019 (N_13019,N_12873,N_12950);
nand U13020 (N_13020,N_12949,N_12839);
or U13021 (N_13021,N_12907,N_12821);
nand U13022 (N_13022,N_12911,N_12919);
nor U13023 (N_13023,N_12899,N_12861);
or U13024 (N_13024,N_12850,N_12836);
or U13025 (N_13025,N_12852,N_12916);
and U13026 (N_13026,N_12811,N_12806);
nand U13027 (N_13027,N_12863,N_12804);
or U13028 (N_13028,N_12951,N_12955);
nand U13029 (N_13029,N_12880,N_12927);
or U13030 (N_13030,N_12918,N_12801);
nor U13031 (N_13031,N_12884,N_12892);
xnor U13032 (N_13032,N_12954,N_12921);
xnor U13033 (N_13033,N_12903,N_12936);
or U13034 (N_13034,N_12856,N_12939);
or U13035 (N_13035,N_12937,N_12814);
xor U13036 (N_13036,N_12832,N_12802);
and U13037 (N_13037,N_12848,N_12817);
nor U13038 (N_13038,N_12894,N_12820);
nor U13039 (N_13039,N_12827,N_12876);
xnor U13040 (N_13040,N_12830,N_12845);
or U13041 (N_13041,N_12803,N_12912);
nor U13042 (N_13042,N_12814,N_12881);
nor U13043 (N_13043,N_12818,N_12906);
or U13044 (N_13044,N_12867,N_12892);
nor U13045 (N_13045,N_12801,N_12817);
and U13046 (N_13046,N_12905,N_12897);
nor U13047 (N_13047,N_12860,N_12819);
or U13048 (N_13048,N_12922,N_12857);
or U13049 (N_13049,N_12827,N_12953);
nor U13050 (N_13050,N_12881,N_12856);
nor U13051 (N_13051,N_12886,N_12939);
or U13052 (N_13052,N_12944,N_12809);
or U13053 (N_13053,N_12818,N_12879);
xnor U13054 (N_13054,N_12850,N_12896);
nor U13055 (N_13055,N_12877,N_12845);
or U13056 (N_13056,N_12935,N_12939);
and U13057 (N_13057,N_12848,N_12867);
xnor U13058 (N_13058,N_12954,N_12915);
xor U13059 (N_13059,N_12867,N_12943);
or U13060 (N_13060,N_12890,N_12857);
nor U13061 (N_13061,N_12937,N_12944);
nand U13062 (N_13062,N_12825,N_12871);
or U13063 (N_13063,N_12820,N_12844);
xor U13064 (N_13064,N_12830,N_12882);
and U13065 (N_13065,N_12936,N_12856);
nand U13066 (N_13066,N_12924,N_12830);
or U13067 (N_13067,N_12809,N_12911);
or U13068 (N_13068,N_12808,N_12918);
nand U13069 (N_13069,N_12824,N_12894);
nand U13070 (N_13070,N_12890,N_12900);
and U13071 (N_13071,N_12939,N_12914);
or U13072 (N_13072,N_12867,N_12940);
and U13073 (N_13073,N_12888,N_12819);
nor U13074 (N_13074,N_12883,N_12941);
xnor U13075 (N_13075,N_12925,N_12922);
nand U13076 (N_13076,N_12817,N_12878);
and U13077 (N_13077,N_12943,N_12881);
or U13078 (N_13078,N_12807,N_12841);
or U13079 (N_13079,N_12824,N_12896);
nand U13080 (N_13080,N_12894,N_12877);
nor U13081 (N_13081,N_12834,N_12888);
nor U13082 (N_13082,N_12883,N_12927);
nand U13083 (N_13083,N_12866,N_12887);
and U13084 (N_13084,N_12820,N_12904);
and U13085 (N_13085,N_12826,N_12836);
and U13086 (N_13086,N_12889,N_12936);
and U13087 (N_13087,N_12883,N_12867);
or U13088 (N_13088,N_12887,N_12855);
nand U13089 (N_13089,N_12912,N_12846);
nand U13090 (N_13090,N_12897,N_12941);
xnor U13091 (N_13091,N_12915,N_12834);
and U13092 (N_13092,N_12835,N_12864);
nand U13093 (N_13093,N_12900,N_12926);
xnor U13094 (N_13094,N_12861,N_12866);
and U13095 (N_13095,N_12851,N_12929);
xnor U13096 (N_13096,N_12889,N_12879);
xor U13097 (N_13097,N_12835,N_12927);
or U13098 (N_13098,N_12941,N_12893);
or U13099 (N_13099,N_12845,N_12904);
or U13100 (N_13100,N_12833,N_12904);
or U13101 (N_13101,N_12944,N_12948);
or U13102 (N_13102,N_12887,N_12910);
or U13103 (N_13103,N_12950,N_12955);
nand U13104 (N_13104,N_12931,N_12946);
nand U13105 (N_13105,N_12922,N_12935);
nor U13106 (N_13106,N_12840,N_12836);
and U13107 (N_13107,N_12885,N_12950);
or U13108 (N_13108,N_12927,N_12830);
nand U13109 (N_13109,N_12857,N_12859);
and U13110 (N_13110,N_12954,N_12883);
nand U13111 (N_13111,N_12813,N_12893);
nor U13112 (N_13112,N_12800,N_12835);
xnor U13113 (N_13113,N_12897,N_12846);
nor U13114 (N_13114,N_12895,N_12803);
nand U13115 (N_13115,N_12827,N_12845);
nor U13116 (N_13116,N_12815,N_12811);
or U13117 (N_13117,N_12838,N_12845);
nand U13118 (N_13118,N_12869,N_12802);
nor U13119 (N_13119,N_12955,N_12928);
or U13120 (N_13120,N_13065,N_13045);
and U13121 (N_13121,N_13096,N_13006);
nor U13122 (N_13122,N_13041,N_13026);
xor U13123 (N_13123,N_13049,N_13070);
and U13124 (N_13124,N_13037,N_13066);
and U13125 (N_13125,N_13111,N_13102);
xnor U13126 (N_13126,N_13044,N_13089);
or U13127 (N_13127,N_13003,N_13053);
nor U13128 (N_13128,N_13098,N_12978);
xnor U13129 (N_13129,N_12995,N_13091);
xor U13130 (N_13130,N_13072,N_13063);
nor U13131 (N_13131,N_12969,N_13109);
xnor U13132 (N_13132,N_13068,N_13051);
nand U13133 (N_13133,N_12990,N_13027);
and U13134 (N_13134,N_12992,N_13115);
nor U13135 (N_13135,N_13013,N_12973);
or U13136 (N_13136,N_13087,N_13085);
or U13137 (N_13137,N_13011,N_13009);
nor U13138 (N_13138,N_12998,N_12961);
xor U13139 (N_13139,N_12964,N_12962);
nand U13140 (N_13140,N_13080,N_13038);
nand U13141 (N_13141,N_13046,N_13022);
and U13142 (N_13142,N_13010,N_12960);
or U13143 (N_13143,N_13056,N_12983);
nor U13144 (N_13144,N_13028,N_12996);
nand U13145 (N_13145,N_13039,N_13054);
nor U13146 (N_13146,N_13029,N_12975);
or U13147 (N_13147,N_13103,N_12989);
nand U13148 (N_13148,N_12991,N_13024);
or U13149 (N_13149,N_13099,N_13075);
or U13150 (N_13150,N_13113,N_13033);
nand U13151 (N_13151,N_13016,N_13078);
xor U13152 (N_13152,N_13086,N_13018);
xor U13153 (N_13153,N_12993,N_13000);
or U13154 (N_13154,N_12976,N_13108);
xor U13155 (N_13155,N_12968,N_13032);
or U13156 (N_13156,N_13017,N_12986);
or U13157 (N_13157,N_13074,N_13110);
and U13158 (N_13158,N_13055,N_13047);
and U13159 (N_13159,N_13088,N_12965);
or U13160 (N_13160,N_13090,N_12984);
nor U13161 (N_13161,N_13036,N_12981);
xor U13162 (N_13162,N_12997,N_13077);
and U13163 (N_13163,N_12971,N_12979);
nor U13164 (N_13164,N_13048,N_13002);
nand U13165 (N_13165,N_13060,N_13105);
nand U13166 (N_13166,N_12985,N_13025);
or U13167 (N_13167,N_13107,N_13057);
or U13168 (N_13168,N_13004,N_13112);
nand U13169 (N_13169,N_13093,N_13020);
nand U13170 (N_13170,N_12967,N_13104);
and U13171 (N_13171,N_13034,N_12970);
nor U13172 (N_13172,N_13083,N_13015);
nor U13173 (N_13173,N_13079,N_13043);
or U13174 (N_13174,N_13094,N_12974);
nor U13175 (N_13175,N_13064,N_13067);
nor U13176 (N_13176,N_13073,N_13019);
and U13177 (N_13177,N_13101,N_13106);
or U13178 (N_13178,N_13040,N_13069);
nand U13179 (N_13179,N_13118,N_13001);
or U13180 (N_13180,N_13097,N_13076);
and U13181 (N_13181,N_13095,N_12972);
nand U13182 (N_13182,N_12966,N_12977);
xnor U13183 (N_13183,N_13082,N_13052);
and U13184 (N_13184,N_13062,N_13031);
nand U13185 (N_13185,N_13042,N_13030);
and U13186 (N_13186,N_12963,N_13021);
nand U13187 (N_13187,N_13012,N_12980);
nand U13188 (N_13188,N_13058,N_13050);
nand U13189 (N_13189,N_13084,N_13035);
xor U13190 (N_13190,N_13117,N_12988);
and U13191 (N_13191,N_12982,N_12994);
and U13192 (N_13192,N_13116,N_13119);
or U13193 (N_13193,N_13005,N_13100);
nand U13194 (N_13194,N_13059,N_13061);
and U13195 (N_13195,N_13007,N_12999);
and U13196 (N_13196,N_13014,N_13008);
nand U13197 (N_13197,N_13114,N_13071);
nand U13198 (N_13198,N_12987,N_13081);
and U13199 (N_13199,N_13092,N_13023);
and U13200 (N_13200,N_12972,N_13058);
or U13201 (N_13201,N_13027,N_13005);
and U13202 (N_13202,N_13015,N_13086);
and U13203 (N_13203,N_13013,N_12996);
xor U13204 (N_13204,N_12961,N_13110);
and U13205 (N_13205,N_13079,N_13001);
or U13206 (N_13206,N_13065,N_12990);
and U13207 (N_13207,N_13001,N_13069);
nand U13208 (N_13208,N_13015,N_13007);
nand U13209 (N_13209,N_13097,N_13020);
or U13210 (N_13210,N_12968,N_12982);
xor U13211 (N_13211,N_12985,N_12966);
nand U13212 (N_13212,N_13118,N_13024);
xnor U13213 (N_13213,N_13038,N_13024);
nand U13214 (N_13214,N_13064,N_12992);
or U13215 (N_13215,N_13116,N_12973);
nand U13216 (N_13216,N_12998,N_13119);
nand U13217 (N_13217,N_13113,N_12976);
nor U13218 (N_13218,N_13008,N_13059);
nor U13219 (N_13219,N_13078,N_13099);
xnor U13220 (N_13220,N_12973,N_13081);
xnor U13221 (N_13221,N_12998,N_13099);
xor U13222 (N_13222,N_13106,N_13107);
or U13223 (N_13223,N_13015,N_13023);
xnor U13224 (N_13224,N_13010,N_13016);
or U13225 (N_13225,N_13086,N_13016);
nand U13226 (N_13226,N_13042,N_13060);
xor U13227 (N_13227,N_13048,N_12982);
or U13228 (N_13228,N_13034,N_13094);
xor U13229 (N_13229,N_12975,N_13086);
or U13230 (N_13230,N_12967,N_13008);
nand U13231 (N_13231,N_13001,N_13078);
or U13232 (N_13232,N_12999,N_13063);
and U13233 (N_13233,N_12961,N_13012);
nor U13234 (N_13234,N_12973,N_13034);
nor U13235 (N_13235,N_13079,N_13004);
or U13236 (N_13236,N_13027,N_12963);
nor U13237 (N_13237,N_13019,N_13119);
xnor U13238 (N_13238,N_13064,N_12965);
or U13239 (N_13239,N_13026,N_12963);
and U13240 (N_13240,N_13027,N_13015);
xor U13241 (N_13241,N_12961,N_13117);
and U13242 (N_13242,N_13012,N_13077);
or U13243 (N_13243,N_12983,N_13055);
nor U13244 (N_13244,N_13010,N_13085);
nand U13245 (N_13245,N_13071,N_13102);
xnor U13246 (N_13246,N_13032,N_13100);
nand U13247 (N_13247,N_13113,N_13021);
and U13248 (N_13248,N_13044,N_13112);
nor U13249 (N_13249,N_13032,N_13052);
nor U13250 (N_13250,N_12973,N_13072);
nand U13251 (N_13251,N_13000,N_13004);
nand U13252 (N_13252,N_13019,N_13000);
nor U13253 (N_13253,N_13102,N_13046);
nor U13254 (N_13254,N_13072,N_13047);
or U13255 (N_13255,N_12966,N_13086);
xnor U13256 (N_13256,N_12998,N_13051);
xnor U13257 (N_13257,N_13025,N_13056);
or U13258 (N_13258,N_13005,N_12962);
xnor U13259 (N_13259,N_13070,N_12975);
xnor U13260 (N_13260,N_13031,N_13028);
or U13261 (N_13261,N_13110,N_13017);
xor U13262 (N_13262,N_13038,N_12972);
nand U13263 (N_13263,N_13058,N_12983);
xnor U13264 (N_13264,N_13093,N_12980);
or U13265 (N_13265,N_13004,N_13114);
xor U13266 (N_13266,N_13071,N_13117);
nor U13267 (N_13267,N_13088,N_13067);
and U13268 (N_13268,N_13062,N_13109);
nor U13269 (N_13269,N_13114,N_13080);
nand U13270 (N_13270,N_13086,N_13059);
or U13271 (N_13271,N_13092,N_13063);
xor U13272 (N_13272,N_13069,N_13068);
and U13273 (N_13273,N_13036,N_12997);
or U13274 (N_13274,N_12971,N_13075);
nor U13275 (N_13275,N_13119,N_13034);
xnor U13276 (N_13276,N_12980,N_13008);
nand U13277 (N_13277,N_13114,N_13025);
and U13278 (N_13278,N_12990,N_12993);
nor U13279 (N_13279,N_13055,N_13054);
and U13280 (N_13280,N_13236,N_13141);
or U13281 (N_13281,N_13183,N_13163);
nor U13282 (N_13282,N_13182,N_13208);
or U13283 (N_13283,N_13266,N_13229);
nand U13284 (N_13284,N_13170,N_13224);
or U13285 (N_13285,N_13256,N_13197);
xor U13286 (N_13286,N_13193,N_13184);
or U13287 (N_13287,N_13215,N_13262);
and U13288 (N_13288,N_13278,N_13202);
nand U13289 (N_13289,N_13130,N_13121);
or U13290 (N_13290,N_13210,N_13261);
and U13291 (N_13291,N_13188,N_13156);
or U13292 (N_13292,N_13192,N_13240);
and U13293 (N_13293,N_13169,N_13178);
nor U13294 (N_13294,N_13167,N_13244);
and U13295 (N_13295,N_13195,N_13271);
nand U13296 (N_13296,N_13151,N_13238);
xor U13297 (N_13297,N_13270,N_13205);
xnor U13298 (N_13298,N_13253,N_13129);
xor U13299 (N_13299,N_13218,N_13172);
and U13300 (N_13300,N_13127,N_13199);
nor U13301 (N_13301,N_13264,N_13131);
xnor U13302 (N_13302,N_13123,N_13175);
and U13303 (N_13303,N_13198,N_13171);
xnor U13304 (N_13304,N_13275,N_13150);
nand U13305 (N_13305,N_13137,N_13248);
or U13306 (N_13306,N_13279,N_13157);
nand U13307 (N_13307,N_13273,N_13138);
nor U13308 (N_13308,N_13155,N_13126);
nor U13309 (N_13309,N_13128,N_13153);
or U13310 (N_13310,N_13154,N_13159);
nand U13311 (N_13311,N_13144,N_13190);
or U13312 (N_13312,N_13263,N_13135);
xnor U13313 (N_13313,N_13237,N_13226);
nor U13314 (N_13314,N_13223,N_13255);
nor U13315 (N_13315,N_13276,N_13189);
or U13316 (N_13316,N_13214,N_13158);
nand U13317 (N_13317,N_13232,N_13125);
xnor U13318 (N_13318,N_13139,N_13147);
xnor U13319 (N_13319,N_13246,N_13257);
and U13320 (N_13320,N_13134,N_13140);
xor U13321 (N_13321,N_13164,N_13249);
and U13322 (N_13322,N_13222,N_13259);
nand U13323 (N_13323,N_13200,N_13185);
or U13324 (N_13324,N_13212,N_13133);
and U13325 (N_13325,N_13149,N_13250);
nor U13326 (N_13326,N_13203,N_13165);
or U13327 (N_13327,N_13194,N_13234);
and U13328 (N_13328,N_13220,N_13277);
and U13329 (N_13329,N_13254,N_13181);
xnor U13330 (N_13330,N_13211,N_13148);
xor U13331 (N_13331,N_13132,N_13225);
nor U13332 (N_13332,N_13120,N_13274);
or U13333 (N_13333,N_13176,N_13122);
nand U13334 (N_13334,N_13145,N_13173);
xor U13335 (N_13335,N_13146,N_13213);
or U13336 (N_13336,N_13217,N_13231);
nor U13337 (N_13337,N_13265,N_13228);
or U13338 (N_13338,N_13216,N_13239);
nor U13339 (N_13339,N_13168,N_13221);
nor U13340 (N_13340,N_13242,N_13245);
xor U13341 (N_13341,N_13243,N_13179);
xnor U13342 (N_13342,N_13207,N_13142);
nor U13343 (N_13343,N_13136,N_13227);
and U13344 (N_13344,N_13267,N_13219);
and U13345 (N_13345,N_13233,N_13209);
and U13346 (N_13346,N_13201,N_13152);
nor U13347 (N_13347,N_13196,N_13166);
or U13348 (N_13348,N_13162,N_13241);
and U13349 (N_13349,N_13230,N_13186);
or U13350 (N_13350,N_13272,N_13174);
xor U13351 (N_13351,N_13187,N_13269);
or U13352 (N_13352,N_13252,N_13161);
nor U13353 (N_13353,N_13124,N_13160);
nand U13354 (N_13354,N_13268,N_13206);
or U13355 (N_13355,N_13191,N_13235);
or U13356 (N_13356,N_13260,N_13258);
xor U13357 (N_13357,N_13247,N_13180);
or U13358 (N_13358,N_13251,N_13143);
xor U13359 (N_13359,N_13177,N_13204);
xnor U13360 (N_13360,N_13267,N_13228);
and U13361 (N_13361,N_13125,N_13215);
nor U13362 (N_13362,N_13146,N_13140);
and U13363 (N_13363,N_13272,N_13223);
nand U13364 (N_13364,N_13123,N_13124);
nand U13365 (N_13365,N_13198,N_13131);
nor U13366 (N_13366,N_13150,N_13175);
nor U13367 (N_13367,N_13138,N_13133);
or U13368 (N_13368,N_13165,N_13215);
xor U13369 (N_13369,N_13276,N_13279);
or U13370 (N_13370,N_13190,N_13250);
nand U13371 (N_13371,N_13163,N_13193);
xnor U13372 (N_13372,N_13141,N_13245);
xor U13373 (N_13373,N_13172,N_13143);
and U13374 (N_13374,N_13189,N_13245);
xnor U13375 (N_13375,N_13248,N_13224);
nor U13376 (N_13376,N_13263,N_13152);
xor U13377 (N_13377,N_13142,N_13169);
or U13378 (N_13378,N_13244,N_13251);
xor U13379 (N_13379,N_13213,N_13271);
xnor U13380 (N_13380,N_13255,N_13274);
and U13381 (N_13381,N_13132,N_13216);
xnor U13382 (N_13382,N_13136,N_13217);
nand U13383 (N_13383,N_13261,N_13154);
xnor U13384 (N_13384,N_13186,N_13270);
or U13385 (N_13385,N_13248,N_13221);
xor U13386 (N_13386,N_13279,N_13171);
nor U13387 (N_13387,N_13268,N_13174);
and U13388 (N_13388,N_13192,N_13173);
nor U13389 (N_13389,N_13227,N_13185);
xnor U13390 (N_13390,N_13148,N_13123);
nor U13391 (N_13391,N_13157,N_13278);
nor U13392 (N_13392,N_13172,N_13127);
nor U13393 (N_13393,N_13206,N_13227);
and U13394 (N_13394,N_13270,N_13138);
or U13395 (N_13395,N_13215,N_13171);
nor U13396 (N_13396,N_13126,N_13241);
nor U13397 (N_13397,N_13197,N_13233);
nand U13398 (N_13398,N_13130,N_13267);
xnor U13399 (N_13399,N_13183,N_13199);
nor U13400 (N_13400,N_13180,N_13233);
and U13401 (N_13401,N_13191,N_13271);
or U13402 (N_13402,N_13164,N_13126);
xnor U13403 (N_13403,N_13160,N_13197);
and U13404 (N_13404,N_13244,N_13241);
nand U13405 (N_13405,N_13222,N_13141);
nor U13406 (N_13406,N_13176,N_13185);
or U13407 (N_13407,N_13219,N_13275);
xor U13408 (N_13408,N_13126,N_13231);
nor U13409 (N_13409,N_13153,N_13266);
nor U13410 (N_13410,N_13121,N_13202);
or U13411 (N_13411,N_13216,N_13149);
nor U13412 (N_13412,N_13278,N_13124);
and U13413 (N_13413,N_13122,N_13251);
xor U13414 (N_13414,N_13223,N_13165);
xor U13415 (N_13415,N_13173,N_13149);
xnor U13416 (N_13416,N_13169,N_13272);
nand U13417 (N_13417,N_13239,N_13177);
nand U13418 (N_13418,N_13163,N_13129);
nand U13419 (N_13419,N_13154,N_13242);
nand U13420 (N_13420,N_13124,N_13165);
and U13421 (N_13421,N_13186,N_13202);
nand U13422 (N_13422,N_13154,N_13246);
or U13423 (N_13423,N_13176,N_13212);
and U13424 (N_13424,N_13181,N_13207);
and U13425 (N_13425,N_13268,N_13234);
nor U13426 (N_13426,N_13222,N_13139);
or U13427 (N_13427,N_13196,N_13155);
xor U13428 (N_13428,N_13252,N_13251);
xor U13429 (N_13429,N_13140,N_13198);
and U13430 (N_13430,N_13146,N_13184);
xor U13431 (N_13431,N_13168,N_13140);
nand U13432 (N_13432,N_13275,N_13178);
xor U13433 (N_13433,N_13155,N_13143);
and U13434 (N_13434,N_13173,N_13195);
nand U13435 (N_13435,N_13167,N_13250);
nand U13436 (N_13436,N_13165,N_13211);
nor U13437 (N_13437,N_13124,N_13168);
or U13438 (N_13438,N_13152,N_13120);
or U13439 (N_13439,N_13274,N_13173);
or U13440 (N_13440,N_13432,N_13392);
and U13441 (N_13441,N_13343,N_13342);
nand U13442 (N_13442,N_13345,N_13302);
xor U13443 (N_13443,N_13414,N_13306);
or U13444 (N_13444,N_13395,N_13322);
nand U13445 (N_13445,N_13337,N_13326);
nor U13446 (N_13446,N_13379,N_13391);
nand U13447 (N_13447,N_13358,N_13344);
xnor U13448 (N_13448,N_13433,N_13355);
nor U13449 (N_13449,N_13297,N_13425);
xnor U13450 (N_13450,N_13353,N_13310);
and U13451 (N_13451,N_13399,N_13439);
or U13452 (N_13452,N_13316,N_13348);
xnor U13453 (N_13453,N_13361,N_13331);
nor U13454 (N_13454,N_13285,N_13401);
or U13455 (N_13455,N_13350,N_13370);
nand U13456 (N_13456,N_13312,N_13282);
or U13457 (N_13457,N_13327,N_13308);
nor U13458 (N_13458,N_13287,N_13405);
nand U13459 (N_13459,N_13368,N_13434);
and U13460 (N_13460,N_13280,N_13315);
nor U13461 (N_13461,N_13388,N_13318);
xnor U13462 (N_13462,N_13303,N_13387);
nor U13463 (N_13463,N_13437,N_13410);
nand U13464 (N_13464,N_13288,N_13411);
nor U13465 (N_13465,N_13325,N_13313);
nor U13466 (N_13466,N_13417,N_13426);
and U13467 (N_13467,N_13329,N_13321);
and U13468 (N_13468,N_13336,N_13385);
nor U13469 (N_13469,N_13334,N_13371);
and U13470 (N_13470,N_13422,N_13362);
nand U13471 (N_13471,N_13409,N_13380);
nand U13472 (N_13472,N_13406,N_13438);
nor U13473 (N_13473,N_13291,N_13413);
or U13474 (N_13474,N_13320,N_13430);
or U13475 (N_13475,N_13375,N_13396);
and U13476 (N_13476,N_13415,N_13349);
or U13477 (N_13477,N_13397,N_13364);
or U13478 (N_13478,N_13419,N_13404);
nor U13479 (N_13479,N_13289,N_13347);
or U13480 (N_13480,N_13298,N_13283);
or U13481 (N_13481,N_13319,N_13338);
and U13482 (N_13482,N_13309,N_13435);
nand U13483 (N_13483,N_13335,N_13311);
xnor U13484 (N_13484,N_13324,N_13393);
and U13485 (N_13485,N_13427,N_13389);
and U13486 (N_13486,N_13294,N_13300);
nor U13487 (N_13487,N_13293,N_13317);
nand U13488 (N_13488,N_13418,N_13307);
or U13489 (N_13489,N_13363,N_13412);
and U13490 (N_13490,N_13305,N_13424);
nor U13491 (N_13491,N_13359,N_13402);
and U13492 (N_13492,N_13394,N_13386);
nor U13493 (N_13493,N_13400,N_13367);
or U13494 (N_13494,N_13423,N_13374);
and U13495 (N_13495,N_13352,N_13296);
xnor U13496 (N_13496,N_13384,N_13346);
or U13497 (N_13497,N_13378,N_13286);
and U13498 (N_13498,N_13301,N_13377);
nor U13499 (N_13499,N_13281,N_13383);
and U13500 (N_13500,N_13284,N_13354);
nand U13501 (N_13501,N_13421,N_13431);
xor U13502 (N_13502,N_13408,N_13323);
or U13503 (N_13503,N_13429,N_13420);
nor U13504 (N_13504,N_13381,N_13372);
nor U13505 (N_13505,N_13290,N_13360);
or U13506 (N_13506,N_13376,N_13332);
and U13507 (N_13507,N_13304,N_13390);
xor U13508 (N_13508,N_13341,N_13356);
and U13509 (N_13509,N_13366,N_13340);
nor U13510 (N_13510,N_13333,N_13428);
xor U13511 (N_13511,N_13357,N_13365);
xnor U13512 (N_13512,N_13314,N_13328);
or U13513 (N_13513,N_13416,N_13339);
nand U13514 (N_13514,N_13299,N_13398);
and U13515 (N_13515,N_13295,N_13373);
and U13516 (N_13516,N_13436,N_13351);
or U13517 (N_13517,N_13292,N_13403);
xnor U13518 (N_13518,N_13330,N_13382);
xor U13519 (N_13519,N_13369,N_13407);
nor U13520 (N_13520,N_13403,N_13422);
or U13521 (N_13521,N_13293,N_13395);
xor U13522 (N_13522,N_13285,N_13284);
xnor U13523 (N_13523,N_13414,N_13425);
xnor U13524 (N_13524,N_13377,N_13403);
nor U13525 (N_13525,N_13355,N_13343);
xor U13526 (N_13526,N_13352,N_13288);
nand U13527 (N_13527,N_13333,N_13418);
and U13528 (N_13528,N_13393,N_13305);
nand U13529 (N_13529,N_13384,N_13398);
nand U13530 (N_13530,N_13324,N_13402);
nor U13531 (N_13531,N_13390,N_13310);
nor U13532 (N_13532,N_13419,N_13425);
or U13533 (N_13533,N_13400,N_13397);
nand U13534 (N_13534,N_13400,N_13322);
and U13535 (N_13535,N_13401,N_13352);
nor U13536 (N_13536,N_13364,N_13413);
xnor U13537 (N_13537,N_13414,N_13314);
and U13538 (N_13538,N_13367,N_13299);
nor U13539 (N_13539,N_13362,N_13349);
or U13540 (N_13540,N_13339,N_13329);
nand U13541 (N_13541,N_13330,N_13331);
and U13542 (N_13542,N_13333,N_13302);
and U13543 (N_13543,N_13284,N_13412);
nand U13544 (N_13544,N_13424,N_13354);
nor U13545 (N_13545,N_13432,N_13435);
nand U13546 (N_13546,N_13418,N_13326);
or U13547 (N_13547,N_13407,N_13311);
nand U13548 (N_13548,N_13371,N_13308);
nor U13549 (N_13549,N_13293,N_13287);
and U13550 (N_13550,N_13353,N_13311);
nor U13551 (N_13551,N_13322,N_13392);
or U13552 (N_13552,N_13282,N_13342);
or U13553 (N_13553,N_13286,N_13327);
nand U13554 (N_13554,N_13316,N_13411);
nand U13555 (N_13555,N_13406,N_13384);
and U13556 (N_13556,N_13303,N_13339);
xnor U13557 (N_13557,N_13342,N_13405);
or U13558 (N_13558,N_13295,N_13288);
or U13559 (N_13559,N_13351,N_13377);
xnor U13560 (N_13560,N_13360,N_13361);
nor U13561 (N_13561,N_13339,N_13407);
nor U13562 (N_13562,N_13318,N_13376);
xor U13563 (N_13563,N_13338,N_13406);
and U13564 (N_13564,N_13400,N_13340);
and U13565 (N_13565,N_13380,N_13346);
nor U13566 (N_13566,N_13401,N_13299);
nand U13567 (N_13567,N_13304,N_13404);
nor U13568 (N_13568,N_13395,N_13390);
and U13569 (N_13569,N_13291,N_13429);
and U13570 (N_13570,N_13374,N_13307);
xor U13571 (N_13571,N_13413,N_13420);
and U13572 (N_13572,N_13318,N_13363);
and U13573 (N_13573,N_13379,N_13438);
nand U13574 (N_13574,N_13320,N_13344);
and U13575 (N_13575,N_13358,N_13312);
or U13576 (N_13576,N_13438,N_13335);
nand U13577 (N_13577,N_13360,N_13355);
nor U13578 (N_13578,N_13284,N_13333);
and U13579 (N_13579,N_13373,N_13302);
xor U13580 (N_13580,N_13316,N_13327);
nor U13581 (N_13581,N_13393,N_13426);
and U13582 (N_13582,N_13364,N_13297);
and U13583 (N_13583,N_13379,N_13408);
and U13584 (N_13584,N_13296,N_13373);
nor U13585 (N_13585,N_13283,N_13309);
xnor U13586 (N_13586,N_13392,N_13337);
nand U13587 (N_13587,N_13336,N_13298);
nor U13588 (N_13588,N_13344,N_13395);
xnor U13589 (N_13589,N_13425,N_13309);
and U13590 (N_13590,N_13300,N_13411);
xor U13591 (N_13591,N_13311,N_13422);
nand U13592 (N_13592,N_13297,N_13404);
or U13593 (N_13593,N_13435,N_13293);
xnor U13594 (N_13594,N_13404,N_13317);
nor U13595 (N_13595,N_13434,N_13341);
xor U13596 (N_13596,N_13362,N_13352);
and U13597 (N_13597,N_13381,N_13390);
xor U13598 (N_13598,N_13333,N_13385);
and U13599 (N_13599,N_13309,N_13411);
xor U13600 (N_13600,N_13469,N_13464);
nand U13601 (N_13601,N_13487,N_13486);
nor U13602 (N_13602,N_13468,N_13506);
or U13603 (N_13603,N_13503,N_13534);
nor U13604 (N_13604,N_13521,N_13483);
or U13605 (N_13605,N_13575,N_13548);
and U13606 (N_13606,N_13470,N_13457);
or U13607 (N_13607,N_13584,N_13553);
xnor U13608 (N_13608,N_13450,N_13565);
nand U13609 (N_13609,N_13582,N_13489);
nand U13610 (N_13610,N_13474,N_13459);
xor U13611 (N_13611,N_13569,N_13528);
xnor U13612 (N_13612,N_13526,N_13531);
and U13613 (N_13613,N_13445,N_13590);
or U13614 (N_13614,N_13588,N_13440);
nand U13615 (N_13615,N_13578,N_13515);
nand U13616 (N_13616,N_13564,N_13544);
nand U13617 (N_13617,N_13596,N_13480);
nand U13618 (N_13618,N_13586,N_13523);
and U13619 (N_13619,N_13524,N_13455);
xnor U13620 (N_13620,N_13460,N_13516);
xor U13621 (N_13621,N_13494,N_13540);
xor U13622 (N_13622,N_13536,N_13545);
or U13623 (N_13623,N_13583,N_13441);
and U13624 (N_13624,N_13504,N_13466);
xor U13625 (N_13625,N_13488,N_13543);
or U13626 (N_13626,N_13579,N_13567);
and U13627 (N_13627,N_13448,N_13566);
nor U13628 (N_13628,N_13563,N_13500);
nor U13629 (N_13629,N_13472,N_13454);
xnor U13630 (N_13630,N_13491,N_13555);
nand U13631 (N_13631,N_13539,N_13571);
or U13632 (N_13632,N_13541,N_13546);
or U13633 (N_13633,N_13573,N_13576);
or U13634 (N_13634,N_13598,N_13501);
and U13635 (N_13635,N_13499,N_13572);
nor U13636 (N_13636,N_13556,N_13453);
xnor U13637 (N_13637,N_13510,N_13481);
nand U13638 (N_13638,N_13496,N_13595);
or U13639 (N_13639,N_13599,N_13530);
xor U13640 (N_13640,N_13533,N_13444);
and U13641 (N_13641,N_13513,N_13478);
or U13642 (N_13642,N_13592,N_13547);
and U13643 (N_13643,N_13574,N_13559);
xnor U13644 (N_13644,N_13527,N_13519);
or U13645 (N_13645,N_13502,N_13493);
nand U13646 (N_13646,N_13554,N_13458);
nand U13647 (N_13647,N_13456,N_13497);
and U13648 (N_13648,N_13463,N_13475);
and U13649 (N_13649,N_13577,N_13560);
nor U13650 (N_13650,N_13482,N_13462);
nand U13651 (N_13651,N_13511,N_13550);
or U13652 (N_13652,N_13446,N_13551);
xor U13653 (N_13653,N_13538,N_13557);
nor U13654 (N_13654,N_13594,N_13517);
or U13655 (N_13655,N_13490,N_13520);
xor U13656 (N_13656,N_13597,N_13509);
xor U13657 (N_13657,N_13442,N_13508);
or U13658 (N_13658,N_13495,N_13535);
or U13659 (N_13659,N_13537,N_13505);
or U13660 (N_13660,N_13473,N_13461);
nor U13661 (N_13661,N_13587,N_13518);
xor U13662 (N_13662,N_13507,N_13585);
and U13663 (N_13663,N_13465,N_13591);
xor U13664 (N_13664,N_13525,N_13581);
nor U13665 (N_13665,N_13561,N_13447);
or U13666 (N_13666,N_13485,N_13522);
and U13667 (N_13667,N_13529,N_13542);
and U13668 (N_13668,N_13467,N_13549);
nand U13669 (N_13669,N_13471,N_13568);
nand U13670 (N_13670,N_13580,N_13532);
and U13671 (N_13671,N_13451,N_13492);
and U13672 (N_13672,N_13570,N_13593);
and U13673 (N_13673,N_13562,N_13477);
nor U13674 (N_13674,N_13589,N_13479);
xor U13675 (N_13675,N_13452,N_13514);
nand U13676 (N_13676,N_13443,N_13512);
nor U13677 (N_13677,N_13498,N_13449);
nand U13678 (N_13678,N_13476,N_13484);
nand U13679 (N_13679,N_13558,N_13552);
or U13680 (N_13680,N_13571,N_13460);
or U13681 (N_13681,N_13465,N_13559);
nand U13682 (N_13682,N_13581,N_13562);
nand U13683 (N_13683,N_13440,N_13452);
and U13684 (N_13684,N_13507,N_13539);
or U13685 (N_13685,N_13578,N_13522);
nand U13686 (N_13686,N_13489,N_13580);
or U13687 (N_13687,N_13531,N_13516);
nand U13688 (N_13688,N_13470,N_13585);
and U13689 (N_13689,N_13444,N_13595);
nor U13690 (N_13690,N_13519,N_13518);
nor U13691 (N_13691,N_13496,N_13480);
or U13692 (N_13692,N_13521,N_13496);
or U13693 (N_13693,N_13569,N_13591);
and U13694 (N_13694,N_13478,N_13588);
and U13695 (N_13695,N_13572,N_13598);
nor U13696 (N_13696,N_13481,N_13593);
or U13697 (N_13697,N_13598,N_13573);
xnor U13698 (N_13698,N_13504,N_13507);
nor U13699 (N_13699,N_13486,N_13523);
or U13700 (N_13700,N_13468,N_13589);
xnor U13701 (N_13701,N_13507,N_13457);
xnor U13702 (N_13702,N_13504,N_13520);
and U13703 (N_13703,N_13510,N_13508);
nor U13704 (N_13704,N_13454,N_13474);
nor U13705 (N_13705,N_13476,N_13589);
nand U13706 (N_13706,N_13484,N_13490);
and U13707 (N_13707,N_13516,N_13538);
nor U13708 (N_13708,N_13514,N_13459);
nor U13709 (N_13709,N_13528,N_13564);
nor U13710 (N_13710,N_13521,N_13536);
xor U13711 (N_13711,N_13522,N_13456);
and U13712 (N_13712,N_13545,N_13583);
and U13713 (N_13713,N_13568,N_13590);
xor U13714 (N_13714,N_13539,N_13546);
or U13715 (N_13715,N_13526,N_13441);
and U13716 (N_13716,N_13459,N_13527);
xor U13717 (N_13717,N_13583,N_13536);
or U13718 (N_13718,N_13455,N_13507);
or U13719 (N_13719,N_13556,N_13450);
or U13720 (N_13720,N_13498,N_13460);
xor U13721 (N_13721,N_13593,N_13580);
and U13722 (N_13722,N_13474,N_13526);
or U13723 (N_13723,N_13492,N_13488);
and U13724 (N_13724,N_13558,N_13518);
nand U13725 (N_13725,N_13552,N_13586);
and U13726 (N_13726,N_13514,N_13482);
and U13727 (N_13727,N_13551,N_13466);
nor U13728 (N_13728,N_13487,N_13496);
nand U13729 (N_13729,N_13598,N_13512);
nand U13730 (N_13730,N_13588,N_13474);
nor U13731 (N_13731,N_13447,N_13504);
and U13732 (N_13732,N_13519,N_13575);
or U13733 (N_13733,N_13585,N_13548);
nand U13734 (N_13734,N_13488,N_13559);
or U13735 (N_13735,N_13478,N_13482);
nand U13736 (N_13736,N_13584,N_13594);
and U13737 (N_13737,N_13534,N_13483);
and U13738 (N_13738,N_13509,N_13457);
xnor U13739 (N_13739,N_13488,N_13448);
nor U13740 (N_13740,N_13567,N_13532);
xnor U13741 (N_13741,N_13493,N_13531);
and U13742 (N_13742,N_13468,N_13526);
and U13743 (N_13743,N_13564,N_13443);
or U13744 (N_13744,N_13588,N_13591);
nor U13745 (N_13745,N_13494,N_13566);
nor U13746 (N_13746,N_13574,N_13458);
xor U13747 (N_13747,N_13560,N_13573);
and U13748 (N_13748,N_13478,N_13498);
nor U13749 (N_13749,N_13511,N_13573);
or U13750 (N_13750,N_13595,N_13516);
nor U13751 (N_13751,N_13455,N_13596);
xnor U13752 (N_13752,N_13497,N_13563);
or U13753 (N_13753,N_13504,N_13572);
xor U13754 (N_13754,N_13539,N_13552);
xnor U13755 (N_13755,N_13578,N_13597);
nand U13756 (N_13756,N_13517,N_13468);
or U13757 (N_13757,N_13562,N_13507);
nand U13758 (N_13758,N_13450,N_13588);
and U13759 (N_13759,N_13549,N_13456);
nor U13760 (N_13760,N_13626,N_13620);
or U13761 (N_13761,N_13630,N_13696);
and U13762 (N_13762,N_13737,N_13748);
nand U13763 (N_13763,N_13729,N_13745);
and U13764 (N_13764,N_13719,N_13621);
nand U13765 (N_13765,N_13694,N_13676);
nor U13766 (N_13766,N_13644,N_13603);
nor U13767 (N_13767,N_13718,N_13608);
nor U13768 (N_13768,N_13675,N_13628);
or U13769 (N_13769,N_13688,N_13659);
and U13770 (N_13770,N_13652,N_13663);
and U13771 (N_13771,N_13604,N_13758);
nor U13772 (N_13772,N_13636,N_13703);
xor U13773 (N_13773,N_13672,N_13616);
or U13774 (N_13774,N_13623,N_13751);
nand U13775 (N_13775,N_13666,N_13647);
and U13776 (N_13776,N_13726,N_13645);
xnor U13777 (N_13777,N_13640,N_13697);
and U13778 (N_13778,N_13690,N_13759);
and U13779 (N_13779,N_13691,N_13658);
nand U13780 (N_13780,N_13612,N_13730);
nor U13781 (N_13781,N_13749,N_13709);
xor U13782 (N_13782,N_13735,N_13699);
and U13783 (N_13783,N_13680,N_13665);
xnor U13784 (N_13784,N_13629,N_13664);
nand U13785 (N_13785,N_13633,N_13738);
xnor U13786 (N_13786,N_13601,N_13639);
nand U13787 (N_13787,N_13660,N_13602);
or U13788 (N_13788,N_13727,N_13682);
xnor U13789 (N_13789,N_13624,N_13674);
nand U13790 (N_13790,N_13646,N_13705);
xor U13791 (N_13791,N_13704,N_13625);
or U13792 (N_13792,N_13609,N_13707);
nand U13793 (N_13793,N_13638,N_13673);
xor U13794 (N_13794,N_13728,N_13741);
xor U13795 (N_13795,N_13753,N_13740);
and U13796 (N_13796,N_13611,N_13610);
xor U13797 (N_13797,N_13634,N_13668);
xnor U13798 (N_13798,N_13618,N_13736);
nor U13799 (N_13799,N_13606,N_13747);
nand U13800 (N_13800,N_13733,N_13642);
xnor U13801 (N_13801,N_13641,N_13649);
xor U13802 (N_13802,N_13643,N_13706);
xor U13803 (N_13803,N_13677,N_13756);
nand U13804 (N_13804,N_13686,N_13600);
xnor U13805 (N_13805,N_13631,N_13708);
nor U13806 (N_13806,N_13622,N_13655);
xnor U13807 (N_13807,N_13710,N_13698);
nand U13808 (N_13808,N_13742,N_13679);
xnor U13809 (N_13809,N_13656,N_13700);
or U13810 (N_13810,N_13605,N_13750);
and U13811 (N_13811,N_13637,N_13725);
xor U13812 (N_13812,N_13746,N_13661);
xor U13813 (N_13813,N_13662,N_13731);
nand U13814 (N_13814,N_13678,N_13693);
xor U13815 (N_13815,N_13754,N_13739);
and U13816 (N_13816,N_13714,N_13716);
or U13817 (N_13817,N_13724,N_13687);
nand U13818 (N_13818,N_13615,N_13717);
nor U13819 (N_13819,N_13648,N_13752);
xor U13820 (N_13820,N_13721,N_13734);
nand U13821 (N_13821,N_13617,N_13713);
xnor U13822 (N_13822,N_13720,N_13689);
nor U13823 (N_13823,N_13712,N_13743);
nand U13824 (N_13824,N_13723,N_13681);
nand U13825 (N_13825,N_13684,N_13627);
nor U13826 (N_13826,N_13650,N_13692);
or U13827 (N_13827,N_13755,N_13669);
or U13828 (N_13828,N_13632,N_13701);
nand U13829 (N_13829,N_13651,N_13757);
nor U13830 (N_13830,N_13613,N_13695);
nor U13831 (N_13831,N_13715,N_13667);
and U13832 (N_13832,N_13670,N_13732);
and U13833 (N_13833,N_13635,N_13702);
nand U13834 (N_13834,N_13614,N_13607);
and U13835 (N_13835,N_13657,N_13653);
and U13836 (N_13836,N_13654,N_13711);
or U13837 (N_13837,N_13722,N_13671);
or U13838 (N_13838,N_13683,N_13685);
xnor U13839 (N_13839,N_13744,N_13619);
xor U13840 (N_13840,N_13625,N_13729);
nor U13841 (N_13841,N_13690,N_13617);
xnor U13842 (N_13842,N_13703,N_13681);
nand U13843 (N_13843,N_13617,N_13641);
or U13844 (N_13844,N_13624,N_13656);
and U13845 (N_13845,N_13678,N_13676);
nor U13846 (N_13846,N_13661,N_13718);
xnor U13847 (N_13847,N_13658,N_13618);
nor U13848 (N_13848,N_13716,N_13704);
and U13849 (N_13849,N_13648,N_13687);
nand U13850 (N_13850,N_13734,N_13718);
nand U13851 (N_13851,N_13608,N_13754);
nand U13852 (N_13852,N_13750,N_13717);
or U13853 (N_13853,N_13715,N_13707);
nand U13854 (N_13854,N_13732,N_13611);
and U13855 (N_13855,N_13676,N_13747);
nand U13856 (N_13856,N_13744,N_13713);
nor U13857 (N_13857,N_13693,N_13708);
xor U13858 (N_13858,N_13605,N_13618);
xor U13859 (N_13859,N_13718,N_13634);
xnor U13860 (N_13860,N_13686,N_13745);
nor U13861 (N_13861,N_13679,N_13653);
xor U13862 (N_13862,N_13660,N_13719);
or U13863 (N_13863,N_13653,N_13728);
nor U13864 (N_13864,N_13621,N_13631);
nor U13865 (N_13865,N_13705,N_13637);
nand U13866 (N_13866,N_13648,N_13716);
xnor U13867 (N_13867,N_13683,N_13643);
xor U13868 (N_13868,N_13610,N_13658);
nor U13869 (N_13869,N_13701,N_13626);
nand U13870 (N_13870,N_13657,N_13739);
xnor U13871 (N_13871,N_13655,N_13752);
xor U13872 (N_13872,N_13759,N_13661);
xor U13873 (N_13873,N_13666,N_13706);
nand U13874 (N_13874,N_13611,N_13671);
or U13875 (N_13875,N_13629,N_13665);
xnor U13876 (N_13876,N_13714,N_13635);
and U13877 (N_13877,N_13708,N_13698);
and U13878 (N_13878,N_13704,N_13745);
xor U13879 (N_13879,N_13607,N_13709);
or U13880 (N_13880,N_13724,N_13696);
and U13881 (N_13881,N_13706,N_13608);
nor U13882 (N_13882,N_13754,N_13678);
nand U13883 (N_13883,N_13711,N_13698);
nand U13884 (N_13884,N_13635,N_13724);
nor U13885 (N_13885,N_13639,N_13742);
nand U13886 (N_13886,N_13734,N_13654);
nor U13887 (N_13887,N_13624,N_13744);
xnor U13888 (N_13888,N_13641,N_13690);
xor U13889 (N_13889,N_13755,N_13690);
nand U13890 (N_13890,N_13676,N_13748);
nor U13891 (N_13891,N_13750,N_13611);
or U13892 (N_13892,N_13613,N_13744);
and U13893 (N_13893,N_13703,N_13751);
nor U13894 (N_13894,N_13687,N_13682);
and U13895 (N_13895,N_13710,N_13711);
xnor U13896 (N_13896,N_13678,N_13757);
or U13897 (N_13897,N_13696,N_13638);
and U13898 (N_13898,N_13758,N_13745);
or U13899 (N_13899,N_13621,N_13709);
xnor U13900 (N_13900,N_13666,N_13707);
nor U13901 (N_13901,N_13709,N_13604);
nor U13902 (N_13902,N_13695,N_13738);
nor U13903 (N_13903,N_13601,N_13745);
nand U13904 (N_13904,N_13680,N_13627);
nor U13905 (N_13905,N_13648,N_13751);
and U13906 (N_13906,N_13676,N_13742);
or U13907 (N_13907,N_13710,N_13617);
xnor U13908 (N_13908,N_13707,N_13696);
nand U13909 (N_13909,N_13740,N_13628);
nand U13910 (N_13910,N_13617,N_13618);
nor U13911 (N_13911,N_13639,N_13610);
or U13912 (N_13912,N_13753,N_13714);
or U13913 (N_13913,N_13722,N_13615);
xnor U13914 (N_13914,N_13757,N_13719);
and U13915 (N_13915,N_13668,N_13677);
and U13916 (N_13916,N_13638,N_13707);
nand U13917 (N_13917,N_13663,N_13708);
xnor U13918 (N_13918,N_13716,N_13693);
and U13919 (N_13919,N_13618,N_13645);
and U13920 (N_13920,N_13880,N_13890);
xor U13921 (N_13921,N_13877,N_13798);
nor U13922 (N_13922,N_13769,N_13886);
and U13923 (N_13923,N_13825,N_13796);
nor U13924 (N_13924,N_13838,N_13811);
or U13925 (N_13925,N_13818,N_13774);
and U13926 (N_13926,N_13810,N_13815);
xnor U13927 (N_13927,N_13834,N_13804);
or U13928 (N_13928,N_13816,N_13782);
nor U13929 (N_13929,N_13775,N_13882);
or U13930 (N_13930,N_13794,N_13917);
or U13931 (N_13931,N_13845,N_13913);
xnor U13932 (N_13932,N_13781,N_13809);
or U13933 (N_13933,N_13916,N_13808);
nor U13934 (N_13934,N_13885,N_13849);
or U13935 (N_13935,N_13918,N_13822);
xnor U13936 (N_13936,N_13773,N_13907);
or U13937 (N_13937,N_13869,N_13832);
and U13938 (N_13938,N_13912,N_13883);
or U13939 (N_13939,N_13836,N_13891);
or U13940 (N_13940,N_13864,N_13771);
nand U13941 (N_13941,N_13813,N_13821);
and U13942 (N_13942,N_13795,N_13820);
xnor U13943 (N_13943,N_13814,N_13896);
nand U13944 (N_13944,N_13805,N_13862);
and U13945 (N_13945,N_13835,N_13853);
nor U13946 (N_13946,N_13860,N_13904);
xor U13947 (N_13947,N_13833,N_13839);
or U13948 (N_13948,N_13910,N_13841);
xnor U13949 (N_13949,N_13830,N_13766);
and U13950 (N_13950,N_13915,N_13878);
and U13951 (N_13951,N_13761,N_13800);
xor U13952 (N_13952,N_13779,N_13863);
nand U13953 (N_13953,N_13851,N_13899);
nor U13954 (N_13954,N_13884,N_13888);
nor U13955 (N_13955,N_13843,N_13777);
and U13956 (N_13956,N_13797,N_13789);
nand U13957 (N_13957,N_13889,N_13760);
or U13958 (N_13958,N_13778,N_13776);
and U13959 (N_13959,N_13859,N_13892);
nor U13960 (N_13960,N_13844,N_13850);
and U13961 (N_13961,N_13876,N_13903);
or U13962 (N_13962,N_13770,N_13823);
nor U13963 (N_13963,N_13764,N_13780);
or U13964 (N_13964,N_13765,N_13772);
xor U13965 (N_13965,N_13858,N_13799);
xnor U13966 (N_13966,N_13868,N_13829);
and U13967 (N_13967,N_13879,N_13897);
xor U13968 (N_13968,N_13763,N_13909);
nor U13969 (N_13969,N_13855,N_13906);
nand U13970 (N_13970,N_13865,N_13802);
nor U13971 (N_13971,N_13826,N_13828);
and U13972 (N_13972,N_13817,N_13872);
xnor U13973 (N_13973,N_13846,N_13900);
and U13974 (N_13974,N_13898,N_13807);
nand U13975 (N_13975,N_13827,N_13848);
and U13976 (N_13976,N_13783,N_13866);
and U13977 (N_13977,N_13852,N_13785);
and U13978 (N_13978,N_13875,N_13819);
or U13979 (N_13979,N_13831,N_13902);
nand U13980 (N_13980,N_13837,N_13840);
nand U13981 (N_13981,N_13905,N_13847);
nor U13982 (N_13982,N_13786,N_13914);
or U13983 (N_13983,N_13893,N_13801);
nand U13984 (N_13984,N_13856,N_13824);
and U13985 (N_13985,N_13842,N_13871);
nand U13986 (N_13986,N_13870,N_13867);
nand U13987 (N_13987,N_13887,N_13854);
nand U13988 (N_13988,N_13908,N_13787);
nand U13989 (N_13989,N_13767,N_13857);
and U13990 (N_13990,N_13874,N_13911);
or U13991 (N_13991,N_13790,N_13901);
nor U13992 (N_13992,N_13812,N_13803);
xnor U13993 (N_13993,N_13784,N_13881);
nor U13994 (N_13994,N_13919,N_13894);
nand U13995 (N_13995,N_13792,N_13788);
and U13996 (N_13996,N_13793,N_13861);
xnor U13997 (N_13997,N_13768,N_13873);
nor U13998 (N_13998,N_13791,N_13806);
or U13999 (N_13999,N_13762,N_13895);
nor U14000 (N_14000,N_13823,N_13887);
and U14001 (N_14001,N_13838,N_13877);
and U14002 (N_14002,N_13843,N_13895);
nor U14003 (N_14003,N_13919,N_13828);
and U14004 (N_14004,N_13851,N_13826);
or U14005 (N_14005,N_13913,N_13799);
nor U14006 (N_14006,N_13773,N_13803);
nor U14007 (N_14007,N_13814,N_13907);
or U14008 (N_14008,N_13915,N_13817);
and U14009 (N_14009,N_13872,N_13847);
xnor U14010 (N_14010,N_13864,N_13809);
xor U14011 (N_14011,N_13897,N_13878);
or U14012 (N_14012,N_13778,N_13780);
nand U14013 (N_14013,N_13888,N_13770);
nand U14014 (N_14014,N_13845,N_13912);
xor U14015 (N_14015,N_13843,N_13915);
xnor U14016 (N_14016,N_13856,N_13833);
nand U14017 (N_14017,N_13894,N_13804);
nand U14018 (N_14018,N_13826,N_13816);
or U14019 (N_14019,N_13911,N_13787);
nand U14020 (N_14020,N_13859,N_13867);
or U14021 (N_14021,N_13850,N_13900);
or U14022 (N_14022,N_13818,N_13847);
xor U14023 (N_14023,N_13806,N_13881);
nor U14024 (N_14024,N_13835,N_13818);
nand U14025 (N_14025,N_13794,N_13798);
xnor U14026 (N_14026,N_13879,N_13849);
nor U14027 (N_14027,N_13784,N_13913);
nand U14028 (N_14028,N_13839,N_13835);
nand U14029 (N_14029,N_13798,N_13766);
nand U14030 (N_14030,N_13864,N_13867);
or U14031 (N_14031,N_13892,N_13876);
xnor U14032 (N_14032,N_13794,N_13904);
nor U14033 (N_14033,N_13785,N_13881);
xnor U14034 (N_14034,N_13772,N_13784);
or U14035 (N_14035,N_13854,N_13828);
and U14036 (N_14036,N_13798,N_13800);
and U14037 (N_14037,N_13783,N_13775);
xnor U14038 (N_14038,N_13776,N_13831);
or U14039 (N_14039,N_13829,N_13828);
and U14040 (N_14040,N_13846,N_13843);
nor U14041 (N_14041,N_13788,N_13786);
and U14042 (N_14042,N_13808,N_13896);
nand U14043 (N_14043,N_13794,N_13902);
and U14044 (N_14044,N_13917,N_13835);
or U14045 (N_14045,N_13879,N_13885);
xor U14046 (N_14046,N_13795,N_13868);
nand U14047 (N_14047,N_13869,N_13833);
xnor U14048 (N_14048,N_13881,N_13850);
and U14049 (N_14049,N_13766,N_13867);
or U14050 (N_14050,N_13767,N_13788);
nand U14051 (N_14051,N_13846,N_13905);
or U14052 (N_14052,N_13851,N_13883);
xor U14053 (N_14053,N_13839,N_13773);
and U14054 (N_14054,N_13831,N_13843);
and U14055 (N_14055,N_13819,N_13844);
nand U14056 (N_14056,N_13895,N_13847);
or U14057 (N_14057,N_13766,N_13906);
nor U14058 (N_14058,N_13859,N_13804);
nor U14059 (N_14059,N_13873,N_13898);
nand U14060 (N_14060,N_13862,N_13760);
and U14061 (N_14061,N_13809,N_13896);
or U14062 (N_14062,N_13884,N_13900);
nor U14063 (N_14063,N_13901,N_13767);
nor U14064 (N_14064,N_13845,N_13849);
nand U14065 (N_14065,N_13806,N_13900);
or U14066 (N_14066,N_13837,N_13791);
nand U14067 (N_14067,N_13889,N_13894);
nor U14068 (N_14068,N_13843,N_13793);
nand U14069 (N_14069,N_13889,N_13814);
nand U14070 (N_14070,N_13862,N_13874);
xnor U14071 (N_14071,N_13821,N_13830);
or U14072 (N_14072,N_13885,N_13800);
and U14073 (N_14073,N_13834,N_13777);
or U14074 (N_14074,N_13776,N_13892);
and U14075 (N_14075,N_13824,N_13886);
or U14076 (N_14076,N_13821,N_13774);
xor U14077 (N_14077,N_13874,N_13842);
and U14078 (N_14078,N_13813,N_13860);
nand U14079 (N_14079,N_13866,N_13877);
xor U14080 (N_14080,N_13962,N_14055);
xnor U14081 (N_14081,N_14064,N_14015);
and U14082 (N_14082,N_14025,N_14047);
or U14083 (N_14083,N_13949,N_14040);
xor U14084 (N_14084,N_13994,N_14078);
nor U14085 (N_14085,N_13995,N_13991);
xnor U14086 (N_14086,N_13933,N_13986);
nand U14087 (N_14087,N_14039,N_13940);
and U14088 (N_14088,N_13980,N_13938);
nand U14089 (N_14089,N_14036,N_14062);
or U14090 (N_14090,N_13989,N_13961);
nor U14091 (N_14091,N_13957,N_14073);
nor U14092 (N_14092,N_14066,N_14071);
and U14093 (N_14093,N_14075,N_14049);
or U14094 (N_14094,N_13974,N_14001);
or U14095 (N_14095,N_14045,N_14021);
xor U14096 (N_14096,N_13985,N_14000);
or U14097 (N_14097,N_13999,N_14059);
nand U14098 (N_14098,N_14027,N_13956);
xor U14099 (N_14099,N_13976,N_14005);
nand U14100 (N_14100,N_14060,N_13923);
nor U14101 (N_14101,N_13955,N_14028);
xnor U14102 (N_14102,N_13947,N_14011);
xor U14103 (N_14103,N_14004,N_13964);
nand U14104 (N_14104,N_14032,N_14031);
or U14105 (N_14105,N_13936,N_14044);
and U14106 (N_14106,N_14019,N_13987);
nand U14107 (N_14107,N_13992,N_14070);
xnor U14108 (N_14108,N_14042,N_13941);
or U14109 (N_14109,N_14053,N_13968);
xnor U14110 (N_14110,N_14034,N_13982);
and U14111 (N_14111,N_13973,N_13939);
or U14112 (N_14112,N_14006,N_14043);
nor U14113 (N_14113,N_13942,N_14003);
and U14114 (N_14114,N_13997,N_14010);
nand U14115 (N_14115,N_14013,N_14012);
or U14116 (N_14116,N_14037,N_13981);
nor U14117 (N_14117,N_14018,N_13953);
nand U14118 (N_14118,N_14016,N_13934);
or U14119 (N_14119,N_13998,N_13978);
xnor U14120 (N_14120,N_14033,N_13963);
or U14121 (N_14121,N_13931,N_13935);
nor U14122 (N_14122,N_14020,N_14052);
nand U14123 (N_14123,N_14035,N_14029);
and U14124 (N_14124,N_14023,N_14007);
and U14125 (N_14125,N_14058,N_14076);
nor U14126 (N_14126,N_13924,N_13946);
nand U14127 (N_14127,N_13959,N_13966);
nand U14128 (N_14128,N_14079,N_13990);
nand U14129 (N_14129,N_13920,N_14061);
nand U14130 (N_14130,N_13951,N_13928);
or U14131 (N_14131,N_13970,N_14051);
nand U14132 (N_14132,N_13950,N_14014);
nor U14133 (N_14133,N_13943,N_14024);
and U14134 (N_14134,N_13922,N_14069);
nand U14135 (N_14135,N_13979,N_14065);
and U14136 (N_14136,N_13977,N_14017);
and U14137 (N_14137,N_14009,N_13948);
xnor U14138 (N_14138,N_13929,N_14072);
xnor U14139 (N_14139,N_13952,N_13958);
or U14140 (N_14140,N_13954,N_14074);
or U14141 (N_14141,N_14008,N_14057);
xor U14142 (N_14142,N_13927,N_13971);
nor U14143 (N_14143,N_13969,N_13993);
nand U14144 (N_14144,N_13975,N_14022);
or U14145 (N_14145,N_14038,N_13972);
nand U14146 (N_14146,N_13988,N_14054);
xor U14147 (N_14147,N_14067,N_14002);
or U14148 (N_14148,N_14068,N_13926);
nor U14149 (N_14149,N_13983,N_13965);
nor U14150 (N_14150,N_14077,N_14056);
or U14151 (N_14151,N_14063,N_13984);
nor U14152 (N_14152,N_13925,N_13932);
nand U14153 (N_14153,N_13960,N_14026);
xor U14154 (N_14154,N_14048,N_13996);
or U14155 (N_14155,N_13921,N_13930);
and U14156 (N_14156,N_13944,N_14046);
and U14157 (N_14157,N_13967,N_14050);
and U14158 (N_14158,N_14041,N_13945);
and U14159 (N_14159,N_14030,N_13937);
or U14160 (N_14160,N_14079,N_13962);
xnor U14161 (N_14161,N_14064,N_14046);
nor U14162 (N_14162,N_13994,N_13926);
and U14163 (N_14163,N_13984,N_14079);
nor U14164 (N_14164,N_13929,N_14006);
or U14165 (N_14165,N_13992,N_13930);
nor U14166 (N_14166,N_14045,N_13990);
xor U14167 (N_14167,N_13972,N_13926);
xor U14168 (N_14168,N_13944,N_13926);
xnor U14169 (N_14169,N_14064,N_14014);
xnor U14170 (N_14170,N_13999,N_14000);
nand U14171 (N_14171,N_14025,N_14029);
or U14172 (N_14172,N_14045,N_14054);
nor U14173 (N_14173,N_13941,N_13932);
and U14174 (N_14174,N_13979,N_14030);
xnor U14175 (N_14175,N_14053,N_13959);
xor U14176 (N_14176,N_14008,N_13988);
xnor U14177 (N_14177,N_14017,N_14041);
nand U14178 (N_14178,N_14072,N_14048);
nand U14179 (N_14179,N_14050,N_14063);
nand U14180 (N_14180,N_13922,N_13989);
nor U14181 (N_14181,N_13954,N_13955);
or U14182 (N_14182,N_13979,N_13991);
and U14183 (N_14183,N_13921,N_13936);
and U14184 (N_14184,N_14012,N_13959);
xor U14185 (N_14185,N_13922,N_13951);
nand U14186 (N_14186,N_14021,N_13962);
nand U14187 (N_14187,N_14051,N_13995);
nor U14188 (N_14188,N_14055,N_13968);
xnor U14189 (N_14189,N_14074,N_14041);
nor U14190 (N_14190,N_13988,N_13924);
xor U14191 (N_14191,N_14002,N_13989);
nor U14192 (N_14192,N_14041,N_13998);
nor U14193 (N_14193,N_14046,N_14026);
xnor U14194 (N_14194,N_13945,N_13957);
xnor U14195 (N_14195,N_14008,N_14000);
nor U14196 (N_14196,N_14039,N_14010);
and U14197 (N_14197,N_13996,N_14067);
nand U14198 (N_14198,N_13975,N_13924);
nand U14199 (N_14199,N_14007,N_14043);
nor U14200 (N_14200,N_13982,N_13959);
and U14201 (N_14201,N_14027,N_13948);
nand U14202 (N_14202,N_13938,N_14013);
and U14203 (N_14203,N_13947,N_13988);
xnor U14204 (N_14204,N_13938,N_14021);
or U14205 (N_14205,N_14059,N_13940);
nor U14206 (N_14206,N_14004,N_14074);
and U14207 (N_14207,N_14009,N_14078);
nor U14208 (N_14208,N_13973,N_14008);
xnor U14209 (N_14209,N_14023,N_14046);
and U14210 (N_14210,N_13928,N_14010);
or U14211 (N_14211,N_13991,N_13949);
and U14212 (N_14212,N_13966,N_13930);
and U14213 (N_14213,N_13951,N_14059);
nor U14214 (N_14214,N_13986,N_14059);
and U14215 (N_14215,N_14025,N_14056);
or U14216 (N_14216,N_14074,N_13928);
or U14217 (N_14217,N_13921,N_14019);
nand U14218 (N_14218,N_14066,N_14057);
nor U14219 (N_14219,N_14025,N_13925);
nand U14220 (N_14220,N_14059,N_14063);
and U14221 (N_14221,N_13927,N_13949);
xor U14222 (N_14222,N_13979,N_13946);
and U14223 (N_14223,N_13964,N_13972);
xnor U14224 (N_14224,N_13981,N_13931);
and U14225 (N_14225,N_14069,N_14038);
nor U14226 (N_14226,N_13990,N_14011);
or U14227 (N_14227,N_14052,N_14058);
or U14228 (N_14228,N_13994,N_14067);
or U14229 (N_14229,N_14002,N_14036);
xnor U14230 (N_14230,N_13925,N_13946);
and U14231 (N_14231,N_14013,N_13950);
or U14232 (N_14232,N_14013,N_14007);
or U14233 (N_14233,N_13988,N_13954);
and U14234 (N_14234,N_13944,N_13975);
and U14235 (N_14235,N_14021,N_13922);
and U14236 (N_14236,N_13956,N_13921);
or U14237 (N_14237,N_14049,N_14042);
or U14238 (N_14238,N_14029,N_13968);
and U14239 (N_14239,N_13987,N_14075);
xnor U14240 (N_14240,N_14111,N_14167);
and U14241 (N_14241,N_14122,N_14196);
nand U14242 (N_14242,N_14164,N_14114);
and U14243 (N_14243,N_14177,N_14084);
xnor U14244 (N_14244,N_14113,N_14104);
nand U14245 (N_14245,N_14232,N_14217);
or U14246 (N_14246,N_14187,N_14168);
or U14247 (N_14247,N_14159,N_14179);
and U14248 (N_14248,N_14185,N_14192);
nor U14249 (N_14249,N_14086,N_14216);
and U14250 (N_14250,N_14172,N_14095);
nor U14251 (N_14251,N_14207,N_14153);
xor U14252 (N_14252,N_14118,N_14218);
xor U14253 (N_14253,N_14098,N_14150);
nor U14254 (N_14254,N_14091,N_14125);
or U14255 (N_14255,N_14169,N_14230);
or U14256 (N_14256,N_14180,N_14120);
or U14257 (N_14257,N_14092,N_14204);
nor U14258 (N_14258,N_14239,N_14210);
and U14259 (N_14259,N_14191,N_14189);
nor U14260 (N_14260,N_14213,N_14130);
and U14261 (N_14261,N_14165,N_14119);
nor U14262 (N_14262,N_14101,N_14214);
and U14263 (N_14263,N_14158,N_14188);
nand U14264 (N_14264,N_14147,N_14211);
and U14265 (N_14265,N_14176,N_14121);
and U14266 (N_14266,N_14154,N_14134);
and U14267 (N_14267,N_14083,N_14144);
nand U14268 (N_14268,N_14112,N_14182);
nor U14269 (N_14269,N_14234,N_14199);
nand U14270 (N_14270,N_14116,N_14103);
or U14271 (N_14271,N_14190,N_14227);
nor U14272 (N_14272,N_14161,N_14221);
or U14273 (N_14273,N_14142,N_14094);
nand U14274 (N_14274,N_14110,N_14215);
or U14275 (N_14275,N_14096,N_14184);
xnor U14276 (N_14276,N_14115,N_14152);
or U14277 (N_14277,N_14198,N_14133);
xor U14278 (N_14278,N_14146,N_14219);
nand U14279 (N_14279,N_14089,N_14206);
nor U14280 (N_14280,N_14123,N_14201);
nor U14281 (N_14281,N_14195,N_14229);
or U14282 (N_14282,N_14151,N_14223);
nor U14283 (N_14283,N_14212,N_14193);
or U14284 (N_14284,N_14108,N_14238);
xnor U14285 (N_14285,N_14087,N_14107);
nor U14286 (N_14286,N_14131,N_14170);
nand U14287 (N_14287,N_14178,N_14203);
nor U14288 (N_14288,N_14208,N_14156);
xnor U14289 (N_14289,N_14149,N_14132);
and U14290 (N_14290,N_14231,N_14085);
nor U14291 (N_14291,N_14126,N_14162);
or U14292 (N_14292,N_14127,N_14102);
nor U14293 (N_14293,N_14175,N_14090);
xor U14294 (N_14294,N_14171,N_14093);
or U14295 (N_14295,N_14088,N_14155);
nor U14296 (N_14296,N_14138,N_14200);
or U14297 (N_14297,N_14140,N_14143);
xor U14298 (N_14298,N_14100,N_14157);
or U14299 (N_14299,N_14181,N_14137);
nand U14300 (N_14300,N_14237,N_14222);
nor U14301 (N_14301,N_14124,N_14233);
nand U14302 (N_14302,N_14082,N_14080);
xnor U14303 (N_14303,N_14183,N_14148);
or U14304 (N_14304,N_14174,N_14141);
and U14305 (N_14305,N_14235,N_14106);
xor U14306 (N_14306,N_14197,N_14186);
and U14307 (N_14307,N_14224,N_14117);
and U14308 (N_14308,N_14135,N_14097);
or U14309 (N_14309,N_14139,N_14166);
nor U14310 (N_14310,N_14081,N_14220);
or U14311 (N_14311,N_14226,N_14173);
nand U14312 (N_14312,N_14209,N_14160);
nor U14313 (N_14313,N_14099,N_14202);
or U14314 (N_14314,N_14145,N_14136);
or U14315 (N_14315,N_14105,N_14236);
or U14316 (N_14316,N_14228,N_14109);
xor U14317 (N_14317,N_14194,N_14128);
or U14318 (N_14318,N_14129,N_14225);
nor U14319 (N_14319,N_14205,N_14163);
xor U14320 (N_14320,N_14209,N_14094);
xor U14321 (N_14321,N_14147,N_14121);
xnor U14322 (N_14322,N_14141,N_14100);
nor U14323 (N_14323,N_14139,N_14099);
nor U14324 (N_14324,N_14234,N_14119);
nand U14325 (N_14325,N_14203,N_14091);
xnor U14326 (N_14326,N_14108,N_14136);
xor U14327 (N_14327,N_14217,N_14210);
nand U14328 (N_14328,N_14131,N_14081);
and U14329 (N_14329,N_14201,N_14228);
or U14330 (N_14330,N_14099,N_14130);
xor U14331 (N_14331,N_14206,N_14136);
xor U14332 (N_14332,N_14112,N_14217);
and U14333 (N_14333,N_14169,N_14104);
and U14334 (N_14334,N_14145,N_14088);
nand U14335 (N_14335,N_14174,N_14084);
nor U14336 (N_14336,N_14151,N_14081);
and U14337 (N_14337,N_14165,N_14204);
nor U14338 (N_14338,N_14173,N_14238);
xnor U14339 (N_14339,N_14160,N_14101);
nand U14340 (N_14340,N_14133,N_14222);
or U14341 (N_14341,N_14239,N_14182);
nand U14342 (N_14342,N_14173,N_14108);
nor U14343 (N_14343,N_14169,N_14194);
or U14344 (N_14344,N_14219,N_14091);
xor U14345 (N_14345,N_14080,N_14171);
xnor U14346 (N_14346,N_14096,N_14165);
nor U14347 (N_14347,N_14089,N_14098);
or U14348 (N_14348,N_14209,N_14132);
or U14349 (N_14349,N_14124,N_14173);
xor U14350 (N_14350,N_14186,N_14204);
nand U14351 (N_14351,N_14114,N_14120);
xnor U14352 (N_14352,N_14153,N_14084);
nand U14353 (N_14353,N_14173,N_14214);
nor U14354 (N_14354,N_14086,N_14225);
nor U14355 (N_14355,N_14153,N_14156);
and U14356 (N_14356,N_14140,N_14198);
or U14357 (N_14357,N_14190,N_14153);
nor U14358 (N_14358,N_14136,N_14097);
nor U14359 (N_14359,N_14170,N_14195);
xor U14360 (N_14360,N_14165,N_14170);
nor U14361 (N_14361,N_14158,N_14183);
nor U14362 (N_14362,N_14153,N_14214);
xor U14363 (N_14363,N_14136,N_14153);
or U14364 (N_14364,N_14239,N_14216);
xor U14365 (N_14365,N_14164,N_14174);
nor U14366 (N_14366,N_14230,N_14107);
nand U14367 (N_14367,N_14082,N_14215);
or U14368 (N_14368,N_14112,N_14239);
nand U14369 (N_14369,N_14218,N_14096);
nor U14370 (N_14370,N_14227,N_14103);
and U14371 (N_14371,N_14133,N_14197);
or U14372 (N_14372,N_14227,N_14200);
and U14373 (N_14373,N_14113,N_14091);
nor U14374 (N_14374,N_14198,N_14232);
and U14375 (N_14375,N_14085,N_14176);
nor U14376 (N_14376,N_14138,N_14207);
nor U14377 (N_14377,N_14101,N_14121);
nand U14378 (N_14378,N_14122,N_14157);
or U14379 (N_14379,N_14144,N_14200);
nor U14380 (N_14380,N_14110,N_14235);
and U14381 (N_14381,N_14202,N_14085);
nor U14382 (N_14382,N_14156,N_14080);
nor U14383 (N_14383,N_14144,N_14127);
nor U14384 (N_14384,N_14194,N_14157);
nor U14385 (N_14385,N_14080,N_14089);
nand U14386 (N_14386,N_14208,N_14179);
xor U14387 (N_14387,N_14121,N_14143);
nand U14388 (N_14388,N_14107,N_14102);
nand U14389 (N_14389,N_14132,N_14082);
xnor U14390 (N_14390,N_14127,N_14105);
nand U14391 (N_14391,N_14090,N_14181);
and U14392 (N_14392,N_14195,N_14096);
nor U14393 (N_14393,N_14233,N_14112);
and U14394 (N_14394,N_14115,N_14220);
nor U14395 (N_14395,N_14153,N_14192);
nor U14396 (N_14396,N_14092,N_14120);
or U14397 (N_14397,N_14192,N_14152);
nand U14398 (N_14398,N_14171,N_14221);
and U14399 (N_14399,N_14138,N_14120);
xor U14400 (N_14400,N_14263,N_14338);
nand U14401 (N_14401,N_14315,N_14290);
nand U14402 (N_14402,N_14308,N_14339);
xnor U14403 (N_14403,N_14346,N_14318);
nor U14404 (N_14404,N_14387,N_14385);
or U14405 (N_14405,N_14324,N_14395);
and U14406 (N_14406,N_14382,N_14342);
xnor U14407 (N_14407,N_14357,N_14379);
and U14408 (N_14408,N_14270,N_14278);
and U14409 (N_14409,N_14283,N_14310);
nor U14410 (N_14410,N_14241,N_14302);
nor U14411 (N_14411,N_14266,N_14358);
xor U14412 (N_14412,N_14394,N_14343);
nand U14413 (N_14413,N_14336,N_14361);
or U14414 (N_14414,N_14363,N_14299);
or U14415 (N_14415,N_14288,N_14389);
xor U14416 (N_14416,N_14268,N_14260);
xor U14417 (N_14417,N_14304,N_14291);
nor U14418 (N_14418,N_14255,N_14269);
and U14419 (N_14419,N_14327,N_14275);
nor U14420 (N_14420,N_14261,N_14352);
nor U14421 (N_14421,N_14254,N_14284);
and U14422 (N_14422,N_14277,N_14380);
nand U14423 (N_14423,N_14355,N_14370);
nor U14424 (N_14424,N_14372,N_14320);
and U14425 (N_14425,N_14319,N_14386);
nand U14426 (N_14426,N_14248,N_14313);
nand U14427 (N_14427,N_14341,N_14398);
xor U14428 (N_14428,N_14340,N_14331);
and U14429 (N_14429,N_14337,N_14276);
nor U14430 (N_14430,N_14396,N_14374);
or U14431 (N_14431,N_14371,N_14246);
xnor U14432 (N_14432,N_14264,N_14292);
nand U14433 (N_14433,N_14345,N_14381);
and U14434 (N_14434,N_14303,N_14383);
or U14435 (N_14435,N_14256,N_14328);
or U14436 (N_14436,N_14362,N_14258);
nor U14437 (N_14437,N_14306,N_14344);
and U14438 (N_14438,N_14273,N_14294);
xnor U14439 (N_14439,N_14356,N_14243);
or U14440 (N_14440,N_14373,N_14347);
nor U14441 (N_14441,N_14271,N_14330);
xor U14442 (N_14442,N_14287,N_14250);
and U14443 (N_14443,N_14388,N_14390);
or U14444 (N_14444,N_14274,N_14242);
xnor U14445 (N_14445,N_14350,N_14399);
and U14446 (N_14446,N_14296,N_14323);
xnor U14447 (N_14447,N_14349,N_14384);
nor U14448 (N_14448,N_14367,N_14392);
nor U14449 (N_14449,N_14314,N_14280);
nor U14450 (N_14450,N_14249,N_14240);
or U14451 (N_14451,N_14368,N_14348);
nand U14452 (N_14452,N_14316,N_14251);
nand U14453 (N_14453,N_14311,N_14245);
and U14454 (N_14454,N_14285,N_14282);
or U14455 (N_14455,N_14317,N_14378);
nor U14456 (N_14456,N_14393,N_14300);
nor U14457 (N_14457,N_14253,N_14360);
nor U14458 (N_14458,N_14369,N_14377);
nand U14459 (N_14459,N_14321,N_14259);
nand U14460 (N_14460,N_14325,N_14295);
xnor U14461 (N_14461,N_14365,N_14333);
and U14462 (N_14462,N_14329,N_14257);
nor U14463 (N_14463,N_14322,N_14289);
xnor U14464 (N_14464,N_14305,N_14359);
xor U14465 (N_14465,N_14297,N_14334);
and U14466 (N_14466,N_14351,N_14279);
nor U14467 (N_14467,N_14286,N_14312);
nor U14468 (N_14468,N_14281,N_14353);
nor U14469 (N_14469,N_14244,N_14332);
xor U14470 (N_14470,N_14298,N_14364);
nor U14471 (N_14471,N_14307,N_14301);
or U14472 (N_14472,N_14267,N_14293);
xnor U14473 (N_14473,N_14375,N_14265);
or U14474 (N_14474,N_14354,N_14252);
or U14475 (N_14475,N_14272,N_14366);
nor U14476 (N_14476,N_14391,N_14247);
and U14477 (N_14477,N_14376,N_14262);
nand U14478 (N_14478,N_14326,N_14335);
or U14479 (N_14479,N_14309,N_14397);
xnor U14480 (N_14480,N_14332,N_14272);
xnor U14481 (N_14481,N_14325,N_14393);
nand U14482 (N_14482,N_14265,N_14250);
and U14483 (N_14483,N_14387,N_14395);
and U14484 (N_14484,N_14319,N_14314);
or U14485 (N_14485,N_14326,N_14371);
xnor U14486 (N_14486,N_14294,N_14355);
xnor U14487 (N_14487,N_14279,N_14369);
and U14488 (N_14488,N_14330,N_14354);
or U14489 (N_14489,N_14372,N_14306);
nor U14490 (N_14490,N_14254,N_14299);
or U14491 (N_14491,N_14360,N_14359);
and U14492 (N_14492,N_14256,N_14370);
nand U14493 (N_14493,N_14351,N_14395);
nand U14494 (N_14494,N_14317,N_14341);
xnor U14495 (N_14495,N_14376,N_14365);
and U14496 (N_14496,N_14267,N_14278);
nor U14497 (N_14497,N_14332,N_14273);
or U14498 (N_14498,N_14246,N_14381);
nand U14499 (N_14499,N_14359,N_14346);
and U14500 (N_14500,N_14396,N_14335);
xnor U14501 (N_14501,N_14272,N_14373);
nand U14502 (N_14502,N_14318,N_14244);
or U14503 (N_14503,N_14312,N_14278);
nand U14504 (N_14504,N_14259,N_14283);
nor U14505 (N_14505,N_14271,N_14389);
nor U14506 (N_14506,N_14333,N_14334);
and U14507 (N_14507,N_14263,N_14349);
xor U14508 (N_14508,N_14246,N_14263);
nor U14509 (N_14509,N_14331,N_14303);
or U14510 (N_14510,N_14370,N_14251);
nand U14511 (N_14511,N_14274,N_14359);
and U14512 (N_14512,N_14390,N_14357);
xor U14513 (N_14513,N_14306,N_14362);
nand U14514 (N_14514,N_14343,N_14384);
or U14515 (N_14515,N_14282,N_14362);
or U14516 (N_14516,N_14269,N_14274);
nand U14517 (N_14517,N_14285,N_14399);
nand U14518 (N_14518,N_14332,N_14361);
or U14519 (N_14519,N_14345,N_14256);
nand U14520 (N_14520,N_14272,N_14276);
or U14521 (N_14521,N_14283,N_14247);
xor U14522 (N_14522,N_14388,N_14365);
nand U14523 (N_14523,N_14339,N_14269);
xor U14524 (N_14524,N_14363,N_14379);
xor U14525 (N_14525,N_14322,N_14395);
or U14526 (N_14526,N_14269,N_14320);
nor U14527 (N_14527,N_14370,N_14399);
nand U14528 (N_14528,N_14326,N_14266);
nor U14529 (N_14529,N_14309,N_14248);
or U14530 (N_14530,N_14331,N_14338);
nor U14531 (N_14531,N_14376,N_14395);
or U14532 (N_14532,N_14295,N_14284);
or U14533 (N_14533,N_14328,N_14245);
and U14534 (N_14534,N_14248,N_14302);
and U14535 (N_14535,N_14304,N_14311);
nand U14536 (N_14536,N_14268,N_14395);
xor U14537 (N_14537,N_14364,N_14294);
and U14538 (N_14538,N_14320,N_14356);
nand U14539 (N_14539,N_14245,N_14333);
xnor U14540 (N_14540,N_14329,N_14343);
nor U14541 (N_14541,N_14299,N_14351);
xor U14542 (N_14542,N_14244,N_14387);
nand U14543 (N_14543,N_14275,N_14355);
xor U14544 (N_14544,N_14250,N_14320);
nor U14545 (N_14545,N_14372,N_14387);
xnor U14546 (N_14546,N_14349,N_14335);
nor U14547 (N_14547,N_14290,N_14287);
nor U14548 (N_14548,N_14355,N_14263);
or U14549 (N_14549,N_14305,N_14243);
nor U14550 (N_14550,N_14340,N_14319);
xnor U14551 (N_14551,N_14303,N_14282);
nand U14552 (N_14552,N_14298,N_14390);
xor U14553 (N_14553,N_14261,N_14365);
and U14554 (N_14554,N_14343,N_14291);
nand U14555 (N_14555,N_14269,N_14342);
nand U14556 (N_14556,N_14386,N_14331);
xnor U14557 (N_14557,N_14398,N_14389);
nand U14558 (N_14558,N_14380,N_14370);
xnor U14559 (N_14559,N_14290,N_14362);
xor U14560 (N_14560,N_14403,N_14421);
nor U14561 (N_14561,N_14446,N_14441);
nor U14562 (N_14562,N_14555,N_14419);
or U14563 (N_14563,N_14401,N_14556);
nor U14564 (N_14564,N_14461,N_14542);
nand U14565 (N_14565,N_14482,N_14536);
and U14566 (N_14566,N_14510,N_14455);
xnor U14567 (N_14567,N_14504,N_14491);
and U14568 (N_14568,N_14520,N_14554);
nor U14569 (N_14569,N_14474,N_14532);
nor U14570 (N_14570,N_14503,N_14518);
xor U14571 (N_14571,N_14546,N_14457);
nor U14572 (N_14572,N_14407,N_14488);
nor U14573 (N_14573,N_14534,N_14456);
nor U14574 (N_14574,N_14438,N_14454);
nand U14575 (N_14575,N_14436,N_14423);
nor U14576 (N_14576,N_14558,N_14526);
xnor U14577 (N_14577,N_14535,N_14462);
nor U14578 (N_14578,N_14525,N_14434);
xnor U14579 (N_14579,N_14411,N_14402);
nor U14580 (N_14580,N_14447,N_14553);
nand U14581 (N_14581,N_14527,N_14501);
and U14582 (N_14582,N_14524,N_14470);
xnor U14583 (N_14583,N_14549,N_14418);
nand U14584 (N_14584,N_14499,N_14439);
and U14585 (N_14585,N_14404,N_14494);
xnor U14586 (N_14586,N_14475,N_14471);
xor U14587 (N_14587,N_14519,N_14427);
nor U14588 (N_14588,N_14417,N_14481);
and U14589 (N_14589,N_14548,N_14483);
xnor U14590 (N_14590,N_14522,N_14550);
xnor U14591 (N_14591,N_14523,N_14476);
or U14592 (N_14592,N_14502,N_14517);
nor U14593 (N_14593,N_14493,N_14409);
and U14594 (N_14594,N_14406,N_14500);
and U14595 (N_14595,N_14508,N_14511);
and U14596 (N_14596,N_14528,N_14521);
nor U14597 (N_14597,N_14533,N_14452);
nor U14598 (N_14598,N_14413,N_14453);
nor U14599 (N_14599,N_14405,N_14431);
or U14600 (N_14600,N_14540,N_14420);
or U14601 (N_14601,N_14465,N_14435);
nor U14602 (N_14602,N_14545,N_14486);
or U14603 (N_14603,N_14530,N_14450);
xor U14604 (N_14604,N_14469,N_14551);
nand U14605 (N_14605,N_14468,N_14505);
nor U14606 (N_14606,N_14445,N_14480);
nand U14607 (N_14607,N_14492,N_14425);
nand U14608 (N_14608,N_14464,N_14539);
xor U14609 (N_14609,N_14489,N_14490);
or U14610 (N_14610,N_14440,N_14408);
nand U14611 (N_14611,N_14544,N_14463);
xor U14612 (N_14612,N_14498,N_14484);
nor U14613 (N_14613,N_14430,N_14429);
and U14614 (N_14614,N_14459,N_14538);
nand U14615 (N_14615,N_14444,N_14414);
nor U14616 (N_14616,N_14516,N_14443);
nand U14617 (N_14617,N_14478,N_14412);
and U14618 (N_14618,N_14426,N_14437);
nand U14619 (N_14619,N_14410,N_14433);
or U14620 (N_14620,N_14416,N_14557);
or U14621 (N_14621,N_14541,N_14424);
or U14622 (N_14622,N_14537,N_14448);
and U14623 (N_14623,N_14509,N_14473);
or U14624 (N_14624,N_14496,N_14479);
and U14625 (N_14625,N_14458,N_14497);
or U14626 (N_14626,N_14531,N_14547);
and U14627 (N_14627,N_14506,N_14472);
and U14628 (N_14628,N_14400,N_14477);
and U14629 (N_14629,N_14422,N_14559);
xnor U14630 (N_14630,N_14466,N_14507);
nor U14631 (N_14631,N_14529,N_14449);
or U14632 (N_14632,N_14467,N_14543);
or U14633 (N_14633,N_14432,N_14442);
and U14634 (N_14634,N_14485,N_14487);
and U14635 (N_14635,N_14428,N_14495);
or U14636 (N_14636,N_14451,N_14552);
nand U14637 (N_14637,N_14515,N_14415);
or U14638 (N_14638,N_14513,N_14514);
xnor U14639 (N_14639,N_14460,N_14512);
and U14640 (N_14640,N_14542,N_14423);
nand U14641 (N_14641,N_14537,N_14457);
xnor U14642 (N_14642,N_14522,N_14475);
nor U14643 (N_14643,N_14439,N_14447);
or U14644 (N_14644,N_14444,N_14408);
and U14645 (N_14645,N_14557,N_14403);
or U14646 (N_14646,N_14445,N_14476);
nand U14647 (N_14647,N_14425,N_14548);
nand U14648 (N_14648,N_14559,N_14410);
and U14649 (N_14649,N_14511,N_14457);
nor U14650 (N_14650,N_14415,N_14445);
or U14651 (N_14651,N_14461,N_14467);
nand U14652 (N_14652,N_14412,N_14502);
xnor U14653 (N_14653,N_14475,N_14553);
xor U14654 (N_14654,N_14441,N_14480);
nand U14655 (N_14655,N_14544,N_14551);
nand U14656 (N_14656,N_14503,N_14400);
xor U14657 (N_14657,N_14553,N_14403);
xor U14658 (N_14658,N_14492,N_14484);
and U14659 (N_14659,N_14464,N_14482);
xor U14660 (N_14660,N_14541,N_14418);
and U14661 (N_14661,N_14435,N_14424);
nor U14662 (N_14662,N_14494,N_14512);
and U14663 (N_14663,N_14409,N_14503);
and U14664 (N_14664,N_14454,N_14494);
nand U14665 (N_14665,N_14500,N_14534);
nand U14666 (N_14666,N_14427,N_14453);
nor U14667 (N_14667,N_14427,N_14523);
or U14668 (N_14668,N_14523,N_14401);
xor U14669 (N_14669,N_14414,N_14526);
xnor U14670 (N_14670,N_14474,N_14468);
nor U14671 (N_14671,N_14457,N_14544);
nor U14672 (N_14672,N_14439,N_14479);
nor U14673 (N_14673,N_14492,N_14541);
xor U14674 (N_14674,N_14467,N_14435);
or U14675 (N_14675,N_14408,N_14506);
nand U14676 (N_14676,N_14403,N_14521);
and U14677 (N_14677,N_14425,N_14428);
xor U14678 (N_14678,N_14444,N_14485);
or U14679 (N_14679,N_14483,N_14501);
xor U14680 (N_14680,N_14529,N_14465);
or U14681 (N_14681,N_14495,N_14453);
nor U14682 (N_14682,N_14444,N_14508);
xnor U14683 (N_14683,N_14415,N_14418);
xnor U14684 (N_14684,N_14541,N_14537);
xnor U14685 (N_14685,N_14440,N_14555);
or U14686 (N_14686,N_14511,N_14435);
xnor U14687 (N_14687,N_14467,N_14405);
xor U14688 (N_14688,N_14475,N_14412);
nor U14689 (N_14689,N_14495,N_14450);
or U14690 (N_14690,N_14430,N_14444);
xor U14691 (N_14691,N_14454,N_14474);
nor U14692 (N_14692,N_14452,N_14407);
nor U14693 (N_14693,N_14522,N_14414);
and U14694 (N_14694,N_14403,N_14428);
nor U14695 (N_14695,N_14531,N_14522);
or U14696 (N_14696,N_14541,N_14426);
or U14697 (N_14697,N_14461,N_14451);
or U14698 (N_14698,N_14515,N_14411);
and U14699 (N_14699,N_14415,N_14484);
nand U14700 (N_14700,N_14440,N_14409);
nor U14701 (N_14701,N_14485,N_14537);
nand U14702 (N_14702,N_14441,N_14431);
and U14703 (N_14703,N_14518,N_14549);
nand U14704 (N_14704,N_14549,N_14450);
nand U14705 (N_14705,N_14454,N_14487);
and U14706 (N_14706,N_14480,N_14541);
nand U14707 (N_14707,N_14423,N_14553);
or U14708 (N_14708,N_14447,N_14516);
and U14709 (N_14709,N_14544,N_14489);
or U14710 (N_14710,N_14428,N_14555);
nor U14711 (N_14711,N_14524,N_14441);
nor U14712 (N_14712,N_14443,N_14401);
and U14713 (N_14713,N_14467,N_14422);
xor U14714 (N_14714,N_14519,N_14438);
or U14715 (N_14715,N_14464,N_14433);
xor U14716 (N_14716,N_14550,N_14427);
xnor U14717 (N_14717,N_14474,N_14535);
or U14718 (N_14718,N_14533,N_14416);
or U14719 (N_14719,N_14510,N_14547);
nand U14720 (N_14720,N_14607,N_14567);
nor U14721 (N_14721,N_14584,N_14697);
xnor U14722 (N_14722,N_14678,N_14649);
or U14723 (N_14723,N_14666,N_14653);
nand U14724 (N_14724,N_14562,N_14589);
xor U14725 (N_14725,N_14673,N_14675);
and U14726 (N_14726,N_14591,N_14686);
nor U14727 (N_14727,N_14652,N_14705);
nor U14728 (N_14728,N_14648,N_14624);
and U14729 (N_14729,N_14651,N_14617);
or U14730 (N_14730,N_14590,N_14681);
nand U14731 (N_14731,N_14599,N_14560);
nor U14732 (N_14732,N_14667,N_14682);
xor U14733 (N_14733,N_14684,N_14677);
nand U14734 (N_14734,N_14632,N_14661);
nor U14735 (N_14735,N_14615,N_14602);
or U14736 (N_14736,N_14646,N_14610);
nand U14737 (N_14737,N_14644,N_14659);
nand U14738 (N_14738,N_14637,N_14628);
and U14739 (N_14739,N_14620,N_14575);
nand U14740 (N_14740,N_14596,N_14627);
nand U14741 (N_14741,N_14573,N_14647);
and U14742 (N_14742,N_14626,N_14657);
and U14743 (N_14743,N_14695,N_14709);
and U14744 (N_14744,N_14712,N_14664);
xor U14745 (N_14745,N_14604,N_14605);
or U14746 (N_14746,N_14708,N_14564);
and U14747 (N_14747,N_14582,N_14565);
and U14748 (N_14748,N_14656,N_14691);
nand U14749 (N_14749,N_14593,N_14635);
and U14750 (N_14750,N_14578,N_14702);
or U14751 (N_14751,N_14609,N_14690);
and U14752 (N_14752,N_14629,N_14685);
xnor U14753 (N_14753,N_14694,N_14561);
and U14754 (N_14754,N_14570,N_14600);
nand U14755 (N_14755,N_14580,N_14687);
nand U14756 (N_14756,N_14689,N_14710);
and U14757 (N_14757,N_14583,N_14704);
nor U14758 (N_14758,N_14700,N_14594);
and U14759 (N_14759,N_14699,N_14631);
nand U14760 (N_14760,N_14707,N_14608);
nor U14761 (N_14761,N_14693,N_14623);
nor U14762 (N_14762,N_14585,N_14668);
nand U14763 (N_14763,N_14574,N_14606);
or U14764 (N_14764,N_14641,N_14645);
nand U14765 (N_14765,N_14566,N_14670);
or U14766 (N_14766,N_14618,N_14718);
nor U14767 (N_14767,N_14688,N_14662);
and U14768 (N_14768,N_14569,N_14625);
nand U14769 (N_14769,N_14660,N_14692);
xor U14770 (N_14770,N_14633,N_14665);
nand U14771 (N_14771,N_14669,N_14683);
xor U14772 (N_14772,N_14579,N_14601);
nand U14773 (N_14773,N_14676,N_14576);
nor U14774 (N_14774,N_14577,N_14630);
xor U14775 (N_14775,N_14571,N_14701);
nor U14776 (N_14776,N_14655,N_14642);
nor U14777 (N_14777,N_14715,N_14614);
nand U14778 (N_14778,N_14696,N_14588);
nor U14779 (N_14779,N_14586,N_14612);
or U14780 (N_14780,N_14703,N_14658);
nand U14781 (N_14781,N_14597,N_14716);
and U14782 (N_14782,N_14711,N_14714);
xor U14783 (N_14783,N_14706,N_14572);
and U14784 (N_14784,N_14679,N_14671);
and U14785 (N_14785,N_14621,N_14680);
or U14786 (N_14786,N_14639,N_14650);
and U14787 (N_14787,N_14713,N_14643);
and U14788 (N_14788,N_14611,N_14595);
and U14789 (N_14789,N_14698,N_14619);
nand U14790 (N_14790,N_14563,N_14674);
nand U14791 (N_14791,N_14719,N_14603);
or U14792 (N_14792,N_14636,N_14634);
nor U14793 (N_14793,N_14581,N_14598);
nand U14794 (N_14794,N_14654,N_14638);
or U14795 (N_14795,N_14640,N_14616);
or U14796 (N_14796,N_14568,N_14622);
nor U14797 (N_14797,N_14672,N_14717);
nand U14798 (N_14798,N_14592,N_14613);
or U14799 (N_14799,N_14587,N_14663);
and U14800 (N_14800,N_14651,N_14672);
nor U14801 (N_14801,N_14715,N_14616);
xnor U14802 (N_14802,N_14622,N_14600);
or U14803 (N_14803,N_14715,N_14659);
or U14804 (N_14804,N_14620,N_14584);
or U14805 (N_14805,N_14716,N_14695);
or U14806 (N_14806,N_14610,N_14560);
nor U14807 (N_14807,N_14693,N_14589);
nor U14808 (N_14808,N_14698,N_14617);
or U14809 (N_14809,N_14670,N_14612);
nand U14810 (N_14810,N_14707,N_14648);
and U14811 (N_14811,N_14683,N_14568);
xor U14812 (N_14812,N_14603,N_14666);
xor U14813 (N_14813,N_14661,N_14633);
and U14814 (N_14814,N_14570,N_14677);
and U14815 (N_14815,N_14589,N_14584);
nand U14816 (N_14816,N_14640,N_14654);
xnor U14817 (N_14817,N_14686,N_14612);
nand U14818 (N_14818,N_14644,N_14668);
and U14819 (N_14819,N_14647,N_14570);
xor U14820 (N_14820,N_14639,N_14660);
and U14821 (N_14821,N_14652,N_14562);
or U14822 (N_14822,N_14648,N_14619);
xnor U14823 (N_14823,N_14645,N_14708);
nand U14824 (N_14824,N_14664,N_14611);
xor U14825 (N_14825,N_14643,N_14680);
nand U14826 (N_14826,N_14695,N_14569);
nor U14827 (N_14827,N_14712,N_14626);
nor U14828 (N_14828,N_14578,N_14670);
and U14829 (N_14829,N_14608,N_14610);
nor U14830 (N_14830,N_14578,N_14607);
or U14831 (N_14831,N_14628,N_14664);
xnor U14832 (N_14832,N_14628,N_14709);
nand U14833 (N_14833,N_14653,N_14607);
and U14834 (N_14834,N_14713,N_14586);
or U14835 (N_14835,N_14599,N_14593);
nor U14836 (N_14836,N_14696,N_14635);
and U14837 (N_14837,N_14697,N_14638);
xor U14838 (N_14838,N_14655,N_14678);
and U14839 (N_14839,N_14719,N_14624);
nor U14840 (N_14840,N_14708,N_14700);
xnor U14841 (N_14841,N_14715,N_14586);
or U14842 (N_14842,N_14715,N_14590);
or U14843 (N_14843,N_14616,N_14588);
xnor U14844 (N_14844,N_14648,N_14672);
or U14845 (N_14845,N_14646,N_14708);
nand U14846 (N_14846,N_14594,N_14628);
nand U14847 (N_14847,N_14649,N_14662);
and U14848 (N_14848,N_14625,N_14676);
or U14849 (N_14849,N_14642,N_14652);
nor U14850 (N_14850,N_14597,N_14648);
nand U14851 (N_14851,N_14670,N_14719);
nand U14852 (N_14852,N_14576,N_14595);
or U14853 (N_14853,N_14664,N_14601);
nor U14854 (N_14854,N_14670,N_14704);
nand U14855 (N_14855,N_14657,N_14584);
nor U14856 (N_14856,N_14647,N_14643);
and U14857 (N_14857,N_14619,N_14667);
nand U14858 (N_14858,N_14634,N_14598);
nor U14859 (N_14859,N_14676,N_14708);
nor U14860 (N_14860,N_14681,N_14663);
xnor U14861 (N_14861,N_14565,N_14661);
nor U14862 (N_14862,N_14673,N_14591);
nor U14863 (N_14863,N_14592,N_14652);
nor U14864 (N_14864,N_14605,N_14706);
nand U14865 (N_14865,N_14701,N_14695);
and U14866 (N_14866,N_14576,N_14579);
and U14867 (N_14867,N_14640,N_14576);
nor U14868 (N_14868,N_14656,N_14663);
or U14869 (N_14869,N_14604,N_14679);
nor U14870 (N_14870,N_14615,N_14578);
xor U14871 (N_14871,N_14621,N_14631);
nand U14872 (N_14872,N_14698,N_14682);
nor U14873 (N_14873,N_14643,N_14610);
nor U14874 (N_14874,N_14599,N_14681);
or U14875 (N_14875,N_14613,N_14713);
and U14876 (N_14876,N_14684,N_14716);
or U14877 (N_14877,N_14665,N_14657);
nor U14878 (N_14878,N_14576,N_14673);
nand U14879 (N_14879,N_14622,N_14703);
or U14880 (N_14880,N_14760,N_14731);
xor U14881 (N_14881,N_14860,N_14834);
or U14882 (N_14882,N_14761,N_14773);
or U14883 (N_14883,N_14783,N_14867);
xnor U14884 (N_14884,N_14824,N_14722);
xnor U14885 (N_14885,N_14791,N_14794);
nand U14886 (N_14886,N_14798,N_14819);
xor U14887 (N_14887,N_14725,N_14737);
and U14888 (N_14888,N_14822,N_14841);
or U14889 (N_14889,N_14818,N_14729);
and U14890 (N_14890,N_14821,N_14876);
and U14891 (N_14891,N_14872,N_14733);
or U14892 (N_14892,N_14865,N_14820);
nand U14893 (N_14893,N_14763,N_14800);
and U14894 (N_14894,N_14856,N_14752);
xnor U14895 (N_14895,N_14835,N_14804);
nor U14896 (N_14896,N_14764,N_14726);
xor U14897 (N_14897,N_14779,N_14817);
xor U14898 (N_14898,N_14793,N_14810);
or U14899 (N_14899,N_14740,N_14766);
nand U14900 (N_14900,N_14721,N_14812);
nand U14901 (N_14901,N_14836,N_14861);
and U14902 (N_14902,N_14744,N_14866);
nand U14903 (N_14903,N_14801,N_14723);
nor U14904 (N_14904,N_14772,N_14748);
xnor U14905 (N_14905,N_14862,N_14785);
nor U14906 (N_14906,N_14751,N_14728);
nand U14907 (N_14907,N_14879,N_14857);
and U14908 (N_14908,N_14853,N_14758);
nand U14909 (N_14909,N_14808,N_14738);
xnor U14910 (N_14910,N_14747,N_14803);
nor U14911 (N_14911,N_14849,N_14755);
xnor U14912 (N_14912,N_14765,N_14850);
nor U14913 (N_14913,N_14756,N_14805);
xor U14914 (N_14914,N_14734,N_14843);
nor U14915 (N_14915,N_14851,N_14769);
or U14916 (N_14916,N_14863,N_14746);
or U14917 (N_14917,N_14753,N_14855);
xor U14918 (N_14918,N_14739,N_14816);
and U14919 (N_14919,N_14781,N_14759);
xor U14920 (N_14920,N_14775,N_14724);
nor U14921 (N_14921,N_14839,N_14784);
nor U14922 (N_14922,N_14854,N_14768);
nor U14923 (N_14923,N_14829,N_14757);
and U14924 (N_14924,N_14869,N_14786);
nand U14925 (N_14925,N_14782,N_14811);
and U14926 (N_14926,N_14742,N_14833);
xor U14927 (N_14927,N_14868,N_14727);
xor U14928 (N_14928,N_14838,N_14845);
nand U14929 (N_14929,N_14846,N_14827);
or U14930 (N_14930,N_14825,N_14788);
nand U14931 (N_14931,N_14848,N_14802);
xor U14932 (N_14932,N_14875,N_14823);
nand U14933 (N_14933,N_14780,N_14807);
xnor U14934 (N_14934,N_14743,N_14736);
or U14935 (N_14935,N_14750,N_14815);
nor U14936 (N_14936,N_14795,N_14762);
or U14937 (N_14937,N_14813,N_14770);
nor U14938 (N_14938,N_14720,N_14789);
or U14939 (N_14939,N_14870,N_14877);
and U14940 (N_14940,N_14878,N_14797);
nand U14941 (N_14941,N_14826,N_14814);
and U14942 (N_14942,N_14837,N_14730);
or U14943 (N_14943,N_14792,N_14847);
or U14944 (N_14944,N_14874,N_14754);
xor U14945 (N_14945,N_14840,N_14828);
xnor U14946 (N_14946,N_14778,N_14796);
or U14947 (N_14947,N_14832,N_14809);
xor U14948 (N_14948,N_14830,N_14787);
and U14949 (N_14949,N_14771,N_14735);
and U14950 (N_14950,N_14776,N_14806);
or U14951 (N_14951,N_14831,N_14732);
xor U14952 (N_14952,N_14864,N_14777);
nand U14953 (N_14953,N_14858,N_14844);
or U14954 (N_14954,N_14741,N_14842);
or U14955 (N_14955,N_14871,N_14852);
or U14956 (N_14956,N_14790,N_14767);
xor U14957 (N_14957,N_14745,N_14873);
xor U14958 (N_14958,N_14774,N_14749);
xnor U14959 (N_14959,N_14799,N_14859);
and U14960 (N_14960,N_14779,N_14789);
xnor U14961 (N_14961,N_14813,N_14791);
and U14962 (N_14962,N_14843,N_14862);
nor U14963 (N_14963,N_14826,N_14834);
and U14964 (N_14964,N_14802,N_14834);
or U14965 (N_14965,N_14739,N_14722);
and U14966 (N_14966,N_14770,N_14872);
and U14967 (N_14967,N_14844,N_14854);
nor U14968 (N_14968,N_14744,N_14722);
nor U14969 (N_14969,N_14733,N_14720);
nand U14970 (N_14970,N_14790,N_14827);
or U14971 (N_14971,N_14870,N_14720);
or U14972 (N_14972,N_14840,N_14765);
and U14973 (N_14973,N_14862,N_14863);
nor U14974 (N_14974,N_14736,N_14798);
and U14975 (N_14975,N_14737,N_14745);
nand U14976 (N_14976,N_14870,N_14844);
nor U14977 (N_14977,N_14757,N_14749);
xor U14978 (N_14978,N_14774,N_14790);
xnor U14979 (N_14979,N_14837,N_14875);
nand U14980 (N_14980,N_14779,N_14788);
and U14981 (N_14981,N_14818,N_14870);
nand U14982 (N_14982,N_14874,N_14866);
nand U14983 (N_14983,N_14786,N_14730);
xnor U14984 (N_14984,N_14811,N_14804);
or U14985 (N_14985,N_14877,N_14803);
nand U14986 (N_14986,N_14851,N_14801);
and U14987 (N_14987,N_14798,N_14810);
or U14988 (N_14988,N_14755,N_14800);
nor U14989 (N_14989,N_14792,N_14835);
or U14990 (N_14990,N_14728,N_14752);
nand U14991 (N_14991,N_14784,N_14866);
and U14992 (N_14992,N_14801,N_14864);
nand U14993 (N_14993,N_14842,N_14771);
or U14994 (N_14994,N_14767,N_14789);
xnor U14995 (N_14995,N_14775,N_14762);
and U14996 (N_14996,N_14773,N_14816);
xor U14997 (N_14997,N_14831,N_14874);
nand U14998 (N_14998,N_14845,N_14812);
xnor U14999 (N_14999,N_14866,N_14815);
nor U15000 (N_15000,N_14850,N_14780);
xor U15001 (N_15001,N_14734,N_14748);
xnor U15002 (N_15002,N_14871,N_14773);
and U15003 (N_15003,N_14756,N_14819);
xor U15004 (N_15004,N_14733,N_14826);
or U15005 (N_15005,N_14781,N_14849);
or U15006 (N_15006,N_14851,N_14854);
nor U15007 (N_15007,N_14788,N_14781);
nand U15008 (N_15008,N_14747,N_14843);
nor U15009 (N_15009,N_14753,N_14822);
or U15010 (N_15010,N_14840,N_14767);
xnor U15011 (N_15011,N_14835,N_14860);
and U15012 (N_15012,N_14824,N_14814);
xor U15013 (N_15013,N_14790,N_14861);
or U15014 (N_15014,N_14771,N_14745);
xor U15015 (N_15015,N_14864,N_14840);
and U15016 (N_15016,N_14730,N_14825);
or U15017 (N_15017,N_14774,N_14778);
or U15018 (N_15018,N_14831,N_14748);
nand U15019 (N_15019,N_14762,N_14769);
and U15020 (N_15020,N_14746,N_14730);
nand U15021 (N_15021,N_14753,N_14795);
or U15022 (N_15022,N_14800,N_14858);
and U15023 (N_15023,N_14782,N_14758);
or U15024 (N_15024,N_14733,N_14827);
nand U15025 (N_15025,N_14732,N_14725);
xor U15026 (N_15026,N_14764,N_14834);
or U15027 (N_15027,N_14773,N_14786);
nor U15028 (N_15028,N_14863,N_14732);
nor U15029 (N_15029,N_14863,N_14872);
nor U15030 (N_15030,N_14833,N_14793);
nand U15031 (N_15031,N_14836,N_14850);
nor U15032 (N_15032,N_14865,N_14809);
xnor U15033 (N_15033,N_14875,N_14860);
and U15034 (N_15034,N_14742,N_14841);
or U15035 (N_15035,N_14776,N_14781);
or U15036 (N_15036,N_14768,N_14839);
or U15037 (N_15037,N_14854,N_14777);
xnor U15038 (N_15038,N_14721,N_14773);
or U15039 (N_15039,N_14826,N_14825);
or U15040 (N_15040,N_14968,N_14917);
and U15041 (N_15041,N_14976,N_14962);
nor U15042 (N_15042,N_15024,N_14926);
or U15043 (N_15043,N_14920,N_14937);
xor U15044 (N_15044,N_14965,N_15009);
nor U15045 (N_15045,N_14948,N_14933);
xor U15046 (N_15046,N_15012,N_15005);
nor U15047 (N_15047,N_14930,N_14996);
or U15048 (N_15048,N_15032,N_15002);
and U15049 (N_15049,N_14922,N_14901);
nand U15050 (N_15050,N_14942,N_14974);
nand U15051 (N_15051,N_14950,N_15021);
nand U15052 (N_15052,N_15000,N_15025);
or U15053 (N_15053,N_14961,N_14889);
and U15054 (N_15054,N_14985,N_15038);
and U15055 (N_15055,N_14987,N_14909);
nand U15056 (N_15056,N_14929,N_14888);
nand U15057 (N_15057,N_14893,N_14954);
xor U15058 (N_15058,N_15010,N_14891);
and U15059 (N_15059,N_15035,N_15022);
or U15060 (N_15060,N_14898,N_14881);
or U15061 (N_15061,N_15014,N_14927);
nor U15062 (N_15062,N_14936,N_14964);
nor U15063 (N_15063,N_14931,N_14986);
and U15064 (N_15064,N_14955,N_15036);
nor U15065 (N_15065,N_14975,N_15006);
and U15066 (N_15066,N_14886,N_15020);
xnor U15067 (N_15067,N_14945,N_14953);
and U15068 (N_15068,N_15030,N_14949);
and U15069 (N_15069,N_14957,N_14910);
nand U15070 (N_15070,N_14912,N_14978);
or U15071 (N_15071,N_14916,N_14982);
nand U15072 (N_15072,N_14915,N_14963);
or U15073 (N_15073,N_14947,N_14967);
nand U15074 (N_15074,N_15023,N_15019);
nand U15075 (N_15075,N_14972,N_14983);
nor U15076 (N_15076,N_14921,N_14984);
xnor U15077 (N_15077,N_15011,N_14977);
nand U15078 (N_15078,N_15017,N_14896);
nand U15079 (N_15079,N_14911,N_14993);
nand U15080 (N_15080,N_14992,N_14995);
nor U15081 (N_15081,N_14928,N_15007);
and U15082 (N_15082,N_15015,N_14900);
nand U15083 (N_15083,N_14918,N_14880);
and U15084 (N_15084,N_14895,N_14994);
or U15085 (N_15085,N_15031,N_14894);
nor U15086 (N_15086,N_14956,N_14907);
and U15087 (N_15087,N_15013,N_15037);
and U15088 (N_15088,N_14960,N_14946);
or U15089 (N_15089,N_14914,N_14980);
and U15090 (N_15090,N_14932,N_14951);
and U15091 (N_15091,N_14944,N_14905);
and U15092 (N_15092,N_14925,N_14885);
or U15093 (N_15093,N_14902,N_14882);
nor U15094 (N_15094,N_14981,N_14940);
nand U15095 (N_15095,N_14919,N_14899);
and U15096 (N_15096,N_14908,N_14969);
nor U15097 (N_15097,N_15039,N_14913);
nor U15098 (N_15098,N_14924,N_14939);
and U15099 (N_15099,N_14952,N_15008);
nor U15100 (N_15100,N_14959,N_15034);
nand U15101 (N_15101,N_14884,N_14999);
and U15102 (N_15102,N_15029,N_14890);
or U15103 (N_15103,N_14989,N_14892);
nor U15104 (N_15104,N_14887,N_14904);
or U15105 (N_15105,N_14943,N_14970);
nor U15106 (N_15106,N_15001,N_14935);
xor U15107 (N_15107,N_14938,N_15004);
xnor U15108 (N_15108,N_14988,N_14973);
or U15109 (N_15109,N_15003,N_14897);
and U15110 (N_15110,N_15018,N_15028);
or U15111 (N_15111,N_14966,N_15027);
or U15112 (N_15112,N_14991,N_14923);
nand U15113 (N_15113,N_14958,N_14990);
nor U15114 (N_15114,N_14997,N_14979);
nand U15115 (N_15115,N_14941,N_14903);
nor U15116 (N_15116,N_14971,N_15026);
xor U15117 (N_15117,N_14883,N_15033);
nand U15118 (N_15118,N_14906,N_14934);
and U15119 (N_15119,N_14998,N_15016);
or U15120 (N_15120,N_14934,N_14976);
and U15121 (N_15121,N_14933,N_14908);
and U15122 (N_15122,N_14938,N_14903);
nand U15123 (N_15123,N_15029,N_14967);
or U15124 (N_15124,N_14952,N_14963);
nor U15125 (N_15125,N_14890,N_14909);
or U15126 (N_15126,N_14917,N_14940);
nor U15127 (N_15127,N_14907,N_14979);
nand U15128 (N_15128,N_14917,N_14989);
nand U15129 (N_15129,N_14942,N_14933);
xor U15130 (N_15130,N_14979,N_14983);
nor U15131 (N_15131,N_15012,N_14973);
nor U15132 (N_15132,N_15017,N_14882);
or U15133 (N_15133,N_15033,N_14981);
and U15134 (N_15134,N_14993,N_14984);
nand U15135 (N_15135,N_14983,N_14962);
and U15136 (N_15136,N_14983,N_14899);
xnor U15137 (N_15137,N_14898,N_14910);
nor U15138 (N_15138,N_15025,N_15002);
xnor U15139 (N_15139,N_14964,N_14914);
or U15140 (N_15140,N_15034,N_15023);
xnor U15141 (N_15141,N_14992,N_14883);
nor U15142 (N_15142,N_14989,N_14997);
nor U15143 (N_15143,N_14897,N_14886);
nand U15144 (N_15144,N_15004,N_14983);
and U15145 (N_15145,N_14993,N_14977);
xor U15146 (N_15146,N_14969,N_14989);
or U15147 (N_15147,N_14990,N_15019);
nand U15148 (N_15148,N_14990,N_14911);
and U15149 (N_15149,N_14919,N_15022);
nand U15150 (N_15150,N_14905,N_14949);
nor U15151 (N_15151,N_14945,N_14928);
and U15152 (N_15152,N_15037,N_14953);
and U15153 (N_15153,N_14976,N_15025);
and U15154 (N_15154,N_14922,N_15001);
nor U15155 (N_15155,N_15020,N_14889);
nor U15156 (N_15156,N_14979,N_14998);
nand U15157 (N_15157,N_15023,N_14982);
nand U15158 (N_15158,N_14939,N_15024);
nand U15159 (N_15159,N_14977,N_14943);
nor U15160 (N_15160,N_15039,N_14902);
nor U15161 (N_15161,N_14915,N_14945);
xor U15162 (N_15162,N_14930,N_14946);
and U15163 (N_15163,N_14886,N_15010);
xnor U15164 (N_15164,N_14972,N_14955);
or U15165 (N_15165,N_14909,N_14945);
and U15166 (N_15166,N_15014,N_15031);
nor U15167 (N_15167,N_14897,N_14916);
nand U15168 (N_15168,N_14891,N_15004);
nor U15169 (N_15169,N_15002,N_14905);
nor U15170 (N_15170,N_14950,N_14889);
or U15171 (N_15171,N_15028,N_15001);
or U15172 (N_15172,N_14955,N_14977);
and U15173 (N_15173,N_14881,N_14937);
nand U15174 (N_15174,N_15008,N_14926);
and U15175 (N_15175,N_14949,N_15008);
nor U15176 (N_15176,N_14933,N_15036);
or U15177 (N_15177,N_14998,N_14914);
xnor U15178 (N_15178,N_14986,N_14885);
and U15179 (N_15179,N_14924,N_14970);
nor U15180 (N_15180,N_15007,N_15004);
and U15181 (N_15181,N_14965,N_15025);
nor U15182 (N_15182,N_14891,N_14998);
xnor U15183 (N_15183,N_14917,N_14910);
and U15184 (N_15184,N_14966,N_14997);
and U15185 (N_15185,N_14988,N_14979);
xnor U15186 (N_15186,N_14958,N_14892);
or U15187 (N_15187,N_15005,N_15038);
or U15188 (N_15188,N_15009,N_15016);
and U15189 (N_15189,N_14991,N_15033);
nor U15190 (N_15190,N_14940,N_14890);
nand U15191 (N_15191,N_15032,N_14904);
nor U15192 (N_15192,N_14892,N_14904);
or U15193 (N_15193,N_14901,N_14965);
nor U15194 (N_15194,N_14939,N_15004);
or U15195 (N_15195,N_15023,N_14927);
or U15196 (N_15196,N_14916,N_14969);
or U15197 (N_15197,N_14986,N_14922);
and U15198 (N_15198,N_14972,N_15001);
xor U15199 (N_15199,N_14898,N_14939);
or U15200 (N_15200,N_15045,N_15131);
or U15201 (N_15201,N_15089,N_15125);
nand U15202 (N_15202,N_15063,N_15123);
and U15203 (N_15203,N_15145,N_15062);
and U15204 (N_15204,N_15106,N_15064);
or U15205 (N_15205,N_15116,N_15159);
nor U15206 (N_15206,N_15068,N_15076);
xnor U15207 (N_15207,N_15170,N_15110);
xnor U15208 (N_15208,N_15071,N_15185);
nand U15209 (N_15209,N_15085,N_15065);
and U15210 (N_15210,N_15138,N_15048);
xor U15211 (N_15211,N_15199,N_15186);
nor U15212 (N_15212,N_15053,N_15134);
nand U15213 (N_15213,N_15103,N_15080);
xnor U15214 (N_15214,N_15121,N_15152);
xnor U15215 (N_15215,N_15174,N_15178);
xor U15216 (N_15216,N_15099,N_15165);
and U15217 (N_15217,N_15082,N_15043);
nor U15218 (N_15218,N_15059,N_15177);
xor U15219 (N_15219,N_15070,N_15191);
or U15220 (N_15220,N_15135,N_15166);
and U15221 (N_15221,N_15057,N_15126);
and U15222 (N_15222,N_15194,N_15179);
and U15223 (N_15223,N_15074,N_15142);
nand U15224 (N_15224,N_15197,N_15148);
nand U15225 (N_15225,N_15051,N_15127);
or U15226 (N_15226,N_15144,N_15146);
and U15227 (N_15227,N_15184,N_15078);
xnor U15228 (N_15228,N_15181,N_15128);
xnor U15229 (N_15229,N_15073,N_15122);
nor U15230 (N_15230,N_15111,N_15072);
or U15231 (N_15231,N_15081,N_15094);
or U15232 (N_15232,N_15050,N_15167);
nand U15233 (N_15233,N_15158,N_15092);
nand U15234 (N_15234,N_15155,N_15056);
xnor U15235 (N_15235,N_15100,N_15173);
nand U15236 (N_15236,N_15147,N_15150);
nand U15237 (N_15237,N_15151,N_15115);
or U15238 (N_15238,N_15187,N_15091);
or U15239 (N_15239,N_15108,N_15084);
and U15240 (N_15240,N_15182,N_15118);
or U15241 (N_15241,N_15044,N_15069);
nor U15242 (N_15242,N_15183,N_15101);
xnor U15243 (N_15243,N_15086,N_15054);
nand U15244 (N_15244,N_15157,N_15117);
and U15245 (N_15245,N_15052,N_15124);
or U15246 (N_15246,N_15090,N_15162);
or U15247 (N_15247,N_15047,N_15176);
and U15248 (N_15248,N_15061,N_15175);
and U15249 (N_15249,N_15049,N_15098);
xnor U15250 (N_15250,N_15113,N_15107);
xnor U15251 (N_15251,N_15196,N_15190);
nand U15252 (N_15252,N_15041,N_15193);
xor U15253 (N_15253,N_15163,N_15087);
and U15254 (N_15254,N_15171,N_15130);
nand U15255 (N_15255,N_15133,N_15060);
or U15256 (N_15256,N_15189,N_15067);
nor U15257 (N_15257,N_15172,N_15156);
nor U15258 (N_15258,N_15169,N_15161);
nor U15259 (N_15259,N_15079,N_15046);
and U15260 (N_15260,N_15129,N_15096);
nor U15261 (N_15261,N_15137,N_15164);
nand U15262 (N_15262,N_15136,N_15192);
or U15263 (N_15263,N_15109,N_15083);
xnor U15264 (N_15264,N_15195,N_15102);
nor U15265 (N_15265,N_15119,N_15153);
nor U15266 (N_15266,N_15058,N_15143);
nand U15267 (N_15267,N_15055,N_15141);
nand U15268 (N_15268,N_15168,N_15088);
or U15269 (N_15269,N_15077,N_15112);
xor U15270 (N_15270,N_15075,N_15093);
and U15271 (N_15271,N_15042,N_15095);
nor U15272 (N_15272,N_15120,N_15188);
or U15273 (N_15273,N_15154,N_15140);
nor U15274 (N_15274,N_15097,N_15114);
or U15275 (N_15275,N_15149,N_15160);
nor U15276 (N_15276,N_15180,N_15132);
xnor U15277 (N_15277,N_15066,N_15198);
nor U15278 (N_15278,N_15105,N_15104);
nand U15279 (N_15279,N_15139,N_15040);
nand U15280 (N_15280,N_15162,N_15193);
nor U15281 (N_15281,N_15095,N_15105);
nor U15282 (N_15282,N_15076,N_15070);
or U15283 (N_15283,N_15096,N_15040);
or U15284 (N_15284,N_15129,N_15188);
nor U15285 (N_15285,N_15086,N_15166);
nand U15286 (N_15286,N_15158,N_15090);
nand U15287 (N_15287,N_15072,N_15086);
and U15288 (N_15288,N_15194,N_15067);
xnor U15289 (N_15289,N_15067,N_15103);
and U15290 (N_15290,N_15119,N_15090);
nand U15291 (N_15291,N_15186,N_15059);
nor U15292 (N_15292,N_15147,N_15091);
nor U15293 (N_15293,N_15049,N_15181);
or U15294 (N_15294,N_15097,N_15152);
and U15295 (N_15295,N_15148,N_15060);
nand U15296 (N_15296,N_15180,N_15117);
nand U15297 (N_15297,N_15048,N_15061);
nor U15298 (N_15298,N_15160,N_15098);
or U15299 (N_15299,N_15091,N_15094);
and U15300 (N_15300,N_15076,N_15100);
nand U15301 (N_15301,N_15086,N_15160);
nor U15302 (N_15302,N_15162,N_15083);
nor U15303 (N_15303,N_15094,N_15171);
or U15304 (N_15304,N_15093,N_15165);
xor U15305 (N_15305,N_15063,N_15066);
or U15306 (N_15306,N_15130,N_15094);
nand U15307 (N_15307,N_15079,N_15129);
nand U15308 (N_15308,N_15118,N_15059);
nor U15309 (N_15309,N_15109,N_15080);
and U15310 (N_15310,N_15145,N_15174);
or U15311 (N_15311,N_15140,N_15118);
nor U15312 (N_15312,N_15064,N_15117);
or U15313 (N_15313,N_15057,N_15146);
or U15314 (N_15314,N_15103,N_15041);
nor U15315 (N_15315,N_15098,N_15040);
and U15316 (N_15316,N_15071,N_15152);
nor U15317 (N_15317,N_15089,N_15120);
nor U15318 (N_15318,N_15074,N_15105);
xor U15319 (N_15319,N_15197,N_15168);
and U15320 (N_15320,N_15126,N_15079);
nand U15321 (N_15321,N_15041,N_15118);
and U15322 (N_15322,N_15091,N_15104);
and U15323 (N_15323,N_15124,N_15126);
and U15324 (N_15324,N_15185,N_15091);
or U15325 (N_15325,N_15144,N_15071);
xnor U15326 (N_15326,N_15099,N_15116);
xor U15327 (N_15327,N_15093,N_15049);
xor U15328 (N_15328,N_15187,N_15189);
and U15329 (N_15329,N_15158,N_15131);
or U15330 (N_15330,N_15185,N_15137);
and U15331 (N_15331,N_15096,N_15082);
nand U15332 (N_15332,N_15137,N_15178);
or U15333 (N_15333,N_15060,N_15166);
and U15334 (N_15334,N_15088,N_15173);
xnor U15335 (N_15335,N_15152,N_15187);
nand U15336 (N_15336,N_15111,N_15177);
nand U15337 (N_15337,N_15048,N_15057);
or U15338 (N_15338,N_15180,N_15126);
xnor U15339 (N_15339,N_15065,N_15190);
nand U15340 (N_15340,N_15056,N_15184);
and U15341 (N_15341,N_15182,N_15107);
nor U15342 (N_15342,N_15187,N_15051);
nand U15343 (N_15343,N_15087,N_15134);
or U15344 (N_15344,N_15058,N_15152);
nor U15345 (N_15345,N_15044,N_15061);
or U15346 (N_15346,N_15184,N_15195);
nor U15347 (N_15347,N_15067,N_15111);
nor U15348 (N_15348,N_15073,N_15176);
nor U15349 (N_15349,N_15098,N_15183);
nand U15350 (N_15350,N_15044,N_15068);
xor U15351 (N_15351,N_15133,N_15153);
nor U15352 (N_15352,N_15145,N_15164);
and U15353 (N_15353,N_15123,N_15155);
nand U15354 (N_15354,N_15142,N_15182);
and U15355 (N_15355,N_15153,N_15162);
nand U15356 (N_15356,N_15138,N_15055);
nor U15357 (N_15357,N_15182,N_15131);
nand U15358 (N_15358,N_15061,N_15049);
xnor U15359 (N_15359,N_15140,N_15161);
nand U15360 (N_15360,N_15245,N_15220);
or U15361 (N_15361,N_15352,N_15259);
nand U15362 (N_15362,N_15200,N_15243);
nand U15363 (N_15363,N_15276,N_15298);
or U15364 (N_15364,N_15270,N_15279);
nor U15365 (N_15365,N_15254,N_15321);
and U15366 (N_15366,N_15231,N_15212);
and U15367 (N_15367,N_15335,N_15304);
and U15368 (N_15368,N_15219,N_15296);
or U15369 (N_15369,N_15286,N_15206);
and U15370 (N_15370,N_15271,N_15244);
and U15371 (N_15371,N_15232,N_15263);
nand U15372 (N_15372,N_15309,N_15305);
xor U15373 (N_15373,N_15295,N_15236);
nor U15374 (N_15374,N_15273,N_15327);
nor U15375 (N_15375,N_15234,N_15233);
nor U15376 (N_15376,N_15247,N_15238);
nand U15377 (N_15377,N_15275,N_15357);
nand U15378 (N_15378,N_15336,N_15297);
nand U15379 (N_15379,N_15223,N_15339);
xnor U15380 (N_15380,N_15340,N_15218);
xor U15381 (N_15381,N_15307,N_15319);
xnor U15382 (N_15382,N_15288,N_15282);
or U15383 (N_15383,N_15242,N_15338);
nand U15384 (N_15384,N_15353,N_15253);
xnor U15385 (N_15385,N_15355,N_15255);
xor U15386 (N_15386,N_15303,N_15269);
xnor U15387 (N_15387,N_15333,N_15264);
nor U15388 (N_15388,N_15207,N_15331);
or U15389 (N_15389,N_15344,N_15274);
xor U15390 (N_15390,N_15235,N_15320);
and U15391 (N_15391,N_15241,N_15334);
xnor U15392 (N_15392,N_15287,N_15211);
or U15393 (N_15393,N_15332,N_15323);
and U15394 (N_15394,N_15248,N_15289);
or U15395 (N_15395,N_15329,N_15285);
xor U15396 (N_15396,N_15291,N_15315);
or U15397 (N_15397,N_15227,N_15308);
and U15398 (N_15398,N_15330,N_15351);
nand U15399 (N_15399,N_15251,N_15358);
and U15400 (N_15400,N_15209,N_15312);
nor U15401 (N_15401,N_15267,N_15346);
xnor U15402 (N_15402,N_15350,N_15348);
nor U15403 (N_15403,N_15301,N_15283);
xnor U15404 (N_15404,N_15237,N_15222);
or U15405 (N_15405,N_15356,N_15208);
nand U15406 (N_15406,N_15210,N_15202);
nand U15407 (N_15407,N_15224,N_15326);
xor U15408 (N_15408,N_15203,N_15225);
nand U15409 (N_15409,N_15205,N_15316);
or U15410 (N_15410,N_15300,N_15325);
nand U15411 (N_15411,N_15347,N_15354);
xor U15412 (N_15412,N_15239,N_15221);
xnor U15413 (N_15413,N_15215,N_15328);
or U15414 (N_15414,N_15250,N_15260);
xnor U15415 (N_15415,N_15256,N_15280);
xor U15416 (N_15416,N_15306,N_15246);
nand U15417 (N_15417,N_15324,N_15204);
and U15418 (N_15418,N_15349,N_15302);
or U15419 (N_15419,N_15217,N_15201);
xor U15420 (N_15420,N_15213,N_15314);
nor U15421 (N_15421,N_15226,N_15261);
or U15422 (N_15422,N_15281,N_15277);
nor U15423 (N_15423,N_15266,N_15284);
and U15424 (N_15424,N_15252,N_15341);
and U15425 (N_15425,N_15268,N_15342);
xor U15426 (N_15426,N_15337,N_15292);
or U15427 (N_15427,N_15311,N_15228);
and U15428 (N_15428,N_15240,N_15216);
nand U15429 (N_15429,N_15230,N_15249);
and U15430 (N_15430,N_15214,N_15262);
or U15431 (N_15431,N_15265,N_15258);
and U15432 (N_15432,N_15317,N_15310);
nor U15433 (N_15433,N_15299,N_15272);
nor U15434 (N_15434,N_15322,N_15294);
nand U15435 (N_15435,N_15345,N_15278);
and U15436 (N_15436,N_15229,N_15313);
xnor U15437 (N_15437,N_15257,N_15318);
nor U15438 (N_15438,N_15343,N_15359);
or U15439 (N_15439,N_15293,N_15290);
nand U15440 (N_15440,N_15216,N_15277);
and U15441 (N_15441,N_15304,N_15353);
or U15442 (N_15442,N_15258,N_15241);
or U15443 (N_15443,N_15241,N_15326);
and U15444 (N_15444,N_15264,N_15244);
nand U15445 (N_15445,N_15252,N_15307);
xnor U15446 (N_15446,N_15210,N_15344);
or U15447 (N_15447,N_15293,N_15235);
and U15448 (N_15448,N_15326,N_15252);
and U15449 (N_15449,N_15227,N_15234);
and U15450 (N_15450,N_15230,N_15234);
and U15451 (N_15451,N_15334,N_15236);
or U15452 (N_15452,N_15247,N_15308);
xnor U15453 (N_15453,N_15330,N_15340);
nor U15454 (N_15454,N_15219,N_15258);
xnor U15455 (N_15455,N_15286,N_15257);
nand U15456 (N_15456,N_15327,N_15255);
and U15457 (N_15457,N_15315,N_15323);
xor U15458 (N_15458,N_15315,N_15215);
nor U15459 (N_15459,N_15356,N_15214);
nor U15460 (N_15460,N_15204,N_15310);
nand U15461 (N_15461,N_15261,N_15278);
or U15462 (N_15462,N_15249,N_15318);
or U15463 (N_15463,N_15351,N_15333);
or U15464 (N_15464,N_15209,N_15235);
nor U15465 (N_15465,N_15292,N_15211);
xor U15466 (N_15466,N_15352,N_15246);
and U15467 (N_15467,N_15250,N_15218);
nor U15468 (N_15468,N_15238,N_15276);
or U15469 (N_15469,N_15266,N_15327);
xor U15470 (N_15470,N_15236,N_15328);
xnor U15471 (N_15471,N_15282,N_15250);
and U15472 (N_15472,N_15255,N_15285);
xnor U15473 (N_15473,N_15297,N_15204);
nor U15474 (N_15474,N_15303,N_15297);
xnor U15475 (N_15475,N_15267,N_15303);
or U15476 (N_15476,N_15343,N_15354);
xnor U15477 (N_15477,N_15308,N_15337);
xor U15478 (N_15478,N_15253,N_15340);
nor U15479 (N_15479,N_15265,N_15346);
nand U15480 (N_15480,N_15246,N_15283);
xnor U15481 (N_15481,N_15207,N_15288);
nor U15482 (N_15482,N_15356,N_15266);
and U15483 (N_15483,N_15275,N_15208);
xnor U15484 (N_15484,N_15280,N_15340);
nor U15485 (N_15485,N_15344,N_15200);
xor U15486 (N_15486,N_15339,N_15287);
or U15487 (N_15487,N_15344,N_15245);
nand U15488 (N_15488,N_15244,N_15222);
nand U15489 (N_15489,N_15249,N_15342);
xnor U15490 (N_15490,N_15354,N_15234);
or U15491 (N_15491,N_15338,N_15332);
nor U15492 (N_15492,N_15219,N_15285);
nand U15493 (N_15493,N_15301,N_15322);
and U15494 (N_15494,N_15291,N_15264);
xor U15495 (N_15495,N_15213,N_15231);
nor U15496 (N_15496,N_15284,N_15322);
or U15497 (N_15497,N_15316,N_15245);
nand U15498 (N_15498,N_15297,N_15258);
or U15499 (N_15499,N_15302,N_15221);
nor U15500 (N_15500,N_15342,N_15325);
and U15501 (N_15501,N_15318,N_15215);
nand U15502 (N_15502,N_15224,N_15277);
nand U15503 (N_15503,N_15315,N_15210);
or U15504 (N_15504,N_15241,N_15344);
nand U15505 (N_15505,N_15258,N_15337);
or U15506 (N_15506,N_15247,N_15299);
nor U15507 (N_15507,N_15331,N_15218);
and U15508 (N_15508,N_15220,N_15321);
and U15509 (N_15509,N_15267,N_15277);
nor U15510 (N_15510,N_15323,N_15290);
xnor U15511 (N_15511,N_15236,N_15319);
nand U15512 (N_15512,N_15262,N_15240);
and U15513 (N_15513,N_15297,N_15228);
nor U15514 (N_15514,N_15348,N_15221);
or U15515 (N_15515,N_15327,N_15252);
nand U15516 (N_15516,N_15236,N_15255);
xnor U15517 (N_15517,N_15239,N_15323);
or U15518 (N_15518,N_15342,N_15218);
and U15519 (N_15519,N_15265,N_15243);
or U15520 (N_15520,N_15478,N_15434);
and U15521 (N_15521,N_15377,N_15458);
nand U15522 (N_15522,N_15512,N_15486);
or U15523 (N_15523,N_15474,N_15495);
and U15524 (N_15524,N_15461,N_15380);
nand U15525 (N_15525,N_15439,N_15360);
nand U15526 (N_15526,N_15504,N_15488);
nor U15527 (N_15527,N_15436,N_15418);
and U15528 (N_15528,N_15484,N_15515);
nand U15529 (N_15529,N_15361,N_15496);
and U15530 (N_15530,N_15501,N_15410);
and U15531 (N_15531,N_15468,N_15456);
and U15532 (N_15532,N_15422,N_15362);
nand U15533 (N_15533,N_15369,N_15384);
and U15534 (N_15534,N_15457,N_15412);
nand U15535 (N_15535,N_15413,N_15498);
nor U15536 (N_15536,N_15453,N_15397);
nor U15537 (N_15537,N_15414,N_15404);
nor U15538 (N_15538,N_15394,N_15409);
xor U15539 (N_15539,N_15416,N_15455);
nand U15540 (N_15540,N_15438,N_15464);
xor U15541 (N_15541,N_15403,N_15463);
xnor U15542 (N_15542,N_15406,N_15367);
and U15543 (N_15543,N_15505,N_15450);
nand U15544 (N_15544,N_15408,N_15502);
nor U15545 (N_15545,N_15480,N_15451);
nor U15546 (N_15546,N_15402,N_15460);
nand U15547 (N_15547,N_15473,N_15385);
and U15548 (N_15548,N_15508,N_15363);
nor U15549 (N_15549,N_15419,N_15382);
or U15550 (N_15550,N_15469,N_15395);
nor U15551 (N_15551,N_15454,N_15424);
or U15552 (N_15552,N_15481,N_15411);
xor U15553 (N_15553,N_15388,N_15491);
nor U15554 (N_15554,N_15400,N_15396);
and U15555 (N_15555,N_15373,N_15368);
or U15556 (N_15556,N_15393,N_15381);
or U15557 (N_15557,N_15421,N_15429);
xor U15558 (N_15558,N_15433,N_15405);
xnor U15559 (N_15559,N_15392,N_15516);
nor U15560 (N_15560,N_15383,N_15482);
xnor U15561 (N_15561,N_15445,N_15499);
and U15562 (N_15562,N_15378,N_15446);
xor U15563 (N_15563,N_15447,N_15431);
nand U15564 (N_15564,N_15374,N_15466);
xnor U15565 (N_15565,N_15441,N_15494);
xor U15566 (N_15566,N_15449,N_15376);
xor U15567 (N_15567,N_15513,N_15430);
xor U15568 (N_15568,N_15500,N_15389);
nor U15569 (N_15569,N_15391,N_15475);
nor U15570 (N_15570,N_15379,N_15426);
nand U15571 (N_15571,N_15372,N_15398);
nand U15572 (N_15572,N_15489,N_15479);
xnor U15573 (N_15573,N_15470,N_15443);
nor U15574 (N_15574,N_15514,N_15448);
xnor U15575 (N_15575,N_15437,N_15401);
nand U15576 (N_15576,N_15407,N_15497);
nand U15577 (N_15577,N_15390,N_15440);
and U15578 (N_15578,N_15365,N_15428);
xor U15579 (N_15579,N_15427,N_15425);
nand U15580 (N_15580,N_15477,N_15487);
or U15581 (N_15581,N_15517,N_15510);
nor U15582 (N_15582,N_15492,N_15518);
or U15583 (N_15583,N_15509,N_15476);
xnor U15584 (N_15584,N_15386,N_15371);
nor U15585 (N_15585,N_15485,N_15444);
nand U15586 (N_15586,N_15506,N_15370);
or U15587 (N_15587,N_15507,N_15471);
and U15588 (N_15588,N_15462,N_15465);
nor U15589 (N_15589,N_15493,N_15387);
nand U15590 (N_15590,N_15399,N_15503);
and U15591 (N_15591,N_15415,N_15366);
nand U15592 (N_15592,N_15364,N_15483);
nand U15593 (N_15593,N_15423,N_15511);
or U15594 (N_15594,N_15490,N_15459);
or U15595 (N_15595,N_15467,N_15435);
xor U15596 (N_15596,N_15375,N_15519);
xnor U15597 (N_15597,N_15432,N_15417);
xor U15598 (N_15598,N_15442,N_15452);
nor U15599 (N_15599,N_15472,N_15420);
or U15600 (N_15600,N_15376,N_15506);
nand U15601 (N_15601,N_15387,N_15460);
or U15602 (N_15602,N_15445,N_15485);
xnor U15603 (N_15603,N_15396,N_15429);
nand U15604 (N_15604,N_15427,N_15368);
or U15605 (N_15605,N_15429,N_15493);
and U15606 (N_15606,N_15441,N_15408);
xnor U15607 (N_15607,N_15393,N_15452);
nand U15608 (N_15608,N_15469,N_15413);
nand U15609 (N_15609,N_15393,N_15428);
xnor U15610 (N_15610,N_15429,N_15389);
xnor U15611 (N_15611,N_15441,N_15403);
and U15612 (N_15612,N_15463,N_15437);
nand U15613 (N_15613,N_15368,N_15508);
xor U15614 (N_15614,N_15360,N_15412);
and U15615 (N_15615,N_15366,N_15452);
and U15616 (N_15616,N_15394,N_15433);
nand U15617 (N_15617,N_15498,N_15407);
nor U15618 (N_15618,N_15456,N_15518);
or U15619 (N_15619,N_15495,N_15466);
and U15620 (N_15620,N_15453,N_15364);
nand U15621 (N_15621,N_15386,N_15410);
and U15622 (N_15622,N_15455,N_15465);
and U15623 (N_15623,N_15518,N_15471);
nand U15624 (N_15624,N_15371,N_15388);
nor U15625 (N_15625,N_15410,N_15400);
or U15626 (N_15626,N_15447,N_15506);
xor U15627 (N_15627,N_15487,N_15510);
nor U15628 (N_15628,N_15414,N_15451);
and U15629 (N_15629,N_15400,N_15518);
nor U15630 (N_15630,N_15418,N_15362);
nand U15631 (N_15631,N_15406,N_15438);
nor U15632 (N_15632,N_15444,N_15511);
nor U15633 (N_15633,N_15418,N_15415);
nor U15634 (N_15634,N_15460,N_15422);
nand U15635 (N_15635,N_15416,N_15445);
or U15636 (N_15636,N_15388,N_15365);
nand U15637 (N_15637,N_15430,N_15421);
nand U15638 (N_15638,N_15488,N_15453);
nor U15639 (N_15639,N_15452,N_15518);
xor U15640 (N_15640,N_15450,N_15515);
and U15641 (N_15641,N_15439,N_15465);
nor U15642 (N_15642,N_15445,N_15366);
xor U15643 (N_15643,N_15363,N_15362);
nor U15644 (N_15644,N_15460,N_15443);
xnor U15645 (N_15645,N_15364,N_15425);
or U15646 (N_15646,N_15503,N_15462);
or U15647 (N_15647,N_15478,N_15444);
or U15648 (N_15648,N_15512,N_15515);
and U15649 (N_15649,N_15514,N_15439);
and U15650 (N_15650,N_15381,N_15476);
xor U15651 (N_15651,N_15389,N_15408);
nor U15652 (N_15652,N_15393,N_15385);
or U15653 (N_15653,N_15514,N_15404);
and U15654 (N_15654,N_15393,N_15371);
or U15655 (N_15655,N_15464,N_15448);
or U15656 (N_15656,N_15498,N_15446);
nand U15657 (N_15657,N_15510,N_15374);
nor U15658 (N_15658,N_15437,N_15486);
nor U15659 (N_15659,N_15442,N_15478);
nor U15660 (N_15660,N_15370,N_15415);
xor U15661 (N_15661,N_15465,N_15406);
and U15662 (N_15662,N_15498,N_15372);
or U15663 (N_15663,N_15476,N_15411);
xor U15664 (N_15664,N_15426,N_15479);
nand U15665 (N_15665,N_15377,N_15370);
xor U15666 (N_15666,N_15465,N_15512);
or U15667 (N_15667,N_15435,N_15455);
or U15668 (N_15668,N_15459,N_15442);
xnor U15669 (N_15669,N_15378,N_15501);
nor U15670 (N_15670,N_15492,N_15393);
and U15671 (N_15671,N_15400,N_15432);
nand U15672 (N_15672,N_15400,N_15494);
and U15673 (N_15673,N_15435,N_15461);
or U15674 (N_15674,N_15400,N_15446);
nor U15675 (N_15675,N_15467,N_15366);
and U15676 (N_15676,N_15445,N_15463);
xnor U15677 (N_15677,N_15496,N_15453);
nand U15678 (N_15678,N_15418,N_15380);
xor U15679 (N_15679,N_15484,N_15430);
nand U15680 (N_15680,N_15561,N_15637);
xnor U15681 (N_15681,N_15549,N_15532);
or U15682 (N_15682,N_15536,N_15626);
nor U15683 (N_15683,N_15607,N_15648);
or U15684 (N_15684,N_15547,N_15534);
xor U15685 (N_15685,N_15624,N_15669);
nor U15686 (N_15686,N_15642,N_15550);
xnor U15687 (N_15687,N_15552,N_15655);
or U15688 (N_15688,N_15528,N_15596);
xnor U15689 (N_15689,N_15543,N_15618);
xnor U15690 (N_15690,N_15546,N_15523);
xor U15691 (N_15691,N_15621,N_15551);
nand U15692 (N_15692,N_15651,N_15629);
nand U15693 (N_15693,N_15526,N_15527);
or U15694 (N_15694,N_15628,N_15557);
nor U15695 (N_15695,N_15612,N_15679);
or U15696 (N_15696,N_15559,N_15582);
nor U15697 (N_15697,N_15524,N_15520);
or U15698 (N_15698,N_15593,N_15563);
nor U15699 (N_15699,N_15592,N_15545);
or U15700 (N_15700,N_15649,N_15539);
xor U15701 (N_15701,N_15652,N_15560);
or U15702 (N_15702,N_15619,N_15564);
nor U15703 (N_15703,N_15646,N_15615);
or U15704 (N_15704,N_15661,N_15583);
nand U15705 (N_15705,N_15673,N_15535);
xor U15706 (N_15706,N_15617,N_15627);
nor U15707 (N_15707,N_15558,N_15657);
nand U15708 (N_15708,N_15633,N_15672);
and U15709 (N_15709,N_15533,N_15554);
or U15710 (N_15710,N_15571,N_15634);
xnor U15711 (N_15711,N_15538,N_15663);
or U15712 (N_15712,N_15668,N_15574);
nand U15713 (N_15713,N_15670,N_15521);
or U15714 (N_15714,N_15556,N_15638);
xnor U15715 (N_15715,N_15529,N_15594);
nor U15716 (N_15716,N_15620,N_15553);
xnor U15717 (N_15717,N_15678,N_15581);
or U15718 (N_15718,N_15664,N_15537);
nand U15719 (N_15719,N_15650,N_15671);
and U15720 (N_15720,N_15542,N_15573);
and U15721 (N_15721,N_15614,N_15608);
xor U15722 (N_15722,N_15606,N_15665);
nand U15723 (N_15723,N_15604,N_15609);
or U15724 (N_15724,N_15610,N_15625);
and U15725 (N_15725,N_15676,N_15565);
nand U15726 (N_15726,N_15643,N_15659);
nor U15727 (N_15727,N_15584,N_15639);
or U15728 (N_15728,N_15569,N_15613);
and U15729 (N_15729,N_15544,N_15570);
nor U15730 (N_15730,N_15635,N_15675);
xnor U15731 (N_15731,N_15595,N_15654);
xnor U15732 (N_15732,N_15576,N_15616);
nand U15733 (N_15733,N_15656,N_15631);
nor U15734 (N_15734,N_15653,N_15555);
xor U15735 (N_15735,N_15644,N_15568);
and U15736 (N_15736,N_15611,N_15522);
nand U15737 (N_15737,N_15575,N_15590);
and U15738 (N_15738,N_15600,N_15640);
and U15739 (N_15739,N_15597,N_15599);
or U15740 (N_15740,N_15667,N_15602);
and U15741 (N_15741,N_15562,N_15588);
nand U15742 (N_15742,N_15601,N_15622);
xnor U15743 (N_15743,N_15603,N_15578);
xnor U15744 (N_15744,N_15666,N_15623);
xor U15745 (N_15745,N_15540,N_15589);
and U15746 (N_15746,N_15662,N_15632);
or U15747 (N_15747,N_15566,N_15548);
or U15748 (N_15748,N_15530,N_15579);
and U15749 (N_15749,N_15641,N_15567);
nor U15750 (N_15750,N_15605,N_15647);
nor U15751 (N_15751,N_15630,N_15636);
or U15752 (N_15752,N_15598,N_15525);
nand U15753 (N_15753,N_15587,N_15660);
or U15754 (N_15754,N_15572,N_15591);
nor U15755 (N_15755,N_15585,N_15541);
xnor U15756 (N_15756,N_15531,N_15658);
nor U15757 (N_15757,N_15645,N_15674);
and U15758 (N_15758,N_15577,N_15586);
or U15759 (N_15759,N_15580,N_15677);
and U15760 (N_15760,N_15529,N_15575);
and U15761 (N_15761,N_15540,N_15628);
nand U15762 (N_15762,N_15627,N_15588);
and U15763 (N_15763,N_15558,N_15648);
nor U15764 (N_15764,N_15527,N_15594);
or U15765 (N_15765,N_15646,N_15644);
and U15766 (N_15766,N_15581,N_15649);
nor U15767 (N_15767,N_15578,N_15634);
and U15768 (N_15768,N_15540,N_15666);
nand U15769 (N_15769,N_15626,N_15634);
xor U15770 (N_15770,N_15591,N_15666);
and U15771 (N_15771,N_15560,N_15549);
and U15772 (N_15772,N_15620,N_15659);
nor U15773 (N_15773,N_15612,N_15530);
nor U15774 (N_15774,N_15620,N_15651);
or U15775 (N_15775,N_15665,N_15575);
nand U15776 (N_15776,N_15526,N_15651);
or U15777 (N_15777,N_15601,N_15547);
xnor U15778 (N_15778,N_15520,N_15550);
nand U15779 (N_15779,N_15577,N_15607);
xor U15780 (N_15780,N_15621,N_15641);
nor U15781 (N_15781,N_15611,N_15607);
and U15782 (N_15782,N_15605,N_15572);
nor U15783 (N_15783,N_15569,N_15542);
and U15784 (N_15784,N_15671,N_15532);
nand U15785 (N_15785,N_15652,N_15678);
xnor U15786 (N_15786,N_15585,N_15593);
nor U15787 (N_15787,N_15583,N_15541);
nor U15788 (N_15788,N_15592,N_15616);
and U15789 (N_15789,N_15586,N_15580);
nand U15790 (N_15790,N_15678,N_15547);
or U15791 (N_15791,N_15673,N_15609);
and U15792 (N_15792,N_15554,N_15590);
nand U15793 (N_15793,N_15640,N_15522);
nand U15794 (N_15794,N_15522,N_15591);
nor U15795 (N_15795,N_15584,N_15662);
nor U15796 (N_15796,N_15596,N_15569);
nor U15797 (N_15797,N_15556,N_15605);
and U15798 (N_15798,N_15618,N_15670);
xnor U15799 (N_15799,N_15555,N_15522);
or U15800 (N_15800,N_15572,N_15637);
nor U15801 (N_15801,N_15678,N_15535);
xor U15802 (N_15802,N_15583,N_15643);
nor U15803 (N_15803,N_15548,N_15573);
nand U15804 (N_15804,N_15589,N_15674);
and U15805 (N_15805,N_15632,N_15646);
nor U15806 (N_15806,N_15641,N_15543);
or U15807 (N_15807,N_15546,N_15619);
nand U15808 (N_15808,N_15650,N_15624);
nor U15809 (N_15809,N_15581,N_15617);
and U15810 (N_15810,N_15552,N_15560);
xnor U15811 (N_15811,N_15595,N_15585);
or U15812 (N_15812,N_15556,N_15531);
nor U15813 (N_15813,N_15568,N_15637);
nor U15814 (N_15814,N_15534,N_15563);
nor U15815 (N_15815,N_15589,N_15651);
xnor U15816 (N_15816,N_15578,N_15622);
xnor U15817 (N_15817,N_15676,N_15645);
or U15818 (N_15818,N_15646,N_15549);
xnor U15819 (N_15819,N_15619,N_15554);
nor U15820 (N_15820,N_15543,N_15551);
and U15821 (N_15821,N_15562,N_15569);
xnor U15822 (N_15822,N_15669,N_15576);
and U15823 (N_15823,N_15593,N_15679);
nor U15824 (N_15824,N_15593,N_15595);
and U15825 (N_15825,N_15572,N_15574);
or U15826 (N_15826,N_15581,N_15606);
nor U15827 (N_15827,N_15628,N_15601);
and U15828 (N_15828,N_15616,N_15585);
xnor U15829 (N_15829,N_15666,N_15575);
or U15830 (N_15830,N_15585,N_15642);
nand U15831 (N_15831,N_15617,N_15532);
xor U15832 (N_15832,N_15580,N_15596);
xnor U15833 (N_15833,N_15573,N_15616);
nand U15834 (N_15834,N_15588,N_15522);
and U15835 (N_15835,N_15666,N_15578);
or U15836 (N_15836,N_15614,N_15615);
or U15837 (N_15837,N_15586,N_15538);
and U15838 (N_15838,N_15621,N_15544);
xnor U15839 (N_15839,N_15645,N_15660);
nand U15840 (N_15840,N_15701,N_15779);
or U15841 (N_15841,N_15760,N_15727);
xor U15842 (N_15842,N_15773,N_15733);
nand U15843 (N_15843,N_15761,N_15832);
or U15844 (N_15844,N_15793,N_15835);
or U15845 (N_15845,N_15752,N_15713);
nor U15846 (N_15846,N_15771,N_15694);
or U15847 (N_15847,N_15783,N_15756);
or U15848 (N_15848,N_15794,N_15681);
and U15849 (N_15849,N_15730,N_15750);
or U15850 (N_15850,N_15768,N_15812);
or U15851 (N_15851,N_15800,N_15709);
xor U15852 (N_15852,N_15719,N_15821);
and U15853 (N_15853,N_15763,N_15827);
nor U15854 (N_15854,N_15767,N_15703);
or U15855 (N_15855,N_15803,N_15697);
xor U15856 (N_15856,N_15829,N_15690);
or U15857 (N_15857,N_15819,N_15755);
nor U15858 (N_15858,N_15789,N_15804);
and U15859 (N_15859,N_15687,N_15809);
nand U15860 (N_15860,N_15784,N_15785);
xor U15861 (N_15861,N_15836,N_15818);
xnor U15862 (N_15862,N_15838,N_15739);
xor U15863 (N_15863,N_15828,N_15743);
or U15864 (N_15864,N_15788,N_15738);
and U15865 (N_15865,N_15751,N_15740);
and U15866 (N_15866,N_15728,N_15698);
and U15867 (N_15867,N_15778,N_15712);
nand U15868 (N_15868,N_15782,N_15805);
or U15869 (N_15869,N_15754,N_15820);
nand U15870 (N_15870,N_15683,N_15765);
xor U15871 (N_15871,N_15688,N_15815);
or U15872 (N_15872,N_15834,N_15684);
nand U15873 (N_15873,N_15797,N_15776);
nor U15874 (N_15874,N_15796,N_15721);
and U15875 (N_15875,N_15737,N_15708);
nor U15876 (N_15876,N_15723,N_15731);
nand U15877 (N_15877,N_15724,N_15706);
xnor U15878 (N_15878,N_15748,N_15718);
or U15879 (N_15879,N_15839,N_15813);
or U15880 (N_15880,N_15814,N_15770);
nor U15881 (N_15881,N_15810,N_15833);
xor U15882 (N_15882,N_15746,N_15799);
and U15883 (N_15883,N_15682,N_15747);
and U15884 (N_15884,N_15823,N_15753);
and U15885 (N_15885,N_15759,N_15802);
or U15886 (N_15886,N_15826,N_15736);
nand U15887 (N_15887,N_15774,N_15705);
or U15888 (N_15888,N_15741,N_15685);
xor U15889 (N_15889,N_15807,N_15787);
and U15890 (N_15890,N_15786,N_15790);
and U15891 (N_15891,N_15830,N_15792);
nand U15892 (N_15892,N_15714,N_15734);
and U15893 (N_15893,N_15717,N_15816);
xor U15894 (N_15894,N_15825,N_15795);
or U15895 (N_15895,N_15689,N_15725);
nor U15896 (N_15896,N_15729,N_15680);
or U15897 (N_15897,N_15811,N_15686);
or U15898 (N_15898,N_15780,N_15742);
and U15899 (N_15899,N_15716,N_15817);
nand U15900 (N_15900,N_15693,N_15831);
xor U15901 (N_15901,N_15700,N_15824);
and U15902 (N_15902,N_15691,N_15769);
xnor U15903 (N_15903,N_15798,N_15837);
xnor U15904 (N_15904,N_15692,N_15749);
or U15905 (N_15905,N_15710,N_15711);
or U15906 (N_15906,N_15757,N_15696);
and U15907 (N_15907,N_15745,N_15707);
nand U15908 (N_15908,N_15715,N_15806);
nor U15909 (N_15909,N_15722,N_15702);
xor U15910 (N_15910,N_15762,N_15764);
xnor U15911 (N_15911,N_15732,N_15791);
or U15912 (N_15912,N_15777,N_15766);
xor U15913 (N_15913,N_15808,N_15735);
and U15914 (N_15914,N_15704,N_15726);
xnor U15915 (N_15915,N_15720,N_15781);
and U15916 (N_15916,N_15744,N_15775);
nand U15917 (N_15917,N_15758,N_15699);
nand U15918 (N_15918,N_15822,N_15801);
or U15919 (N_15919,N_15772,N_15695);
and U15920 (N_15920,N_15825,N_15774);
nor U15921 (N_15921,N_15814,N_15722);
nand U15922 (N_15922,N_15826,N_15775);
and U15923 (N_15923,N_15760,N_15703);
nand U15924 (N_15924,N_15755,N_15716);
and U15925 (N_15925,N_15742,N_15835);
nand U15926 (N_15926,N_15760,N_15712);
and U15927 (N_15927,N_15754,N_15839);
xor U15928 (N_15928,N_15762,N_15806);
and U15929 (N_15929,N_15757,N_15760);
or U15930 (N_15930,N_15812,N_15690);
nor U15931 (N_15931,N_15795,N_15778);
nor U15932 (N_15932,N_15837,N_15713);
and U15933 (N_15933,N_15792,N_15796);
nor U15934 (N_15934,N_15782,N_15749);
or U15935 (N_15935,N_15739,N_15681);
xnor U15936 (N_15936,N_15704,N_15747);
nand U15937 (N_15937,N_15692,N_15795);
xor U15938 (N_15938,N_15703,N_15734);
xnor U15939 (N_15939,N_15758,N_15777);
xnor U15940 (N_15940,N_15780,N_15774);
and U15941 (N_15941,N_15789,N_15817);
and U15942 (N_15942,N_15735,N_15702);
nand U15943 (N_15943,N_15743,N_15815);
xnor U15944 (N_15944,N_15781,N_15751);
or U15945 (N_15945,N_15779,N_15825);
xnor U15946 (N_15946,N_15710,N_15749);
nor U15947 (N_15947,N_15782,N_15712);
and U15948 (N_15948,N_15768,N_15749);
xnor U15949 (N_15949,N_15789,N_15744);
nand U15950 (N_15950,N_15734,N_15755);
and U15951 (N_15951,N_15763,N_15728);
nor U15952 (N_15952,N_15691,N_15731);
nand U15953 (N_15953,N_15786,N_15698);
or U15954 (N_15954,N_15821,N_15817);
or U15955 (N_15955,N_15723,N_15783);
or U15956 (N_15956,N_15739,N_15779);
nand U15957 (N_15957,N_15831,N_15825);
nor U15958 (N_15958,N_15695,N_15706);
nor U15959 (N_15959,N_15739,N_15750);
nand U15960 (N_15960,N_15821,N_15714);
nor U15961 (N_15961,N_15817,N_15830);
nor U15962 (N_15962,N_15810,N_15790);
nand U15963 (N_15963,N_15782,N_15730);
nor U15964 (N_15964,N_15782,N_15704);
nand U15965 (N_15965,N_15695,N_15715);
nand U15966 (N_15966,N_15817,N_15757);
nor U15967 (N_15967,N_15707,N_15734);
nor U15968 (N_15968,N_15696,N_15717);
and U15969 (N_15969,N_15710,N_15783);
xor U15970 (N_15970,N_15815,N_15838);
xor U15971 (N_15971,N_15686,N_15688);
xor U15972 (N_15972,N_15798,N_15801);
and U15973 (N_15973,N_15777,N_15749);
or U15974 (N_15974,N_15697,N_15794);
nor U15975 (N_15975,N_15745,N_15728);
xnor U15976 (N_15976,N_15808,N_15688);
nand U15977 (N_15977,N_15812,N_15777);
or U15978 (N_15978,N_15709,N_15819);
xor U15979 (N_15979,N_15689,N_15801);
nand U15980 (N_15980,N_15728,N_15834);
nand U15981 (N_15981,N_15806,N_15685);
or U15982 (N_15982,N_15831,N_15782);
xnor U15983 (N_15983,N_15734,N_15766);
nand U15984 (N_15984,N_15762,N_15696);
or U15985 (N_15985,N_15761,N_15749);
or U15986 (N_15986,N_15831,N_15828);
xnor U15987 (N_15987,N_15818,N_15798);
and U15988 (N_15988,N_15710,N_15782);
or U15989 (N_15989,N_15731,N_15715);
nor U15990 (N_15990,N_15740,N_15735);
nand U15991 (N_15991,N_15773,N_15750);
and U15992 (N_15992,N_15834,N_15817);
xnor U15993 (N_15993,N_15758,N_15811);
or U15994 (N_15994,N_15691,N_15760);
nand U15995 (N_15995,N_15832,N_15788);
and U15996 (N_15996,N_15708,N_15750);
xor U15997 (N_15997,N_15681,N_15783);
and U15998 (N_15998,N_15748,N_15771);
xor U15999 (N_15999,N_15795,N_15754);
and U16000 (N_16000,N_15960,N_15930);
or U16001 (N_16001,N_15994,N_15847);
nand U16002 (N_16002,N_15969,N_15944);
and U16003 (N_16003,N_15995,N_15842);
and U16004 (N_16004,N_15937,N_15895);
nor U16005 (N_16005,N_15891,N_15855);
nor U16006 (N_16006,N_15975,N_15907);
or U16007 (N_16007,N_15902,N_15840);
nor U16008 (N_16008,N_15971,N_15862);
xor U16009 (N_16009,N_15924,N_15997);
xor U16010 (N_16010,N_15892,N_15938);
nor U16011 (N_16011,N_15906,N_15950);
and U16012 (N_16012,N_15955,N_15933);
and U16013 (N_16013,N_15874,N_15935);
nand U16014 (N_16014,N_15999,N_15977);
nor U16015 (N_16015,N_15945,N_15851);
and U16016 (N_16016,N_15972,N_15867);
xnor U16017 (N_16017,N_15910,N_15913);
nand U16018 (N_16018,N_15954,N_15959);
nor U16019 (N_16019,N_15992,N_15989);
or U16020 (N_16020,N_15889,N_15864);
xnor U16021 (N_16021,N_15878,N_15883);
and U16022 (N_16022,N_15923,N_15958);
or U16023 (N_16023,N_15908,N_15856);
nand U16024 (N_16024,N_15849,N_15979);
xnor U16025 (N_16025,N_15934,N_15964);
and U16026 (N_16026,N_15888,N_15848);
nand U16027 (N_16027,N_15911,N_15914);
or U16028 (N_16028,N_15931,N_15904);
nand U16029 (N_16029,N_15976,N_15980);
and U16030 (N_16030,N_15900,N_15860);
and U16031 (N_16031,N_15841,N_15857);
nand U16032 (N_16032,N_15915,N_15854);
or U16033 (N_16033,N_15876,N_15939);
or U16034 (N_16034,N_15925,N_15927);
nor U16035 (N_16035,N_15880,N_15920);
nor U16036 (N_16036,N_15897,N_15973);
nor U16037 (N_16037,N_15918,N_15881);
nor U16038 (N_16038,N_15877,N_15863);
nor U16039 (N_16039,N_15943,N_15947);
xnor U16040 (N_16040,N_15896,N_15861);
or U16041 (N_16041,N_15919,N_15993);
or U16042 (N_16042,N_15879,N_15853);
nor U16043 (N_16043,N_15988,N_15875);
nor U16044 (N_16044,N_15957,N_15982);
or U16045 (N_16045,N_15885,N_15845);
or U16046 (N_16046,N_15991,N_15872);
and U16047 (N_16047,N_15963,N_15985);
nor U16048 (N_16048,N_15894,N_15865);
or U16049 (N_16049,N_15868,N_15893);
and U16050 (N_16050,N_15996,N_15974);
nor U16051 (N_16051,N_15952,N_15898);
nor U16052 (N_16052,N_15951,N_15887);
nand U16053 (N_16053,N_15941,N_15882);
or U16054 (N_16054,N_15871,N_15984);
nand U16055 (N_16055,N_15940,N_15899);
nand U16056 (N_16056,N_15953,N_15990);
nand U16057 (N_16057,N_15843,N_15962);
nor U16058 (N_16058,N_15981,N_15932);
or U16059 (N_16059,N_15948,N_15986);
and U16060 (N_16060,N_15978,N_15873);
nor U16061 (N_16061,N_15869,N_15850);
or U16062 (N_16062,N_15965,N_15909);
nand U16063 (N_16063,N_15921,N_15928);
or U16064 (N_16064,N_15967,N_15942);
or U16065 (N_16065,N_15912,N_15946);
and U16066 (N_16066,N_15929,N_15961);
and U16067 (N_16067,N_15936,N_15852);
and U16068 (N_16068,N_15983,N_15859);
or U16069 (N_16069,N_15956,N_15916);
xnor U16070 (N_16070,N_15870,N_15844);
nand U16071 (N_16071,N_15968,N_15998);
xor U16072 (N_16072,N_15884,N_15905);
xnor U16073 (N_16073,N_15987,N_15846);
nor U16074 (N_16074,N_15926,N_15922);
xor U16075 (N_16075,N_15890,N_15886);
xnor U16076 (N_16076,N_15917,N_15970);
and U16077 (N_16077,N_15903,N_15866);
or U16078 (N_16078,N_15949,N_15901);
nand U16079 (N_16079,N_15858,N_15966);
nor U16080 (N_16080,N_15869,N_15941);
and U16081 (N_16081,N_15905,N_15970);
or U16082 (N_16082,N_15893,N_15955);
or U16083 (N_16083,N_15978,N_15880);
nor U16084 (N_16084,N_15935,N_15958);
nand U16085 (N_16085,N_15840,N_15964);
xor U16086 (N_16086,N_15923,N_15999);
nor U16087 (N_16087,N_15866,N_15948);
xnor U16088 (N_16088,N_15901,N_15898);
nor U16089 (N_16089,N_15855,N_15956);
xnor U16090 (N_16090,N_15973,N_15876);
xor U16091 (N_16091,N_15966,N_15943);
nor U16092 (N_16092,N_15908,N_15903);
or U16093 (N_16093,N_15906,N_15881);
and U16094 (N_16094,N_15920,N_15964);
and U16095 (N_16095,N_15933,N_15880);
and U16096 (N_16096,N_15895,N_15869);
or U16097 (N_16097,N_15873,N_15885);
or U16098 (N_16098,N_15863,N_15925);
and U16099 (N_16099,N_15958,N_15950);
nand U16100 (N_16100,N_15943,N_15863);
nand U16101 (N_16101,N_15995,N_15941);
nor U16102 (N_16102,N_15967,N_15887);
nand U16103 (N_16103,N_15847,N_15927);
nand U16104 (N_16104,N_15951,N_15920);
or U16105 (N_16105,N_15862,N_15983);
nor U16106 (N_16106,N_15953,N_15879);
or U16107 (N_16107,N_15943,N_15938);
and U16108 (N_16108,N_15888,N_15990);
nand U16109 (N_16109,N_15877,N_15997);
or U16110 (N_16110,N_15941,N_15892);
nand U16111 (N_16111,N_15928,N_15957);
or U16112 (N_16112,N_15972,N_15903);
xor U16113 (N_16113,N_15946,N_15887);
nor U16114 (N_16114,N_15998,N_15983);
nand U16115 (N_16115,N_15912,N_15967);
xor U16116 (N_16116,N_15893,N_15871);
or U16117 (N_16117,N_15895,N_15977);
or U16118 (N_16118,N_15973,N_15915);
and U16119 (N_16119,N_15901,N_15982);
nor U16120 (N_16120,N_15879,N_15886);
and U16121 (N_16121,N_15970,N_15962);
nand U16122 (N_16122,N_15935,N_15850);
and U16123 (N_16123,N_15911,N_15846);
or U16124 (N_16124,N_15979,N_15899);
and U16125 (N_16125,N_15982,N_15892);
xnor U16126 (N_16126,N_15900,N_15935);
nand U16127 (N_16127,N_15890,N_15865);
and U16128 (N_16128,N_15871,N_15915);
and U16129 (N_16129,N_15905,N_15851);
or U16130 (N_16130,N_15961,N_15913);
and U16131 (N_16131,N_15943,N_15900);
nor U16132 (N_16132,N_15961,N_15940);
and U16133 (N_16133,N_15862,N_15843);
or U16134 (N_16134,N_15973,N_15993);
nand U16135 (N_16135,N_15924,N_15985);
and U16136 (N_16136,N_15846,N_15845);
nand U16137 (N_16137,N_15913,N_15879);
and U16138 (N_16138,N_15914,N_15938);
nand U16139 (N_16139,N_15868,N_15981);
nor U16140 (N_16140,N_15992,N_15960);
nand U16141 (N_16141,N_15861,N_15892);
xor U16142 (N_16142,N_15857,N_15846);
or U16143 (N_16143,N_15902,N_15914);
or U16144 (N_16144,N_15965,N_15975);
nand U16145 (N_16145,N_15908,N_15995);
nor U16146 (N_16146,N_15896,N_15939);
nand U16147 (N_16147,N_15959,N_15953);
nor U16148 (N_16148,N_15973,N_15972);
nand U16149 (N_16149,N_15986,N_15975);
nand U16150 (N_16150,N_15898,N_15907);
and U16151 (N_16151,N_15862,N_15966);
or U16152 (N_16152,N_15857,N_15923);
xor U16153 (N_16153,N_15912,N_15890);
nor U16154 (N_16154,N_15973,N_15916);
nor U16155 (N_16155,N_15927,N_15841);
xnor U16156 (N_16156,N_15982,N_15980);
and U16157 (N_16157,N_15933,N_15964);
xor U16158 (N_16158,N_15855,N_15899);
nand U16159 (N_16159,N_15853,N_15941);
nand U16160 (N_16160,N_16029,N_16061);
or U16161 (N_16161,N_16072,N_16091);
nor U16162 (N_16162,N_16048,N_16124);
and U16163 (N_16163,N_16112,N_16095);
or U16164 (N_16164,N_16100,N_16110);
and U16165 (N_16165,N_16005,N_16001);
nand U16166 (N_16166,N_16036,N_16122);
nor U16167 (N_16167,N_16086,N_16125);
xnor U16168 (N_16168,N_16105,N_16006);
and U16169 (N_16169,N_16157,N_16003);
nor U16170 (N_16170,N_16021,N_16115);
xnor U16171 (N_16171,N_16130,N_16034);
or U16172 (N_16172,N_16056,N_16081);
or U16173 (N_16173,N_16062,N_16129);
and U16174 (N_16174,N_16120,N_16084);
and U16175 (N_16175,N_16015,N_16045);
nand U16176 (N_16176,N_16018,N_16077);
or U16177 (N_16177,N_16136,N_16089);
nand U16178 (N_16178,N_16069,N_16052);
or U16179 (N_16179,N_16108,N_16134);
xor U16180 (N_16180,N_16090,N_16146);
xor U16181 (N_16181,N_16007,N_16153);
xnor U16182 (N_16182,N_16025,N_16002);
nor U16183 (N_16183,N_16082,N_16019);
nor U16184 (N_16184,N_16060,N_16059);
nand U16185 (N_16185,N_16030,N_16123);
or U16186 (N_16186,N_16039,N_16093);
or U16187 (N_16187,N_16079,N_16098);
nor U16188 (N_16188,N_16118,N_16132);
xnor U16189 (N_16189,N_16078,N_16073);
nand U16190 (N_16190,N_16102,N_16088);
nand U16191 (N_16191,N_16070,N_16139);
or U16192 (N_16192,N_16063,N_16028);
or U16193 (N_16193,N_16128,N_16033);
and U16194 (N_16194,N_16023,N_16109);
or U16195 (N_16195,N_16154,N_16092);
or U16196 (N_16196,N_16016,N_16074);
xnor U16197 (N_16197,N_16013,N_16044);
or U16198 (N_16198,N_16131,N_16126);
or U16199 (N_16199,N_16083,N_16011);
nor U16200 (N_16200,N_16049,N_16101);
or U16201 (N_16201,N_16000,N_16155);
xor U16202 (N_16202,N_16087,N_16113);
nor U16203 (N_16203,N_16145,N_16037);
nand U16204 (N_16204,N_16152,N_16046);
nand U16205 (N_16205,N_16156,N_16032);
xor U16206 (N_16206,N_16121,N_16119);
or U16207 (N_16207,N_16064,N_16022);
xor U16208 (N_16208,N_16020,N_16009);
xnor U16209 (N_16209,N_16043,N_16142);
and U16210 (N_16210,N_16097,N_16111);
and U16211 (N_16211,N_16085,N_16104);
and U16212 (N_16212,N_16041,N_16058);
and U16213 (N_16213,N_16107,N_16114);
or U16214 (N_16214,N_16159,N_16158);
or U16215 (N_16215,N_16076,N_16038);
nand U16216 (N_16216,N_16024,N_16099);
and U16217 (N_16217,N_16065,N_16138);
xnor U16218 (N_16218,N_16137,N_16031);
xnor U16219 (N_16219,N_16010,N_16067);
or U16220 (N_16220,N_16055,N_16149);
xor U16221 (N_16221,N_16143,N_16148);
and U16222 (N_16222,N_16094,N_16080);
nor U16223 (N_16223,N_16066,N_16057);
nand U16224 (N_16224,N_16027,N_16147);
and U16225 (N_16225,N_16135,N_16004);
or U16226 (N_16226,N_16047,N_16117);
nor U16227 (N_16227,N_16054,N_16042);
nor U16228 (N_16228,N_16106,N_16144);
or U16229 (N_16229,N_16141,N_16150);
and U16230 (N_16230,N_16103,N_16051);
and U16231 (N_16231,N_16012,N_16133);
nor U16232 (N_16232,N_16140,N_16026);
nand U16233 (N_16233,N_16053,N_16116);
nor U16234 (N_16234,N_16127,N_16008);
nor U16235 (N_16235,N_16017,N_16151);
nand U16236 (N_16236,N_16071,N_16040);
nand U16237 (N_16237,N_16068,N_16035);
nand U16238 (N_16238,N_16050,N_16096);
and U16239 (N_16239,N_16014,N_16075);
xnor U16240 (N_16240,N_16115,N_16066);
or U16241 (N_16241,N_16106,N_16046);
nand U16242 (N_16242,N_16008,N_16114);
or U16243 (N_16243,N_16036,N_16101);
xor U16244 (N_16244,N_16035,N_16012);
and U16245 (N_16245,N_16033,N_16091);
or U16246 (N_16246,N_16106,N_16049);
nor U16247 (N_16247,N_16000,N_16136);
nand U16248 (N_16248,N_16145,N_16129);
nor U16249 (N_16249,N_16088,N_16026);
xor U16250 (N_16250,N_16112,N_16144);
or U16251 (N_16251,N_16060,N_16117);
and U16252 (N_16252,N_16144,N_16129);
and U16253 (N_16253,N_16082,N_16150);
nor U16254 (N_16254,N_16024,N_16156);
and U16255 (N_16255,N_16146,N_16116);
and U16256 (N_16256,N_16055,N_16102);
and U16257 (N_16257,N_16066,N_16098);
xnor U16258 (N_16258,N_16087,N_16110);
and U16259 (N_16259,N_16112,N_16022);
or U16260 (N_16260,N_16075,N_16035);
or U16261 (N_16261,N_16111,N_16011);
or U16262 (N_16262,N_16085,N_16012);
nor U16263 (N_16263,N_16037,N_16003);
nor U16264 (N_16264,N_16094,N_16081);
nand U16265 (N_16265,N_16111,N_16041);
nand U16266 (N_16266,N_16100,N_16133);
nor U16267 (N_16267,N_16140,N_16119);
nand U16268 (N_16268,N_16114,N_16090);
or U16269 (N_16269,N_16087,N_16001);
nand U16270 (N_16270,N_16138,N_16011);
nand U16271 (N_16271,N_16005,N_16034);
nor U16272 (N_16272,N_16128,N_16038);
or U16273 (N_16273,N_16020,N_16158);
nand U16274 (N_16274,N_16066,N_16077);
nand U16275 (N_16275,N_16099,N_16000);
xor U16276 (N_16276,N_16075,N_16026);
or U16277 (N_16277,N_16089,N_16040);
nor U16278 (N_16278,N_16102,N_16082);
nand U16279 (N_16279,N_16137,N_16046);
nor U16280 (N_16280,N_16119,N_16100);
or U16281 (N_16281,N_16125,N_16025);
and U16282 (N_16282,N_16145,N_16137);
or U16283 (N_16283,N_16139,N_16025);
nand U16284 (N_16284,N_16153,N_16043);
nor U16285 (N_16285,N_16139,N_16006);
or U16286 (N_16286,N_16048,N_16098);
nor U16287 (N_16287,N_16071,N_16103);
xnor U16288 (N_16288,N_16105,N_16033);
nor U16289 (N_16289,N_16019,N_16159);
nand U16290 (N_16290,N_16136,N_16142);
xor U16291 (N_16291,N_16156,N_16035);
or U16292 (N_16292,N_16094,N_16060);
and U16293 (N_16293,N_16023,N_16091);
or U16294 (N_16294,N_16085,N_16108);
and U16295 (N_16295,N_16154,N_16128);
nand U16296 (N_16296,N_16091,N_16070);
and U16297 (N_16297,N_16108,N_16084);
xnor U16298 (N_16298,N_16032,N_16015);
nand U16299 (N_16299,N_16032,N_16062);
or U16300 (N_16300,N_16079,N_16063);
or U16301 (N_16301,N_16027,N_16108);
xnor U16302 (N_16302,N_16035,N_16108);
xor U16303 (N_16303,N_16115,N_16080);
xor U16304 (N_16304,N_16123,N_16034);
nor U16305 (N_16305,N_16096,N_16007);
and U16306 (N_16306,N_16132,N_16002);
xnor U16307 (N_16307,N_16034,N_16020);
nor U16308 (N_16308,N_16007,N_16157);
and U16309 (N_16309,N_16059,N_16093);
and U16310 (N_16310,N_16069,N_16050);
nor U16311 (N_16311,N_16005,N_16025);
or U16312 (N_16312,N_16148,N_16050);
or U16313 (N_16313,N_16127,N_16126);
nand U16314 (N_16314,N_16147,N_16034);
or U16315 (N_16315,N_16091,N_16009);
and U16316 (N_16316,N_16066,N_16102);
or U16317 (N_16317,N_16028,N_16036);
nand U16318 (N_16318,N_16101,N_16026);
xor U16319 (N_16319,N_16058,N_16107);
xnor U16320 (N_16320,N_16240,N_16286);
and U16321 (N_16321,N_16207,N_16270);
and U16322 (N_16322,N_16220,N_16250);
and U16323 (N_16323,N_16298,N_16314);
or U16324 (N_16324,N_16266,N_16161);
and U16325 (N_16325,N_16249,N_16305);
or U16326 (N_16326,N_16315,N_16312);
or U16327 (N_16327,N_16313,N_16200);
xor U16328 (N_16328,N_16255,N_16281);
or U16329 (N_16329,N_16204,N_16259);
nand U16330 (N_16330,N_16188,N_16199);
nand U16331 (N_16331,N_16252,N_16191);
or U16332 (N_16332,N_16289,N_16244);
nand U16333 (N_16333,N_16277,N_16183);
nor U16334 (N_16334,N_16318,N_16304);
xnor U16335 (N_16335,N_16301,N_16162);
and U16336 (N_16336,N_16180,N_16216);
xnor U16337 (N_16337,N_16309,N_16310);
xor U16338 (N_16338,N_16170,N_16215);
or U16339 (N_16339,N_16316,N_16175);
nand U16340 (N_16340,N_16168,N_16275);
and U16341 (N_16341,N_16261,N_16218);
and U16342 (N_16342,N_16276,N_16195);
or U16343 (N_16343,N_16299,N_16166);
or U16344 (N_16344,N_16317,N_16272);
or U16345 (N_16345,N_16201,N_16178);
or U16346 (N_16346,N_16292,N_16209);
nand U16347 (N_16347,N_16253,N_16222);
xnor U16348 (N_16348,N_16238,N_16284);
or U16349 (N_16349,N_16193,N_16234);
nor U16350 (N_16350,N_16287,N_16184);
or U16351 (N_16351,N_16221,N_16243);
or U16352 (N_16352,N_16248,N_16293);
or U16353 (N_16353,N_16267,N_16311);
or U16354 (N_16354,N_16273,N_16308);
xor U16355 (N_16355,N_16208,N_16225);
xor U16356 (N_16356,N_16256,N_16290);
xor U16357 (N_16357,N_16260,N_16295);
xnor U16358 (N_16358,N_16210,N_16211);
xor U16359 (N_16359,N_16194,N_16232);
nor U16360 (N_16360,N_16163,N_16227);
nand U16361 (N_16361,N_16202,N_16288);
and U16362 (N_16362,N_16274,N_16294);
nor U16363 (N_16363,N_16177,N_16229);
or U16364 (N_16364,N_16235,N_16206);
and U16365 (N_16365,N_16185,N_16282);
nand U16366 (N_16366,N_16224,N_16291);
nand U16367 (N_16367,N_16176,N_16280);
and U16368 (N_16368,N_16228,N_16283);
or U16369 (N_16369,N_16212,N_16296);
or U16370 (N_16370,N_16262,N_16285);
and U16371 (N_16371,N_16181,N_16197);
or U16372 (N_16372,N_16190,N_16173);
xnor U16373 (N_16373,N_16264,N_16196);
or U16374 (N_16374,N_16236,N_16233);
xor U16375 (N_16375,N_16169,N_16223);
nor U16376 (N_16376,N_16254,N_16306);
xnor U16377 (N_16377,N_16271,N_16319);
or U16378 (N_16378,N_16217,N_16302);
and U16379 (N_16379,N_16268,N_16179);
or U16380 (N_16380,N_16213,N_16205);
and U16381 (N_16381,N_16226,N_16186);
and U16382 (N_16382,N_16279,N_16251);
nor U16383 (N_16383,N_16265,N_16303);
or U16384 (N_16384,N_16297,N_16245);
nand U16385 (N_16385,N_16263,N_16219);
xnor U16386 (N_16386,N_16231,N_16165);
or U16387 (N_16387,N_16278,N_16237);
xnor U16388 (N_16388,N_16203,N_16269);
and U16389 (N_16389,N_16300,N_16242);
and U16390 (N_16390,N_16257,N_16230);
xor U16391 (N_16391,N_16247,N_16182);
and U16392 (N_16392,N_16164,N_16172);
or U16393 (N_16393,N_16241,N_16192);
nor U16394 (N_16394,N_16187,N_16189);
nand U16395 (N_16395,N_16167,N_16198);
nor U16396 (N_16396,N_16174,N_16258);
or U16397 (N_16397,N_16239,N_16160);
or U16398 (N_16398,N_16171,N_16307);
or U16399 (N_16399,N_16214,N_16246);
nor U16400 (N_16400,N_16237,N_16290);
nand U16401 (N_16401,N_16309,N_16255);
nand U16402 (N_16402,N_16258,N_16170);
xor U16403 (N_16403,N_16200,N_16206);
nor U16404 (N_16404,N_16186,N_16308);
and U16405 (N_16405,N_16291,N_16280);
xnor U16406 (N_16406,N_16279,N_16260);
nor U16407 (N_16407,N_16297,N_16269);
and U16408 (N_16408,N_16250,N_16218);
xnor U16409 (N_16409,N_16206,N_16261);
xnor U16410 (N_16410,N_16268,N_16244);
nor U16411 (N_16411,N_16177,N_16305);
nor U16412 (N_16412,N_16218,N_16235);
xnor U16413 (N_16413,N_16319,N_16283);
xor U16414 (N_16414,N_16291,N_16282);
and U16415 (N_16415,N_16168,N_16230);
and U16416 (N_16416,N_16318,N_16296);
xor U16417 (N_16417,N_16216,N_16199);
xnor U16418 (N_16418,N_16206,N_16236);
nand U16419 (N_16419,N_16210,N_16283);
and U16420 (N_16420,N_16263,N_16260);
nand U16421 (N_16421,N_16277,N_16161);
or U16422 (N_16422,N_16316,N_16296);
nor U16423 (N_16423,N_16234,N_16225);
xor U16424 (N_16424,N_16297,N_16224);
xor U16425 (N_16425,N_16235,N_16307);
or U16426 (N_16426,N_16303,N_16213);
or U16427 (N_16427,N_16312,N_16241);
nand U16428 (N_16428,N_16191,N_16208);
or U16429 (N_16429,N_16284,N_16267);
nand U16430 (N_16430,N_16180,N_16204);
or U16431 (N_16431,N_16287,N_16244);
and U16432 (N_16432,N_16274,N_16172);
nor U16433 (N_16433,N_16255,N_16229);
or U16434 (N_16434,N_16236,N_16253);
nor U16435 (N_16435,N_16203,N_16272);
or U16436 (N_16436,N_16213,N_16169);
nand U16437 (N_16437,N_16289,N_16288);
nand U16438 (N_16438,N_16178,N_16192);
nand U16439 (N_16439,N_16288,N_16308);
or U16440 (N_16440,N_16283,N_16306);
xor U16441 (N_16441,N_16242,N_16284);
or U16442 (N_16442,N_16299,N_16195);
or U16443 (N_16443,N_16218,N_16280);
xnor U16444 (N_16444,N_16257,N_16241);
xnor U16445 (N_16445,N_16212,N_16207);
and U16446 (N_16446,N_16191,N_16258);
xor U16447 (N_16447,N_16197,N_16285);
nor U16448 (N_16448,N_16211,N_16310);
xnor U16449 (N_16449,N_16290,N_16194);
and U16450 (N_16450,N_16271,N_16261);
and U16451 (N_16451,N_16182,N_16205);
and U16452 (N_16452,N_16211,N_16307);
and U16453 (N_16453,N_16202,N_16305);
xor U16454 (N_16454,N_16266,N_16251);
nor U16455 (N_16455,N_16196,N_16276);
nand U16456 (N_16456,N_16164,N_16301);
nand U16457 (N_16457,N_16308,N_16213);
nor U16458 (N_16458,N_16290,N_16219);
or U16459 (N_16459,N_16269,N_16274);
nand U16460 (N_16460,N_16196,N_16175);
nand U16461 (N_16461,N_16262,N_16253);
nand U16462 (N_16462,N_16271,N_16215);
nand U16463 (N_16463,N_16188,N_16196);
nor U16464 (N_16464,N_16164,N_16249);
xor U16465 (N_16465,N_16262,N_16304);
and U16466 (N_16466,N_16235,N_16258);
or U16467 (N_16467,N_16173,N_16161);
nor U16468 (N_16468,N_16179,N_16297);
nand U16469 (N_16469,N_16177,N_16306);
xor U16470 (N_16470,N_16272,N_16216);
nor U16471 (N_16471,N_16178,N_16182);
and U16472 (N_16472,N_16229,N_16298);
xor U16473 (N_16473,N_16205,N_16196);
nor U16474 (N_16474,N_16238,N_16216);
or U16475 (N_16475,N_16284,N_16235);
and U16476 (N_16476,N_16184,N_16249);
nor U16477 (N_16477,N_16273,N_16319);
and U16478 (N_16478,N_16184,N_16307);
xor U16479 (N_16479,N_16309,N_16161);
and U16480 (N_16480,N_16344,N_16413);
xnor U16481 (N_16481,N_16334,N_16401);
and U16482 (N_16482,N_16351,N_16391);
xor U16483 (N_16483,N_16365,N_16336);
and U16484 (N_16484,N_16468,N_16352);
nand U16485 (N_16485,N_16458,N_16361);
xor U16486 (N_16486,N_16476,N_16337);
or U16487 (N_16487,N_16415,N_16350);
xnor U16488 (N_16488,N_16470,N_16434);
or U16489 (N_16489,N_16385,N_16323);
nand U16490 (N_16490,N_16327,N_16362);
nand U16491 (N_16491,N_16451,N_16399);
nand U16492 (N_16492,N_16417,N_16437);
and U16493 (N_16493,N_16363,N_16338);
nand U16494 (N_16494,N_16364,N_16423);
or U16495 (N_16495,N_16424,N_16340);
xnor U16496 (N_16496,N_16408,N_16456);
and U16497 (N_16497,N_16403,N_16421);
nand U16498 (N_16498,N_16452,N_16325);
nand U16499 (N_16499,N_16371,N_16404);
and U16500 (N_16500,N_16359,N_16477);
nand U16501 (N_16501,N_16430,N_16353);
xnor U16502 (N_16502,N_16422,N_16394);
nand U16503 (N_16503,N_16378,N_16357);
xnor U16504 (N_16504,N_16412,N_16384);
nand U16505 (N_16505,N_16465,N_16383);
or U16506 (N_16506,N_16374,N_16464);
xnor U16507 (N_16507,N_16478,N_16455);
or U16508 (N_16508,N_16405,N_16380);
and U16509 (N_16509,N_16427,N_16466);
nor U16510 (N_16510,N_16469,N_16400);
nor U16511 (N_16511,N_16441,N_16443);
xnor U16512 (N_16512,N_16360,N_16330);
nor U16513 (N_16513,N_16460,N_16396);
nor U16514 (N_16514,N_16356,N_16348);
and U16515 (N_16515,N_16445,N_16322);
nand U16516 (N_16516,N_16369,N_16388);
or U16517 (N_16517,N_16375,N_16407);
xor U16518 (N_16518,N_16321,N_16471);
nor U16519 (N_16519,N_16345,N_16432);
and U16520 (N_16520,N_16377,N_16475);
nand U16521 (N_16521,N_16370,N_16331);
nand U16522 (N_16522,N_16411,N_16390);
nor U16523 (N_16523,N_16376,N_16347);
and U16524 (N_16524,N_16341,N_16339);
or U16525 (N_16525,N_16395,N_16342);
xor U16526 (N_16526,N_16392,N_16393);
xor U16527 (N_16527,N_16416,N_16436);
nor U16528 (N_16528,N_16387,N_16332);
or U16529 (N_16529,N_16381,N_16473);
nor U16530 (N_16530,N_16439,N_16329);
or U16531 (N_16531,N_16457,N_16409);
and U16532 (N_16532,N_16467,N_16326);
nand U16533 (N_16533,N_16418,N_16435);
nor U16534 (N_16534,N_16397,N_16474);
or U16535 (N_16535,N_16438,N_16410);
xnor U16536 (N_16536,N_16419,N_16442);
nand U16537 (N_16537,N_16453,N_16402);
nor U16538 (N_16538,N_16368,N_16461);
nor U16539 (N_16539,N_16446,N_16354);
xnor U16540 (N_16540,N_16382,N_16349);
nor U16541 (N_16541,N_16450,N_16358);
xnor U16542 (N_16542,N_16428,N_16431);
or U16543 (N_16543,N_16320,N_16444);
xor U16544 (N_16544,N_16429,N_16328);
nor U16545 (N_16545,N_16433,N_16449);
or U16546 (N_16546,N_16367,N_16448);
xnor U16547 (N_16547,N_16386,N_16462);
nand U16548 (N_16548,N_16420,N_16343);
and U16549 (N_16549,N_16459,N_16372);
nand U16550 (N_16550,N_16346,N_16389);
nand U16551 (N_16551,N_16447,N_16373);
or U16552 (N_16552,N_16440,N_16355);
nor U16553 (N_16553,N_16333,N_16324);
or U16554 (N_16554,N_16426,N_16479);
and U16555 (N_16555,N_16454,N_16406);
and U16556 (N_16556,N_16398,N_16379);
or U16557 (N_16557,N_16425,N_16335);
nand U16558 (N_16558,N_16472,N_16463);
nand U16559 (N_16559,N_16366,N_16414);
and U16560 (N_16560,N_16330,N_16410);
and U16561 (N_16561,N_16363,N_16320);
nand U16562 (N_16562,N_16353,N_16435);
nor U16563 (N_16563,N_16322,N_16423);
xnor U16564 (N_16564,N_16395,N_16351);
nor U16565 (N_16565,N_16454,N_16404);
nor U16566 (N_16566,N_16397,N_16420);
nand U16567 (N_16567,N_16444,N_16374);
nand U16568 (N_16568,N_16371,N_16457);
and U16569 (N_16569,N_16339,N_16455);
nor U16570 (N_16570,N_16427,N_16395);
xnor U16571 (N_16571,N_16342,N_16473);
nand U16572 (N_16572,N_16347,N_16450);
and U16573 (N_16573,N_16442,N_16434);
and U16574 (N_16574,N_16336,N_16408);
and U16575 (N_16575,N_16331,N_16343);
and U16576 (N_16576,N_16365,N_16461);
nand U16577 (N_16577,N_16351,N_16386);
or U16578 (N_16578,N_16376,N_16410);
xnor U16579 (N_16579,N_16384,N_16420);
nand U16580 (N_16580,N_16415,N_16454);
nor U16581 (N_16581,N_16373,N_16402);
nand U16582 (N_16582,N_16442,N_16346);
xor U16583 (N_16583,N_16464,N_16357);
nand U16584 (N_16584,N_16406,N_16324);
or U16585 (N_16585,N_16441,N_16440);
and U16586 (N_16586,N_16394,N_16385);
and U16587 (N_16587,N_16384,N_16453);
nand U16588 (N_16588,N_16471,N_16367);
or U16589 (N_16589,N_16337,N_16398);
or U16590 (N_16590,N_16388,N_16477);
and U16591 (N_16591,N_16470,N_16476);
and U16592 (N_16592,N_16445,N_16405);
or U16593 (N_16593,N_16392,N_16330);
nand U16594 (N_16594,N_16393,N_16456);
and U16595 (N_16595,N_16472,N_16398);
nand U16596 (N_16596,N_16401,N_16456);
and U16597 (N_16597,N_16475,N_16419);
nand U16598 (N_16598,N_16392,N_16366);
xor U16599 (N_16599,N_16476,N_16389);
and U16600 (N_16600,N_16383,N_16427);
xnor U16601 (N_16601,N_16394,N_16393);
xnor U16602 (N_16602,N_16457,N_16411);
and U16603 (N_16603,N_16409,N_16325);
nor U16604 (N_16604,N_16359,N_16383);
nand U16605 (N_16605,N_16404,N_16370);
or U16606 (N_16606,N_16413,N_16418);
or U16607 (N_16607,N_16377,N_16430);
xnor U16608 (N_16608,N_16421,N_16325);
or U16609 (N_16609,N_16355,N_16449);
or U16610 (N_16610,N_16461,N_16450);
or U16611 (N_16611,N_16401,N_16454);
nor U16612 (N_16612,N_16478,N_16392);
and U16613 (N_16613,N_16394,N_16392);
or U16614 (N_16614,N_16428,N_16367);
or U16615 (N_16615,N_16428,N_16353);
and U16616 (N_16616,N_16368,N_16402);
nand U16617 (N_16617,N_16386,N_16382);
and U16618 (N_16618,N_16471,N_16475);
nand U16619 (N_16619,N_16325,N_16423);
or U16620 (N_16620,N_16444,N_16426);
nor U16621 (N_16621,N_16413,N_16338);
or U16622 (N_16622,N_16464,N_16355);
or U16623 (N_16623,N_16376,N_16388);
nand U16624 (N_16624,N_16405,N_16458);
xnor U16625 (N_16625,N_16358,N_16337);
xor U16626 (N_16626,N_16478,N_16378);
or U16627 (N_16627,N_16431,N_16406);
nor U16628 (N_16628,N_16369,N_16324);
nor U16629 (N_16629,N_16347,N_16453);
xor U16630 (N_16630,N_16328,N_16447);
and U16631 (N_16631,N_16360,N_16390);
or U16632 (N_16632,N_16393,N_16339);
and U16633 (N_16633,N_16462,N_16334);
xnor U16634 (N_16634,N_16465,N_16330);
xnor U16635 (N_16635,N_16446,N_16469);
or U16636 (N_16636,N_16321,N_16325);
nor U16637 (N_16637,N_16346,N_16429);
nor U16638 (N_16638,N_16471,N_16398);
nand U16639 (N_16639,N_16392,N_16361);
nand U16640 (N_16640,N_16561,N_16630);
or U16641 (N_16641,N_16581,N_16598);
and U16642 (N_16642,N_16636,N_16519);
and U16643 (N_16643,N_16544,N_16570);
and U16644 (N_16644,N_16555,N_16596);
nor U16645 (N_16645,N_16534,N_16616);
nor U16646 (N_16646,N_16484,N_16588);
nand U16647 (N_16647,N_16597,N_16582);
nand U16648 (N_16648,N_16614,N_16559);
nor U16649 (N_16649,N_16612,N_16495);
or U16650 (N_16650,N_16606,N_16575);
or U16651 (N_16651,N_16504,N_16517);
nor U16652 (N_16652,N_16620,N_16590);
and U16653 (N_16653,N_16633,N_16618);
and U16654 (N_16654,N_16586,N_16506);
or U16655 (N_16655,N_16508,N_16584);
xnor U16656 (N_16656,N_16605,N_16615);
or U16657 (N_16657,N_16494,N_16545);
or U16658 (N_16658,N_16591,N_16603);
or U16659 (N_16659,N_16513,N_16604);
xor U16660 (N_16660,N_16485,N_16592);
and U16661 (N_16661,N_16580,N_16543);
nand U16662 (N_16662,N_16481,N_16623);
nand U16663 (N_16663,N_16556,N_16548);
nor U16664 (N_16664,N_16549,N_16602);
xnor U16665 (N_16665,N_16585,N_16574);
nand U16666 (N_16666,N_16516,N_16629);
and U16667 (N_16667,N_16594,N_16572);
nand U16668 (N_16668,N_16530,N_16483);
xor U16669 (N_16669,N_16566,N_16510);
and U16670 (N_16670,N_16635,N_16537);
xnor U16671 (N_16671,N_16627,N_16512);
or U16672 (N_16672,N_16608,N_16610);
xor U16673 (N_16673,N_16571,N_16533);
nand U16674 (N_16674,N_16540,N_16529);
or U16675 (N_16675,N_16563,N_16526);
xor U16676 (N_16676,N_16499,N_16554);
and U16677 (N_16677,N_16500,N_16490);
xor U16678 (N_16678,N_16624,N_16619);
xor U16679 (N_16679,N_16511,N_16520);
or U16680 (N_16680,N_16522,N_16501);
xnor U16681 (N_16681,N_16507,N_16541);
nand U16682 (N_16682,N_16539,N_16637);
nor U16683 (N_16683,N_16480,N_16493);
or U16684 (N_16684,N_16532,N_16577);
xor U16685 (N_16685,N_16565,N_16509);
nor U16686 (N_16686,N_16491,N_16560);
or U16687 (N_16687,N_16515,N_16521);
and U16688 (N_16688,N_16503,N_16492);
nor U16689 (N_16689,N_16578,N_16626);
or U16690 (N_16690,N_16558,N_16525);
or U16691 (N_16691,N_16625,N_16583);
and U16692 (N_16692,N_16498,N_16488);
nand U16693 (N_16693,N_16552,N_16639);
xnor U16694 (N_16694,N_16564,N_16576);
xor U16695 (N_16695,N_16617,N_16514);
nor U16696 (N_16696,N_16579,N_16601);
or U16697 (N_16697,N_16613,N_16611);
nand U16698 (N_16698,N_16551,N_16593);
xor U16699 (N_16699,N_16568,N_16587);
and U16700 (N_16700,N_16524,N_16589);
nand U16701 (N_16701,N_16538,N_16631);
or U16702 (N_16702,N_16609,N_16595);
xnor U16703 (N_16703,N_16567,N_16535);
nor U16704 (N_16704,N_16573,N_16622);
or U16705 (N_16705,N_16628,N_16600);
and U16706 (N_16706,N_16562,N_16527);
nor U16707 (N_16707,N_16542,N_16528);
xnor U16708 (N_16708,N_16557,N_16482);
xor U16709 (N_16709,N_16634,N_16496);
nor U16710 (N_16710,N_16621,N_16638);
or U16711 (N_16711,N_16547,N_16531);
and U16712 (N_16712,N_16546,N_16505);
nand U16713 (N_16713,N_16553,N_16550);
nand U16714 (N_16714,N_16518,N_16536);
and U16715 (N_16715,N_16607,N_16487);
or U16716 (N_16716,N_16497,N_16489);
or U16717 (N_16717,N_16599,N_16632);
or U16718 (N_16718,N_16502,N_16569);
and U16719 (N_16719,N_16486,N_16523);
xnor U16720 (N_16720,N_16508,N_16635);
xnor U16721 (N_16721,N_16488,N_16482);
or U16722 (N_16722,N_16619,N_16627);
or U16723 (N_16723,N_16502,N_16511);
nand U16724 (N_16724,N_16634,N_16504);
xor U16725 (N_16725,N_16547,N_16572);
and U16726 (N_16726,N_16530,N_16480);
and U16727 (N_16727,N_16604,N_16570);
and U16728 (N_16728,N_16497,N_16578);
xnor U16729 (N_16729,N_16591,N_16495);
xnor U16730 (N_16730,N_16514,N_16569);
xor U16731 (N_16731,N_16588,N_16525);
nor U16732 (N_16732,N_16515,N_16628);
and U16733 (N_16733,N_16507,N_16494);
or U16734 (N_16734,N_16614,N_16553);
nor U16735 (N_16735,N_16492,N_16509);
or U16736 (N_16736,N_16638,N_16614);
nor U16737 (N_16737,N_16549,N_16488);
or U16738 (N_16738,N_16533,N_16491);
nor U16739 (N_16739,N_16522,N_16520);
nor U16740 (N_16740,N_16577,N_16531);
or U16741 (N_16741,N_16598,N_16516);
nand U16742 (N_16742,N_16505,N_16606);
nand U16743 (N_16743,N_16566,N_16558);
xnor U16744 (N_16744,N_16587,N_16629);
nor U16745 (N_16745,N_16550,N_16594);
nor U16746 (N_16746,N_16509,N_16607);
nor U16747 (N_16747,N_16626,N_16503);
or U16748 (N_16748,N_16486,N_16585);
xnor U16749 (N_16749,N_16536,N_16555);
and U16750 (N_16750,N_16634,N_16568);
or U16751 (N_16751,N_16513,N_16564);
xor U16752 (N_16752,N_16636,N_16534);
or U16753 (N_16753,N_16483,N_16496);
xnor U16754 (N_16754,N_16618,N_16571);
and U16755 (N_16755,N_16559,N_16627);
xnor U16756 (N_16756,N_16578,N_16491);
nor U16757 (N_16757,N_16584,N_16632);
nor U16758 (N_16758,N_16607,N_16533);
nand U16759 (N_16759,N_16586,N_16582);
and U16760 (N_16760,N_16615,N_16483);
nand U16761 (N_16761,N_16599,N_16567);
nor U16762 (N_16762,N_16494,N_16483);
xnor U16763 (N_16763,N_16588,N_16570);
nor U16764 (N_16764,N_16592,N_16582);
nand U16765 (N_16765,N_16633,N_16630);
nand U16766 (N_16766,N_16560,N_16582);
and U16767 (N_16767,N_16581,N_16521);
nor U16768 (N_16768,N_16591,N_16634);
nand U16769 (N_16769,N_16589,N_16488);
and U16770 (N_16770,N_16554,N_16480);
nor U16771 (N_16771,N_16639,N_16621);
and U16772 (N_16772,N_16542,N_16525);
xnor U16773 (N_16773,N_16526,N_16482);
or U16774 (N_16774,N_16494,N_16603);
and U16775 (N_16775,N_16583,N_16506);
nand U16776 (N_16776,N_16512,N_16589);
xor U16777 (N_16777,N_16484,N_16604);
nor U16778 (N_16778,N_16537,N_16586);
nand U16779 (N_16779,N_16557,N_16628);
or U16780 (N_16780,N_16560,N_16639);
nand U16781 (N_16781,N_16583,N_16517);
nor U16782 (N_16782,N_16575,N_16565);
nor U16783 (N_16783,N_16546,N_16636);
or U16784 (N_16784,N_16550,N_16519);
and U16785 (N_16785,N_16596,N_16573);
and U16786 (N_16786,N_16618,N_16631);
nand U16787 (N_16787,N_16591,N_16579);
or U16788 (N_16788,N_16487,N_16589);
and U16789 (N_16789,N_16487,N_16570);
nand U16790 (N_16790,N_16547,N_16542);
xor U16791 (N_16791,N_16569,N_16487);
xnor U16792 (N_16792,N_16564,N_16610);
or U16793 (N_16793,N_16587,N_16482);
nor U16794 (N_16794,N_16628,N_16553);
nand U16795 (N_16795,N_16541,N_16515);
nor U16796 (N_16796,N_16563,N_16633);
nand U16797 (N_16797,N_16600,N_16504);
and U16798 (N_16798,N_16539,N_16603);
and U16799 (N_16799,N_16635,N_16489);
xnor U16800 (N_16800,N_16722,N_16688);
nor U16801 (N_16801,N_16719,N_16788);
or U16802 (N_16802,N_16693,N_16721);
nor U16803 (N_16803,N_16759,N_16662);
nor U16804 (N_16804,N_16683,N_16757);
or U16805 (N_16805,N_16735,N_16725);
xnor U16806 (N_16806,N_16644,N_16792);
and U16807 (N_16807,N_16713,N_16746);
xnor U16808 (N_16808,N_16652,N_16727);
nor U16809 (N_16809,N_16769,N_16656);
and U16810 (N_16810,N_16730,N_16741);
xnor U16811 (N_16811,N_16655,N_16772);
and U16812 (N_16812,N_16716,N_16763);
xor U16813 (N_16813,N_16791,N_16703);
nor U16814 (N_16814,N_16657,N_16689);
and U16815 (N_16815,N_16756,N_16782);
xnor U16816 (N_16816,N_16723,N_16720);
xnor U16817 (N_16817,N_16715,N_16681);
nand U16818 (N_16818,N_16777,N_16712);
or U16819 (N_16819,N_16669,N_16781);
xnor U16820 (N_16820,N_16642,N_16748);
or U16821 (N_16821,N_16768,N_16761);
or U16822 (N_16822,N_16790,N_16754);
or U16823 (N_16823,N_16700,N_16685);
nand U16824 (N_16824,N_16706,N_16786);
and U16825 (N_16825,N_16701,N_16653);
nor U16826 (N_16826,N_16799,N_16651);
nand U16827 (N_16827,N_16664,N_16784);
nand U16828 (N_16828,N_16677,N_16778);
nand U16829 (N_16829,N_16661,N_16771);
and U16830 (N_16830,N_16707,N_16666);
and U16831 (N_16831,N_16711,N_16663);
xnor U16832 (N_16832,N_16766,N_16789);
or U16833 (N_16833,N_16702,N_16753);
and U16834 (N_16834,N_16783,N_16697);
and U16835 (N_16835,N_16705,N_16650);
nor U16836 (N_16836,N_16647,N_16646);
nand U16837 (N_16837,N_16734,N_16728);
or U16838 (N_16838,N_16641,N_16776);
and U16839 (N_16839,N_16718,N_16667);
and U16840 (N_16840,N_16747,N_16724);
or U16841 (N_16841,N_16774,N_16649);
xor U16842 (N_16842,N_16672,N_16668);
or U16843 (N_16843,N_16744,N_16670);
nand U16844 (N_16844,N_16658,N_16749);
nand U16845 (N_16845,N_16796,N_16704);
nand U16846 (N_16846,N_16676,N_16797);
and U16847 (N_16847,N_16793,N_16764);
nand U16848 (N_16848,N_16737,N_16698);
nor U16849 (N_16849,N_16648,N_16709);
or U16850 (N_16850,N_16751,N_16742);
and U16851 (N_16851,N_16645,N_16752);
nand U16852 (N_16852,N_16695,N_16640);
xnor U16853 (N_16853,N_16692,N_16736);
or U16854 (N_16854,N_16659,N_16767);
and U16855 (N_16855,N_16665,N_16729);
nor U16856 (N_16856,N_16739,N_16750);
nand U16857 (N_16857,N_16762,N_16795);
and U16858 (N_16858,N_16743,N_16680);
nand U16859 (N_16859,N_16765,N_16673);
or U16860 (N_16860,N_16745,N_16732);
xor U16861 (N_16861,N_16733,N_16699);
xnor U16862 (N_16862,N_16780,N_16770);
nand U16863 (N_16863,N_16654,N_16708);
xor U16864 (N_16864,N_16717,N_16775);
xnor U16865 (N_16865,N_16758,N_16760);
and U16866 (N_16866,N_16678,N_16671);
nand U16867 (N_16867,N_16696,N_16691);
or U16868 (N_16868,N_16785,N_16679);
nor U16869 (N_16869,N_16779,N_16690);
nand U16870 (N_16870,N_16773,N_16674);
and U16871 (N_16871,N_16660,N_16687);
and U16872 (N_16872,N_16675,N_16643);
and U16873 (N_16873,N_16694,N_16740);
or U16874 (N_16874,N_16787,N_16794);
and U16875 (N_16875,N_16710,N_16731);
xnor U16876 (N_16876,N_16684,N_16738);
xor U16877 (N_16877,N_16682,N_16726);
or U16878 (N_16878,N_16755,N_16686);
or U16879 (N_16879,N_16798,N_16714);
and U16880 (N_16880,N_16767,N_16678);
nand U16881 (N_16881,N_16743,N_16739);
and U16882 (N_16882,N_16675,N_16724);
xor U16883 (N_16883,N_16641,N_16731);
nand U16884 (N_16884,N_16683,N_16765);
nand U16885 (N_16885,N_16767,N_16754);
xor U16886 (N_16886,N_16790,N_16737);
nor U16887 (N_16887,N_16761,N_16707);
xnor U16888 (N_16888,N_16693,N_16754);
or U16889 (N_16889,N_16695,N_16760);
nor U16890 (N_16890,N_16670,N_16712);
nand U16891 (N_16891,N_16708,N_16702);
or U16892 (N_16892,N_16790,N_16701);
nand U16893 (N_16893,N_16768,N_16643);
xnor U16894 (N_16894,N_16693,N_16684);
nor U16895 (N_16895,N_16723,N_16758);
xnor U16896 (N_16896,N_16670,N_16753);
xnor U16897 (N_16897,N_16720,N_16706);
nand U16898 (N_16898,N_16704,N_16665);
nand U16899 (N_16899,N_16674,N_16718);
and U16900 (N_16900,N_16791,N_16670);
or U16901 (N_16901,N_16779,N_16737);
or U16902 (N_16902,N_16773,N_16681);
and U16903 (N_16903,N_16721,N_16788);
and U16904 (N_16904,N_16641,N_16648);
xor U16905 (N_16905,N_16649,N_16797);
nand U16906 (N_16906,N_16782,N_16742);
and U16907 (N_16907,N_16701,N_16718);
xor U16908 (N_16908,N_16785,N_16666);
nor U16909 (N_16909,N_16771,N_16795);
nand U16910 (N_16910,N_16694,N_16754);
and U16911 (N_16911,N_16740,N_16703);
nor U16912 (N_16912,N_16647,N_16712);
xor U16913 (N_16913,N_16704,N_16737);
nor U16914 (N_16914,N_16687,N_16735);
xor U16915 (N_16915,N_16664,N_16657);
xor U16916 (N_16916,N_16798,N_16774);
nor U16917 (N_16917,N_16746,N_16717);
nand U16918 (N_16918,N_16749,N_16757);
and U16919 (N_16919,N_16746,N_16760);
or U16920 (N_16920,N_16787,N_16700);
and U16921 (N_16921,N_16645,N_16682);
and U16922 (N_16922,N_16661,N_16797);
nand U16923 (N_16923,N_16749,N_16799);
or U16924 (N_16924,N_16679,N_16646);
and U16925 (N_16925,N_16655,N_16689);
xor U16926 (N_16926,N_16655,N_16764);
nand U16927 (N_16927,N_16773,N_16736);
nand U16928 (N_16928,N_16782,N_16675);
or U16929 (N_16929,N_16682,N_16762);
xnor U16930 (N_16930,N_16659,N_16768);
xnor U16931 (N_16931,N_16765,N_16719);
or U16932 (N_16932,N_16675,N_16706);
and U16933 (N_16933,N_16646,N_16750);
or U16934 (N_16934,N_16676,N_16674);
nand U16935 (N_16935,N_16669,N_16672);
nand U16936 (N_16936,N_16751,N_16656);
nand U16937 (N_16937,N_16711,N_16760);
nor U16938 (N_16938,N_16785,N_16677);
and U16939 (N_16939,N_16696,N_16726);
or U16940 (N_16940,N_16728,N_16697);
nand U16941 (N_16941,N_16739,N_16773);
nor U16942 (N_16942,N_16795,N_16640);
xor U16943 (N_16943,N_16656,N_16661);
and U16944 (N_16944,N_16754,N_16781);
nand U16945 (N_16945,N_16790,N_16780);
or U16946 (N_16946,N_16646,N_16712);
nor U16947 (N_16947,N_16654,N_16760);
nor U16948 (N_16948,N_16784,N_16675);
and U16949 (N_16949,N_16689,N_16659);
nand U16950 (N_16950,N_16708,N_16759);
nand U16951 (N_16951,N_16760,N_16673);
or U16952 (N_16952,N_16738,N_16694);
xor U16953 (N_16953,N_16764,N_16710);
xnor U16954 (N_16954,N_16697,N_16759);
nand U16955 (N_16955,N_16722,N_16698);
xor U16956 (N_16956,N_16793,N_16761);
nor U16957 (N_16957,N_16642,N_16735);
and U16958 (N_16958,N_16774,N_16690);
nor U16959 (N_16959,N_16680,N_16651);
or U16960 (N_16960,N_16871,N_16861);
nand U16961 (N_16961,N_16914,N_16919);
nor U16962 (N_16962,N_16959,N_16853);
nor U16963 (N_16963,N_16851,N_16852);
xor U16964 (N_16964,N_16915,N_16907);
nor U16965 (N_16965,N_16880,N_16931);
or U16966 (N_16966,N_16815,N_16885);
or U16967 (N_16967,N_16912,N_16804);
nand U16968 (N_16968,N_16828,N_16820);
nand U16969 (N_16969,N_16857,N_16850);
xnor U16970 (N_16970,N_16887,N_16882);
nand U16971 (N_16971,N_16881,N_16941);
and U16972 (N_16972,N_16903,N_16913);
or U16973 (N_16973,N_16842,N_16895);
and U16974 (N_16974,N_16872,N_16908);
and U16975 (N_16975,N_16856,N_16922);
nand U16976 (N_16976,N_16958,N_16834);
or U16977 (N_16977,N_16848,N_16940);
xor U16978 (N_16978,N_16800,N_16935);
xor U16979 (N_16979,N_16902,N_16909);
xor U16980 (N_16980,N_16899,N_16901);
nor U16981 (N_16981,N_16827,N_16845);
nor U16982 (N_16982,N_16938,N_16832);
nor U16983 (N_16983,N_16929,N_16900);
nand U16984 (N_16984,N_16926,N_16841);
nand U16985 (N_16985,N_16890,N_16886);
or U16986 (N_16986,N_16911,N_16803);
nor U16987 (N_16987,N_16835,N_16936);
xnor U16988 (N_16988,N_16859,N_16821);
xor U16989 (N_16989,N_16802,N_16870);
nand U16990 (N_16990,N_16840,N_16823);
or U16991 (N_16991,N_16874,N_16818);
nand U16992 (N_16992,N_16934,N_16930);
or U16993 (N_16993,N_16817,N_16910);
and U16994 (N_16994,N_16932,N_16819);
nand U16995 (N_16995,N_16809,N_16904);
xor U16996 (N_16996,N_16948,N_16839);
nor U16997 (N_16997,N_16925,N_16924);
xor U16998 (N_16998,N_16893,N_16862);
nand U16999 (N_16999,N_16928,N_16906);
nand U17000 (N_17000,N_16877,N_16825);
xor U17001 (N_17001,N_16891,N_16955);
nor U17002 (N_17002,N_16898,N_16843);
nand U17003 (N_17003,N_16855,N_16918);
xor U17004 (N_17004,N_16943,N_16816);
or U17005 (N_17005,N_16829,N_16946);
xnor U17006 (N_17006,N_16863,N_16812);
xor U17007 (N_17007,N_16879,N_16814);
nand U17008 (N_17008,N_16854,N_16831);
or U17009 (N_17009,N_16866,N_16865);
nand U17010 (N_17010,N_16933,N_16939);
or U17011 (N_17011,N_16883,N_16951);
and U17012 (N_17012,N_16807,N_16847);
nand U17013 (N_17013,N_16923,N_16806);
and U17014 (N_17014,N_16949,N_16921);
or U17015 (N_17015,N_16838,N_16822);
nor U17016 (N_17016,N_16888,N_16876);
and U17017 (N_17017,N_16927,N_16889);
and U17018 (N_17018,N_16858,N_16869);
xnor U17019 (N_17019,N_16896,N_16813);
or U17020 (N_17020,N_16867,N_16916);
nand U17021 (N_17021,N_16894,N_16937);
nand U17022 (N_17022,N_16833,N_16873);
nor U17023 (N_17023,N_16810,N_16884);
or U17024 (N_17024,N_16950,N_16956);
xnor U17025 (N_17025,N_16875,N_16897);
or U17026 (N_17026,N_16878,N_16892);
xor U17027 (N_17027,N_16837,N_16811);
xnor U17028 (N_17028,N_16824,N_16944);
and U17029 (N_17029,N_16920,N_16917);
xor U17030 (N_17030,N_16942,N_16846);
and U17031 (N_17031,N_16947,N_16945);
or U17032 (N_17032,N_16844,N_16836);
or U17033 (N_17033,N_16953,N_16808);
nor U17034 (N_17034,N_16830,N_16860);
xor U17035 (N_17035,N_16868,N_16849);
and U17036 (N_17036,N_16864,N_16905);
xor U17037 (N_17037,N_16957,N_16954);
nor U17038 (N_17038,N_16952,N_16826);
nand U17039 (N_17039,N_16801,N_16805);
or U17040 (N_17040,N_16830,N_16958);
xnor U17041 (N_17041,N_16820,N_16823);
and U17042 (N_17042,N_16953,N_16858);
nor U17043 (N_17043,N_16913,N_16879);
nand U17044 (N_17044,N_16899,N_16930);
or U17045 (N_17045,N_16864,N_16948);
and U17046 (N_17046,N_16848,N_16907);
and U17047 (N_17047,N_16881,N_16928);
nor U17048 (N_17048,N_16918,N_16811);
and U17049 (N_17049,N_16857,N_16945);
nand U17050 (N_17050,N_16827,N_16955);
or U17051 (N_17051,N_16865,N_16873);
xnor U17052 (N_17052,N_16868,N_16854);
nor U17053 (N_17053,N_16830,N_16836);
or U17054 (N_17054,N_16810,N_16824);
nand U17055 (N_17055,N_16894,N_16801);
or U17056 (N_17056,N_16874,N_16926);
xor U17057 (N_17057,N_16953,N_16920);
and U17058 (N_17058,N_16811,N_16908);
nand U17059 (N_17059,N_16820,N_16940);
or U17060 (N_17060,N_16918,N_16952);
nand U17061 (N_17061,N_16855,N_16902);
nand U17062 (N_17062,N_16831,N_16926);
nand U17063 (N_17063,N_16914,N_16804);
and U17064 (N_17064,N_16893,N_16834);
xnor U17065 (N_17065,N_16867,N_16938);
nand U17066 (N_17066,N_16826,N_16860);
and U17067 (N_17067,N_16812,N_16859);
xnor U17068 (N_17068,N_16874,N_16949);
and U17069 (N_17069,N_16917,N_16819);
and U17070 (N_17070,N_16829,N_16906);
and U17071 (N_17071,N_16871,N_16912);
nand U17072 (N_17072,N_16866,N_16871);
and U17073 (N_17073,N_16867,N_16801);
xor U17074 (N_17074,N_16919,N_16956);
or U17075 (N_17075,N_16948,N_16805);
xnor U17076 (N_17076,N_16852,N_16906);
or U17077 (N_17077,N_16872,N_16942);
or U17078 (N_17078,N_16849,N_16834);
or U17079 (N_17079,N_16813,N_16824);
nor U17080 (N_17080,N_16898,N_16893);
xnor U17081 (N_17081,N_16945,N_16924);
nor U17082 (N_17082,N_16857,N_16821);
nand U17083 (N_17083,N_16882,N_16910);
xnor U17084 (N_17084,N_16819,N_16803);
or U17085 (N_17085,N_16904,N_16829);
nor U17086 (N_17086,N_16932,N_16873);
nand U17087 (N_17087,N_16950,N_16875);
nand U17088 (N_17088,N_16925,N_16854);
nor U17089 (N_17089,N_16830,N_16943);
xnor U17090 (N_17090,N_16848,N_16910);
nand U17091 (N_17091,N_16922,N_16822);
xor U17092 (N_17092,N_16844,N_16833);
and U17093 (N_17093,N_16813,N_16830);
xor U17094 (N_17094,N_16889,N_16821);
nor U17095 (N_17095,N_16920,N_16873);
xor U17096 (N_17096,N_16838,N_16917);
nor U17097 (N_17097,N_16939,N_16888);
and U17098 (N_17098,N_16837,N_16825);
nor U17099 (N_17099,N_16894,N_16852);
or U17100 (N_17100,N_16863,N_16848);
nand U17101 (N_17101,N_16914,N_16882);
xnor U17102 (N_17102,N_16924,N_16889);
or U17103 (N_17103,N_16865,N_16811);
and U17104 (N_17104,N_16901,N_16822);
nor U17105 (N_17105,N_16905,N_16836);
and U17106 (N_17106,N_16938,N_16858);
nor U17107 (N_17107,N_16830,N_16913);
nand U17108 (N_17108,N_16958,N_16901);
and U17109 (N_17109,N_16928,N_16857);
or U17110 (N_17110,N_16881,N_16867);
nor U17111 (N_17111,N_16807,N_16854);
and U17112 (N_17112,N_16896,N_16922);
and U17113 (N_17113,N_16955,N_16832);
and U17114 (N_17114,N_16884,N_16926);
and U17115 (N_17115,N_16920,N_16854);
nor U17116 (N_17116,N_16831,N_16932);
xnor U17117 (N_17117,N_16944,N_16911);
nor U17118 (N_17118,N_16829,N_16845);
nand U17119 (N_17119,N_16898,N_16886);
xor U17120 (N_17120,N_16997,N_16987);
xor U17121 (N_17121,N_16986,N_17088);
nor U17122 (N_17122,N_17073,N_17104);
or U17123 (N_17123,N_17110,N_17014);
and U17124 (N_17124,N_16994,N_16979);
or U17125 (N_17125,N_16985,N_17002);
nor U17126 (N_17126,N_17067,N_17048);
or U17127 (N_17127,N_16972,N_17052);
nand U17128 (N_17128,N_17012,N_17107);
and U17129 (N_17129,N_17068,N_17082);
and U17130 (N_17130,N_17035,N_16981);
and U17131 (N_17131,N_16984,N_16998);
and U17132 (N_17132,N_17023,N_17096);
and U17133 (N_17133,N_17029,N_17094);
and U17134 (N_17134,N_17026,N_17041);
nand U17135 (N_17135,N_17013,N_17076);
and U17136 (N_17136,N_17106,N_17060);
and U17137 (N_17137,N_16999,N_17118);
nand U17138 (N_17138,N_16968,N_17000);
and U17139 (N_17139,N_17022,N_17007);
and U17140 (N_17140,N_16976,N_17072);
and U17141 (N_17141,N_16963,N_16961);
or U17142 (N_17142,N_16995,N_17049);
xor U17143 (N_17143,N_17116,N_17086);
or U17144 (N_17144,N_17031,N_17042);
xor U17145 (N_17145,N_17016,N_17055);
nand U17146 (N_17146,N_17114,N_16975);
or U17147 (N_17147,N_17040,N_16973);
and U17148 (N_17148,N_17091,N_17115);
xor U17149 (N_17149,N_17080,N_17044);
or U17150 (N_17150,N_17100,N_16982);
nand U17151 (N_17151,N_17021,N_17066);
xor U17152 (N_17152,N_17101,N_17085);
or U17153 (N_17153,N_16960,N_16964);
nand U17154 (N_17154,N_17050,N_16983);
or U17155 (N_17155,N_17051,N_17005);
and U17156 (N_17156,N_17081,N_16970);
xnor U17157 (N_17157,N_17090,N_17036);
nand U17158 (N_17158,N_16980,N_17071);
and U17159 (N_17159,N_17010,N_16962);
xnor U17160 (N_17160,N_17093,N_17117);
xnor U17161 (N_17161,N_16966,N_17006);
or U17162 (N_17162,N_17039,N_16990);
xnor U17163 (N_17163,N_17112,N_17105);
or U17164 (N_17164,N_17074,N_17038);
or U17165 (N_17165,N_17069,N_17103);
xnor U17166 (N_17166,N_17009,N_16978);
nand U17167 (N_17167,N_17062,N_16967);
or U17168 (N_17168,N_16965,N_17054);
or U17169 (N_17169,N_16977,N_16969);
and U17170 (N_17170,N_17043,N_17059);
nand U17171 (N_17171,N_17056,N_17113);
nand U17172 (N_17172,N_17075,N_17015);
nor U17173 (N_17173,N_17097,N_17092);
xor U17174 (N_17174,N_17017,N_17084);
xor U17175 (N_17175,N_17111,N_16988);
nor U17176 (N_17176,N_17070,N_16993);
and U17177 (N_17177,N_17078,N_16991);
or U17178 (N_17178,N_17025,N_17030);
nor U17179 (N_17179,N_16971,N_17047);
and U17180 (N_17180,N_17102,N_17003);
xor U17181 (N_17181,N_17057,N_17001);
and U17182 (N_17182,N_17028,N_17004);
nor U17183 (N_17183,N_17032,N_16996);
xnor U17184 (N_17184,N_17011,N_17033);
nand U17185 (N_17185,N_17034,N_17108);
nor U17186 (N_17186,N_17095,N_17109);
nand U17187 (N_17187,N_17064,N_17019);
and U17188 (N_17188,N_16974,N_17053);
nand U17189 (N_17189,N_17061,N_17018);
xor U17190 (N_17190,N_17083,N_17079);
nand U17191 (N_17191,N_17027,N_16992);
nand U17192 (N_17192,N_17065,N_17087);
nand U17193 (N_17193,N_17058,N_17024);
nand U17194 (N_17194,N_17089,N_17020);
nor U17195 (N_17195,N_16989,N_17063);
nor U17196 (N_17196,N_17045,N_17099);
nand U17197 (N_17197,N_17046,N_17037);
nor U17198 (N_17198,N_17098,N_17119);
nand U17199 (N_17199,N_17077,N_17008);
and U17200 (N_17200,N_17044,N_17019);
nand U17201 (N_17201,N_17077,N_17020);
nand U17202 (N_17202,N_17053,N_17030);
or U17203 (N_17203,N_17053,N_17037);
nand U17204 (N_17204,N_17009,N_16963);
nor U17205 (N_17205,N_16991,N_17098);
or U17206 (N_17206,N_16990,N_17078);
and U17207 (N_17207,N_16992,N_17069);
and U17208 (N_17208,N_17066,N_17024);
nand U17209 (N_17209,N_17018,N_16964);
xor U17210 (N_17210,N_17079,N_17049);
or U17211 (N_17211,N_17072,N_17049);
xor U17212 (N_17212,N_17057,N_16984);
nand U17213 (N_17213,N_17103,N_17061);
nor U17214 (N_17214,N_16999,N_17015);
or U17215 (N_17215,N_17117,N_16965);
xor U17216 (N_17216,N_17023,N_17076);
and U17217 (N_17217,N_16973,N_16971);
and U17218 (N_17218,N_16981,N_17112);
nand U17219 (N_17219,N_17016,N_17114);
nand U17220 (N_17220,N_17023,N_17017);
xor U17221 (N_17221,N_17049,N_17003);
xnor U17222 (N_17222,N_16997,N_17052);
nor U17223 (N_17223,N_17068,N_17073);
nor U17224 (N_17224,N_17098,N_17083);
and U17225 (N_17225,N_17005,N_17037);
nor U17226 (N_17226,N_16968,N_16997);
xnor U17227 (N_17227,N_17078,N_16989);
xor U17228 (N_17228,N_16998,N_17109);
nand U17229 (N_17229,N_16988,N_17102);
nor U17230 (N_17230,N_16991,N_17033);
and U17231 (N_17231,N_17093,N_17119);
nand U17232 (N_17232,N_17083,N_17059);
or U17233 (N_17233,N_17063,N_16960);
nand U17234 (N_17234,N_17104,N_16972);
or U17235 (N_17235,N_17033,N_17100);
xnor U17236 (N_17236,N_17042,N_16996);
xnor U17237 (N_17237,N_16985,N_17008);
nand U17238 (N_17238,N_17093,N_17099);
nor U17239 (N_17239,N_16967,N_17028);
and U17240 (N_17240,N_17020,N_16970);
nor U17241 (N_17241,N_17052,N_17026);
xor U17242 (N_17242,N_17066,N_17050);
xnor U17243 (N_17243,N_17054,N_17039);
xnor U17244 (N_17244,N_16967,N_16960);
xnor U17245 (N_17245,N_17073,N_17114);
nor U17246 (N_17246,N_16988,N_17064);
or U17247 (N_17247,N_16972,N_17094);
and U17248 (N_17248,N_17072,N_17075);
nor U17249 (N_17249,N_17109,N_17119);
and U17250 (N_17250,N_17096,N_16963);
and U17251 (N_17251,N_17022,N_17074);
or U17252 (N_17252,N_17064,N_17045);
or U17253 (N_17253,N_17092,N_17008);
and U17254 (N_17254,N_17103,N_16981);
xor U17255 (N_17255,N_17049,N_17088);
nor U17256 (N_17256,N_17114,N_17080);
and U17257 (N_17257,N_17075,N_17054);
xnor U17258 (N_17258,N_17046,N_16979);
and U17259 (N_17259,N_17087,N_16993);
nor U17260 (N_17260,N_16985,N_17086);
nand U17261 (N_17261,N_17092,N_17010);
nand U17262 (N_17262,N_16967,N_17006);
nand U17263 (N_17263,N_16988,N_17082);
xnor U17264 (N_17264,N_17027,N_17087);
xor U17265 (N_17265,N_17118,N_17063);
or U17266 (N_17266,N_16996,N_16989);
or U17267 (N_17267,N_17104,N_17077);
or U17268 (N_17268,N_16968,N_17094);
or U17269 (N_17269,N_16974,N_17088);
xor U17270 (N_17270,N_16975,N_17097);
nor U17271 (N_17271,N_16969,N_17031);
nand U17272 (N_17272,N_16985,N_16990);
nor U17273 (N_17273,N_17047,N_17078);
and U17274 (N_17274,N_17029,N_17015);
or U17275 (N_17275,N_17009,N_17091);
nor U17276 (N_17276,N_16964,N_17083);
nor U17277 (N_17277,N_17108,N_17112);
nor U17278 (N_17278,N_16976,N_16983);
nand U17279 (N_17279,N_17010,N_16966);
nor U17280 (N_17280,N_17127,N_17132);
nor U17281 (N_17281,N_17266,N_17172);
nor U17282 (N_17282,N_17145,N_17175);
or U17283 (N_17283,N_17203,N_17272);
nor U17284 (N_17284,N_17246,N_17277);
nand U17285 (N_17285,N_17155,N_17216);
nand U17286 (N_17286,N_17253,N_17279);
nor U17287 (N_17287,N_17170,N_17220);
nand U17288 (N_17288,N_17160,N_17213);
or U17289 (N_17289,N_17255,N_17163);
or U17290 (N_17290,N_17176,N_17259);
nor U17291 (N_17291,N_17248,N_17250);
nand U17292 (N_17292,N_17262,N_17256);
nand U17293 (N_17293,N_17240,N_17239);
and U17294 (N_17294,N_17217,N_17168);
nor U17295 (N_17295,N_17258,N_17171);
and U17296 (N_17296,N_17162,N_17201);
or U17297 (N_17297,N_17167,N_17235);
nor U17298 (N_17298,N_17243,N_17135);
nand U17299 (N_17299,N_17244,N_17183);
nand U17300 (N_17300,N_17234,N_17153);
xnor U17301 (N_17301,N_17249,N_17230);
nor U17302 (N_17302,N_17212,N_17194);
xnor U17303 (N_17303,N_17150,N_17267);
xnor U17304 (N_17304,N_17130,N_17156);
nand U17305 (N_17305,N_17174,N_17227);
xnor U17306 (N_17306,N_17133,N_17208);
and U17307 (N_17307,N_17157,N_17206);
and U17308 (N_17308,N_17238,N_17274);
xnor U17309 (N_17309,N_17236,N_17278);
and U17310 (N_17310,N_17179,N_17232);
or U17311 (N_17311,N_17173,N_17161);
and U17312 (N_17312,N_17148,N_17188);
and U17313 (N_17313,N_17146,N_17224);
nand U17314 (N_17314,N_17260,N_17120);
and U17315 (N_17315,N_17209,N_17191);
nor U17316 (N_17316,N_17257,N_17181);
xnor U17317 (N_17317,N_17143,N_17233);
xnor U17318 (N_17318,N_17214,N_17141);
xnor U17319 (N_17319,N_17159,N_17128);
nand U17320 (N_17320,N_17122,N_17166);
or U17321 (N_17321,N_17142,N_17187);
or U17322 (N_17322,N_17123,N_17237);
nand U17323 (N_17323,N_17198,N_17165);
and U17324 (N_17324,N_17226,N_17247);
xor U17325 (N_17325,N_17215,N_17164);
nor U17326 (N_17326,N_17180,N_17275);
nor U17327 (N_17327,N_17136,N_17154);
and U17328 (N_17328,N_17218,N_17152);
nor U17329 (N_17329,N_17270,N_17131);
and U17330 (N_17330,N_17178,N_17182);
nor U17331 (N_17331,N_17151,N_17222);
nand U17332 (N_17332,N_17190,N_17134);
nor U17333 (N_17333,N_17197,N_17139);
or U17334 (N_17334,N_17193,N_17125);
and U17335 (N_17335,N_17140,N_17137);
nand U17336 (N_17336,N_17254,N_17177);
nand U17337 (N_17337,N_17229,N_17268);
xor U17338 (N_17338,N_17231,N_17273);
nand U17339 (N_17339,N_17207,N_17200);
nor U17340 (N_17340,N_17202,N_17121);
nand U17341 (N_17341,N_17241,N_17204);
and U17342 (N_17342,N_17138,N_17263);
nand U17343 (N_17343,N_17169,N_17269);
or U17344 (N_17344,N_17252,N_17129);
xor U17345 (N_17345,N_17245,N_17219);
nand U17346 (N_17346,N_17144,N_17221);
or U17347 (N_17347,N_17210,N_17186);
nand U17348 (N_17348,N_17158,N_17196);
nor U17349 (N_17349,N_17185,N_17251);
or U17350 (N_17350,N_17265,N_17189);
nor U17351 (N_17351,N_17223,N_17126);
or U17352 (N_17352,N_17192,N_17261);
nor U17353 (N_17353,N_17124,N_17225);
nand U17354 (N_17354,N_17242,N_17205);
xnor U17355 (N_17355,N_17199,N_17195);
and U17356 (N_17356,N_17276,N_17149);
xor U17357 (N_17357,N_17264,N_17228);
xor U17358 (N_17358,N_17271,N_17184);
or U17359 (N_17359,N_17211,N_17147);
or U17360 (N_17360,N_17124,N_17193);
or U17361 (N_17361,N_17165,N_17240);
nor U17362 (N_17362,N_17267,N_17273);
and U17363 (N_17363,N_17142,N_17130);
and U17364 (N_17364,N_17155,N_17192);
and U17365 (N_17365,N_17195,N_17175);
nand U17366 (N_17366,N_17150,N_17154);
nand U17367 (N_17367,N_17189,N_17177);
xor U17368 (N_17368,N_17263,N_17121);
and U17369 (N_17369,N_17152,N_17261);
and U17370 (N_17370,N_17170,N_17128);
and U17371 (N_17371,N_17154,N_17172);
nor U17372 (N_17372,N_17240,N_17178);
and U17373 (N_17373,N_17266,N_17225);
and U17374 (N_17374,N_17195,N_17245);
or U17375 (N_17375,N_17262,N_17194);
or U17376 (N_17376,N_17132,N_17138);
and U17377 (N_17377,N_17135,N_17227);
nand U17378 (N_17378,N_17263,N_17134);
or U17379 (N_17379,N_17149,N_17172);
and U17380 (N_17380,N_17251,N_17159);
xnor U17381 (N_17381,N_17192,N_17278);
nor U17382 (N_17382,N_17173,N_17266);
or U17383 (N_17383,N_17121,N_17161);
nand U17384 (N_17384,N_17206,N_17155);
or U17385 (N_17385,N_17216,N_17268);
or U17386 (N_17386,N_17276,N_17147);
or U17387 (N_17387,N_17211,N_17197);
xor U17388 (N_17388,N_17136,N_17262);
nor U17389 (N_17389,N_17274,N_17257);
nor U17390 (N_17390,N_17192,N_17263);
nand U17391 (N_17391,N_17227,N_17177);
and U17392 (N_17392,N_17223,N_17136);
and U17393 (N_17393,N_17208,N_17260);
xnor U17394 (N_17394,N_17147,N_17251);
nand U17395 (N_17395,N_17207,N_17194);
xnor U17396 (N_17396,N_17212,N_17214);
nor U17397 (N_17397,N_17239,N_17184);
nor U17398 (N_17398,N_17244,N_17236);
or U17399 (N_17399,N_17165,N_17138);
and U17400 (N_17400,N_17226,N_17222);
and U17401 (N_17401,N_17262,N_17190);
or U17402 (N_17402,N_17142,N_17125);
nor U17403 (N_17403,N_17225,N_17125);
xnor U17404 (N_17404,N_17166,N_17221);
nor U17405 (N_17405,N_17129,N_17255);
or U17406 (N_17406,N_17140,N_17243);
or U17407 (N_17407,N_17276,N_17231);
nand U17408 (N_17408,N_17188,N_17220);
nand U17409 (N_17409,N_17136,N_17185);
and U17410 (N_17410,N_17268,N_17211);
or U17411 (N_17411,N_17255,N_17238);
nor U17412 (N_17412,N_17205,N_17276);
or U17413 (N_17413,N_17124,N_17168);
nand U17414 (N_17414,N_17187,N_17178);
nor U17415 (N_17415,N_17257,N_17202);
and U17416 (N_17416,N_17172,N_17215);
or U17417 (N_17417,N_17132,N_17226);
and U17418 (N_17418,N_17214,N_17268);
or U17419 (N_17419,N_17193,N_17128);
xnor U17420 (N_17420,N_17132,N_17267);
and U17421 (N_17421,N_17163,N_17203);
xnor U17422 (N_17422,N_17211,N_17138);
nor U17423 (N_17423,N_17192,N_17279);
xor U17424 (N_17424,N_17279,N_17197);
xnor U17425 (N_17425,N_17178,N_17214);
or U17426 (N_17426,N_17208,N_17247);
xnor U17427 (N_17427,N_17219,N_17121);
and U17428 (N_17428,N_17168,N_17250);
nor U17429 (N_17429,N_17160,N_17196);
and U17430 (N_17430,N_17142,N_17147);
nor U17431 (N_17431,N_17189,N_17140);
nor U17432 (N_17432,N_17238,N_17175);
or U17433 (N_17433,N_17238,N_17254);
xor U17434 (N_17434,N_17170,N_17200);
and U17435 (N_17435,N_17273,N_17227);
and U17436 (N_17436,N_17189,N_17180);
nor U17437 (N_17437,N_17151,N_17268);
nor U17438 (N_17438,N_17146,N_17261);
or U17439 (N_17439,N_17223,N_17159);
nand U17440 (N_17440,N_17350,N_17349);
nand U17441 (N_17441,N_17421,N_17282);
and U17442 (N_17442,N_17397,N_17373);
or U17443 (N_17443,N_17425,N_17291);
xnor U17444 (N_17444,N_17280,N_17384);
and U17445 (N_17445,N_17344,N_17402);
and U17446 (N_17446,N_17369,N_17365);
or U17447 (N_17447,N_17378,N_17375);
or U17448 (N_17448,N_17364,N_17394);
or U17449 (N_17449,N_17381,N_17360);
and U17450 (N_17450,N_17408,N_17393);
and U17451 (N_17451,N_17426,N_17376);
nor U17452 (N_17452,N_17374,N_17337);
or U17453 (N_17453,N_17347,N_17406);
nor U17454 (N_17454,N_17295,N_17331);
nor U17455 (N_17455,N_17314,N_17328);
and U17456 (N_17456,N_17323,N_17368);
xor U17457 (N_17457,N_17439,N_17405);
nand U17458 (N_17458,N_17361,N_17411);
xor U17459 (N_17459,N_17410,N_17399);
nor U17460 (N_17460,N_17428,N_17372);
nand U17461 (N_17461,N_17332,N_17396);
xnor U17462 (N_17462,N_17313,N_17287);
xnor U17463 (N_17463,N_17352,N_17417);
and U17464 (N_17464,N_17329,N_17388);
or U17465 (N_17465,N_17387,N_17336);
or U17466 (N_17466,N_17281,N_17306);
and U17467 (N_17467,N_17298,N_17362);
and U17468 (N_17468,N_17357,N_17345);
and U17469 (N_17469,N_17338,N_17315);
xor U17470 (N_17470,N_17415,N_17305);
nor U17471 (N_17471,N_17392,N_17333);
and U17472 (N_17472,N_17427,N_17339);
nand U17473 (N_17473,N_17430,N_17355);
and U17474 (N_17474,N_17358,N_17308);
nor U17475 (N_17475,N_17431,N_17419);
and U17476 (N_17476,N_17353,N_17432);
xnor U17477 (N_17477,N_17294,N_17412);
xnor U17478 (N_17478,N_17335,N_17312);
or U17479 (N_17479,N_17348,N_17342);
and U17480 (N_17480,N_17404,N_17380);
xor U17481 (N_17481,N_17370,N_17382);
and U17482 (N_17482,N_17398,N_17386);
or U17483 (N_17483,N_17319,N_17371);
xnor U17484 (N_17484,N_17299,N_17334);
or U17485 (N_17485,N_17283,N_17429);
xnor U17486 (N_17486,N_17301,N_17300);
or U17487 (N_17487,N_17379,N_17356);
nor U17488 (N_17488,N_17303,N_17389);
nor U17489 (N_17489,N_17359,N_17346);
nand U17490 (N_17490,N_17422,N_17317);
nand U17491 (N_17491,N_17290,N_17401);
nor U17492 (N_17492,N_17316,N_17321);
nor U17493 (N_17493,N_17395,N_17434);
and U17494 (N_17494,N_17413,N_17286);
or U17495 (N_17495,N_17284,N_17437);
nor U17496 (N_17496,N_17424,N_17391);
or U17497 (N_17497,N_17377,N_17309);
nand U17498 (N_17498,N_17343,N_17322);
xor U17499 (N_17499,N_17438,N_17324);
or U17500 (N_17500,N_17366,N_17326);
and U17501 (N_17501,N_17423,N_17363);
or U17502 (N_17502,N_17351,N_17304);
nand U17503 (N_17503,N_17416,N_17311);
nand U17504 (N_17504,N_17310,N_17320);
nand U17505 (N_17505,N_17292,N_17390);
xnor U17506 (N_17506,N_17285,N_17325);
xor U17507 (N_17507,N_17327,N_17407);
or U17508 (N_17508,N_17433,N_17385);
or U17509 (N_17509,N_17289,N_17418);
or U17510 (N_17510,N_17293,N_17409);
nand U17511 (N_17511,N_17296,N_17288);
nor U17512 (N_17512,N_17354,N_17414);
xnor U17513 (N_17513,N_17367,N_17400);
nor U17514 (N_17514,N_17302,N_17383);
nand U17515 (N_17515,N_17330,N_17435);
nand U17516 (N_17516,N_17307,N_17341);
nand U17517 (N_17517,N_17318,N_17436);
or U17518 (N_17518,N_17340,N_17403);
or U17519 (N_17519,N_17420,N_17297);
nor U17520 (N_17520,N_17343,N_17348);
and U17521 (N_17521,N_17338,N_17412);
nand U17522 (N_17522,N_17282,N_17390);
or U17523 (N_17523,N_17347,N_17417);
nor U17524 (N_17524,N_17392,N_17281);
and U17525 (N_17525,N_17406,N_17312);
or U17526 (N_17526,N_17284,N_17336);
or U17527 (N_17527,N_17363,N_17433);
or U17528 (N_17528,N_17430,N_17343);
nand U17529 (N_17529,N_17410,N_17359);
xnor U17530 (N_17530,N_17313,N_17290);
nor U17531 (N_17531,N_17362,N_17301);
xor U17532 (N_17532,N_17346,N_17393);
nor U17533 (N_17533,N_17302,N_17397);
nor U17534 (N_17534,N_17428,N_17406);
and U17535 (N_17535,N_17331,N_17320);
nand U17536 (N_17536,N_17285,N_17410);
xor U17537 (N_17537,N_17353,N_17335);
xor U17538 (N_17538,N_17326,N_17381);
nand U17539 (N_17539,N_17395,N_17338);
or U17540 (N_17540,N_17415,N_17378);
nor U17541 (N_17541,N_17381,N_17417);
nor U17542 (N_17542,N_17312,N_17435);
nor U17543 (N_17543,N_17319,N_17323);
nor U17544 (N_17544,N_17305,N_17422);
nor U17545 (N_17545,N_17401,N_17317);
nand U17546 (N_17546,N_17378,N_17345);
and U17547 (N_17547,N_17414,N_17352);
nor U17548 (N_17548,N_17364,N_17400);
xnor U17549 (N_17549,N_17317,N_17375);
xnor U17550 (N_17550,N_17433,N_17384);
nand U17551 (N_17551,N_17421,N_17412);
nand U17552 (N_17552,N_17366,N_17349);
and U17553 (N_17553,N_17430,N_17414);
nor U17554 (N_17554,N_17367,N_17300);
or U17555 (N_17555,N_17300,N_17376);
nor U17556 (N_17556,N_17380,N_17305);
nand U17557 (N_17557,N_17437,N_17302);
xor U17558 (N_17558,N_17369,N_17397);
and U17559 (N_17559,N_17368,N_17416);
xor U17560 (N_17560,N_17314,N_17346);
and U17561 (N_17561,N_17288,N_17350);
nand U17562 (N_17562,N_17420,N_17374);
xnor U17563 (N_17563,N_17399,N_17424);
xor U17564 (N_17564,N_17378,N_17330);
nand U17565 (N_17565,N_17379,N_17339);
nand U17566 (N_17566,N_17422,N_17327);
nor U17567 (N_17567,N_17293,N_17350);
and U17568 (N_17568,N_17394,N_17356);
and U17569 (N_17569,N_17392,N_17311);
nor U17570 (N_17570,N_17291,N_17408);
xor U17571 (N_17571,N_17379,N_17353);
nor U17572 (N_17572,N_17427,N_17371);
and U17573 (N_17573,N_17360,N_17310);
xnor U17574 (N_17574,N_17382,N_17404);
xnor U17575 (N_17575,N_17416,N_17409);
nor U17576 (N_17576,N_17317,N_17289);
and U17577 (N_17577,N_17319,N_17286);
nand U17578 (N_17578,N_17337,N_17342);
xor U17579 (N_17579,N_17295,N_17380);
xnor U17580 (N_17580,N_17407,N_17342);
and U17581 (N_17581,N_17402,N_17328);
nand U17582 (N_17582,N_17397,N_17346);
nor U17583 (N_17583,N_17435,N_17292);
or U17584 (N_17584,N_17383,N_17439);
nand U17585 (N_17585,N_17393,N_17395);
and U17586 (N_17586,N_17433,N_17416);
nor U17587 (N_17587,N_17389,N_17312);
or U17588 (N_17588,N_17364,N_17281);
or U17589 (N_17589,N_17395,N_17318);
nand U17590 (N_17590,N_17349,N_17387);
and U17591 (N_17591,N_17286,N_17395);
or U17592 (N_17592,N_17380,N_17281);
xor U17593 (N_17593,N_17372,N_17346);
nand U17594 (N_17594,N_17281,N_17438);
nand U17595 (N_17595,N_17360,N_17374);
or U17596 (N_17596,N_17439,N_17324);
nand U17597 (N_17597,N_17312,N_17319);
nand U17598 (N_17598,N_17380,N_17438);
nor U17599 (N_17599,N_17283,N_17365);
nand U17600 (N_17600,N_17507,N_17449);
nor U17601 (N_17601,N_17571,N_17566);
and U17602 (N_17602,N_17508,N_17477);
or U17603 (N_17603,N_17521,N_17586);
nor U17604 (N_17604,N_17442,N_17550);
nor U17605 (N_17605,N_17472,N_17538);
and U17606 (N_17606,N_17528,N_17565);
nor U17607 (N_17607,N_17518,N_17587);
nand U17608 (N_17608,N_17564,N_17532);
and U17609 (N_17609,N_17500,N_17557);
nor U17610 (N_17610,N_17547,N_17592);
xnor U17611 (N_17611,N_17458,N_17591);
nor U17612 (N_17612,N_17469,N_17468);
or U17613 (N_17613,N_17456,N_17446);
xor U17614 (N_17614,N_17497,N_17567);
xnor U17615 (N_17615,N_17580,N_17542);
nor U17616 (N_17616,N_17479,N_17510);
nand U17617 (N_17617,N_17447,N_17554);
or U17618 (N_17618,N_17473,N_17594);
nand U17619 (N_17619,N_17579,N_17495);
nor U17620 (N_17620,N_17441,N_17552);
nand U17621 (N_17621,N_17525,N_17482);
or U17622 (N_17622,N_17519,N_17520);
and U17623 (N_17623,N_17526,N_17534);
nand U17624 (N_17624,N_17499,N_17509);
or U17625 (N_17625,N_17524,N_17563);
nand U17626 (N_17626,N_17440,N_17590);
nor U17627 (N_17627,N_17502,N_17560);
or U17628 (N_17628,N_17493,N_17513);
nand U17629 (N_17629,N_17569,N_17486);
and U17630 (N_17630,N_17546,N_17540);
nand U17631 (N_17631,N_17582,N_17577);
xnor U17632 (N_17632,N_17464,N_17533);
xor U17633 (N_17633,N_17475,N_17568);
nand U17634 (N_17634,N_17461,N_17460);
nor U17635 (N_17635,N_17529,N_17593);
nand U17636 (N_17636,N_17512,N_17551);
nand U17637 (N_17637,N_17573,N_17559);
nand U17638 (N_17638,N_17466,N_17536);
nor U17639 (N_17639,N_17583,N_17553);
and U17640 (N_17640,N_17492,N_17596);
xnor U17641 (N_17641,N_17496,N_17505);
xor U17642 (N_17642,N_17467,N_17498);
nand U17643 (N_17643,N_17489,N_17451);
xor U17644 (N_17644,N_17535,N_17531);
nand U17645 (N_17645,N_17450,N_17478);
or U17646 (N_17646,N_17514,N_17516);
xnor U17647 (N_17647,N_17455,N_17462);
and U17648 (N_17648,N_17595,N_17448);
nand U17649 (N_17649,N_17453,N_17454);
nand U17650 (N_17650,N_17556,N_17459);
xnor U17651 (N_17651,N_17543,N_17549);
and U17652 (N_17652,N_17517,N_17480);
nand U17653 (N_17653,N_17465,N_17470);
or U17654 (N_17654,N_17452,N_17488);
nand U17655 (N_17655,N_17537,N_17555);
nand U17656 (N_17656,N_17474,N_17599);
nand U17657 (N_17657,N_17584,N_17494);
nor U17658 (N_17658,N_17445,N_17545);
or U17659 (N_17659,N_17598,N_17522);
and U17660 (N_17660,N_17484,N_17504);
xor U17661 (N_17661,N_17562,N_17515);
and U17662 (N_17662,N_17444,N_17544);
nand U17663 (N_17663,N_17481,N_17539);
nand U17664 (N_17664,N_17443,N_17575);
or U17665 (N_17665,N_17585,N_17561);
and U17666 (N_17666,N_17490,N_17483);
nor U17667 (N_17667,N_17485,N_17597);
xnor U17668 (N_17668,N_17581,N_17476);
nand U17669 (N_17669,N_17572,N_17491);
nand U17670 (N_17670,N_17487,N_17548);
xnor U17671 (N_17671,N_17574,N_17523);
nand U17672 (N_17672,N_17541,N_17530);
nand U17673 (N_17673,N_17506,N_17501);
xor U17674 (N_17674,N_17463,N_17588);
nand U17675 (N_17675,N_17503,N_17589);
and U17676 (N_17676,N_17511,N_17578);
xor U17677 (N_17677,N_17527,N_17558);
and U17678 (N_17678,N_17471,N_17457);
xnor U17679 (N_17679,N_17570,N_17576);
nor U17680 (N_17680,N_17466,N_17530);
nand U17681 (N_17681,N_17505,N_17518);
or U17682 (N_17682,N_17447,N_17445);
or U17683 (N_17683,N_17597,N_17520);
nor U17684 (N_17684,N_17529,N_17581);
xnor U17685 (N_17685,N_17444,N_17560);
nor U17686 (N_17686,N_17592,N_17444);
nor U17687 (N_17687,N_17556,N_17561);
xor U17688 (N_17688,N_17521,N_17585);
or U17689 (N_17689,N_17529,N_17526);
nor U17690 (N_17690,N_17480,N_17497);
xnor U17691 (N_17691,N_17464,N_17450);
and U17692 (N_17692,N_17528,N_17535);
nand U17693 (N_17693,N_17494,N_17452);
xnor U17694 (N_17694,N_17494,N_17491);
or U17695 (N_17695,N_17485,N_17491);
nor U17696 (N_17696,N_17492,N_17535);
nor U17697 (N_17697,N_17568,N_17515);
nor U17698 (N_17698,N_17576,N_17588);
and U17699 (N_17699,N_17468,N_17494);
xnor U17700 (N_17700,N_17443,N_17596);
nor U17701 (N_17701,N_17443,N_17472);
nand U17702 (N_17702,N_17563,N_17568);
and U17703 (N_17703,N_17524,N_17572);
or U17704 (N_17704,N_17509,N_17567);
xnor U17705 (N_17705,N_17566,N_17521);
and U17706 (N_17706,N_17557,N_17473);
nand U17707 (N_17707,N_17587,N_17568);
nand U17708 (N_17708,N_17514,N_17448);
nor U17709 (N_17709,N_17441,N_17529);
nand U17710 (N_17710,N_17489,N_17509);
nand U17711 (N_17711,N_17501,N_17517);
or U17712 (N_17712,N_17462,N_17443);
nand U17713 (N_17713,N_17596,N_17548);
and U17714 (N_17714,N_17597,N_17568);
or U17715 (N_17715,N_17527,N_17523);
nand U17716 (N_17716,N_17520,N_17453);
xnor U17717 (N_17717,N_17454,N_17576);
and U17718 (N_17718,N_17442,N_17475);
or U17719 (N_17719,N_17536,N_17599);
nand U17720 (N_17720,N_17523,N_17520);
xnor U17721 (N_17721,N_17511,N_17443);
xnor U17722 (N_17722,N_17557,N_17560);
or U17723 (N_17723,N_17598,N_17508);
and U17724 (N_17724,N_17599,N_17520);
and U17725 (N_17725,N_17592,N_17452);
or U17726 (N_17726,N_17500,N_17528);
xnor U17727 (N_17727,N_17496,N_17531);
and U17728 (N_17728,N_17517,N_17445);
nor U17729 (N_17729,N_17519,N_17513);
xor U17730 (N_17730,N_17567,N_17452);
nor U17731 (N_17731,N_17591,N_17468);
and U17732 (N_17732,N_17449,N_17553);
xnor U17733 (N_17733,N_17541,N_17585);
xor U17734 (N_17734,N_17467,N_17569);
and U17735 (N_17735,N_17527,N_17536);
xnor U17736 (N_17736,N_17570,N_17494);
nor U17737 (N_17737,N_17553,N_17566);
nor U17738 (N_17738,N_17462,N_17507);
xor U17739 (N_17739,N_17484,N_17571);
nand U17740 (N_17740,N_17590,N_17485);
and U17741 (N_17741,N_17547,N_17501);
or U17742 (N_17742,N_17535,N_17581);
xnor U17743 (N_17743,N_17449,N_17492);
or U17744 (N_17744,N_17583,N_17527);
xnor U17745 (N_17745,N_17471,N_17511);
nor U17746 (N_17746,N_17492,N_17597);
nand U17747 (N_17747,N_17458,N_17507);
xor U17748 (N_17748,N_17528,N_17507);
and U17749 (N_17749,N_17558,N_17470);
nor U17750 (N_17750,N_17567,N_17515);
or U17751 (N_17751,N_17588,N_17584);
nor U17752 (N_17752,N_17552,N_17508);
or U17753 (N_17753,N_17477,N_17479);
nand U17754 (N_17754,N_17464,N_17532);
or U17755 (N_17755,N_17562,N_17595);
or U17756 (N_17756,N_17596,N_17451);
and U17757 (N_17757,N_17452,N_17571);
nor U17758 (N_17758,N_17446,N_17473);
or U17759 (N_17759,N_17576,N_17510);
xor U17760 (N_17760,N_17623,N_17697);
xnor U17761 (N_17761,N_17678,N_17700);
or U17762 (N_17762,N_17707,N_17632);
or U17763 (N_17763,N_17675,N_17759);
nor U17764 (N_17764,N_17742,N_17748);
nor U17765 (N_17765,N_17755,N_17730);
xnor U17766 (N_17766,N_17680,N_17640);
xor U17767 (N_17767,N_17658,N_17741);
xnor U17768 (N_17768,N_17715,N_17643);
nand U17769 (N_17769,N_17743,N_17684);
or U17770 (N_17770,N_17674,N_17687);
xnor U17771 (N_17771,N_17711,N_17745);
nor U17772 (N_17772,N_17717,N_17616);
xor U17773 (N_17773,N_17624,N_17628);
and U17774 (N_17774,N_17671,N_17676);
xnor U17775 (N_17775,N_17663,N_17627);
xor U17776 (N_17776,N_17653,N_17729);
nor U17777 (N_17777,N_17716,N_17656);
nand U17778 (N_17778,N_17622,N_17669);
nand U17779 (N_17779,N_17751,N_17696);
or U17780 (N_17780,N_17689,N_17756);
nor U17781 (N_17781,N_17629,N_17737);
or U17782 (N_17782,N_17692,N_17733);
and U17783 (N_17783,N_17703,N_17665);
or U17784 (N_17784,N_17735,N_17668);
nand U17785 (N_17785,N_17723,N_17608);
or U17786 (N_17786,N_17673,N_17638);
or U17787 (N_17787,N_17602,N_17708);
or U17788 (N_17788,N_17609,N_17618);
or U17789 (N_17789,N_17718,N_17636);
or U17790 (N_17790,N_17637,N_17648);
xnor U17791 (N_17791,N_17709,N_17650);
nand U17792 (N_17792,N_17605,N_17641);
nor U17793 (N_17793,N_17639,N_17734);
nor U17794 (N_17794,N_17630,N_17651);
xnor U17795 (N_17795,N_17647,N_17615);
nor U17796 (N_17796,N_17726,N_17683);
nor U17797 (N_17797,N_17661,N_17625);
nor U17798 (N_17798,N_17659,N_17613);
xnor U17799 (N_17799,N_17631,N_17739);
or U17800 (N_17800,N_17621,N_17603);
xnor U17801 (N_17801,N_17740,N_17691);
or U17802 (N_17802,N_17649,N_17682);
nand U17803 (N_17803,N_17705,N_17744);
nand U17804 (N_17804,N_17706,N_17654);
xnor U17805 (N_17805,N_17695,N_17617);
nand U17806 (N_17806,N_17644,N_17614);
nand U17807 (N_17807,N_17719,N_17610);
nor U17808 (N_17808,N_17746,N_17657);
or U17809 (N_17809,N_17664,N_17601);
nor U17810 (N_17810,N_17660,N_17600);
or U17811 (N_17811,N_17724,N_17611);
xor U17812 (N_17812,N_17633,N_17732);
or U17813 (N_17813,N_17606,N_17714);
nand U17814 (N_17814,N_17677,N_17704);
nand U17815 (N_17815,N_17727,N_17731);
or U17816 (N_17816,N_17750,N_17701);
or U17817 (N_17817,N_17679,N_17694);
and U17818 (N_17818,N_17642,N_17712);
or U17819 (N_17819,N_17713,N_17688);
xor U17820 (N_17820,N_17753,N_17725);
and U17821 (N_17821,N_17754,N_17710);
or U17822 (N_17822,N_17619,N_17607);
nand U17823 (N_17823,N_17604,N_17752);
nor U17824 (N_17824,N_17626,N_17690);
nor U17825 (N_17825,N_17655,N_17634);
xnor U17826 (N_17826,N_17620,N_17749);
nand U17827 (N_17827,N_17736,N_17662);
nand U17828 (N_17828,N_17685,N_17670);
or U17829 (N_17829,N_17699,N_17747);
or U17830 (N_17830,N_17721,N_17635);
nor U17831 (N_17831,N_17722,N_17612);
xnor U17832 (N_17832,N_17667,N_17738);
nand U17833 (N_17833,N_17681,N_17645);
and U17834 (N_17834,N_17698,N_17686);
xor U17835 (N_17835,N_17672,N_17702);
and U17836 (N_17836,N_17666,N_17693);
or U17837 (N_17837,N_17646,N_17728);
and U17838 (N_17838,N_17758,N_17720);
nand U17839 (N_17839,N_17757,N_17652);
or U17840 (N_17840,N_17605,N_17625);
and U17841 (N_17841,N_17614,N_17651);
xor U17842 (N_17842,N_17626,N_17749);
or U17843 (N_17843,N_17627,N_17727);
nor U17844 (N_17844,N_17613,N_17750);
or U17845 (N_17845,N_17672,N_17681);
nor U17846 (N_17846,N_17738,N_17677);
nand U17847 (N_17847,N_17690,N_17610);
nand U17848 (N_17848,N_17641,N_17601);
nor U17849 (N_17849,N_17700,N_17684);
or U17850 (N_17850,N_17696,N_17732);
nor U17851 (N_17851,N_17618,N_17712);
nor U17852 (N_17852,N_17613,N_17686);
nand U17853 (N_17853,N_17636,N_17620);
nor U17854 (N_17854,N_17627,N_17745);
and U17855 (N_17855,N_17750,N_17699);
and U17856 (N_17856,N_17743,N_17609);
nor U17857 (N_17857,N_17646,N_17672);
nor U17858 (N_17858,N_17613,N_17736);
or U17859 (N_17859,N_17722,N_17645);
xnor U17860 (N_17860,N_17637,N_17703);
nor U17861 (N_17861,N_17702,N_17697);
nand U17862 (N_17862,N_17744,N_17694);
xnor U17863 (N_17863,N_17645,N_17724);
nand U17864 (N_17864,N_17611,N_17655);
nand U17865 (N_17865,N_17711,N_17627);
xnor U17866 (N_17866,N_17661,N_17683);
xnor U17867 (N_17867,N_17626,N_17732);
nor U17868 (N_17868,N_17663,N_17666);
or U17869 (N_17869,N_17636,N_17710);
xnor U17870 (N_17870,N_17634,N_17605);
nand U17871 (N_17871,N_17628,N_17756);
xor U17872 (N_17872,N_17612,N_17737);
nor U17873 (N_17873,N_17715,N_17709);
nand U17874 (N_17874,N_17725,N_17744);
or U17875 (N_17875,N_17733,N_17699);
and U17876 (N_17876,N_17728,N_17752);
and U17877 (N_17877,N_17675,N_17742);
xor U17878 (N_17878,N_17694,N_17668);
xnor U17879 (N_17879,N_17650,N_17641);
xor U17880 (N_17880,N_17662,N_17605);
nor U17881 (N_17881,N_17701,N_17622);
nor U17882 (N_17882,N_17693,N_17619);
and U17883 (N_17883,N_17703,N_17643);
or U17884 (N_17884,N_17662,N_17699);
nand U17885 (N_17885,N_17690,N_17651);
nand U17886 (N_17886,N_17717,N_17638);
xor U17887 (N_17887,N_17614,N_17673);
xnor U17888 (N_17888,N_17603,N_17729);
or U17889 (N_17889,N_17687,N_17670);
nor U17890 (N_17890,N_17727,N_17699);
nor U17891 (N_17891,N_17744,N_17685);
xnor U17892 (N_17892,N_17652,N_17704);
and U17893 (N_17893,N_17744,N_17717);
or U17894 (N_17894,N_17681,N_17743);
and U17895 (N_17895,N_17724,N_17756);
nand U17896 (N_17896,N_17679,N_17687);
xnor U17897 (N_17897,N_17617,N_17612);
and U17898 (N_17898,N_17607,N_17665);
xor U17899 (N_17899,N_17754,N_17617);
and U17900 (N_17900,N_17700,N_17606);
nor U17901 (N_17901,N_17659,N_17675);
xnor U17902 (N_17902,N_17680,N_17711);
nand U17903 (N_17903,N_17680,N_17722);
nor U17904 (N_17904,N_17652,N_17656);
nor U17905 (N_17905,N_17728,N_17759);
or U17906 (N_17906,N_17755,N_17687);
nor U17907 (N_17907,N_17622,N_17608);
xnor U17908 (N_17908,N_17674,N_17694);
nor U17909 (N_17909,N_17745,N_17646);
nor U17910 (N_17910,N_17613,N_17643);
or U17911 (N_17911,N_17612,N_17707);
nand U17912 (N_17912,N_17755,N_17664);
nand U17913 (N_17913,N_17684,N_17676);
xnor U17914 (N_17914,N_17637,N_17616);
or U17915 (N_17915,N_17620,N_17719);
or U17916 (N_17916,N_17684,N_17688);
xor U17917 (N_17917,N_17686,N_17600);
or U17918 (N_17918,N_17695,N_17747);
or U17919 (N_17919,N_17680,N_17740);
or U17920 (N_17920,N_17878,N_17820);
nand U17921 (N_17921,N_17803,N_17845);
nand U17922 (N_17922,N_17791,N_17855);
and U17923 (N_17923,N_17870,N_17764);
nor U17924 (N_17924,N_17874,N_17818);
or U17925 (N_17925,N_17768,N_17843);
nor U17926 (N_17926,N_17807,N_17915);
nand U17927 (N_17927,N_17821,N_17904);
nor U17928 (N_17928,N_17873,N_17798);
or U17929 (N_17929,N_17912,N_17861);
and U17930 (N_17930,N_17899,N_17856);
nand U17931 (N_17931,N_17771,N_17852);
and U17932 (N_17932,N_17853,N_17892);
or U17933 (N_17933,N_17827,N_17787);
xnor U17934 (N_17934,N_17869,N_17863);
and U17935 (N_17935,N_17829,N_17761);
and U17936 (N_17936,N_17871,N_17882);
and U17937 (N_17937,N_17822,N_17781);
nand U17938 (N_17938,N_17819,N_17824);
nor U17939 (N_17939,N_17888,N_17877);
or U17940 (N_17940,N_17913,N_17770);
nor U17941 (N_17941,N_17766,N_17801);
and U17942 (N_17942,N_17907,N_17910);
and U17943 (N_17943,N_17898,N_17808);
nand U17944 (N_17944,N_17812,N_17867);
nor U17945 (N_17945,N_17901,N_17826);
nor U17946 (N_17946,N_17794,N_17846);
nor U17947 (N_17947,N_17914,N_17885);
or U17948 (N_17948,N_17793,N_17847);
nand U17949 (N_17949,N_17780,N_17891);
nor U17950 (N_17950,N_17893,N_17817);
and U17951 (N_17951,N_17851,N_17919);
xnor U17952 (N_17952,N_17916,N_17876);
nand U17953 (N_17953,N_17868,N_17850);
xor U17954 (N_17954,N_17864,N_17903);
xor U17955 (N_17955,N_17783,N_17835);
nor U17956 (N_17956,N_17767,N_17894);
or U17957 (N_17957,N_17834,N_17862);
xnor U17958 (N_17958,N_17779,N_17790);
nor U17959 (N_17959,N_17830,N_17879);
and U17960 (N_17960,N_17800,N_17763);
nand U17961 (N_17961,N_17796,N_17859);
and U17962 (N_17962,N_17906,N_17762);
nand U17963 (N_17963,N_17823,N_17809);
xnor U17964 (N_17964,N_17909,N_17782);
xnor U17965 (N_17965,N_17875,N_17806);
or U17966 (N_17966,N_17848,N_17816);
or U17967 (N_17967,N_17775,N_17917);
or U17968 (N_17968,N_17777,N_17857);
nor U17969 (N_17969,N_17837,N_17849);
and U17970 (N_17970,N_17802,N_17805);
nand U17971 (N_17971,N_17908,N_17840);
or U17972 (N_17972,N_17905,N_17902);
nand U17973 (N_17973,N_17833,N_17831);
xnor U17974 (N_17974,N_17784,N_17866);
nand U17975 (N_17975,N_17832,N_17839);
xnor U17976 (N_17976,N_17883,N_17785);
xor U17977 (N_17977,N_17838,N_17911);
nand U17978 (N_17978,N_17900,N_17890);
or U17979 (N_17979,N_17765,N_17760);
xor U17980 (N_17980,N_17789,N_17773);
nor U17981 (N_17981,N_17844,N_17842);
xor U17982 (N_17982,N_17792,N_17797);
xnor U17983 (N_17983,N_17776,N_17825);
and U17984 (N_17984,N_17774,N_17815);
or U17985 (N_17985,N_17880,N_17865);
or U17986 (N_17986,N_17786,N_17884);
nand U17987 (N_17987,N_17881,N_17887);
xor U17988 (N_17988,N_17788,N_17854);
or U17989 (N_17989,N_17814,N_17828);
nor U17990 (N_17990,N_17872,N_17804);
nand U17991 (N_17991,N_17897,N_17810);
and U17992 (N_17992,N_17841,N_17858);
and U17993 (N_17993,N_17895,N_17896);
nor U17994 (N_17994,N_17795,N_17918);
and U17995 (N_17995,N_17769,N_17778);
xor U17996 (N_17996,N_17886,N_17813);
and U17997 (N_17997,N_17836,N_17889);
and U17998 (N_17998,N_17860,N_17799);
and U17999 (N_17999,N_17811,N_17772);
nor U18000 (N_18000,N_17781,N_17808);
or U18001 (N_18001,N_17839,N_17876);
nor U18002 (N_18002,N_17771,N_17804);
xnor U18003 (N_18003,N_17898,N_17880);
or U18004 (N_18004,N_17809,N_17804);
nor U18005 (N_18005,N_17776,N_17804);
nand U18006 (N_18006,N_17882,N_17844);
nor U18007 (N_18007,N_17785,N_17766);
or U18008 (N_18008,N_17893,N_17884);
and U18009 (N_18009,N_17789,N_17782);
xor U18010 (N_18010,N_17900,N_17785);
nand U18011 (N_18011,N_17785,N_17802);
xor U18012 (N_18012,N_17787,N_17822);
or U18013 (N_18013,N_17902,N_17818);
nand U18014 (N_18014,N_17777,N_17795);
or U18015 (N_18015,N_17870,N_17823);
nor U18016 (N_18016,N_17870,N_17832);
or U18017 (N_18017,N_17854,N_17829);
nor U18018 (N_18018,N_17848,N_17782);
and U18019 (N_18019,N_17766,N_17877);
nor U18020 (N_18020,N_17838,N_17885);
and U18021 (N_18021,N_17829,N_17862);
and U18022 (N_18022,N_17784,N_17845);
xor U18023 (N_18023,N_17848,N_17811);
and U18024 (N_18024,N_17788,N_17873);
xnor U18025 (N_18025,N_17772,N_17843);
or U18026 (N_18026,N_17848,N_17807);
nand U18027 (N_18027,N_17815,N_17780);
xnor U18028 (N_18028,N_17901,N_17805);
and U18029 (N_18029,N_17845,N_17819);
or U18030 (N_18030,N_17831,N_17904);
nor U18031 (N_18031,N_17859,N_17856);
xnor U18032 (N_18032,N_17869,N_17771);
and U18033 (N_18033,N_17801,N_17871);
nand U18034 (N_18034,N_17802,N_17845);
xor U18035 (N_18035,N_17879,N_17890);
nor U18036 (N_18036,N_17805,N_17835);
nor U18037 (N_18037,N_17830,N_17776);
nor U18038 (N_18038,N_17808,N_17913);
or U18039 (N_18039,N_17834,N_17826);
and U18040 (N_18040,N_17911,N_17762);
or U18041 (N_18041,N_17797,N_17774);
or U18042 (N_18042,N_17897,N_17918);
nor U18043 (N_18043,N_17786,N_17904);
nand U18044 (N_18044,N_17796,N_17840);
xor U18045 (N_18045,N_17779,N_17886);
and U18046 (N_18046,N_17887,N_17914);
nand U18047 (N_18047,N_17763,N_17894);
and U18048 (N_18048,N_17838,N_17842);
or U18049 (N_18049,N_17886,N_17843);
xor U18050 (N_18050,N_17763,N_17772);
nand U18051 (N_18051,N_17898,N_17907);
xnor U18052 (N_18052,N_17765,N_17892);
nand U18053 (N_18053,N_17843,N_17916);
nand U18054 (N_18054,N_17860,N_17859);
xnor U18055 (N_18055,N_17871,N_17770);
nand U18056 (N_18056,N_17906,N_17865);
nand U18057 (N_18057,N_17856,N_17763);
nand U18058 (N_18058,N_17789,N_17835);
nand U18059 (N_18059,N_17766,N_17822);
and U18060 (N_18060,N_17892,N_17824);
nand U18061 (N_18061,N_17903,N_17792);
nand U18062 (N_18062,N_17827,N_17860);
and U18063 (N_18063,N_17912,N_17770);
nor U18064 (N_18064,N_17798,N_17885);
nor U18065 (N_18065,N_17784,N_17840);
xnor U18066 (N_18066,N_17892,N_17867);
and U18067 (N_18067,N_17808,N_17844);
xor U18068 (N_18068,N_17809,N_17884);
and U18069 (N_18069,N_17800,N_17876);
nand U18070 (N_18070,N_17810,N_17773);
and U18071 (N_18071,N_17832,N_17818);
or U18072 (N_18072,N_17830,N_17911);
or U18073 (N_18073,N_17795,N_17811);
or U18074 (N_18074,N_17852,N_17891);
or U18075 (N_18075,N_17797,N_17885);
nor U18076 (N_18076,N_17766,N_17910);
and U18077 (N_18077,N_17887,N_17858);
and U18078 (N_18078,N_17796,N_17788);
nor U18079 (N_18079,N_17837,N_17782);
nor U18080 (N_18080,N_18030,N_18079);
nor U18081 (N_18081,N_17935,N_17939);
nor U18082 (N_18082,N_17987,N_17920);
or U18083 (N_18083,N_17997,N_17990);
and U18084 (N_18084,N_18020,N_18006);
or U18085 (N_18085,N_17937,N_18011);
or U18086 (N_18086,N_17960,N_17929);
or U18087 (N_18087,N_17977,N_17928);
or U18088 (N_18088,N_18071,N_18037);
or U18089 (N_18089,N_18038,N_17976);
or U18090 (N_18090,N_17953,N_17978);
or U18091 (N_18091,N_18035,N_17991);
nand U18092 (N_18092,N_17951,N_17947);
and U18093 (N_18093,N_18048,N_18056);
nor U18094 (N_18094,N_17925,N_18027);
nor U18095 (N_18095,N_17934,N_18062);
xor U18096 (N_18096,N_17957,N_17962);
and U18097 (N_18097,N_18078,N_18044);
nor U18098 (N_18098,N_18065,N_17942);
or U18099 (N_18099,N_17946,N_17943);
and U18100 (N_18100,N_18018,N_18054);
or U18101 (N_18101,N_17989,N_17998);
or U18102 (N_18102,N_17958,N_18049);
or U18103 (N_18103,N_18001,N_18047);
nor U18104 (N_18104,N_18064,N_18069);
and U18105 (N_18105,N_18009,N_17992);
xor U18106 (N_18106,N_17954,N_18063);
and U18107 (N_18107,N_17959,N_18015);
nor U18108 (N_18108,N_17921,N_17982);
nand U18109 (N_18109,N_17974,N_18002);
nor U18110 (N_18110,N_17988,N_18026);
xor U18111 (N_18111,N_18042,N_17994);
nor U18112 (N_18112,N_18036,N_18032);
nand U18113 (N_18113,N_17964,N_17986);
nand U18114 (N_18114,N_18031,N_18068);
or U18115 (N_18115,N_18010,N_17993);
and U18116 (N_18116,N_17969,N_18014);
and U18117 (N_18117,N_17981,N_17965);
and U18118 (N_18118,N_18057,N_18041);
and U18119 (N_18119,N_18004,N_18033);
or U18120 (N_18120,N_18007,N_17999);
and U18121 (N_18121,N_17948,N_18008);
and U18122 (N_18122,N_17995,N_18058);
xor U18123 (N_18123,N_17955,N_17966);
or U18124 (N_18124,N_17963,N_18055);
nand U18125 (N_18125,N_17950,N_17936);
or U18126 (N_18126,N_17973,N_17952);
or U18127 (N_18127,N_18073,N_17975);
and U18128 (N_18128,N_17968,N_17985);
or U18129 (N_18129,N_17979,N_17944);
nor U18130 (N_18130,N_17961,N_18019);
nand U18131 (N_18131,N_18046,N_18012);
and U18132 (N_18132,N_18005,N_17924);
nand U18133 (N_18133,N_18003,N_18039);
and U18134 (N_18134,N_18021,N_17996);
and U18135 (N_18135,N_18077,N_17941);
xor U18136 (N_18136,N_18067,N_18060);
and U18137 (N_18137,N_18022,N_17956);
nand U18138 (N_18138,N_17983,N_18070);
nand U18139 (N_18139,N_18072,N_18045);
xnor U18140 (N_18140,N_17949,N_18040);
nor U18141 (N_18141,N_17945,N_18023);
xor U18142 (N_18142,N_18052,N_17970);
xor U18143 (N_18143,N_18025,N_17930);
xor U18144 (N_18144,N_17971,N_17932);
nand U18145 (N_18145,N_18061,N_17984);
nand U18146 (N_18146,N_17923,N_18016);
and U18147 (N_18147,N_18043,N_17931);
nor U18148 (N_18148,N_18000,N_18024);
or U18149 (N_18149,N_18017,N_17967);
nand U18150 (N_18150,N_18029,N_18050);
nand U18151 (N_18151,N_18076,N_17922);
nand U18152 (N_18152,N_18028,N_17927);
nor U18153 (N_18153,N_17933,N_18034);
and U18154 (N_18154,N_17980,N_18075);
nor U18155 (N_18155,N_18053,N_18074);
xor U18156 (N_18156,N_17938,N_18059);
and U18157 (N_18157,N_18051,N_18013);
nor U18158 (N_18158,N_17972,N_17940);
and U18159 (N_18159,N_17926,N_18066);
nor U18160 (N_18160,N_17993,N_18028);
nand U18161 (N_18161,N_17988,N_17970);
or U18162 (N_18162,N_17929,N_17996);
nand U18163 (N_18163,N_18030,N_17976);
nor U18164 (N_18164,N_17932,N_17934);
nand U18165 (N_18165,N_18072,N_17992);
xnor U18166 (N_18166,N_17996,N_18035);
xnor U18167 (N_18167,N_18054,N_17988);
and U18168 (N_18168,N_18071,N_17975);
and U18169 (N_18169,N_17993,N_17954);
and U18170 (N_18170,N_17981,N_18075);
nand U18171 (N_18171,N_17940,N_18060);
xor U18172 (N_18172,N_18000,N_18064);
nor U18173 (N_18173,N_18074,N_17926);
or U18174 (N_18174,N_18011,N_17922);
or U18175 (N_18175,N_17933,N_18036);
nand U18176 (N_18176,N_17977,N_17930);
xor U18177 (N_18177,N_18008,N_18015);
nand U18178 (N_18178,N_17994,N_18025);
and U18179 (N_18179,N_18019,N_18023);
and U18180 (N_18180,N_17937,N_17953);
and U18181 (N_18181,N_17975,N_17931);
nor U18182 (N_18182,N_18078,N_18023);
nand U18183 (N_18183,N_17975,N_17976);
nand U18184 (N_18184,N_17988,N_17942);
or U18185 (N_18185,N_17931,N_18013);
nor U18186 (N_18186,N_18058,N_17984);
or U18187 (N_18187,N_17980,N_18054);
or U18188 (N_18188,N_17958,N_17974);
nor U18189 (N_18189,N_17951,N_17922);
or U18190 (N_18190,N_18027,N_18002);
or U18191 (N_18191,N_18050,N_18011);
xor U18192 (N_18192,N_18078,N_18076);
nand U18193 (N_18193,N_17940,N_17958);
and U18194 (N_18194,N_17932,N_18000);
nor U18195 (N_18195,N_18063,N_17957);
xnor U18196 (N_18196,N_18065,N_17977);
nand U18197 (N_18197,N_17964,N_17930);
or U18198 (N_18198,N_18057,N_17986);
and U18199 (N_18199,N_17967,N_17926);
xor U18200 (N_18200,N_17981,N_18039);
nor U18201 (N_18201,N_18018,N_17983);
nand U18202 (N_18202,N_17973,N_17989);
and U18203 (N_18203,N_17956,N_18045);
xnor U18204 (N_18204,N_18073,N_18012);
or U18205 (N_18205,N_18071,N_18040);
nor U18206 (N_18206,N_17993,N_18016);
nand U18207 (N_18207,N_17958,N_18004);
xor U18208 (N_18208,N_18079,N_17926);
nor U18209 (N_18209,N_17966,N_18064);
or U18210 (N_18210,N_17987,N_17960);
and U18211 (N_18211,N_18039,N_18025);
xnor U18212 (N_18212,N_18014,N_17929);
or U18213 (N_18213,N_18015,N_17936);
and U18214 (N_18214,N_17970,N_17952);
nand U18215 (N_18215,N_18053,N_17972);
nor U18216 (N_18216,N_17970,N_17950);
xnor U18217 (N_18217,N_17991,N_17986);
and U18218 (N_18218,N_17971,N_17924);
and U18219 (N_18219,N_17987,N_18030);
nand U18220 (N_18220,N_18003,N_17994);
and U18221 (N_18221,N_17961,N_17959);
and U18222 (N_18222,N_17944,N_17976);
nand U18223 (N_18223,N_18068,N_18015);
and U18224 (N_18224,N_17974,N_18038);
and U18225 (N_18225,N_18033,N_17965);
nand U18226 (N_18226,N_18043,N_18049);
nand U18227 (N_18227,N_17945,N_18038);
or U18228 (N_18228,N_18053,N_18032);
and U18229 (N_18229,N_17967,N_18067);
nor U18230 (N_18230,N_18022,N_17997);
nand U18231 (N_18231,N_18001,N_18029);
or U18232 (N_18232,N_17946,N_17947);
nor U18233 (N_18233,N_17998,N_17965);
nand U18234 (N_18234,N_18046,N_17971);
xor U18235 (N_18235,N_18034,N_18021);
xnor U18236 (N_18236,N_17968,N_18031);
nand U18237 (N_18237,N_18064,N_18007);
and U18238 (N_18238,N_17999,N_17936);
or U18239 (N_18239,N_17993,N_18001);
xor U18240 (N_18240,N_18177,N_18195);
xnor U18241 (N_18241,N_18209,N_18113);
and U18242 (N_18242,N_18109,N_18198);
and U18243 (N_18243,N_18120,N_18167);
xor U18244 (N_18244,N_18197,N_18080);
or U18245 (N_18245,N_18122,N_18175);
nand U18246 (N_18246,N_18235,N_18233);
and U18247 (N_18247,N_18130,N_18126);
nand U18248 (N_18248,N_18119,N_18155);
or U18249 (N_18249,N_18215,N_18117);
xor U18250 (N_18250,N_18129,N_18230);
or U18251 (N_18251,N_18218,N_18161);
and U18252 (N_18252,N_18153,N_18173);
and U18253 (N_18253,N_18157,N_18221);
xnor U18254 (N_18254,N_18094,N_18170);
xnor U18255 (N_18255,N_18100,N_18135);
and U18256 (N_18256,N_18144,N_18115);
nand U18257 (N_18257,N_18099,N_18185);
xor U18258 (N_18258,N_18238,N_18140);
nand U18259 (N_18259,N_18166,N_18211);
or U18260 (N_18260,N_18159,N_18183);
xnor U18261 (N_18261,N_18156,N_18200);
and U18262 (N_18262,N_18133,N_18207);
nor U18263 (N_18263,N_18106,N_18160);
nand U18264 (N_18264,N_18108,N_18188);
and U18265 (N_18265,N_18237,N_18182);
or U18266 (N_18266,N_18220,N_18138);
xor U18267 (N_18267,N_18102,N_18189);
or U18268 (N_18268,N_18151,N_18158);
and U18269 (N_18269,N_18227,N_18229);
nand U18270 (N_18270,N_18148,N_18191);
xor U18271 (N_18271,N_18104,N_18093);
nor U18272 (N_18272,N_18083,N_18194);
nor U18273 (N_18273,N_18168,N_18095);
or U18274 (N_18274,N_18199,N_18234);
nand U18275 (N_18275,N_18097,N_18201);
or U18276 (N_18276,N_18223,N_18134);
nor U18277 (N_18277,N_18136,N_18084);
nand U18278 (N_18278,N_18181,N_18121);
or U18279 (N_18279,N_18162,N_18184);
or U18280 (N_18280,N_18226,N_18087);
xnor U18281 (N_18281,N_18096,N_18210);
nand U18282 (N_18282,N_18163,N_18179);
xor U18283 (N_18283,N_18149,N_18204);
xnor U18284 (N_18284,N_18088,N_18196);
nand U18285 (N_18285,N_18111,N_18239);
nor U18286 (N_18286,N_18110,N_18090);
xor U18287 (N_18287,N_18082,N_18085);
xnor U18288 (N_18288,N_18164,N_18139);
nor U18289 (N_18289,N_18118,N_18174);
xnor U18290 (N_18290,N_18101,N_18142);
and U18291 (N_18291,N_18086,N_18137);
and U18292 (N_18292,N_18219,N_18127);
or U18293 (N_18293,N_18092,N_18205);
xnor U18294 (N_18294,N_18228,N_18212);
nor U18295 (N_18295,N_18180,N_18232);
and U18296 (N_18296,N_18213,N_18150);
xnor U18297 (N_18297,N_18143,N_18116);
or U18298 (N_18298,N_18128,N_18091);
nor U18299 (N_18299,N_18187,N_18114);
or U18300 (N_18300,N_18217,N_18169);
or U18301 (N_18301,N_18172,N_18231);
or U18302 (N_18302,N_18123,N_18112);
nor U18303 (N_18303,N_18202,N_18222);
xor U18304 (N_18304,N_18146,N_18098);
or U18305 (N_18305,N_18089,N_18208);
and U18306 (N_18306,N_18176,N_18192);
nor U18307 (N_18307,N_18190,N_18165);
xnor U18308 (N_18308,N_18236,N_18103);
or U18309 (N_18309,N_18081,N_18224);
or U18310 (N_18310,N_18145,N_18132);
nor U18311 (N_18311,N_18225,N_18186);
nand U18312 (N_18312,N_18125,N_18107);
nand U18313 (N_18313,N_18216,N_18124);
nor U18314 (N_18314,N_18193,N_18203);
xnor U18315 (N_18315,N_18105,N_18178);
nand U18316 (N_18316,N_18131,N_18152);
xor U18317 (N_18317,N_18214,N_18171);
and U18318 (N_18318,N_18147,N_18141);
or U18319 (N_18319,N_18206,N_18154);
nand U18320 (N_18320,N_18222,N_18165);
xnor U18321 (N_18321,N_18237,N_18098);
nand U18322 (N_18322,N_18101,N_18237);
xnor U18323 (N_18323,N_18173,N_18148);
xor U18324 (N_18324,N_18170,N_18201);
nand U18325 (N_18325,N_18139,N_18178);
or U18326 (N_18326,N_18184,N_18190);
or U18327 (N_18327,N_18159,N_18157);
nor U18328 (N_18328,N_18115,N_18105);
and U18329 (N_18329,N_18220,N_18218);
or U18330 (N_18330,N_18121,N_18140);
xnor U18331 (N_18331,N_18089,N_18239);
xnor U18332 (N_18332,N_18164,N_18158);
or U18333 (N_18333,N_18220,N_18202);
xor U18334 (N_18334,N_18212,N_18213);
and U18335 (N_18335,N_18184,N_18088);
nand U18336 (N_18336,N_18201,N_18114);
and U18337 (N_18337,N_18213,N_18226);
and U18338 (N_18338,N_18224,N_18152);
and U18339 (N_18339,N_18080,N_18090);
nand U18340 (N_18340,N_18089,N_18087);
nor U18341 (N_18341,N_18235,N_18161);
or U18342 (N_18342,N_18086,N_18218);
nor U18343 (N_18343,N_18169,N_18183);
xor U18344 (N_18344,N_18236,N_18208);
nand U18345 (N_18345,N_18227,N_18230);
or U18346 (N_18346,N_18212,N_18129);
nor U18347 (N_18347,N_18095,N_18226);
and U18348 (N_18348,N_18147,N_18184);
nand U18349 (N_18349,N_18221,N_18084);
xnor U18350 (N_18350,N_18131,N_18217);
and U18351 (N_18351,N_18088,N_18188);
nor U18352 (N_18352,N_18208,N_18202);
and U18353 (N_18353,N_18099,N_18142);
nor U18354 (N_18354,N_18147,N_18107);
xnor U18355 (N_18355,N_18083,N_18239);
xnor U18356 (N_18356,N_18154,N_18099);
or U18357 (N_18357,N_18176,N_18111);
and U18358 (N_18358,N_18137,N_18199);
nor U18359 (N_18359,N_18199,N_18151);
or U18360 (N_18360,N_18123,N_18202);
nor U18361 (N_18361,N_18093,N_18098);
or U18362 (N_18362,N_18189,N_18085);
or U18363 (N_18363,N_18232,N_18112);
xor U18364 (N_18364,N_18200,N_18098);
and U18365 (N_18365,N_18168,N_18194);
xnor U18366 (N_18366,N_18081,N_18118);
nand U18367 (N_18367,N_18116,N_18236);
nand U18368 (N_18368,N_18205,N_18139);
and U18369 (N_18369,N_18160,N_18147);
nor U18370 (N_18370,N_18082,N_18144);
or U18371 (N_18371,N_18117,N_18192);
or U18372 (N_18372,N_18207,N_18092);
or U18373 (N_18373,N_18103,N_18162);
and U18374 (N_18374,N_18188,N_18191);
nor U18375 (N_18375,N_18206,N_18151);
and U18376 (N_18376,N_18160,N_18118);
xnor U18377 (N_18377,N_18115,N_18141);
xor U18378 (N_18378,N_18211,N_18213);
nor U18379 (N_18379,N_18230,N_18164);
or U18380 (N_18380,N_18085,N_18162);
and U18381 (N_18381,N_18117,N_18119);
nand U18382 (N_18382,N_18097,N_18197);
nand U18383 (N_18383,N_18099,N_18137);
nand U18384 (N_18384,N_18237,N_18208);
xnor U18385 (N_18385,N_18167,N_18119);
nor U18386 (N_18386,N_18121,N_18088);
nand U18387 (N_18387,N_18171,N_18224);
and U18388 (N_18388,N_18211,N_18145);
or U18389 (N_18389,N_18231,N_18180);
or U18390 (N_18390,N_18097,N_18110);
xor U18391 (N_18391,N_18171,N_18092);
or U18392 (N_18392,N_18218,N_18199);
and U18393 (N_18393,N_18188,N_18175);
nand U18394 (N_18394,N_18214,N_18156);
or U18395 (N_18395,N_18198,N_18130);
and U18396 (N_18396,N_18211,N_18216);
and U18397 (N_18397,N_18154,N_18109);
xor U18398 (N_18398,N_18228,N_18189);
nand U18399 (N_18399,N_18127,N_18159);
nor U18400 (N_18400,N_18345,N_18244);
nand U18401 (N_18401,N_18250,N_18278);
and U18402 (N_18402,N_18290,N_18320);
xor U18403 (N_18403,N_18266,N_18394);
and U18404 (N_18404,N_18315,N_18264);
nand U18405 (N_18405,N_18327,N_18254);
nor U18406 (N_18406,N_18241,N_18387);
nor U18407 (N_18407,N_18322,N_18393);
and U18408 (N_18408,N_18294,N_18304);
xor U18409 (N_18409,N_18319,N_18312);
and U18410 (N_18410,N_18340,N_18374);
nor U18411 (N_18411,N_18251,N_18314);
and U18412 (N_18412,N_18279,N_18333);
nand U18413 (N_18413,N_18260,N_18318);
nand U18414 (N_18414,N_18396,N_18391);
or U18415 (N_18415,N_18325,N_18270);
nand U18416 (N_18416,N_18317,N_18363);
or U18417 (N_18417,N_18328,N_18259);
and U18418 (N_18418,N_18330,N_18375);
xnor U18419 (N_18419,N_18397,N_18267);
xnor U18420 (N_18420,N_18338,N_18305);
nand U18421 (N_18421,N_18337,N_18326);
and U18422 (N_18422,N_18356,N_18347);
nand U18423 (N_18423,N_18274,N_18306);
xnor U18424 (N_18424,N_18395,N_18298);
nand U18425 (N_18425,N_18369,N_18355);
nand U18426 (N_18426,N_18303,N_18370);
and U18427 (N_18427,N_18358,N_18308);
nand U18428 (N_18428,N_18362,N_18247);
or U18429 (N_18429,N_18342,N_18242);
nand U18430 (N_18430,N_18353,N_18292);
nor U18431 (N_18431,N_18385,N_18386);
nand U18432 (N_18432,N_18299,N_18357);
nand U18433 (N_18433,N_18390,N_18344);
nand U18434 (N_18434,N_18336,N_18268);
and U18435 (N_18435,N_18379,N_18271);
or U18436 (N_18436,N_18243,N_18332);
nand U18437 (N_18437,N_18366,N_18360);
nand U18438 (N_18438,N_18291,N_18288);
and U18439 (N_18439,N_18301,N_18389);
and U18440 (N_18440,N_18372,N_18311);
nor U18441 (N_18441,N_18316,N_18349);
nand U18442 (N_18442,N_18359,N_18329);
or U18443 (N_18443,N_18295,N_18252);
xor U18444 (N_18444,N_18354,N_18263);
and U18445 (N_18445,N_18383,N_18348);
and U18446 (N_18446,N_18368,N_18388);
or U18447 (N_18447,N_18261,N_18346);
or U18448 (N_18448,N_18367,N_18399);
or U18449 (N_18449,N_18245,N_18287);
nor U18450 (N_18450,N_18249,N_18309);
and U18451 (N_18451,N_18398,N_18286);
or U18452 (N_18452,N_18257,N_18341);
nand U18453 (N_18453,N_18350,N_18273);
and U18454 (N_18454,N_18331,N_18302);
nor U18455 (N_18455,N_18275,N_18246);
or U18456 (N_18456,N_18365,N_18285);
or U18457 (N_18457,N_18280,N_18256);
xnor U18458 (N_18458,N_18293,N_18339);
and U18459 (N_18459,N_18381,N_18371);
or U18460 (N_18460,N_18262,N_18276);
and U18461 (N_18461,N_18253,N_18343);
nor U18462 (N_18462,N_18380,N_18255);
nor U18463 (N_18463,N_18281,N_18364);
nor U18464 (N_18464,N_18352,N_18384);
or U18465 (N_18465,N_18300,N_18351);
xnor U18466 (N_18466,N_18248,N_18258);
nand U18467 (N_18467,N_18283,N_18335);
and U18468 (N_18468,N_18361,N_18378);
or U18469 (N_18469,N_18297,N_18334);
xor U18470 (N_18470,N_18282,N_18307);
nor U18471 (N_18471,N_18272,N_18321);
nor U18472 (N_18472,N_18377,N_18240);
or U18473 (N_18473,N_18265,N_18310);
or U18474 (N_18474,N_18324,N_18382);
and U18475 (N_18475,N_18313,N_18269);
nor U18476 (N_18476,N_18392,N_18277);
nand U18477 (N_18477,N_18296,N_18289);
xnor U18478 (N_18478,N_18323,N_18376);
nor U18479 (N_18479,N_18284,N_18373);
nand U18480 (N_18480,N_18297,N_18338);
xnor U18481 (N_18481,N_18334,N_18242);
xor U18482 (N_18482,N_18310,N_18381);
and U18483 (N_18483,N_18280,N_18336);
nand U18484 (N_18484,N_18393,N_18385);
nor U18485 (N_18485,N_18392,N_18388);
and U18486 (N_18486,N_18285,N_18275);
xor U18487 (N_18487,N_18267,N_18326);
and U18488 (N_18488,N_18372,N_18284);
or U18489 (N_18489,N_18392,N_18395);
and U18490 (N_18490,N_18302,N_18304);
xor U18491 (N_18491,N_18293,N_18335);
and U18492 (N_18492,N_18325,N_18386);
nor U18493 (N_18493,N_18370,N_18311);
xnor U18494 (N_18494,N_18272,N_18358);
and U18495 (N_18495,N_18393,N_18276);
xor U18496 (N_18496,N_18378,N_18394);
or U18497 (N_18497,N_18259,N_18279);
nor U18498 (N_18498,N_18344,N_18328);
or U18499 (N_18499,N_18366,N_18267);
nand U18500 (N_18500,N_18369,N_18306);
or U18501 (N_18501,N_18285,N_18387);
xor U18502 (N_18502,N_18302,N_18326);
nor U18503 (N_18503,N_18279,N_18334);
nand U18504 (N_18504,N_18249,N_18262);
nand U18505 (N_18505,N_18294,N_18246);
nand U18506 (N_18506,N_18329,N_18285);
xnor U18507 (N_18507,N_18314,N_18241);
nor U18508 (N_18508,N_18388,N_18321);
nor U18509 (N_18509,N_18350,N_18362);
and U18510 (N_18510,N_18264,N_18299);
and U18511 (N_18511,N_18327,N_18283);
xnor U18512 (N_18512,N_18249,N_18393);
nand U18513 (N_18513,N_18360,N_18399);
xor U18514 (N_18514,N_18264,N_18378);
xor U18515 (N_18515,N_18318,N_18262);
xor U18516 (N_18516,N_18353,N_18338);
and U18517 (N_18517,N_18378,N_18368);
and U18518 (N_18518,N_18359,N_18395);
nor U18519 (N_18519,N_18360,N_18368);
nand U18520 (N_18520,N_18251,N_18365);
and U18521 (N_18521,N_18323,N_18365);
nor U18522 (N_18522,N_18255,N_18370);
and U18523 (N_18523,N_18366,N_18308);
nand U18524 (N_18524,N_18305,N_18388);
and U18525 (N_18525,N_18250,N_18243);
nand U18526 (N_18526,N_18286,N_18342);
and U18527 (N_18527,N_18321,N_18278);
and U18528 (N_18528,N_18381,N_18337);
and U18529 (N_18529,N_18266,N_18323);
xnor U18530 (N_18530,N_18318,N_18322);
nand U18531 (N_18531,N_18346,N_18303);
and U18532 (N_18532,N_18303,N_18332);
xnor U18533 (N_18533,N_18324,N_18377);
or U18534 (N_18534,N_18282,N_18357);
and U18535 (N_18535,N_18326,N_18339);
nor U18536 (N_18536,N_18383,N_18290);
nand U18537 (N_18537,N_18367,N_18372);
xnor U18538 (N_18538,N_18249,N_18392);
or U18539 (N_18539,N_18360,N_18362);
xnor U18540 (N_18540,N_18390,N_18346);
xor U18541 (N_18541,N_18283,N_18339);
or U18542 (N_18542,N_18339,N_18269);
or U18543 (N_18543,N_18274,N_18365);
nor U18544 (N_18544,N_18264,N_18256);
and U18545 (N_18545,N_18318,N_18240);
nand U18546 (N_18546,N_18328,N_18287);
or U18547 (N_18547,N_18298,N_18254);
nor U18548 (N_18548,N_18280,N_18349);
nor U18549 (N_18549,N_18320,N_18396);
or U18550 (N_18550,N_18276,N_18312);
and U18551 (N_18551,N_18377,N_18276);
or U18552 (N_18552,N_18379,N_18368);
nor U18553 (N_18553,N_18310,N_18293);
nand U18554 (N_18554,N_18276,N_18244);
nand U18555 (N_18555,N_18277,N_18382);
and U18556 (N_18556,N_18306,N_18364);
and U18557 (N_18557,N_18338,N_18242);
nor U18558 (N_18558,N_18275,N_18346);
and U18559 (N_18559,N_18287,N_18380);
or U18560 (N_18560,N_18488,N_18400);
nor U18561 (N_18561,N_18419,N_18480);
and U18562 (N_18562,N_18461,N_18489);
nand U18563 (N_18563,N_18433,N_18472);
or U18564 (N_18564,N_18492,N_18463);
or U18565 (N_18565,N_18430,N_18431);
or U18566 (N_18566,N_18432,N_18415);
xnor U18567 (N_18567,N_18558,N_18478);
and U18568 (N_18568,N_18505,N_18538);
nand U18569 (N_18569,N_18493,N_18508);
nor U18570 (N_18570,N_18531,N_18451);
and U18571 (N_18571,N_18479,N_18513);
nor U18572 (N_18572,N_18462,N_18526);
and U18573 (N_18573,N_18555,N_18522);
or U18574 (N_18574,N_18436,N_18409);
or U18575 (N_18575,N_18429,N_18426);
and U18576 (N_18576,N_18427,N_18511);
or U18577 (N_18577,N_18536,N_18425);
nand U18578 (N_18578,N_18404,N_18546);
or U18579 (N_18579,N_18456,N_18403);
xor U18580 (N_18580,N_18541,N_18539);
nand U18581 (N_18581,N_18442,N_18540);
xor U18582 (N_18582,N_18501,N_18500);
nand U18583 (N_18583,N_18533,N_18527);
or U18584 (N_18584,N_18421,N_18552);
and U18585 (N_18585,N_18422,N_18407);
nand U18586 (N_18586,N_18460,N_18510);
or U18587 (N_18587,N_18498,N_18455);
nand U18588 (N_18588,N_18499,N_18543);
and U18589 (N_18589,N_18506,N_18524);
and U18590 (N_18590,N_18514,N_18444);
or U18591 (N_18591,N_18529,N_18483);
nand U18592 (N_18592,N_18475,N_18466);
and U18593 (N_18593,N_18532,N_18523);
and U18594 (N_18594,N_18509,N_18447);
nand U18595 (N_18595,N_18520,N_18530);
nor U18596 (N_18596,N_18474,N_18502);
nor U18597 (N_18597,N_18519,N_18553);
or U18598 (N_18598,N_18458,N_18402);
or U18599 (N_18599,N_18469,N_18438);
nor U18600 (N_18600,N_18428,N_18481);
nand U18601 (N_18601,N_18476,N_18494);
xor U18602 (N_18602,N_18468,N_18551);
or U18603 (N_18603,N_18534,N_18512);
xnor U18604 (N_18604,N_18441,N_18401);
and U18605 (N_18605,N_18547,N_18549);
and U18606 (N_18606,N_18504,N_18424);
or U18607 (N_18607,N_18423,N_18477);
and U18608 (N_18608,N_18414,N_18454);
nor U18609 (N_18609,N_18471,N_18515);
nor U18610 (N_18610,N_18443,N_18557);
and U18611 (N_18611,N_18491,N_18405);
nor U18612 (N_18612,N_18434,N_18452);
xor U18613 (N_18613,N_18417,N_18503);
nand U18614 (N_18614,N_18554,N_18449);
nand U18615 (N_18615,N_18459,N_18495);
nand U18616 (N_18616,N_18559,N_18440);
and U18617 (N_18617,N_18439,N_18545);
xor U18618 (N_18618,N_18418,N_18446);
or U18619 (N_18619,N_18420,N_18516);
xnor U18620 (N_18620,N_18408,N_18416);
and U18621 (N_18621,N_18537,N_18435);
or U18622 (N_18622,N_18437,N_18486);
or U18623 (N_18623,N_18517,N_18411);
or U18624 (N_18624,N_18482,N_18556);
xor U18625 (N_18625,N_18535,N_18490);
xor U18626 (N_18626,N_18542,N_18487);
nor U18627 (N_18627,N_18485,N_18496);
or U18628 (N_18628,N_18484,N_18550);
nand U18629 (N_18629,N_18445,N_18521);
nor U18630 (N_18630,N_18470,N_18548);
nand U18631 (N_18631,N_18413,N_18473);
xor U18632 (N_18632,N_18497,N_18518);
or U18633 (N_18633,N_18450,N_18457);
nor U18634 (N_18634,N_18448,N_18453);
xor U18635 (N_18635,N_18406,N_18410);
or U18636 (N_18636,N_18465,N_18544);
and U18637 (N_18637,N_18528,N_18467);
xor U18638 (N_18638,N_18525,N_18507);
or U18639 (N_18639,N_18412,N_18464);
or U18640 (N_18640,N_18533,N_18455);
and U18641 (N_18641,N_18513,N_18550);
and U18642 (N_18642,N_18469,N_18543);
nor U18643 (N_18643,N_18501,N_18516);
nand U18644 (N_18644,N_18464,N_18523);
and U18645 (N_18645,N_18455,N_18479);
and U18646 (N_18646,N_18552,N_18485);
nand U18647 (N_18647,N_18460,N_18526);
nor U18648 (N_18648,N_18469,N_18478);
nand U18649 (N_18649,N_18540,N_18553);
and U18650 (N_18650,N_18442,N_18420);
or U18651 (N_18651,N_18526,N_18466);
nor U18652 (N_18652,N_18458,N_18559);
nand U18653 (N_18653,N_18546,N_18540);
xor U18654 (N_18654,N_18478,N_18551);
or U18655 (N_18655,N_18503,N_18532);
nand U18656 (N_18656,N_18480,N_18497);
nand U18657 (N_18657,N_18508,N_18464);
nand U18658 (N_18658,N_18408,N_18449);
nand U18659 (N_18659,N_18540,N_18491);
nand U18660 (N_18660,N_18554,N_18513);
and U18661 (N_18661,N_18512,N_18432);
xor U18662 (N_18662,N_18431,N_18505);
nand U18663 (N_18663,N_18537,N_18510);
nor U18664 (N_18664,N_18519,N_18449);
and U18665 (N_18665,N_18463,N_18493);
nand U18666 (N_18666,N_18550,N_18482);
nand U18667 (N_18667,N_18462,N_18520);
or U18668 (N_18668,N_18523,N_18429);
and U18669 (N_18669,N_18461,N_18439);
and U18670 (N_18670,N_18548,N_18433);
or U18671 (N_18671,N_18438,N_18459);
and U18672 (N_18672,N_18548,N_18450);
xnor U18673 (N_18673,N_18419,N_18453);
nand U18674 (N_18674,N_18479,N_18459);
nor U18675 (N_18675,N_18455,N_18435);
or U18676 (N_18676,N_18452,N_18464);
or U18677 (N_18677,N_18442,N_18498);
or U18678 (N_18678,N_18446,N_18413);
nand U18679 (N_18679,N_18539,N_18402);
nand U18680 (N_18680,N_18485,N_18459);
nor U18681 (N_18681,N_18473,N_18509);
and U18682 (N_18682,N_18493,N_18435);
nand U18683 (N_18683,N_18445,N_18449);
nand U18684 (N_18684,N_18495,N_18468);
nand U18685 (N_18685,N_18459,N_18491);
nor U18686 (N_18686,N_18423,N_18531);
nor U18687 (N_18687,N_18531,N_18407);
or U18688 (N_18688,N_18514,N_18441);
or U18689 (N_18689,N_18483,N_18445);
xor U18690 (N_18690,N_18427,N_18463);
xor U18691 (N_18691,N_18443,N_18452);
and U18692 (N_18692,N_18511,N_18433);
nand U18693 (N_18693,N_18471,N_18434);
nand U18694 (N_18694,N_18486,N_18533);
and U18695 (N_18695,N_18414,N_18499);
nor U18696 (N_18696,N_18400,N_18489);
and U18697 (N_18697,N_18423,N_18408);
nor U18698 (N_18698,N_18539,N_18520);
nand U18699 (N_18699,N_18446,N_18435);
nor U18700 (N_18700,N_18484,N_18437);
and U18701 (N_18701,N_18536,N_18498);
xnor U18702 (N_18702,N_18486,N_18464);
xor U18703 (N_18703,N_18557,N_18543);
nand U18704 (N_18704,N_18480,N_18435);
and U18705 (N_18705,N_18427,N_18496);
or U18706 (N_18706,N_18504,N_18463);
nand U18707 (N_18707,N_18555,N_18501);
nor U18708 (N_18708,N_18494,N_18418);
xnor U18709 (N_18709,N_18547,N_18545);
or U18710 (N_18710,N_18414,N_18400);
xor U18711 (N_18711,N_18526,N_18489);
and U18712 (N_18712,N_18417,N_18536);
xor U18713 (N_18713,N_18476,N_18479);
and U18714 (N_18714,N_18553,N_18460);
or U18715 (N_18715,N_18514,N_18557);
or U18716 (N_18716,N_18479,N_18526);
nand U18717 (N_18717,N_18551,N_18500);
nor U18718 (N_18718,N_18446,N_18491);
or U18719 (N_18719,N_18443,N_18459);
or U18720 (N_18720,N_18596,N_18647);
xnor U18721 (N_18721,N_18671,N_18636);
or U18722 (N_18722,N_18687,N_18682);
and U18723 (N_18723,N_18608,N_18703);
xor U18724 (N_18724,N_18628,N_18654);
or U18725 (N_18725,N_18649,N_18572);
and U18726 (N_18726,N_18640,N_18614);
xnor U18727 (N_18727,N_18639,N_18663);
and U18728 (N_18728,N_18587,N_18627);
or U18729 (N_18729,N_18561,N_18588);
nor U18730 (N_18730,N_18610,N_18659);
and U18731 (N_18731,N_18668,N_18599);
xor U18732 (N_18732,N_18680,N_18714);
xnor U18733 (N_18733,N_18672,N_18591);
nor U18734 (N_18734,N_18667,N_18597);
nand U18735 (N_18735,N_18602,N_18645);
and U18736 (N_18736,N_18616,N_18653);
nor U18737 (N_18737,N_18716,N_18704);
and U18738 (N_18738,N_18643,N_18692);
xor U18739 (N_18739,N_18590,N_18560);
xnor U18740 (N_18740,N_18658,N_18573);
and U18741 (N_18741,N_18575,N_18635);
nand U18742 (N_18742,N_18622,N_18691);
and U18743 (N_18743,N_18706,N_18710);
xor U18744 (N_18744,N_18630,N_18601);
nor U18745 (N_18745,N_18565,N_18581);
xnor U18746 (N_18746,N_18656,N_18702);
nand U18747 (N_18747,N_18563,N_18583);
xnor U18748 (N_18748,N_18626,N_18567);
xor U18749 (N_18749,N_18677,N_18688);
and U18750 (N_18750,N_18638,N_18634);
xnor U18751 (N_18751,N_18684,N_18611);
nor U18752 (N_18752,N_18662,N_18718);
xor U18753 (N_18753,N_18595,N_18582);
or U18754 (N_18754,N_18679,N_18577);
and U18755 (N_18755,N_18644,N_18570);
or U18756 (N_18756,N_18696,N_18642);
and U18757 (N_18757,N_18629,N_18651);
and U18758 (N_18758,N_18600,N_18632);
and U18759 (N_18759,N_18661,N_18657);
nand U18760 (N_18760,N_18619,N_18613);
xnor U18761 (N_18761,N_18631,N_18686);
nand U18762 (N_18762,N_18604,N_18695);
and U18763 (N_18763,N_18670,N_18697);
or U18764 (N_18764,N_18675,N_18719);
or U18765 (N_18765,N_18698,N_18579);
nor U18766 (N_18766,N_18689,N_18593);
nor U18767 (N_18767,N_18641,N_18609);
nor U18768 (N_18768,N_18694,N_18574);
or U18769 (N_18769,N_18566,N_18598);
nand U18770 (N_18770,N_18650,N_18713);
or U18771 (N_18771,N_18664,N_18625);
nor U18772 (N_18772,N_18615,N_18646);
nand U18773 (N_18773,N_18594,N_18683);
or U18774 (N_18774,N_18569,N_18711);
nand U18775 (N_18775,N_18568,N_18621);
or U18776 (N_18776,N_18580,N_18701);
or U18777 (N_18777,N_18674,N_18633);
nor U18778 (N_18778,N_18578,N_18617);
or U18779 (N_18779,N_18709,N_18612);
nor U18780 (N_18780,N_18584,N_18715);
xor U18781 (N_18781,N_18623,N_18571);
nand U18782 (N_18782,N_18707,N_18652);
or U18783 (N_18783,N_18592,N_18589);
nor U18784 (N_18784,N_18562,N_18690);
and U18785 (N_18785,N_18607,N_18576);
nor U18786 (N_18786,N_18685,N_18666);
and U18787 (N_18787,N_18673,N_18693);
nor U18788 (N_18788,N_18681,N_18606);
and U18789 (N_18789,N_18669,N_18564);
nand U18790 (N_18790,N_18605,N_18603);
or U18791 (N_18791,N_18708,N_18717);
and U18792 (N_18792,N_18678,N_18676);
nor U18793 (N_18793,N_18637,N_18699);
nand U18794 (N_18794,N_18655,N_18712);
nand U18795 (N_18795,N_18660,N_18665);
and U18796 (N_18796,N_18624,N_18705);
and U18797 (N_18797,N_18585,N_18618);
nand U18798 (N_18798,N_18648,N_18620);
or U18799 (N_18799,N_18586,N_18700);
or U18800 (N_18800,N_18638,N_18664);
and U18801 (N_18801,N_18688,N_18692);
xor U18802 (N_18802,N_18673,N_18698);
nand U18803 (N_18803,N_18568,N_18676);
and U18804 (N_18804,N_18659,N_18626);
or U18805 (N_18805,N_18633,N_18699);
nor U18806 (N_18806,N_18684,N_18705);
nor U18807 (N_18807,N_18675,N_18708);
nand U18808 (N_18808,N_18688,N_18681);
and U18809 (N_18809,N_18622,N_18583);
and U18810 (N_18810,N_18628,N_18588);
nand U18811 (N_18811,N_18719,N_18563);
nor U18812 (N_18812,N_18655,N_18647);
nand U18813 (N_18813,N_18690,N_18564);
and U18814 (N_18814,N_18571,N_18583);
nand U18815 (N_18815,N_18675,N_18693);
or U18816 (N_18816,N_18634,N_18665);
nor U18817 (N_18817,N_18582,N_18692);
or U18818 (N_18818,N_18611,N_18695);
nor U18819 (N_18819,N_18567,N_18584);
nand U18820 (N_18820,N_18659,N_18604);
xor U18821 (N_18821,N_18682,N_18681);
nand U18822 (N_18822,N_18574,N_18699);
nand U18823 (N_18823,N_18650,N_18702);
and U18824 (N_18824,N_18564,N_18573);
and U18825 (N_18825,N_18580,N_18606);
and U18826 (N_18826,N_18677,N_18691);
nand U18827 (N_18827,N_18642,N_18662);
xnor U18828 (N_18828,N_18644,N_18718);
xor U18829 (N_18829,N_18707,N_18702);
or U18830 (N_18830,N_18689,N_18647);
or U18831 (N_18831,N_18677,N_18681);
or U18832 (N_18832,N_18701,N_18647);
xnor U18833 (N_18833,N_18637,N_18687);
and U18834 (N_18834,N_18628,N_18580);
or U18835 (N_18835,N_18687,N_18719);
or U18836 (N_18836,N_18581,N_18677);
nand U18837 (N_18837,N_18688,N_18575);
and U18838 (N_18838,N_18613,N_18576);
or U18839 (N_18839,N_18644,N_18686);
xnor U18840 (N_18840,N_18621,N_18678);
nor U18841 (N_18841,N_18638,N_18609);
or U18842 (N_18842,N_18686,N_18650);
nand U18843 (N_18843,N_18614,N_18587);
and U18844 (N_18844,N_18653,N_18602);
nor U18845 (N_18845,N_18564,N_18707);
nand U18846 (N_18846,N_18675,N_18646);
xor U18847 (N_18847,N_18639,N_18568);
or U18848 (N_18848,N_18582,N_18625);
nand U18849 (N_18849,N_18660,N_18565);
xor U18850 (N_18850,N_18575,N_18578);
xnor U18851 (N_18851,N_18697,N_18690);
xnor U18852 (N_18852,N_18610,N_18572);
nor U18853 (N_18853,N_18592,N_18658);
nand U18854 (N_18854,N_18586,N_18689);
or U18855 (N_18855,N_18574,N_18580);
nand U18856 (N_18856,N_18641,N_18677);
and U18857 (N_18857,N_18639,N_18681);
nand U18858 (N_18858,N_18572,N_18655);
xnor U18859 (N_18859,N_18680,N_18657);
nand U18860 (N_18860,N_18587,N_18694);
and U18861 (N_18861,N_18632,N_18634);
xor U18862 (N_18862,N_18696,N_18677);
or U18863 (N_18863,N_18663,N_18570);
and U18864 (N_18864,N_18560,N_18602);
nand U18865 (N_18865,N_18605,N_18571);
xor U18866 (N_18866,N_18597,N_18633);
nor U18867 (N_18867,N_18570,N_18667);
or U18868 (N_18868,N_18609,N_18656);
and U18869 (N_18869,N_18585,N_18604);
nor U18870 (N_18870,N_18601,N_18684);
nor U18871 (N_18871,N_18601,N_18636);
nand U18872 (N_18872,N_18573,N_18630);
or U18873 (N_18873,N_18707,N_18649);
and U18874 (N_18874,N_18641,N_18570);
xnor U18875 (N_18875,N_18596,N_18650);
xnor U18876 (N_18876,N_18697,N_18604);
xnor U18877 (N_18877,N_18682,N_18656);
xor U18878 (N_18878,N_18598,N_18692);
and U18879 (N_18879,N_18594,N_18573);
xor U18880 (N_18880,N_18819,N_18755);
nand U18881 (N_18881,N_18802,N_18879);
or U18882 (N_18882,N_18731,N_18836);
nand U18883 (N_18883,N_18835,N_18740);
nand U18884 (N_18884,N_18831,N_18815);
and U18885 (N_18885,N_18871,N_18766);
xor U18886 (N_18886,N_18807,N_18813);
and U18887 (N_18887,N_18775,N_18735);
and U18888 (N_18888,N_18850,N_18805);
nand U18889 (N_18889,N_18771,N_18856);
and U18890 (N_18890,N_18841,N_18812);
nor U18891 (N_18891,N_18840,N_18722);
nand U18892 (N_18892,N_18876,N_18833);
nor U18893 (N_18893,N_18866,N_18848);
nor U18894 (N_18894,N_18846,N_18858);
xor U18895 (N_18895,N_18830,N_18769);
or U18896 (N_18896,N_18875,N_18809);
nand U18897 (N_18897,N_18730,N_18758);
or U18898 (N_18898,N_18803,N_18794);
or U18899 (N_18899,N_18847,N_18745);
nand U18900 (N_18900,N_18791,N_18763);
nor U18901 (N_18901,N_18768,N_18734);
or U18902 (N_18902,N_18726,N_18754);
and U18903 (N_18903,N_18849,N_18743);
xnor U18904 (N_18904,N_18787,N_18720);
and U18905 (N_18905,N_18783,N_18786);
or U18906 (N_18906,N_18854,N_18877);
or U18907 (N_18907,N_18762,N_18798);
nand U18908 (N_18908,N_18744,N_18861);
and U18909 (N_18909,N_18764,N_18761);
xor U18910 (N_18910,N_18772,N_18864);
nand U18911 (N_18911,N_18827,N_18778);
nand U18912 (N_18912,N_18739,N_18797);
nor U18913 (N_18913,N_18808,N_18873);
nor U18914 (N_18914,N_18752,N_18865);
nand U18915 (N_18915,N_18723,N_18855);
nand U18916 (N_18916,N_18821,N_18784);
nand U18917 (N_18917,N_18837,N_18795);
nor U18918 (N_18918,N_18838,N_18728);
nand U18919 (N_18919,N_18851,N_18878);
nand U18920 (N_18920,N_18776,N_18779);
nor U18921 (N_18921,N_18828,N_18750);
nand U18922 (N_18922,N_18844,N_18818);
nand U18923 (N_18923,N_18814,N_18872);
or U18924 (N_18924,N_18843,N_18780);
and U18925 (N_18925,N_18868,N_18767);
nor U18926 (N_18926,N_18816,N_18825);
and U18927 (N_18927,N_18742,N_18770);
and U18928 (N_18928,N_18870,N_18845);
and U18929 (N_18929,N_18773,N_18806);
or U18930 (N_18930,N_18792,N_18869);
or U18931 (N_18931,N_18777,N_18810);
nand U18932 (N_18932,N_18747,N_18824);
nand U18933 (N_18933,N_18751,N_18832);
nand U18934 (N_18934,N_18748,N_18817);
and U18935 (N_18935,N_18721,N_18741);
and U18936 (N_18936,N_18732,N_18782);
and U18937 (N_18937,N_18829,N_18863);
and U18938 (N_18938,N_18725,N_18799);
nand U18939 (N_18939,N_18826,N_18834);
xnor U18940 (N_18940,N_18800,N_18867);
xor U18941 (N_18941,N_18811,N_18781);
xnor U18942 (N_18942,N_18862,N_18796);
nand U18943 (N_18943,N_18839,N_18760);
xor U18944 (N_18944,N_18729,N_18790);
or U18945 (N_18945,N_18789,N_18765);
nand U18946 (N_18946,N_18853,N_18727);
and U18947 (N_18947,N_18820,N_18822);
xor U18948 (N_18948,N_18801,N_18874);
nand U18949 (N_18949,N_18860,N_18736);
nor U18950 (N_18950,N_18737,N_18774);
and U18951 (N_18951,N_18788,N_18759);
nand U18952 (N_18952,N_18738,N_18746);
xor U18953 (N_18953,N_18842,N_18757);
xor U18954 (N_18954,N_18804,N_18859);
or U18955 (N_18955,N_18733,N_18857);
nor U18956 (N_18956,N_18753,N_18852);
nor U18957 (N_18957,N_18756,N_18785);
and U18958 (N_18958,N_18793,N_18823);
nand U18959 (N_18959,N_18724,N_18749);
and U18960 (N_18960,N_18730,N_18774);
xor U18961 (N_18961,N_18873,N_18737);
or U18962 (N_18962,N_18777,N_18747);
nand U18963 (N_18963,N_18869,N_18722);
and U18964 (N_18964,N_18763,N_18752);
nor U18965 (N_18965,N_18744,N_18803);
nor U18966 (N_18966,N_18741,N_18846);
or U18967 (N_18967,N_18815,N_18724);
xnor U18968 (N_18968,N_18733,N_18753);
xor U18969 (N_18969,N_18766,N_18764);
nor U18970 (N_18970,N_18842,N_18847);
or U18971 (N_18971,N_18821,N_18741);
xnor U18972 (N_18972,N_18857,N_18798);
or U18973 (N_18973,N_18876,N_18840);
or U18974 (N_18974,N_18751,N_18782);
nor U18975 (N_18975,N_18832,N_18868);
xor U18976 (N_18976,N_18760,N_18816);
nand U18977 (N_18977,N_18860,N_18829);
nor U18978 (N_18978,N_18867,N_18725);
nor U18979 (N_18979,N_18747,N_18796);
nand U18980 (N_18980,N_18806,N_18805);
nor U18981 (N_18981,N_18817,N_18874);
nor U18982 (N_18982,N_18835,N_18879);
xnor U18983 (N_18983,N_18721,N_18764);
xnor U18984 (N_18984,N_18856,N_18871);
nand U18985 (N_18985,N_18862,N_18764);
nor U18986 (N_18986,N_18740,N_18727);
and U18987 (N_18987,N_18720,N_18868);
nand U18988 (N_18988,N_18811,N_18775);
and U18989 (N_18989,N_18792,N_18764);
nor U18990 (N_18990,N_18872,N_18746);
nand U18991 (N_18991,N_18761,N_18871);
nand U18992 (N_18992,N_18841,N_18824);
and U18993 (N_18993,N_18848,N_18741);
nand U18994 (N_18994,N_18766,N_18787);
nand U18995 (N_18995,N_18879,N_18763);
nand U18996 (N_18996,N_18841,N_18783);
nor U18997 (N_18997,N_18827,N_18742);
xor U18998 (N_18998,N_18820,N_18831);
and U18999 (N_18999,N_18814,N_18840);
xor U19000 (N_19000,N_18796,N_18746);
xor U19001 (N_19001,N_18833,N_18838);
and U19002 (N_19002,N_18783,N_18772);
xnor U19003 (N_19003,N_18843,N_18728);
nand U19004 (N_19004,N_18869,N_18859);
and U19005 (N_19005,N_18856,N_18861);
and U19006 (N_19006,N_18781,N_18834);
and U19007 (N_19007,N_18869,N_18841);
and U19008 (N_19008,N_18854,N_18773);
or U19009 (N_19009,N_18753,N_18799);
xor U19010 (N_19010,N_18750,N_18729);
nor U19011 (N_19011,N_18814,N_18861);
or U19012 (N_19012,N_18741,N_18793);
nand U19013 (N_19013,N_18753,N_18853);
and U19014 (N_19014,N_18759,N_18800);
xnor U19015 (N_19015,N_18732,N_18791);
nand U19016 (N_19016,N_18760,N_18815);
nor U19017 (N_19017,N_18848,N_18726);
xor U19018 (N_19018,N_18850,N_18843);
nand U19019 (N_19019,N_18826,N_18798);
xor U19020 (N_19020,N_18845,N_18774);
nor U19021 (N_19021,N_18768,N_18826);
nand U19022 (N_19022,N_18757,N_18722);
or U19023 (N_19023,N_18850,N_18724);
nand U19024 (N_19024,N_18748,N_18862);
xor U19025 (N_19025,N_18774,N_18781);
nand U19026 (N_19026,N_18871,N_18767);
or U19027 (N_19027,N_18792,N_18850);
nor U19028 (N_19028,N_18811,N_18821);
and U19029 (N_19029,N_18857,N_18800);
or U19030 (N_19030,N_18864,N_18855);
nand U19031 (N_19031,N_18793,N_18865);
xor U19032 (N_19032,N_18849,N_18729);
nand U19033 (N_19033,N_18851,N_18854);
and U19034 (N_19034,N_18833,N_18866);
nand U19035 (N_19035,N_18820,N_18836);
and U19036 (N_19036,N_18866,N_18786);
and U19037 (N_19037,N_18750,N_18831);
xnor U19038 (N_19038,N_18733,N_18800);
nand U19039 (N_19039,N_18839,N_18837);
or U19040 (N_19040,N_18972,N_19035);
and U19041 (N_19041,N_19030,N_18883);
nor U19042 (N_19042,N_18931,N_19023);
xor U19043 (N_19043,N_18955,N_19033);
xnor U19044 (N_19044,N_18950,N_19034);
nor U19045 (N_19045,N_18942,N_18916);
or U19046 (N_19046,N_18983,N_18894);
nand U19047 (N_19047,N_18893,N_18964);
and U19048 (N_19048,N_18949,N_19018);
and U19049 (N_19049,N_18988,N_18882);
nand U19050 (N_19050,N_18938,N_18901);
and U19051 (N_19051,N_19012,N_19022);
nand U19052 (N_19052,N_18929,N_18923);
nand U19053 (N_19053,N_18948,N_18935);
nor U19054 (N_19054,N_19020,N_18885);
xnor U19055 (N_19055,N_18984,N_18939);
and U19056 (N_19056,N_19006,N_18921);
or U19057 (N_19057,N_18937,N_18986);
and U19058 (N_19058,N_18928,N_18979);
nand U19059 (N_19059,N_18903,N_19039);
nand U19060 (N_19060,N_18975,N_19038);
nor U19061 (N_19061,N_19010,N_18902);
nand U19062 (N_19062,N_18973,N_19029);
xor U19063 (N_19063,N_19005,N_18980);
or U19064 (N_19064,N_18884,N_18998);
or U19065 (N_19065,N_18989,N_18914);
or U19066 (N_19066,N_18888,N_18974);
nand U19067 (N_19067,N_18995,N_18991);
nand U19068 (N_19068,N_18992,N_19032);
xnor U19069 (N_19069,N_18907,N_18892);
nor U19070 (N_19070,N_18904,N_18911);
or U19071 (N_19071,N_18943,N_18970);
xnor U19072 (N_19072,N_18999,N_18997);
nor U19073 (N_19073,N_18971,N_18957);
nand U19074 (N_19074,N_19013,N_18941);
xnor U19075 (N_19075,N_18954,N_18908);
and U19076 (N_19076,N_18951,N_18880);
nand U19077 (N_19077,N_18946,N_18889);
nand U19078 (N_19078,N_18944,N_18900);
nand U19079 (N_19079,N_18982,N_18912);
xor U19080 (N_19080,N_19003,N_18936);
xor U19081 (N_19081,N_18963,N_18994);
nor U19082 (N_19082,N_19000,N_19021);
xnor U19083 (N_19083,N_18961,N_19031);
or U19084 (N_19084,N_18958,N_18952);
nor U19085 (N_19085,N_18940,N_18966);
or U19086 (N_19086,N_18917,N_18896);
or U19087 (N_19087,N_18985,N_19009);
or U19088 (N_19088,N_19004,N_18990);
and U19089 (N_19089,N_18897,N_19037);
xor U19090 (N_19090,N_18967,N_18932);
and U19091 (N_19091,N_18947,N_18898);
nor U19092 (N_19092,N_18993,N_19008);
xnor U19093 (N_19093,N_18996,N_18881);
xnor U19094 (N_19094,N_18913,N_18906);
or U19095 (N_19095,N_18905,N_18977);
nand U19096 (N_19096,N_18981,N_19026);
nor U19097 (N_19097,N_18925,N_18895);
xor U19098 (N_19098,N_18926,N_19019);
and U19099 (N_19099,N_18969,N_18959);
or U19100 (N_19100,N_18956,N_19015);
nand U19101 (N_19101,N_18945,N_19007);
xnor U19102 (N_19102,N_18978,N_18930);
nand U19103 (N_19103,N_18909,N_18953);
and U19104 (N_19104,N_18960,N_19017);
or U19105 (N_19105,N_18927,N_18968);
or U19106 (N_19106,N_18976,N_18899);
and U19107 (N_19107,N_18933,N_18924);
nand U19108 (N_19108,N_19001,N_19011);
and U19109 (N_19109,N_18887,N_19002);
and U19110 (N_19110,N_19025,N_18918);
nor U19111 (N_19111,N_19036,N_18886);
or U19112 (N_19112,N_18987,N_18934);
nand U19113 (N_19113,N_18890,N_18965);
xnor U19114 (N_19114,N_19024,N_18915);
and U19115 (N_19115,N_18920,N_18922);
xor U19116 (N_19116,N_18910,N_19028);
and U19117 (N_19117,N_19016,N_18962);
and U19118 (N_19118,N_18919,N_19027);
xnor U19119 (N_19119,N_18891,N_19014);
nand U19120 (N_19120,N_18888,N_18905);
xnor U19121 (N_19121,N_18910,N_18971);
and U19122 (N_19122,N_18883,N_18956);
xnor U19123 (N_19123,N_18917,N_18890);
and U19124 (N_19124,N_18897,N_18918);
or U19125 (N_19125,N_19031,N_18948);
and U19126 (N_19126,N_18914,N_18983);
and U19127 (N_19127,N_18886,N_18909);
xnor U19128 (N_19128,N_18902,N_18919);
nor U19129 (N_19129,N_18896,N_18890);
and U19130 (N_19130,N_18884,N_19028);
and U19131 (N_19131,N_18927,N_18956);
or U19132 (N_19132,N_18962,N_18928);
xnor U19133 (N_19133,N_18910,N_18949);
nor U19134 (N_19134,N_19010,N_18917);
and U19135 (N_19135,N_18900,N_19013);
or U19136 (N_19136,N_19024,N_18972);
xor U19137 (N_19137,N_19014,N_19019);
xnor U19138 (N_19138,N_18883,N_18932);
and U19139 (N_19139,N_18962,N_18947);
nor U19140 (N_19140,N_18890,N_18969);
xor U19141 (N_19141,N_18923,N_18987);
and U19142 (N_19142,N_18948,N_18921);
xnor U19143 (N_19143,N_18982,N_18927);
nand U19144 (N_19144,N_18985,N_18995);
and U19145 (N_19145,N_18957,N_18953);
nor U19146 (N_19146,N_18956,N_19003);
or U19147 (N_19147,N_19016,N_19018);
and U19148 (N_19148,N_18988,N_18935);
and U19149 (N_19149,N_18940,N_19035);
or U19150 (N_19150,N_18924,N_18935);
and U19151 (N_19151,N_18933,N_18943);
nand U19152 (N_19152,N_18929,N_18920);
nand U19153 (N_19153,N_18899,N_19037);
nand U19154 (N_19154,N_19018,N_19035);
or U19155 (N_19155,N_19007,N_19010);
or U19156 (N_19156,N_18896,N_18971);
and U19157 (N_19157,N_19014,N_19023);
nor U19158 (N_19158,N_19002,N_18948);
and U19159 (N_19159,N_19018,N_18957);
nor U19160 (N_19160,N_18896,N_18898);
or U19161 (N_19161,N_18901,N_18956);
or U19162 (N_19162,N_18988,N_19008);
nor U19163 (N_19163,N_19006,N_18991);
nor U19164 (N_19164,N_18964,N_18892);
nor U19165 (N_19165,N_18956,N_18947);
and U19166 (N_19166,N_18896,N_19010);
or U19167 (N_19167,N_18924,N_18990);
or U19168 (N_19168,N_18888,N_18967);
and U19169 (N_19169,N_18994,N_18940);
and U19170 (N_19170,N_18916,N_19035);
nand U19171 (N_19171,N_18919,N_18896);
and U19172 (N_19172,N_18982,N_18963);
and U19173 (N_19173,N_19000,N_18881);
and U19174 (N_19174,N_19008,N_18927);
nand U19175 (N_19175,N_18933,N_18955);
nor U19176 (N_19176,N_18978,N_18894);
xor U19177 (N_19177,N_19030,N_19024);
nor U19178 (N_19178,N_19014,N_19021);
or U19179 (N_19179,N_18967,N_19004);
and U19180 (N_19180,N_18934,N_19027);
and U19181 (N_19181,N_19000,N_18928);
and U19182 (N_19182,N_18927,N_18967);
nor U19183 (N_19183,N_19022,N_18907);
nor U19184 (N_19184,N_18989,N_19027);
nor U19185 (N_19185,N_18901,N_18898);
nand U19186 (N_19186,N_18889,N_18988);
nand U19187 (N_19187,N_18969,N_18988);
or U19188 (N_19188,N_18976,N_18926);
or U19189 (N_19189,N_19001,N_18941);
and U19190 (N_19190,N_18947,N_18914);
nor U19191 (N_19191,N_18963,N_19036);
nor U19192 (N_19192,N_18913,N_18961);
and U19193 (N_19193,N_18882,N_18912);
or U19194 (N_19194,N_18965,N_18975);
nand U19195 (N_19195,N_18881,N_18956);
or U19196 (N_19196,N_19014,N_18903);
xnor U19197 (N_19197,N_19003,N_18891);
and U19198 (N_19198,N_18903,N_19033);
or U19199 (N_19199,N_18981,N_18888);
nor U19200 (N_19200,N_19152,N_19055);
xnor U19201 (N_19201,N_19138,N_19048);
and U19202 (N_19202,N_19060,N_19093);
or U19203 (N_19203,N_19092,N_19086);
nor U19204 (N_19204,N_19102,N_19095);
xnor U19205 (N_19205,N_19044,N_19190);
and U19206 (N_19206,N_19150,N_19160);
nand U19207 (N_19207,N_19064,N_19046);
or U19208 (N_19208,N_19181,N_19121);
nand U19209 (N_19209,N_19104,N_19079);
xnor U19210 (N_19210,N_19103,N_19156);
nand U19211 (N_19211,N_19041,N_19059);
xnor U19212 (N_19212,N_19110,N_19051);
or U19213 (N_19213,N_19134,N_19089);
nand U19214 (N_19214,N_19180,N_19067);
and U19215 (N_19215,N_19128,N_19042);
xnor U19216 (N_19216,N_19197,N_19189);
xor U19217 (N_19217,N_19198,N_19132);
nand U19218 (N_19218,N_19043,N_19107);
and U19219 (N_19219,N_19083,N_19053);
xnor U19220 (N_19220,N_19122,N_19179);
nand U19221 (N_19221,N_19177,N_19074);
xor U19222 (N_19222,N_19101,N_19169);
nand U19223 (N_19223,N_19070,N_19105);
xor U19224 (N_19224,N_19106,N_19173);
or U19225 (N_19225,N_19088,N_19145);
nand U19226 (N_19226,N_19141,N_19115);
nor U19227 (N_19227,N_19172,N_19084);
and U19228 (N_19228,N_19195,N_19191);
and U19229 (N_19229,N_19148,N_19127);
nor U19230 (N_19230,N_19072,N_19183);
xor U19231 (N_19231,N_19096,N_19058);
nor U19232 (N_19232,N_19186,N_19119);
nor U19233 (N_19233,N_19192,N_19056);
nor U19234 (N_19234,N_19117,N_19123);
xor U19235 (N_19235,N_19143,N_19168);
nand U19236 (N_19236,N_19185,N_19193);
and U19237 (N_19237,N_19126,N_19176);
nand U19238 (N_19238,N_19184,N_19052);
nand U19239 (N_19239,N_19163,N_19165);
and U19240 (N_19240,N_19171,N_19111);
and U19241 (N_19241,N_19054,N_19133);
nand U19242 (N_19242,N_19050,N_19112);
xnor U19243 (N_19243,N_19114,N_19157);
and U19244 (N_19244,N_19175,N_19124);
nor U19245 (N_19245,N_19164,N_19167);
or U19246 (N_19246,N_19151,N_19071);
and U19247 (N_19247,N_19090,N_19142);
nand U19248 (N_19248,N_19049,N_19076);
and U19249 (N_19249,N_19188,N_19047);
or U19250 (N_19250,N_19129,N_19144);
xnor U19251 (N_19251,N_19108,N_19174);
nand U19252 (N_19252,N_19149,N_19097);
and U19253 (N_19253,N_19146,N_19082);
and U19254 (N_19254,N_19068,N_19136);
and U19255 (N_19255,N_19099,N_19194);
and U19256 (N_19256,N_19087,N_19199);
and U19257 (N_19257,N_19085,N_19120);
nand U19258 (N_19258,N_19061,N_19130);
nor U19259 (N_19259,N_19094,N_19118);
or U19260 (N_19260,N_19182,N_19062);
or U19261 (N_19261,N_19159,N_19131);
nand U19262 (N_19262,N_19081,N_19154);
or U19263 (N_19263,N_19073,N_19137);
nor U19264 (N_19264,N_19069,N_19066);
nor U19265 (N_19265,N_19116,N_19155);
xor U19266 (N_19266,N_19187,N_19153);
or U19267 (N_19267,N_19063,N_19077);
and U19268 (N_19268,N_19040,N_19078);
xnor U19269 (N_19269,N_19080,N_19139);
or U19270 (N_19270,N_19091,N_19170);
or U19271 (N_19271,N_19100,N_19065);
or U19272 (N_19272,N_19161,N_19140);
and U19273 (N_19273,N_19045,N_19098);
nor U19274 (N_19274,N_19135,N_19166);
nor U19275 (N_19275,N_19178,N_19057);
nand U19276 (N_19276,N_19113,N_19162);
nand U19277 (N_19277,N_19147,N_19196);
and U19278 (N_19278,N_19109,N_19158);
nand U19279 (N_19279,N_19125,N_19075);
or U19280 (N_19280,N_19182,N_19043);
nand U19281 (N_19281,N_19102,N_19176);
nor U19282 (N_19282,N_19123,N_19118);
or U19283 (N_19283,N_19152,N_19057);
nand U19284 (N_19284,N_19110,N_19149);
or U19285 (N_19285,N_19160,N_19133);
xnor U19286 (N_19286,N_19175,N_19057);
or U19287 (N_19287,N_19161,N_19047);
nor U19288 (N_19288,N_19073,N_19069);
nor U19289 (N_19289,N_19126,N_19046);
nand U19290 (N_19290,N_19194,N_19117);
xnor U19291 (N_19291,N_19087,N_19041);
nand U19292 (N_19292,N_19131,N_19079);
or U19293 (N_19293,N_19183,N_19171);
and U19294 (N_19294,N_19136,N_19140);
xor U19295 (N_19295,N_19146,N_19115);
nor U19296 (N_19296,N_19058,N_19044);
and U19297 (N_19297,N_19170,N_19080);
nor U19298 (N_19298,N_19090,N_19148);
or U19299 (N_19299,N_19189,N_19169);
xnor U19300 (N_19300,N_19155,N_19080);
or U19301 (N_19301,N_19043,N_19116);
nand U19302 (N_19302,N_19187,N_19127);
nand U19303 (N_19303,N_19095,N_19104);
nor U19304 (N_19304,N_19199,N_19133);
or U19305 (N_19305,N_19128,N_19052);
or U19306 (N_19306,N_19155,N_19118);
nand U19307 (N_19307,N_19099,N_19115);
nand U19308 (N_19308,N_19115,N_19118);
nand U19309 (N_19309,N_19150,N_19144);
and U19310 (N_19310,N_19195,N_19102);
nor U19311 (N_19311,N_19156,N_19145);
and U19312 (N_19312,N_19112,N_19148);
or U19313 (N_19313,N_19110,N_19132);
or U19314 (N_19314,N_19121,N_19095);
nor U19315 (N_19315,N_19139,N_19134);
or U19316 (N_19316,N_19151,N_19177);
xor U19317 (N_19317,N_19148,N_19098);
nand U19318 (N_19318,N_19156,N_19166);
or U19319 (N_19319,N_19127,N_19107);
or U19320 (N_19320,N_19141,N_19088);
or U19321 (N_19321,N_19068,N_19097);
xor U19322 (N_19322,N_19109,N_19071);
or U19323 (N_19323,N_19061,N_19164);
and U19324 (N_19324,N_19095,N_19120);
and U19325 (N_19325,N_19185,N_19198);
or U19326 (N_19326,N_19057,N_19136);
and U19327 (N_19327,N_19067,N_19171);
nand U19328 (N_19328,N_19155,N_19112);
nor U19329 (N_19329,N_19191,N_19141);
and U19330 (N_19330,N_19136,N_19073);
nand U19331 (N_19331,N_19110,N_19157);
xnor U19332 (N_19332,N_19188,N_19127);
nor U19333 (N_19333,N_19098,N_19140);
or U19334 (N_19334,N_19192,N_19092);
nand U19335 (N_19335,N_19049,N_19091);
and U19336 (N_19336,N_19165,N_19082);
nor U19337 (N_19337,N_19192,N_19102);
and U19338 (N_19338,N_19146,N_19085);
xnor U19339 (N_19339,N_19192,N_19141);
xor U19340 (N_19340,N_19075,N_19189);
nand U19341 (N_19341,N_19057,N_19142);
and U19342 (N_19342,N_19152,N_19150);
and U19343 (N_19343,N_19157,N_19072);
and U19344 (N_19344,N_19071,N_19063);
or U19345 (N_19345,N_19105,N_19107);
and U19346 (N_19346,N_19096,N_19126);
xnor U19347 (N_19347,N_19196,N_19091);
or U19348 (N_19348,N_19149,N_19045);
and U19349 (N_19349,N_19185,N_19124);
and U19350 (N_19350,N_19133,N_19155);
or U19351 (N_19351,N_19187,N_19170);
or U19352 (N_19352,N_19158,N_19195);
xor U19353 (N_19353,N_19158,N_19067);
or U19354 (N_19354,N_19051,N_19177);
nor U19355 (N_19355,N_19181,N_19103);
nand U19356 (N_19356,N_19077,N_19118);
xor U19357 (N_19357,N_19080,N_19082);
and U19358 (N_19358,N_19125,N_19139);
or U19359 (N_19359,N_19157,N_19084);
nand U19360 (N_19360,N_19290,N_19272);
or U19361 (N_19361,N_19234,N_19304);
or U19362 (N_19362,N_19230,N_19232);
nor U19363 (N_19363,N_19204,N_19352);
nor U19364 (N_19364,N_19329,N_19240);
or U19365 (N_19365,N_19346,N_19217);
nor U19366 (N_19366,N_19300,N_19246);
xor U19367 (N_19367,N_19330,N_19296);
and U19368 (N_19368,N_19212,N_19309);
or U19369 (N_19369,N_19323,N_19356);
or U19370 (N_19370,N_19209,N_19202);
nor U19371 (N_19371,N_19292,N_19299);
xnor U19372 (N_19372,N_19201,N_19318);
nand U19373 (N_19373,N_19287,N_19255);
and U19374 (N_19374,N_19314,N_19275);
or U19375 (N_19375,N_19313,N_19263);
or U19376 (N_19376,N_19259,N_19281);
nor U19377 (N_19377,N_19359,N_19260);
nand U19378 (N_19378,N_19220,N_19307);
nand U19379 (N_19379,N_19301,N_19328);
or U19380 (N_19380,N_19336,N_19271);
xnor U19381 (N_19381,N_19327,N_19315);
nand U19382 (N_19382,N_19231,N_19208);
xnor U19383 (N_19383,N_19284,N_19344);
and U19384 (N_19384,N_19306,N_19278);
nand U19385 (N_19385,N_19256,N_19215);
xor U19386 (N_19386,N_19253,N_19289);
xnor U19387 (N_19387,N_19266,N_19236);
or U19388 (N_19388,N_19302,N_19250);
nor U19389 (N_19389,N_19214,N_19228);
xor U19390 (N_19390,N_19241,N_19316);
nand U19391 (N_19391,N_19244,N_19280);
or U19392 (N_19392,N_19324,N_19249);
and U19393 (N_19393,N_19252,N_19293);
xor U19394 (N_19394,N_19288,N_19226);
or U19395 (N_19395,N_19351,N_19229);
or U19396 (N_19396,N_19340,N_19218);
nor U19397 (N_19397,N_19305,N_19235);
xor U19398 (N_19398,N_19213,N_19274);
and U19399 (N_19399,N_19206,N_19276);
xnor U19400 (N_19400,N_19261,N_19343);
nand U19401 (N_19401,N_19283,N_19279);
nor U19402 (N_19402,N_19342,N_19354);
xnor U19403 (N_19403,N_19298,N_19303);
or U19404 (N_19404,N_19297,N_19291);
xnor U19405 (N_19405,N_19210,N_19270);
and U19406 (N_19406,N_19257,N_19319);
and U19407 (N_19407,N_19203,N_19326);
and U19408 (N_19408,N_19321,N_19233);
and U19409 (N_19409,N_19200,N_19358);
xnor U19410 (N_19410,N_19320,N_19339);
xnor U19411 (N_19411,N_19222,N_19221);
nand U19412 (N_19412,N_19338,N_19286);
or U19413 (N_19413,N_19251,N_19245);
xnor U19414 (N_19414,N_19267,N_19294);
nand U19415 (N_19415,N_19317,N_19282);
nor U19416 (N_19416,N_19337,N_19247);
nand U19417 (N_19417,N_19262,N_19269);
or U19418 (N_19418,N_19207,N_19225);
xnor U19419 (N_19419,N_19341,N_19322);
and U19420 (N_19420,N_19308,N_19285);
and U19421 (N_19421,N_19205,N_19237);
or U19422 (N_19422,N_19277,N_19312);
or U19423 (N_19423,N_19227,N_19254);
nand U19424 (N_19424,N_19310,N_19349);
or U19425 (N_19425,N_19355,N_19347);
and U19426 (N_19426,N_19243,N_19265);
nor U19427 (N_19427,N_19264,N_19334);
or U19428 (N_19428,N_19348,N_19219);
nand U19429 (N_19429,N_19242,N_19332);
nor U19430 (N_19430,N_19357,N_19350);
and U19431 (N_19431,N_19353,N_19335);
nand U19432 (N_19432,N_19331,N_19223);
or U19433 (N_19433,N_19211,N_19311);
or U19434 (N_19434,N_19258,N_19224);
nand U19435 (N_19435,N_19216,N_19333);
nand U19436 (N_19436,N_19295,N_19268);
and U19437 (N_19437,N_19345,N_19273);
and U19438 (N_19438,N_19239,N_19325);
and U19439 (N_19439,N_19248,N_19238);
or U19440 (N_19440,N_19250,N_19347);
and U19441 (N_19441,N_19211,N_19356);
nand U19442 (N_19442,N_19215,N_19337);
xor U19443 (N_19443,N_19224,N_19298);
or U19444 (N_19444,N_19272,N_19245);
nand U19445 (N_19445,N_19282,N_19268);
or U19446 (N_19446,N_19358,N_19334);
or U19447 (N_19447,N_19334,N_19301);
nand U19448 (N_19448,N_19355,N_19310);
nor U19449 (N_19449,N_19230,N_19346);
or U19450 (N_19450,N_19205,N_19332);
xor U19451 (N_19451,N_19211,N_19287);
or U19452 (N_19452,N_19201,N_19346);
xor U19453 (N_19453,N_19279,N_19294);
nand U19454 (N_19454,N_19238,N_19324);
nor U19455 (N_19455,N_19265,N_19305);
or U19456 (N_19456,N_19287,N_19343);
or U19457 (N_19457,N_19205,N_19259);
or U19458 (N_19458,N_19336,N_19293);
nand U19459 (N_19459,N_19230,N_19338);
nand U19460 (N_19460,N_19278,N_19297);
xnor U19461 (N_19461,N_19202,N_19318);
nand U19462 (N_19462,N_19223,N_19317);
nor U19463 (N_19463,N_19342,N_19220);
or U19464 (N_19464,N_19345,N_19322);
or U19465 (N_19465,N_19306,N_19300);
nand U19466 (N_19466,N_19348,N_19246);
or U19467 (N_19467,N_19204,N_19215);
and U19468 (N_19468,N_19293,N_19341);
xnor U19469 (N_19469,N_19356,N_19349);
nand U19470 (N_19470,N_19345,N_19258);
xor U19471 (N_19471,N_19256,N_19252);
or U19472 (N_19472,N_19240,N_19334);
and U19473 (N_19473,N_19337,N_19320);
xor U19474 (N_19474,N_19261,N_19331);
and U19475 (N_19475,N_19324,N_19230);
nand U19476 (N_19476,N_19209,N_19223);
nand U19477 (N_19477,N_19219,N_19248);
or U19478 (N_19478,N_19217,N_19260);
and U19479 (N_19479,N_19284,N_19240);
and U19480 (N_19480,N_19264,N_19261);
or U19481 (N_19481,N_19239,N_19216);
xor U19482 (N_19482,N_19215,N_19276);
xor U19483 (N_19483,N_19328,N_19302);
nand U19484 (N_19484,N_19260,N_19303);
or U19485 (N_19485,N_19269,N_19299);
nor U19486 (N_19486,N_19284,N_19225);
nor U19487 (N_19487,N_19336,N_19255);
or U19488 (N_19488,N_19346,N_19274);
xor U19489 (N_19489,N_19305,N_19245);
nor U19490 (N_19490,N_19335,N_19336);
and U19491 (N_19491,N_19335,N_19300);
nor U19492 (N_19492,N_19267,N_19236);
nor U19493 (N_19493,N_19213,N_19201);
or U19494 (N_19494,N_19346,N_19275);
and U19495 (N_19495,N_19246,N_19229);
and U19496 (N_19496,N_19262,N_19357);
nand U19497 (N_19497,N_19275,N_19253);
or U19498 (N_19498,N_19213,N_19244);
and U19499 (N_19499,N_19208,N_19268);
nor U19500 (N_19500,N_19352,N_19209);
nor U19501 (N_19501,N_19273,N_19356);
xor U19502 (N_19502,N_19275,N_19264);
xor U19503 (N_19503,N_19325,N_19326);
and U19504 (N_19504,N_19283,N_19216);
or U19505 (N_19505,N_19261,N_19355);
xor U19506 (N_19506,N_19290,N_19238);
nand U19507 (N_19507,N_19215,N_19354);
nand U19508 (N_19508,N_19255,N_19241);
nand U19509 (N_19509,N_19335,N_19355);
and U19510 (N_19510,N_19284,N_19305);
xor U19511 (N_19511,N_19262,N_19246);
or U19512 (N_19512,N_19333,N_19222);
or U19513 (N_19513,N_19310,N_19339);
xnor U19514 (N_19514,N_19253,N_19323);
nand U19515 (N_19515,N_19355,N_19215);
nor U19516 (N_19516,N_19249,N_19358);
nand U19517 (N_19517,N_19298,N_19215);
nand U19518 (N_19518,N_19281,N_19246);
or U19519 (N_19519,N_19320,N_19231);
and U19520 (N_19520,N_19418,N_19476);
and U19521 (N_19521,N_19485,N_19513);
nand U19522 (N_19522,N_19398,N_19475);
xnor U19523 (N_19523,N_19480,N_19396);
xnor U19524 (N_19524,N_19364,N_19362);
nor U19525 (N_19525,N_19507,N_19372);
nand U19526 (N_19526,N_19450,N_19386);
nand U19527 (N_19527,N_19518,N_19394);
xnor U19528 (N_19528,N_19406,N_19432);
nand U19529 (N_19529,N_19483,N_19460);
nor U19530 (N_19530,N_19429,N_19481);
nand U19531 (N_19531,N_19435,N_19446);
or U19532 (N_19532,N_19445,N_19452);
nor U19533 (N_19533,N_19436,N_19447);
xnor U19534 (N_19534,N_19457,N_19409);
or U19535 (N_19535,N_19421,N_19495);
or U19536 (N_19536,N_19401,N_19374);
and U19537 (N_19537,N_19441,N_19405);
nor U19538 (N_19538,N_19387,N_19408);
xor U19539 (N_19539,N_19430,N_19390);
nand U19540 (N_19540,N_19515,N_19517);
nor U19541 (N_19541,N_19461,N_19464);
and U19542 (N_19542,N_19369,N_19376);
nand U19543 (N_19543,N_19428,N_19504);
nand U19544 (N_19544,N_19455,N_19443);
or U19545 (N_19545,N_19462,N_19425);
xnor U19546 (N_19546,N_19360,N_19392);
and U19547 (N_19547,N_19484,N_19471);
nor U19548 (N_19548,N_19442,N_19380);
xnor U19549 (N_19549,N_19426,N_19415);
nor U19550 (N_19550,N_19466,N_19377);
nor U19551 (N_19551,N_19417,N_19459);
xnor U19552 (N_19552,N_19371,N_19375);
and U19553 (N_19553,N_19497,N_19411);
and U19554 (N_19554,N_19416,N_19368);
and U19555 (N_19555,N_19395,N_19506);
or U19556 (N_19556,N_19391,N_19410);
nor U19557 (N_19557,N_19420,N_19512);
or U19558 (N_19558,N_19399,N_19519);
nor U19559 (N_19559,N_19487,N_19486);
nor U19560 (N_19560,N_19403,N_19448);
nand U19561 (N_19561,N_19470,N_19427);
or U19562 (N_19562,N_19503,N_19492);
and U19563 (N_19563,N_19488,N_19516);
xnor U19564 (N_19564,N_19373,N_19490);
nand U19565 (N_19565,N_19367,N_19393);
xor U19566 (N_19566,N_19453,N_19501);
nand U19567 (N_19567,N_19511,N_19477);
nand U19568 (N_19568,N_19438,N_19465);
xor U19569 (N_19569,N_19440,N_19456);
and U19570 (N_19570,N_19413,N_19510);
or U19571 (N_19571,N_19400,N_19444);
xor U19572 (N_19572,N_19467,N_19412);
nand U19573 (N_19573,N_19383,N_19463);
nor U19574 (N_19574,N_19451,N_19378);
nor U19575 (N_19575,N_19505,N_19433);
xnor U19576 (N_19576,N_19449,N_19502);
or U19577 (N_19577,N_19489,N_19434);
nor U19578 (N_19578,N_19402,N_19422);
nand U19579 (N_19579,N_19424,N_19498);
or U19580 (N_19580,N_19404,N_19474);
nor U19581 (N_19581,N_19397,N_19509);
or U19582 (N_19582,N_19473,N_19500);
nand U19583 (N_19583,N_19479,N_19496);
nor U19584 (N_19584,N_19365,N_19366);
nor U19585 (N_19585,N_19458,N_19494);
xor U19586 (N_19586,N_19472,N_19363);
nand U19587 (N_19587,N_19407,N_19454);
xnor U19588 (N_19588,N_19439,N_19468);
and U19589 (N_19589,N_19381,N_19431);
nor U19590 (N_19590,N_19419,N_19423);
and U19591 (N_19591,N_19414,N_19478);
or U19592 (N_19592,N_19384,N_19514);
or U19593 (N_19593,N_19382,N_19491);
nand U19594 (N_19594,N_19493,N_19499);
and U19595 (N_19595,N_19469,N_19370);
xnor U19596 (N_19596,N_19379,N_19482);
nor U19597 (N_19597,N_19388,N_19437);
or U19598 (N_19598,N_19508,N_19361);
nand U19599 (N_19599,N_19389,N_19385);
nand U19600 (N_19600,N_19503,N_19371);
or U19601 (N_19601,N_19513,N_19413);
nand U19602 (N_19602,N_19458,N_19472);
or U19603 (N_19603,N_19516,N_19397);
xor U19604 (N_19604,N_19386,N_19473);
nand U19605 (N_19605,N_19400,N_19379);
xnor U19606 (N_19606,N_19365,N_19451);
xnor U19607 (N_19607,N_19434,N_19366);
and U19608 (N_19608,N_19434,N_19410);
nor U19609 (N_19609,N_19439,N_19458);
nand U19610 (N_19610,N_19392,N_19420);
and U19611 (N_19611,N_19462,N_19479);
xnor U19612 (N_19612,N_19373,N_19367);
nand U19613 (N_19613,N_19472,N_19454);
and U19614 (N_19614,N_19491,N_19429);
nand U19615 (N_19615,N_19456,N_19360);
xor U19616 (N_19616,N_19491,N_19388);
nand U19617 (N_19617,N_19462,N_19408);
nand U19618 (N_19618,N_19425,N_19426);
nor U19619 (N_19619,N_19511,N_19497);
nand U19620 (N_19620,N_19362,N_19448);
nand U19621 (N_19621,N_19364,N_19385);
nor U19622 (N_19622,N_19474,N_19497);
nor U19623 (N_19623,N_19489,N_19409);
xor U19624 (N_19624,N_19482,N_19400);
xnor U19625 (N_19625,N_19403,N_19434);
xor U19626 (N_19626,N_19369,N_19467);
and U19627 (N_19627,N_19444,N_19391);
and U19628 (N_19628,N_19409,N_19509);
xor U19629 (N_19629,N_19468,N_19497);
nand U19630 (N_19630,N_19453,N_19455);
xnor U19631 (N_19631,N_19449,N_19486);
or U19632 (N_19632,N_19444,N_19440);
xnor U19633 (N_19633,N_19501,N_19387);
nor U19634 (N_19634,N_19514,N_19497);
xor U19635 (N_19635,N_19458,N_19489);
xor U19636 (N_19636,N_19430,N_19451);
and U19637 (N_19637,N_19457,N_19486);
nand U19638 (N_19638,N_19369,N_19407);
nand U19639 (N_19639,N_19486,N_19418);
nor U19640 (N_19640,N_19382,N_19437);
or U19641 (N_19641,N_19503,N_19421);
and U19642 (N_19642,N_19420,N_19478);
xor U19643 (N_19643,N_19472,N_19386);
nor U19644 (N_19644,N_19447,N_19399);
or U19645 (N_19645,N_19495,N_19465);
nor U19646 (N_19646,N_19372,N_19425);
xnor U19647 (N_19647,N_19365,N_19494);
or U19648 (N_19648,N_19404,N_19435);
nand U19649 (N_19649,N_19365,N_19382);
nor U19650 (N_19650,N_19439,N_19384);
nor U19651 (N_19651,N_19388,N_19368);
or U19652 (N_19652,N_19458,N_19453);
or U19653 (N_19653,N_19470,N_19404);
nor U19654 (N_19654,N_19409,N_19435);
nor U19655 (N_19655,N_19432,N_19417);
xnor U19656 (N_19656,N_19463,N_19485);
or U19657 (N_19657,N_19371,N_19442);
or U19658 (N_19658,N_19453,N_19449);
or U19659 (N_19659,N_19389,N_19378);
nand U19660 (N_19660,N_19386,N_19431);
and U19661 (N_19661,N_19428,N_19381);
nor U19662 (N_19662,N_19501,N_19486);
and U19663 (N_19663,N_19500,N_19432);
and U19664 (N_19664,N_19474,N_19438);
or U19665 (N_19665,N_19508,N_19379);
or U19666 (N_19666,N_19514,N_19517);
nor U19667 (N_19667,N_19376,N_19487);
xor U19668 (N_19668,N_19379,N_19391);
xor U19669 (N_19669,N_19377,N_19485);
or U19670 (N_19670,N_19479,N_19484);
nand U19671 (N_19671,N_19382,N_19501);
nand U19672 (N_19672,N_19373,N_19436);
xnor U19673 (N_19673,N_19509,N_19478);
or U19674 (N_19674,N_19411,N_19473);
or U19675 (N_19675,N_19424,N_19426);
and U19676 (N_19676,N_19456,N_19487);
and U19677 (N_19677,N_19466,N_19404);
nand U19678 (N_19678,N_19367,N_19496);
xor U19679 (N_19679,N_19423,N_19363);
nor U19680 (N_19680,N_19614,N_19532);
nor U19681 (N_19681,N_19631,N_19671);
or U19682 (N_19682,N_19597,N_19591);
or U19683 (N_19683,N_19646,N_19544);
nor U19684 (N_19684,N_19590,N_19575);
nor U19685 (N_19685,N_19558,N_19662);
nand U19686 (N_19686,N_19542,N_19615);
and U19687 (N_19687,N_19521,N_19530);
nand U19688 (N_19688,N_19525,N_19579);
and U19689 (N_19689,N_19621,N_19537);
or U19690 (N_19690,N_19635,N_19653);
and U19691 (N_19691,N_19523,N_19654);
xnor U19692 (N_19692,N_19651,N_19586);
nor U19693 (N_19693,N_19632,N_19554);
nand U19694 (N_19694,N_19607,N_19677);
xnor U19695 (N_19695,N_19593,N_19650);
or U19696 (N_19696,N_19624,N_19636);
nand U19697 (N_19697,N_19678,N_19612);
nor U19698 (N_19698,N_19642,N_19600);
nand U19699 (N_19699,N_19553,N_19664);
nor U19700 (N_19700,N_19659,N_19524);
xnor U19701 (N_19701,N_19598,N_19547);
nor U19702 (N_19702,N_19626,N_19549);
nor U19703 (N_19703,N_19522,N_19675);
nor U19704 (N_19704,N_19584,N_19572);
or U19705 (N_19705,N_19603,N_19596);
or U19706 (N_19706,N_19641,N_19588);
xor U19707 (N_19707,N_19630,N_19566);
nor U19708 (N_19708,N_19567,N_19625);
xnor U19709 (N_19709,N_19585,N_19568);
or U19710 (N_19710,N_19529,N_19546);
xor U19711 (N_19711,N_19548,N_19648);
or U19712 (N_19712,N_19556,N_19602);
nor U19713 (N_19713,N_19649,N_19656);
nor U19714 (N_19714,N_19540,N_19652);
nand U19715 (N_19715,N_19643,N_19628);
or U19716 (N_19716,N_19665,N_19595);
or U19717 (N_19717,N_19616,N_19552);
nor U19718 (N_19718,N_19535,N_19557);
nor U19719 (N_19719,N_19620,N_19528);
nand U19720 (N_19720,N_19644,N_19594);
nand U19721 (N_19721,N_19543,N_19629);
and U19722 (N_19722,N_19564,N_19583);
and U19723 (N_19723,N_19527,N_19580);
nor U19724 (N_19724,N_19610,N_19673);
nor U19725 (N_19725,N_19676,N_19539);
nand U19726 (N_19726,N_19573,N_19570);
or U19727 (N_19727,N_19618,N_19633);
nand U19728 (N_19728,N_19639,N_19560);
nand U19729 (N_19729,N_19647,N_19668);
nand U19730 (N_19730,N_19599,N_19658);
xor U19731 (N_19731,N_19605,N_19619);
nor U19732 (N_19732,N_19663,N_19637);
nand U19733 (N_19733,N_19622,N_19606);
nand U19734 (N_19734,N_19582,N_19617);
xnor U19735 (N_19735,N_19550,N_19592);
and U19736 (N_19736,N_19661,N_19638);
nor U19737 (N_19737,N_19623,N_19561);
nor U19738 (N_19738,N_19551,N_19601);
or U19739 (N_19739,N_19526,N_19541);
or U19740 (N_19740,N_19577,N_19563);
or U19741 (N_19741,N_19666,N_19627);
or U19742 (N_19742,N_19645,N_19672);
nor U19743 (N_19743,N_19533,N_19657);
or U19744 (N_19744,N_19604,N_19669);
nor U19745 (N_19745,N_19609,N_19531);
nand U19746 (N_19746,N_19562,N_19536);
nor U19747 (N_19747,N_19634,N_19611);
nand U19748 (N_19748,N_19534,N_19587);
nor U19749 (N_19749,N_19655,N_19581);
nand U19750 (N_19750,N_19538,N_19640);
nand U19751 (N_19751,N_19571,N_19660);
nor U19752 (N_19752,N_19670,N_19520);
nor U19753 (N_19753,N_19667,N_19578);
nor U19754 (N_19754,N_19574,N_19555);
or U19755 (N_19755,N_19674,N_19569);
nor U19756 (N_19756,N_19589,N_19613);
or U19757 (N_19757,N_19608,N_19565);
xnor U19758 (N_19758,N_19679,N_19559);
nor U19759 (N_19759,N_19545,N_19576);
nand U19760 (N_19760,N_19669,N_19536);
nand U19761 (N_19761,N_19531,N_19639);
nor U19762 (N_19762,N_19658,N_19670);
xor U19763 (N_19763,N_19579,N_19531);
and U19764 (N_19764,N_19555,N_19575);
nor U19765 (N_19765,N_19600,N_19540);
nor U19766 (N_19766,N_19627,N_19572);
or U19767 (N_19767,N_19536,N_19635);
or U19768 (N_19768,N_19559,N_19601);
xnor U19769 (N_19769,N_19572,N_19659);
and U19770 (N_19770,N_19661,N_19635);
xor U19771 (N_19771,N_19573,N_19534);
xor U19772 (N_19772,N_19677,N_19675);
and U19773 (N_19773,N_19617,N_19612);
and U19774 (N_19774,N_19611,N_19613);
nor U19775 (N_19775,N_19528,N_19561);
and U19776 (N_19776,N_19590,N_19593);
xor U19777 (N_19777,N_19671,N_19550);
or U19778 (N_19778,N_19533,N_19597);
and U19779 (N_19779,N_19666,N_19626);
nor U19780 (N_19780,N_19530,N_19646);
nor U19781 (N_19781,N_19611,N_19601);
nand U19782 (N_19782,N_19523,N_19611);
xor U19783 (N_19783,N_19589,N_19663);
nand U19784 (N_19784,N_19616,N_19562);
and U19785 (N_19785,N_19542,N_19551);
or U19786 (N_19786,N_19564,N_19661);
and U19787 (N_19787,N_19582,N_19566);
and U19788 (N_19788,N_19530,N_19549);
nor U19789 (N_19789,N_19536,N_19660);
or U19790 (N_19790,N_19637,N_19658);
nand U19791 (N_19791,N_19619,N_19674);
nand U19792 (N_19792,N_19654,N_19602);
nor U19793 (N_19793,N_19563,N_19637);
nor U19794 (N_19794,N_19527,N_19665);
nand U19795 (N_19795,N_19580,N_19679);
nand U19796 (N_19796,N_19585,N_19668);
nand U19797 (N_19797,N_19623,N_19583);
and U19798 (N_19798,N_19548,N_19570);
and U19799 (N_19799,N_19624,N_19679);
or U19800 (N_19800,N_19521,N_19607);
or U19801 (N_19801,N_19539,N_19641);
xnor U19802 (N_19802,N_19525,N_19640);
nor U19803 (N_19803,N_19631,N_19567);
xnor U19804 (N_19804,N_19530,N_19568);
nand U19805 (N_19805,N_19610,N_19608);
xor U19806 (N_19806,N_19663,N_19639);
or U19807 (N_19807,N_19597,N_19599);
xor U19808 (N_19808,N_19587,N_19609);
nand U19809 (N_19809,N_19623,N_19619);
or U19810 (N_19810,N_19602,N_19530);
nor U19811 (N_19811,N_19541,N_19587);
nor U19812 (N_19812,N_19570,N_19533);
or U19813 (N_19813,N_19564,N_19655);
xor U19814 (N_19814,N_19595,N_19612);
and U19815 (N_19815,N_19574,N_19533);
xor U19816 (N_19816,N_19652,N_19598);
nand U19817 (N_19817,N_19543,N_19595);
or U19818 (N_19818,N_19527,N_19651);
xor U19819 (N_19819,N_19666,N_19642);
xnor U19820 (N_19820,N_19625,N_19521);
nand U19821 (N_19821,N_19605,N_19653);
or U19822 (N_19822,N_19667,N_19540);
or U19823 (N_19823,N_19531,N_19570);
nor U19824 (N_19824,N_19619,N_19560);
nand U19825 (N_19825,N_19553,N_19534);
or U19826 (N_19826,N_19631,N_19633);
nor U19827 (N_19827,N_19639,N_19538);
nor U19828 (N_19828,N_19649,N_19613);
nor U19829 (N_19829,N_19545,N_19537);
nand U19830 (N_19830,N_19601,N_19544);
and U19831 (N_19831,N_19598,N_19526);
or U19832 (N_19832,N_19671,N_19620);
and U19833 (N_19833,N_19535,N_19593);
nand U19834 (N_19834,N_19625,N_19520);
xor U19835 (N_19835,N_19562,N_19675);
nand U19836 (N_19836,N_19574,N_19543);
xnor U19837 (N_19837,N_19678,N_19530);
xnor U19838 (N_19838,N_19591,N_19666);
or U19839 (N_19839,N_19525,N_19663);
nor U19840 (N_19840,N_19750,N_19748);
nor U19841 (N_19841,N_19793,N_19766);
xor U19842 (N_19842,N_19811,N_19685);
or U19843 (N_19843,N_19779,N_19717);
and U19844 (N_19844,N_19714,N_19777);
nand U19845 (N_19845,N_19704,N_19693);
nor U19846 (N_19846,N_19770,N_19754);
nand U19847 (N_19847,N_19711,N_19795);
nand U19848 (N_19848,N_19746,N_19780);
nand U19849 (N_19849,N_19764,N_19813);
nand U19850 (N_19850,N_19701,N_19719);
xnor U19851 (N_19851,N_19775,N_19721);
xor U19852 (N_19852,N_19781,N_19707);
xnor U19853 (N_19853,N_19745,N_19822);
or U19854 (N_19854,N_19792,N_19807);
nor U19855 (N_19855,N_19725,N_19739);
xor U19856 (N_19856,N_19755,N_19819);
and U19857 (N_19857,N_19835,N_19757);
xor U19858 (N_19858,N_19839,N_19826);
or U19859 (N_19859,N_19751,N_19829);
nor U19860 (N_19860,N_19689,N_19747);
xor U19861 (N_19861,N_19809,N_19786);
nor U19862 (N_19862,N_19761,N_19697);
nand U19863 (N_19863,N_19735,N_19688);
and U19864 (N_19864,N_19728,N_19709);
and U19865 (N_19865,N_19759,N_19742);
nand U19866 (N_19866,N_19756,N_19737);
nand U19867 (N_19867,N_19708,N_19686);
nor U19868 (N_19868,N_19767,N_19713);
xnor U19869 (N_19869,N_19718,N_19799);
xnor U19870 (N_19870,N_19763,N_19836);
xnor U19871 (N_19871,N_19831,N_19692);
xor U19872 (N_19872,N_19682,N_19765);
xor U19873 (N_19873,N_19700,N_19696);
nand U19874 (N_19874,N_19726,N_19791);
xnor U19875 (N_19875,N_19771,N_19712);
or U19876 (N_19876,N_19695,N_19821);
and U19877 (N_19877,N_19825,N_19806);
and U19878 (N_19878,N_19790,N_19818);
and U19879 (N_19879,N_19834,N_19823);
and U19880 (N_19880,N_19740,N_19743);
nor U19881 (N_19881,N_19812,N_19773);
and U19882 (N_19882,N_19752,N_19758);
xnor U19883 (N_19883,N_19699,N_19706);
and U19884 (N_19884,N_19733,N_19736);
or U19885 (N_19885,N_19798,N_19817);
or U19886 (N_19886,N_19797,N_19832);
nand U19887 (N_19887,N_19808,N_19827);
or U19888 (N_19888,N_19716,N_19824);
nor U19889 (N_19889,N_19837,N_19694);
nor U19890 (N_19890,N_19690,N_19724);
and U19891 (N_19891,N_19768,N_19710);
and U19892 (N_19892,N_19816,N_19789);
xnor U19893 (N_19893,N_19731,N_19749);
and U19894 (N_19894,N_19683,N_19784);
nand U19895 (N_19895,N_19684,N_19732);
nor U19896 (N_19896,N_19800,N_19776);
nand U19897 (N_19897,N_19702,N_19687);
xor U19898 (N_19898,N_19802,N_19774);
nand U19899 (N_19899,N_19734,N_19803);
or U19900 (N_19900,N_19703,N_19722);
and U19901 (N_19901,N_19727,N_19810);
xor U19902 (N_19902,N_19794,N_19788);
nand U19903 (N_19903,N_19715,N_19796);
nand U19904 (N_19904,N_19738,N_19681);
nand U19905 (N_19905,N_19830,N_19782);
and U19906 (N_19906,N_19787,N_19691);
nor U19907 (N_19907,N_19723,N_19801);
and U19908 (N_19908,N_19762,N_19729);
nor U19909 (N_19909,N_19785,N_19778);
xnor U19910 (N_19910,N_19753,N_19741);
or U19911 (N_19911,N_19698,N_19744);
or U19912 (N_19912,N_19814,N_19838);
or U19913 (N_19913,N_19804,N_19783);
and U19914 (N_19914,N_19805,N_19833);
or U19915 (N_19915,N_19705,N_19760);
or U19916 (N_19916,N_19815,N_19730);
and U19917 (N_19917,N_19772,N_19720);
xor U19918 (N_19918,N_19820,N_19828);
nand U19919 (N_19919,N_19680,N_19769);
nor U19920 (N_19920,N_19759,N_19763);
or U19921 (N_19921,N_19739,N_19778);
and U19922 (N_19922,N_19700,N_19724);
nand U19923 (N_19923,N_19749,N_19815);
nand U19924 (N_19924,N_19781,N_19727);
nor U19925 (N_19925,N_19780,N_19806);
xor U19926 (N_19926,N_19769,N_19831);
and U19927 (N_19927,N_19782,N_19708);
and U19928 (N_19928,N_19834,N_19793);
xor U19929 (N_19929,N_19804,N_19713);
xnor U19930 (N_19930,N_19718,N_19695);
and U19931 (N_19931,N_19778,N_19697);
xor U19932 (N_19932,N_19762,N_19755);
nor U19933 (N_19933,N_19702,N_19778);
nand U19934 (N_19934,N_19745,N_19826);
nand U19935 (N_19935,N_19790,N_19784);
or U19936 (N_19936,N_19785,N_19802);
nand U19937 (N_19937,N_19693,N_19688);
xor U19938 (N_19938,N_19800,N_19825);
nor U19939 (N_19939,N_19733,N_19741);
nor U19940 (N_19940,N_19783,N_19800);
nor U19941 (N_19941,N_19731,N_19821);
nor U19942 (N_19942,N_19698,N_19696);
and U19943 (N_19943,N_19833,N_19685);
or U19944 (N_19944,N_19801,N_19797);
nand U19945 (N_19945,N_19743,N_19705);
and U19946 (N_19946,N_19754,N_19709);
nand U19947 (N_19947,N_19811,N_19792);
nand U19948 (N_19948,N_19822,N_19689);
nand U19949 (N_19949,N_19733,N_19791);
and U19950 (N_19950,N_19692,N_19700);
or U19951 (N_19951,N_19787,N_19735);
or U19952 (N_19952,N_19830,N_19767);
nand U19953 (N_19953,N_19702,N_19786);
nor U19954 (N_19954,N_19813,N_19681);
nor U19955 (N_19955,N_19698,N_19786);
and U19956 (N_19956,N_19755,N_19737);
nor U19957 (N_19957,N_19705,N_19747);
or U19958 (N_19958,N_19819,N_19827);
or U19959 (N_19959,N_19800,N_19795);
or U19960 (N_19960,N_19782,N_19831);
nor U19961 (N_19961,N_19722,N_19749);
xnor U19962 (N_19962,N_19830,N_19819);
and U19963 (N_19963,N_19813,N_19798);
nand U19964 (N_19964,N_19798,N_19693);
nor U19965 (N_19965,N_19754,N_19831);
or U19966 (N_19966,N_19782,N_19750);
and U19967 (N_19967,N_19796,N_19766);
and U19968 (N_19968,N_19686,N_19778);
nand U19969 (N_19969,N_19681,N_19833);
nor U19970 (N_19970,N_19761,N_19710);
nor U19971 (N_19971,N_19783,N_19728);
and U19972 (N_19972,N_19770,N_19720);
and U19973 (N_19973,N_19803,N_19778);
and U19974 (N_19974,N_19826,N_19796);
and U19975 (N_19975,N_19750,N_19786);
nand U19976 (N_19976,N_19687,N_19754);
or U19977 (N_19977,N_19829,N_19726);
xor U19978 (N_19978,N_19712,N_19830);
or U19979 (N_19979,N_19772,N_19753);
nor U19980 (N_19980,N_19731,N_19757);
xor U19981 (N_19981,N_19715,N_19754);
and U19982 (N_19982,N_19740,N_19715);
nand U19983 (N_19983,N_19827,N_19713);
xnor U19984 (N_19984,N_19758,N_19734);
nor U19985 (N_19985,N_19740,N_19788);
nand U19986 (N_19986,N_19725,N_19806);
or U19987 (N_19987,N_19800,N_19834);
xor U19988 (N_19988,N_19786,N_19823);
nor U19989 (N_19989,N_19695,N_19723);
xor U19990 (N_19990,N_19699,N_19835);
nand U19991 (N_19991,N_19685,N_19709);
and U19992 (N_19992,N_19728,N_19836);
xnor U19993 (N_19993,N_19767,N_19719);
nand U19994 (N_19994,N_19727,N_19784);
nand U19995 (N_19995,N_19689,N_19721);
and U19996 (N_19996,N_19774,N_19782);
or U19997 (N_19997,N_19764,N_19748);
nor U19998 (N_19998,N_19794,N_19735);
nor U19999 (N_19999,N_19819,N_19722);
or UO_0 (O_0,N_19898,N_19858);
nor UO_1 (O_1,N_19933,N_19991);
or UO_2 (O_2,N_19856,N_19997);
nand UO_3 (O_3,N_19896,N_19921);
or UO_4 (O_4,N_19956,N_19873);
nand UO_5 (O_5,N_19930,N_19941);
nand UO_6 (O_6,N_19995,N_19934);
nor UO_7 (O_7,N_19889,N_19977);
xor UO_8 (O_8,N_19984,N_19970);
or UO_9 (O_9,N_19845,N_19998);
nand UO_10 (O_10,N_19892,N_19869);
or UO_11 (O_11,N_19911,N_19925);
nand UO_12 (O_12,N_19861,N_19910);
xor UO_13 (O_13,N_19986,N_19992);
or UO_14 (O_14,N_19978,N_19987);
xnor UO_15 (O_15,N_19915,N_19870);
or UO_16 (O_16,N_19893,N_19851);
nor UO_17 (O_17,N_19854,N_19928);
nor UO_18 (O_18,N_19864,N_19878);
or UO_19 (O_19,N_19907,N_19939);
nor UO_20 (O_20,N_19981,N_19899);
xor UO_21 (O_21,N_19968,N_19953);
or UO_22 (O_22,N_19875,N_19926);
or UO_23 (O_23,N_19975,N_19983);
or UO_24 (O_24,N_19848,N_19883);
or UO_25 (O_25,N_19877,N_19863);
or UO_26 (O_26,N_19843,N_19890);
nor UO_27 (O_27,N_19901,N_19924);
nor UO_28 (O_28,N_19958,N_19887);
or UO_29 (O_29,N_19846,N_19857);
xnor UO_30 (O_30,N_19865,N_19912);
nor UO_31 (O_31,N_19982,N_19868);
xnor UO_32 (O_32,N_19881,N_19882);
nor UO_33 (O_33,N_19951,N_19944);
nand UO_34 (O_34,N_19913,N_19917);
or UO_35 (O_35,N_19876,N_19867);
and UO_36 (O_36,N_19996,N_19872);
and UO_37 (O_37,N_19849,N_19965);
nand UO_38 (O_38,N_19855,N_19866);
nand UO_39 (O_39,N_19966,N_19943);
nand UO_40 (O_40,N_19922,N_19879);
and UO_41 (O_41,N_19841,N_19960);
or UO_42 (O_42,N_19957,N_19874);
or UO_43 (O_43,N_19905,N_19999);
or UO_44 (O_44,N_19903,N_19959);
and UO_45 (O_45,N_19871,N_19971);
and UO_46 (O_46,N_19918,N_19885);
or UO_47 (O_47,N_19988,N_19847);
and UO_48 (O_48,N_19840,N_19976);
nand UO_49 (O_49,N_19969,N_19947);
nand UO_50 (O_50,N_19859,N_19949);
or UO_51 (O_51,N_19842,N_19929);
nor UO_52 (O_52,N_19946,N_19989);
and UO_53 (O_53,N_19963,N_19894);
nand UO_54 (O_54,N_19850,N_19914);
nand UO_55 (O_55,N_19994,N_19916);
and UO_56 (O_56,N_19906,N_19937);
nand UO_57 (O_57,N_19897,N_19886);
or UO_58 (O_58,N_19952,N_19932);
nand UO_59 (O_59,N_19974,N_19940);
xor UO_60 (O_60,N_19936,N_19927);
and UO_61 (O_61,N_19923,N_19852);
and UO_62 (O_62,N_19950,N_19985);
nand UO_63 (O_63,N_19967,N_19979);
xor UO_64 (O_64,N_19860,N_19884);
and UO_65 (O_65,N_19908,N_19909);
xor UO_66 (O_66,N_19990,N_19945);
xor UO_67 (O_67,N_19902,N_19980);
nor UO_68 (O_68,N_19938,N_19972);
nor UO_69 (O_69,N_19862,N_19891);
and UO_70 (O_70,N_19973,N_19853);
xor UO_71 (O_71,N_19919,N_19920);
or UO_72 (O_72,N_19964,N_19993);
and UO_73 (O_73,N_19954,N_19888);
nor UO_74 (O_74,N_19935,N_19962);
nor UO_75 (O_75,N_19961,N_19955);
or UO_76 (O_76,N_19844,N_19948);
or UO_77 (O_77,N_19895,N_19900);
nand UO_78 (O_78,N_19931,N_19942);
and UO_79 (O_79,N_19880,N_19904);
nor UO_80 (O_80,N_19893,N_19917);
or UO_81 (O_81,N_19969,N_19842);
and UO_82 (O_82,N_19908,N_19858);
nor UO_83 (O_83,N_19952,N_19844);
nor UO_84 (O_84,N_19993,N_19927);
nand UO_85 (O_85,N_19899,N_19880);
nor UO_86 (O_86,N_19954,N_19972);
xor UO_87 (O_87,N_19994,N_19868);
xnor UO_88 (O_88,N_19960,N_19996);
or UO_89 (O_89,N_19847,N_19931);
xnor UO_90 (O_90,N_19860,N_19873);
nor UO_91 (O_91,N_19862,N_19928);
nand UO_92 (O_92,N_19840,N_19843);
nor UO_93 (O_93,N_19842,N_19874);
nand UO_94 (O_94,N_19908,N_19889);
and UO_95 (O_95,N_19878,N_19940);
xnor UO_96 (O_96,N_19887,N_19869);
or UO_97 (O_97,N_19844,N_19961);
xor UO_98 (O_98,N_19910,N_19974);
xor UO_99 (O_99,N_19867,N_19920);
or UO_100 (O_100,N_19869,N_19955);
or UO_101 (O_101,N_19994,N_19906);
nor UO_102 (O_102,N_19999,N_19982);
or UO_103 (O_103,N_19967,N_19917);
and UO_104 (O_104,N_19867,N_19840);
or UO_105 (O_105,N_19921,N_19949);
nand UO_106 (O_106,N_19872,N_19850);
and UO_107 (O_107,N_19904,N_19868);
nand UO_108 (O_108,N_19874,N_19920);
nand UO_109 (O_109,N_19907,N_19952);
and UO_110 (O_110,N_19873,N_19888);
or UO_111 (O_111,N_19842,N_19868);
nor UO_112 (O_112,N_19954,N_19846);
xnor UO_113 (O_113,N_19947,N_19920);
and UO_114 (O_114,N_19949,N_19883);
nand UO_115 (O_115,N_19992,N_19980);
and UO_116 (O_116,N_19886,N_19909);
and UO_117 (O_117,N_19905,N_19943);
nand UO_118 (O_118,N_19971,N_19917);
xnor UO_119 (O_119,N_19842,N_19962);
nand UO_120 (O_120,N_19919,N_19933);
and UO_121 (O_121,N_19874,N_19866);
nor UO_122 (O_122,N_19865,N_19991);
or UO_123 (O_123,N_19986,N_19841);
and UO_124 (O_124,N_19894,N_19881);
or UO_125 (O_125,N_19893,N_19929);
and UO_126 (O_126,N_19960,N_19981);
nor UO_127 (O_127,N_19879,N_19850);
or UO_128 (O_128,N_19927,N_19866);
and UO_129 (O_129,N_19916,N_19925);
or UO_130 (O_130,N_19969,N_19844);
nor UO_131 (O_131,N_19963,N_19920);
xnor UO_132 (O_132,N_19933,N_19882);
nand UO_133 (O_133,N_19911,N_19922);
xnor UO_134 (O_134,N_19868,N_19961);
nand UO_135 (O_135,N_19977,N_19873);
nand UO_136 (O_136,N_19929,N_19974);
or UO_137 (O_137,N_19915,N_19978);
or UO_138 (O_138,N_19881,N_19945);
and UO_139 (O_139,N_19871,N_19845);
and UO_140 (O_140,N_19845,N_19940);
nand UO_141 (O_141,N_19915,N_19854);
nand UO_142 (O_142,N_19943,N_19967);
nor UO_143 (O_143,N_19888,N_19893);
nand UO_144 (O_144,N_19986,N_19922);
nand UO_145 (O_145,N_19875,N_19932);
xnor UO_146 (O_146,N_19873,N_19908);
and UO_147 (O_147,N_19908,N_19864);
nor UO_148 (O_148,N_19949,N_19869);
nand UO_149 (O_149,N_19853,N_19870);
xor UO_150 (O_150,N_19875,N_19927);
and UO_151 (O_151,N_19936,N_19903);
nand UO_152 (O_152,N_19929,N_19972);
xnor UO_153 (O_153,N_19951,N_19972);
xnor UO_154 (O_154,N_19890,N_19950);
xor UO_155 (O_155,N_19955,N_19903);
and UO_156 (O_156,N_19993,N_19941);
nor UO_157 (O_157,N_19911,N_19878);
nand UO_158 (O_158,N_19849,N_19969);
xnor UO_159 (O_159,N_19885,N_19860);
or UO_160 (O_160,N_19855,N_19967);
nor UO_161 (O_161,N_19871,N_19937);
xnor UO_162 (O_162,N_19853,N_19946);
xor UO_163 (O_163,N_19917,N_19875);
or UO_164 (O_164,N_19999,N_19978);
xor UO_165 (O_165,N_19919,N_19967);
and UO_166 (O_166,N_19992,N_19889);
and UO_167 (O_167,N_19890,N_19944);
or UO_168 (O_168,N_19912,N_19872);
and UO_169 (O_169,N_19919,N_19842);
xor UO_170 (O_170,N_19971,N_19965);
nor UO_171 (O_171,N_19934,N_19998);
nand UO_172 (O_172,N_19968,N_19947);
nor UO_173 (O_173,N_19980,N_19947);
nor UO_174 (O_174,N_19924,N_19932);
xnor UO_175 (O_175,N_19940,N_19897);
nor UO_176 (O_176,N_19939,N_19840);
nor UO_177 (O_177,N_19899,N_19885);
or UO_178 (O_178,N_19851,N_19899);
nor UO_179 (O_179,N_19860,N_19960);
and UO_180 (O_180,N_19910,N_19891);
and UO_181 (O_181,N_19963,N_19951);
xor UO_182 (O_182,N_19989,N_19982);
or UO_183 (O_183,N_19939,N_19956);
nor UO_184 (O_184,N_19851,N_19901);
and UO_185 (O_185,N_19994,N_19984);
and UO_186 (O_186,N_19931,N_19991);
nand UO_187 (O_187,N_19996,N_19998);
or UO_188 (O_188,N_19863,N_19924);
xnor UO_189 (O_189,N_19857,N_19995);
xor UO_190 (O_190,N_19953,N_19969);
and UO_191 (O_191,N_19998,N_19863);
or UO_192 (O_192,N_19872,N_19968);
nand UO_193 (O_193,N_19863,N_19906);
nand UO_194 (O_194,N_19969,N_19914);
xnor UO_195 (O_195,N_19988,N_19970);
nand UO_196 (O_196,N_19922,N_19972);
and UO_197 (O_197,N_19889,N_19938);
or UO_198 (O_198,N_19983,N_19960);
or UO_199 (O_199,N_19938,N_19944);
nor UO_200 (O_200,N_19903,N_19875);
nand UO_201 (O_201,N_19953,N_19893);
and UO_202 (O_202,N_19920,N_19899);
nor UO_203 (O_203,N_19875,N_19935);
nor UO_204 (O_204,N_19961,N_19954);
nand UO_205 (O_205,N_19940,N_19976);
and UO_206 (O_206,N_19918,N_19921);
and UO_207 (O_207,N_19948,N_19912);
nor UO_208 (O_208,N_19987,N_19845);
nand UO_209 (O_209,N_19887,N_19976);
and UO_210 (O_210,N_19865,N_19849);
nor UO_211 (O_211,N_19846,N_19913);
and UO_212 (O_212,N_19896,N_19841);
nor UO_213 (O_213,N_19939,N_19859);
nand UO_214 (O_214,N_19935,N_19958);
and UO_215 (O_215,N_19863,N_19981);
or UO_216 (O_216,N_19926,N_19870);
nand UO_217 (O_217,N_19872,N_19974);
nor UO_218 (O_218,N_19950,N_19895);
nand UO_219 (O_219,N_19990,N_19991);
xnor UO_220 (O_220,N_19906,N_19923);
or UO_221 (O_221,N_19988,N_19945);
nand UO_222 (O_222,N_19845,N_19877);
and UO_223 (O_223,N_19866,N_19983);
and UO_224 (O_224,N_19902,N_19883);
nor UO_225 (O_225,N_19973,N_19891);
and UO_226 (O_226,N_19957,N_19941);
nor UO_227 (O_227,N_19934,N_19900);
nand UO_228 (O_228,N_19875,N_19978);
xnor UO_229 (O_229,N_19956,N_19920);
and UO_230 (O_230,N_19971,N_19905);
and UO_231 (O_231,N_19903,N_19873);
or UO_232 (O_232,N_19867,N_19945);
nor UO_233 (O_233,N_19898,N_19935);
or UO_234 (O_234,N_19861,N_19919);
or UO_235 (O_235,N_19902,N_19932);
and UO_236 (O_236,N_19885,N_19962);
or UO_237 (O_237,N_19918,N_19954);
xnor UO_238 (O_238,N_19906,N_19943);
and UO_239 (O_239,N_19884,N_19843);
nor UO_240 (O_240,N_19945,N_19951);
nand UO_241 (O_241,N_19909,N_19849);
xor UO_242 (O_242,N_19909,N_19853);
nand UO_243 (O_243,N_19865,N_19969);
xnor UO_244 (O_244,N_19941,N_19948);
xor UO_245 (O_245,N_19964,N_19999);
nand UO_246 (O_246,N_19857,N_19961);
or UO_247 (O_247,N_19983,N_19871);
xor UO_248 (O_248,N_19944,N_19918);
nor UO_249 (O_249,N_19905,N_19844);
nand UO_250 (O_250,N_19951,N_19900);
nor UO_251 (O_251,N_19992,N_19982);
nand UO_252 (O_252,N_19947,N_19938);
or UO_253 (O_253,N_19995,N_19872);
nand UO_254 (O_254,N_19954,N_19903);
and UO_255 (O_255,N_19914,N_19892);
and UO_256 (O_256,N_19920,N_19954);
nand UO_257 (O_257,N_19962,N_19848);
and UO_258 (O_258,N_19844,N_19916);
xnor UO_259 (O_259,N_19975,N_19931);
nand UO_260 (O_260,N_19840,N_19988);
nor UO_261 (O_261,N_19863,N_19932);
or UO_262 (O_262,N_19933,N_19950);
and UO_263 (O_263,N_19917,N_19970);
xor UO_264 (O_264,N_19941,N_19911);
nor UO_265 (O_265,N_19998,N_19974);
and UO_266 (O_266,N_19912,N_19968);
or UO_267 (O_267,N_19953,N_19882);
and UO_268 (O_268,N_19998,N_19997);
and UO_269 (O_269,N_19870,N_19967);
nand UO_270 (O_270,N_19883,N_19913);
nand UO_271 (O_271,N_19928,N_19840);
or UO_272 (O_272,N_19855,N_19917);
or UO_273 (O_273,N_19872,N_19921);
nand UO_274 (O_274,N_19963,N_19944);
nor UO_275 (O_275,N_19859,N_19973);
or UO_276 (O_276,N_19981,N_19933);
and UO_277 (O_277,N_19865,N_19896);
nor UO_278 (O_278,N_19955,N_19984);
or UO_279 (O_279,N_19887,N_19860);
xor UO_280 (O_280,N_19848,N_19872);
nor UO_281 (O_281,N_19927,N_19899);
and UO_282 (O_282,N_19883,N_19937);
or UO_283 (O_283,N_19934,N_19950);
or UO_284 (O_284,N_19979,N_19932);
and UO_285 (O_285,N_19870,N_19860);
nor UO_286 (O_286,N_19866,N_19957);
xnor UO_287 (O_287,N_19977,N_19996);
nor UO_288 (O_288,N_19988,N_19898);
or UO_289 (O_289,N_19906,N_19944);
nor UO_290 (O_290,N_19880,N_19874);
nand UO_291 (O_291,N_19875,N_19915);
and UO_292 (O_292,N_19984,N_19918);
nand UO_293 (O_293,N_19961,N_19878);
and UO_294 (O_294,N_19989,N_19841);
xor UO_295 (O_295,N_19908,N_19884);
and UO_296 (O_296,N_19902,N_19943);
and UO_297 (O_297,N_19864,N_19934);
nand UO_298 (O_298,N_19956,N_19885);
nand UO_299 (O_299,N_19961,N_19881);
nand UO_300 (O_300,N_19887,N_19882);
nor UO_301 (O_301,N_19863,N_19875);
nor UO_302 (O_302,N_19895,N_19946);
xnor UO_303 (O_303,N_19907,N_19927);
and UO_304 (O_304,N_19934,N_19962);
or UO_305 (O_305,N_19891,N_19960);
nor UO_306 (O_306,N_19912,N_19890);
nand UO_307 (O_307,N_19970,N_19861);
and UO_308 (O_308,N_19886,N_19915);
xnor UO_309 (O_309,N_19849,N_19973);
xor UO_310 (O_310,N_19990,N_19901);
and UO_311 (O_311,N_19853,N_19875);
and UO_312 (O_312,N_19960,N_19843);
nor UO_313 (O_313,N_19957,N_19891);
nand UO_314 (O_314,N_19894,N_19854);
or UO_315 (O_315,N_19855,N_19972);
nand UO_316 (O_316,N_19935,N_19873);
or UO_317 (O_317,N_19967,N_19964);
nor UO_318 (O_318,N_19963,N_19913);
or UO_319 (O_319,N_19860,N_19965);
nor UO_320 (O_320,N_19905,N_19920);
and UO_321 (O_321,N_19845,N_19900);
or UO_322 (O_322,N_19940,N_19852);
or UO_323 (O_323,N_19998,N_19890);
nand UO_324 (O_324,N_19893,N_19879);
nor UO_325 (O_325,N_19924,N_19951);
nor UO_326 (O_326,N_19868,N_19978);
or UO_327 (O_327,N_19999,N_19957);
nor UO_328 (O_328,N_19866,N_19926);
nand UO_329 (O_329,N_19982,N_19936);
nand UO_330 (O_330,N_19963,N_19880);
nand UO_331 (O_331,N_19931,N_19840);
and UO_332 (O_332,N_19960,N_19938);
nand UO_333 (O_333,N_19890,N_19898);
nor UO_334 (O_334,N_19870,N_19871);
nand UO_335 (O_335,N_19967,N_19952);
nand UO_336 (O_336,N_19880,N_19863);
nor UO_337 (O_337,N_19926,N_19967);
and UO_338 (O_338,N_19862,N_19961);
nand UO_339 (O_339,N_19895,N_19998);
and UO_340 (O_340,N_19962,N_19920);
xor UO_341 (O_341,N_19936,N_19852);
and UO_342 (O_342,N_19904,N_19978);
and UO_343 (O_343,N_19860,N_19973);
and UO_344 (O_344,N_19895,N_19993);
and UO_345 (O_345,N_19998,N_19916);
or UO_346 (O_346,N_19994,N_19877);
nand UO_347 (O_347,N_19843,N_19900);
xnor UO_348 (O_348,N_19917,N_19999);
xor UO_349 (O_349,N_19995,N_19899);
nand UO_350 (O_350,N_19988,N_19924);
and UO_351 (O_351,N_19901,N_19928);
xnor UO_352 (O_352,N_19980,N_19948);
and UO_353 (O_353,N_19938,N_19941);
nand UO_354 (O_354,N_19847,N_19888);
xor UO_355 (O_355,N_19997,N_19859);
nand UO_356 (O_356,N_19979,N_19955);
or UO_357 (O_357,N_19899,N_19844);
nand UO_358 (O_358,N_19885,N_19928);
nand UO_359 (O_359,N_19955,N_19998);
xnor UO_360 (O_360,N_19853,N_19989);
or UO_361 (O_361,N_19911,N_19853);
or UO_362 (O_362,N_19977,N_19975);
nor UO_363 (O_363,N_19871,N_19880);
and UO_364 (O_364,N_19916,N_19930);
and UO_365 (O_365,N_19984,N_19894);
xnor UO_366 (O_366,N_19981,N_19995);
nor UO_367 (O_367,N_19897,N_19978);
and UO_368 (O_368,N_19878,N_19919);
nor UO_369 (O_369,N_19852,N_19943);
and UO_370 (O_370,N_19970,N_19933);
nand UO_371 (O_371,N_19880,N_19910);
xor UO_372 (O_372,N_19890,N_19976);
and UO_373 (O_373,N_19843,N_19877);
or UO_374 (O_374,N_19850,N_19989);
xor UO_375 (O_375,N_19913,N_19840);
xor UO_376 (O_376,N_19897,N_19980);
nor UO_377 (O_377,N_19949,N_19918);
and UO_378 (O_378,N_19897,N_19859);
nor UO_379 (O_379,N_19974,N_19905);
nor UO_380 (O_380,N_19938,N_19986);
nand UO_381 (O_381,N_19921,N_19868);
xor UO_382 (O_382,N_19995,N_19844);
xnor UO_383 (O_383,N_19911,N_19936);
or UO_384 (O_384,N_19960,N_19965);
and UO_385 (O_385,N_19900,N_19857);
and UO_386 (O_386,N_19968,N_19985);
nor UO_387 (O_387,N_19844,N_19992);
nand UO_388 (O_388,N_19986,N_19963);
or UO_389 (O_389,N_19987,N_19924);
nor UO_390 (O_390,N_19941,N_19900);
and UO_391 (O_391,N_19861,N_19929);
and UO_392 (O_392,N_19884,N_19941);
nand UO_393 (O_393,N_19883,N_19886);
nor UO_394 (O_394,N_19985,N_19924);
nor UO_395 (O_395,N_19976,N_19853);
xnor UO_396 (O_396,N_19970,N_19925);
nor UO_397 (O_397,N_19903,N_19979);
nor UO_398 (O_398,N_19928,N_19984);
xnor UO_399 (O_399,N_19840,N_19903);
xor UO_400 (O_400,N_19954,N_19842);
and UO_401 (O_401,N_19961,N_19971);
xor UO_402 (O_402,N_19930,N_19879);
or UO_403 (O_403,N_19915,N_19872);
or UO_404 (O_404,N_19986,N_19991);
and UO_405 (O_405,N_19914,N_19861);
and UO_406 (O_406,N_19887,N_19926);
or UO_407 (O_407,N_19979,N_19976);
or UO_408 (O_408,N_19990,N_19976);
nor UO_409 (O_409,N_19930,N_19843);
and UO_410 (O_410,N_19902,N_19857);
and UO_411 (O_411,N_19961,N_19879);
nand UO_412 (O_412,N_19928,N_19980);
and UO_413 (O_413,N_19917,N_19883);
nor UO_414 (O_414,N_19918,N_19935);
and UO_415 (O_415,N_19910,N_19926);
nor UO_416 (O_416,N_19934,N_19957);
and UO_417 (O_417,N_19946,N_19840);
nand UO_418 (O_418,N_19871,N_19942);
nand UO_419 (O_419,N_19974,N_19964);
nand UO_420 (O_420,N_19993,N_19912);
nor UO_421 (O_421,N_19918,N_19870);
and UO_422 (O_422,N_19906,N_19875);
and UO_423 (O_423,N_19946,N_19849);
and UO_424 (O_424,N_19916,N_19890);
and UO_425 (O_425,N_19966,N_19956);
and UO_426 (O_426,N_19876,N_19848);
nor UO_427 (O_427,N_19948,N_19944);
xor UO_428 (O_428,N_19882,N_19998);
nand UO_429 (O_429,N_19944,N_19846);
or UO_430 (O_430,N_19980,N_19841);
nand UO_431 (O_431,N_19955,N_19856);
or UO_432 (O_432,N_19872,N_19933);
and UO_433 (O_433,N_19845,N_19985);
or UO_434 (O_434,N_19912,N_19995);
and UO_435 (O_435,N_19945,N_19893);
and UO_436 (O_436,N_19843,N_19893);
nand UO_437 (O_437,N_19918,N_19952);
nor UO_438 (O_438,N_19910,N_19950);
nor UO_439 (O_439,N_19983,N_19874);
and UO_440 (O_440,N_19845,N_19926);
nor UO_441 (O_441,N_19877,N_19921);
xor UO_442 (O_442,N_19958,N_19864);
xnor UO_443 (O_443,N_19935,N_19998);
and UO_444 (O_444,N_19845,N_19993);
xnor UO_445 (O_445,N_19932,N_19994);
or UO_446 (O_446,N_19929,N_19986);
nor UO_447 (O_447,N_19978,N_19935);
nor UO_448 (O_448,N_19928,N_19859);
nor UO_449 (O_449,N_19917,N_19870);
xnor UO_450 (O_450,N_19952,N_19988);
xor UO_451 (O_451,N_19889,N_19990);
nor UO_452 (O_452,N_19942,N_19916);
nand UO_453 (O_453,N_19913,N_19931);
or UO_454 (O_454,N_19955,N_19940);
nand UO_455 (O_455,N_19960,N_19963);
nor UO_456 (O_456,N_19980,N_19896);
or UO_457 (O_457,N_19911,N_19995);
or UO_458 (O_458,N_19939,N_19926);
xnor UO_459 (O_459,N_19862,N_19877);
or UO_460 (O_460,N_19864,N_19929);
nor UO_461 (O_461,N_19956,N_19953);
nor UO_462 (O_462,N_19955,N_19857);
nor UO_463 (O_463,N_19968,N_19905);
nor UO_464 (O_464,N_19988,N_19893);
and UO_465 (O_465,N_19926,N_19913);
nand UO_466 (O_466,N_19999,N_19943);
nand UO_467 (O_467,N_19852,N_19988);
nand UO_468 (O_468,N_19854,N_19985);
nand UO_469 (O_469,N_19949,N_19992);
or UO_470 (O_470,N_19977,N_19952);
nor UO_471 (O_471,N_19891,N_19871);
nor UO_472 (O_472,N_19987,N_19936);
xnor UO_473 (O_473,N_19869,N_19893);
nor UO_474 (O_474,N_19958,N_19843);
nand UO_475 (O_475,N_19858,N_19889);
nand UO_476 (O_476,N_19861,N_19882);
xnor UO_477 (O_477,N_19917,N_19881);
nor UO_478 (O_478,N_19852,N_19960);
or UO_479 (O_479,N_19995,N_19895);
nand UO_480 (O_480,N_19983,N_19882);
or UO_481 (O_481,N_19886,N_19937);
and UO_482 (O_482,N_19992,N_19918);
or UO_483 (O_483,N_19913,N_19922);
or UO_484 (O_484,N_19841,N_19929);
or UO_485 (O_485,N_19871,N_19849);
nor UO_486 (O_486,N_19848,N_19925);
nor UO_487 (O_487,N_19937,N_19842);
nor UO_488 (O_488,N_19847,N_19913);
xor UO_489 (O_489,N_19981,N_19920);
and UO_490 (O_490,N_19872,N_19900);
and UO_491 (O_491,N_19890,N_19906);
nand UO_492 (O_492,N_19886,N_19942);
nor UO_493 (O_493,N_19920,N_19861);
and UO_494 (O_494,N_19845,N_19905);
or UO_495 (O_495,N_19951,N_19953);
or UO_496 (O_496,N_19923,N_19858);
xor UO_497 (O_497,N_19916,N_19978);
and UO_498 (O_498,N_19991,N_19930);
or UO_499 (O_499,N_19990,N_19959);
xnor UO_500 (O_500,N_19848,N_19895);
nor UO_501 (O_501,N_19991,N_19891);
nor UO_502 (O_502,N_19963,N_19896);
xnor UO_503 (O_503,N_19869,N_19878);
xnor UO_504 (O_504,N_19891,N_19951);
and UO_505 (O_505,N_19933,N_19922);
or UO_506 (O_506,N_19964,N_19862);
and UO_507 (O_507,N_19953,N_19938);
or UO_508 (O_508,N_19949,N_19951);
and UO_509 (O_509,N_19943,N_19850);
xor UO_510 (O_510,N_19947,N_19952);
and UO_511 (O_511,N_19878,N_19922);
or UO_512 (O_512,N_19925,N_19995);
nor UO_513 (O_513,N_19847,N_19967);
and UO_514 (O_514,N_19975,N_19997);
xnor UO_515 (O_515,N_19892,N_19891);
nand UO_516 (O_516,N_19880,N_19978);
xnor UO_517 (O_517,N_19928,N_19989);
nor UO_518 (O_518,N_19870,N_19861);
xor UO_519 (O_519,N_19852,N_19947);
or UO_520 (O_520,N_19938,N_19933);
nand UO_521 (O_521,N_19866,N_19966);
xor UO_522 (O_522,N_19852,N_19863);
or UO_523 (O_523,N_19935,N_19890);
nor UO_524 (O_524,N_19983,N_19896);
and UO_525 (O_525,N_19872,N_19987);
nor UO_526 (O_526,N_19900,N_19914);
nor UO_527 (O_527,N_19856,N_19907);
or UO_528 (O_528,N_19988,N_19888);
and UO_529 (O_529,N_19864,N_19931);
or UO_530 (O_530,N_19889,N_19924);
or UO_531 (O_531,N_19905,N_19848);
nand UO_532 (O_532,N_19962,N_19864);
nor UO_533 (O_533,N_19993,N_19891);
and UO_534 (O_534,N_19883,N_19870);
and UO_535 (O_535,N_19844,N_19906);
xor UO_536 (O_536,N_19951,N_19923);
nand UO_537 (O_537,N_19913,N_19871);
nor UO_538 (O_538,N_19947,N_19937);
xor UO_539 (O_539,N_19885,N_19862);
or UO_540 (O_540,N_19987,N_19935);
xor UO_541 (O_541,N_19961,N_19901);
nand UO_542 (O_542,N_19950,N_19929);
nor UO_543 (O_543,N_19935,N_19925);
nand UO_544 (O_544,N_19951,N_19964);
nor UO_545 (O_545,N_19913,N_19949);
or UO_546 (O_546,N_19922,N_19899);
and UO_547 (O_547,N_19973,N_19972);
nor UO_548 (O_548,N_19862,N_19956);
or UO_549 (O_549,N_19962,N_19843);
nor UO_550 (O_550,N_19901,N_19849);
and UO_551 (O_551,N_19961,N_19937);
and UO_552 (O_552,N_19947,N_19978);
nor UO_553 (O_553,N_19924,N_19981);
xor UO_554 (O_554,N_19911,N_19986);
nor UO_555 (O_555,N_19900,N_19949);
xor UO_556 (O_556,N_19881,N_19977);
or UO_557 (O_557,N_19946,N_19874);
xor UO_558 (O_558,N_19847,N_19851);
or UO_559 (O_559,N_19953,N_19853);
xnor UO_560 (O_560,N_19871,N_19877);
nor UO_561 (O_561,N_19955,N_19890);
or UO_562 (O_562,N_19881,N_19998);
nor UO_563 (O_563,N_19854,N_19962);
and UO_564 (O_564,N_19882,N_19937);
nand UO_565 (O_565,N_19873,N_19985);
xnor UO_566 (O_566,N_19924,N_19984);
nand UO_567 (O_567,N_19923,N_19908);
xor UO_568 (O_568,N_19907,N_19857);
xnor UO_569 (O_569,N_19969,N_19876);
nand UO_570 (O_570,N_19947,N_19941);
or UO_571 (O_571,N_19986,N_19863);
nor UO_572 (O_572,N_19915,N_19861);
nand UO_573 (O_573,N_19864,N_19842);
xnor UO_574 (O_574,N_19861,N_19985);
or UO_575 (O_575,N_19998,N_19880);
xnor UO_576 (O_576,N_19908,N_19929);
nor UO_577 (O_577,N_19846,N_19972);
and UO_578 (O_578,N_19923,N_19857);
nor UO_579 (O_579,N_19944,N_19877);
or UO_580 (O_580,N_19960,N_19887);
nor UO_581 (O_581,N_19986,N_19924);
xor UO_582 (O_582,N_19912,N_19965);
and UO_583 (O_583,N_19884,N_19863);
nand UO_584 (O_584,N_19858,N_19867);
nand UO_585 (O_585,N_19981,N_19999);
or UO_586 (O_586,N_19944,N_19858);
nand UO_587 (O_587,N_19984,N_19872);
or UO_588 (O_588,N_19960,N_19875);
or UO_589 (O_589,N_19890,N_19846);
and UO_590 (O_590,N_19877,N_19970);
nor UO_591 (O_591,N_19962,N_19985);
nor UO_592 (O_592,N_19954,N_19932);
xor UO_593 (O_593,N_19886,N_19968);
or UO_594 (O_594,N_19948,N_19888);
xnor UO_595 (O_595,N_19978,N_19857);
xnor UO_596 (O_596,N_19933,N_19959);
xor UO_597 (O_597,N_19954,N_19885);
xnor UO_598 (O_598,N_19992,N_19946);
nand UO_599 (O_599,N_19857,N_19882);
and UO_600 (O_600,N_19936,N_19849);
nand UO_601 (O_601,N_19874,N_19974);
nor UO_602 (O_602,N_19983,N_19997);
xor UO_603 (O_603,N_19989,N_19937);
and UO_604 (O_604,N_19858,N_19978);
and UO_605 (O_605,N_19910,N_19878);
and UO_606 (O_606,N_19991,N_19866);
and UO_607 (O_607,N_19849,N_19925);
nor UO_608 (O_608,N_19983,N_19872);
nor UO_609 (O_609,N_19935,N_19905);
and UO_610 (O_610,N_19843,N_19910);
and UO_611 (O_611,N_19845,N_19930);
nor UO_612 (O_612,N_19906,N_19991);
or UO_613 (O_613,N_19957,N_19844);
and UO_614 (O_614,N_19917,N_19904);
and UO_615 (O_615,N_19910,N_19870);
and UO_616 (O_616,N_19939,N_19960);
or UO_617 (O_617,N_19952,N_19992);
xor UO_618 (O_618,N_19895,N_19931);
nor UO_619 (O_619,N_19931,N_19974);
nor UO_620 (O_620,N_19900,N_19860);
nand UO_621 (O_621,N_19985,N_19933);
nand UO_622 (O_622,N_19904,N_19854);
xor UO_623 (O_623,N_19900,N_19964);
and UO_624 (O_624,N_19965,N_19954);
and UO_625 (O_625,N_19973,N_19966);
nor UO_626 (O_626,N_19893,N_19914);
xnor UO_627 (O_627,N_19980,N_19925);
nor UO_628 (O_628,N_19968,N_19960);
or UO_629 (O_629,N_19999,N_19847);
xnor UO_630 (O_630,N_19889,N_19840);
and UO_631 (O_631,N_19859,N_19924);
or UO_632 (O_632,N_19909,N_19866);
and UO_633 (O_633,N_19985,N_19998);
and UO_634 (O_634,N_19841,N_19935);
xor UO_635 (O_635,N_19905,N_19994);
xor UO_636 (O_636,N_19877,N_19991);
nor UO_637 (O_637,N_19903,N_19924);
xnor UO_638 (O_638,N_19983,N_19923);
nand UO_639 (O_639,N_19932,N_19846);
and UO_640 (O_640,N_19925,N_19892);
or UO_641 (O_641,N_19864,N_19913);
or UO_642 (O_642,N_19856,N_19987);
nor UO_643 (O_643,N_19907,N_19910);
or UO_644 (O_644,N_19923,N_19961);
or UO_645 (O_645,N_19850,N_19970);
or UO_646 (O_646,N_19862,N_19967);
nor UO_647 (O_647,N_19979,N_19843);
xnor UO_648 (O_648,N_19985,N_19944);
or UO_649 (O_649,N_19847,N_19893);
xor UO_650 (O_650,N_19956,N_19965);
or UO_651 (O_651,N_19900,N_19929);
nand UO_652 (O_652,N_19985,N_19874);
xor UO_653 (O_653,N_19906,N_19990);
nor UO_654 (O_654,N_19909,N_19929);
or UO_655 (O_655,N_19924,N_19888);
nor UO_656 (O_656,N_19990,N_19930);
nor UO_657 (O_657,N_19879,N_19845);
nand UO_658 (O_658,N_19910,N_19865);
or UO_659 (O_659,N_19931,N_19910);
nand UO_660 (O_660,N_19936,N_19899);
and UO_661 (O_661,N_19878,N_19951);
nand UO_662 (O_662,N_19956,N_19964);
xnor UO_663 (O_663,N_19916,N_19949);
nand UO_664 (O_664,N_19998,N_19956);
and UO_665 (O_665,N_19976,N_19893);
and UO_666 (O_666,N_19922,N_19872);
xnor UO_667 (O_667,N_19862,N_19889);
nand UO_668 (O_668,N_19978,N_19926);
nand UO_669 (O_669,N_19925,N_19899);
nand UO_670 (O_670,N_19862,N_19918);
nand UO_671 (O_671,N_19928,N_19954);
or UO_672 (O_672,N_19928,N_19946);
or UO_673 (O_673,N_19972,N_19971);
xnor UO_674 (O_674,N_19997,N_19973);
nor UO_675 (O_675,N_19880,N_19979);
or UO_676 (O_676,N_19879,N_19897);
or UO_677 (O_677,N_19900,N_19931);
and UO_678 (O_678,N_19948,N_19870);
xor UO_679 (O_679,N_19868,N_19911);
xnor UO_680 (O_680,N_19977,N_19915);
or UO_681 (O_681,N_19984,N_19986);
and UO_682 (O_682,N_19924,N_19850);
xnor UO_683 (O_683,N_19960,N_19940);
xor UO_684 (O_684,N_19995,N_19993);
nand UO_685 (O_685,N_19908,N_19902);
or UO_686 (O_686,N_19929,N_19992);
nor UO_687 (O_687,N_19941,N_19895);
and UO_688 (O_688,N_19849,N_19931);
nor UO_689 (O_689,N_19977,N_19954);
xor UO_690 (O_690,N_19841,N_19906);
xnor UO_691 (O_691,N_19854,N_19940);
or UO_692 (O_692,N_19989,N_19969);
nor UO_693 (O_693,N_19897,N_19969);
and UO_694 (O_694,N_19983,N_19979);
xor UO_695 (O_695,N_19977,N_19852);
nand UO_696 (O_696,N_19971,N_19846);
nor UO_697 (O_697,N_19906,N_19931);
nand UO_698 (O_698,N_19939,N_19974);
nor UO_699 (O_699,N_19935,N_19957);
xor UO_700 (O_700,N_19885,N_19842);
nor UO_701 (O_701,N_19856,N_19891);
and UO_702 (O_702,N_19937,N_19884);
nand UO_703 (O_703,N_19996,N_19922);
nor UO_704 (O_704,N_19976,N_19981);
nand UO_705 (O_705,N_19970,N_19888);
nand UO_706 (O_706,N_19878,N_19917);
nand UO_707 (O_707,N_19852,N_19991);
xnor UO_708 (O_708,N_19880,N_19944);
xnor UO_709 (O_709,N_19947,N_19981);
nor UO_710 (O_710,N_19871,N_19847);
xnor UO_711 (O_711,N_19863,N_19908);
nand UO_712 (O_712,N_19889,N_19927);
nand UO_713 (O_713,N_19946,N_19971);
and UO_714 (O_714,N_19949,N_19940);
nand UO_715 (O_715,N_19973,N_19888);
nand UO_716 (O_716,N_19980,N_19949);
nor UO_717 (O_717,N_19861,N_19999);
xor UO_718 (O_718,N_19918,N_19865);
nor UO_719 (O_719,N_19879,N_19931);
nand UO_720 (O_720,N_19848,N_19916);
xor UO_721 (O_721,N_19940,N_19907);
nand UO_722 (O_722,N_19902,N_19921);
nand UO_723 (O_723,N_19991,N_19968);
or UO_724 (O_724,N_19850,N_19954);
nor UO_725 (O_725,N_19894,N_19883);
xnor UO_726 (O_726,N_19903,N_19967);
and UO_727 (O_727,N_19983,N_19856);
or UO_728 (O_728,N_19908,N_19983);
and UO_729 (O_729,N_19953,N_19851);
nor UO_730 (O_730,N_19952,N_19841);
nand UO_731 (O_731,N_19854,N_19848);
xnor UO_732 (O_732,N_19963,N_19916);
nand UO_733 (O_733,N_19940,N_19891);
and UO_734 (O_734,N_19943,N_19986);
nand UO_735 (O_735,N_19843,N_19957);
and UO_736 (O_736,N_19869,N_19853);
nand UO_737 (O_737,N_19970,N_19847);
nand UO_738 (O_738,N_19860,N_19946);
xnor UO_739 (O_739,N_19942,N_19969);
nand UO_740 (O_740,N_19890,N_19975);
or UO_741 (O_741,N_19986,N_19871);
xnor UO_742 (O_742,N_19973,N_19921);
xor UO_743 (O_743,N_19955,N_19910);
nor UO_744 (O_744,N_19932,N_19931);
xnor UO_745 (O_745,N_19852,N_19972);
xor UO_746 (O_746,N_19970,N_19996);
xor UO_747 (O_747,N_19909,N_19951);
xnor UO_748 (O_748,N_19937,N_19907);
nor UO_749 (O_749,N_19988,N_19947);
nand UO_750 (O_750,N_19976,N_19995);
and UO_751 (O_751,N_19883,N_19920);
nand UO_752 (O_752,N_19884,N_19877);
nand UO_753 (O_753,N_19855,N_19907);
and UO_754 (O_754,N_19931,N_19899);
or UO_755 (O_755,N_19906,N_19929);
nor UO_756 (O_756,N_19906,N_19877);
and UO_757 (O_757,N_19840,N_19972);
nor UO_758 (O_758,N_19936,N_19930);
xor UO_759 (O_759,N_19923,N_19988);
or UO_760 (O_760,N_19985,N_19903);
nand UO_761 (O_761,N_19940,N_19939);
nor UO_762 (O_762,N_19885,N_19905);
nand UO_763 (O_763,N_19949,N_19874);
xnor UO_764 (O_764,N_19944,N_19888);
and UO_765 (O_765,N_19892,N_19970);
xnor UO_766 (O_766,N_19949,N_19977);
nor UO_767 (O_767,N_19849,N_19899);
or UO_768 (O_768,N_19877,N_19989);
or UO_769 (O_769,N_19840,N_19997);
nand UO_770 (O_770,N_19894,N_19893);
xnor UO_771 (O_771,N_19956,N_19858);
nand UO_772 (O_772,N_19990,N_19957);
and UO_773 (O_773,N_19845,N_19958);
or UO_774 (O_774,N_19966,N_19945);
and UO_775 (O_775,N_19963,N_19965);
and UO_776 (O_776,N_19978,N_19854);
or UO_777 (O_777,N_19918,N_19863);
xnor UO_778 (O_778,N_19921,N_19857);
xor UO_779 (O_779,N_19931,N_19904);
and UO_780 (O_780,N_19942,N_19918);
and UO_781 (O_781,N_19890,N_19971);
xnor UO_782 (O_782,N_19862,N_19934);
nor UO_783 (O_783,N_19919,N_19859);
nor UO_784 (O_784,N_19903,N_19956);
and UO_785 (O_785,N_19975,N_19893);
nor UO_786 (O_786,N_19883,N_19914);
nand UO_787 (O_787,N_19846,N_19872);
or UO_788 (O_788,N_19947,N_19998);
nand UO_789 (O_789,N_19855,N_19898);
and UO_790 (O_790,N_19951,N_19941);
or UO_791 (O_791,N_19955,N_19938);
or UO_792 (O_792,N_19902,N_19886);
nand UO_793 (O_793,N_19855,N_19924);
and UO_794 (O_794,N_19930,N_19872);
nand UO_795 (O_795,N_19930,N_19946);
nor UO_796 (O_796,N_19979,N_19981);
nor UO_797 (O_797,N_19932,N_19991);
xor UO_798 (O_798,N_19900,N_19885);
nor UO_799 (O_799,N_19946,N_19993);
or UO_800 (O_800,N_19851,N_19916);
or UO_801 (O_801,N_19947,N_19915);
xnor UO_802 (O_802,N_19865,N_19925);
or UO_803 (O_803,N_19932,N_19986);
xnor UO_804 (O_804,N_19884,N_19895);
xnor UO_805 (O_805,N_19882,N_19931);
nand UO_806 (O_806,N_19873,N_19984);
xnor UO_807 (O_807,N_19950,N_19866);
or UO_808 (O_808,N_19877,N_19886);
nor UO_809 (O_809,N_19953,N_19950);
xnor UO_810 (O_810,N_19874,N_19868);
nor UO_811 (O_811,N_19860,N_19943);
nor UO_812 (O_812,N_19965,N_19990);
nor UO_813 (O_813,N_19897,N_19913);
and UO_814 (O_814,N_19869,N_19923);
or UO_815 (O_815,N_19901,N_19878);
nand UO_816 (O_816,N_19994,N_19985);
and UO_817 (O_817,N_19913,N_19955);
nor UO_818 (O_818,N_19998,N_19960);
xor UO_819 (O_819,N_19946,N_19891);
nor UO_820 (O_820,N_19980,N_19853);
nand UO_821 (O_821,N_19938,N_19968);
nor UO_822 (O_822,N_19911,N_19996);
nor UO_823 (O_823,N_19853,N_19987);
nor UO_824 (O_824,N_19997,N_19845);
or UO_825 (O_825,N_19979,N_19972);
and UO_826 (O_826,N_19957,N_19895);
xor UO_827 (O_827,N_19946,N_19995);
nand UO_828 (O_828,N_19908,N_19918);
xnor UO_829 (O_829,N_19842,N_19893);
or UO_830 (O_830,N_19953,N_19954);
nor UO_831 (O_831,N_19971,N_19988);
and UO_832 (O_832,N_19977,N_19953);
xor UO_833 (O_833,N_19930,N_19864);
nor UO_834 (O_834,N_19889,N_19886);
nor UO_835 (O_835,N_19872,N_19920);
and UO_836 (O_836,N_19985,N_19940);
nand UO_837 (O_837,N_19845,N_19936);
nor UO_838 (O_838,N_19905,N_19946);
nor UO_839 (O_839,N_19877,N_19982);
xor UO_840 (O_840,N_19941,N_19866);
or UO_841 (O_841,N_19893,N_19904);
xor UO_842 (O_842,N_19967,N_19970);
and UO_843 (O_843,N_19848,N_19941);
nand UO_844 (O_844,N_19849,N_19944);
or UO_845 (O_845,N_19985,N_19902);
and UO_846 (O_846,N_19907,N_19874);
xnor UO_847 (O_847,N_19865,N_19869);
and UO_848 (O_848,N_19921,N_19843);
nor UO_849 (O_849,N_19957,N_19847);
xnor UO_850 (O_850,N_19971,N_19840);
xnor UO_851 (O_851,N_19983,N_19888);
nand UO_852 (O_852,N_19978,N_19996);
nor UO_853 (O_853,N_19914,N_19992);
or UO_854 (O_854,N_19856,N_19941);
nor UO_855 (O_855,N_19868,N_19936);
or UO_856 (O_856,N_19922,N_19897);
xor UO_857 (O_857,N_19853,N_19879);
xor UO_858 (O_858,N_19876,N_19953);
nor UO_859 (O_859,N_19990,N_19999);
nor UO_860 (O_860,N_19851,N_19959);
and UO_861 (O_861,N_19900,N_19894);
nor UO_862 (O_862,N_19951,N_19934);
nand UO_863 (O_863,N_19925,N_19857);
or UO_864 (O_864,N_19966,N_19960);
xnor UO_865 (O_865,N_19971,N_19881);
xnor UO_866 (O_866,N_19881,N_19940);
and UO_867 (O_867,N_19840,N_19932);
nand UO_868 (O_868,N_19894,N_19862);
or UO_869 (O_869,N_19884,N_19851);
or UO_870 (O_870,N_19979,N_19988);
or UO_871 (O_871,N_19848,N_19871);
and UO_872 (O_872,N_19862,N_19994);
or UO_873 (O_873,N_19871,N_19974);
xor UO_874 (O_874,N_19998,N_19898);
or UO_875 (O_875,N_19935,N_19856);
or UO_876 (O_876,N_19949,N_19860);
and UO_877 (O_877,N_19883,N_19868);
xor UO_878 (O_878,N_19853,N_19855);
xor UO_879 (O_879,N_19956,N_19843);
and UO_880 (O_880,N_19948,N_19851);
or UO_881 (O_881,N_19859,N_19999);
nand UO_882 (O_882,N_19864,N_19967);
xor UO_883 (O_883,N_19935,N_19926);
nand UO_884 (O_884,N_19931,N_19902);
nor UO_885 (O_885,N_19951,N_19916);
and UO_886 (O_886,N_19964,N_19998);
and UO_887 (O_887,N_19859,N_19969);
xor UO_888 (O_888,N_19915,N_19844);
nand UO_889 (O_889,N_19998,N_19920);
or UO_890 (O_890,N_19912,N_19935);
nor UO_891 (O_891,N_19995,N_19875);
or UO_892 (O_892,N_19865,N_19908);
or UO_893 (O_893,N_19861,N_19978);
and UO_894 (O_894,N_19913,N_19905);
nor UO_895 (O_895,N_19847,N_19983);
xnor UO_896 (O_896,N_19991,N_19977);
nor UO_897 (O_897,N_19845,N_19978);
and UO_898 (O_898,N_19970,N_19945);
xor UO_899 (O_899,N_19860,N_19902);
or UO_900 (O_900,N_19952,N_19849);
or UO_901 (O_901,N_19982,N_19953);
nor UO_902 (O_902,N_19900,N_19975);
xor UO_903 (O_903,N_19962,N_19923);
nand UO_904 (O_904,N_19906,N_19861);
nor UO_905 (O_905,N_19902,N_19917);
xnor UO_906 (O_906,N_19975,N_19923);
nand UO_907 (O_907,N_19959,N_19970);
xnor UO_908 (O_908,N_19877,N_19856);
nor UO_909 (O_909,N_19922,N_19952);
and UO_910 (O_910,N_19976,N_19954);
nor UO_911 (O_911,N_19896,N_19904);
and UO_912 (O_912,N_19928,N_19935);
or UO_913 (O_913,N_19893,N_19906);
or UO_914 (O_914,N_19882,N_19897);
xor UO_915 (O_915,N_19918,N_19967);
xnor UO_916 (O_916,N_19886,N_19932);
xnor UO_917 (O_917,N_19934,N_19880);
nand UO_918 (O_918,N_19840,N_19989);
and UO_919 (O_919,N_19937,N_19874);
or UO_920 (O_920,N_19912,N_19878);
nor UO_921 (O_921,N_19888,N_19932);
xor UO_922 (O_922,N_19898,N_19872);
and UO_923 (O_923,N_19964,N_19898);
nor UO_924 (O_924,N_19897,N_19941);
xor UO_925 (O_925,N_19874,N_19916);
and UO_926 (O_926,N_19948,N_19957);
nor UO_927 (O_927,N_19994,N_19876);
nand UO_928 (O_928,N_19904,N_19944);
and UO_929 (O_929,N_19884,N_19881);
nor UO_930 (O_930,N_19858,N_19881);
nand UO_931 (O_931,N_19962,N_19907);
or UO_932 (O_932,N_19857,N_19911);
nor UO_933 (O_933,N_19890,N_19925);
nand UO_934 (O_934,N_19898,N_19955);
or UO_935 (O_935,N_19863,N_19977);
nor UO_936 (O_936,N_19932,N_19946);
nand UO_937 (O_937,N_19894,N_19960);
and UO_938 (O_938,N_19964,N_19882);
or UO_939 (O_939,N_19992,N_19875);
nor UO_940 (O_940,N_19941,N_19894);
nand UO_941 (O_941,N_19990,N_19857);
nand UO_942 (O_942,N_19908,N_19972);
nor UO_943 (O_943,N_19857,N_19952);
or UO_944 (O_944,N_19999,N_19913);
and UO_945 (O_945,N_19896,N_19928);
nor UO_946 (O_946,N_19989,N_19890);
nor UO_947 (O_947,N_19926,N_19928);
or UO_948 (O_948,N_19934,N_19861);
xor UO_949 (O_949,N_19951,N_19989);
or UO_950 (O_950,N_19856,N_19841);
and UO_951 (O_951,N_19875,N_19962);
xnor UO_952 (O_952,N_19909,N_19942);
and UO_953 (O_953,N_19926,N_19994);
nor UO_954 (O_954,N_19847,N_19862);
and UO_955 (O_955,N_19981,N_19927);
or UO_956 (O_956,N_19845,N_19876);
and UO_957 (O_957,N_19863,N_19915);
and UO_958 (O_958,N_19895,N_19927);
xor UO_959 (O_959,N_19932,N_19921);
and UO_960 (O_960,N_19896,N_19948);
nor UO_961 (O_961,N_19969,N_19863);
or UO_962 (O_962,N_19980,N_19910);
and UO_963 (O_963,N_19931,N_19908);
xnor UO_964 (O_964,N_19876,N_19913);
nand UO_965 (O_965,N_19859,N_19947);
nor UO_966 (O_966,N_19879,N_19854);
and UO_967 (O_967,N_19865,N_19858);
or UO_968 (O_968,N_19982,N_19867);
or UO_969 (O_969,N_19897,N_19858);
nand UO_970 (O_970,N_19846,N_19902);
nand UO_971 (O_971,N_19887,N_19987);
or UO_972 (O_972,N_19848,N_19852);
or UO_973 (O_973,N_19918,N_19948);
xor UO_974 (O_974,N_19911,N_19972);
nor UO_975 (O_975,N_19929,N_19997);
and UO_976 (O_976,N_19988,N_19998);
nand UO_977 (O_977,N_19969,N_19901);
nand UO_978 (O_978,N_19929,N_19886);
xor UO_979 (O_979,N_19894,N_19967);
nand UO_980 (O_980,N_19964,N_19908);
and UO_981 (O_981,N_19992,N_19975);
nand UO_982 (O_982,N_19895,N_19872);
nand UO_983 (O_983,N_19977,N_19872);
nor UO_984 (O_984,N_19847,N_19865);
and UO_985 (O_985,N_19861,N_19860);
or UO_986 (O_986,N_19994,N_19875);
xnor UO_987 (O_987,N_19903,N_19901);
nand UO_988 (O_988,N_19872,N_19887);
or UO_989 (O_989,N_19905,N_19898);
and UO_990 (O_990,N_19848,N_19995);
xor UO_991 (O_991,N_19891,N_19852);
nor UO_992 (O_992,N_19853,N_19913);
nor UO_993 (O_993,N_19854,N_19959);
nor UO_994 (O_994,N_19843,N_19969);
nor UO_995 (O_995,N_19973,N_19920);
or UO_996 (O_996,N_19841,N_19939);
nand UO_997 (O_997,N_19945,N_19946);
nor UO_998 (O_998,N_19905,N_19969);
xor UO_999 (O_999,N_19997,N_19940);
or UO_1000 (O_1000,N_19999,N_19942);
or UO_1001 (O_1001,N_19954,N_19950);
and UO_1002 (O_1002,N_19997,N_19937);
or UO_1003 (O_1003,N_19894,N_19950);
xnor UO_1004 (O_1004,N_19920,N_19850);
nor UO_1005 (O_1005,N_19918,N_19998);
nor UO_1006 (O_1006,N_19914,N_19932);
nand UO_1007 (O_1007,N_19913,N_19909);
or UO_1008 (O_1008,N_19961,N_19993);
and UO_1009 (O_1009,N_19979,N_19973);
nand UO_1010 (O_1010,N_19951,N_19979);
and UO_1011 (O_1011,N_19958,N_19882);
nor UO_1012 (O_1012,N_19907,N_19999);
or UO_1013 (O_1013,N_19997,N_19902);
nand UO_1014 (O_1014,N_19910,N_19908);
or UO_1015 (O_1015,N_19906,N_19866);
and UO_1016 (O_1016,N_19895,N_19847);
nand UO_1017 (O_1017,N_19920,N_19889);
xnor UO_1018 (O_1018,N_19973,N_19876);
nor UO_1019 (O_1019,N_19985,N_19949);
xnor UO_1020 (O_1020,N_19976,N_19917);
or UO_1021 (O_1021,N_19921,N_19926);
or UO_1022 (O_1022,N_19943,N_19855);
nor UO_1023 (O_1023,N_19878,N_19942);
and UO_1024 (O_1024,N_19915,N_19937);
xor UO_1025 (O_1025,N_19889,N_19913);
xnor UO_1026 (O_1026,N_19871,N_19864);
nor UO_1027 (O_1027,N_19970,N_19930);
or UO_1028 (O_1028,N_19923,N_19998);
nand UO_1029 (O_1029,N_19960,N_19877);
nor UO_1030 (O_1030,N_19910,N_19845);
xor UO_1031 (O_1031,N_19850,N_19847);
nand UO_1032 (O_1032,N_19856,N_19869);
nor UO_1033 (O_1033,N_19898,N_19906);
xnor UO_1034 (O_1034,N_19873,N_19898);
or UO_1035 (O_1035,N_19987,N_19871);
nand UO_1036 (O_1036,N_19953,N_19936);
xnor UO_1037 (O_1037,N_19972,N_19968);
and UO_1038 (O_1038,N_19966,N_19948);
or UO_1039 (O_1039,N_19966,N_19996);
nand UO_1040 (O_1040,N_19878,N_19890);
or UO_1041 (O_1041,N_19860,N_19845);
or UO_1042 (O_1042,N_19902,N_19906);
and UO_1043 (O_1043,N_19905,N_19917);
nor UO_1044 (O_1044,N_19923,N_19912);
nand UO_1045 (O_1045,N_19889,N_19863);
xor UO_1046 (O_1046,N_19962,N_19879);
and UO_1047 (O_1047,N_19857,N_19985);
and UO_1048 (O_1048,N_19972,N_19948);
nor UO_1049 (O_1049,N_19957,N_19908);
xnor UO_1050 (O_1050,N_19919,N_19979);
or UO_1051 (O_1051,N_19898,N_19939);
nand UO_1052 (O_1052,N_19998,N_19888);
nand UO_1053 (O_1053,N_19854,N_19954);
and UO_1054 (O_1054,N_19998,N_19846);
or UO_1055 (O_1055,N_19963,N_19949);
and UO_1056 (O_1056,N_19982,N_19897);
nand UO_1057 (O_1057,N_19893,N_19858);
or UO_1058 (O_1058,N_19946,N_19977);
nand UO_1059 (O_1059,N_19891,N_19939);
and UO_1060 (O_1060,N_19939,N_19983);
nand UO_1061 (O_1061,N_19934,N_19920);
and UO_1062 (O_1062,N_19859,N_19946);
nor UO_1063 (O_1063,N_19863,N_19879);
nand UO_1064 (O_1064,N_19949,N_19919);
and UO_1065 (O_1065,N_19986,N_19959);
nor UO_1066 (O_1066,N_19895,N_19976);
nand UO_1067 (O_1067,N_19855,N_19878);
xnor UO_1068 (O_1068,N_19845,N_19960);
nand UO_1069 (O_1069,N_19977,N_19901);
nor UO_1070 (O_1070,N_19964,N_19860);
and UO_1071 (O_1071,N_19993,N_19877);
nand UO_1072 (O_1072,N_19888,N_19971);
nor UO_1073 (O_1073,N_19867,N_19910);
and UO_1074 (O_1074,N_19940,N_19892);
or UO_1075 (O_1075,N_19966,N_19909);
or UO_1076 (O_1076,N_19867,N_19970);
or UO_1077 (O_1077,N_19900,N_19992);
nor UO_1078 (O_1078,N_19875,N_19940);
or UO_1079 (O_1079,N_19850,N_19950);
or UO_1080 (O_1080,N_19874,N_19979);
nand UO_1081 (O_1081,N_19977,N_19919);
xor UO_1082 (O_1082,N_19890,N_19956);
and UO_1083 (O_1083,N_19934,N_19953);
or UO_1084 (O_1084,N_19878,N_19955);
nand UO_1085 (O_1085,N_19883,N_19874);
nor UO_1086 (O_1086,N_19959,N_19879);
nand UO_1087 (O_1087,N_19856,N_19926);
nor UO_1088 (O_1088,N_19960,N_19947);
nand UO_1089 (O_1089,N_19883,N_19924);
nand UO_1090 (O_1090,N_19909,N_19893);
or UO_1091 (O_1091,N_19906,N_19969);
nand UO_1092 (O_1092,N_19853,N_19881);
xor UO_1093 (O_1093,N_19966,N_19900);
nand UO_1094 (O_1094,N_19862,N_19896);
xor UO_1095 (O_1095,N_19878,N_19994);
and UO_1096 (O_1096,N_19863,N_19956);
nand UO_1097 (O_1097,N_19896,N_19886);
or UO_1098 (O_1098,N_19853,N_19923);
nand UO_1099 (O_1099,N_19860,N_19978);
or UO_1100 (O_1100,N_19994,N_19991);
nor UO_1101 (O_1101,N_19863,N_19878);
nand UO_1102 (O_1102,N_19892,N_19921);
or UO_1103 (O_1103,N_19861,N_19890);
or UO_1104 (O_1104,N_19923,N_19891);
nand UO_1105 (O_1105,N_19990,N_19973);
and UO_1106 (O_1106,N_19952,N_19917);
nor UO_1107 (O_1107,N_19965,N_19855);
xor UO_1108 (O_1108,N_19925,N_19895);
xnor UO_1109 (O_1109,N_19920,N_19893);
nand UO_1110 (O_1110,N_19937,N_19944);
or UO_1111 (O_1111,N_19935,N_19896);
nor UO_1112 (O_1112,N_19926,N_19851);
or UO_1113 (O_1113,N_19898,N_19877);
xor UO_1114 (O_1114,N_19943,N_19931);
nor UO_1115 (O_1115,N_19940,N_19933);
xnor UO_1116 (O_1116,N_19993,N_19908);
nor UO_1117 (O_1117,N_19918,N_19920);
nand UO_1118 (O_1118,N_19912,N_19934);
nor UO_1119 (O_1119,N_19925,N_19955);
nor UO_1120 (O_1120,N_19949,N_19888);
nand UO_1121 (O_1121,N_19917,N_19968);
nor UO_1122 (O_1122,N_19987,N_19873);
and UO_1123 (O_1123,N_19850,N_19840);
or UO_1124 (O_1124,N_19855,N_19873);
or UO_1125 (O_1125,N_19961,N_19866);
or UO_1126 (O_1126,N_19897,N_19889);
nor UO_1127 (O_1127,N_19951,N_19936);
xor UO_1128 (O_1128,N_19932,N_19858);
nand UO_1129 (O_1129,N_19973,N_19887);
xor UO_1130 (O_1130,N_19856,N_19970);
nand UO_1131 (O_1131,N_19844,N_19954);
and UO_1132 (O_1132,N_19949,N_19922);
nand UO_1133 (O_1133,N_19872,N_19875);
or UO_1134 (O_1134,N_19983,N_19895);
or UO_1135 (O_1135,N_19901,N_19921);
nand UO_1136 (O_1136,N_19956,N_19878);
nor UO_1137 (O_1137,N_19848,N_19940);
nand UO_1138 (O_1138,N_19863,N_19979);
or UO_1139 (O_1139,N_19884,N_19973);
nor UO_1140 (O_1140,N_19841,N_19847);
nor UO_1141 (O_1141,N_19917,N_19897);
xnor UO_1142 (O_1142,N_19980,N_19915);
or UO_1143 (O_1143,N_19965,N_19988);
nor UO_1144 (O_1144,N_19902,N_19942);
or UO_1145 (O_1145,N_19883,N_19903);
xnor UO_1146 (O_1146,N_19842,N_19970);
nor UO_1147 (O_1147,N_19926,N_19914);
nor UO_1148 (O_1148,N_19873,N_19998);
xor UO_1149 (O_1149,N_19856,N_19992);
xor UO_1150 (O_1150,N_19868,N_19970);
xor UO_1151 (O_1151,N_19931,N_19990);
or UO_1152 (O_1152,N_19936,N_19909);
and UO_1153 (O_1153,N_19943,N_19971);
xnor UO_1154 (O_1154,N_19930,N_19934);
nor UO_1155 (O_1155,N_19957,N_19986);
or UO_1156 (O_1156,N_19842,N_19945);
xor UO_1157 (O_1157,N_19888,N_19984);
xnor UO_1158 (O_1158,N_19975,N_19870);
and UO_1159 (O_1159,N_19913,N_19858);
xnor UO_1160 (O_1160,N_19891,N_19958);
nand UO_1161 (O_1161,N_19955,N_19919);
and UO_1162 (O_1162,N_19873,N_19961);
xnor UO_1163 (O_1163,N_19979,N_19931);
nor UO_1164 (O_1164,N_19980,N_19957);
xnor UO_1165 (O_1165,N_19873,N_19885);
or UO_1166 (O_1166,N_19903,N_19915);
nand UO_1167 (O_1167,N_19848,N_19923);
or UO_1168 (O_1168,N_19889,N_19943);
xor UO_1169 (O_1169,N_19924,N_19845);
nor UO_1170 (O_1170,N_19882,N_19873);
nor UO_1171 (O_1171,N_19960,N_19982);
and UO_1172 (O_1172,N_19931,N_19859);
nand UO_1173 (O_1173,N_19880,N_19866);
nor UO_1174 (O_1174,N_19846,N_19919);
or UO_1175 (O_1175,N_19930,N_19932);
nand UO_1176 (O_1176,N_19976,N_19843);
or UO_1177 (O_1177,N_19965,N_19936);
xor UO_1178 (O_1178,N_19878,N_19904);
nand UO_1179 (O_1179,N_19844,N_19977);
and UO_1180 (O_1180,N_19904,N_19927);
nand UO_1181 (O_1181,N_19894,N_19993);
and UO_1182 (O_1182,N_19880,N_19938);
and UO_1183 (O_1183,N_19992,N_19840);
and UO_1184 (O_1184,N_19847,N_19979);
xor UO_1185 (O_1185,N_19912,N_19858);
nand UO_1186 (O_1186,N_19875,N_19902);
nand UO_1187 (O_1187,N_19928,N_19951);
xnor UO_1188 (O_1188,N_19938,N_19914);
nand UO_1189 (O_1189,N_19947,N_19986);
xor UO_1190 (O_1190,N_19965,N_19893);
and UO_1191 (O_1191,N_19969,N_19988);
nand UO_1192 (O_1192,N_19876,N_19959);
nand UO_1193 (O_1193,N_19927,N_19975);
nor UO_1194 (O_1194,N_19998,N_19883);
and UO_1195 (O_1195,N_19849,N_19932);
xnor UO_1196 (O_1196,N_19994,N_19967);
nand UO_1197 (O_1197,N_19904,N_19972);
or UO_1198 (O_1198,N_19896,N_19910);
or UO_1199 (O_1199,N_19946,N_19887);
nor UO_1200 (O_1200,N_19993,N_19933);
nand UO_1201 (O_1201,N_19893,N_19862);
and UO_1202 (O_1202,N_19916,N_19850);
nand UO_1203 (O_1203,N_19918,N_19896);
or UO_1204 (O_1204,N_19863,N_19872);
or UO_1205 (O_1205,N_19891,N_19842);
xor UO_1206 (O_1206,N_19866,N_19942);
nand UO_1207 (O_1207,N_19983,N_19976);
or UO_1208 (O_1208,N_19873,N_19946);
nor UO_1209 (O_1209,N_19911,N_19877);
nand UO_1210 (O_1210,N_19860,N_19855);
xnor UO_1211 (O_1211,N_19930,N_19866);
or UO_1212 (O_1212,N_19966,N_19875);
nor UO_1213 (O_1213,N_19908,N_19911);
and UO_1214 (O_1214,N_19870,N_19889);
xor UO_1215 (O_1215,N_19941,N_19923);
xor UO_1216 (O_1216,N_19903,N_19870);
and UO_1217 (O_1217,N_19999,N_19937);
or UO_1218 (O_1218,N_19841,N_19912);
xnor UO_1219 (O_1219,N_19857,N_19885);
nor UO_1220 (O_1220,N_19937,N_19843);
nand UO_1221 (O_1221,N_19855,N_19904);
or UO_1222 (O_1222,N_19918,N_19955);
nor UO_1223 (O_1223,N_19859,N_19953);
xnor UO_1224 (O_1224,N_19910,N_19912);
and UO_1225 (O_1225,N_19914,N_19924);
and UO_1226 (O_1226,N_19938,N_19845);
and UO_1227 (O_1227,N_19976,N_19878);
nand UO_1228 (O_1228,N_19870,N_19923);
xor UO_1229 (O_1229,N_19921,N_19944);
nor UO_1230 (O_1230,N_19909,N_19931);
nand UO_1231 (O_1231,N_19849,N_19917);
nor UO_1232 (O_1232,N_19936,N_19980);
nand UO_1233 (O_1233,N_19840,N_19980);
nor UO_1234 (O_1234,N_19850,N_19952);
or UO_1235 (O_1235,N_19896,N_19848);
and UO_1236 (O_1236,N_19996,N_19983);
and UO_1237 (O_1237,N_19989,N_19992);
or UO_1238 (O_1238,N_19966,N_19968);
xor UO_1239 (O_1239,N_19870,N_19851);
and UO_1240 (O_1240,N_19868,N_19928);
or UO_1241 (O_1241,N_19994,N_19968);
or UO_1242 (O_1242,N_19842,N_19872);
nand UO_1243 (O_1243,N_19895,N_19960);
xor UO_1244 (O_1244,N_19923,N_19967);
nor UO_1245 (O_1245,N_19983,N_19990);
xnor UO_1246 (O_1246,N_19990,N_19905);
nand UO_1247 (O_1247,N_19909,N_19848);
or UO_1248 (O_1248,N_19853,N_19856);
and UO_1249 (O_1249,N_19874,N_19855);
nand UO_1250 (O_1250,N_19997,N_19893);
xnor UO_1251 (O_1251,N_19844,N_19917);
or UO_1252 (O_1252,N_19981,N_19913);
xnor UO_1253 (O_1253,N_19858,N_19986);
nor UO_1254 (O_1254,N_19871,N_19928);
or UO_1255 (O_1255,N_19866,N_19876);
and UO_1256 (O_1256,N_19874,N_19859);
xnor UO_1257 (O_1257,N_19974,N_19876);
xnor UO_1258 (O_1258,N_19964,N_19937);
nand UO_1259 (O_1259,N_19957,N_19905);
and UO_1260 (O_1260,N_19904,N_19915);
nand UO_1261 (O_1261,N_19932,N_19934);
xor UO_1262 (O_1262,N_19869,N_19863);
xor UO_1263 (O_1263,N_19852,N_19884);
nor UO_1264 (O_1264,N_19898,N_19869);
and UO_1265 (O_1265,N_19973,N_19901);
or UO_1266 (O_1266,N_19992,N_19898);
or UO_1267 (O_1267,N_19983,N_19840);
and UO_1268 (O_1268,N_19881,N_19923);
nor UO_1269 (O_1269,N_19957,N_19910);
xor UO_1270 (O_1270,N_19845,N_19981);
nor UO_1271 (O_1271,N_19930,N_19951);
nor UO_1272 (O_1272,N_19955,N_19875);
nand UO_1273 (O_1273,N_19942,N_19845);
or UO_1274 (O_1274,N_19986,N_19939);
and UO_1275 (O_1275,N_19926,N_19944);
or UO_1276 (O_1276,N_19852,N_19908);
nand UO_1277 (O_1277,N_19880,N_19940);
or UO_1278 (O_1278,N_19993,N_19929);
or UO_1279 (O_1279,N_19875,N_19916);
nor UO_1280 (O_1280,N_19985,N_19892);
nor UO_1281 (O_1281,N_19854,N_19982);
and UO_1282 (O_1282,N_19885,N_19848);
xor UO_1283 (O_1283,N_19983,N_19937);
xor UO_1284 (O_1284,N_19902,N_19995);
or UO_1285 (O_1285,N_19864,N_19982);
and UO_1286 (O_1286,N_19926,N_19982);
xor UO_1287 (O_1287,N_19979,N_19962);
nor UO_1288 (O_1288,N_19928,N_19890);
nand UO_1289 (O_1289,N_19872,N_19985);
xor UO_1290 (O_1290,N_19999,N_19887);
or UO_1291 (O_1291,N_19898,N_19904);
nand UO_1292 (O_1292,N_19942,N_19885);
nand UO_1293 (O_1293,N_19920,N_19932);
xnor UO_1294 (O_1294,N_19857,N_19916);
nand UO_1295 (O_1295,N_19975,N_19845);
xor UO_1296 (O_1296,N_19903,N_19962);
xnor UO_1297 (O_1297,N_19868,N_19951);
nor UO_1298 (O_1298,N_19982,N_19899);
or UO_1299 (O_1299,N_19920,N_19978);
or UO_1300 (O_1300,N_19929,N_19891);
and UO_1301 (O_1301,N_19939,N_19982);
and UO_1302 (O_1302,N_19899,N_19863);
or UO_1303 (O_1303,N_19841,N_19904);
xor UO_1304 (O_1304,N_19908,N_19956);
and UO_1305 (O_1305,N_19884,N_19891);
or UO_1306 (O_1306,N_19952,N_19866);
nand UO_1307 (O_1307,N_19950,N_19971);
nor UO_1308 (O_1308,N_19943,N_19962);
and UO_1309 (O_1309,N_19945,N_19911);
and UO_1310 (O_1310,N_19980,N_19982);
or UO_1311 (O_1311,N_19987,N_19993);
nand UO_1312 (O_1312,N_19956,N_19979);
nor UO_1313 (O_1313,N_19985,N_19928);
or UO_1314 (O_1314,N_19866,N_19867);
or UO_1315 (O_1315,N_19869,N_19855);
nand UO_1316 (O_1316,N_19877,N_19881);
or UO_1317 (O_1317,N_19847,N_19945);
nand UO_1318 (O_1318,N_19909,N_19992);
nor UO_1319 (O_1319,N_19924,N_19937);
nand UO_1320 (O_1320,N_19989,N_19844);
or UO_1321 (O_1321,N_19909,N_19892);
nor UO_1322 (O_1322,N_19981,N_19921);
nand UO_1323 (O_1323,N_19959,N_19885);
xor UO_1324 (O_1324,N_19941,N_19857);
xor UO_1325 (O_1325,N_19863,N_19965);
nor UO_1326 (O_1326,N_19899,N_19990);
and UO_1327 (O_1327,N_19911,N_19899);
and UO_1328 (O_1328,N_19999,N_19880);
nor UO_1329 (O_1329,N_19865,N_19897);
or UO_1330 (O_1330,N_19919,N_19845);
and UO_1331 (O_1331,N_19922,N_19968);
xor UO_1332 (O_1332,N_19962,N_19840);
or UO_1333 (O_1333,N_19989,N_19936);
and UO_1334 (O_1334,N_19845,N_19862);
nand UO_1335 (O_1335,N_19939,N_19901);
nor UO_1336 (O_1336,N_19960,N_19920);
nand UO_1337 (O_1337,N_19958,N_19933);
nand UO_1338 (O_1338,N_19973,N_19946);
xnor UO_1339 (O_1339,N_19840,N_19978);
nor UO_1340 (O_1340,N_19937,N_19972);
nand UO_1341 (O_1341,N_19911,N_19864);
nand UO_1342 (O_1342,N_19840,N_19948);
nand UO_1343 (O_1343,N_19864,N_19914);
or UO_1344 (O_1344,N_19941,N_19983);
nor UO_1345 (O_1345,N_19865,N_19900);
and UO_1346 (O_1346,N_19912,N_19947);
nor UO_1347 (O_1347,N_19992,N_19962);
nor UO_1348 (O_1348,N_19937,N_19988);
nand UO_1349 (O_1349,N_19993,N_19988);
nor UO_1350 (O_1350,N_19847,N_19927);
xor UO_1351 (O_1351,N_19917,N_19936);
and UO_1352 (O_1352,N_19942,N_19940);
nor UO_1353 (O_1353,N_19995,N_19938);
nor UO_1354 (O_1354,N_19940,N_19902);
nor UO_1355 (O_1355,N_19944,N_19965);
nor UO_1356 (O_1356,N_19899,N_19965);
nor UO_1357 (O_1357,N_19843,N_19847);
or UO_1358 (O_1358,N_19925,N_19907);
and UO_1359 (O_1359,N_19975,N_19859);
or UO_1360 (O_1360,N_19948,N_19959);
or UO_1361 (O_1361,N_19898,N_19948);
and UO_1362 (O_1362,N_19914,N_19998);
nor UO_1363 (O_1363,N_19920,N_19857);
and UO_1364 (O_1364,N_19968,N_19928);
or UO_1365 (O_1365,N_19862,N_19946);
xor UO_1366 (O_1366,N_19999,N_19879);
nand UO_1367 (O_1367,N_19989,N_19962);
xor UO_1368 (O_1368,N_19984,N_19909);
or UO_1369 (O_1369,N_19974,N_19875);
nor UO_1370 (O_1370,N_19846,N_19917);
and UO_1371 (O_1371,N_19886,N_19914);
xnor UO_1372 (O_1372,N_19993,N_19849);
nor UO_1373 (O_1373,N_19964,N_19955);
xor UO_1374 (O_1374,N_19846,N_19862);
nand UO_1375 (O_1375,N_19937,N_19951);
or UO_1376 (O_1376,N_19914,N_19860);
and UO_1377 (O_1377,N_19845,N_19927);
nand UO_1378 (O_1378,N_19850,N_19936);
nor UO_1379 (O_1379,N_19904,N_19970);
or UO_1380 (O_1380,N_19956,N_19948);
nand UO_1381 (O_1381,N_19911,N_19965);
xor UO_1382 (O_1382,N_19947,N_19871);
xnor UO_1383 (O_1383,N_19896,N_19863);
xnor UO_1384 (O_1384,N_19862,N_19943);
xnor UO_1385 (O_1385,N_19880,N_19972);
and UO_1386 (O_1386,N_19857,N_19964);
and UO_1387 (O_1387,N_19991,N_19888);
nor UO_1388 (O_1388,N_19922,N_19846);
nor UO_1389 (O_1389,N_19886,N_19976);
or UO_1390 (O_1390,N_19975,N_19896);
nor UO_1391 (O_1391,N_19961,N_19999);
nand UO_1392 (O_1392,N_19931,N_19948);
xor UO_1393 (O_1393,N_19981,N_19984);
or UO_1394 (O_1394,N_19869,N_19850);
xnor UO_1395 (O_1395,N_19870,N_19944);
nand UO_1396 (O_1396,N_19936,N_19856);
xor UO_1397 (O_1397,N_19866,N_19974);
xor UO_1398 (O_1398,N_19953,N_19916);
or UO_1399 (O_1399,N_19967,N_19939);
xnor UO_1400 (O_1400,N_19926,N_19975);
xor UO_1401 (O_1401,N_19924,N_19875);
nor UO_1402 (O_1402,N_19958,N_19941);
nor UO_1403 (O_1403,N_19876,N_19911);
xnor UO_1404 (O_1404,N_19922,N_19967);
nor UO_1405 (O_1405,N_19991,N_19923);
nand UO_1406 (O_1406,N_19867,N_19940);
and UO_1407 (O_1407,N_19909,N_19948);
or UO_1408 (O_1408,N_19997,N_19925);
xor UO_1409 (O_1409,N_19894,N_19899);
or UO_1410 (O_1410,N_19922,N_19934);
nor UO_1411 (O_1411,N_19886,N_19994);
and UO_1412 (O_1412,N_19925,N_19986);
nand UO_1413 (O_1413,N_19863,N_19909);
or UO_1414 (O_1414,N_19955,N_19905);
and UO_1415 (O_1415,N_19978,N_19905);
or UO_1416 (O_1416,N_19962,N_19928);
or UO_1417 (O_1417,N_19841,N_19984);
or UO_1418 (O_1418,N_19873,N_19994);
or UO_1419 (O_1419,N_19945,N_19841);
and UO_1420 (O_1420,N_19975,N_19942);
xor UO_1421 (O_1421,N_19938,N_19901);
nand UO_1422 (O_1422,N_19959,N_19880);
nand UO_1423 (O_1423,N_19868,N_19927);
or UO_1424 (O_1424,N_19896,N_19959);
xor UO_1425 (O_1425,N_19979,N_19959);
and UO_1426 (O_1426,N_19870,N_19895);
or UO_1427 (O_1427,N_19882,N_19982);
nor UO_1428 (O_1428,N_19909,N_19918);
xor UO_1429 (O_1429,N_19875,N_19972);
and UO_1430 (O_1430,N_19848,N_19998);
xor UO_1431 (O_1431,N_19965,N_19931);
nor UO_1432 (O_1432,N_19882,N_19959);
nor UO_1433 (O_1433,N_19847,N_19936);
or UO_1434 (O_1434,N_19894,N_19896);
nand UO_1435 (O_1435,N_19950,N_19909);
nor UO_1436 (O_1436,N_19900,N_19897);
and UO_1437 (O_1437,N_19930,N_19899);
xor UO_1438 (O_1438,N_19842,N_19951);
nand UO_1439 (O_1439,N_19899,N_19989);
and UO_1440 (O_1440,N_19942,N_19864);
nor UO_1441 (O_1441,N_19934,N_19927);
nand UO_1442 (O_1442,N_19840,N_19888);
and UO_1443 (O_1443,N_19983,N_19899);
nor UO_1444 (O_1444,N_19976,N_19907);
xnor UO_1445 (O_1445,N_19977,N_19950);
nor UO_1446 (O_1446,N_19951,N_19986);
nor UO_1447 (O_1447,N_19863,N_19993);
xnor UO_1448 (O_1448,N_19850,N_19856);
xnor UO_1449 (O_1449,N_19949,N_19914);
nand UO_1450 (O_1450,N_19982,N_19984);
or UO_1451 (O_1451,N_19876,N_19854);
xor UO_1452 (O_1452,N_19902,N_19933);
or UO_1453 (O_1453,N_19872,N_19859);
or UO_1454 (O_1454,N_19840,N_19959);
or UO_1455 (O_1455,N_19907,N_19909);
xnor UO_1456 (O_1456,N_19972,N_19883);
or UO_1457 (O_1457,N_19913,N_19979);
nor UO_1458 (O_1458,N_19885,N_19979);
or UO_1459 (O_1459,N_19897,N_19884);
and UO_1460 (O_1460,N_19975,N_19969);
or UO_1461 (O_1461,N_19872,N_19982);
or UO_1462 (O_1462,N_19942,N_19920);
nand UO_1463 (O_1463,N_19876,N_19917);
nand UO_1464 (O_1464,N_19978,N_19939);
xor UO_1465 (O_1465,N_19903,N_19892);
or UO_1466 (O_1466,N_19840,N_19859);
nor UO_1467 (O_1467,N_19846,N_19869);
xor UO_1468 (O_1468,N_19997,N_19995);
nor UO_1469 (O_1469,N_19996,N_19863);
and UO_1470 (O_1470,N_19854,N_19852);
and UO_1471 (O_1471,N_19957,N_19997);
nand UO_1472 (O_1472,N_19887,N_19995);
nor UO_1473 (O_1473,N_19993,N_19971);
nand UO_1474 (O_1474,N_19842,N_19850);
or UO_1475 (O_1475,N_19998,N_19973);
nor UO_1476 (O_1476,N_19977,N_19842);
nor UO_1477 (O_1477,N_19891,N_19895);
xnor UO_1478 (O_1478,N_19915,N_19845);
nor UO_1479 (O_1479,N_19874,N_19915);
and UO_1480 (O_1480,N_19869,N_19871);
xnor UO_1481 (O_1481,N_19968,N_19918);
and UO_1482 (O_1482,N_19864,N_19857);
and UO_1483 (O_1483,N_19924,N_19843);
and UO_1484 (O_1484,N_19891,N_19921);
or UO_1485 (O_1485,N_19924,N_19900);
nor UO_1486 (O_1486,N_19968,N_19974);
nand UO_1487 (O_1487,N_19884,N_19929);
or UO_1488 (O_1488,N_19976,N_19901);
and UO_1489 (O_1489,N_19863,N_19907);
xnor UO_1490 (O_1490,N_19997,N_19871);
nor UO_1491 (O_1491,N_19960,N_19992);
and UO_1492 (O_1492,N_19970,N_19999);
xnor UO_1493 (O_1493,N_19847,N_19844);
and UO_1494 (O_1494,N_19983,N_19946);
and UO_1495 (O_1495,N_19871,N_19904);
or UO_1496 (O_1496,N_19881,N_19942);
nor UO_1497 (O_1497,N_19989,N_19934);
or UO_1498 (O_1498,N_19942,N_19879);
nor UO_1499 (O_1499,N_19901,N_19949);
nor UO_1500 (O_1500,N_19987,N_19968);
or UO_1501 (O_1501,N_19948,N_19908);
or UO_1502 (O_1502,N_19840,N_19854);
nand UO_1503 (O_1503,N_19847,N_19937);
nor UO_1504 (O_1504,N_19929,N_19850);
nor UO_1505 (O_1505,N_19916,N_19865);
and UO_1506 (O_1506,N_19922,N_19860);
and UO_1507 (O_1507,N_19880,N_19914);
nand UO_1508 (O_1508,N_19949,N_19854);
and UO_1509 (O_1509,N_19951,N_19861);
and UO_1510 (O_1510,N_19893,N_19938);
xor UO_1511 (O_1511,N_19919,N_19931);
and UO_1512 (O_1512,N_19980,N_19862);
or UO_1513 (O_1513,N_19933,N_19906);
nand UO_1514 (O_1514,N_19898,N_19853);
nor UO_1515 (O_1515,N_19872,N_19852);
and UO_1516 (O_1516,N_19935,N_19930);
nand UO_1517 (O_1517,N_19921,N_19959);
nor UO_1518 (O_1518,N_19860,N_19985);
nor UO_1519 (O_1519,N_19976,N_19938);
or UO_1520 (O_1520,N_19955,N_19914);
or UO_1521 (O_1521,N_19925,N_19874);
xnor UO_1522 (O_1522,N_19867,N_19875);
nand UO_1523 (O_1523,N_19895,N_19915);
xor UO_1524 (O_1524,N_19917,N_19977);
xor UO_1525 (O_1525,N_19962,N_19984);
or UO_1526 (O_1526,N_19954,N_19892);
or UO_1527 (O_1527,N_19917,N_19990);
or UO_1528 (O_1528,N_19953,N_19937);
xor UO_1529 (O_1529,N_19957,N_19871);
nand UO_1530 (O_1530,N_19880,N_19858);
xor UO_1531 (O_1531,N_19994,N_19957);
or UO_1532 (O_1532,N_19927,N_19843);
and UO_1533 (O_1533,N_19896,N_19888);
or UO_1534 (O_1534,N_19968,N_19908);
xnor UO_1535 (O_1535,N_19944,N_19866);
nor UO_1536 (O_1536,N_19953,N_19981);
nand UO_1537 (O_1537,N_19918,N_19911);
nand UO_1538 (O_1538,N_19880,N_19991);
xnor UO_1539 (O_1539,N_19960,N_19954);
or UO_1540 (O_1540,N_19958,N_19924);
and UO_1541 (O_1541,N_19860,N_19998);
xor UO_1542 (O_1542,N_19891,N_19983);
xor UO_1543 (O_1543,N_19979,N_19986);
nand UO_1544 (O_1544,N_19907,N_19980);
xor UO_1545 (O_1545,N_19865,N_19980);
nor UO_1546 (O_1546,N_19937,N_19995);
nand UO_1547 (O_1547,N_19953,N_19840);
nor UO_1548 (O_1548,N_19998,N_19903);
or UO_1549 (O_1549,N_19888,N_19996);
or UO_1550 (O_1550,N_19899,N_19929);
and UO_1551 (O_1551,N_19907,N_19972);
or UO_1552 (O_1552,N_19988,N_19972);
or UO_1553 (O_1553,N_19907,N_19913);
or UO_1554 (O_1554,N_19887,N_19908);
nor UO_1555 (O_1555,N_19847,N_19975);
nor UO_1556 (O_1556,N_19934,N_19882);
and UO_1557 (O_1557,N_19902,N_19840);
or UO_1558 (O_1558,N_19937,N_19916);
or UO_1559 (O_1559,N_19942,N_19948);
xor UO_1560 (O_1560,N_19998,N_19904);
nor UO_1561 (O_1561,N_19940,N_19910);
or UO_1562 (O_1562,N_19861,N_19869);
or UO_1563 (O_1563,N_19852,N_19956);
xnor UO_1564 (O_1564,N_19983,N_19999);
or UO_1565 (O_1565,N_19950,N_19855);
nand UO_1566 (O_1566,N_19920,N_19900);
nor UO_1567 (O_1567,N_19884,N_19967);
xnor UO_1568 (O_1568,N_19910,N_19874);
or UO_1569 (O_1569,N_19914,N_19916);
and UO_1570 (O_1570,N_19919,N_19882);
xnor UO_1571 (O_1571,N_19847,N_19968);
or UO_1572 (O_1572,N_19940,N_19893);
and UO_1573 (O_1573,N_19899,N_19883);
and UO_1574 (O_1574,N_19883,N_19851);
nand UO_1575 (O_1575,N_19877,N_19841);
and UO_1576 (O_1576,N_19975,N_19909);
or UO_1577 (O_1577,N_19928,N_19902);
or UO_1578 (O_1578,N_19924,N_19848);
nor UO_1579 (O_1579,N_19913,N_19988);
nor UO_1580 (O_1580,N_19903,N_19986);
nor UO_1581 (O_1581,N_19863,N_19845);
xor UO_1582 (O_1582,N_19884,N_19904);
xor UO_1583 (O_1583,N_19962,N_19905);
and UO_1584 (O_1584,N_19919,N_19963);
and UO_1585 (O_1585,N_19896,N_19924);
xnor UO_1586 (O_1586,N_19953,N_19864);
nor UO_1587 (O_1587,N_19911,N_19914);
nand UO_1588 (O_1588,N_19906,N_19904);
nor UO_1589 (O_1589,N_19979,N_19881);
or UO_1590 (O_1590,N_19852,N_19894);
nor UO_1591 (O_1591,N_19963,N_19908);
xor UO_1592 (O_1592,N_19970,N_19890);
nand UO_1593 (O_1593,N_19980,N_19913);
or UO_1594 (O_1594,N_19892,N_19973);
nor UO_1595 (O_1595,N_19937,N_19996);
and UO_1596 (O_1596,N_19971,N_19964);
or UO_1597 (O_1597,N_19917,N_19997);
nor UO_1598 (O_1598,N_19884,N_19944);
and UO_1599 (O_1599,N_19923,N_19889);
nand UO_1600 (O_1600,N_19999,N_19956);
and UO_1601 (O_1601,N_19961,N_19875);
nor UO_1602 (O_1602,N_19876,N_19908);
xnor UO_1603 (O_1603,N_19998,N_19905);
nor UO_1604 (O_1604,N_19878,N_19915);
nor UO_1605 (O_1605,N_19911,N_19975);
nor UO_1606 (O_1606,N_19996,N_19947);
and UO_1607 (O_1607,N_19858,N_19915);
xnor UO_1608 (O_1608,N_19999,N_19844);
nor UO_1609 (O_1609,N_19899,N_19907);
or UO_1610 (O_1610,N_19955,N_19973);
or UO_1611 (O_1611,N_19934,N_19872);
xnor UO_1612 (O_1612,N_19870,N_19939);
nor UO_1613 (O_1613,N_19928,N_19905);
and UO_1614 (O_1614,N_19977,N_19860);
nor UO_1615 (O_1615,N_19981,N_19950);
xnor UO_1616 (O_1616,N_19934,N_19948);
and UO_1617 (O_1617,N_19996,N_19965);
xor UO_1618 (O_1618,N_19907,N_19885);
xnor UO_1619 (O_1619,N_19959,N_19848);
nor UO_1620 (O_1620,N_19986,N_19975);
nor UO_1621 (O_1621,N_19871,N_19943);
or UO_1622 (O_1622,N_19870,N_19956);
nand UO_1623 (O_1623,N_19907,N_19843);
nor UO_1624 (O_1624,N_19879,N_19969);
or UO_1625 (O_1625,N_19871,N_19960);
nor UO_1626 (O_1626,N_19979,N_19957);
and UO_1627 (O_1627,N_19872,N_19909);
or UO_1628 (O_1628,N_19867,N_19957);
nor UO_1629 (O_1629,N_19923,N_19944);
or UO_1630 (O_1630,N_19844,N_19923);
or UO_1631 (O_1631,N_19905,N_19866);
nor UO_1632 (O_1632,N_19895,N_19930);
nor UO_1633 (O_1633,N_19867,N_19921);
nand UO_1634 (O_1634,N_19919,N_19938);
xnor UO_1635 (O_1635,N_19961,N_19896);
nand UO_1636 (O_1636,N_19847,N_19969);
nand UO_1637 (O_1637,N_19931,N_19992);
or UO_1638 (O_1638,N_19994,N_19940);
xor UO_1639 (O_1639,N_19844,N_19943);
nand UO_1640 (O_1640,N_19902,N_19895);
nor UO_1641 (O_1641,N_19917,N_19887);
or UO_1642 (O_1642,N_19932,N_19933);
and UO_1643 (O_1643,N_19996,N_19865);
or UO_1644 (O_1644,N_19855,N_19974);
nand UO_1645 (O_1645,N_19916,N_19934);
nor UO_1646 (O_1646,N_19984,N_19953);
nand UO_1647 (O_1647,N_19855,N_19854);
or UO_1648 (O_1648,N_19903,N_19891);
xor UO_1649 (O_1649,N_19840,N_19856);
and UO_1650 (O_1650,N_19985,N_19866);
nor UO_1651 (O_1651,N_19935,N_19919);
xor UO_1652 (O_1652,N_19889,N_19849);
or UO_1653 (O_1653,N_19959,N_19873);
or UO_1654 (O_1654,N_19980,N_19941);
nor UO_1655 (O_1655,N_19844,N_19978);
and UO_1656 (O_1656,N_19884,N_19892);
xnor UO_1657 (O_1657,N_19845,N_19980);
and UO_1658 (O_1658,N_19849,N_19985);
nor UO_1659 (O_1659,N_19980,N_19893);
nand UO_1660 (O_1660,N_19939,N_19883);
nor UO_1661 (O_1661,N_19858,N_19994);
nand UO_1662 (O_1662,N_19870,N_19885);
xnor UO_1663 (O_1663,N_19990,N_19926);
nand UO_1664 (O_1664,N_19866,N_19856);
and UO_1665 (O_1665,N_19861,N_19946);
and UO_1666 (O_1666,N_19862,N_19850);
nor UO_1667 (O_1667,N_19959,N_19928);
or UO_1668 (O_1668,N_19881,N_19928);
nand UO_1669 (O_1669,N_19866,N_19872);
or UO_1670 (O_1670,N_19942,N_19884);
and UO_1671 (O_1671,N_19863,N_19902);
or UO_1672 (O_1672,N_19890,N_19910);
xor UO_1673 (O_1673,N_19875,N_19841);
and UO_1674 (O_1674,N_19955,N_19933);
and UO_1675 (O_1675,N_19892,N_19928);
and UO_1676 (O_1676,N_19850,N_19870);
or UO_1677 (O_1677,N_19964,N_19912);
nor UO_1678 (O_1678,N_19906,N_19947);
nand UO_1679 (O_1679,N_19939,N_19945);
or UO_1680 (O_1680,N_19926,N_19878);
and UO_1681 (O_1681,N_19999,N_19989);
nand UO_1682 (O_1682,N_19866,N_19843);
xnor UO_1683 (O_1683,N_19986,N_19856);
nand UO_1684 (O_1684,N_19945,N_19916);
and UO_1685 (O_1685,N_19881,N_19866);
xor UO_1686 (O_1686,N_19929,N_19920);
and UO_1687 (O_1687,N_19849,N_19893);
nor UO_1688 (O_1688,N_19962,N_19915);
nor UO_1689 (O_1689,N_19895,N_19910);
nor UO_1690 (O_1690,N_19889,N_19951);
nor UO_1691 (O_1691,N_19880,N_19903);
nand UO_1692 (O_1692,N_19976,N_19852);
xnor UO_1693 (O_1693,N_19856,N_19908);
and UO_1694 (O_1694,N_19944,N_19992);
or UO_1695 (O_1695,N_19889,N_19852);
and UO_1696 (O_1696,N_19848,N_19863);
nand UO_1697 (O_1697,N_19997,N_19897);
and UO_1698 (O_1698,N_19844,N_19919);
xor UO_1699 (O_1699,N_19862,N_19907);
or UO_1700 (O_1700,N_19897,N_19996);
nor UO_1701 (O_1701,N_19928,N_19992);
nor UO_1702 (O_1702,N_19864,N_19885);
or UO_1703 (O_1703,N_19874,N_19966);
xor UO_1704 (O_1704,N_19877,N_19908);
or UO_1705 (O_1705,N_19975,N_19935);
nor UO_1706 (O_1706,N_19955,N_19854);
and UO_1707 (O_1707,N_19928,N_19861);
and UO_1708 (O_1708,N_19992,N_19956);
nand UO_1709 (O_1709,N_19932,N_19974);
nand UO_1710 (O_1710,N_19856,N_19883);
nor UO_1711 (O_1711,N_19994,N_19915);
nand UO_1712 (O_1712,N_19996,N_19972);
xnor UO_1713 (O_1713,N_19854,N_19945);
nand UO_1714 (O_1714,N_19882,N_19979);
nor UO_1715 (O_1715,N_19890,N_19867);
nand UO_1716 (O_1716,N_19960,N_19876);
nor UO_1717 (O_1717,N_19876,N_19898);
xor UO_1718 (O_1718,N_19976,N_19899);
xnor UO_1719 (O_1719,N_19841,N_19997);
xnor UO_1720 (O_1720,N_19889,N_19890);
xor UO_1721 (O_1721,N_19865,N_19905);
nand UO_1722 (O_1722,N_19951,N_19952);
nand UO_1723 (O_1723,N_19993,N_19852);
xnor UO_1724 (O_1724,N_19954,N_19945);
xnor UO_1725 (O_1725,N_19871,N_19868);
or UO_1726 (O_1726,N_19917,N_19939);
or UO_1727 (O_1727,N_19895,N_19859);
nand UO_1728 (O_1728,N_19855,N_19988);
and UO_1729 (O_1729,N_19980,N_19938);
nand UO_1730 (O_1730,N_19904,N_19926);
and UO_1731 (O_1731,N_19876,N_19975);
nor UO_1732 (O_1732,N_19840,N_19914);
nand UO_1733 (O_1733,N_19858,N_19917);
or UO_1734 (O_1734,N_19986,N_19904);
or UO_1735 (O_1735,N_19854,N_19967);
and UO_1736 (O_1736,N_19997,N_19990);
or UO_1737 (O_1737,N_19981,N_19902);
nor UO_1738 (O_1738,N_19899,N_19897);
nand UO_1739 (O_1739,N_19999,N_19918);
and UO_1740 (O_1740,N_19894,N_19855);
xnor UO_1741 (O_1741,N_19874,N_19950);
or UO_1742 (O_1742,N_19855,N_19944);
nor UO_1743 (O_1743,N_19924,N_19941);
and UO_1744 (O_1744,N_19981,N_19843);
xor UO_1745 (O_1745,N_19884,N_19845);
nor UO_1746 (O_1746,N_19902,N_19973);
and UO_1747 (O_1747,N_19896,N_19967);
nor UO_1748 (O_1748,N_19887,N_19985);
or UO_1749 (O_1749,N_19969,N_19856);
nor UO_1750 (O_1750,N_19980,N_19959);
xor UO_1751 (O_1751,N_19984,N_19908);
nand UO_1752 (O_1752,N_19882,N_19858);
xnor UO_1753 (O_1753,N_19985,N_19862);
nor UO_1754 (O_1754,N_19869,N_19999);
or UO_1755 (O_1755,N_19897,N_19915);
or UO_1756 (O_1756,N_19937,N_19948);
and UO_1757 (O_1757,N_19957,N_19909);
or UO_1758 (O_1758,N_19995,N_19898);
nand UO_1759 (O_1759,N_19907,N_19870);
nand UO_1760 (O_1760,N_19901,N_19930);
nand UO_1761 (O_1761,N_19972,N_19942);
xnor UO_1762 (O_1762,N_19997,N_19882);
nor UO_1763 (O_1763,N_19910,N_19850);
xnor UO_1764 (O_1764,N_19996,N_19846);
nand UO_1765 (O_1765,N_19860,N_19863);
nor UO_1766 (O_1766,N_19884,N_19925);
or UO_1767 (O_1767,N_19890,N_19892);
or UO_1768 (O_1768,N_19851,N_19922);
and UO_1769 (O_1769,N_19885,N_19896);
xor UO_1770 (O_1770,N_19905,N_19904);
xnor UO_1771 (O_1771,N_19878,N_19905);
nand UO_1772 (O_1772,N_19859,N_19881);
nand UO_1773 (O_1773,N_19878,N_19931);
nor UO_1774 (O_1774,N_19948,N_19952);
or UO_1775 (O_1775,N_19867,N_19894);
nor UO_1776 (O_1776,N_19899,N_19850);
nor UO_1777 (O_1777,N_19974,N_19996);
xor UO_1778 (O_1778,N_19886,N_19961);
nand UO_1779 (O_1779,N_19924,N_19849);
nor UO_1780 (O_1780,N_19874,N_19980);
and UO_1781 (O_1781,N_19863,N_19959);
nand UO_1782 (O_1782,N_19941,N_19935);
nand UO_1783 (O_1783,N_19925,N_19846);
nand UO_1784 (O_1784,N_19993,N_19842);
nand UO_1785 (O_1785,N_19953,N_19908);
xnor UO_1786 (O_1786,N_19957,N_19963);
nor UO_1787 (O_1787,N_19847,N_19941);
or UO_1788 (O_1788,N_19868,N_19919);
nor UO_1789 (O_1789,N_19942,N_19973);
nor UO_1790 (O_1790,N_19941,N_19840);
or UO_1791 (O_1791,N_19862,N_19981);
nand UO_1792 (O_1792,N_19925,N_19902);
nand UO_1793 (O_1793,N_19960,N_19987);
nor UO_1794 (O_1794,N_19871,N_19841);
nor UO_1795 (O_1795,N_19876,N_19957);
or UO_1796 (O_1796,N_19929,N_19868);
xor UO_1797 (O_1797,N_19989,N_19970);
and UO_1798 (O_1798,N_19961,N_19898);
nand UO_1799 (O_1799,N_19959,N_19934);
and UO_1800 (O_1800,N_19993,N_19973);
nand UO_1801 (O_1801,N_19901,N_19908);
xnor UO_1802 (O_1802,N_19928,N_19979);
xor UO_1803 (O_1803,N_19869,N_19977);
or UO_1804 (O_1804,N_19905,N_19922);
and UO_1805 (O_1805,N_19945,N_19935);
xnor UO_1806 (O_1806,N_19941,N_19944);
and UO_1807 (O_1807,N_19934,N_19840);
and UO_1808 (O_1808,N_19945,N_19981);
nor UO_1809 (O_1809,N_19858,N_19959);
nand UO_1810 (O_1810,N_19853,N_19900);
and UO_1811 (O_1811,N_19974,N_19999);
or UO_1812 (O_1812,N_19921,N_19870);
or UO_1813 (O_1813,N_19971,N_19951);
xnor UO_1814 (O_1814,N_19910,N_19922);
and UO_1815 (O_1815,N_19955,N_19967);
or UO_1816 (O_1816,N_19921,N_19992);
nor UO_1817 (O_1817,N_19862,N_19886);
and UO_1818 (O_1818,N_19843,N_19994);
xnor UO_1819 (O_1819,N_19950,N_19958);
and UO_1820 (O_1820,N_19995,N_19849);
or UO_1821 (O_1821,N_19936,N_19884);
nand UO_1822 (O_1822,N_19906,N_19843);
and UO_1823 (O_1823,N_19905,N_19950);
or UO_1824 (O_1824,N_19961,N_19903);
nor UO_1825 (O_1825,N_19971,N_19906);
xor UO_1826 (O_1826,N_19935,N_19992);
or UO_1827 (O_1827,N_19966,N_19961);
nor UO_1828 (O_1828,N_19870,N_19963);
nand UO_1829 (O_1829,N_19844,N_19933);
or UO_1830 (O_1830,N_19995,N_19900);
and UO_1831 (O_1831,N_19892,N_19924);
nor UO_1832 (O_1832,N_19946,N_19996);
xor UO_1833 (O_1833,N_19858,N_19927);
xor UO_1834 (O_1834,N_19973,N_19890);
or UO_1835 (O_1835,N_19906,N_19853);
xor UO_1836 (O_1836,N_19949,N_19931);
or UO_1837 (O_1837,N_19865,N_19851);
nand UO_1838 (O_1838,N_19919,N_19902);
nand UO_1839 (O_1839,N_19934,N_19981);
xnor UO_1840 (O_1840,N_19980,N_19872);
nand UO_1841 (O_1841,N_19852,N_19942);
nor UO_1842 (O_1842,N_19982,N_19943);
xnor UO_1843 (O_1843,N_19911,N_19969);
xnor UO_1844 (O_1844,N_19971,N_19918);
xor UO_1845 (O_1845,N_19968,N_19914);
and UO_1846 (O_1846,N_19897,N_19991);
nor UO_1847 (O_1847,N_19939,N_19947);
and UO_1848 (O_1848,N_19942,N_19998);
nor UO_1849 (O_1849,N_19923,N_19885);
or UO_1850 (O_1850,N_19948,N_19999);
nor UO_1851 (O_1851,N_19911,N_19952);
nand UO_1852 (O_1852,N_19878,N_19907);
nor UO_1853 (O_1853,N_19873,N_19958);
nor UO_1854 (O_1854,N_19944,N_19969);
nor UO_1855 (O_1855,N_19919,N_19999);
or UO_1856 (O_1856,N_19886,N_19933);
nand UO_1857 (O_1857,N_19858,N_19962);
xor UO_1858 (O_1858,N_19876,N_19982);
and UO_1859 (O_1859,N_19895,N_19852);
xnor UO_1860 (O_1860,N_19977,N_19895);
nand UO_1861 (O_1861,N_19913,N_19903);
xnor UO_1862 (O_1862,N_19937,N_19893);
and UO_1863 (O_1863,N_19952,N_19906);
nor UO_1864 (O_1864,N_19854,N_19867);
or UO_1865 (O_1865,N_19930,N_19919);
nor UO_1866 (O_1866,N_19880,N_19922);
xnor UO_1867 (O_1867,N_19861,N_19911);
and UO_1868 (O_1868,N_19950,N_19919);
nand UO_1869 (O_1869,N_19851,N_19929);
and UO_1870 (O_1870,N_19899,N_19901);
xor UO_1871 (O_1871,N_19980,N_19956);
or UO_1872 (O_1872,N_19953,N_19903);
xnor UO_1873 (O_1873,N_19897,N_19896);
or UO_1874 (O_1874,N_19871,N_19961);
nand UO_1875 (O_1875,N_19982,N_19848);
or UO_1876 (O_1876,N_19977,N_19896);
nor UO_1877 (O_1877,N_19858,N_19875);
nand UO_1878 (O_1878,N_19994,N_19874);
and UO_1879 (O_1879,N_19872,N_19889);
xnor UO_1880 (O_1880,N_19860,N_19976);
nand UO_1881 (O_1881,N_19986,N_19958);
or UO_1882 (O_1882,N_19860,N_19899);
and UO_1883 (O_1883,N_19960,N_19919);
nand UO_1884 (O_1884,N_19898,N_19880);
or UO_1885 (O_1885,N_19862,N_19997);
nand UO_1886 (O_1886,N_19898,N_19997);
or UO_1887 (O_1887,N_19913,N_19879);
and UO_1888 (O_1888,N_19916,N_19983);
xnor UO_1889 (O_1889,N_19847,N_19987);
and UO_1890 (O_1890,N_19960,N_19926);
nor UO_1891 (O_1891,N_19901,N_19912);
and UO_1892 (O_1892,N_19858,N_19862);
and UO_1893 (O_1893,N_19901,N_19943);
or UO_1894 (O_1894,N_19996,N_19871);
or UO_1895 (O_1895,N_19970,N_19902);
or UO_1896 (O_1896,N_19869,N_19990);
nand UO_1897 (O_1897,N_19854,N_19856);
nor UO_1898 (O_1898,N_19887,N_19873);
xor UO_1899 (O_1899,N_19964,N_19920);
or UO_1900 (O_1900,N_19878,N_19954);
xor UO_1901 (O_1901,N_19841,N_19848);
and UO_1902 (O_1902,N_19993,N_19909);
nor UO_1903 (O_1903,N_19900,N_19898);
and UO_1904 (O_1904,N_19975,N_19938);
and UO_1905 (O_1905,N_19971,N_19983);
nand UO_1906 (O_1906,N_19912,N_19894);
nand UO_1907 (O_1907,N_19978,N_19955);
nand UO_1908 (O_1908,N_19867,N_19898);
and UO_1909 (O_1909,N_19985,N_19971);
nand UO_1910 (O_1910,N_19928,N_19994);
nand UO_1911 (O_1911,N_19895,N_19871);
nand UO_1912 (O_1912,N_19930,N_19871);
and UO_1913 (O_1913,N_19978,N_19948);
xor UO_1914 (O_1914,N_19888,N_19850);
and UO_1915 (O_1915,N_19845,N_19982);
or UO_1916 (O_1916,N_19994,N_19889);
or UO_1917 (O_1917,N_19963,N_19985);
nor UO_1918 (O_1918,N_19951,N_19877);
or UO_1919 (O_1919,N_19870,N_19953);
nand UO_1920 (O_1920,N_19961,N_19931);
nor UO_1921 (O_1921,N_19941,N_19878);
xnor UO_1922 (O_1922,N_19938,N_19945);
nand UO_1923 (O_1923,N_19870,N_19849);
or UO_1924 (O_1924,N_19894,N_19877);
xnor UO_1925 (O_1925,N_19976,N_19882);
and UO_1926 (O_1926,N_19942,N_19872);
or UO_1927 (O_1927,N_19995,N_19930);
or UO_1928 (O_1928,N_19860,N_19972);
xor UO_1929 (O_1929,N_19943,N_19958);
or UO_1930 (O_1930,N_19881,N_19944);
or UO_1931 (O_1931,N_19911,N_19862);
xor UO_1932 (O_1932,N_19987,N_19974);
and UO_1933 (O_1933,N_19923,N_19903);
nand UO_1934 (O_1934,N_19840,N_19951);
or UO_1935 (O_1935,N_19889,N_19846);
nor UO_1936 (O_1936,N_19989,N_19906);
or UO_1937 (O_1937,N_19900,N_19952);
xor UO_1938 (O_1938,N_19908,N_19969);
xor UO_1939 (O_1939,N_19854,N_19927);
nand UO_1940 (O_1940,N_19976,N_19942);
nor UO_1941 (O_1941,N_19959,N_19912);
or UO_1942 (O_1942,N_19863,N_19849);
or UO_1943 (O_1943,N_19964,N_19938);
nor UO_1944 (O_1944,N_19983,N_19848);
nand UO_1945 (O_1945,N_19859,N_19910);
and UO_1946 (O_1946,N_19971,N_19855);
and UO_1947 (O_1947,N_19961,N_19927);
xnor UO_1948 (O_1948,N_19880,N_19872);
or UO_1949 (O_1949,N_19932,N_19885);
and UO_1950 (O_1950,N_19973,N_19918);
xnor UO_1951 (O_1951,N_19949,N_19865);
or UO_1952 (O_1952,N_19900,N_19909);
nand UO_1953 (O_1953,N_19880,N_19984);
xor UO_1954 (O_1954,N_19848,N_19846);
nor UO_1955 (O_1955,N_19852,N_19878);
nor UO_1956 (O_1956,N_19883,N_19857);
nor UO_1957 (O_1957,N_19945,N_19999);
nand UO_1958 (O_1958,N_19963,N_19864);
and UO_1959 (O_1959,N_19863,N_19891);
nor UO_1960 (O_1960,N_19872,N_19841);
and UO_1961 (O_1961,N_19864,N_19845);
and UO_1962 (O_1962,N_19965,N_19921);
xor UO_1963 (O_1963,N_19996,N_19893);
or UO_1964 (O_1964,N_19957,N_19845);
nor UO_1965 (O_1965,N_19884,N_19961);
nand UO_1966 (O_1966,N_19847,N_19940);
and UO_1967 (O_1967,N_19915,N_19883);
nand UO_1968 (O_1968,N_19922,N_19885);
xnor UO_1969 (O_1969,N_19938,N_19872);
nand UO_1970 (O_1970,N_19997,N_19979);
nor UO_1971 (O_1971,N_19863,N_19999);
xor UO_1972 (O_1972,N_19872,N_19879);
nor UO_1973 (O_1973,N_19877,N_19861);
or UO_1974 (O_1974,N_19926,N_19971);
or UO_1975 (O_1975,N_19994,N_19853);
xor UO_1976 (O_1976,N_19855,N_19914);
nor UO_1977 (O_1977,N_19903,N_19884);
nand UO_1978 (O_1978,N_19999,N_19984);
nand UO_1979 (O_1979,N_19888,N_19844);
and UO_1980 (O_1980,N_19999,N_19896);
nand UO_1981 (O_1981,N_19858,N_19841);
xor UO_1982 (O_1982,N_19852,N_19997);
and UO_1983 (O_1983,N_19856,N_19963);
or UO_1984 (O_1984,N_19846,N_19965);
xnor UO_1985 (O_1985,N_19979,N_19888);
nand UO_1986 (O_1986,N_19893,N_19915);
and UO_1987 (O_1987,N_19869,N_19917);
nand UO_1988 (O_1988,N_19922,N_19915);
xor UO_1989 (O_1989,N_19957,N_19968);
xor UO_1990 (O_1990,N_19937,N_19868);
nand UO_1991 (O_1991,N_19934,N_19853);
and UO_1992 (O_1992,N_19976,N_19903);
and UO_1993 (O_1993,N_19874,N_19843);
or UO_1994 (O_1994,N_19910,N_19888);
xor UO_1995 (O_1995,N_19850,N_19906);
nor UO_1996 (O_1996,N_19961,N_19975);
nand UO_1997 (O_1997,N_19904,N_19994);
or UO_1998 (O_1998,N_19892,N_19889);
and UO_1999 (O_1999,N_19919,N_19954);
nor UO_2000 (O_2000,N_19959,N_19877);
nor UO_2001 (O_2001,N_19853,N_19886);
nor UO_2002 (O_2002,N_19870,N_19931);
xnor UO_2003 (O_2003,N_19953,N_19909);
or UO_2004 (O_2004,N_19951,N_19919);
xor UO_2005 (O_2005,N_19907,N_19847);
nor UO_2006 (O_2006,N_19924,N_19862);
and UO_2007 (O_2007,N_19973,N_19954);
nand UO_2008 (O_2008,N_19854,N_19902);
nand UO_2009 (O_2009,N_19874,N_19850);
or UO_2010 (O_2010,N_19945,N_19862);
nand UO_2011 (O_2011,N_19971,N_19898);
and UO_2012 (O_2012,N_19934,N_19850);
nand UO_2013 (O_2013,N_19922,N_19982);
and UO_2014 (O_2014,N_19957,N_19946);
and UO_2015 (O_2015,N_19846,N_19928);
xnor UO_2016 (O_2016,N_19939,N_19865);
nor UO_2017 (O_2017,N_19860,N_19881);
and UO_2018 (O_2018,N_19921,N_19929);
and UO_2019 (O_2019,N_19981,N_19968);
nand UO_2020 (O_2020,N_19897,N_19962);
nand UO_2021 (O_2021,N_19890,N_19968);
and UO_2022 (O_2022,N_19966,N_19937);
nor UO_2023 (O_2023,N_19894,N_19985);
and UO_2024 (O_2024,N_19866,N_19923);
and UO_2025 (O_2025,N_19852,N_19925);
nor UO_2026 (O_2026,N_19967,N_19981);
nand UO_2027 (O_2027,N_19887,N_19972);
or UO_2028 (O_2028,N_19954,N_19911);
nor UO_2029 (O_2029,N_19960,N_19896);
nor UO_2030 (O_2030,N_19958,N_19940);
nor UO_2031 (O_2031,N_19955,N_19908);
and UO_2032 (O_2032,N_19877,N_19946);
nand UO_2033 (O_2033,N_19854,N_19934);
nor UO_2034 (O_2034,N_19913,N_19859);
nand UO_2035 (O_2035,N_19845,N_19908);
and UO_2036 (O_2036,N_19932,N_19847);
or UO_2037 (O_2037,N_19984,N_19939);
nand UO_2038 (O_2038,N_19889,N_19988);
xor UO_2039 (O_2039,N_19974,N_19903);
xor UO_2040 (O_2040,N_19875,N_19976);
xnor UO_2041 (O_2041,N_19889,N_19928);
or UO_2042 (O_2042,N_19862,N_19899);
nand UO_2043 (O_2043,N_19970,N_19948);
and UO_2044 (O_2044,N_19874,N_19981);
and UO_2045 (O_2045,N_19985,N_19847);
xor UO_2046 (O_2046,N_19869,N_19845);
xor UO_2047 (O_2047,N_19848,N_19856);
nor UO_2048 (O_2048,N_19992,N_19886);
nand UO_2049 (O_2049,N_19924,N_19921);
or UO_2050 (O_2050,N_19865,N_19937);
or UO_2051 (O_2051,N_19895,N_19955);
nor UO_2052 (O_2052,N_19979,N_19964);
nor UO_2053 (O_2053,N_19990,N_19915);
and UO_2054 (O_2054,N_19985,N_19951);
nand UO_2055 (O_2055,N_19926,N_19976);
and UO_2056 (O_2056,N_19969,N_19927);
xor UO_2057 (O_2057,N_19957,N_19937);
or UO_2058 (O_2058,N_19941,N_19920);
xor UO_2059 (O_2059,N_19882,N_19963);
xnor UO_2060 (O_2060,N_19862,N_19866);
and UO_2061 (O_2061,N_19933,N_19892);
nand UO_2062 (O_2062,N_19935,N_19887);
nand UO_2063 (O_2063,N_19924,N_19935);
xnor UO_2064 (O_2064,N_19959,N_19847);
xor UO_2065 (O_2065,N_19903,N_19948);
or UO_2066 (O_2066,N_19875,N_19934);
and UO_2067 (O_2067,N_19996,N_19862);
nand UO_2068 (O_2068,N_19981,N_19844);
nor UO_2069 (O_2069,N_19909,N_19974);
nand UO_2070 (O_2070,N_19959,N_19955);
nor UO_2071 (O_2071,N_19880,N_19997);
xor UO_2072 (O_2072,N_19925,N_19941);
nand UO_2073 (O_2073,N_19944,N_19857);
or UO_2074 (O_2074,N_19862,N_19913);
and UO_2075 (O_2075,N_19924,N_19867);
nand UO_2076 (O_2076,N_19972,N_19864);
nand UO_2077 (O_2077,N_19905,N_19958);
nand UO_2078 (O_2078,N_19996,N_19931);
or UO_2079 (O_2079,N_19847,N_19917);
xnor UO_2080 (O_2080,N_19888,N_19963);
and UO_2081 (O_2081,N_19916,N_19988);
nand UO_2082 (O_2082,N_19949,N_19915);
and UO_2083 (O_2083,N_19859,N_19847);
xor UO_2084 (O_2084,N_19957,N_19977);
nand UO_2085 (O_2085,N_19992,N_19912);
nor UO_2086 (O_2086,N_19856,N_19874);
or UO_2087 (O_2087,N_19922,N_19844);
nand UO_2088 (O_2088,N_19934,N_19931);
or UO_2089 (O_2089,N_19852,N_19857);
and UO_2090 (O_2090,N_19878,N_19889);
and UO_2091 (O_2091,N_19938,N_19985);
and UO_2092 (O_2092,N_19893,N_19933);
nand UO_2093 (O_2093,N_19912,N_19961);
or UO_2094 (O_2094,N_19953,N_19924);
xor UO_2095 (O_2095,N_19987,N_19990);
xnor UO_2096 (O_2096,N_19853,N_19925);
nor UO_2097 (O_2097,N_19938,N_19926);
and UO_2098 (O_2098,N_19970,N_19897);
or UO_2099 (O_2099,N_19853,N_19937);
xor UO_2100 (O_2100,N_19896,N_19994);
nor UO_2101 (O_2101,N_19914,N_19940);
and UO_2102 (O_2102,N_19961,N_19856);
nand UO_2103 (O_2103,N_19874,N_19991);
or UO_2104 (O_2104,N_19842,N_19940);
and UO_2105 (O_2105,N_19954,N_19865);
and UO_2106 (O_2106,N_19858,N_19984);
and UO_2107 (O_2107,N_19993,N_19913);
nand UO_2108 (O_2108,N_19961,N_19997);
or UO_2109 (O_2109,N_19998,N_19858);
nand UO_2110 (O_2110,N_19919,N_19888);
or UO_2111 (O_2111,N_19864,N_19949);
nand UO_2112 (O_2112,N_19986,N_19998);
and UO_2113 (O_2113,N_19995,N_19842);
and UO_2114 (O_2114,N_19893,N_19961);
nor UO_2115 (O_2115,N_19849,N_19953);
nand UO_2116 (O_2116,N_19847,N_19997);
xor UO_2117 (O_2117,N_19912,N_19950);
or UO_2118 (O_2118,N_19861,N_19840);
nand UO_2119 (O_2119,N_19930,N_19874);
xnor UO_2120 (O_2120,N_19909,N_19846);
xor UO_2121 (O_2121,N_19901,N_19850);
nor UO_2122 (O_2122,N_19845,N_19922);
or UO_2123 (O_2123,N_19895,N_19935);
xor UO_2124 (O_2124,N_19945,N_19910);
nand UO_2125 (O_2125,N_19840,N_19876);
or UO_2126 (O_2126,N_19867,N_19963);
and UO_2127 (O_2127,N_19984,N_19862);
xnor UO_2128 (O_2128,N_19914,N_19933);
and UO_2129 (O_2129,N_19983,N_19849);
xor UO_2130 (O_2130,N_19914,N_19920);
or UO_2131 (O_2131,N_19964,N_19910);
and UO_2132 (O_2132,N_19892,N_19840);
or UO_2133 (O_2133,N_19873,N_19865);
and UO_2134 (O_2134,N_19875,N_19931);
nor UO_2135 (O_2135,N_19964,N_19958);
and UO_2136 (O_2136,N_19981,N_19989);
nand UO_2137 (O_2137,N_19892,N_19942);
nor UO_2138 (O_2138,N_19985,N_19972);
nand UO_2139 (O_2139,N_19945,N_19989);
nor UO_2140 (O_2140,N_19855,N_19861);
or UO_2141 (O_2141,N_19852,N_19870);
and UO_2142 (O_2142,N_19870,N_19848);
and UO_2143 (O_2143,N_19940,N_19946);
nand UO_2144 (O_2144,N_19929,N_19887);
and UO_2145 (O_2145,N_19954,N_19849);
and UO_2146 (O_2146,N_19862,N_19922);
or UO_2147 (O_2147,N_19850,N_19857);
or UO_2148 (O_2148,N_19915,N_19961);
nand UO_2149 (O_2149,N_19951,N_19983);
and UO_2150 (O_2150,N_19881,N_19994);
and UO_2151 (O_2151,N_19842,N_19863);
or UO_2152 (O_2152,N_19940,N_19999);
or UO_2153 (O_2153,N_19888,N_19943);
nand UO_2154 (O_2154,N_19864,N_19841);
and UO_2155 (O_2155,N_19846,N_19914);
and UO_2156 (O_2156,N_19892,N_19946);
nand UO_2157 (O_2157,N_19954,N_19975);
nor UO_2158 (O_2158,N_19857,N_19841);
nand UO_2159 (O_2159,N_19963,N_19847);
nand UO_2160 (O_2160,N_19999,N_19916);
nand UO_2161 (O_2161,N_19954,N_19896);
and UO_2162 (O_2162,N_19892,N_19995);
nand UO_2163 (O_2163,N_19932,N_19955);
xnor UO_2164 (O_2164,N_19914,N_19931);
and UO_2165 (O_2165,N_19951,N_19959);
xnor UO_2166 (O_2166,N_19870,N_19925);
xor UO_2167 (O_2167,N_19989,N_19852);
nand UO_2168 (O_2168,N_19922,N_19951);
and UO_2169 (O_2169,N_19945,N_19962);
and UO_2170 (O_2170,N_19925,N_19961);
and UO_2171 (O_2171,N_19898,N_19923);
nor UO_2172 (O_2172,N_19858,N_19977);
and UO_2173 (O_2173,N_19874,N_19871);
xnor UO_2174 (O_2174,N_19956,N_19991);
nor UO_2175 (O_2175,N_19965,N_19845);
xor UO_2176 (O_2176,N_19951,N_19940);
nor UO_2177 (O_2177,N_19876,N_19955);
xnor UO_2178 (O_2178,N_19858,N_19964);
nand UO_2179 (O_2179,N_19906,N_19936);
or UO_2180 (O_2180,N_19878,N_19974);
nor UO_2181 (O_2181,N_19944,N_19861);
xor UO_2182 (O_2182,N_19844,N_19903);
xor UO_2183 (O_2183,N_19999,N_19998);
xnor UO_2184 (O_2184,N_19922,N_19993);
and UO_2185 (O_2185,N_19975,N_19882);
xor UO_2186 (O_2186,N_19937,N_19952);
and UO_2187 (O_2187,N_19947,N_19970);
xnor UO_2188 (O_2188,N_19935,N_19900);
nor UO_2189 (O_2189,N_19859,N_19869);
nand UO_2190 (O_2190,N_19968,N_19916);
nand UO_2191 (O_2191,N_19997,N_19844);
nor UO_2192 (O_2192,N_19954,N_19863);
nand UO_2193 (O_2193,N_19901,N_19857);
nor UO_2194 (O_2194,N_19949,N_19906);
nor UO_2195 (O_2195,N_19842,N_19964);
and UO_2196 (O_2196,N_19945,N_19908);
and UO_2197 (O_2197,N_19915,N_19972);
xnor UO_2198 (O_2198,N_19995,N_19921);
nor UO_2199 (O_2199,N_19955,N_19867);
or UO_2200 (O_2200,N_19877,N_19973);
nand UO_2201 (O_2201,N_19933,N_19863);
or UO_2202 (O_2202,N_19949,N_19909);
and UO_2203 (O_2203,N_19867,N_19864);
nand UO_2204 (O_2204,N_19966,N_19999);
nor UO_2205 (O_2205,N_19997,N_19966);
and UO_2206 (O_2206,N_19867,N_19986);
nor UO_2207 (O_2207,N_19901,N_19989);
xor UO_2208 (O_2208,N_19992,N_19841);
nand UO_2209 (O_2209,N_19840,N_19872);
or UO_2210 (O_2210,N_19980,N_19975);
xnor UO_2211 (O_2211,N_19902,N_19843);
xor UO_2212 (O_2212,N_19936,N_19869);
nor UO_2213 (O_2213,N_19876,N_19877);
xor UO_2214 (O_2214,N_19966,N_19969);
nand UO_2215 (O_2215,N_19850,N_19935);
and UO_2216 (O_2216,N_19877,N_19864);
nand UO_2217 (O_2217,N_19995,N_19959);
nor UO_2218 (O_2218,N_19933,N_19897);
nand UO_2219 (O_2219,N_19896,N_19992);
nor UO_2220 (O_2220,N_19920,N_19907);
xnor UO_2221 (O_2221,N_19840,N_19956);
nand UO_2222 (O_2222,N_19869,N_19992);
nor UO_2223 (O_2223,N_19877,N_19890);
nor UO_2224 (O_2224,N_19985,N_19989);
or UO_2225 (O_2225,N_19932,N_19855);
xnor UO_2226 (O_2226,N_19896,N_19891);
and UO_2227 (O_2227,N_19848,N_19850);
xnor UO_2228 (O_2228,N_19847,N_19961);
nor UO_2229 (O_2229,N_19941,N_19887);
nand UO_2230 (O_2230,N_19952,N_19980);
and UO_2231 (O_2231,N_19905,N_19929);
nor UO_2232 (O_2232,N_19985,N_19921);
xnor UO_2233 (O_2233,N_19978,N_19883);
or UO_2234 (O_2234,N_19934,N_19869);
or UO_2235 (O_2235,N_19879,N_19940);
nand UO_2236 (O_2236,N_19906,N_19935);
nand UO_2237 (O_2237,N_19909,N_19921);
xnor UO_2238 (O_2238,N_19877,N_19901);
xor UO_2239 (O_2239,N_19976,N_19933);
xnor UO_2240 (O_2240,N_19933,N_19889);
nand UO_2241 (O_2241,N_19982,N_19875);
nand UO_2242 (O_2242,N_19929,N_19949);
and UO_2243 (O_2243,N_19951,N_19871);
nor UO_2244 (O_2244,N_19966,N_19864);
xor UO_2245 (O_2245,N_19916,N_19995);
nand UO_2246 (O_2246,N_19849,N_19997);
nand UO_2247 (O_2247,N_19978,N_19956);
or UO_2248 (O_2248,N_19889,N_19855);
or UO_2249 (O_2249,N_19845,N_19977);
or UO_2250 (O_2250,N_19997,N_19922);
and UO_2251 (O_2251,N_19950,N_19880);
or UO_2252 (O_2252,N_19969,N_19929);
nand UO_2253 (O_2253,N_19844,N_19972);
nand UO_2254 (O_2254,N_19914,N_19863);
nor UO_2255 (O_2255,N_19924,N_19851);
nand UO_2256 (O_2256,N_19926,N_19877);
nor UO_2257 (O_2257,N_19961,N_19883);
xor UO_2258 (O_2258,N_19965,N_19916);
xnor UO_2259 (O_2259,N_19990,N_19858);
xor UO_2260 (O_2260,N_19897,N_19972);
nor UO_2261 (O_2261,N_19991,N_19936);
and UO_2262 (O_2262,N_19973,N_19889);
nand UO_2263 (O_2263,N_19936,N_19939);
or UO_2264 (O_2264,N_19901,N_19984);
or UO_2265 (O_2265,N_19883,N_19882);
or UO_2266 (O_2266,N_19961,N_19970);
nand UO_2267 (O_2267,N_19925,N_19963);
nor UO_2268 (O_2268,N_19912,N_19867);
xnor UO_2269 (O_2269,N_19901,N_19873);
nor UO_2270 (O_2270,N_19934,N_19844);
or UO_2271 (O_2271,N_19964,N_19948);
nor UO_2272 (O_2272,N_19884,N_19938);
and UO_2273 (O_2273,N_19908,N_19986);
nand UO_2274 (O_2274,N_19852,N_19986);
nand UO_2275 (O_2275,N_19964,N_19915);
xnor UO_2276 (O_2276,N_19967,N_19993);
or UO_2277 (O_2277,N_19964,N_19843);
or UO_2278 (O_2278,N_19906,N_19909);
nor UO_2279 (O_2279,N_19912,N_19903);
or UO_2280 (O_2280,N_19855,N_19883);
xor UO_2281 (O_2281,N_19859,N_19956);
nor UO_2282 (O_2282,N_19969,N_19960);
xnor UO_2283 (O_2283,N_19980,N_19852);
xnor UO_2284 (O_2284,N_19962,N_19893);
and UO_2285 (O_2285,N_19987,N_19852);
and UO_2286 (O_2286,N_19912,N_19885);
or UO_2287 (O_2287,N_19988,N_19895);
nand UO_2288 (O_2288,N_19867,N_19914);
nand UO_2289 (O_2289,N_19866,N_19844);
xor UO_2290 (O_2290,N_19994,N_19969);
nor UO_2291 (O_2291,N_19945,N_19937);
and UO_2292 (O_2292,N_19925,N_19877);
xnor UO_2293 (O_2293,N_19846,N_19934);
xnor UO_2294 (O_2294,N_19940,N_19987);
or UO_2295 (O_2295,N_19989,N_19872);
nor UO_2296 (O_2296,N_19991,N_19997);
nor UO_2297 (O_2297,N_19843,N_19842);
nand UO_2298 (O_2298,N_19847,N_19898);
nor UO_2299 (O_2299,N_19991,N_19869);
and UO_2300 (O_2300,N_19860,N_19987);
and UO_2301 (O_2301,N_19999,N_19986);
nor UO_2302 (O_2302,N_19880,N_19976);
and UO_2303 (O_2303,N_19966,N_19988);
nand UO_2304 (O_2304,N_19879,N_19953);
nand UO_2305 (O_2305,N_19967,N_19849);
xor UO_2306 (O_2306,N_19999,N_19881);
xnor UO_2307 (O_2307,N_19960,N_19886);
or UO_2308 (O_2308,N_19843,N_19978);
nand UO_2309 (O_2309,N_19874,N_19928);
or UO_2310 (O_2310,N_19993,N_19935);
nand UO_2311 (O_2311,N_19846,N_19858);
or UO_2312 (O_2312,N_19860,N_19897);
nand UO_2313 (O_2313,N_19900,N_19967);
nor UO_2314 (O_2314,N_19851,N_19878);
xnor UO_2315 (O_2315,N_19864,N_19970);
nand UO_2316 (O_2316,N_19879,N_19886);
xnor UO_2317 (O_2317,N_19895,N_19875);
nor UO_2318 (O_2318,N_19978,N_19991);
nor UO_2319 (O_2319,N_19879,N_19934);
or UO_2320 (O_2320,N_19905,N_19937);
nor UO_2321 (O_2321,N_19964,N_19847);
nor UO_2322 (O_2322,N_19975,N_19875);
nor UO_2323 (O_2323,N_19905,N_19841);
nand UO_2324 (O_2324,N_19856,N_19861);
and UO_2325 (O_2325,N_19895,N_19969);
nand UO_2326 (O_2326,N_19943,N_19941);
nor UO_2327 (O_2327,N_19947,N_19940);
and UO_2328 (O_2328,N_19880,N_19855);
nand UO_2329 (O_2329,N_19940,N_19923);
xnor UO_2330 (O_2330,N_19925,N_19998);
nand UO_2331 (O_2331,N_19978,N_19871);
or UO_2332 (O_2332,N_19902,N_19954);
nand UO_2333 (O_2333,N_19904,N_19856);
or UO_2334 (O_2334,N_19871,N_19925);
xnor UO_2335 (O_2335,N_19999,N_19866);
nand UO_2336 (O_2336,N_19843,N_19887);
nor UO_2337 (O_2337,N_19969,N_19923);
and UO_2338 (O_2338,N_19930,N_19967);
nor UO_2339 (O_2339,N_19901,N_19968);
xnor UO_2340 (O_2340,N_19944,N_19882);
and UO_2341 (O_2341,N_19888,N_19980);
or UO_2342 (O_2342,N_19892,N_19998);
nand UO_2343 (O_2343,N_19864,N_19872);
and UO_2344 (O_2344,N_19967,N_19907);
nor UO_2345 (O_2345,N_19976,N_19915);
nor UO_2346 (O_2346,N_19905,N_19995);
and UO_2347 (O_2347,N_19842,N_19987);
and UO_2348 (O_2348,N_19987,N_19952);
and UO_2349 (O_2349,N_19894,N_19980);
xor UO_2350 (O_2350,N_19873,N_19972);
or UO_2351 (O_2351,N_19908,N_19846);
xnor UO_2352 (O_2352,N_19993,N_19896);
xor UO_2353 (O_2353,N_19978,N_19921);
or UO_2354 (O_2354,N_19891,N_19912);
and UO_2355 (O_2355,N_19878,N_19953);
nor UO_2356 (O_2356,N_19897,N_19904);
or UO_2357 (O_2357,N_19885,N_19972);
nand UO_2358 (O_2358,N_19847,N_19981);
and UO_2359 (O_2359,N_19966,N_19897);
and UO_2360 (O_2360,N_19942,N_19939);
nand UO_2361 (O_2361,N_19922,N_19858);
nand UO_2362 (O_2362,N_19852,N_19969);
nand UO_2363 (O_2363,N_19864,N_19901);
or UO_2364 (O_2364,N_19935,N_19977);
and UO_2365 (O_2365,N_19953,N_19926);
nand UO_2366 (O_2366,N_19895,N_19938);
xor UO_2367 (O_2367,N_19932,N_19890);
nor UO_2368 (O_2368,N_19938,N_19841);
nor UO_2369 (O_2369,N_19863,N_19840);
or UO_2370 (O_2370,N_19994,N_19937);
nand UO_2371 (O_2371,N_19878,N_19881);
nand UO_2372 (O_2372,N_19933,N_19998);
nor UO_2373 (O_2373,N_19907,N_19882);
nor UO_2374 (O_2374,N_19970,N_19939);
or UO_2375 (O_2375,N_19884,N_19971);
and UO_2376 (O_2376,N_19882,N_19889);
nor UO_2377 (O_2377,N_19973,N_19931);
or UO_2378 (O_2378,N_19859,N_19938);
xor UO_2379 (O_2379,N_19909,N_19962);
and UO_2380 (O_2380,N_19889,N_19935);
nor UO_2381 (O_2381,N_19972,N_19982);
nor UO_2382 (O_2382,N_19939,N_19959);
and UO_2383 (O_2383,N_19927,N_19902);
nor UO_2384 (O_2384,N_19946,N_19939);
nand UO_2385 (O_2385,N_19881,N_19992);
and UO_2386 (O_2386,N_19857,N_19974);
and UO_2387 (O_2387,N_19923,N_19847);
nor UO_2388 (O_2388,N_19975,N_19989);
xnor UO_2389 (O_2389,N_19908,N_19940);
nor UO_2390 (O_2390,N_19923,N_19904);
and UO_2391 (O_2391,N_19925,N_19973);
nor UO_2392 (O_2392,N_19854,N_19883);
xor UO_2393 (O_2393,N_19922,N_19882);
nor UO_2394 (O_2394,N_19886,N_19840);
nor UO_2395 (O_2395,N_19897,N_19846);
xor UO_2396 (O_2396,N_19991,N_19917);
or UO_2397 (O_2397,N_19867,N_19917);
and UO_2398 (O_2398,N_19988,N_19903);
or UO_2399 (O_2399,N_19953,N_19930);
nand UO_2400 (O_2400,N_19999,N_19944);
xnor UO_2401 (O_2401,N_19975,N_19960);
and UO_2402 (O_2402,N_19920,N_19863);
nand UO_2403 (O_2403,N_19967,N_19987);
and UO_2404 (O_2404,N_19920,N_19969);
xor UO_2405 (O_2405,N_19925,N_19988);
and UO_2406 (O_2406,N_19854,N_19905);
or UO_2407 (O_2407,N_19854,N_19913);
nor UO_2408 (O_2408,N_19962,N_19921);
nand UO_2409 (O_2409,N_19966,N_19957);
and UO_2410 (O_2410,N_19850,N_19939);
or UO_2411 (O_2411,N_19851,N_19863);
xnor UO_2412 (O_2412,N_19953,N_19846);
nor UO_2413 (O_2413,N_19876,N_19860);
and UO_2414 (O_2414,N_19890,N_19972);
xnor UO_2415 (O_2415,N_19864,N_19881);
nor UO_2416 (O_2416,N_19979,N_19917);
nor UO_2417 (O_2417,N_19978,N_19957);
and UO_2418 (O_2418,N_19959,N_19960);
nand UO_2419 (O_2419,N_19891,N_19931);
nor UO_2420 (O_2420,N_19889,N_19981);
and UO_2421 (O_2421,N_19924,N_19887);
and UO_2422 (O_2422,N_19840,N_19995);
nor UO_2423 (O_2423,N_19864,N_19965);
xnor UO_2424 (O_2424,N_19954,N_19981);
nand UO_2425 (O_2425,N_19844,N_19842);
or UO_2426 (O_2426,N_19985,N_19934);
and UO_2427 (O_2427,N_19864,N_19984);
nor UO_2428 (O_2428,N_19967,N_19980);
nor UO_2429 (O_2429,N_19987,N_19882);
and UO_2430 (O_2430,N_19962,N_19867);
nor UO_2431 (O_2431,N_19864,N_19909);
nor UO_2432 (O_2432,N_19890,N_19974);
nor UO_2433 (O_2433,N_19953,N_19991);
nor UO_2434 (O_2434,N_19981,N_19949);
and UO_2435 (O_2435,N_19984,N_19985);
xor UO_2436 (O_2436,N_19942,N_19894);
xor UO_2437 (O_2437,N_19960,N_19909);
or UO_2438 (O_2438,N_19915,N_19950);
or UO_2439 (O_2439,N_19971,N_19851);
and UO_2440 (O_2440,N_19968,N_19983);
xnor UO_2441 (O_2441,N_19997,N_19941);
xor UO_2442 (O_2442,N_19842,N_19934);
and UO_2443 (O_2443,N_19849,N_19888);
nor UO_2444 (O_2444,N_19873,N_19931);
nand UO_2445 (O_2445,N_19863,N_19995);
and UO_2446 (O_2446,N_19944,N_19897);
or UO_2447 (O_2447,N_19911,N_19870);
nor UO_2448 (O_2448,N_19845,N_19943);
nor UO_2449 (O_2449,N_19903,N_19916);
xnor UO_2450 (O_2450,N_19966,N_19886);
nand UO_2451 (O_2451,N_19913,N_19850);
nor UO_2452 (O_2452,N_19916,N_19892);
and UO_2453 (O_2453,N_19945,N_19974);
nor UO_2454 (O_2454,N_19916,N_19985);
and UO_2455 (O_2455,N_19959,N_19849);
or UO_2456 (O_2456,N_19958,N_19971);
nor UO_2457 (O_2457,N_19881,N_19861);
xnor UO_2458 (O_2458,N_19949,N_19991);
xor UO_2459 (O_2459,N_19919,N_19956);
and UO_2460 (O_2460,N_19889,N_19964);
and UO_2461 (O_2461,N_19945,N_19995);
and UO_2462 (O_2462,N_19951,N_19899);
xor UO_2463 (O_2463,N_19978,N_19881);
and UO_2464 (O_2464,N_19881,N_19880);
and UO_2465 (O_2465,N_19866,N_19997);
or UO_2466 (O_2466,N_19993,N_19905);
or UO_2467 (O_2467,N_19950,N_19851);
nor UO_2468 (O_2468,N_19897,N_19898);
nand UO_2469 (O_2469,N_19913,N_19878);
or UO_2470 (O_2470,N_19928,N_19917);
xor UO_2471 (O_2471,N_19900,N_19955);
nor UO_2472 (O_2472,N_19873,N_19872);
nor UO_2473 (O_2473,N_19931,N_19911);
xnor UO_2474 (O_2474,N_19846,N_19866);
nor UO_2475 (O_2475,N_19959,N_19981);
xor UO_2476 (O_2476,N_19993,N_19928);
nor UO_2477 (O_2477,N_19944,N_19868);
nand UO_2478 (O_2478,N_19850,N_19894);
and UO_2479 (O_2479,N_19977,N_19980);
or UO_2480 (O_2480,N_19971,N_19948);
and UO_2481 (O_2481,N_19902,N_19912);
xnor UO_2482 (O_2482,N_19918,N_19907);
nor UO_2483 (O_2483,N_19970,N_19875);
nor UO_2484 (O_2484,N_19860,N_19858);
nand UO_2485 (O_2485,N_19996,N_19857);
xnor UO_2486 (O_2486,N_19857,N_19946);
nor UO_2487 (O_2487,N_19924,N_19930);
xor UO_2488 (O_2488,N_19997,N_19976);
nor UO_2489 (O_2489,N_19853,N_19979);
or UO_2490 (O_2490,N_19948,N_19865);
nor UO_2491 (O_2491,N_19997,N_19999);
and UO_2492 (O_2492,N_19906,N_19959);
or UO_2493 (O_2493,N_19866,N_19864);
or UO_2494 (O_2494,N_19913,N_19896);
xnor UO_2495 (O_2495,N_19918,N_19977);
xnor UO_2496 (O_2496,N_19935,N_19979);
and UO_2497 (O_2497,N_19871,N_19955);
and UO_2498 (O_2498,N_19926,N_19900);
nand UO_2499 (O_2499,N_19979,N_19992);
endmodule