module basic_500_3000_500_5_levels_5xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_101,In_61);
or U1 (N_1,In_435,In_88);
nand U2 (N_2,In_400,In_191);
nand U3 (N_3,In_465,In_215);
nor U4 (N_4,In_351,In_488);
and U5 (N_5,In_125,In_29);
nor U6 (N_6,In_431,In_376);
or U7 (N_7,In_179,In_200);
and U8 (N_8,In_18,In_277);
or U9 (N_9,In_313,In_19);
nor U10 (N_10,In_109,In_487);
nand U11 (N_11,In_76,In_437);
or U12 (N_12,In_104,In_228);
or U13 (N_13,In_159,In_151);
nor U14 (N_14,In_442,In_95);
and U15 (N_15,In_260,In_403);
or U16 (N_16,In_486,In_312);
nand U17 (N_17,In_327,In_479);
nand U18 (N_18,In_378,In_42);
and U19 (N_19,In_340,In_234);
or U20 (N_20,In_254,In_248);
nor U21 (N_21,In_337,In_441);
and U22 (N_22,In_48,In_387);
and U23 (N_23,In_147,In_55);
or U24 (N_24,In_362,In_396);
or U25 (N_25,In_3,In_302);
and U26 (N_26,In_91,In_252);
nor U27 (N_27,In_132,In_350);
nand U28 (N_28,In_402,In_165);
and U29 (N_29,In_107,In_23);
and U30 (N_30,In_253,In_294);
nor U31 (N_31,In_453,In_37);
nand U32 (N_32,In_212,In_461);
nor U33 (N_33,In_390,In_137);
nand U34 (N_34,In_304,In_177);
nor U35 (N_35,In_381,In_231);
and U36 (N_36,In_291,In_448);
nand U37 (N_37,In_17,In_349);
nand U38 (N_38,In_113,In_345);
or U39 (N_39,In_459,In_389);
xor U40 (N_40,In_194,In_422);
and U41 (N_41,In_261,In_183);
nand U42 (N_42,In_222,In_343);
xor U43 (N_43,In_22,In_6);
nor U44 (N_44,In_369,In_67);
or U45 (N_45,In_344,In_8);
or U46 (N_46,In_464,In_146);
or U47 (N_47,In_280,In_223);
nand U48 (N_48,In_54,In_341);
and U49 (N_49,In_237,In_120);
nor U50 (N_50,In_462,In_385);
nor U51 (N_51,In_279,In_450);
nor U52 (N_52,In_423,In_227);
nor U53 (N_53,In_148,In_404);
or U54 (N_54,In_59,In_356);
nand U55 (N_55,In_264,In_289);
nor U56 (N_56,In_5,In_474);
or U57 (N_57,In_367,In_131);
or U58 (N_58,In_92,In_308);
nand U59 (N_59,In_152,In_34);
nor U60 (N_60,In_229,In_207);
nand U61 (N_61,In_499,In_50);
nor U62 (N_62,In_243,In_53);
or U63 (N_63,In_210,In_103);
xor U64 (N_64,In_314,In_161);
nand U65 (N_65,In_320,In_173);
and U66 (N_66,In_399,In_436);
xnor U67 (N_67,In_495,In_489);
nor U68 (N_68,In_43,In_144);
or U69 (N_69,In_418,In_319);
and U70 (N_70,In_143,In_218);
xor U71 (N_71,In_365,In_150);
and U72 (N_72,In_116,In_51);
nor U73 (N_73,In_374,In_384);
nor U74 (N_74,In_130,In_438);
and U75 (N_75,In_174,In_273);
or U76 (N_76,In_219,In_25);
and U77 (N_77,In_117,In_310);
nor U78 (N_78,In_298,In_155);
or U79 (N_79,In_316,In_241);
or U80 (N_80,In_286,In_11);
nand U81 (N_81,In_21,In_110);
nor U82 (N_82,In_469,In_373);
or U83 (N_83,In_138,In_186);
nor U84 (N_84,In_26,In_326);
and U85 (N_85,In_456,In_30);
and U86 (N_86,In_145,In_202);
nand U87 (N_87,In_256,In_409);
nand U88 (N_88,In_424,In_41);
and U89 (N_89,In_49,In_129);
or U90 (N_90,In_375,In_299);
nand U91 (N_91,In_392,In_250);
and U92 (N_92,In_370,In_239);
nand U93 (N_93,In_70,In_328);
nor U94 (N_94,In_108,In_301);
nor U95 (N_95,In_100,In_318);
and U96 (N_96,In_309,In_172);
xnor U97 (N_97,In_245,In_226);
and U98 (N_98,In_342,In_154);
nand U99 (N_99,In_334,In_364);
nor U100 (N_100,In_188,In_336);
and U101 (N_101,In_171,In_262);
nand U102 (N_102,In_307,In_168);
or U103 (N_103,In_118,In_458);
or U104 (N_104,In_346,In_122);
nor U105 (N_105,In_230,In_80);
nor U106 (N_106,In_156,In_139);
nor U107 (N_107,In_325,In_322);
nand U108 (N_108,In_235,In_283);
or U109 (N_109,In_20,In_493);
and U110 (N_110,In_244,In_251);
xor U111 (N_111,In_208,In_447);
nor U112 (N_112,In_394,In_359);
nor U113 (N_113,In_112,In_428);
nand U114 (N_114,In_169,In_383);
or U115 (N_115,In_164,In_170);
nor U116 (N_116,In_380,In_57);
nand U117 (N_117,In_491,In_247);
nor U118 (N_118,In_463,In_119);
xor U119 (N_119,In_472,In_481);
or U120 (N_120,In_457,In_121);
nor U121 (N_121,In_195,In_444);
or U122 (N_122,In_429,In_217);
nand U123 (N_123,In_176,In_377);
and U124 (N_124,In_84,In_124);
or U125 (N_125,In_68,In_204);
nand U126 (N_126,In_240,In_303);
nand U127 (N_127,In_335,In_282);
or U128 (N_128,In_31,In_315);
nor U129 (N_129,In_97,In_232);
and U130 (N_130,In_274,In_216);
or U131 (N_131,In_166,In_93);
or U132 (N_132,In_321,In_87);
and U133 (N_133,In_106,In_269);
nor U134 (N_134,In_407,In_15);
and U135 (N_135,In_77,In_290);
and U136 (N_136,In_178,In_192);
and U137 (N_137,In_85,In_347);
nor U138 (N_138,In_439,In_79);
nor U139 (N_139,In_366,In_111);
or U140 (N_140,In_470,In_323);
nor U141 (N_141,In_368,In_203);
nor U142 (N_142,In_127,In_379);
nor U143 (N_143,In_133,In_467);
and U144 (N_144,In_430,In_187);
nand U145 (N_145,In_311,In_348);
nor U146 (N_146,In_83,In_485);
or U147 (N_147,In_484,In_496);
nand U148 (N_148,In_329,In_4);
xor U149 (N_149,In_278,In_184);
or U150 (N_150,In_24,In_466);
nor U151 (N_151,In_38,In_398);
nand U152 (N_152,In_71,In_405);
nor U153 (N_153,In_288,In_393);
nand U154 (N_154,In_421,In_449);
nand U155 (N_155,In_175,In_333);
and U156 (N_156,In_331,In_63);
nand U157 (N_157,In_445,In_427);
and U158 (N_158,In_89,In_12);
or U159 (N_159,In_236,In_480);
and U160 (N_160,In_454,In_432);
and U161 (N_161,In_416,In_300);
xor U162 (N_162,In_406,In_141);
nor U163 (N_163,In_358,In_1);
nand U164 (N_164,In_136,In_72);
and U165 (N_165,In_397,In_206);
nor U166 (N_166,In_305,In_440);
and U167 (N_167,In_45,In_263);
nand U168 (N_168,In_411,In_413);
and U169 (N_169,In_426,In_296);
or U170 (N_170,In_265,In_47);
nand U171 (N_171,In_477,In_99);
or U172 (N_172,In_455,In_267);
nand U173 (N_173,In_75,In_352);
or U174 (N_174,In_193,In_199);
xnor U175 (N_175,In_190,In_0);
and U176 (N_176,In_180,In_473);
nand U177 (N_177,In_233,In_214);
xnor U178 (N_178,In_443,In_490);
and U179 (N_179,In_293,In_98);
or U180 (N_180,In_255,In_297);
and U181 (N_181,In_324,In_246);
nor U182 (N_182,In_287,In_33);
xnor U183 (N_183,In_13,In_153);
nand U184 (N_184,In_478,In_242);
and U185 (N_185,In_39,In_382);
nor U186 (N_186,In_46,In_306);
or U187 (N_187,In_167,In_205);
or U188 (N_188,In_64,In_7);
and U189 (N_189,In_483,In_275);
nor U190 (N_190,In_281,In_257);
xnor U191 (N_191,In_209,In_238);
nor U192 (N_192,In_330,In_163);
nand U193 (N_193,In_14,In_44);
xor U194 (N_194,In_420,In_94);
and U195 (N_195,In_58,In_52);
nand U196 (N_196,In_419,In_388);
or U197 (N_197,In_73,In_434);
nand U198 (N_198,In_35,In_96);
and U199 (N_199,In_213,In_357);
and U200 (N_200,In_317,In_198);
and U201 (N_201,In_471,In_10);
or U202 (N_202,In_285,In_276);
xor U203 (N_203,In_140,In_82);
or U204 (N_204,In_224,In_149);
nor U205 (N_205,In_258,In_211);
nand U206 (N_206,In_9,In_115);
nand U207 (N_207,In_102,In_182);
and U208 (N_208,In_446,In_189);
or U209 (N_209,In_69,In_408);
or U210 (N_210,In_391,In_414);
nand U211 (N_211,In_401,In_355);
and U212 (N_212,In_332,In_492);
xor U213 (N_213,In_135,In_412);
and U214 (N_214,In_158,In_460);
or U215 (N_215,In_482,In_386);
or U216 (N_216,In_16,In_249);
nand U217 (N_217,In_185,In_498);
xor U218 (N_218,In_295,In_225);
and U219 (N_219,In_268,In_338);
and U220 (N_220,In_181,In_468);
nor U221 (N_221,In_157,In_86);
and U222 (N_222,In_270,In_221);
or U223 (N_223,In_128,In_105);
or U224 (N_224,In_284,In_271);
and U225 (N_225,In_201,In_60);
or U226 (N_226,In_65,In_415);
and U227 (N_227,In_494,In_56);
and U228 (N_228,In_32,In_36);
nor U229 (N_229,In_259,In_66);
xnor U230 (N_230,In_220,In_360);
and U231 (N_231,In_40,In_162);
nand U232 (N_232,In_417,In_114);
or U233 (N_233,In_134,In_90);
and U234 (N_234,In_272,In_363);
nand U235 (N_235,In_410,In_81);
or U236 (N_236,In_395,In_353);
and U237 (N_237,In_292,In_371);
or U238 (N_238,In_126,In_476);
or U239 (N_239,In_475,In_451);
and U240 (N_240,In_142,In_372);
or U241 (N_241,In_160,In_354);
nor U242 (N_242,In_497,In_78);
or U243 (N_243,In_123,In_27);
nand U244 (N_244,In_433,In_28);
nor U245 (N_245,In_266,In_361);
or U246 (N_246,In_196,In_452);
nor U247 (N_247,In_2,In_62);
and U248 (N_248,In_197,In_425);
nor U249 (N_249,In_74,In_339);
nor U250 (N_250,In_339,In_8);
and U251 (N_251,In_63,In_27);
xor U252 (N_252,In_309,In_90);
or U253 (N_253,In_142,In_3);
xnor U254 (N_254,In_422,In_427);
and U255 (N_255,In_295,In_421);
and U256 (N_256,In_161,In_480);
and U257 (N_257,In_459,In_259);
nor U258 (N_258,In_216,In_411);
and U259 (N_259,In_470,In_75);
and U260 (N_260,In_385,In_467);
nor U261 (N_261,In_376,In_140);
and U262 (N_262,In_455,In_286);
xnor U263 (N_263,In_262,In_209);
or U264 (N_264,In_31,In_232);
nor U265 (N_265,In_11,In_448);
and U266 (N_266,In_365,In_494);
or U267 (N_267,In_392,In_315);
nand U268 (N_268,In_144,In_154);
nand U269 (N_269,In_354,In_97);
or U270 (N_270,In_228,In_131);
or U271 (N_271,In_480,In_183);
or U272 (N_272,In_73,In_188);
xnor U273 (N_273,In_361,In_138);
nor U274 (N_274,In_421,In_90);
or U275 (N_275,In_57,In_103);
or U276 (N_276,In_112,In_439);
nand U277 (N_277,In_190,In_61);
and U278 (N_278,In_447,In_112);
xnor U279 (N_279,In_346,In_123);
and U280 (N_280,In_132,In_154);
or U281 (N_281,In_37,In_64);
or U282 (N_282,In_354,In_241);
nor U283 (N_283,In_253,In_173);
nor U284 (N_284,In_64,In_149);
and U285 (N_285,In_264,In_352);
nand U286 (N_286,In_400,In_133);
and U287 (N_287,In_274,In_281);
nand U288 (N_288,In_122,In_344);
or U289 (N_289,In_51,In_494);
nor U290 (N_290,In_231,In_245);
and U291 (N_291,In_169,In_159);
nor U292 (N_292,In_369,In_287);
or U293 (N_293,In_231,In_89);
and U294 (N_294,In_44,In_89);
nor U295 (N_295,In_162,In_122);
nor U296 (N_296,In_397,In_82);
or U297 (N_297,In_359,In_228);
or U298 (N_298,In_213,In_18);
nor U299 (N_299,In_70,In_37);
nor U300 (N_300,In_95,In_15);
nor U301 (N_301,In_94,In_431);
nand U302 (N_302,In_174,In_23);
nor U303 (N_303,In_176,In_494);
xnor U304 (N_304,In_353,In_476);
or U305 (N_305,In_456,In_257);
nand U306 (N_306,In_98,In_135);
and U307 (N_307,In_77,In_11);
or U308 (N_308,In_98,In_424);
xnor U309 (N_309,In_225,In_93);
or U310 (N_310,In_192,In_257);
or U311 (N_311,In_462,In_163);
nand U312 (N_312,In_29,In_132);
nand U313 (N_313,In_294,In_98);
nor U314 (N_314,In_266,In_343);
nor U315 (N_315,In_341,In_423);
and U316 (N_316,In_299,In_199);
nor U317 (N_317,In_395,In_49);
or U318 (N_318,In_211,In_260);
nor U319 (N_319,In_4,In_496);
nor U320 (N_320,In_171,In_42);
or U321 (N_321,In_441,In_467);
and U322 (N_322,In_140,In_119);
nand U323 (N_323,In_137,In_172);
nor U324 (N_324,In_242,In_316);
xnor U325 (N_325,In_391,In_100);
nor U326 (N_326,In_157,In_209);
and U327 (N_327,In_305,In_422);
nor U328 (N_328,In_448,In_24);
and U329 (N_329,In_204,In_305);
nor U330 (N_330,In_448,In_218);
and U331 (N_331,In_326,In_212);
nor U332 (N_332,In_211,In_438);
nand U333 (N_333,In_463,In_123);
nand U334 (N_334,In_250,In_223);
and U335 (N_335,In_299,In_349);
nand U336 (N_336,In_379,In_436);
and U337 (N_337,In_489,In_148);
nand U338 (N_338,In_269,In_147);
or U339 (N_339,In_45,In_238);
and U340 (N_340,In_499,In_34);
or U341 (N_341,In_253,In_126);
nand U342 (N_342,In_138,In_54);
or U343 (N_343,In_433,In_237);
and U344 (N_344,In_413,In_31);
and U345 (N_345,In_95,In_266);
or U346 (N_346,In_63,In_151);
nor U347 (N_347,In_139,In_439);
nor U348 (N_348,In_463,In_295);
and U349 (N_349,In_451,In_230);
nand U350 (N_350,In_476,In_94);
nor U351 (N_351,In_235,In_58);
or U352 (N_352,In_172,In_152);
and U353 (N_353,In_33,In_328);
or U354 (N_354,In_216,In_83);
xnor U355 (N_355,In_151,In_128);
or U356 (N_356,In_379,In_36);
or U357 (N_357,In_323,In_351);
or U358 (N_358,In_387,In_85);
or U359 (N_359,In_206,In_292);
or U360 (N_360,In_275,In_322);
or U361 (N_361,In_417,In_12);
xnor U362 (N_362,In_487,In_104);
and U363 (N_363,In_344,In_29);
xor U364 (N_364,In_486,In_145);
or U365 (N_365,In_499,In_186);
and U366 (N_366,In_454,In_80);
xnor U367 (N_367,In_44,In_40);
or U368 (N_368,In_111,In_52);
nand U369 (N_369,In_426,In_391);
and U370 (N_370,In_128,In_348);
or U371 (N_371,In_267,In_12);
and U372 (N_372,In_423,In_149);
or U373 (N_373,In_172,In_66);
or U374 (N_374,In_443,In_206);
or U375 (N_375,In_463,In_323);
nor U376 (N_376,In_349,In_125);
or U377 (N_377,In_45,In_336);
nor U378 (N_378,In_460,In_2);
nor U379 (N_379,In_365,In_238);
and U380 (N_380,In_342,In_451);
nand U381 (N_381,In_355,In_314);
or U382 (N_382,In_108,In_307);
nand U383 (N_383,In_75,In_210);
or U384 (N_384,In_131,In_300);
nand U385 (N_385,In_187,In_160);
or U386 (N_386,In_79,In_127);
and U387 (N_387,In_325,In_344);
or U388 (N_388,In_497,In_405);
nand U389 (N_389,In_357,In_323);
or U390 (N_390,In_244,In_462);
nand U391 (N_391,In_4,In_362);
nor U392 (N_392,In_279,In_194);
xnor U393 (N_393,In_356,In_472);
nor U394 (N_394,In_213,In_23);
or U395 (N_395,In_358,In_288);
nor U396 (N_396,In_249,In_298);
xnor U397 (N_397,In_258,In_165);
or U398 (N_398,In_358,In_120);
nor U399 (N_399,In_453,In_447);
xnor U400 (N_400,In_273,In_405);
nand U401 (N_401,In_1,In_479);
xnor U402 (N_402,In_455,In_87);
nand U403 (N_403,In_376,In_33);
xor U404 (N_404,In_223,In_218);
nor U405 (N_405,In_340,In_357);
nor U406 (N_406,In_430,In_295);
nor U407 (N_407,In_200,In_489);
nor U408 (N_408,In_206,In_42);
and U409 (N_409,In_381,In_105);
or U410 (N_410,In_431,In_485);
nor U411 (N_411,In_337,In_193);
nand U412 (N_412,In_166,In_352);
nor U413 (N_413,In_126,In_343);
xnor U414 (N_414,In_27,In_283);
nor U415 (N_415,In_413,In_244);
nand U416 (N_416,In_435,In_289);
and U417 (N_417,In_106,In_330);
nand U418 (N_418,In_48,In_132);
nand U419 (N_419,In_15,In_102);
or U420 (N_420,In_236,In_142);
nand U421 (N_421,In_317,In_423);
nand U422 (N_422,In_365,In_268);
xor U423 (N_423,In_375,In_391);
nand U424 (N_424,In_481,In_131);
or U425 (N_425,In_232,In_157);
or U426 (N_426,In_213,In_328);
nor U427 (N_427,In_100,In_70);
or U428 (N_428,In_358,In_133);
or U429 (N_429,In_476,In_477);
nor U430 (N_430,In_13,In_130);
or U431 (N_431,In_62,In_84);
nand U432 (N_432,In_192,In_101);
nor U433 (N_433,In_343,In_301);
or U434 (N_434,In_201,In_125);
nand U435 (N_435,In_461,In_90);
xnor U436 (N_436,In_372,In_252);
nor U437 (N_437,In_380,In_362);
nand U438 (N_438,In_85,In_280);
nand U439 (N_439,In_45,In_314);
xor U440 (N_440,In_444,In_112);
and U441 (N_441,In_435,In_125);
nand U442 (N_442,In_348,In_388);
or U443 (N_443,In_7,In_37);
nor U444 (N_444,In_41,In_465);
and U445 (N_445,In_390,In_442);
nand U446 (N_446,In_407,In_472);
nand U447 (N_447,In_204,In_304);
nand U448 (N_448,In_130,In_185);
and U449 (N_449,In_144,In_423);
nand U450 (N_450,In_441,In_463);
xnor U451 (N_451,In_314,In_444);
xnor U452 (N_452,In_302,In_226);
nor U453 (N_453,In_243,In_33);
and U454 (N_454,In_156,In_425);
and U455 (N_455,In_200,In_258);
nor U456 (N_456,In_456,In_37);
xnor U457 (N_457,In_5,In_228);
nand U458 (N_458,In_253,In_451);
and U459 (N_459,In_438,In_482);
or U460 (N_460,In_255,In_375);
and U461 (N_461,In_43,In_240);
nand U462 (N_462,In_397,In_443);
or U463 (N_463,In_471,In_22);
or U464 (N_464,In_198,In_362);
or U465 (N_465,In_211,In_83);
xor U466 (N_466,In_60,In_409);
nand U467 (N_467,In_179,In_203);
nor U468 (N_468,In_366,In_275);
nand U469 (N_469,In_272,In_328);
or U470 (N_470,In_12,In_20);
xor U471 (N_471,In_118,In_297);
nand U472 (N_472,In_391,In_125);
and U473 (N_473,In_41,In_323);
xor U474 (N_474,In_294,In_177);
nor U475 (N_475,In_234,In_406);
nor U476 (N_476,In_468,In_236);
or U477 (N_477,In_251,In_113);
and U478 (N_478,In_222,In_199);
xor U479 (N_479,In_404,In_355);
nand U480 (N_480,In_383,In_326);
and U481 (N_481,In_439,In_55);
nand U482 (N_482,In_173,In_411);
nor U483 (N_483,In_188,In_269);
and U484 (N_484,In_240,In_312);
or U485 (N_485,In_497,In_32);
nand U486 (N_486,In_216,In_397);
or U487 (N_487,In_10,In_91);
and U488 (N_488,In_489,In_202);
nand U489 (N_489,In_251,In_215);
nor U490 (N_490,In_308,In_415);
nor U491 (N_491,In_43,In_248);
or U492 (N_492,In_128,In_150);
and U493 (N_493,In_32,In_333);
xnor U494 (N_494,In_215,In_488);
nor U495 (N_495,In_28,In_375);
nor U496 (N_496,In_12,In_396);
or U497 (N_497,In_195,In_133);
xnor U498 (N_498,In_77,In_42);
nor U499 (N_499,In_351,In_451);
or U500 (N_500,In_263,In_111);
xor U501 (N_501,In_237,In_324);
and U502 (N_502,In_152,In_344);
and U503 (N_503,In_255,In_291);
and U504 (N_504,In_400,In_307);
xnor U505 (N_505,In_442,In_271);
and U506 (N_506,In_36,In_178);
or U507 (N_507,In_377,In_222);
or U508 (N_508,In_483,In_158);
or U509 (N_509,In_129,In_471);
nand U510 (N_510,In_202,In_344);
nor U511 (N_511,In_268,In_382);
or U512 (N_512,In_443,In_239);
and U513 (N_513,In_262,In_94);
nand U514 (N_514,In_247,In_230);
and U515 (N_515,In_426,In_9);
nand U516 (N_516,In_355,In_58);
and U517 (N_517,In_335,In_336);
nand U518 (N_518,In_389,In_126);
nand U519 (N_519,In_138,In_225);
nand U520 (N_520,In_449,In_420);
and U521 (N_521,In_133,In_264);
and U522 (N_522,In_212,In_175);
or U523 (N_523,In_102,In_189);
or U524 (N_524,In_212,In_54);
or U525 (N_525,In_71,In_4);
and U526 (N_526,In_153,In_242);
nand U527 (N_527,In_240,In_300);
nand U528 (N_528,In_248,In_403);
nor U529 (N_529,In_152,In_64);
nand U530 (N_530,In_345,In_341);
and U531 (N_531,In_203,In_26);
nand U532 (N_532,In_147,In_37);
xnor U533 (N_533,In_337,In_215);
or U534 (N_534,In_291,In_464);
or U535 (N_535,In_364,In_450);
nor U536 (N_536,In_448,In_315);
and U537 (N_537,In_421,In_341);
nand U538 (N_538,In_445,In_110);
and U539 (N_539,In_387,In_332);
and U540 (N_540,In_384,In_440);
or U541 (N_541,In_331,In_98);
xor U542 (N_542,In_369,In_391);
or U543 (N_543,In_494,In_14);
nor U544 (N_544,In_88,In_477);
nand U545 (N_545,In_267,In_446);
nand U546 (N_546,In_209,In_357);
nand U547 (N_547,In_176,In_456);
nor U548 (N_548,In_230,In_167);
nor U549 (N_549,In_164,In_317);
nor U550 (N_550,In_116,In_262);
nand U551 (N_551,In_38,In_99);
and U552 (N_552,In_51,In_274);
nor U553 (N_553,In_377,In_119);
nor U554 (N_554,In_171,In_343);
nand U555 (N_555,In_53,In_319);
or U556 (N_556,In_27,In_0);
or U557 (N_557,In_314,In_134);
nand U558 (N_558,In_395,In_394);
or U559 (N_559,In_375,In_65);
or U560 (N_560,In_185,In_390);
and U561 (N_561,In_450,In_14);
xor U562 (N_562,In_340,In_325);
nor U563 (N_563,In_96,In_280);
or U564 (N_564,In_245,In_99);
nor U565 (N_565,In_12,In_485);
nor U566 (N_566,In_226,In_74);
nor U567 (N_567,In_189,In_469);
nand U568 (N_568,In_93,In_101);
and U569 (N_569,In_476,In_9);
xnor U570 (N_570,In_375,In_292);
nand U571 (N_571,In_404,In_243);
nor U572 (N_572,In_376,In_152);
nor U573 (N_573,In_447,In_48);
nand U574 (N_574,In_51,In_37);
nor U575 (N_575,In_163,In_303);
xor U576 (N_576,In_296,In_146);
nand U577 (N_577,In_3,In_435);
xor U578 (N_578,In_160,In_479);
and U579 (N_579,In_8,In_67);
nor U580 (N_580,In_380,In_9);
or U581 (N_581,In_101,In_318);
and U582 (N_582,In_283,In_322);
nand U583 (N_583,In_420,In_252);
or U584 (N_584,In_387,In_138);
nand U585 (N_585,In_16,In_229);
and U586 (N_586,In_84,In_61);
xor U587 (N_587,In_391,In_219);
nand U588 (N_588,In_148,In_384);
or U589 (N_589,In_383,In_144);
nor U590 (N_590,In_490,In_377);
or U591 (N_591,In_422,In_243);
nand U592 (N_592,In_170,In_179);
and U593 (N_593,In_77,In_93);
or U594 (N_594,In_31,In_85);
or U595 (N_595,In_274,In_375);
nor U596 (N_596,In_370,In_268);
xnor U597 (N_597,In_428,In_482);
xor U598 (N_598,In_47,In_224);
and U599 (N_599,In_60,In_275);
nand U600 (N_600,N_501,N_25);
and U601 (N_601,N_303,N_284);
or U602 (N_602,N_368,N_396);
and U603 (N_603,N_174,N_183);
nand U604 (N_604,N_186,N_397);
xnor U605 (N_605,N_99,N_263);
xnor U606 (N_606,N_209,N_522);
or U607 (N_607,N_0,N_155);
and U608 (N_608,N_227,N_567);
nand U609 (N_609,N_67,N_509);
nor U610 (N_610,N_170,N_257);
nand U611 (N_611,N_167,N_282);
or U612 (N_612,N_456,N_125);
nand U613 (N_613,N_553,N_446);
or U614 (N_614,N_423,N_458);
nand U615 (N_615,N_535,N_225);
nor U616 (N_616,N_376,N_544);
and U617 (N_617,N_547,N_109);
nor U618 (N_618,N_461,N_586);
and U619 (N_619,N_517,N_96);
and U620 (N_620,N_374,N_28);
or U621 (N_621,N_215,N_416);
or U622 (N_622,N_502,N_80);
or U623 (N_623,N_430,N_298);
nor U624 (N_624,N_372,N_74);
nand U625 (N_625,N_415,N_217);
nand U626 (N_626,N_105,N_71);
or U627 (N_627,N_178,N_45);
xor U628 (N_628,N_244,N_400);
and U629 (N_629,N_543,N_271);
or U630 (N_630,N_579,N_134);
nand U631 (N_631,N_56,N_288);
or U632 (N_632,N_47,N_537);
nand U633 (N_633,N_349,N_171);
nand U634 (N_634,N_32,N_103);
nand U635 (N_635,N_172,N_525);
nor U636 (N_636,N_164,N_503);
or U637 (N_637,N_440,N_43);
nor U638 (N_638,N_432,N_393);
nor U639 (N_639,N_68,N_532);
or U640 (N_640,N_574,N_39);
xor U641 (N_641,N_294,N_431);
nor U642 (N_642,N_422,N_580);
nor U643 (N_643,N_314,N_79);
xnor U644 (N_644,N_165,N_255);
or U645 (N_645,N_561,N_587);
or U646 (N_646,N_569,N_573);
or U647 (N_647,N_312,N_38);
or U648 (N_648,N_233,N_176);
nand U649 (N_649,N_281,N_272);
xnor U650 (N_650,N_6,N_98);
nand U651 (N_651,N_588,N_520);
and U652 (N_652,N_146,N_31);
nand U653 (N_653,N_50,N_427);
nor U654 (N_654,N_3,N_137);
nand U655 (N_655,N_229,N_319);
nand U656 (N_656,N_131,N_21);
nand U657 (N_657,N_381,N_377);
or U658 (N_658,N_492,N_221);
and U659 (N_659,N_55,N_191);
and U660 (N_660,N_141,N_121);
nor U661 (N_661,N_127,N_259);
and U662 (N_662,N_292,N_285);
xnor U663 (N_663,N_213,N_526);
or U664 (N_664,N_447,N_538);
nor U665 (N_665,N_250,N_139);
nor U666 (N_666,N_414,N_524);
and U667 (N_667,N_265,N_241);
nand U668 (N_668,N_253,N_455);
nand U669 (N_669,N_236,N_471);
and U670 (N_670,N_407,N_582);
and U671 (N_671,N_404,N_113);
xor U672 (N_672,N_578,N_505);
or U673 (N_673,N_344,N_287);
or U674 (N_674,N_486,N_19);
nor U675 (N_675,N_504,N_453);
xor U676 (N_676,N_110,N_142);
or U677 (N_677,N_514,N_20);
nor U678 (N_678,N_118,N_360);
or U679 (N_679,N_89,N_307);
and U680 (N_680,N_570,N_267);
nand U681 (N_681,N_136,N_340);
and U682 (N_682,N_380,N_460);
and U683 (N_683,N_548,N_278);
nand U684 (N_684,N_402,N_168);
nor U685 (N_685,N_410,N_302);
nand U686 (N_686,N_5,N_391);
or U687 (N_687,N_339,N_40);
nor U688 (N_688,N_104,N_470);
or U689 (N_689,N_334,N_388);
or U690 (N_690,N_9,N_370);
and U691 (N_691,N_92,N_246);
xor U692 (N_692,N_270,N_87);
xnor U693 (N_693,N_542,N_333);
nand U694 (N_694,N_466,N_192);
and U695 (N_695,N_266,N_264);
or U696 (N_696,N_448,N_143);
and U697 (N_697,N_348,N_85);
xor U698 (N_698,N_498,N_315);
nor U699 (N_699,N_474,N_595);
nand U700 (N_700,N_383,N_316);
or U701 (N_701,N_434,N_290);
or U702 (N_702,N_488,N_452);
nand U703 (N_703,N_232,N_478);
and U704 (N_704,N_403,N_584);
or U705 (N_705,N_210,N_425);
nand U706 (N_706,N_347,N_590);
nor U707 (N_707,N_289,N_507);
nand U708 (N_708,N_301,N_467);
nor U709 (N_709,N_169,N_36);
nor U710 (N_710,N_500,N_534);
or U711 (N_711,N_433,N_539);
and U712 (N_712,N_426,N_328);
and U713 (N_713,N_489,N_107);
and U714 (N_714,N_247,N_585);
nor U715 (N_715,N_119,N_30);
nand U716 (N_716,N_592,N_18);
xor U717 (N_717,N_378,N_511);
xnor U718 (N_718,N_476,N_275);
nand U719 (N_719,N_224,N_516);
nor U720 (N_720,N_220,N_256);
or U721 (N_721,N_366,N_490);
and U722 (N_722,N_346,N_386);
nand U723 (N_723,N_81,N_343);
or U724 (N_724,N_419,N_231);
or U725 (N_725,N_297,N_1);
and U726 (N_726,N_219,N_196);
nor U727 (N_727,N_442,N_100);
and U728 (N_728,N_269,N_313);
nor U729 (N_729,N_565,N_394);
nand U730 (N_730,N_166,N_480);
and U731 (N_731,N_154,N_205);
and U732 (N_732,N_296,N_12);
nand U733 (N_733,N_518,N_599);
or U734 (N_734,N_338,N_276);
nand U735 (N_735,N_550,N_559);
nor U736 (N_736,N_162,N_258);
or U737 (N_737,N_175,N_60);
and U738 (N_738,N_536,N_300);
xnor U739 (N_739,N_17,N_35);
nor U740 (N_740,N_412,N_305);
nor U741 (N_741,N_75,N_306);
nand U742 (N_742,N_77,N_126);
nor U743 (N_743,N_475,N_52);
xor U744 (N_744,N_411,N_558);
nor U745 (N_745,N_23,N_353);
and U746 (N_746,N_53,N_223);
and U747 (N_747,N_521,N_180);
nor U748 (N_748,N_150,N_251);
and U749 (N_749,N_530,N_88);
or U750 (N_750,N_323,N_95);
nor U751 (N_751,N_44,N_260);
or U752 (N_752,N_441,N_8);
nand U753 (N_753,N_352,N_409);
nor U754 (N_754,N_133,N_280);
or U755 (N_755,N_373,N_576);
or U756 (N_756,N_128,N_188);
and U757 (N_757,N_234,N_10);
xnor U758 (N_758,N_159,N_462);
nand U759 (N_759,N_214,N_112);
or U760 (N_760,N_345,N_435);
nand U761 (N_761,N_156,N_401);
and U762 (N_762,N_443,N_465);
or U763 (N_763,N_444,N_291);
nor U764 (N_764,N_459,N_204);
nor U765 (N_765,N_384,N_197);
or U766 (N_766,N_274,N_329);
and U767 (N_767,N_22,N_310);
nand U768 (N_768,N_405,N_332);
or U769 (N_769,N_541,N_207);
nor U770 (N_770,N_326,N_575);
nor U771 (N_771,N_212,N_506);
nand U772 (N_772,N_76,N_392);
and U773 (N_773,N_62,N_493);
nor U774 (N_774,N_320,N_322);
xor U775 (N_775,N_571,N_367);
nand U776 (N_776,N_324,N_330);
nand U777 (N_777,N_57,N_439);
xor U778 (N_778,N_240,N_11);
or U779 (N_779,N_54,N_589);
and U780 (N_780,N_37,N_91);
or U781 (N_781,N_140,N_252);
nor U782 (N_782,N_235,N_596);
nor U783 (N_783,N_243,N_515);
or U784 (N_784,N_200,N_108);
xor U785 (N_785,N_46,N_369);
and U786 (N_786,N_293,N_115);
nor U787 (N_787,N_408,N_429);
or U788 (N_788,N_230,N_325);
nand U789 (N_789,N_239,N_563);
nor U790 (N_790,N_189,N_84);
nand U791 (N_791,N_557,N_304);
nor U792 (N_792,N_485,N_318);
xnor U793 (N_793,N_149,N_457);
or U794 (N_794,N_41,N_286);
or U795 (N_795,N_163,N_195);
nand U796 (N_796,N_193,N_202);
or U797 (N_797,N_469,N_523);
or U798 (N_798,N_187,N_577);
or U799 (N_799,N_496,N_158);
and U800 (N_800,N_327,N_375);
or U801 (N_801,N_273,N_237);
nand U802 (N_802,N_116,N_132);
nor U803 (N_803,N_148,N_495);
and U804 (N_804,N_173,N_111);
or U805 (N_805,N_120,N_389);
and U806 (N_806,N_185,N_184);
or U807 (N_807,N_382,N_33);
and U808 (N_808,N_519,N_199);
nor U809 (N_809,N_597,N_24);
or U810 (N_810,N_153,N_211);
nand U811 (N_811,N_61,N_513);
nand U812 (N_812,N_198,N_66);
nor U813 (N_813,N_413,N_365);
or U814 (N_814,N_398,N_331);
nor U815 (N_815,N_179,N_487);
or U816 (N_816,N_445,N_568);
or U817 (N_817,N_145,N_248);
and U818 (N_818,N_437,N_48);
nor U819 (N_819,N_424,N_591);
nand U820 (N_820,N_7,N_182);
nor U821 (N_821,N_72,N_49);
and U822 (N_822,N_529,N_151);
and U823 (N_823,N_463,N_598);
xnor U824 (N_824,N_390,N_510);
nand U825 (N_825,N_560,N_94);
or U826 (N_826,N_546,N_26);
nand U827 (N_827,N_123,N_362);
and U828 (N_828,N_63,N_279);
or U829 (N_829,N_70,N_545);
xnor U830 (N_830,N_566,N_551);
xor U831 (N_831,N_262,N_554);
or U832 (N_832,N_385,N_238);
and U833 (N_833,N_436,N_283);
nand U834 (N_834,N_484,N_473);
nand U835 (N_835,N_117,N_194);
nor U836 (N_836,N_572,N_552);
or U837 (N_837,N_438,N_203);
xnor U838 (N_838,N_152,N_421);
nand U839 (N_839,N_309,N_16);
or U840 (N_840,N_479,N_64);
nand U841 (N_841,N_78,N_387);
nand U842 (N_842,N_512,N_555);
and U843 (N_843,N_508,N_395);
nand U844 (N_844,N_583,N_218);
nor U845 (N_845,N_135,N_160);
nand U846 (N_846,N_102,N_549);
xnor U847 (N_847,N_228,N_13);
or U848 (N_848,N_69,N_295);
nor U849 (N_849,N_308,N_245);
nand U850 (N_850,N_581,N_124);
and U851 (N_851,N_451,N_14);
nand U852 (N_852,N_482,N_499);
or U853 (N_853,N_216,N_42);
or U854 (N_854,N_190,N_564);
and U855 (N_855,N_356,N_379);
nor U856 (N_856,N_147,N_311);
nor U857 (N_857,N_181,N_468);
nor U858 (N_858,N_201,N_491);
or U859 (N_859,N_277,N_15);
nor U860 (N_860,N_157,N_359);
and U861 (N_861,N_335,N_399);
xnor U862 (N_862,N_106,N_428);
and U863 (N_863,N_351,N_59);
and U864 (N_864,N_406,N_355);
and U865 (N_865,N_363,N_336);
and U866 (N_866,N_472,N_222);
nor U867 (N_867,N_254,N_177);
xnor U868 (N_868,N_34,N_364);
or U869 (N_869,N_450,N_27);
and U870 (N_870,N_122,N_73);
nor U871 (N_871,N_533,N_261);
or U872 (N_872,N_93,N_114);
nand U873 (N_873,N_342,N_51);
xor U874 (N_874,N_129,N_540);
or U875 (N_875,N_418,N_65);
nand U876 (N_876,N_161,N_249);
or U877 (N_877,N_354,N_594);
nor U878 (N_878,N_206,N_29);
and U879 (N_879,N_357,N_82);
nand U880 (N_880,N_481,N_556);
nand U881 (N_881,N_341,N_299);
and U882 (N_882,N_58,N_417);
xor U883 (N_883,N_454,N_83);
nor U884 (N_884,N_226,N_562);
and U885 (N_885,N_90,N_497);
and U886 (N_886,N_144,N_449);
nand U887 (N_887,N_420,N_483);
or U888 (N_888,N_4,N_97);
nor U889 (N_889,N_350,N_361);
nor U890 (N_890,N_86,N_268);
xnor U891 (N_891,N_593,N_464);
nand U892 (N_892,N_208,N_358);
and U893 (N_893,N_138,N_528);
or U894 (N_894,N_371,N_2);
nand U895 (N_895,N_531,N_494);
or U896 (N_896,N_477,N_337);
nand U897 (N_897,N_527,N_242);
and U898 (N_898,N_130,N_321);
or U899 (N_899,N_101,N_317);
and U900 (N_900,N_395,N_348);
nor U901 (N_901,N_488,N_121);
nand U902 (N_902,N_546,N_334);
or U903 (N_903,N_409,N_459);
xor U904 (N_904,N_544,N_393);
nand U905 (N_905,N_269,N_443);
nand U906 (N_906,N_445,N_86);
or U907 (N_907,N_243,N_139);
nor U908 (N_908,N_10,N_146);
nor U909 (N_909,N_457,N_374);
nor U910 (N_910,N_309,N_300);
and U911 (N_911,N_549,N_377);
nand U912 (N_912,N_244,N_415);
nand U913 (N_913,N_312,N_387);
or U914 (N_914,N_297,N_290);
xnor U915 (N_915,N_386,N_29);
xnor U916 (N_916,N_519,N_506);
or U917 (N_917,N_464,N_556);
and U918 (N_918,N_392,N_149);
and U919 (N_919,N_4,N_37);
or U920 (N_920,N_203,N_490);
and U921 (N_921,N_357,N_403);
nand U922 (N_922,N_483,N_103);
nand U923 (N_923,N_103,N_161);
and U924 (N_924,N_262,N_274);
or U925 (N_925,N_191,N_291);
and U926 (N_926,N_42,N_19);
nor U927 (N_927,N_164,N_196);
or U928 (N_928,N_431,N_289);
nor U929 (N_929,N_107,N_519);
or U930 (N_930,N_563,N_211);
xnor U931 (N_931,N_483,N_59);
or U932 (N_932,N_5,N_33);
nor U933 (N_933,N_298,N_469);
and U934 (N_934,N_281,N_198);
nor U935 (N_935,N_405,N_386);
and U936 (N_936,N_157,N_340);
and U937 (N_937,N_273,N_378);
nor U938 (N_938,N_599,N_14);
and U939 (N_939,N_304,N_300);
and U940 (N_940,N_375,N_495);
nand U941 (N_941,N_482,N_29);
xor U942 (N_942,N_55,N_466);
and U943 (N_943,N_86,N_54);
nand U944 (N_944,N_374,N_357);
nand U945 (N_945,N_180,N_186);
and U946 (N_946,N_99,N_435);
nand U947 (N_947,N_592,N_107);
and U948 (N_948,N_95,N_160);
nand U949 (N_949,N_594,N_330);
nor U950 (N_950,N_366,N_180);
nand U951 (N_951,N_353,N_462);
xor U952 (N_952,N_374,N_196);
or U953 (N_953,N_209,N_442);
nand U954 (N_954,N_431,N_327);
or U955 (N_955,N_582,N_452);
or U956 (N_956,N_142,N_118);
nor U957 (N_957,N_459,N_116);
xnor U958 (N_958,N_196,N_191);
nand U959 (N_959,N_67,N_491);
nand U960 (N_960,N_211,N_332);
nand U961 (N_961,N_483,N_49);
and U962 (N_962,N_128,N_115);
nor U963 (N_963,N_304,N_85);
and U964 (N_964,N_167,N_16);
and U965 (N_965,N_13,N_220);
or U966 (N_966,N_449,N_67);
nor U967 (N_967,N_122,N_559);
and U968 (N_968,N_89,N_364);
or U969 (N_969,N_311,N_466);
nand U970 (N_970,N_150,N_591);
nand U971 (N_971,N_503,N_502);
xor U972 (N_972,N_522,N_216);
and U973 (N_973,N_508,N_43);
or U974 (N_974,N_422,N_161);
or U975 (N_975,N_311,N_537);
or U976 (N_976,N_533,N_226);
or U977 (N_977,N_276,N_211);
and U978 (N_978,N_12,N_16);
and U979 (N_979,N_467,N_122);
nor U980 (N_980,N_403,N_295);
or U981 (N_981,N_383,N_586);
nor U982 (N_982,N_565,N_253);
nand U983 (N_983,N_259,N_365);
xnor U984 (N_984,N_245,N_39);
nand U985 (N_985,N_32,N_572);
and U986 (N_986,N_92,N_186);
and U987 (N_987,N_127,N_499);
or U988 (N_988,N_134,N_577);
nand U989 (N_989,N_77,N_433);
nand U990 (N_990,N_96,N_71);
and U991 (N_991,N_293,N_432);
xnor U992 (N_992,N_178,N_120);
or U993 (N_993,N_337,N_321);
nand U994 (N_994,N_429,N_541);
nor U995 (N_995,N_388,N_294);
and U996 (N_996,N_363,N_116);
xnor U997 (N_997,N_197,N_576);
xnor U998 (N_998,N_303,N_130);
and U999 (N_999,N_281,N_389);
xor U1000 (N_1000,N_61,N_70);
nor U1001 (N_1001,N_512,N_445);
and U1002 (N_1002,N_478,N_441);
nor U1003 (N_1003,N_399,N_585);
nor U1004 (N_1004,N_503,N_465);
nand U1005 (N_1005,N_398,N_158);
xnor U1006 (N_1006,N_5,N_78);
xor U1007 (N_1007,N_187,N_78);
nor U1008 (N_1008,N_474,N_566);
or U1009 (N_1009,N_548,N_275);
or U1010 (N_1010,N_339,N_580);
or U1011 (N_1011,N_291,N_86);
nor U1012 (N_1012,N_0,N_360);
or U1013 (N_1013,N_529,N_65);
nor U1014 (N_1014,N_521,N_590);
nor U1015 (N_1015,N_281,N_346);
nand U1016 (N_1016,N_507,N_476);
nor U1017 (N_1017,N_449,N_103);
nor U1018 (N_1018,N_78,N_111);
and U1019 (N_1019,N_197,N_370);
and U1020 (N_1020,N_390,N_386);
nand U1021 (N_1021,N_565,N_203);
nand U1022 (N_1022,N_70,N_194);
xnor U1023 (N_1023,N_221,N_296);
nand U1024 (N_1024,N_556,N_32);
nor U1025 (N_1025,N_371,N_159);
and U1026 (N_1026,N_302,N_218);
and U1027 (N_1027,N_309,N_415);
and U1028 (N_1028,N_472,N_417);
nor U1029 (N_1029,N_191,N_539);
nand U1030 (N_1030,N_322,N_394);
and U1031 (N_1031,N_194,N_429);
nand U1032 (N_1032,N_161,N_590);
and U1033 (N_1033,N_487,N_208);
nand U1034 (N_1034,N_319,N_191);
nand U1035 (N_1035,N_218,N_472);
nand U1036 (N_1036,N_483,N_448);
nor U1037 (N_1037,N_469,N_491);
or U1038 (N_1038,N_579,N_143);
xnor U1039 (N_1039,N_598,N_474);
nor U1040 (N_1040,N_136,N_193);
or U1041 (N_1041,N_363,N_184);
nor U1042 (N_1042,N_74,N_535);
nor U1043 (N_1043,N_258,N_287);
and U1044 (N_1044,N_110,N_509);
or U1045 (N_1045,N_333,N_590);
and U1046 (N_1046,N_112,N_310);
or U1047 (N_1047,N_64,N_17);
and U1048 (N_1048,N_517,N_459);
and U1049 (N_1049,N_114,N_168);
nor U1050 (N_1050,N_434,N_88);
nand U1051 (N_1051,N_127,N_377);
or U1052 (N_1052,N_294,N_567);
and U1053 (N_1053,N_362,N_451);
nor U1054 (N_1054,N_397,N_596);
and U1055 (N_1055,N_374,N_461);
nor U1056 (N_1056,N_230,N_195);
and U1057 (N_1057,N_505,N_15);
or U1058 (N_1058,N_32,N_593);
nand U1059 (N_1059,N_160,N_178);
nand U1060 (N_1060,N_1,N_489);
nand U1061 (N_1061,N_292,N_505);
nor U1062 (N_1062,N_173,N_179);
and U1063 (N_1063,N_241,N_203);
nor U1064 (N_1064,N_233,N_256);
nor U1065 (N_1065,N_268,N_227);
or U1066 (N_1066,N_331,N_239);
or U1067 (N_1067,N_488,N_372);
nand U1068 (N_1068,N_281,N_357);
nor U1069 (N_1069,N_81,N_568);
nor U1070 (N_1070,N_236,N_353);
nor U1071 (N_1071,N_58,N_553);
or U1072 (N_1072,N_333,N_495);
and U1073 (N_1073,N_231,N_548);
and U1074 (N_1074,N_409,N_127);
nand U1075 (N_1075,N_95,N_367);
or U1076 (N_1076,N_90,N_364);
or U1077 (N_1077,N_166,N_540);
xnor U1078 (N_1078,N_520,N_157);
nor U1079 (N_1079,N_234,N_525);
and U1080 (N_1080,N_111,N_357);
and U1081 (N_1081,N_487,N_347);
nor U1082 (N_1082,N_491,N_115);
nor U1083 (N_1083,N_468,N_308);
nand U1084 (N_1084,N_50,N_231);
nand U1085 (N_1085,N_187,N_174);
xnor U1086 (N_1086,N_405,N_144);
and U1087 (N_1087,N_568,N_231);
nand U1088 (N_1088,N_31,N_527);
or U1089 (N_1089,N_540,N_36);
xnor U1090 (N_1090,N_585,N_26);
xor U1091 (N_1091,N_181,N_375);
nor U1092 (N_1092,N_291,N_465);
or U1093 (N_1093,N_472,N_176);
or U1094 (N_1094,N_180,N_117);
nand U1095 (N_1095,N_399,N_290);
or U1096 (N_1096,N_515,N_129);
nor U1097 (N_1097,N_352,N_534);
nor U1098 (N_1098,N_113,N_28);
nor U1099 (N_1099,N_410,N_87);
or U1100 (N_1100,N_286,N_403);
nand U1101 (N_1101,N_45,N_140);
and U1102 (N_1102,N_213,N_173);
and U1103 (N_1103,N_360,N_321);
xor U1104 (N_1104,N_501,N_128);
and U1105 (N_1105,N_504,N_573);
and U1106 (N_1106,N_207,N_405);
nor U1107 (N_1107,N_67,N_380);
nor U1108 (N_1108,N_305,N_584);
nand U1109 (N_1109,N_73,N_119);
or U1110 (N_1110,N_157,N_241);
or U1111 (N_1111,N_258,N_530);
nand U1112 (N_1112,N_105,N_113);
nor U1113 (N_1113,N_102,N_325);
nand U1114 (N_1114,N_563,N_119);
nand U1115 (N_1115,N_400,N_435);
and U1116 (N_1116,N_69,N_270);
or U1117 (N_1117,N_263,N_255);
nand U1118 (N_1118,N_166,N_430);
nand U1119 (N_1119,N_467,N_438);
and U1120 (N_1120,N_580,N_596);
and U1121 (N_1121,N_544,N_470);
and U1122 (N_1122,N_588,N_489);
or U1123 (N_1123,N_94,N_119);
nor U1124 (N_1124,N_111,N_134);
nor U1125 (N_1125,N_220,N_265);
nor U1126 (N_1126,N_455,N_448);
nor U1127 (N_1127,N_508,N_24);
xnor U1128 (N_1128,N_220,N_403);
nor U1129 (N_1129,N_84,N_197);
and U1130 (N_1130,N_238,N_173);
nand U1131 (N_1131,N_174,N_17);
or U1132 (N_1132,N_296,N_183);
nand U1133 (N_1133,N_260,N_477);
nand U1134 (N_1134,N_180,N_184);
xnor U1135 (N_1135,N_57,N_114);
nor U1136 (N_1136,N_585,N_99);
nand U1137 (N_1137,N_322,N_407);
nor U1138 (N_1138,N_584,N_90);
or U1139 (N_1139,N_484,N_373);
nor U1140 (N_1140,N_336,N_581);
nor U1141 (N_1141,N_142,N_239);
and U1142 (N_1142,N_341,N_520);
nor U1143 (N_1143,N_592,N_178);
and U1144 (N_1144,N_10,N_370);
or U1145 (N_1145,N_341,N_63);
nor U1146 (N_1146,N_589,N_319);
xor U1147 (N_1147,N_464,N_589);
nor U1148 (N_1148,N_573,N_58);
nand U1149 (N_1149,N_161,N_307);
and U1150 (N_1150,N_121,N_407);
or U1151 (N_1151,N_97,N_202);
nand U1152 (N_1152,N_453,N_30);
and U1153 (N_1153,N_367,N_365);
or U1154 (N_1154,N_454,N_115);
nor U1155 (N_1155,N_181,N_44);
or U1156 (N_1156,N_406,N_523);
or U1157 (N_1157,N_545,N_282);
or U1158 (N_1158,N_116,N_549);
and U1159 (N_1159,N_52,N_74);
and U1160 (N_1160,N_140,N_70);
nand U1161 (N_1161,N_192,N_343);
and U1162 (N_1162,N_254,N_5);
and U1163 (N_1163,N_432,N_51);
nand U1164 (N_1164,N_227,N_154);
nand U1165 (N_1165,N_30,N_102);
or U1166 (N_1166,N_373,N_256);
nor U1167 (N_1167,N_477,N_489);
nand U1168 (N_1168,N_33,N_308);
nor U1169 (N_1169,N_192,N_542);
xor U1170 (N_1170,N_297,N_35);
and U1171 (N_1171,N_79,N_499);
or U1172 (N_1172,N_143,N_271);
and U1173 (N_1173,N_288,N_53);
and U1174 (N_1174,N_237,N_567);
or U1175 (N_1175,N_356,N_479);
or U1176 (N_1176,N_318,N_339);
nor U1177 (N_1177,N_435,N_147);
nor U1178 (N_1178,N_381,N_1);
and U1179 (N_1179,N_247,N_311);
and U1180 (N_1180,N_195,N_470);
and U1181 (N_1181,N_589,N_207);
nand U1182 (N_1182,N_466,N_251);
nor U1183 (N_1183,N_154,N_289);
nand U1184 (N_1184,N_354,N_131);
or U1185 (N_1185,N_515,N_413);
or U1186 (N_1186,N_227,N_164);
xor U1187 (N_1187,N_104,N_49);
xnor U1188 (N_1188,N_466,N_115);
nor U1189 (N_1189,N_100,N_8);
or U1190 (N_1190,N_541,N_227);
and U1191 (N_1191,N_15,N_472);
or U1192 (N_1192,N_433,N_103);
xor U1193 (N_1193,N_442,N_159);
nand U1194 (N_1194,N_229,N_420);
nor U1195 (N_1195,N_365,N_20);
nand U1196 (N_1196,N_545,N_370);
xnor U1197 (N_1197,N_584,N_575);
nand U1198 (N_1198,N_353,N_423);
nor U1199 (N_1199,N_474,N_240);
nor U1200 (N_1200,N_624,N_1011);
nor U1201 (N_1201,N_869,N_983);
or U1202 (N_1202,N_1057,N_769);
nand U1203 (N_1203,N_877,N_1186);
nor U1204 (N_1204,N_787,N_826);
xnor U1205 (N_1205,N_924,N_1121);
or U1206 (N_1206,N_1196,N_1104);
nand U1207 (N_1207,N_821,N_674);
and U1208 (N_1208,N_1005,N_1066);
nor U1209 (N_1209,N_991,N_839);
xnor U1210 (N_1210,N_1063,N_962);
nor U1211 (N_1211,N_794,N_854);
and U1212 (N_1212,N_1188,N_1030);
nand U1213 (N_1213,N_785,N_670);
or U1214 (N_1214,N_691,N_711);
and U1215 (N_1215,N_848,N_1013);
nand U1216 (N_1216,N_1032,N_1071);
and U1217 (N_1217,N_1118,N_742);
nor U1218 (N_1218,N_705,N_887);
nand U1219 (N_1219,N_775,N_954);
nand U1220 (N_1220,N_1152,N_653);
and U1221 (N_1221,N_707,N_1038);
xnor U1222 (N_1222,N_626,N_881);
nand U1223 (N_1223,N_849,N_765);
and U1224 (N_1224,N_733,N_757);
or U1225 (N_1225,N_762,N_992);
xnor U1226 (N_1226,N_885,N_1167);
and U1227 (N_1227,N_1181,N_1019);
and U1228 (N_1228,N_946,N_642);
or U1229 (N_1229,N_684,N_929);
nor U1230 (N_1230,N_1076,N_1045);
and U1231 (N_1231,N_1153,N_884);
nand U1232 (N_1232,N_802,N_857);
and U1233 (N_1233,N_1026,N_867);
nor U1234 (N_1234,N_996,N_970);
nand U1235 (N_1235,N_1033,N_1164);
or U1236 (N_1236,N_795,N_641);
nor U1237 (N_1237,N_1025,N_678);
xor U1238 (N_1238,N_644,N_660);
or U1239 (N_1239,N_815,N_915);
and U1240 (N_1240,N_955,N_753);
or U1241 (N_1241,N_824,N_1146);
and U1242 (N_1242,N_1069,N_783);
and U1243 (N_1243,N_1093,N_865);
xor U1244 (N_1244,N_1168,N_817);
and U1245 (N_1245,N_693,N_1106);
nand U1246 (N_1246,N_902,N_702);
nor U1247 (N_1247,N_1149,N_966);
and U1248 (N_1248,N_667,N_1178);
and U1249 (N_1249,N_1086,N_859);
nand U1250 (N_1250,N_1022,N_1097);
nand U1251 (N_1251,N_1091,N_916);
or U1252 (N_1252,N_1128,N_947);
and U1253 (N_1253,N_629,N_662);
nor U1254 (N_1254,N_889,N_994);
and U1255 (N_1255,N_1092,N_1112);
nand U1256 (N_1256,N_975,N_825);
and U1257 (N_1257,N_784,N_838);
or U1258 (N_1258,N_722,N_716);
or U1259 (N_1259,N_739,N_761);
or U1260 (N_1260,N_1198,N_935);
or U1261 (N_1261,N_949,N_957);
nor U1262 (N_1262,N_974,N_1171);
or U1263 (N_1263,N_1184,N_770);
nand U1264 (N_1264,N_862,N_1132);
nand U1265 (N_1265,N_984,N_646);
or U1266 (N_1266,N_998,N_628);
or U1267 (N_1267,N_615,N_995);
xnor U1268 (N_1268,N_1035,N_1080);
or U1269 (N_1269,N_730,N_688);
nor U1270 (N_1270,N_1039,N_1044);
or U1271 (N_1271,N_976,N_788);
or U1272 (N_1272,N_1048,N_724);
and U1273 (N_1273,N_806,N_792);
and U1274 (N_1274,N_749,N_1084);
nand U1275 (N_1275,N_1111,N_1054);
nor U1276 (N_1276,N_923,N_829);
nor U1277 (N_1277,N_763,N_799);
and U1278 (N_1278,N_797,N_696);
nand U1279 (N_1279,N_987,N_1177);
nor U1280 (N_1280,N_782,N_1162);
nand U1281 (N_1281,N_728,N_1006);
and U1282 (N_1282,N_618,N_936);
or U1283 (N_1283,N_1157,N_771);
nand U1284 (N_1284,N_1159,N_779);
or U1285 (N_1285,N_967,N_1062);
nand U1286 (N_1286,N_969,N_1094);
and U1287 (N_1287,N_1183,N_964);
and U1288 (N_1288,N_1105,N_1108);
and U1289 (N_1289,N_1142,N_1154);
or U1290 (N_1290,N_1075,N_681);
nand U1291 (N_1291,N_1089,N_961);
nor U1292 (N_1292,N_1135,N_1020);
nor U1293 (N_1293,N_842,N_989);
nand U1294 (N_1294,N_639,N_893);
nand U1295 (N_1295,N_700,N_813);
nor U1296 (N_1296,N_719,N_827);
or U1297 (N_1297,N_958,N_1015);
or U1298 (N_1298,N_870,N_1009);
nor U1299 (N_1299,N_883,N_843);
and U1300 (N_1300,N_1139,N_781);
nand U1301 (N_1301,N_927,N_837);
nor U1302 (N_1302,N_1189,N_743);
nor U1303 (N_1303,N_1150,N_951);
nor U1304 (N_1304,N_1070,N_1014);
or U1305 (N_1305,N_971,N_1147);
and U1306 (N_1306,N_1083,N_844);
and U1307 (N_1307,N_1141,N_965);
or U1308 (N_1308,N_942,N_816);
and U1309 (N_1309,N_1095,N_898);
and U1310 (N_1310,N_863,N_773);
nand U1311 (N_1311,N_1156,N_820);
nand U1312 (N_1312,N_841,N_822);
nand U1313 (N_1313,N_745,N_1129);
nor U1314 (N_1314,N_993,N_944);
or U1315 (N_1315,N_875,N_1099);
nor U1316 (N_1316,N_963,N_651);
or U1317 (N_1317,N_752,N_834);
and U1318 (N_1318,N_1031,N_686);
nor U1319 (N_1319,N_1002,N_680);
and U1320 (N_1320,N_868,N_1018);
nor U1321 (N_1321,N_832,N_748);
and U1322 (N_1322,N_909,N_1180);
nand U1323 (N_1323,N_1029,N_830);
and U1324 (N_1324,N_897,N_634);
nor U1325 (N_1325,N_921,N_847);
or U1326 (N_1326,N_741,N_727);
nand U1327 (N_1327,N_637,N_819);
nand U1328 (N_1328,N_731,N_647);
nor U1329 (N_1329,N_712,N_718);
xnor U1330 (N_1330,N_932,N_720);
and U1331 (N_1331,N_791,N_1037);
or U1332 (N_1332,N_1179,N_697);
nor U1333 (N_1333,N_694,N_677);
nor U1334 (N_1334,N_635,N_851);
nand U1335 (N_1335,N_602,N_603);
and U1336 (N_1336,N_988,N_1125);
nor U1337 (N_1337,N_698,N_945);
nand U1338 (N_1338,N_910,N_1074);
nand U1339 (N_1339,N_1034,N_760);
and U1340 (N_1340,N_1163,N_655);
or U1341 (N_1341,N_845,N_1138);
or U1342 (N_1342,N_943,N_650);
and U1343 (N_1343,N_903,N_860);
nor U1344 (N_1344,N_928,N_872);
or U1345 (N_1345,N_1116,N_682);
and U1346 (N_1346,N_803,N_810);
or U1347 (N_1347,N_1043,N_1068);
nor U1348 (N_1348,N_836,N_981);
xor U1349 (N_1349,N_654,N_1098);
or U1350 (N_1350,N_866,N_701);
nor U1351 (N_1351,N_1140,N_1073);
and U1352 (N_1352,N_933,N_1117);
xor U1353 (N_1353,N_941,N_960);
xor U1354 (N_1354,N_1148,N_710);
nor U1355 (N_1355,N_751,N_895);
nor U1356 (N_1356,N_675,N_612);
or U1357 (N_1357,N_1166,N_764);
or U1358 (N_1358,N_892,N_894);
and U1359 (N_1359,N_687,N_699);
or U1360 (N_1360,N_1001,N_1134);
nor U1361 (N_1361,N_768,N_917);
or U1362 (N_1362,N_940,N_1010);
xor U1363 (N_1363,N_798,N_997);
nor U1364 (N_1364,N_1199,N_1110);
nor U1365 (N_1365,N_676,N_664);
nor U1366 (N_1366,N_818,N_1107);
xor U1367 (N_1367,N_977,N_774);
xor U1368 (N_1368,N_619,N_786);
or U1369 (N_1369,N_657,N_1145);
nand U1370 (N_1370,N_918,N_850);
xor U1371 (N_1371,N_1072,N_1079);
nor U1372 (N_1372,N_1155,N_1016);
or U1373 (N_1373,N_609,N_807);
or U1374 (N_1374,N_911,N_715);
or U1375 (N_1375,N_1096,N_1023);
or U1376 (N_1376,N_1017,N_692);
nor U1377 (N_1377,N_756,N_919);
nand U1378 (N_1378,N_1040,N_750);
or U1379 (N_1379,N_890,N_671);
nand U1380 (N_1380,N_789,N_858);
or U1381 (N_1381,N_1182,N_925);
or U1382 (N_1382,N_1126,N_968);
nor U1383 (N_1383,N_601,N_1059);
nand U1384 (N_1384,N_900,N_864);
nand U1385 (N_1385,N_708,N_616);
xnor U1386 (N_1386,N_1165,N_1085);
nor U1387 (N_1387,N_886,N_1161);
nor U1388 (N_1388,N_907,N_922);
nand U1389 (N_1389,N_908,N_980);
and U1390 (N_1390,N_878,N_638);
nor U1391 (N_1391,N_800,N_939);
nor U1392 (N_1392,N_1103,N_1119);
nor U1393 (N_1393,N_906,N_1101);
or U1394 (N_1394,N_645,N_1187);
nor U1395 (N_1395,N_623,N_1194);
nor U1396 (N_1396,N_717,N_611);
and U1397 (N_1397,N_1061,N_882);
or U1398 (N_1398,N_614,N_648);
or U1399 (N_1399,N_621,N_871);
nor U1400 (N_1400,N_833,N_835);
or U1401 (N_1401,N_874,N_778);
and U1402 (N_1402,N_673,N_796);
and U1403 (N_1403,N_901,N_1007);
nand U1404 (N_1404,N_663,N_1053);
nand U1405 (N_1405,N_668,N_1131);
nand U1406 (N_1406,N_904,N_1133);
nand U1407 (N_1407,N_1047,N_656);
nand U1408 (N_1408,N_683,N_605);
nor U1409 (N_1409,N_1090,N_1176);
or U1410 (N_1410,N_658,N_793);
and U1411 (N_1411,N_1008,N_659);
nand U1412 (N_1412,N_772,N_607);
xor U1413 (N_1413,N_1081,N_780);
nand U1414 (N_1414,N_1088,N_734);
or U1415 (N_1415,N_852,N_600);
and U1416 (N_1416,N_812,N_685);
and U1417 (N_1417,N_914,N_861);
and U1418 (N_1418,N_1051,N_880);
nor U1419 (N_1419,N_754,N_608);
nor U1420 (N_1420,N_1003,N_759);
nand U1421 (N_1421,N_876,N_652);
and U1422 (N_1422,N_758,N_990);
or U1423 (N_1423,N_622,N_956);
nand U1424 (N_1424,N_610,N_709);
or U1425 (N_1425,N_747,N_776);
or U1426 (N_1426,N_1082,N_1050);
nand U1427 (N_1427,N_1060,N_1115);
nor U1428 (N_1428,N_736,N_704);
or U1429 (N_1429,N_1056,N_811);
and U1430 (N_1430,N_856,N_855);
and U1431 (N_1431,N_804,N_1065);
xor U1432 (N_1432,N_665,N_672);
nand U1433 (N_1433,N_952,N_1102);
or U1434 (N_1434,N_1077,N_1114);
and U1435 (N_1435,N_627,N_938);
and U1436 (N_1436,N_633,N_986);
and U1437 (N_1437,N_1137,N_613);
or U1438 (N_1438,N_1078,N_1174);
nand U1439 (N_1439,N_643,N_926);
nor U1440 (N_1440,N_726,N_666);
nor U1441 (N_1441,N_979,N_1143);
nand U1442 (N_1442,N_1191,N_735);
or U1443 (N_1443,N_1042,N_959);
xnor U1444 (N_1444,N_1064,N_1197);
nor U1445 (N_1445,N_1046,N_953);
nor U1446 (N_1446,N_713,N_690);
xor U1447 (N_1447,N_808,N_934);
nand U1448 (N_1448,N_669,N_1127);
xnor U1449 (N_1449,N_640,N_1036);
nor U1450 (N_1450,N_1058,N_1021);
nand U1451 (N_1451,N_695,N_1027);
or U1452 (N_1452,N_999,N_1087);
and U1453 (N_1453,N_1122,N_723);
or U1454 (N_1454,N_1192,N_985);
and U1455 (N_1455,N_625,N_630);
nor U1456 (N_1456,N_948,N_1190);
nand U1457 (N_1457,N_679,N_649);
nor U1458 (N_1458,N_1144,N_1113);
or U1459 (N_1459,N_912,N_1193);
and U1460 (N_1460,N_767,N_1012);
nand U1461 (N_1461,N_896,N_814);
nor U1462 (N_1462,N_746,N_809);
and U1463 (N_1463,N_1195,N_950);
nand U1464 (N_1464,N_1041,N_853);
and U1465 (N_1465,N_846,N_905);
nor U1466 (N_1466,N_1123,N_714);
nor U1467 (N_1467,N_732,N_1175);
nand U1468 (N_1468,N_738,N_1158);
and U1469 (N_1469,N_879,N_631);
or U1470 (N_1470,N_766,N_1100);
nand U1471 (N_1471,N_1185,N_777);
nand U1472 (N_1472,N_617,N_805);
nor U1473 (N_1473,N_606,N_1000);
and U1474 (N_1474,N_1120,N_729);
nor U1475 (N_1475,N_978,N_706);
or U1476 (N_1476,N_891,N_873);
nor U1477 (N_1477,N_740,N_1130);
nand U1478 (N_1478,N_899,N_1173);
nand U1479 (N_1479,N_744,N_604);
nor U1480 (N_1480,N_636,N_661);
nand U1481 (N_1481,N_1160,N_632);
or U1482 (N_1482,N_937,N_931);
nor U1483 (N_1483,N_913,N_823);
and U1484 (N_1484,N_828,N_1004);
nand U1485 (N_1485,N_1151,N_1067);
nand U1486 (N_1486,N_737,N_1170);
nor U1487 (N_1487,N_1028,N_1169);
or U1488 (N_1488,N_930,N_1172);
nor U1489 (N_1489,N_801,N_1124);
or U1490 (N_1490,N_1136,N_1109);
xor U1491 (N_1491,N_1024,N_725);
or U1492 (N_1492,N_1052,N_755);
nor U1493 (N_1493,N_620,N_703);
and U1494 (N_1494,N_689,N_982);
nor U1495 (N_1495,N_721,N_1049);
nor U1496 (N_1496,N_1055,N_888);
nand U1497 (N_1497,N_972,N_831);
and U1498 (N_1498,N_920,N_840);
and U1499 (N_1499,N_790,N_973);
nand U1500 (N_1500,N_801,N_661);
or U1501 (N_1501,N_1091,N_1163);
or U1502 (N_1502,N_837,N_1080);
nand U1503 (N_1503,N_1118,N_774);
nand U1504 (N_1504,N_888,N_1123);
or U1505 (N_1505,N_1006,N_1000);
or U1506 (N_1506,N_615,N_982);
xnor U1507 (N_1507,N_1104,N_1129);
nand U1508 (N_1508,N_719,N_1127);
nor U1509 (N_1509,N_1141,N_619);
nor U1510 (N_1510,N_755,N_945);
or U1511 (N_1511,N_935,N_1158);
nand U1512 (N_1512,N_959,N_1074);
xnor U1513 (N_1513,N_1122,N_979);
xnor U1514 (N_1514,N_1063,N_736);
nor U1515 (N_1515,N_966,N_941);
and U1516 (N_1516,N_937,N_670);
nand U1517 (N_1517,N_1160,N_936);
and U1518 (N_1518,N_1024,N_776);
nand U1519 (N_1519,N_980,N_841);
nand U1520 (N_1520,N_1074,N_678);
or U1521 (N_1521,N_1114,N_840);
nor U1522 (N_1522,N_997,N_1160);
xnor U1523 (N_1523,N_901,N_768);
or U1524 (N_1524,N_1074,N_842);
and U1525 (N_1525,N_917,N_1184);
nand U1526 (N_1526,N_1055,N_766);
and U1527 (N_1527,N_607,N_1018);
nand U1528 (N_1528,N_894,N_865);
xnor U1529 (N_1529,N_667,N_1166);
nand U1530 (N_1530,N_894,N_1159);
or U1531 (N_1531,N_894,N_982);
and U1532 (N_1532,N_673,N_788);
or U1533 (N_1533,N_617,N_716);
xnor U1534 (N_1534,N_1027,N_1107);
and U1535 (N_1535,N_627,N_975);
nor U1536 (N_1536,N_1101,N_1070);
nand U1537 (N_1537,N_1179,N_864);
or U1538 (N_1538,N_825,N_746);
nor U1539 (N_1539,N_622,N_909);
and U1540 (N_1540,N_877,N_873);
nand U1541 (N_1541,N_1109,N_794);
and U1542 (N_1542,N_762,N_783);
nand U1543 (N_1543,N_1064,N_609);
xnor U1544 (N_1544,N_1114,N_1165);
or U1545 (N_1545,N_872,N_947);
xor U1546 (N_1546,N_1069,N_885);
and U1547 (N_1547,N_838,N_1125);
or U1548 (N_1548,N_1110,N_999);
nand U1549 (N_1549,N_1134,N_987);
nor U1550 (N_1550,N_938,N_846);
nand U1551 (N_1551,N_707,N_914);
xnor U1552 (N_1552,N_1085,N_1127);
nor U1553 (N_1553,N_1131,N_824);
or U1554 (N_1554,N_804,N_1109);
and U1555 (N_1555,N_874,N_791);
nor U1556 (N_1556,N_670,N_941);
nand U1557 (N_1557,N_1195,N_915);
nand U1558 (N_1558,N_1026,N_1116);
nand U1559 (N_1559,N_1186,N_737);
nand U1560 (N_1560,N_666,N_894);
nor U1561 (N_1561,N_790,N_901);
nor U1562 (N_1562,N_891,N_1037);
or U1563 (N_1563,N_1077,N_988);
or U1564 (N_1564,N_814,N_684);
nor U1565 (N_1565,N_981,N_890);
nor U1566 (N_1566,N_1016,N_1162);
or U1567 (N_1567,N_1147,N_900);
nand U1568 (N_1568,N_1135,N_608);
xor U1569 (N_1569,N_859,N_763);
xnor U1570 (N_1570,N_1093,N_1100);
nor U1571 (N_1571,N_1118,N_1124);
or U1572 (N_1572,N_882,N_1179);
nand U1573 (N_1573,N_826,N_1000);
and U1574 (N_1574,N_659,N_767);
xor U1575 (N_1575,N_882,N_1147);
nor U1576 (N_1576,N_938,N_1189);
nand U1577 (N_1577,N_1041,N_804);
xnor U1578 (N_1578,N_797,N_1039);
nor U1579 (N_1579,N_953,N_1166);
and U1580 (N_1580,N_810,N_988);
or U1581 (N_1581,N_853,N_724);
or U1582 (N_1582,N_1144,N_1072);
nor U1583 (N_1583,N_790,N_971);
or U1584 (N_1584,N_1193,N_898);
xor U1585 (N_1585,N_1009,N_662);
and U1586 (N_1586,N_985,N_674);
and U1587 (N_1587,N_863,N_1051);
nand U1588 (N_1588,N_1075,N_1086);
or U1589 (N_1589,N_952,N_1176);
and U1590 (N_1590,N_1083,N_867);
or U1591 (N_1591,N_993,N_1140);
and U1592 (N_1592,N_798,N_686);
nand U1593 (N_1593,N_816,N_1000);
and U1594 (N_1594,N_614,N_782);
and U1595 (N_1595,N_1164,N_780);
or U1596 (N_1596,N_672,N_1088);
nand U1597 (N_1597,N_649,N_891);
and U1598 (N_1598,N_910,N_1032);
and U1599 (N_1599,N_669,N_1135);
nor U1600 (N_1600,N_885,N_777);
xnor U1601 (N_1601,N_1178,N_1028);
and U1602 (N_1602,N_1034,N_924);
or U1603 (N_1603,N_903,N_1122);
nand U1604 (N_1604,N_906,N_1126);
xnor U1605 (N_1605,N_758,N_1085);
or U1606 (N_1606,N_1076,N_745);
and U1607 (N_1607,N_1074,N_1118);
nand U1608 (N_1608,N_932,N_1117);
and U1609 (N_1609,N_624,N_1171);
nand U1610 (N_1610,N_969,N_1160);
nor U1611 (N_1611,N_746,N_1135);
nor U1612 (N_1612,N_684,N_1029);
nor U1613 (N_1613,N_1162,N_1021);
nand U1614 (N_1614,N_1093,N_1120);
and U1615 (N_1615,N_1092,N_954);
nor U1616 (N_1616,N_688,N_610);
nor U1617 (N_1617,N_1105,N_724);
nand U1618 (N_1618,N_1170,N_1044);
xor U1619 (N_1619,N_868,N_1078);
nand U1620 (N_1620,N_1005,N_795);
or U1621 (N_1621,N_924,N_972);
nor U1622 (N_1622,N_696,N_1061);
and U1623 (N_1623,N_920,N_874);
nor U1624 (N_1624,N_672,N_912);
nand U1625 (N_1625,N_757,N_1175);
and U1626 (N_1626,N_969,N_820);
nor U1627 (N_1627,N_691,N_1121);
or U1628 (N_1628,N_1070,N_1168);
or U1629 (N_1629,N_934,N_1120);
nor U1630 (N_1630,N_788,N_683);
nor U1631 (N_1631,N_812,N_1055);
nand U1632 (N_1632,N_1175,N_885);
nand U1633 (N_1633,N_1018,N_899);
nand U1634 (N_1634,N_983,N_682);
nor U1635 (N_1635,N_692,N_1028);
nand U1636 (N_1636,N_685,N_873);
nor U1637 (N_1637,N_1197,N_964);
or U1638 (N_1638,N_996,N_604);
nor U1639 (N_1639,N_1073,N_1100);
nor U1640 (N_1640,N_1153,N_1010);
and U1641 (N_1641,N_1034,N_861);
nor U1642 (N_1642,N_902,N_774);
nor U1643 (N_1643,N_810,N_668);
nand U1644 (N_1644,N_721,N_1056);
nor U1645 (N_1645,N_1166,N_982);
or U1646 (N_1646,N_729,N_926);
nor U1647 (N_1647,N_843,N_1192);
or U1648 (N_1648,N_705,N_1041);
nor U1649 (N_1649,N_682,N_873);
or U1650 (N_1650,N_1097,N_670);
nor U1651 (N_1651,N_828,N_650);
nor U1652 (N_1652,N_634,N_761);
xnor U1653 (N_1653,N_725,N_991);
or U1654 (N_1654,N_653,N_804);
or U1655 (N_1655,N_839,N_990);
xnor U1656 (N_1656,N_856,N_1183);
nand U1657 (N_1657,N_1139,N_601);
nor U1658 (N_1658,N_770,N_812);
nor U1659 (N_1659,N_854,N_1176);
nand U1660 (N_1660,N_948,N_739);
nor U1661 (N_1661,N_771,N_1073);
and U1662 (N_1662,N_1116,N_804);
nor U1663 (N_1663,N_1063,N_641);
nand U1664 (N_1664,N_925,N_776);
nor U1665 (N_1665,N_955,N_606);
nand U1666 (N_1666,N_1029,N_716);
nand U1667 (N_1667,N_815,N_816);
and U1668 (N_1668,N_903,N_619);
and U1669 (N_1669,N_739,N_968);
nor U1670 (N_1670,N_746,N_1042);
or U1671 (N_1671,N_855,N_866);
and U1672 (N_1672,N_798,N_711);
or U1673 (N_1673,N_910,N_600);
nand U1674 (N_1674,N_1110,N_603);
nor U1675 (N_1675,N_615,N_813);
nor U1676 (N_1676,N_1102,N_1017);
nor U1677 (N_1677,N_757,N_702);
nand U1678 (N_1678,N_1106,N_622);
nor U1679 (N_1679,N_1171,N_648);
and U1680 (N_1680,N_963,N_765);
and U1681 (N_1681,N_858,N_1143);
and U1682 (N_1682,N_949,N_985);
nand U1683 (N_1683,N_707,N_603);
and U1684 (N_1684,N_819,N_607);
and U1685 (N_1685,N_832,N_762);
nor U1686 (N_1686,N_1075,N_992);
nand U1687 (N_1687,N_882,N_683);
or U1688 (N_1688,N_1180,N_900);
nand U1689 (N_1689,N_1035,N_646);
nor U1690 (N_1690,N_979,N_1171);
and U1691 (N_1691,N_951,N_831);
nand U1692 (N_1692,N_854,N_921);
nor U1693 (N_1693,N_766,N_1197);
nor U1694 (N_1694,N_1119,N_1166);
nor U1695 (N_1695,N_1064,N_604);
and U1696 (N_1696,N_754,N_824);
and U1697 (N_1697,N_994,N_606);
or U1698 (N_1698,N_726,N_1172);
nor U1699 (N_1699,N_960,N_888);
nand U1700 (N_1700,N_1071,N_1168);
nor U1701 (N_1701,N_849,N_965);
or U1702 (N_1702,N_1102,N_1064);
or U1703 (N_1703,N_972,N_1015);
nand U1704 (N_1704,N_786,N_799);
nor U1705 (N_1705,N_771,N_813);
nor U1706 (N_1706,N_1192,N_1005);
nand U1707 (N_1707,N_998,N_999);
xnor U1708 (N_1708,N_1188,N_981);
and U1709 (N_1709,N_695,N_764);
or U1710 (N_1710,N_905,N_921);
nand U1711 (N_1711,N_1022,N_788);
and U1712 (N_1712,N_955,N_1043);
nand U1713 (N_1713,N_1123,N_663);
and U1714 (N_1714,N_1083,N_921);
nand U1715 (N_1715,N_1016,N_940);
and U1716 (N_1716,N_951,N_953);
and U1717 (N_1717,N_979,N_848);
or U1718 (N_1718,N_687,N_1029);
or U1719 (N_1719,N_1117,N_920);
xor U1720 (N_1720,N_983,N_817);
nand U1721 (N_1721,N_1177,N_1159);
and U1722 (N_1722,N_922,N_652);
and U1723 (N_1723,N_641,N_874);
and U1724 (N_1724,N_877,N_783);
nand U1725 (N_1725,N_602,N_709);
nand U1726 (N_1726,N_721,N_739);
nand U1727 (N_1727,N_669,N_702);
and U1728 (N_1728,N_787,N_758);
and U1729 (N_1729,N_632,N_1116);
nor U1730 (N_1730,N_1114,N_704);
or U1731 (N_1731,N_911,N_1111);
nand U1732 (N_1732,N_759,N_1048);
or U1733 (N_1733,N_915,N_1196);
or U1734 (N_1734,N_1064,N_672);
and U1735 (N_1735,N_613,N_674);
and U1736 (N_1736,N_993,N_758);
nand U1737 (N_1737,N_932,N_971);
or U1738 (N_1738,N_895,N_1017);
xnor U1739 (N_1739,N_662,N_794);
and U1740 (N_1740,N_680,N_815);
nor U1741 (N_1741,N_609,N_1114);
nand U1742 (N_1742,N_920,N_753);
nand U1743 (N_1743,N_1093,N_1062);
nor U1744 (N_1744,N_710,N_748);
xor U1745 (N_1745,N_635,N_926);
nand U1746 (N_1746,N_1139,N_722);
nor U1747 (N_1747,N_1120,N_1007);
or U1748 (N_1748,N_998,N_1134);
or U1749 (N_1749,N_1102,N_714);
and U1750 (N_1750,N_833,N_610);
nand U1751 (N_1751,N_812,N_806);
nor U1752 (N_1752,N_1032,N_663);
nand U1753 (N_1753,N_858,N_771);
nor U1754 (N_1754,N_1004,N_1137);
xor U1755 (N_1755,N_1009,N_1077);
or U1756 (N_1756,N_986,N_859);
nor U1757 (N_1757,N_875,N_846);
or U1758 (N_1758,N_801,N_602);
xor U1759 (N_1759,N_1181,N_1008);
nor U1760 (N_1760,N_1183,N_1182);
nand U1761 (N_1761,N_724,N_1006);
or U1762 (N_1762,N_758,N_714);
nor U1763 (N_1763,N_806,N_1102);
xor U1764 (N_1764,N_1187,N_608);
and U1765 (N_1765,N_771,N_1045);
and U1766 (N_1766,N_641,N_606);
and U1767 (N_1767,N_1084,N_772);
or U1768 (N_1768,N_905,N_747);
xnor U1769 (N_1769,N_1053,N_919);
or U1770 (N_1770,N_769,N_1084);
and U1771 (N_1771,N_708,N_735);
and U1772 (N_1772,N_693,N_1152);
and U1773 (N_1773,N_1043,N_764);
or U1774 (N_1774,N_1166,N_779);
or U1775 (N_1775,N_622,N_831);
nor U1776 (N_1776,N_805,N_1080);
nor U1777 (N_1777,N_863,N_1082);
or U1778 (N_1778,N_993,N_690);
and U1779 (N_1779,N_883,N_1023);
and U1780 (N_1780,N_743,N_1168);
nor U1781 (N_1781,N_1092,N_668);
nor U1782 (N_1782,N_874,N_783);
xnor U1783 (N_1783,N_762,N_734);
nor U1784 (N_1784,N_1126,N_705);
nand U1785 (N_1785,N_1154,N_707);
and U1786 (N_1786,N_998,N_927);
nor U1787 (N_1787,N_658,N_903);
and U1788 (N_1788,N_647,N_1161);
or U1789 (N_1789,N_1006,N_764);
and U1790 (N_1790,N_1085,N_865);
or U1791 (N_1791,N_1104,N_1185);
or U1792 (N_1792,N_1080,N_734);
nand U1793 (N_1793,N_973,N_707);
nor U1794 (N_1794,N_840,N_631);
nand U1795 (N_1795,N_1068,N_655);
and U1796 (N_1796,N_714,N_730);
xnor U1797 (N_1797,N_1059,N_683);
and U1798 (N_1798,N_658,N_770);
xnor U1799 (N_1799,N_786,N_1194);
or U1800 (N_1800,N_1323,N_1468);
nor U1801 (N_1801,N_1303,N_1219);
and U1802 (N_1802,N_1593,N_1212);
nor U1803 (N_1803,N_1719,N_1714);
and U1804 (N_1804,N_1704,N_1353);
nor U1805 (N_1805,N_1239,N_1292);
nor U1806 (N_1806,N_1206,N_1531);
nand U1807 (N_1807,N_1545,N_1419);
xnor U1808 (N_1808,N_1508,N_1474);
nand U1809 (N_1809,N_1767,N_1382);
xor U1810 (N_1810,N_1305,N_1499);
or U1811 (N_1811,N_1253,N_1678);
nand U1812 (N_1812,N_1698,N_1534);
nand U1813 (N_1813,N_1222,N_1426);
or U1814 (N_1814,N_1481,N_1682);
nand U1815 (N_1815,N_1715,N_1590);
or U1816 (N_1816,N_1317,N_1777);
and U1817 (N_1817,N_1209,N_1226);
xnor U1818 (N_1818,N_1725,N_1575);
nand U1819 (N_1819,N_1307,N_1768);
and U1820 (N_1820,N_1797,N_1446);
and U1821 (N_1821,N_1564,N_1556);
nor U1822 (N_1822,N_1223,N_1410);
nand U1823 (N_1823,N_1256,N_1211);
and U1824 (N_1824,N_1731,N_1229);
nor U1825 (N_1825,N_1670,N_1782);
and U1826 (N_1826,N_1755,N_1561);
or U1827 (N_1827,N_1739,N_1512);
and U1828 (N_1828,N_1260,N_1763);
nor U1829 (N_1829,N_1627,N_1537);
nor U1830 (N_1830,N_1663,N_1326);
and U1831 (N_1831,N_1742,N_1337);
and U1832 (N_1832,N_1503,N_1553);
and U1833 (N_1833,N_1334,N_1373);
or U1834 (N_1834,N_1313,N_1336);
xnor U1835 (N_1835,N_1362,N_1559);
nand U1836 (N_1836,N_1280,N_1366);
nor U1837 (N_1837,N_1751,N_1683);
or U1838 (N_1838,N_1467,N_1754);
nand U1839 (N_1839,N_1721,N_1412);
or U1840 (N_1840,N_1498,N_1210);
and U1841 (N_1841,N_1708,N_1315);
or U1842 (N_1842,N_1737,N_1271);
nor U1843 (N_1843,N_1230,N_1519);
nor U1844 (N_1844,N_1579,N_1557);
nor U1845 (N_1845,N_1729,N_1732);
and U1846 (N_1846,N_1378,N_1504);
and U1847 (N_1847,N_1584,N_1756);
and U1848 (N_1848,N_1706,N_1447);
nor U1849 (N_1849,N_1327,N_1527);
nand U1850 (N_1850,N_1322,N_1591);
and U1851 (N_1851,N_1248,N_1486);
xnor U1852 (N_1852,N_1651,N_1655);
nand U1853 (N_1853,N_1453,N_1371);
xnor U1854 (N_1854,N_1726,N_1489);
nand U1855 (N_1855,N_1513,N_1781);
nand U1856 (N_1856,N_1775,N_1300);
nand U1857 (N_1857,N_1638,N_1705);
and U1858 (N_1858,N_1532,N_1455);
and U1859 (N_1859,N_1623,N_1214);
or U1860 (N_1860,N_1244,N_1381);
and U1861 (N_1861,N_1662,N_1743);
nand U1862 (N_1862,N_1372,N_1771);
and U1863 (N_1863,N_1398,N_1505);
or U1864 (N_1864,N_1367,N_1783);
nor U1865 (N_1865,N_1484,N_1434);
nand U1866 (N_1866,N_1785,N_1583);
nand U1867 (N_1867,N_1409,N_1476);
and U1868 (N_1868,N_1680,N_1444);
or U1869 (N_1869,N_1351,N_1243);
nand U1870 (N_1870,N_1535,N_1495);
nand U1871 (N_1871,N_1795,N_1776);
xor U1872 (N_1872,N_1369,N_1414);
nand U1873 (N_1873,N_1297,N_1363);
nand U1874 (N_1874,N_1483,N_1437);
nand U1875 (N_1875,N_1450,N_1740);
or U1876 (N_1876,N_1541,N_1749);
nor U1877 (N_1877,N_1786,N_1270);
nor U1878 (N_1878,N_1202,N_1462);
and U1879 (N_1879,N_1261,N_1760);
nand U1880 (N_1880,N_1666,N_1547);
nand U1881 (N_1881,N_1452,N_1659);
or U1882 (N_1882,N_1676,N_1458);
nor U1883 (N_1883,N_1496,N_1386);
xor U1884 (N_1884,N_1562,N_1360);
nor U1885 (N_1885,N_1594,N_1511);
or U1886 (N_1886,N_1718,N_1459);
nand U1887 (N_1887,N_1478,N_1710);
nand U1888 (N_1888,N_1546,N_1679);
nand U1889 (N_1889,N_1661,N_1449);
xor U1890 (N_1890,N_1791,N_1293);
xor U1891 (N_1891,N_1276,N_1424);
nand U1892 (N_1892,N_1330,N_1431);
xnor U1893 (N_1893,N_1473,N_1724);
nand U1894 (N_1894,N_1430,N_1636);
nor U1895 (N_1895,N_1611,N_1766);
nor U1896 (N_1896,N_1578,N_1521);
nor U1897 (N_1897,N_1649,N_1626);
nand U1898 (N_1898,N_1275,N_1668);
and U1899 (N_1899,N_1707,N_1722);
nand U1900 (N_1900,N_1543,N_1418);
or U1901 (N_1901,N_1341,N_1701);
or U1902 (N_1902,N_1475,N_1648);
nor U1903 (N_1903,N_1520,N_1402);
nor U1904 (N_1904,N_1405,N_1238);
xnor U1905 (N_1905,N_1650,N_1298);
nor U1906 (N_1906,N_1657,N_1457);
and U1907 (N_1907,N_1227,N_1263);
and U1908 (N_1908,N_1438,N_1370);
and U1909 (N_1909,N_1355,N_1538);
nand U1910 (N_1910,N_1262,N_1234);
nor U1911 (N_1911,N_1577,N_1314);
or U1912 (N_1912,N_1340,N_1279);
or U1913 (N_1913,N_1441,N_1773);
and U1914 (N_1914,N_1586,N_1616);
nand U1915 (N_1915,N_1778,N_1712);
nand U1916 (N_1916,N_1493,N_1342);
and U1917 (N_1917,N_1357,N_1388);
or U1918 (N_1918,N_1730,N_1460);
and U1919 (N_1919,N_1607,N_1617);
or U1920 (N_1920,N_1569,N_1632);
and U1921 (N_1921,N_1612,N_1788);
or U1922 (N_1922,N_1633,N_1745);
nor U1923 (N_1923,N_1523,N_1242);
nand U1924 (N_1924,N_1560,N_1479);
nor U1925 (N_1925,N_1554,N_1637);
nor U1926 (N_1926,N_1377,N_1762);
nand U1927 (N_1927,N_1660,N_1390);
nand U1928 (N_1928,N_1602,N_1671);
nand U1929 (N_1929,N_1765,N_1618);
nor U1930 (N_1930,N_1622,N_1203);
nand U1931 (N_1931,N_1752,N_1325);
nor U1932 (N_1932,N_1673,N_1551);
and U1933 (N_1933,N_1364,N_1779);
and U1934 (N_1934,N_1379,N_1759);
and U1935 (N_1935,N_1416,N_1272);
and U1936 (N_1936,N_1522,N_1425);
xor U1937 (N_1937,N_1393,N_1385);
nand U1938 (N_1938,N_1615,N_1658);
nand U1939 (N_1939,N_1613,N_1524);
and U1940 (N_1940,N_1744,N_1231);
and U1941 (N_1941,N_1610,N_1669);
or U1942 (N_1942,N_1422,N_1290);
nor U1943 (N_1943,N_1343,N_1757);
or U1944 (N_1944,N_1589,N_1235);
xnor U1945 (N_1945,N_1713,N_1601);
nand U1946 (N_1946,N_1396,N_1792);
nand U1947 (N_1947,N_1686,N_1251);
nand U1948 (N_1948,N_1585,N_1690);
or U1949 (N_1949,N_1687,N_1558);
and U1950 (N_1950,N_1443,N_1772);
or U1951 (N_1951,N_1536,N_1699);
nor U1952 (N_1952,N_1681,N_1753);
nor U1953 (N_1953,N_1354,N_1790);
nand U1954 (N_1954,N_1491,N_1580);
and U1955 (N_1955,N_1224,N_1345);
nor U1956 (N_1956,N_1406,N_1324);
nand U1957 (N_1957,N_1750,N_1482);
nand U1958 (N_1958,N_1494,N_1304);
nand U1959 (N_1959,N_1735,N_1514);
nand U1960 (N_1960,N_1727,N_1605);
or U1961 (N_1961,N_1429,N_1629);
xor U1962 (N_1962,N_1287,N_1692);
nor U1963 (N_1963,N_1549,N_1625);
nand U1964 (N_1964,N_1634,N_1654);
nand U1965 (N_1965,N_1228,N_1728);
or U1966 (N_1966,N_1201,N_1647);
nand U1967 (N_1967,N_1675,N_1758);
xnor U1968 (N_1968,N_1335,N_1321);
nand U1969 (N_1969,N_1338,N_1597);
and U1970 (N_1970,N_1672,N_1525);
nand U1971 (N_1971,N_1273,N_1774);
and U1972 (N_1972,N_1507,N_1665);
nand U1973 (N_1973,N_1208,N_1497);
nand U1974 (N_1974,N_1247,N_1588);
xnor U1975 (N_1975,N_1267,N_1375);
and U1976 (N_1976,N_1288,N_1245);
nor U1977 (N_1977,N_1466,N_1320);
or U1978 (N_1978,N_1352,N_1282);
or U1979 (N_1979,N_1492,N_1696);
and U1980 (N_1980,N_1448,N_1299);
or U1981 (N_1981,N_1472,N_1582);
nand U1982 (N_1982,N_1308,N_1454);
nand U1983 (N_1983,N_1463,N_1542);
or U1984 (N_1984,N_1787,N_1257);
and U1985 (N_1985,N_1316,N_1281);
or U1986 (N_1986,N_1347,N_1798);
nor U1987 (N_1987,N_1358,N_1480);
nor U1988 (N_1988,N_1384,N_1769);
or U1989 (N_1989,N_1506,N_1296);
and U1990 (N_1990,N_1677,N_1796);
or U1991 (N_1991,N_1359,N_1394);
nor U1992 (N_1992,N_1286,N_1278);
and U1993 (N_1993,N_1574,N_1249);
and U1994 (N_1994,N_1509,N_1421);
xnor U1995 (N_1995,N_1642,N_1391);
and U1996 (N_1996,N_1259,N_1411);
and U1997 (N_1997,N_1723,N_1387);
nand U1998 (N_1998,N_1641,N_1417);
and U1999 (N_1999,N_1487,N_1456);
nor U2000 (N_2000,N_1310,N_1596);
nand U2001 (N_2001,N_1439,N_1770);
nand U2002 (N_2002,N_1709,N_1311);
nor U2003 (N_2003,N_1664,N_1397);
nor U2004 (N_2004,N_1530,N_1603);
nor U2005 (N_2005,N_1252,N_1552);
nor U2006 (N_2006,N_1399,N_1436);
or U2007 (N_2007,N_1312,N_1628);
nand U2008 (N_2008,N_1599,N_1268);
nand U2009 (N_2009,N_1218,N_1216);
or U2010 (N_2010,N_1517,N_1794);
nor U2011 (N_2011,N_1277,N_1433);
nand U2012 (N_2012,N_1695,N_1741);
and U2013 (N_2013,N_1350,N_1274);
and U2014 (N_2014,N_1600,N_1395);
nor U2015 (N_2015,N_1265,N_1652);
and U2016 (N_2016,N_1368,N_1464);
or U2017 (N_2017,N_1736,N_1346);
nor U2018 (N_2018,N_1383,N_1415);
nand U2019 (N_2019,N_1331,N_1734);
nand U2020 (N_2020,N_1501,N_1403);
xor U2021 (N_2021,N_1285,N_1747);
and U2022 (N_2022,N_1258,N_1780);
or U2023 (N_2023,N_1576,N_1392);
xnor U2024 (N_2024,N_1717,N_1689);
or U2025 (N_2025,N_1428,N_1624);
or U2026 (N_2026,N_1619,N_1643);
and U2027 (N_2027,N_1309,N_1236);
xnor U2028 (N_2028,N_1469,N_1306);
and U2029 (N_2029,N_1356,N_1215);
and U2030 (N_2030,N_1573,N_1207);
xor U2031 (N_2031,N_1205,N_1233);
nand U2032 (N_2032,N_1488,N_1301);
nand U2033 (N_2033,N_1400,N_1241);
nand U2034 (N_2034,N_1614,N_1528);
or U2035 (N_2035,N_1567,N_1328);
nand U2036 (N_2036,N_1471,N_1420);
nand U2037 (N_2037,N_1571,N_1639);
and U2038 (N_2038,N_1461,N_1711);
or U2039 (N_2039,N_1339,N_1269);
or U2040 (N_2040,N_1684,N_1606);
and U2041 (N_2041,N_1240,N_1451);
xnor U2042 (N_2042,N_1568,N_1595);
nor U2043 (N_2043,N_1380,N_1635);
or U2044 (N_2044,N_1544,N_1349);
nand U2045 (N_2045,N_1477,N_1365);
and U2046 (N_2046,N_1685,N_1609);
nor U2047 (N_2047,N_1516,N_1700);
xor U2048 (N_2048,N_1200,N_1413);
xor U2049 (N_2049,N_1592,N_1720);
nand U2050 (N_2050,N_1702,N_1329);
nor U2051 (N_2051,N_1319,N_1254);
and U2052 (N_2052,N_1550,N_1548);
nand U2053 (N_2053,N_1738,N_1716);
nor U2054 (N_2054,N_1407,N_1529);
nor U2055 (N_2055,N_1748,N_1799);
nor U2056 (N_2056,N_1237,N_1295);
nand U2057 (N_2057,N_1656,N_1217);
nand U2058 (N_2058,N_1318,N_1691);
nor U2059 (N_2059,N_1440,N_1401);
or U2060 (N_2060,N_1733,N_1502);
and U2061 (N_2061,N_1572,N_1789);
nand U2062 (N_2062,N_1255,N_1630);
nand U2063 (N_2063,N_1674,N_1565);
or U2064 (N_2064,N_1566,N_1374);
and U2065 (N_2065,N_1640,N_1500);
and U2066 (N_2066,N_1621,N_1423);
and U2067 (N_2067,N_1348,N_1526);
and U2068 (N_2068,N_1221,N_1465);
nand U2069 (N_2069,N_1703,N_1264);
and U2070 (N_2070,N_1570,N_1246);
nand U2071 (N_2071,N_1344,N_1225);
or U2072 (N_2072,N_1563,N_1442);
nor U2073 (N_2073,N_1631,N_1485);
or U2074 (N_2074,N_1213,N_1250);
and U2075 (N_2075,N_1539,N_1784);
or U2076 (N_2076,N_1220,N_1555);
nor U2077 (N_2077,N_1694,N_1510);
or U2078 (N_2078,N_1266,N_1404);
nand U2079 (N_2079,N_1435,N_1291);
or U2080 (N_2080,N_1302,N_1333);
nor U2081 (N_2081,N_1620,N_1515);
or U2082 (N_2082,N_1232,N_1540);
xnor U2083 (N_2083,N_1289,N_1693);
and U2084 (N_2084,N_1389,N_1646);
xnor U2085 (N_2085,N_1688,N_1533);
nor U2086 (N_2086,N_1332,N_1361);
nor U2087 (N_2087,N_1667,N_1294);
nand U2088 (N_2088,N_1490,N_1518);
or U2089 (N_2089,N_1283,N_1697);
or U2090 (N_2090,N_1427,N_1645);
nand U2091 (N_2091,N_1284,N_1445);
and U2092 (N_2092,N_1764,N_1432);
and U2093 (N_2093,N_1204,N_1587);
or U2094 (N_2094,N_1581,N_1793);
nand U2095 (N_2095,N_1470,N_1598);
and U2096 (N_2096,N_1376,N_1604);
nor U2097 (N_2097,N_1746,N_1761);
or U2098 (N_2098,N_1408,N_1653);
nand U2099 (N_2099,N_1608,N_1644);
xor U2100 (N_2100,N_1529,N_1787);
nor U2101 (N_2101,N_1443,N_1329);
nor U2102 (N_2102,N_1203,N_1746);
nor U2103 (N_2103,N_1769,N_1332);
or U2104 (N_2104,N_1708,N_1665);
and U2105 (N_2105,N_1729,N_1416);
xnor U2106 (N_2106,N_1331,N_1345);
and U2107 (N_2107,N_1665,N_1223);
nor U2108 (N_2108,N_1205,N_1404);
xor U2109 (N_2109,N_1639,N_1664);
and U2110 (N_2110,N_1235,N_1704);
nor U2111 (N_2111,N_1541,N_1306);
xor U2112 (N_2112,N_1450,N_1663);
nand U2113 (N_2113,N_1496,N_1632);
or U2114 (N_2114,N_1484,N_1753);
nand U2115 (N_2115,N_1380,N_1422);
and U2116 (N_2116,N_1502,N_1633);
or U2117 (N_2117,N_1729,N_1780);
and U2118 (N_2118,N_1315,N_1631);
nor U2119 (N_2119,N_1585,N_1376);
nor U2120 (N_2120,N_1763,N_1371);
and U2121 (N_2121,N_1266,N_1405);
nand U2122 (N_2122,N_1710,N_1664);
nand U2123 (N_2123,N_1261,N_1354);
nor U2124 (N_2124,N_1572,N_1544);
nor U2125 (N_2125,N_1585,N_1295);
and U2126 (N_2126,N_1743,N_1465);
or U2127 (N_2127,N_1555,N_1381);
or U2128 (N_2128,N_1753,N_1607);
nor U2129 (N_2129,N_1764,N_1666);
nor U2130 (N_2130,N_1554,N_1346);
nor U2131 (N_2131,N_1407,N_1557);
nor U2132 (N_2132,N_1514,N_1609);
and U2133 (N_2133,N_1284,N_1486);
nor U2134 (N_2134,N_1583,N_1362);
nor U2135 (N_2135,N_1318,N_1629);
nand U2136 (N_2136,N_1596,N_1642);
and U2137 (N_2137,N_1479,N_1499);
nand U2138 (N_2138,N_1208,N_1692);
nor U2139 (N_2139,N_1254,N_1205);
and U2140 (N_2140,N_1788,N_1390);
or U2141 (N_2141,N_1716,N_1379);
nand U2142 (N_2142,N_1460,N_1646);
or U2143 (N_2143,N_1704,N_1552);
or U2144 (N_2144,N_1539,N_1702);
and U2145 (N_2145,N_1698,N_1689);
xor U2146 (N_2146,N_1621,N_1321);
nor U2147 (N_2147,N_1543,N_1730);
nor U2148 (N_2148,N_1216,N_1572);
xor U2149 (N_2149,N_1750,N_1245);
nor U2150 (N_2150,N_1245,N_1793);
and U2151 (N_2151,N_1237,N_1266);
nor U2152 (N_2152,N_1643,N_1699);
or U2153 (N_2153,N_1749,N_1373);
or U2154 (N_2154,N_1306,N_1571);
nand U2155 (N_2155,N_1590,N_1297);
or U2156 (N_2156,N_1692,N_1219);
nand U2157 (N_2157,N_1356,N_1507);
or U2158 (N_2158,N_1498,N_1478);
nor U2159 (N_2159,N_1644,N_1220);
nor U2160 (N_2160,N_1223,N_1560);
nor U2161 (N_2161,N_1397,N_1565);
nand U2162 (N_2162,N_1406,N_1299);
nor U2163 (N_2163,N_1412,N_1331);
or U2164 (N_2164,N_1439,N_1535);
nor U2165 (N_2165,N_1355,N_1676);
nor U2166 (N_2166,N_1584,N_1275);
nand U2167 (N_2167,N_1777,N_1632);
and U2168 (N_2168,N_1522,N_1765);
xor U2169 (N_2169,N_1361,N_1388);
nor U2170 (N_2170,N_1270,N_1791);
nand U2171 (N_2171,N_1502,N_1215);
or U2172 (N_2172,N_1686,N_1512);
nor U2173 (N_2173,N_1624,N_1336);
nand U2174 (N_2174,N_1272,N_1539);
xnor U2175 (N_2175,N_1398,N_1485);
and U2176 (N_2176,N_1288,N_1388);
nand U2177 (N_2177,N_1473,N_1680);
nand U2178 (N_2178,N_1487,N_1392);
and U2179 (N_2179,N_1508,N_1599);
and U2180 (N_2180,N_1492,N_1672);
and U2181 (N_2181,N_1795,N_1503);
and U2182 (N_2182,N_1525,N_1200);
nand U2183 (N_2183,N_1383,N_1755);
nand U2184 (N_2184,N_1761,N_1432);
and U2185 (N_2185,N_1621,N_1786);
nand U2186 (N_2186,N_1448,N_1370);
and U2187 (N_2187,N_1432,N_1780);
or U2188 (N_2188,N_1442,N_1784);
nor U2189 (N_2189,N_1251,N_1262);
nor U2190 (N_2190,N_1489,N_1648);
nor U2191 (N_2191,N_1384,N_1221);
nor U2192 (N_2192,N_1363,N_1621);
or U2193 (N_2193,N_1531,N_1731);
or U2194 (N_2194,N_1430,N_1484);
and U2195 (N_2195,N_1494,N_1799);
or U2196 (N_2196,N_1487,N_1734);
and U2197 (N_2197,N_1377,N_1281);
or U2198 (N_2198,N_1722,N_1674);
or U2199 (N_2199,N_1349,N_1606);
nor U2200 (N_2200,N_1331,N_1532);
nand U2201 (N_2201,N_1546,N_1755);
nor U2202 (N_2202,N_1467,N_1755);
and U2203 (N_2203,N_1551,N_1338);
nand U2204 (N_2204,N_1610,N_1412);
xnor U2205 (N_2205,N_1241,N_1788);
nor U2206 (N_2206,N_1214,N_1279);
and U2207 (N_2207,N_1507,N_1308);
nand U2208 (N_2208,N_1408,N_1308);
or U2209 (N_2209,N_1339,N_1448);
nand U2210 (N_2210,N_1527,N_1641);
nor U2211 (N_2211,N_1368,N_1529);
nor U2212 (N_2212,N_1393,N_1412);
nand U2213 (N_2213,N_1444,N_1717);
xnor U2214 (N_2214,N_1624,N_1574);
nand U2215 (N_2215,N_1786,N_1554);
xor U2216 (N_2216,N_1686,N_1609);
nor U2217 (N_2217,N_1343,N_1671);
nor U2218 (N_2218,N_1508,N_1784);
or U2219 (N_2219,N_1462,N_1405);
or U2220 (N_2220,N_1203,N_1789);
nand U2221 (N_2221,N_1563,N_1338);
and U2222 (N_2222,N_1642,N_1404);
nor U2223 (N_2223,N_1300,N_1262);
nor U2224 (N_2224,N_1572,N_1579);
nor U2225 (N_2225,N_1379,N_1746);
or U2226 (N_2226,N_1618,N_1736);
or U2227 (N_2227,N_1437,N_1425);
and U2228 (N_2228,N_1336,N_1284);
and U2229 (N_2229,N_1263,N_1468);
xor U2230 (N_2230,N_1720,N_1408);
or U2231 (N_2231,N_1518,N_1426);
or U2232 (N_2232,N_1490,N_1746);
nor U2233 (N_2233,N_1448,N_1530);
nand U2234 (N_2234,N_1493,N_1423);
nor U2235 (N_2235,N_1506,N_1286);
nand U2236 (N_2236,N_1607,N_1280);
and U2237 (N_2237,N_1297,N_1301);
xnor U2238 (N_2238,N_1744,N_1244);
and U2239 (N_2239,N_1481,N_1334);
or U2240 (N_2240,N_1326,N_1587);
nand U2241 (N_2241,N_1365,N_1506);
nand U2242 (N_2242,N_1661,N_1591);
or U2243 (N_2243,N_1281,N_1346);
or U2244 (N_2244,N_1285,N_1566);
nand U2245 (N_2245,N_1612,N_1657);
or U2246 (N_2246,N_1784,N_1449);
and U2247 (N_2247,N_1743,N_1740);
and U2248 (N_2248,N_1222,N_1420);
nand U2249 (N_2249,N_1724,N_1694);
and U2250 (N_2250,N_1366,N_1792);
xnor U2251 (N_2251,N_1657,N_1383);
or U2252 (N_2252,N_1645,N_1532);
nand U2253 (N_2253,N_1300,N_1590);
or U2254 (N_2254,N_1453,N_1511);
nor U2255 (N_2255,N_1406,N_1582);
and U2256 (N_2256,N_1779,N_1259);
nand U2257 (N_2257,N_1402,N_1257);
nor U2258 (N_2258,N_1610,N_1719);
nand U2259 (N_2259,N_1207,N_1712);
nor U2260 (N_2260,N_1530,N_1244);
xor U2261 (N_2261,N_1606,N_1637);
nand U2262 (N_2262,N_1339,N_1536);
and U2263 (N_2263,N_1347,N_1752);
nand U2264 (N_2264,N_1781,N_1300);
and U2265 (N_2265,N_1513,N_1731);
and U2266 (N_2266,N_1511,N_1704);
xor U2267 (N_2267,N_1205,N_1604);
nor U2268 (N_2268,N_1317,N_1769);
and U2269 (N_2269,N_1626,N_1243);
or U2270 (N_2270,N_1350,N_1445);
and U2271 (N_2271,N_1762,N_1480);
nor U2272 (N_2272,N_1646,N_1636);
or U2273 (N_2273,N_1378,N_1369);
or U2274 (N_2274,N_1257,N_1631);
nor U2275 (N_2275,N_1513,N_1485);
or U2276 (N_2276,N_1486,N_1763);
nand U2277 (N_2277,N_1750,N_1220);
and U2278 (N_2278,N_1331,N_1772);
nor U2279 (N_2279,N_1246,N_1565);
or U2280 (N_2280,N_1664,N_1549);
and U2281 (N_2281,N_1758,N_1725);
nand U2282 (N_2282,N_1219,N_1776);
nor U2283 (N_2283,N_1450,N_1577);
xnor U2284 (N_2284,N_1741,N_1454);
and U2285 (N_2285,N_1290,N_1743);
or U2286 (N_2286,N_1747,N_1568);
or U2287 (N_2287,N_1653,N_1589);
nor U2288 (N_2288,N_1528,N_1504);
or U2289 (N_2289,N_1511,N_1670);
nand U2290 (N_2290,N_1611,N_1208);
or U2291 (N_2291,N_1617,N_1527);
xor U2292 (N_2292,N_1719,N_1641);
and U2293 (N_2293,N_1596,N_1497);
or U2294 (N_2294,N_1780,N_1549);
or U2295 (N_2295,N_1390,N_1772);
nand U2296 (N_2296,N_1349,N_1663);
or U2297 (N_2297,N_1316,N_1439);
and U2298 (N_2298,N_1467,N_1719);
nor U2299 (N_2299,N_1673,N_1692);
or U2300 (N_2300,N_1383,N_1405);
or U2301 (N_2301,N_1259,N_1261);
nor U2302 (N_2302,N_1313,N_1363);
nand U2303 (N_2303,N_1261,N_1751);
and U2304 (N_2304,N_1353,N_1485);
or U2305 (N_2305,N_1590,N_1524);
nand U2306 (N_2306,N_1408,N_1476);
nor U2307 (N_2307,N_1480,N_1273);
nand U2308 (N_2308,N_1206,N_1243);
and U2309 (N_2309,N_1272,N_1688);
nand U2310 (N_2310,N_1434,N_1469);
and U2311 (N_2311,N_1575,N_1457);
or U2312 (N_2312,N_1420,N_1727);
and U2313 (N_2313,N_1706,N_1339);
xnor U2314 (N_2314,N_1456,N_1688);
nand U2315 (N_2315,N_1757,N_1254);
nor U2316 (N_2316,N_1548,N_1219);
and U2317 (N_2317,N_1542,N_1324);
or U2318 (N_2318,N_1509,N_1266);
nand U2319 (N_2319,N_1615,N_1211);
or U2320 (N_2320,N_1545,N_1456);
and U2321 (N_2321,N_1452,N_1513);
xor U2322 (N_2322,N_1654,N_1522);
and U2323 (N_2323,N_1665,N_1447);
xnor U2324 (N_2324,N_1602,N_1523);
xnor U2325 (N_2325,N_1698,N_1251);
xnor U2326 (N_2326,N_1298,N_1211);
and U2327 (N_2327,N_1373,N_1214);
nand U2328 (N_2328,N_1569,N_1323);
nor U2329 (N_2329,N_1202,N_1319);
nor U2330 (N_2330,N_1211,N_1790);
nor U2331 (N_2331,N_1710,N_1607);
nand U2332 (N_2332,N_1226,N_1385);
xor U2333 (N_2333,N_1461,N_1598);
nand U2334 (N_2334,N_1252,N_1353);
or U2335 (N_2335,N_1251,N_1248);
xnor U2336 (N_2336,N_1776,N_1634);
and U2337 (N_2337,N_1468,N_1395);
nand U2338 (N_2338,N_1703,N_1597);
and U2339 (N_2339,N_1239,N_1362);
nand U2340 (N_2340,N_1675,N_1613);
nand U2341 (N_2341,N_1323,N_1515);
or U2342 (N_2342,N_1587,N_1311);
or U2343 (N_2343,N_1566,N_1539);
nand U2344 (N_2344,N_1696,N_1625);
nor U2345 (N_2345,N_1539,N_1280);
nor U2346 (N_2346,N_1632,N_1554);
and U2347 (N_2347,N_1345,N_1703);
or U2348 (N_2348,N_1255,N_1485);
or U2349 (N_2349,N_1473,N_1450);
xor U2350 (N_2350,N_1233,N_1449);
or U2351 (N_2351,N_1404,N_1238);
nor U2352 (N_2352,N_1605,N_1628);
nand U2353 (N_2353,N_1217,N_1473);
and U2354 (N_2354,N_1535,N_1416);
nor U2355 (N_2355,N_1231,N_1521);
nor U2356 (N_2356,N_1636,N_1622);
and U2357 (N_2357,N_1527,N_1242);
and U2358 (N_2358,N_1514,N_1277);
xor U2359 (N_2359,N_1617,N_1649);
nor U2360 (N_2360,N_1321,N_1634);
or U2361 (N_2361,N_1721,N_1436);
nand U2362 (N_2362,N_1771,N_1757);
nor U2363 (N_2363,N_1772,N_1761);
nand U2364 (N_2364,N_1230,N_1531);
nand U2365 (N_2365,N_1740,N_1367);
nand U2366 (N_2366,N_1332,N_1740);
nor U2367 (N_2367,N_1353,N_1202);
xnor U2368 (N_2368,N_1363,N_1606);
nor U2369 (N_2369,N_1447,N_1379);
or U2370 (N_2370,N_1763,N_1530);
nand U2371 (N_2371,N_1523,N_1775);
nand U2372 (N_2372,N_1429,N_1755);
xnor U2373 (N_2373,N_1745,N_1521);
or U2374 (N_2374,N_1711,N_1420);
or U2375 (N_2375,N_1359,N_1735);
nand U2376 (N_2376,N_1296,N_1206);
xor U2377 (N_2377,N_1582,N_1326);
nor U2378 (N_2378,N_1791,N_1523);
nand U2379 (N_2379,N_1387,N_1673);
and U2380 (N_2380,N_1586,N_1528);
nor U2381 (N_2381,N_1579,N_1651);
nor U2382 (N_2382,N_1664,N_1654);
xor U2383 (N_2383,N_1565,N_1301);
nor U2384 (N_2384,N_1781,N_1623);
nor U2385 (N_2385,N_1577,N_1423);
xnor U2386 (N_2386,N_1455,N_1275);
nor U2387 (N_2387,N_1570,N_1647);
nor U2388 (N_2388,N_1756,N_1523);
or U2389 (N_2389,N_1206,N_1701);
nor U2390 (N_2390,N_1755,N_1703);
nor U2391 (N_2391,N_1641,N_1419);
or U2392 (N_2392,N_1522,N_1715);
nor U2393 (N_2393,N_1480,N_1508);
nor U2394 (N_2394,N_1444,N_1623);
or U2395 (N_2395,N_1338,N_1434);
xor U2396 (N_2396,N_1256,N_1311);
or U2397 (N_2397,N_1764,N_1631);
xor U2398 (N_2398,N_1416,N_1489);
or U2399 (N_2399,N_1429,N_1641);
nand U2400 (N_2400,N_2208,N_2267);
and U2401 (N_2401,N_1958,N_1994);
and U2402 (N_2402,N_1921,N_2109);
or U2403 (N_2403,N_1952,N_1863);
nor U2404 (N_2404,N_2232,N_2356);
nand U2405 (N_2405,N_2257,N_2057);
nor U2406 (N_2406,N_2096,N_1846);
or U2407 (N_2407,N_2065,N_2207);
nor U2408 (N_2408,N_1947,N_2119);
nand U2409 (N_2409,N_2392,N_1929);
and U2410 (N_2410,N_2358,N_1883);
and U2411 (N_2411,N_1961,N_2372);
nor U2412 (N_2412,N_1881,N_1829);
nor U2413 (N_2413,N_2366,N_2038);
or U2414 (N_2414,N_2317,N_2310);
and U2415 (N_2415,N_2399,N_2188);
or U2416 (N_2416,N_1977,N_2325);
xor U2417 (N_2417,N_2221,N_1923);
or U2418 (N_2418,N_2082,N_2297);
nor U2419 (N_2419,N_2084,N_2365);
nand U2420 (N_2420,N_1871,N_2278);
and U2421 (N_2421,N_2004,N_2281);
nor U2422 (N_2422,N_1817,N_2003);
nor U2423 (N_2423,N_2239,N_1950);
nand U2424 (N_2424,N_2313,N_2088);
nor U2425 (N_2425,N_1990,N_1896);
or U2426 (N_2426,N_1976,N_1967);
or U2427 (N_2427,N_1922,N_1866);
nand U2428 (N_2428,N_1802,N_2253);
nand U2429 (N_2429,N_2203,N_2319);
or U2430 (N_2430,N_2078,N_1848);
and U2431 (N_2431,N_2008,N_2064);
nor U2432 (N_2432,N_2315,N_1930);
nor U2433 (N_2433,N_2213,N_2070);
and U2434 (N_2434,N_2052,N_2206);
and U2435 (N_2435,N_1832,N_1833);
nor U2436 (N_2436,N_1862,N_1910);
nand U2437 (N_2437,N_2099,N_2229);
nor U2438 (N_2438,N_1854,N_2047);
xor U2439 (N_2439,N_2370,N_2246);
or U2440 (N_2440,N_2385,N_2039);
nand U2441 (N_2441,N_2153,N_2123);
or U2442 (N_2442,N_2383,N_2046);
nor U2443 (N_2443,N_2196,N_1877);
and U2444 (N_2444,N_2294,N_2201);
or U2445 (N_2445,N_2049,N_2388);
nor U2446 (N_2446,N_1805,N_2058);
nand U2447 (N_2447,N_2160,N_2181);
nand U2448 (N_2448,N_1864,N_2115);
nor U2449 (N_2449,N_2241,N_1996);
xor U2450 (N_2450,N_1853,N_1814);
and U2451 (N_2451,N_2093,N_2311);
xnor U2452 (N_2452,N_1999,N_1925);
or U2453 (N_2453,N_2216,N_2338);
nand U2454 (N_2454,N_2176,N_1978);
or U2455 (N_2455,N_1908,N_2265);
nor U2456 (N_2456,N_2116,N_2304);
nor U2457 (N_2457,N_1918,N_2056);
nor U2458 (N_2458,N_1931,N_2044);
nor U2459 (N_2459,N_2217,N_2318);
and U2460 (N_2460,N_1836,N_2354);
or U2461 (N_2461,N_2022,N_2118);
nor U2462 (N_2462,N_2136,N_2306);
nand U2463 (N_2463,N_2105,N_2301);
nand U2464 (N_2464,N_1948,N_2290);
nand U2465 (N_2465,N_1876,N_2337);
and U2466 (N_2466,N_1828,N_1882);
nand U2467 (N_2467,N_2296,N_1825);
nand U2468 (N_2468,N_1894,N_2156);
xor U2469 (N_2469,N_2390,N_2261);
or U2470 (N_2470,N_2215,N_2353);
xnor U2471 (N_2471,N_2134,N_1818);
and U2472 (N_2472,N_1974,N_1808);
or U2473 (N_2473,N_2340,N_1955);
nor U2474 (N_2474,N_1801,N_1949);
and U2475 (N_2475,N_2132,N_1819);
and U2476 (N_2476,N_1806,N_2226);
and U2477 (N_2477,N_2050,N_2351);
nand U2478 (N_2478,N_2314,N_2187);
or U2479 (N_2479,N_2143,N_2369);
nand U2480 (N_2480,N_2194,N_2270);
nor U2481 (N_2481,N_2086,N_1951);
xnor U2482 (N_2482,N_2076,N_1823);
nor U2483 (N_2483,N_2083,N_2193);
or U2484 (N_2484,N_1979,N_2066);
nor U2485 (N_2485,N_2240,N_1970);
xnor U2486 (N_2486,N_2191,N_2259);
and U2487 (N_2487,N_1956,N_2129);
nand U2488 (N_2488,N_1913,N_1867);
and U2489 (N_2489,N_2299,N_2378);
nor U2490 (N_2490,N_1892,N_2379);
or U2491 (N_2491,N_2072,N_2043);
nor U2492 (N_2492,N_2167,N_2382);
and U2493 (N_2493,N_2189,N_1984);
or U2494 (N_2494,N_2137,N_1803);
and U2495 (N_2495,N_1957,N_2026);
and U2496 (N_2496,N_2042,N_1932);
nor U2497 (N_2497,N_2100,N_2202);
nor U2498 (N_2498,N_2352,N_2092);
nand U2499 (N_2499,N_1900,N_2179);
nor U2500 (N_2500,N_2291,N_2178);
or U2501 (N_2501,N_2140,N_2211);
or U2502 (N_2502,N_2359,N_2108);
nor U2503 (N_2503,N_2157,N_2371);
and U2504 (N_2504,N_1945,N_1826);
and U2505 (N_2505,N_2081,N_2238);
nand U2506 (N_2506,N_2341,N_2329);
xor U2507 (N_2507,N_2235,N_1991);
nand U2508 (N_2508,N_1875,N_2219);
nand U2509 (N_2509,N_2210,N_1972);
xnor U2510 (N_2510,N_2288,N_2102);
or U2511 (N_2511,N_2074,N_2012);
nand U2512 (N_2512,N_1965,N_1981);
nor U2513 (N_2513,N_1917,N_1909);
xnor U2514 (N_2514,N_1860,N_2316);
nand U2515 (N_2515,N_2139,N_2249);
and U2516 (N_2516,N_2251,N_2032);
nor U2517 (N_2517,N_2357,N_1964);
nor U2518 (N_2518,N_2300,N_2247);
and U2519 (N_2519,N_1834,N_2060);
and U2520 (N_2520,N_2274,N_2151);
and U2521 (N_2521,N_2040,N_2225);
and U2522 (N_2522,N_2391,N_1988);
nand U2523 (N_2523,N_1904,N_2230);
or U2524 (N_2524,N_1901,N_1983);
nand U2525 (N_2525,N_1946,N_2333);
nor U2526 (N_2526,N_2200,N_2104);
or U2527 (N_2527,N_2381,N_2085);
xor U2528 (N_2528,N_2033,N_1940);
nor U2529 (N_2529,N_2166,N_1907);
nand U2530 (N_2530,N_1928,N_2069);
nor U2531 (N_2531,N_1812,N_1880);
and U2532 (N_2532,N_2283,N_2293);
nand U2533 (N_2533,N_2346,N_2113);
or U2534 (N_2534,N_2162,N_2159);
and U2535 (N_2535,N_2110,N_1912);
and U2536 (N_2536,N_2131,N_1858);
and U2537 (N_2537,N_1810,N_1998);
nand U2538 (N_2538,N_2007,N_2377);
and U2539 (N_2539,N_2095,N_2106);
nor U2540 (N_2540,N_1851,N_2209);
nand U2541 (N_2541,N_2360,N_2334);
nand U2542 (N_2542,N_2295,N_1869);
and U2543 (N_2543,N_2037,N_1980);
and U2544 (N_2544,N_1903,N_2326);
nor U2545 (N_2545,N_2255,N_2017);
xor U2546 (N_2546,N_1992,N_1830);
xor U2547 (N_2547,N_2324,N_2011);
or U2548 (N_2548,N_2089,N_1879);
nand U2549 (N_2549,N_2397,N_1822);
nand U2550 (N_2550,N_2393,N_2344);
nor U2551 (N_2551,N_1852,N_2073);
or U2552 (N_2552,N_2158,N_2126);
nor U2553 (N_2553,N_2248,N_2124);
and U2554 (N_2554,N_2266,N_2330);
xor U2555 (N_2555,N_1884,N_2094);
nor U2556 (N_2556,N_2015,N_2000);
and U2557 (N_2557,N_2091,N_2282);
or U2558 (N_2558,N_2260,N_2080);
and U2559 (N_2559,N_1926,N_1888);
nor U2560 (N_2560,N_2172,N_1827);
and U2561 (N_2561,N_1898,N_2234);
and U2562 (N_2562,N_2171,N_2336);
xnor U2563 (N_2563,N_2250,N_2263);
nor U2564 (N_2564,N_2205,N_2138);
nor U2565 (N_2565,N_2079,N_1989);
nor U2566 (N_2566,N_2059,N_2224);
or U2567 (N_2567,N_2002,N_2186);
nand U2568 (N_2568,N_2307,N_2231);
or U2569 (N_2569,N_1886,N_2036);
or U2570 (N_2570,N_2024,N_2025);
nand U2571 (N_2571,N_2114,N_1963);
or U2572 (N_2572,N_2305,N_1843);
nor U2573 (N_2573,N_1933,N_2192);
or U2574 (N_2574,N_2244,N_2214);
nor U2575 (N_2575,N_2063,N_2068);
nand U2576 (N_2576,N_1995,N_2242);
or U2577 (N_2577,N_1850,N_2130);
and U2578 (N_2578,N_1915,N_2394);
and U2579 (N_2579,N_2271,N_1820);
or U2580 (N_2580,N_2133,N_2165);
nor U2581 (N_2581,N_2031,N_2212);
nand U2582 (N_2582,N_1811,N_2269);
nand U2583 (N_2583,N_1845,N_2355);
xor U2584 (N_2584,N_2389,N_2125);
nand U2585 (N_2585,N_1835,N_1902);
nand U2586 (N_2586,N_2041,N_2141);
nor U2587 (N_2587,N_2312,N_2264);
nor U2588 (N_2588,N_1944,N_2335);
nand U2589 (N_2589,N_2331,N_2164);
and U2590 (N_2590,N_2256,N_2273);
and U2591 (N_2591,N_2175,N_1893);
nand U2592 (N_2592,N_1856,N_2289);
nand U2593 (N_2593,N_2021,N_1861);
nor U2594 (N_2594,N_2034,N_1914);
or U2595 (N_2595,N_1844,N_1924);
and U2596 (N_2596,N_1954,N_2062);
nor U2597 (N_2597,N_1973,N_1889);
or U2598 (N_2598,N_2161,N_1800);
nand U2599 (N_2599,N_2275,N_1953);
or U2600 (N_2600,N_2009,N_2035);
nor U2601 (N_2601,N_1920,N_2112);
nor U2602 (N_2602,N_2395,N_1857);
nor U2603 (N_2603,N_2376,N_2322);
nor U2604 (N_2604,N_2183,N_2195);
and U2605 (N_2605,N_2343,N_2236);
nand U2606 (N_2606,N_1872,N_1966);
nand U2607 (N_2607,N_2280,N_2148);
nor U2608 (N_2608,N_2097,N_2198);
or U2609 (N_2609,N_2152,N_2107);
nor U2610 (N_2610,N_2154,N_2010);
xnor U2611 (N_2611,N_2218,N_1878);
or U2612 (N_2612,N_1987,N_1935);
nor U2613 (N_2613,N_2228,N_2276);
and U2614 (N_2614,N_1985,N_2308);
nand U2615 (N_2615,N_2128,N_1824);
or U2616 (N_2616,N_2233,N_2163);
nor U2617 (N_2617,N_2197,N_2170);
and U2618 (N_2618,N_1982,N_2071);
nor U2619 (N_2619,N_2380,N_2286);
nor U2620 (N_2620,N_1865,N_1868);
nand U2621 (N_2621,N_2190,N_2364);
nor U2622 (N_2622,N_2292,N_2090);
nand U2623 (N_2623,N_1859,N_2268);
xor U2624 (N_2624,N_2347,N_2384);
nor U2625 (N_2625,N_2386,N_1942);
and U2626 (N_2626,N_1840,N_2019);
nand U2627 (N_2627,N_1962,N_2048);
or U2628 (N_2628,N_2030,N_1897);
or U2629 (N_2629,N_2054,N_2150);
and U2630 (N_2630,N_2342,N_2272);
and U2631 (N_2631,N_1887,N_1821);
nand U2632 (N_2632,N_1939,N_1938);
or U2633 (N_2633,N_1895,N_2028);
nand U2634 (N_2634,N_2145,N_2285);
and U2635 (N_2635,N_2362,N_1831);
nor U2636 (N_2636,N_2168,N_2016);
and U2637 (N_2637,N_1816,N_1911);
xnor U2638 (N_2638,N_2245,N_2349);
or U2639 (N_2639,N_1993,N_2323);
and U2640 (N_2640,N_2174,N_2006);
nand U2641 (N_2641,N_1943,N_2029);
nand U2642 (N_2642,N_2243,N_1937);
and U2643 (N_2643,N_2117,N_2339);
xor U2644 (N_2644,N_1804,N_2279);
xor U2645 (N_2645,N_2098,N_2184);
xor U2646 (N_2646,N_2001,N_1986);
nor U2647 (N_2647,N_2121,N_2014);
and U2648 (N_2648,N_2177,N_2332);
xnor U2649 (N_2649,N_2027,N_1837);
xor U2650 (N_2650,N_2142,N_2005);
and U2651 (N_2651,N_2222,N_2368);
nand U2652 (N_2652,N_1927,N_2396);
and U2653 (N_2653,N_1815,N_2302);
nand U2654 (N_2654,N_1891,N_1919);
or U2655 (N_2655,N_1969,N_2363);
nor U2656 (N_2656,N_2051,N_1874);
nand U2657 (N_2657,N_2398,N_2127);
nor U2658 (N_2658,N_2147,N_1809);
and U2659 (N_2659,N_2254,N_1870);
or U2660 (N_2660,N_2327,N_2237);
and U2661 (N_2661,N_2287,N_2077);
or U2662 (N_2662,N_2111,N_2173);
and U2663 (N_2663,N_1813,N_1842);
nand U2664 (N_2664,N_2373,N_2220);
nor U2665 (N_2665,N_2013,N_2185);
nor U2666 (N_2666,N_1906,N_2067);
nor U2667 (N_2667,N_2144,N_1847);
or U2668 (N_2668,N_2227,N_2321);
nand U2669 (N_2669,N_2061,N_2345);
or U2670 (N_2670,N_2284,N_1934);
nand U2671 (N_2671,N_2180,N_1849);
and U2672 (N_2672,N_1971,N_1916);
and U2673 (N_2673,N_2277,N_2149);
nand U2674 (N_2674,N_2387,N_1905);
nand U2675 (N_2675,N_2298,N_1890);
nor U2676 (N_2676,N_2374,N_2020);
or U2677 (N_2677,N_1997,N_2350);
or U2678 (N_2678,N_1838,N_2303);
and U2679 (N_2679,N_2262,N_2252);
nor U2680 (N_2680,N_1841,N_2146);
nand U2681 (N_2681,N_1941,N_2120);
nor U2682 (N_2682,N_2258,N_1873);
nor U2683 (N_2683,N_1839,N_2101);
xnor U2684 (N_2684,N_2223,N_1968);
nor U2685 (N_2685,N_2348,N_2155);
or U2686 (N_2686,N_2023,N_2182);
nand U2687 (N_2687,N_1936,N_2087);
or U2688 (N_2688,N_2103,N_2309);
or U2689 (N_2689,N_2135,N_2367);
or U2690 (N_2690,N_2122,N_2204);
nand U2691 (N_2691,N_2199,N_2075);
nand U2692 (N_2692,N_2328,N_1959);
and U2693 (N_2693,N_1899,N_1807);
and U2694 (N_2694,N_2320,N_2361);
nor U2695 (N_2695,N_1960,N_2053);
and U2696 (N_2696,N_2018,N_1855);
nand U2697 (N_2697,N_1975,N_2169);
or U2698 (N_2698,N_2375,N_2045);
nand U2699 (N_2699,N_2055,N_1885);
nand U2700 (N_2700,N_1940,N_2078);
nor U2701 (N_2701,N_1823,N_1952);
or U2702 (N_2702,N_1930,N_1923);
and U2703 (N_2703,N_2279,N_1864);
and U2704 (N_2704,N_1805,N_1924);
and U2705 (N_2705,N_1982,N_1900);
or U2706 (N_2706,N_2157,N_2369);
or U2707 (N_2707,N_1920,N_1978);
or U2708 (N_2708,N_2266,N_2392);
and U2709 (N_2709,N_2152,N_2287);
nand U2710 (N_2710,N_2272,N_1819);
xnor U2711 (N_2711,N_1810,N_2029);
or U2712 (N_2712,N_2027,N_2339);
or U2713 (N_2713,N_2095,N_1816);
nand U2714 (N_2714,N_2046,N_2325);
and U2715 (N_2715,N_2296,N_2362);
or U2716 (N_2716,N_2103,N_2294);
nor U2717 (N_2717,N_2055,N_1873);
and U2718 (N_2718,N_2035,N_2228);
nor U2719 (N_2719,N_1959,N_2096);
nor U2720 (N_2720,N_2211,N_2283);
xor U2721 (N_2721,N_1994,N_1940);
or U2722 (N_2722,N_1917,N_2307);
or U2723 (N_2723,N_2122,N_2079);
nor U2724 (N_2724,N_2396,N_2308);
and U2725 (N_2725,N_1813,N_1935);
nand U2726 (N_2726,N_2291,N_2046);
nand U2727 (N_2727,N_1855,N_2305);
nor U2728 (N_2728,N_1876,N_1970);
nor U2729 (N_2729,N_2369,N_2041);
nor U2730 (N_2730,N_2331,N_2126);
or U2731 (N_2731,N_2083,N_2219);
and U2732 (N_2732,N_1977,N_1864);
and U2733 (N_2733,N_2074,N_1869);
nand U2734 (N_2734,N_1935,N_2221);
nand U2735 (N_2735,N_2320,N_2113);
and U2736 (N_2736,N_2309,N_2106);
nor U2737 (N_2737,N_2016,N_2004);
nand U2738 (N_2738,N_2130,N_2375);
and U2739 (N_2739,N_1930,N_2242);
and U2740 (N_2740,N_1821,N_1944);
and U2741 (N_2741,N_2318,N_2345);
nor U2742 (N_2742,N_2151,N_1913);
nor U2743 (N_2743,N_1836,N_2217);
nor U2744 (N_2744,N_1870,N_2156);
or U2745 (N_2745,N_2096,N_2340);
nand U2746 (N_2746,N_2306,N_2008);
and U2747 (N_2747,N_2106,N_2352);
and U2748 (N_2748,N_2166,N_1846);
nand U2749 (N_2749,N_1934,N_2099);
and U2750 (N_2750,N_1947,N_2320);
or U2751 (N_2751,N_1926,N_2250);
and U2752 (N_2752,N_1932,N_2266);
xor U2753 (N_2753,N_2317,N_2019);
nor U2754 (N_2754,N_2101,N_2086);
nand U2755 (N_2755,N_2249,N_2126);
and U2756 (N_2756,N_2260,N_2241);
and U2757 (N_2757,N_1949,N_1902);
and U2758 (N_2758,N_2316,N_1825);
nor U2759 (N_2759,N_2057,N_2060);
nand U2760 (N_2760,N_1932,N_2179);
nand U2761 (N_2761,N_2309,N_2149);
and U2762 (N_2762,N_2051,N_1822);
nor U2763 (N_2763,N_2354,N_1952);
or U2764 (N_2764,N_2130,N_2100);
and U2765 (N_2765,N_2151,N_1936);
nor U2766 (N_2766,N_2288,N_2313);
or U2767 (N_2767,N_1915,N_2164);
or U2768 (N_2768,N_2339,N_2215);
and U2769 (N_2769,N_2002,N_2233);
or U2770 (N_2770,N_1937,N_2129);
nand U2771 (N_2771,N_2058,N_2090);
and U2772 (N_2772,N_2099,N_2144);
nand U2773 (N_2773,N_2169,N_2040);
and U2774 (N_2774,N_1970,N_1817);
or U2775 (N_2775,N_2100,N_2372);
nand U2776 (N_2776,N_1818,N_1829);
nor U2777 (N_2777,N_1940,N_2165);
nand U2778 (N_2778,N_1931,N_2207);
nand U2779 (N_2779,N_1901,N_1981);
and U2780 (N_2780,N_1883,N_2159);
or U2781 (N_2781,N_2078,N_1929);
nor U2782 (N_2782,N_2130,N_2002);
xnor U2783 (N_2783,N_2336,N_2146);
or U2784 (N_2784,N_2272,N_2388);
nand U2785 (N_2785,N_2375,N_2106);
and U2786 (N_2786,N_1965,N_2305);
xnor U2787 (N_2787,N_2395,N_2155);
and U2788 (N_2788,N_1983,N_2329);
and U2789 (N_2789,N_1870,N_2387);
and U2790 (N_2790,N_2383,N_1984);
nand U2791 (N_2791,N_2271,N_2346);
nand U2792 (N_2792,N_2044,N_1817);
or U2793 (N_2793,N_2283,N_2009);
nand U2794 (N_2794,N_2249,N_1823);
xnor U2795 (N_2795,N_2349,N_1872);
xnor U2796 (N_2796,N_2379,N_2020);
or U2797 (N_2797,N_1989,N_1971);
nor U2798 (N_2798,N_2329,N_2334);
nand U2799 (N_2799,N_2198,N_1926);
or U2800 (N_2800,N_2333,N_1934);
nor U2801 (N_2801,N_2059,N_2294);
nand U2802 (N_2802,N_2257,N_2006);
nand U2803 (N_2803,N_2058,N_1999);
and U2804 (N_2804,N_2249,N_2290);
nand U2805 (N_2805,N_2085,N_2232);
and U2806 (N_2806,N_2127,N_2358);
nor U2807 (N_2807,N_1865,N_2123);
and U2808 (N_2808,N_2266,N_2059);
and U2809 (N_2809,N_2332,N_2235);
and U2810 (N_2810,N_1852,N_2246);
nor U2811 (N_2811,N_2091,N_1981);
nand U2812 (N_2812,N_2033,N_2107);
nand U2813 (N_2813,N_2250,N_1925);
nor U2814 (N_2814,N_2071,N_2384);
or U2815 (N_2815,N_2259,N_1871);
or U2816 (N_2816,N_2083,N_1890);
nor U2817 (N_2817,N_2142,N_2221);
or U2818 (N_2818,N_2093,N_2136);
nor U2819 (N_2819,N_2120,N_1888);
nand U2820 (N_2820,N_1950,N_1810);
and U2821 (N_2821,N_2147,N_2324);
nand U2822 (N_2822,N_1862,N_2224);
and U2823 (N_2823,N_2216,N_2191);
and U2824 (N_2824,N_2361,N_1924);
nor U2825 (N_2825,N_2075,N_2329);
or U2826 (N_2826,N_2054,N_2229);
or U2827 (N_2827,N_1865,N_1938);
or U2828 (N_2828,N_2159,N_2236);
or U2829 (N_2829,N_1914,N_2313);
and U2830 (N_2830,N_2154,N_1889);
nand U2831 (N_2831,N_1991,N_1910);
and U2832 (N_2832,N_2275,N_2150);
nor U2833 (N_2833,N_2161,N_1811);
nand U2834 (N_2834,N_2338,N_1906);
or U2835 (N_2835,N_1811,N_2104);
nand U2836 (N_2836,N_1964,N_2048);
nand U2837 (N_2837,N_2303,N_2121);
nand U2838 (N_2838,N_1887,N_2112);
and U2839 (N_2839,N_2339,N_2244);
nand U2840 (N_2840,N_2163,N_1800);
or U2841 (N_2841,N_2109,N_2387);
or U2842 (N_2842,N_2221,N_2246);
or U2843 (N_2843,N_2079,N_2073);
nand U2844 (N_2844,N_1837,N_2113);
or U2845 (N_2845,N_1849,N_1894);
nor U2846 (N_2846,N_1950,N_2306);
and U2847 (N_2847,N_1831,N_2323);
nand U2848 (N_2848,N_2053,N_2150);
and U2849 (N_2849,N_1944,N_2142);
or U2850 (N_2850,N_2134,N_2355);
and U2851 (N_2851,N_2263,N_2093);
and U2852 (N_2852,N_2340,N_2022);
xnor U2853 (N_2853,N_2309,N_1844);
nor U2854 (N_2854,N_2315,N_1904);
or U2855 (N_2855,N_1856,N_2171);
and U2856 (N_2856,N_2299,N_1925);
or U2857 (N_2857,N_1925,N_2369);
nor U2858 (N_2858,N_2037,N_1947);
nor U2859 (N_2859,N_1917,N_2297);
xnor U2860 (N_2860,N_2392,N_1999);
xnor U2861 (N_2861,N_2124,N_2294);
nand U2862 (N_2862,N_2304,N_1912);
or U2863 (N_2863,N_2319,N_2173);
nor U2864 (N_2864,N_2199,N_2277);
nand U2865 (N_2865,N_1800,N_1842);
nand U2866 (N_2866,N_1859,N_2039);
or U2867 (N_2867,N_2178,N_2363);
nor U2868 (N_2868,N_2237,N_2336);
nor U2869 (N_2869,N_2305,N_2131);
or U2870 (N_2870,N_2182,N_2088);
and U2871 (N_2871,N_2326,N_2345);
nor U2872 (N_2872,N_1858,N_1812);
nor U2873 (N_2873,N_1935,N_2092);
nand U2874 (N_2874,N_2305,N_1972);
and U2875 (N_2875,N_2008,N_2028);
xor U2876 (N_2876,N_2212,N_1944);
xnor U2877 (N_2877,N_1852,N_1807);
and U2878 (N_2878,N_2116,N_2312);
and U2879 (N_2879,N_2354,N_1893);
and U2880 (N_2880,N_1919,N_2346);
nand U2881 (N_2881,N_1824,N_2189);
nor U2882 (N_2882,N_1804,N_2182);
or U2883 (N_2883,N_2361,N_2132);
and U2884 (N_2884,N_1865,N_1901);
nor U2885 (N_2885,N_2168,N_2124);
or U2886 (N_2886,N_1812,N_2015);
or U2887 (N_2887,N_1805,N_1997);
nand U2888 (N_2888,N_2152,N_2211);
nor U2889 (N_2889,N_1871,N_2351);
nor U2890 (N_2890,N_2374,N_2255);
and U2891 (N_2891,N_2348,N_2091);
and U2892 (N_2892,N_2345,N_2056);
and U2893 (N_2893,N_2334,N_1867);
or U2894 (N_2894,N_2379,N_1942);
or U2895 (N_2895,N_2031,N_2225);
nand U2896 (N_2896,N_2333,N_2086);
xnor U2897 (N_2897,N_2049,N_2250);
and U2898 (N_2898,N_2139,N_1924);
nor U2899 (N_2899,N_2000,N_2136);
or U2900 (N_2900,N_2152,N_2003);
and U2901 (N_2901,N_2081,N_1959);
nor U2902 (N_2902,N_2239,N_2282);
and U2903 (N_2903,N_2224,N_2175);
nand U2904 (N_2904,N_1876,N_2266);
nand U2905 (N_2905,N_1990,N_1886);
and U2906 (N_2906,N_2346,N_2265);
nand U2907 (N_2907,N_1953,N_2052);
or U2908 (N_2908,N_2086,N_2043);
or U2909 (N_2909,N_2117,N_2317);
nand U2910 (N_2910,N_1960,N_2140);
nor U2911 (N_2911,N_2229,N_2389);
or U2912 (N_2912,N_2366,N_2285);
or U2913 (N_2913,N_1962,N_2372);
or U2914 (N_2914,N_2359,N_1858);
nor U2915 (N_2915,N_2064,N_1924);
and U2916 (N_2916,N_2132,N_1878);
xnor U2917 (N_2917,N_1985,N_1917);
or U2918 (N_2918,N_2014,N_1887);
nor U2919 (N_2919,N_2225,N_1985);
xor U2920 (N_2920,N_1842,N_1957);
nand U2921 (N_2921,N_1914,N_1847);
nor U2922 (N_2922,N_2241,N_2096);
xor U2923 (N_2923,N_2211,N_1873);
nand U2924 (N_2924,N_2025,N_2075);
nor U2925 (N_2925,N_2175,N_1848);
and U2926 (N_2926,N_2179,N_2332);
or U2927 (N_2927,N_2049,N_2214);
or U2928 (N_2928,N_2109,N_2380);
or U2929 (N_2929,N_2279,N_2287);
xor U2930 (N_2930,N_2085,N_2114);
nand U2931 (N_2931,N_2231,N_2338);
nand U2932 (N_2932,N_1868,N_1812);
nor U2933 (N_2933,N_1971,N_2217);
nand U2934 (N_2934,N_1989,N_2341);
and U2935 (N_2935,N_2122,N_1898);
and U2936 (N_2936,N_1817,N_2178);
nor U2937 (N_2937,N_2261,N_1972);
nand U2938 (N_2938,N_1970,N_1961);
and U2939 (N_2939,N_2387,N_2220);
and U2940 (N_2940,N_2152,N_2244);
and U2941 (N_2941,N_2010,N_2218);
or U2942 (N_2942,N_1949,N_2187);
or U2943 (N_2943,N_1890,N_2099);
nand U2944 (N_2944,N_2162,N_2356);
nor U2945 (N_2945,N_2386,N_1839);
nand U2946 (N_2946,N_1964,N_1931);
and U2947 (N_2947,N_2382,N_2113);
or U2948 (N_2948,N_2071,N_2063);
and U2949 (N_2949,N_1852,N_2235);
nand U2950 (N_2950,N_1819,N_2178);
and U2951 (N_2951,N_2160,N_2162);
or U2952 (N_2952,N_1898,N_2185);
and U2953 (N_2953,N_1980,N_2278);
nor U2954 (N_2954,N_1879,N_2325);
and U2955 (N_2955,N_2115,N_2312);
nand U2956 (N_2956,N_1985,N_2038);
nand U2957 (N_2957,N_1925,N_2186);
and U2958 (N_2958,N_1814,N_2371);
nand U2959 (N_2959,N_2143,N_2137);
nand U2960 (N_2960,N_1889,N_1974);
nand U2961 (N_2961,N_2184,N_1805);
nand U2962 (N_2962,N_1939,N_2343);
nand U2963 (N_2963,N_2034,N_2242);
and U2964 (N_2964,N_1807,N_2192);
and U2965 (N_2965,N_2323,N_1843);
nor U2966 (N_2966,N_1942,N_2029);
nor U2967 (N_2967,N_2181,N_2092);
nand U2968 (N_2968,N_2373,N_2079);
xor U2969 (N_2969,N_1895,N_2283);
or U2970 (N_2970,N_2218,N_1950);
or U2971 (N_2971,N_1956,N_2331);
and U2972 (N_2972,N_2255,N_2152);
nand U2973 (N_2973,N_1965,N_1972);
and U2974 (N_2974,N_2133,N_2275);
nand U2975 (N_2975,N_2018,N_2383);
or U2976 (N_2976,N_2074,N_1817);
and U2977 (N_2977,N_1933,N_2249);
nor U2978 (N_2978,N_1975,N_2376);
xor U2979 (N_2979,N_2240,N_1826);
nand U2980 (N_2980,N_2011,N_2126);
or U2981 (N_2981,N_2243,N_2138);
nor U2982 (N_2982,N_2383,N_1951);
nand U2983 (N_2983,N_2324,N_2180);
or U2984 (N_2984,N_2072,N_2193);
and U2985 (N_2985,N_1903,N_2029);
nand U2986 (N_2986,N_2229,N_2381);
and U2987 (N_2987,N_2178,N_1995);
nand U2988 (N_2988,N_2200,N_1967);
and U2989 (N_2989,N_2032,N_2144);
or U2990 (N_2990,N_2010,N_1940);
and U2991 (N_2991,N_2200,N_2390);
and U2992 (N_2992,N_2362,N_2304);
or U2993 (N_2993,N_1943,N_1827);
nor U2994 (N_2994,N_2335,N_1836);
or U2995 (N_2995,N_2169,N_2259);
nand U2996 (N_2996,N_2042,N_1849);
xor U2997 (N_2997,N_2066,N_2263);
nor U2998 (N_2998,N_2060,N_2320);
nand U2999 (N_2999,N_1823,N_1824);
or UO_0 (O_0,N_2655,N_2413);
nand UO_1 (O_1,N_2934,N_2817);
and UO_2 (O_2,N_2879,N_2599);
and UO_3 (O_3,N_2444,N_2972);
and UO_4 (O_4,N_2797,N_2981);
or UO_5 (O_5,N_2710,N_2932);
nor UO_6 (O_6,N_2490,N_2585);
nand UO_7 (O_7,N_2827,N_2813);
nor UO_8 (O_8,N_2952,N_2892);
or UO_9 (O_9,N_2753,N_2534);
and UO_10 (O_10,N_2890,N_2909);
nand UO_11 (O_11,N_2808,N_2623);
nor UO_12 (O_12,N_2885,N_2537);
or UO_13 (O_13,N_2662,N_2888);
and UO_14 (O_14,N_2525,N_2842);
nor UO_15 (O_15,N_2877,N_2510);
and UO_16 (O_16,N_2939,N_2648);
nand UO_17 (O_17,N_2647,N_2938);
or UO_18 (O_18,N_2872,N_2796);
or UO_19 (O_19,N_2994,N_2806);
nor UO_20 (O_20,N_2705,N_2670);
xnor UO_21 (O_21,N_2787,N_2450);
and UO_22 (O_22,N_2673,N_2788);
nor UO_23 (O_23,N_2959,N_2677);
or UO_24 (O_24,N_2503,N_2911);
xnor UO_25 (O_25,N_2804,N_2401);
nor UO_26 (O_26,N_2702,N_2881);
nor UO_27 (O_27,N_2426,N_2604);
nor UO_28 (O_28,N_2828,N_2697);
xnor UO_29 (O_29,N_2699,N_2531);
and UO_30 (O_30,N_2491,N_2843);
and UO_31 (O_31,N_2567,N_2955);
nor UO_32 (O_32,N_2584,N_2935);
nand UO_33 (O_33,N_2402,N_2529);
and UO_34 (O_34,N_2887,N_2763);
or UO_35 (O_35,N_2985,N_2860);
nor UO_36 (O_36,N_2743,N_2722);
and UO_37 (O_37,N_2865,N_2666);
xnor UO_38 (O_38,N_2875,N_2632);
xor UO_39 (O_39,N_2993,N_2975);
nand UO_40 (O_40,N_2807,N_2476);
nand UO_41 (O_41,N_2597,N_2509);
or UO_42 (O_42,N_2578,N_2992);
nor UO_43 (O_43,N_2618,N_2580);
nor UO_44 (O_44,N_2498,N_2547);
nor UO_45 (O_45,N_2989,N_2668);
nor UO_46 (O_46,N_2999,N_2447);
nor UO_47 (O_47,N_2424,N_2969);
nand UO_48 (O_48,N_2440,N_2484);
nand UO_49 (O_49,N_2944,N_2453);
nor UO_50 (O_50,N_2431,N_2734);
or UO_51 (O_51,N_2683,N_2583);
nand UO_52 (O_52,N_2507,N_2778);
nor UO_53 (O_53,N_2433,N_2575);
nand UO_54 (O_54,N_2684,N_2949);
xor UO_55 (O_55,N_2940,N_2415);
and UO_56 (O_56,N_2965,N_2620);
nor UO_57 (O_57,N_2518,N_2732);
nor UO_58 (O_58,N_2884,N_2953);
nor UO_59 (O_59,N_2707,N_2590);
nor UO_60 (O_60,N_2750,N_2492);
nor UO_61 (O_61,N_2480,N_2400);
nand UO_62 (O_62,N_2915,N_2644);
nand UO_63 (O_63,N_2499,N_2463);
nor UO_64 (O_64,N_2616,N_2669);
and UO_65 (O_65,N_2641,N_2443);
nand UO_66 (O_66,N_2967,N_2728);
or UO_67 (O_67,N_2589,N_2675);
and UO_68 (O_68,N_2595,N_2445);
xnor UO_69 (O_69,N_2749,N_2452);
or UO_70 (O_70,N_2626,N_2792);
xnor UO_71 (O_71,N_2504,N_2555);
xor UO_72 (O_72,N_2614,N_2550);
and UO_73 (O_73,N_2466,N_2624);
or UO_74 (O_74,N_2682,N_2726);
or UO_75 (O_75,N_2645,N_2947);
nand UO_76 (O_76,N_2689,N_2736);
nand UO_77 (O_77,N_2837,N_2962);
nand UO_78 (O_78,N_2783,N_2556);
nand UO_79 (O_79,N_2448,N_2824);
nor UO_80 (O_80,N_2945,N_2630);
nand UO_81 (O_81,N_2990,N_2766);
and UO_82 (O_82,N_2869,N_2970);
nor UO_83 (O_83,N_2536,N_2759);
or UO_84 (O_84,N_2619,N_2846);
nor UO_85 (O_85,N_2698,N_2554);
nand UO_86 (O_86,N_2781,N_2951);
and UO_87 (O_87,N_2652,N_2470);
xnor UO_88 (O_88,N_2936,N_2421);
and UO_89 (O_89,N_2876,N_2716);
nand UO_90 (O_90,N_2977,N_2795);
and UO_91 (O_91,N_2637,N_2408);
nor UO_92 (O_92,N_2891,N_2995);
nor UO_93 (O_93,N_2956,N_2658);
or UO_94 (O_94,N_2775,N_2786);
and UO_95 (O_95,N_2568,N_2929);
and UO_96 (O_96,N_2600,N_2727);
or UO_97 (O_97,N_2908,N_2686);
nor UO_98 (O_98,N_2617,N_2570);
xor UO_99 (O_99,N_2767,N_2744);
xnor UO_100 (O_100,N_2719,N_2678);
xor UO_101 (O_101,N_2672,N_2449);
and UO_102 (O_102,N_2712,N_2609);
nor UO_103 (O_103,N_2986,N_2416);
xor UO_104 (O_104,N_2411,N_2920);
and UO_105 (O_105,N_2454,N_2690);
nor UO_106 (O_106,N_2560,N_2591);
xnor UO_107 (O_107,N_2695,N_2906);
and UO_108 (O_108,N_2841,N_2883);
and UO_109 (O_109,N_2954,N_2847);
nor UO_110 (O_110,N_2825,N_2897);
nand UO_111 (O_111,N_2487,N_2901);
and UO_112 (O_112,N_2810,N_2533);
and UO_113 (O_113,N_2918,N_2552);
nand UO_114 (O_114,N_2653,N_2541);
nand UO_115 (O_115,N_2500,N_2638);
and UO_116 (O_116,N_2755,N_2823);
nor UO_117 (O_117,N_2611,N_2714);
and UO_118 (O_118,N_2966,N_2866);
nor UO_119 (O_119,N_2905,N_2765);
and UO_120 (O_120,N_2709,N_2627);
nand UO_121 (O_121,N_2571,N_2545);
nand UO_122 (O_122,N_2809,N_2943);
nand UO_123 (O_123,N_2548,N_2687);
xor UO_124 (O_124,N_2640,N_2770);
and UO_125 (O_125,N_2403,N_2826);
or UO_126 (O_126,N_2631,N_2665);
nand UO_127 (O_127,N_2458,N_2838);
nand UO_128 (O_128,N_2873,N_2963);
or UO_129 (O_129,N_2691,N_2871);
or UO_130 (O_130,N_2671,N_2633);
nor UO_131 (O_131,N_2815,N_2836);
nor UO_132 (O_132,N_2622,N_2978);
or UO_133 (O_133,N_2798,N_2853);
nand UO_134 (O_134,N_2835,N_2907);
and UO_135 (O_135,N_2729,N_2696);
nand UO_136 (O_136,N_2814,N_2680);
or UO_137 (O_137,N_2464,N_2667);
nand UO_138 (O_138,N_2980,N_2864);
nand UO_139 (O_139,N_2852,N_2832);
or UO_140 (O_140,N_2708,N_2868);
and UO_141 (O_141,N_2418,N_2979);
nor UO_142 (O_142,N_2894,N_2780);
xor UO_143 (O_143,N_2818,N_2922);
nand UO_144 (O_144,N_2473,N_2654);
nor UO_145 (O_145,N_2478,N_2521);
xnor UO_146 (O_146,N_2557,N_2742);
xnor UO_147 (O_147,N_2844,N_2880);
nand UO_148 (O_148,N_2479,N_2776);
or UO_149 (O_149,N_2739,N_2629);
or UO_150 (O_150,N_2405,N_2855);
nor UO_151 (O_151,N_2800,N_2506);
and UO_152 (O_152,N_2738,N_2694);
nor UO_153 (O_153,N_2982,N_2700);
xor UO_154 (O_154,N_2659,N_2477);
nor UO_155 (O_155,N_2779,N_2974);
nand UO_156 (O_156,N_2586,N_2520);
or UO_157 (O_157,N_2820,N_2542);
nor UO_158 (O_158,N_2451,N_2486);
and UO_159 (O_159,N_2983,N_2931);
nor UO_160 (O_160,N_2467,N_2751);
and UO_161 (O_161,N_2756,N_2651);
and UO_162 (O_162,N_2957,N_2829);
or UO_163 (O_163,N_2893,N_2497);
and UO_164 (O_164,N_2927,N_2522);
and UO_165 (O_165,N_2886,N_2960);
nand UO_166 (O_166,N_2482,N_2515);
and UO_167 (O_167,N_2771,N_2845);
and UO_168 (O_168,N_2821,N_2532);
nor UO_169 (O_169,N_2693,N_2688);
nand UO_170 (O_170,N_2976,N_2946);
nor UO_171 (O_171,N_2928,N_2715);
nand UO_172 (O_172,N_2774,N_2530);
and UO_173 (O_173,N_2642,N_2914);
nand UO_174 (O_174,N_2471,N_2441);
and UO_175 (O_175,N_2551,N_2527);
nand UO_176 (O_176,N_2538,N_2754);
nor UO_177 (O_177,N_2519,N_2540);
and UO_178 (O_178,N_2725,N_2895);
and UO_179 (O_179,N_2535,N_2916);
and UO_180 (O_180,N_2636,N_2588);
nor UO_181 (O_181,N_2816,N_2839);
or UO_182 (O_182,N_2941,N_2747);
or UO_183 (O_183,N_2723,N_2517);
or UO_184 (O_184,N_2442,N_2997);
nor UO_185 (O_185,N_2410,N_2831);
or UO_186 (O_186,N_2475,N_2602);
nor UO_187 (O_187,N_2730,N_2679);
nand UO_188 (O_188,N_2516,N_2528);
nor UO_189 (O_189,N_2582,N_2576);
and UO_190 (O_190,N_2917,N_2446);
xnor UO_191 (O_191,N_2802,N_2713);
nor UO_192 (O_192,N_2437,N_2791);
or UO_193 (O_193,N_2737,N_2858);
nand UO_194 (O_194,N_2925,N_2439);
and UO_195 (O_195,N_2805,N_2769);
or UO_196 (O_196,N_2973,N_2812);
nand UO_197 (O_197,N_2903,N_2502);
xor UO_198 (O_198,N_2513,N_2924);
or UO_199 (O_199,N_2564,N_2902);
xor UO_200 (O_200,N_2933,N_2762);
xnor UO_201 (O_201,N_2711,N_2427);
nor UO_202 (O_202,N_2610,N_2561);
xor UO_203 (O_203,N_2745,N_2608);
or UO_204 (O_204,N_2988,N_2607);
nor UO_205 (O_205,N_2472,N_2462);
nor UO_206 (O_206,N_2596,N_2857);
and UO_207 (O_207,N_2434,N_2919);
nor UO_208 (O_208,N_2674,N_2758);
nand UO_209 (O_209,N_2848,N_2573);
nor UO_210 (O_210,N_2468,N_2459);
and UO_211 (O_211,N_2457,N_2628);
and UO_212 (O_212,N_2469,N_2495);
or UO_213 (O_213,N_2741,N_2834);
nor UO_214 (O_214,N_2731,N_2899);
or UO_215 (O_215,N_2593,N_2692);
and UO_216 (O_216,N_2921,N_2950);
or UO_217 (O_217,N_2910,N_2489);
nand UO_218 (O_218,N_2508,N_2579);
or UO_219 (O_219,N_2456,N_2904);
nor UO_220 (O_220,N_2874,N_2773);
nor UO_221 (O_221,N_2615,N_2870);
xor UO_222 (O_222,N_2748,N_2664);
or UO_223 (O_223,N_2819,N_2438);
or UO_224 (O_224,N_2889,N_2942);
nor UO_225 (O_225,N_2937,N_2811);
nand UO_226 (O_226,N_2423,N_2801);
xnor UO_227 (O_227,N_2681,N_2577);
and UO_228 (O_228,N_2514,N_2840);
nor UO_229 (O_229,N_2958,N_2996);
or UO_230 (O_230,N_2496,N_2803);
nor UO_231 (O_231,N_2526,N_2882);
or UO_232 (O_232,N_2948,N_2488);
xor UO_233 (O_233,N_2420,N_2740);
nand UO_234 (O_234,N_2833,N_2603);
or UO_235 (O_235,N_2856,N_2559);
nand UO_236 (O_236,N_2657,N_2850);
nor UO_237 (O_237,N_2634,N_2785);
nor UO_238 (O_238,N_2572,N_2404);
xor UO_239 (O_239,N_2406,N_2861);
xor UO_240 (O_240,N_2984,N_2761);
or UO_241 (O_241,N_2701,N_2768);
or UO_242 (O_242,N_2505,N_2587);
or UO_243 (O_243,N_2830,N_2598);
nand UO_244 (O_244,N_2563,N_2772);
and UO_245 (O_245,N_2493,N_2913);
or UO_246 (O_246,N_2646,N_2964);
nand UO_247 (O_247,N_2409,N_2436);
and UO_248 (O_248,N_2494,N_2417);
nand UO_249 (O_249,N_2660,N_2923);
nor UO_250 (O_250,N_2912,N_2419);
and UO_251 (O_251,N_2706,N_2724);
nand UO_252 (O_252,N_2435,N_2606);
and UO_253 (O_253,N_2961,N_2625);
nand UO_254 (O_254,N_2549,N_2601);
nand UO_255 (O_255,N_2661,N_2863);
or UO_256 (O_256,N_2483,N_2703);
xor UO_257 (O_257,N_2465,N_2562);
nor UO_258 (O_258,N_2422,N_2764);
and UO_259 (O_259,N_2735,N_2432);
nand UO_260 (O_260,N_2971,N_2720);
or UO_261 (O_261,N_2460,N_2639);
nor UO_262 (O_262,N_2574,N_2746);
and UO_263 (O_263,N_2635,N_2733);
xnor UO_264 (O_264,N_2782,N_2926);
or UO_265 (O_265,N_2429,N_2524);
or UO_266 (O_266,N_2991,N_2663);
nand UO_267 (O_267,N_2501,N_2414);
and UO_268 (O_268,N_2474,N_2704);
and UO_269 (O_269,N_2676,N_2539);
and UO_270 (O_270,N_2643,N_2412);
and UO_271 (O_271,N_2543,N_2425);
and UO_272 (O_272,N_2799,N_2544);
or UO_273 (O_273,N_2718,N_2523);
nand UO_274 (O_274,N_2789,N_2512);
nand UO_275 (O_275,N_2566,N_2553);
xnor UO_276 (O_276,N_2862,N_2565);
xor UO_277 (O_277,N_2594,N_2428);
and UO_278 (O_278,N_2898,N_2777);
nor UO_279 (O_279,N_2407,N_2650);
nor UO_280 (O_280,N_2752,N_2790);
nor UO_281 (O_281,N_2485,N_2649);
or UO_282 (O_282,N_2849,N_2896);
nor UO_283 (O_283,N_2859,N_2784);
nor UO_284 (O_284,N_2546,N_2930);
nand UO_285 (O_285,N_2760,N_2757);
and UO_286 (O_286,N_2878,N_2569);
or UO_287 (O_287,N_2621,N_2998);
nor UO_288 (O_288,N_2511,N_2822);
or UO_289 (O_289,N_2558,N_2612);
and UO_290 (O_290,N_2987,N_2794);
or UO_291 (O_291,N_2717,N_2605);
nor UO_292 (O_292,N_2685,N_2968);
nand UO_293 (O_293,N_2461,N_2430);
and UO_294 (O_294,N_2656,N_2581);
xnor UO_295 (O_295,N_2793,N_2854);
and UO_296 (O_296,N_2900,N_2851);
or UO_297 (O_297,N_2455,N_2721);
nand UO_298 (O_298,N_2592,N_2867);
nand UO_299 (O_299,N_2613,N_2481);
and UO_300 (O_300,N_2687,N_2714);
nand UO_301 (O_301,N_2976,N_2633);
nor UO_302 (O_302,N_2652,N_2765);
and UO_303 (O_303,N_2757,N_2580);
nand UO_304 (O_304,N_2878,N_2960);
nor UO_305 (O_305,N_2910,N_2770);
and UO_306 (O_306,N_2655,N_2962);
nor UO_307 (O_307,N_2951,N_2507);
xor UO_308 (O_308,N_2645,N_2784);
or UO_309 (O_309,N_2823,N_2978);
nand UO_310 (O_310,N_2961,N_2813);
nand UO_311 (O_311,N_2507,N_2936);
or UO_312 (O_312,N_2625,N_2745);
or UO_313 (O_313,N_2436,N_2772);
nand UO_314 (O_314,N_2844,N_2948);
and UO_315 (O_315,N_2945,N_2691);
and UO_316 (O_316,N_2849,N_2612);
and UO_317 (O_317,N_2777,N_2647);
and UO_318 (O_318,N_2953,N_2862);
nor UO_319 (O_319,N_2428,N_2514);
and UO_320 (O_320,N_2849,N_2557);
nand UO_321 (O_321,N_2503,N_2512);
or UO_322 (O_322,N_2490,N_2600);
and UO_323 (O_323,N_2791,N_2522);
nor UO_324 (O_324,N_2805,N_2502);
nand UO_325 (O_325,N_2631,N_2483);
or UO_326 (O_326,N_2521,N_2732);
and UO_327 (O_327,N_2716,N_2480);
and UO_328 (O_328,N_2407,N_2944);
and UO_329 (O_329,N_2454,N_2884);
nor UO_330 (O_330,N_2499,N_2557);
or UO_331 (O_331,N_2594,N_2648);
nor UO_332 (O_332,N_2475,N_2534);
and UO_333 (O_333,N_2805,N_2938);
nand UO_334 (O_334,N_2739,N_2423);
and UO_335 (O_335,N_2791,N_2448);
nand UO_336 (O_336,N_2827,N_2880);
nor UO_337 (O_337,N_2781,N_2593);
or UO_338 (O_338,N_2786,N_2952);
and UO_339 (O_339,N_2770,N_2442);
xnor UO_340 (O_340,N_2652,N_2625);
nand UO_341 (O_341,N_2652,N_2705);
nor UO_342 (O_342,N_2618,N_2594);
and UO_343 (O_343,N_2857,N_2433);
and UO_344 (O_344,N_2686,N_2549);
nor UO_345 (O_345,N_2903,N_2578);
nand UO_346 (O_346,N_2761,N_2974);
or UO_347 (O_347,N_2588,N_2507);
and UO_348 (O_348,N_2539,N_2470);
or UO_349 (O_349,N_2450,N_2675);
nand UO_350 (O_350,N_2692,N_2418);
xor UO_351 (O_351,N_2820,N_2595);
nand UO_352 (O_352,N_2620,N_2530);
or UO_353 (O_353,N_2766,N_2754);
nand UO_354 (O_354,N_2494,N_2925);
or UO_355 (O_355,N_2625,N_2799);
nor UO_356 (O_356,N_2547,N_2617);
nor UO_357 (O_357,N_2870,N_2774);
or UO_358 (O_358,N_2402,N_2755);
or UO_359 (O_359,N_2434,N_2934);
nor UO_360 (O_360,N_2949,N_2479);
or UO_361 (O_361,N_2851,N_2823);
nand UO_362 (O_362,N_2559,N_2446);
or UO_363 (O_363,N_2845,N_2854);
or UO_364 (O_364,N_2958,N_2831);
nand UO_365 (O_365,N_2508,N_2404);
nand UO_366 (O_366,N_2986,N_2617);
nor UO_367 (O_367,N_2521,N_2936);
and UO_368 (O_368,N_2993,N_2899);
nor UO_369 (O_369,N_2654,N_2680);
or UO_370 (O_370,N_2820,N_2503);
or UO_371 (O_371,N_2514,N_2554);
nor UO_372 (O_372,N_2739,N_2995);
xnor UO_373 (O_373,N_2826,N_2442);
or UO_374 (O_374,N_2819,N_2957);
and UO_375 (O_375,N_2435,N_2877);
nor UO_376 (O_376,N_2493,N_2697);
xor UO_377 (O_377,N_2777,N_2827);
nand UO_378 (O_378,N_2507,N_2639);
nand UO_379 (O_379,N_2813,N_2602);
nor UO_380 (O_380,N_2929,N_2981);
and UO_381 (O_381,N_2446,N_2512);
nor UO_382 (O_382,N_2679,N_2444);
nor UO_383 (O_383,N_2776,N_2767);
xnor UO_384 (O_384,N_2858,N_2713);
or UO_385 (O_385,N_2636,N_2700);
xor UO_386 (O_386,N_2779,N_2726);
nor UO_387 (O_387,N_2952,N_2534);
and UO_388 (O_388,N_2860,N_2564);
or UO_389 (O_389,N_2870,N_2737);
or UO_390 (O_390,N_2520,N_2557);
and UO_391 (O_391,N_2657,N_2724);
nor UO_392 (O_392,N_2629,N_2700);
nand UO_393 (O_393,N_2875,N_2816);
nand UO_394 (O_394,N_2815,N_2695);
nor UO_395 (O_395,N_2782,N_2876);
nor UO_396 (O_396,N_2627,N_2897);
nand UO_397 (O_397,N_2676,N_2798);
and UO_398 (O_398,N_2792,N_2655);
or UO_399 (O_399,N_2661,N_2953);
and UO_400 (O_400,N_2772,N_2699);
xnor UO_401 (O_401,N_2568,N_2665);
nor UO_402 (O_402,N_2489,N_2872);
xor UO_403 (O_403,N_2408,N_2548);
nor UO_404 (O_404,N_2925,N_2899);
xnor UO_405 (O_405,N_2824,N_2896);
or UO_406 (O_406,N_2558,N_2564);
nor UO_407 (O_407,N_2669,N_2629);
and UO_408 (O_408,N_2582,N_2493);
and UO_409 (O_409,N_2535,N_2732);
or UO_410 (O_410,N_2971,N_2741);
and UO_411 (O_411,N_2929,N_2514);
and UO_412 (O_412,N_2822,N_2482);
and UO_413 (O_413,N_2812,N_2991);
nor UO_414 (O_414,N_2562,N_2598);
nand UO_415 (O_415,N_2588,N_2799);
nor UO_416 (O_416,N_2958,N_2489);
nor UO_417 (O_417,N_2514,N_2906);
or UO_418 (O_418,N_2417,N_2836);
or UO_419 (O_419,N_2983,N_2445);
nand UO_420 (O_420,N_2719,N_2920);
nand UO_421 (O_421,N_2920,N_2549);
and UO_422 (O_422,N_2417,N_2676);
or UO_423 (O_423,N_2947,N_2711);
nand UO_424 (O_424,N_2789,N_2537);
xnor UO_425 (O_425,N_2836,N_2999);
and UO_426 (O_426,N_2725,N_2533);
nand UO_427 (O_427,N_2594,N_2584);
nand UO_428 (O_428,N_2665,N_2462);
and UO_429 (O_429,N_2699,N_2525);
or UO_430 (O_430,N_2650,N_2857);
nor UO_431 (O_431,N_2935,N_2905);
nand UO_432 (O_432,N_2783,N_2837);
or UO_433 (O_433,N_2586,N_2657);
and UO_434 (O_434,N_2620,N_2472);
nor UO_435 (O_435,N_2606,N_2480);
nand UO_436 (O_436,N_2905,N_2934);
nand UO_437 (O_437,N_2751,N_2443);
nor UO_438 (O_438,N_2675,N_2566);
and UO_439 (O_439,N_2919,N_2520);
and UO_440 (O_440,N_2563,N_2583);
nor UO_441 (O_441,N_2596,N_2716);
xnor UO_442 (O_442,N_2986,N_2597);
nor UO_443 (O_443,N_2863,N_2959);
or UO_444 (O_444,N_2481,N_2545);
and UO_445 (O_445,N_2681,N_2773);
and UO_446 (O_446,N_2777,N_2919);
or UO_447 (O_447,N_2882,N_2946);
and UO_448 (O_448,N_2558,N_2757);
and UO_449 (O_449,N_2467,N_2576);
or UO_450 (O_450,N_2765,N_2740);
and UO_451 (O_451,N_2504,N_2694);
nand UO_452 (O_452,N_2868,N_2980);
and UO_453 (O_453,N_2875,N_2623);
nand UO_454 (O_454,N_2658,N_2901);
nor UO_455 (O_455,N_2620,N_2743);
nand UO_456 (O_456,N_2475,N_2482);
xor UO_457 (O_457,N_2841,N_2442);
nand UO_458 (O_458,N_2515,N_2792);
nor UO_459 (O_459,N_2853,N_2418);
and UO_460 (O_460,N_2434,N_2428);
xnor UO_461 (O_461,N_2890,N_2459);
and UO_462 (O_462,N_2783,N_2811);
and UO_463 (O_463,N_2948,N_2762);
and UO_464 (O_464,N_2453,N_2718);
nand UO_465 (O_465,N_2556,N_2516);
or UO_466 (O_466,N_2618,N_2872);
and UO_467 (O_467,N_2550,N_2463);
and UO_468 (O_468,N_2845,N_2791);
or UO_469 (O_469,N_2702,N_2560);
and UO_470 (O_470,N_2937,N_2816);
nand UO_471 (O_471,N_2998,N_2945);
and UO_472 (O_472,N_2520,N_2411);
nand UO_473 (O_473,N_2975,N_2789);
or UO_474 (O_474,N_2791,N_2533);
nand UO_475 (O_475,N_2568,N_2874);
and UO_476 (O_476,N_2780,N_2711);
nand UO_477 (O_477,N_2883,N_2591);
xnor UO_478 (O_478,N_2586,N_2933);
or UO_479 (O_479,N_2644,N_2499);
nand UO_480 (O_480,N_2502,N_2660);
nand UO_481 (O_481,N_2855,N_2618);
nor UO_482 (O_482,N_2466,N_2931);
nor UO_483 (O_483,N_2567,N_2981);
nor UO_484 (O_484,N_2908,N_2501);
and UO_485 (O_485,N_2590,N_2840);
nor UO_486 (O_486,N_2462,N_2810);
or UO_487 (O_487,N_2993,N_2448);
or UO_488 (O_488,N_2769,N_2586);
nor UO_489 (O_489,N_2680,N_2697);
xnor UO_490 (O_490,N_2727,N_2802);
and UO_491 (O_491,N_2618,N_2746);
or UO_492 (O_492,N_2463,N_2757);
and UO_493 (O_493,N_2669,N_2843);
and UO_494 (O_494,N_2605,N_2651);
nand UO_495 (O_495,N_2487,N_2738);
nand UO_496 (O_496,N_2925,N_2806);
nand UO_497 (O_497,N_2539,N_2987);
nand UO_498 (O_498,N_2580,N_2765);
nand UO_499 (O_499,N_2853,N_2926);
endmodule