module basic_2000_20000_2500_40_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1438,In_1301);
nand U1 (N_1,In_702,In_111);
xor U2 (N_2,In_1667,In_1808);
xor U3 (N_3,In_1799,In_509);
nor U4 (N_4,In_1493,In_1807);
nor U5 (N_5,In_267,In_1423);
nand U6 (N_6,In_335,In_299);
nor U7 (N_7,In_1180,In_633);
and U8 (N_8,In_142,In_1);
nor U9 (N_9,In_1385,In_1855);
nand U10 (N_10,In_1936,In_1823);
nand U11 (N_11,In_1986,In_918);
nor U12 (N_12,In_1514,In_191);
nor U13 (N_13,In_1228,In_1125);
or U14 (N_14,In_1282,In_196);
nand U15 (N_15,In_91,In_1511);
nor U16 (N_16,In_1711,In_1215);
nor U17 (N_17,In_1769,In_210);
nor U18 (N_18,In_1152,In_138);
or U19 (N_19,In_617,In_1346);
nand U20 (N_20,In_1116,In_1285);
or U21 (N_21,In_1941,In_1088);
or U22 (N_22,In_898,In_1457);
nor U23 (N_23,In_480,In_1437);
and U24 (N_24,In_1266,In_1436);
or U25 (N_25,In_1631,In_1107);
nor U26 (N_26,In_1257,In_678);
xnor U27 (N_27,In_1460,In_1742);
xnor U28 (N_28,In_733,In_1970);
or U29 (N_29,In_347,In_51);
nand U30 (N_30,In_1000,In_336);
nor U31 (N_31,In_1313,In_1520);
nand U32 (N_32,In_1656,In_685);
xor U33 (N_33,In_828,In_1448);
nor U34 (N_34,In_893,In_151);
and U35 (N_35,In_1111,In_270);
or U36 (N_36,In_775,In_684);
xnor U37 (N_37,In_1171,In_1381);
xor U38 (N_38,In_739,In_59);
and U39 (N_39,In_653,In_1177);
and U40 (N_40,In_1456,In_533);
and U41 (N_41,In_985,In_1292);
and U42 (N_42,In_174,In_364);
xor U43 (N_43,In_1883,In_885);
nor U44 (N_44,In_557,In_1063);
nor U45 (N_45,In_598,In_212);
nor U46 (N_46,In_49,In_1375);
xor U47 (N_47,In_1622,In_499);
nor U48 (N_48,In_1529,In_322);
nor U49 (N_49,In_376,In_1989);
nand U50 (N_50,In_746,In_200);
nand U51 (N_51,In_1918,In_1492);
nand U52 (N_52,In_1973,In_201);
or U53 (N_53,In_1811,In_492);
xor U54 (N_54,In_1568,In_628);
and U55 (N_55,In_298,In_473);
or U56 (N_56,In_510,In_820);
nand U57 (N_57,In_1078,In_1768);
or U58 (N_58,In_350,In_1021);
xnor U59 (N_59,In_1632,In_120);
nor U60 (N_60,In_1713,In_1519);
xor U61 (N_61,In_1795,In_1666);
xor U62 (N_62,In_1246,In_1148);
nand U63 (N_63,In_253,In_45);
xnor U64 (N_64,In_541,In_891);
nor U65 (N_65,In_221,In_404);
xnor U66 (N_66,In_1310,In_1389);
nor U67 (N_67,In_920,In_538);
and U68 (N_68,In_1422,In_445);
or U69 (N_69,In_469,In_1749);
nand U70 (N_70,In_1383,In_1717);
nand U71 (N_71,In_324,In_103);
nor U72 (N_72,In_965,In_1673);
and U73 (N_73,In_652,In_260);
and U74 (N_74,In_1988,In_1894);
or U75 (N_75,In_147,In_986);
nand U76 (N_76,In_1040,In_1706);
and U77 (N_77,In_622,In_1930);
or U78 (N_78,In_1149,In_1583);
nor U79 (N_79,In_1851,In_709);
nand U80 (N_80,In_1193,In_495);
nand U81 (N_81,In_996,In_358);
xor U82 (N_82,In_1874,In_351);
xnor U83 (N_83,In_719,In_1834);
nor U84 (N_84,In_386,In_454);
or U85 (N_85,In_1934,In_1710);
nor U86 (N_86,In_1562,In_1138);
nor U87 (N_87,In_798,In_231);
nand U88 (N_88,In_1898,In_361);
or U89 (N_89,In_553,In_1353);
nand U90 (N_90,In_136,In_1736);
or U91 (N_91,In_1262,In_356);
nand U92 (N_92,In_214,In_160);
and U93 (N_93,In_794,In_360);
xor U94 (N_94,In_400,In_423);
xnor U95 (N_95,In_688,In_1565);
nand U96 (N_96,In_1600,In_50);
and U97 (N_97,In_512,In_303);
xor U98 (N_98,In_846,In_1143);
nand U99 (N_99,In_1482,In_693);
and U100 (N_100,In_1065,In_888);
and U101 (N_101,In_104,In_836);
and U102 (N_102,In_1951,In_419);
xnor U103 (N_103,In_602,In_814);
and U104 (N_104,In_877,In_326);
or U105 (N_105,In_1850,In_1252);
nor U106 (N_106,In_1651,In_25);
nor U107 (N_107,In_812,In_455);
and U108 (N_108,In_695,In_823);
xor U109 (N_109,In_385,In_525);
and U110 (N_110,In_433,In_1464);
xnor U111 (N_111,In_1269,In_1380);
and U112 (N_112,In_1554,In_1889);
or U113 (N_113,In_1289,In_1860);
nor U114 (N_114,In_1046,In_663);
and U115 (N_115,In_1497,In_242);
nor U116 (N_116,In_611,In_421);
or U117 (N_117,In_1619,In_1868);
or U118 (N_118,In_283,In_1516);
nor U119 (N_119,In_713,In_18);
nand U120 (N_120,In_1053,In_306);
nand U121 (N_121,In_1210,In_1390);
or U122 (N_122,In_964,In_1599);
or U123 (N_123,In_1841,In_1169);
or U124 (N_124,In_981,In_1420);
nor U125 (N_125,In_1196,In_1816);
xnor U126 (N_126,In_970,In_285);
nand U127 (N_127,In_61,In_821);
nor U128 (N_128,In_313,In_62);
xor U129 (N_129,In_873,In_531);
nand U130 (N_130,In_1032,In_268);
nand U131 (N_131,In_1140,In_722);
and U132 (N_132,In_1926,In_573);
xnor U133 (N_133,In_78,In_121);
and U134 (N_134,In_378,In_81);
xor U135 (N_135,In_1567,In_1778);
and U136 (N_136,In_1178,In_184);
xnor U137 (N_137,In_668,In_102);
nor U138 (N_138,In_799,In_671);
nand U139 (N_139,In_758,In_990);
xnor U140 (N_140,In_1638,In_1853);
and U141 (N_141,In_131,In_1703);
nand U142 (N_142,In_1893,In_1294);
and U143 (N_143,In_1818,In_853);
or U144 (N_144,In_1740,In_1245);
nand U145 (N_145,In_521,In_215);
and U146 (N_146,In_1333,In_1884);
xnor U147 (N_147,In_1126,In_1056);
nor U148 (N_148,In_1837,In_323);
nor U149 (N_149,In_1344,In_1549);
or U150 (N_150,In_1879,In_12);
and U151 (N_151,In_883,In_1185);
nor U152 (N_152,In_1683,In_1428);
nor U153 (N_153,In_5,In_1015);
nor U154 (N_154,In_367,In_900);
xnor U155 (N_155,In_1253,In_278);
xor U156 (N_156,In_1907,In_1560);
xnor U157 (N_157,In_1888,In_1017);
and U158 (N_158,In_987,In_676);
nor U159 (N_159,In_1872,In_1163);
nor U160 (N_160,In_320,In_730);
xor U161 (N_161,In_932,In_570);
nor U162 (N_162,In_1357,In_1668);
or U163 (N_163,In_281,In_1770);
xnor U164 (N_164,In_1098,In_1956);
nand U165 (N_165,In_664,In_2);
nor U166 (N_166,In_884,In_641);
and U167 (N_167,In_1296,In_337);
nand U168 (N_168,In_1960,In_1787);
nand U169 (N_169,In_1329,In_1038);
xnor U170 (N_170,In_631,In_763);
xor U171 (N_171,In_489,In_1513);
and U172 (N_172,In_1217,In_610);
nor U173 (N_173,In_1101,In_1755);
or U174 (N_174,In_1203,In_1582);
nand U175 (N_175,In_672,In_1862);
xor U176 (N_176,In_272,In_1921);
xor U177 (N_177,In_1722,In_46);
or U178 (N_178,In_575,In_437);
xnor U179 (N_179,In_946,In_1904);
nand U180 (N_180,In_694,In_529);
and U181 (N_181,In_408,In_186);
nor U182 (N_182,In_1280,In_971);
nand U183 (N_183,In_1763,In_349);
nand U184 (N_184,In_1084,In_1812);
or U185 (N_185,In_1335,In_1972);
nor U186 (N_186,In_863,In_1489);
nor U187 (N_187,In_235,In_1544);
and U188 (N_188,In_1935,In_57);
nor U189 (N_189,In_1451,In_600);
xor U190 (N_190,In_861,In_982);
xnor U191 (N_191,In_1601,In_1320);
xor U192 (N_192,In_1961,In_1848);
nor U193 (N_193,In_697,In_1846);
xnor U194 (N_194,In_1629,In_1539);
and U195 (N_195,In_983,In_1355);
xnor U196 (N_196,In_1446,In_872);
nor U197 (N_197,In_1145,In_485);
and U198 (N_198,In_618,In_84);
and U199 (N_199,In_545,In_1096);
xnor U200 (N_200,In_569,In_774);
or U201 (N_201,In_205,In_113);
or U202 (N_202,In_657,In_745);
nor U203 (N_203,In_917,In_647);
xnor U204 (N_204,In_804,In_751);
nand U205 (N_205,In_339,In_319);
nand U206 (N_206,In_1982,In_1068);
nand U207 (N_207,In_1892,In_208);
xor U208 (N_208,In_583,In_457);
xor U209 (N_209,In_706,In_1831);
nor U210 (N_210,In_1728,In_170);
xor U211 (N_211,In_1662,In_1166);
nor U212 (N_212,In_301,In_1009);
nor U213 (N_213,In_1449,In_241);
nand U214 (N_214,In_844,In_162);
nor U215 (N_215,In_1877,In_1933);
and U216 (N_216,In_118,In_422);
nor U217 (N_217,In_345,In_1351);
nand U218 (N_218,In_1114,In_1942);
and U219 (N_219,In_183,In_239);
or U220 (N_220,In_795,In_1358);
nor U221 (N_221,In_1275,In_659);
nand U222 (N_222,In_1596,In_166);
or U223 (N_223,In_937,In_773);
nor U224 (N_224,In_238,In_1043);
and U225 (N_225,In_1191,In_651);
or U226 (N_226,In_1238,In_1917);
or U227 (N_227,In_851,In_1546);
xor U228 (N_228,In_86,In_383);
or U229 (N_229,In_699,In_1240);
nand U230 (N_230,In_1517,In_1429);
nor U231 (N_231,In_309,In_998);
nand U232 (N_232,In_27,In_686);
nand U233 (N_233,In_802,In_466);
xnor U234 (N_234,In_1966,In_670);
nand U235 (N_235,In_1427,In_1815);
nor U236 (N_236,In_137,In_1648);
xnor U237 (N_237,In_1223,In_748);
or U238 (N_238,In_737,In_1750);
xor U239 (N_239,In_1397,In_950);
and U240 (N_240,In_691,In_951);
and U241 (N_241,In_1532,In_537);
xnor U242 (N_242,In_910,In_1241);
nand U243 (N_243,In_1198,In_771);
nand U244 (N_244,In_1827,In_188);
nand U245 (N_245,In_744,In_1655);
nor U246 (N_246,In_1391,In_82);
and U247 (N_247,In_1665,In_1268);
xnor U248 (N_248,In_551,In_467);
and U249 (N_249,In_1573,In_426);
or U250 (N_250,In_225,In_1500);
nand U251 (N_251,In_1331,In_742);
xnor U252 (N_252,In_1521,In_587);
or U253 (N_253,In_1412,In_895);
nand U254 (N_254,In_752,In_16);
or U255 (N_255,In_1471,In_148);
and U256 (N_256,In_1479,In_70);
nand U257 (N_257,In_593,In_1948);
or U258 (N_258,In_1336,In_89);
and U259 (N_259,In_1943,In_585);
xnor U260 (N_260,In_1817,In_1641);
nand U261 (N_261,In_1744,In_1552);
nor U262 (N_262,In_178,In_714);
nor U263 (N_263,In_958,In_1415);
nand U264 (N_264,In_346,In_978);
nand U265 (N_265,In_1356,In_829);
nor U266 (N_266,In_1099,In_54);
nand U267 (N_267,In_390,In_1897);
nand U268 (N_268,In_1974,In_439);
xor U269 (N_269,In_332,In_1833);
xor U270 (N_270,In_1944,In_1488);
or U271 (N_271,In_1503,In_348);
and U272 (N_272,In_441,In_1709);
or U273 (N_273,In_747,In_517);
nor U274 (N_274,In_394,In_479);
nand U275 (N_275,In_743,In_247);
or U276 (N_276,In_1653,In_1175);
xor U277 (N_277,In_1129,In_1782);
and U278 (N_278,In_406,In_1213);
xnor U279 (N_279,In_1558,In_1737);
or U280 (N_280,In_584,In_740);
nand U281 (N_281,In_1663,In_1761);
and U282 (N_282,In_1279,In_1866);
nand U283 (N_283,In_1458,In_667);
or U284 (N_284,In_988,In_172);
and U285 (N_285,In_444,In_734);
nor U286 (N_286,In_1146,In_1259);
xnor U287 (N_287,In_705,In_1077);
xnor U288 (N_288,In_1105,In_892);
xnor U289 (N_289,In_616,In_446);
nor U290 (N_290,In_1743,In_416);
nand U291 (N_291,In_399,In_1528);
xnor U292 (N_292,In_607,In_1142);
or U293 (N_293,In_374,In_1055);
nand U294 (N_294,In_26,In_32);
xnor U295 (N_295,In_44,In_805);
nand U296 (N_296,In_757,In_1263);
and U297 (N_297,In_1414,In_604);
nor U298 (N_298,In_152,In_357);
nor U299 (N_299,In_109,In_1954);
and U300 (N_300,In_377,In_803);
nand U301 (N_301,In_1490,In_1875);
nand U302 (N_302,In_126,In_1480);
xor U303 (N_303,In_199,In_1929);
and U304 (N_304,In_1192,In_721);
or U305 (N_305,In_1374,In_843);
and U306 (N_306,In_1165,In_1463);
and U307 (N_307,In_848,In_1589);
nand U308 (N_308,In_1396,In_1216);
and U309 (N_309,In_1157,In_1920);
nor U310 (N_310,In_1388,In_1571);
or U311 (N_311,In_1677,In_1977);
nand U312 (N_312,In_219,In_655);
nor U313 (N_313,In_24,In_1825);
xnor U314 (N_314,In_1981,In_98);
xnor U315 (N_315,In_720,In_1797);
nand U316 (N_316,In_1630,In_1908);
or U317 (N_317,In_1221,In_1845);
xor U318 (N_318,In_902,In_761);
nand U319 (N_319,In_468,In_1828);
nand U320 (N_320,In_1802,In_430);
and U321 (N_321,In_601,In_1510);
xor U322 (N_322,In_52,In_881);
nor U323 (N_323,In_770,In_535);
or U324 (N_324,In_1820,In_933);
nand U325 (N_325,In_1117,In_1739);
nand U326 (N_326,In_1945,In_680);
and U327 (N_327,In_262,In_966);
nand U328 (N_328,In_603,In_1996);
nor U329 (N_329,In_1407,In_1435);
nand U330 (N_330,In_882,In_236);
and U331 (N_331,In_1804,In_1564);
nand U332 (N_332,In_943,In_269);
and U333 (N_333,In_1984,In_1729);
or U334 (N_334,In_286,In_1450);
nor U335 (N_335,In_198,In_1037);
nor U336 (N_336,In_108,In_976);
nor U337 (N_337,In_418,In_1591);
nand U338 (N_338,In_1167,In_935);
xor U339 (N_339,In_340,In_1234);
xor U340 (N_340,In_1443,In_67);
nand U341 (N_341,In_154,In_1604);
nor U342 (N_342,In_329,In_3);
nand U343 (N_343,In_591,In_658);
xor U344 (N_344,In_1326,In_627);
or U345 (N_345,In_1071,In_776);
xor U346 (N_346,In_1012,In_1870);
or U347 (N_347,In_1712,In_1311);
xnor U348 (N_348,In_187,In_1179);
nand U349 (N_349,In_1515,In_769);
xnor U350 (N_350,In_1258,In_1295);
nand U351 (N_351,In_1971,In_1212);
and U352 (N_352,In_963,In_19);
xor U353 (N_353,In_1849,In_632);
nor U354 (N_354,In_1990,In_107);
and U355 (N_355,In_330,In_1686);
and U356 (N_356,In_1161,In_831);
nand U357 (N_357,In_1647,In_417);
nor U358 (N_358,In_195,In_1014);
or U359 (N_359,In_1556,In_487);
nand U360 (N_360,In_650,In_1890);
or U361 (N_361,In_393,In_99);
xnor U362 (N_362,In_732,In_1242);
nor U363 (N_363,In_1139,In_1752);
nor U364 (N_364,In_1200,In_37);
or U365 (N_365,In_503,In_167);
nor U366 (N_366,In_265,In_700);
or U367 (N_367,In_1983,In_646);
nor U368 (N_368,In_1350,In_424);
nor U369 (N_369,In_576,In_1994);
nor U370 (N_370,In_547,In_1170);
nand U371 (N_371,In_1939,In_42);
nor U372 (N_372,In_133,In_994);
nor U373 (N_373,In_755,In_334);
nand U374 (N_374,In_1657,In_1110);
xnor U375 (N_375,In_1847,In_405);
and U376 (N_376,In_88,In_1688);
xor U377 (N_377,In_1337,In_481);
xor U378 (N_378,In_922,In_1016);
nor U379 (N_379,In_431,In_486);
and U380 (N_380,In_1792,In_1617);
nand U381 (N_381,In_915,In_500);
nor U382 (N_382,In_1842,In_930);
or U383 (N_383,In_1303,In_150);
or U384 (N_384,In_991,In_1704);
nand U385 (N_385,In_683,In_1483);
and U386 (N_386,In_905,In_1635);
nand U387 (N_387,In_343,In_1074);
xor U388 (N_388,In_1810,In_1964);
xnor U389 (N_389,In_925,In_1222);
or U390 (N_390,In_291,In_1499);
nor U391 (N_391,In_724,In_497);
and U392 (N_392,In_380,In_862);
or U393 (N_393,In_1230,In_1132);
or U394 (N_394,In_13,In_1976);
or U395 (N_395,In_279,In_1880);
and U396 (N_396,In_1524,In_692);
or U397 (N_397,In_972,In_682);
and U398 (N_398,In_169,In_1602);
nand U399 (N_399,In_1474,In_1551);
or U400 (N_400,In_245,In_984);
or U401 (N_401,In_85,In_1540);
xnor U402 (N_402,In_728,In_1590);
nand U403 (N_403,In_827,In_1181);
xor U404 (N_404,In_588,In_1561);
and U405 (N_405,In_1211,In_155);
xnor U406 (N_406,In_1720,In_1621);
or U407 (N_407,In_1923,In_1518);
nor U408 (N_408,In_555,In_1727);
xnor U409 (N_409,In_928,In_858);
and U410 (N_410,In_1027,In_1962);
nand U411 (N_411,In_1579,In_665);
and U412 (N_412,In_384,In_211);
or U413 (N_413,In_66,In_1433);
or U414 (N_414,In_163,In_540);
or U415 (N_415,In_1477,In_562);
nand U416 (N_416,In_1594,In_1857);
or U417 (N_417,In_1530,In_302);
or U418 (N_418,In_1119,In_252);
and U419 (N_419,In_1865,In_1618);
xnor U420 (N_420,In_673,In_944);
nand U421 (N_421,In_472,In_741);
nand U422 (N_422,In_780,In_941);
nand U423 (N_423,In_1566,In_300);
nand U424 (N_424,In_1867,In_55);
and U425 (N_425,In_1283,In_161);
or U426 (N_426,In_271,In_1045);
and U427 (N_427,In_1398,In_127);
xnor U428 (N_428,In_203,In_1419);
nor U429 (N_429,In_1542,In_1735);
nand U430 (N_430,In_599,In_1302);
and U431 (N_431,In_1751,In_274);
and U432 (N_432,In_577,In_927);
nand U433 (N_433,In_1620,In_1975);
xor U434 (N_434,In_619,In_1771);
nor U435 (N_435,In_1915,In_1122);
xnor U436 (N_436,In_797,In_1224);
or U437 (N_437,In_666,In_36);
nand U438 (N_438,In_243,In_629);
or U439 (N_439,In_75,In_234);
or U440 (N_440,In_228,In_114);
nor U441 (N_441,In_1286,In_1035);
or U442 (N_442,In_1254,In_1156);
and U443 (N_443,In_11,In_1784);
and U444 (N_444,In_1343,In_1592);
nor U445 (N_445,In_766,In_1284);
nand U446 (N_446,In_310,In_173);
nor U447 (N_447,In_609,In_608);
or U448 (N_448,In_936,In_1059);
xor U449 (N_449,In_559,In_975);
nor U450 (N_450,In_777,In_402);
nor U451 (N_451,In_463,In_572);
nor U452 (N_452,In_1066,In_96);
or U453 (N_453,In_560,In_1197);
and U454 (N_454,In_564,In_1475);
nand U455 (N_455,In_1327,In_40);
xor U456 (N_456,In_428,In_914);
nor U457 (N_457,In_1644,In_1937);
and U458 (N_458,In_738,In_1553);
nand U459 (N_459,In_817,In_1288);
xor U460 (N_460,In_1010,In_206);
nand U461 (N_461,In_1642,In_362);
and U462 (N_462,In_217,In_1723);
xor U463 (N_463,In_122,In_842);
nand U464 (N_464,In_879,In_22);
or U465 (N_465,In_1376,In_1793);
and U466 (N_466,In_674,In_1947);
nor U467 (N_467,In_185,In_1229);
or U468 (N_468,In_1330,In_1840);
xor U469 (N_469,In_1495,In_635);
nand U470 (N_470,In_623,In_1664);
xor U471 (N_471,In_1725,In_1349);
xnor U472 (N_472,In_139,In_1698);
xnor U473 (N_473,In_952,In_1109);
and U474 (N_474,In_1931,In_909);
nand U475 (N_475,In_876,In_1721);
and U476 (N_476,In_1031,In_1512);
nand U477 (N_477,In_707,In_1593);
and U478 (N_478,In_1748,In_95);
xnor U479 (N_479,In_1575,In_1758);
and U480 (N_480,In_1762,In_115);
nor U481 (N_481,In_1025,In_1083);
xor U482 (N_482,In_1441,In_589);
or U483 (N_483,In_1069,In_1261);
nor U484 (N_484,In_1048,In_1745);
nor U485 (N_485,In_1123,In_387);
xor U486 (N_486,In_840,In_425);
nand U487 (N_487,In_1946,In_193);
and U488 (N_488,In_1442,In_259);
nor U489 (N_489,In_1580,In_1626);
nor U490 (N_490,In_865,In_341);
and U491 (N_491,In_1886,In_352);
and U492 (N_492,In_913,In_237);
and U493 (N_493,In_1226,In_207);
or U494 (N_494,In_294,In_1603);
xor U495 (N_495,In_1522,In_1154);
or U496 (N_496,In_100,In_1406);
and U497 (N_497,In_940,In_1715);
xnor U498 (N_498,In_1121,In_415);
nand U499 (N_499,In_1563,In_548);
xnor U500 (N_500,N_96,N_265);
and U501 (N_501,N_150,N_287);
xnor U502 (N_502,In_1627,N_400);
or U503 (N_503,In_1255,N_203);
nand U504 (N_504,In_783,In_491);
nand U505 (N_505,N_40,In_1650);
nor U506 (N_506,N_484,In_1678);
or U507 (N_507,N_87,In_1318);
nand U508 (N_508,In_209,In_396);
nand U509 (N_509,In_1608,In_1455);
and U510 (N_510,In_1424,N_389);
nand U511 (N_511,In_1696,In_894);
nand U512 (N_512,In_838,In_477);
or U513 (N_513,In_867,In_64);
xnor U514 (N_514,N_470,In_33);
and U515 (N_515,N_312,In_165);
or U516 (N_516,In_1791,In_703);
or U517 (N_517,In_1136,In_1260);
nand U518 (N_518,In_369,N_384);
xnor U519 (N_519,In_1033,In_822);
or U520 (N_520,In_1537,In_449);
nand U521 (N_521,In_1141,In_566);
and U522 (N_522,In_1218,In_344);
and U523 (N_523,In_1001,In_1274);
or U524 (N_524,In_1578,N_156);
and U525 (N_525,In_1669,In_1120);
nand U526 (N_526,N_410,In_1328);
xor U527 (N_527,In_496,In_516);
and U528 (N_528,N_187,N_390);
xor U529 (N_529,In_1271,In_871);
nor U530 (N_530,In_29,In_164);
or U531 (N_531,In_801,N_401);
xor U532 (N_532,In_1876,N_252);
nor U533 (N_533,N_320,In_1369);
or U534 (N_534,In_875,N_221);
nor U535 (N_535,In_168,N_446);
xor U536 (N_536,N_223,In_788);
nor U537 (N_537,N_309,In_1029);
and U538 (N_538,N_109,N_247);
or U539 (N_539,In_1790,N_119);
nand U540 (N_540,In_621,In_1298);
xnor U541 (N_541,In_1836,N_245);
nand U542 (N_542,In_955,N_378);
xnor U543 (N_543,In_1023,N_84);
nand U544 (N_544,In_727,N_367);
or U545 (N_545,N_493,In_660);
xor U546 (N_546,In_420,In_263);
and U547 (N_547,In_90,In_1718);
xnor U548 (N_548,N_167,In_1363);
xor U549 (N_549,In_554,In_786);
and U550 (N_550,In_1018,In_511);
nand U551 (N_551,N_339,In_1155);
nand U552 (N_552,In_1891,In_501);
xnor U553 (N_553,In_1339,In_6);
and U554 (N_554,N_362,N_462);
or U555 (N_555,N_424,In_1885);
or U556 (N_556,In_149,N_127);
nor U557 (N_557,In_1487,In_1624);
nor U558 (N_558,N_475,N_435);
xor U559 (N_559,N_409,In_23);
and U560 (N_560,In_1277,N_440);
and U561 (N_561,In_1201,In_954);
xor U562 (N_562,N_59,In_1095);
nand U563 (N_563,N_170,In_857);
or U564 (N_564,N_26,In_389);
nand U565 (N_565,In_1411,In_712);
and U566 (N_566,In_1965,In_926);
xor U567 (N_567,In_257,In_440);
xor U568 (N_568,In_1468,In_992);
and U569 (N_569,In_1072,In_1679);
and U570 (N_570,In_125,In_1425);
xnor U571 (N_571,In_1076,In_1094);
and U572 (N_572,In_789,N_215);
and U573 (N_573,In_1452,In_837);
xnor U574 (N_574,N_193,In_1950);
nor U575 (N_575,N_169,N_295);
nand U576 (N_576,N_464,N_492);
xnor U577 (N_577,N_259,In_471);
or U578 (N_578,In_961,In_1801);
nor U579 (N_579,In_474,In_1979);
and U580 (N_580,In_931,In_379);
nand U581 (N_581,N_382,In_1633);
nand U582 (N_582,N_346,N_455);
xnor U583 (N_583,In_287,In_305);
xor U584 (N_584,In_307,In_1133);
nor U585 (N_585,In_662,In_534);
nand U586 (N_586,In_1124,In_764);
and U587 (N_587,In_1645,In_856);
xnor U588 (N_588,In_1237,In_1293);
and U589 (N_589,N_113,N_11);
and U590 (N_590,N_333,In_850);
or U591 (N_591,N_107,In_597);
or U592 (N_592,N_199,In_1087);
xor U593 (N_593,N_327,In_1584);
nor U594 (N_594,In_1684,In_1176);
or U595 (N_595,In_292,In_197);
nor U596 (N_596,In_1305,In_813);
and U597 (N_597,N_148,In_1239);
nor U598 (N_598,In_21,In_1634);
nand U599 (N_599,N_176,In_502);
xor U600 (N_600,In_1097,In_1545);
nor U601 (N_601,In_1922,In_896);
or U602 (N_602,In_1674,In_1912);
and U603 (N_603,N_190,N_64);
xnor U604 (N_604,N_31,In_453);
nor U605 (N_605,N_108,N_73);
xnor U606 (N_606,N_208,In_48);
or U607 (N_607,In_792,In_1643);
xor U608 (N_608,N_388,In_1557);
nor U609 (N_609,In_249,In_1478);
and U610 (N_610,In_395,In_74);
or U611 (N_611,In_959,In_993);
nand U612 (N_612,In_432,In_1534);
or U613 (N_613,N_416,In_580);
and U614 (N_614,N_240,N_386);
nor U615 (N_615,In_498,N_92);
xor U616 (N_616,In_1410,N_430);
nand U617 (N_617,N_284,In_1164);
nor U618 (N_618,N_100,In_407);
nor U619 (N_619,N_488,In_175);
and U620 (N_620,In_452,In_1779);
or U621 (N_621,In_1625,N_103);
nor U622 (N_622,N_68,In_482);
nand U623 (N_623,N_453,N_258);
nand U624 (N_624,In_296,N_10);
nor U625 (N_625,In_1227,In_1135);
and U626 (N_626,In_1134,N_249);
nand U627 (N_627,In_1746,N_291);
or U628 (N_628,In_1306,In_1184);
xnor U629 (N_629,N_229,In_1597);
xnor U630 (N_630,N_336,In_488);
or U631 (N_631,N_352,In_1395);
nor U632 (N_632,In_1409,In_1538);
or U633 (N_633,In_143,In_282);
or U634 (N_634,In_1671,In_436);
nand U635 (N_635,In_465,In_297);
nor U636 (N_636,In_38,In_644);
xnor U637 (N_637,N_374,N_225);
nand U638 (N_638,In_847,N_219);
nor U639 (N_639,In_772,In_79);
nor U640 (N_640,N_306,N_393);
xor U641 (N_641,In_1090,N_13);
or U642 (N_642,In_244,In_768);
nor U643 (N_643,In_1322,In_1467);
and U644 (N_644,In_93,N_448);
xor U645 (N_645,In_119,N_359);
xnor U646 (N_646,In_1439,In_1440);
or U647 (N_647,N_60,In_366);
or U648 (N_648,N_426,In_1186);
xor U649 (N_649,N_341,In_9);
or U650 (N_650,In_1786,N_185);
or U651 (N_651,N_88,In_756);
or U652 (N_652,In_1753,In_1403);
or U653 (N_653,In_1444,In_194);
or U654 (N_654,In_1049,N_348);
nand U655 (N_655,N_330,In_723);
or U656 (N_656,N_372,In_620);
nand U657 (N_657,N_37,In_34);
or U658 (N_658,In_216,In_957);
nand U659 (N_659,N_174,In_859);
nor U660 (N_660,N_271,In_373);
xnor U661 (N_661,In_854,In_130);
or U662 (N_662,N_105,N_179);
nand U663 (N_663,In_1822,In_1764);
nand U664 (N_664,In_832,N_487);
nor U665 (N_665,N_454,N_180);
xnor U666 (N_666,N_160,N_181);
or U667 (N_667,N_282,N_344);
nand U668 (N_668,N_52,N_286);
or U669 (N_669,In_141,In_594);
nor U670 (N_670,N_217,In_227);
xnor U671 (N_671,In_1741,In_967);
xor U672 (N_672,In_1509,N_451);
or U673 (N_673,In_1800,In_1368);
or U674 (N_674,In_0,In_461);
and U675 (N_675,In_565,In_675);
nor U676 (N_676,N_266,N_444);
nand U677 (N_677,In_824,In_226);
nand U678 (N_678,In_1598,In_1334);
nor U679 (N_679,N_204,In_1757);
and U680 (N_680,In_921,In_679);
xnor U681 (N_681,In_1637,N_99);
and U682 (N_682,In_1773,N_421);
nor U683 (N_683,In_1382,N_67);
xnor U684 (N_684,In_785,In_916);
nor U685 (N_685,In_266,N_261);
xnor U686 (N_686,In_949,In_1207);
or U687 (N_687,In_1607,In_1008);
xor U688 (N_688,N_41,In_919);
or U689 (N_689,N_267,In_552);
xor U690 (N_690,N_283,In_1555);
nand U691 (N_691,N_407,In_1691);
nand U692 (N_692,N_294,In_1251);
nor U693 (N_693,In_1308,N_269);
nand U694 (N_694,In_1312,N_315);
nand U695 (N_695,In_1062,In_478);
xor U696 (N_696,In_578,In_1030);
nand U697 (N_697,In_1405,In_736);
nor U698 (N_698,N_276,N_93);
xor U699 (N_699,In_852,In_806);
xor U700 (N_700,In_1916,N_387);
nor U701 (N_701,In_359,N_370);
xor U702 (N_702,N_48,N_21);
nand U703 (N_703,In_135,In_634);
nor U704 (N_704,In_1348,N_1);
xnor U705 (N_705,In_327,N_342);
nor U706 (N_706,N_23,N_355);
nand U707 (N_707,N_325,In_1051);
nand U708 (N_708,In_312,In_1220);
and U709 (N_709,In_1993,In_20);
nor U710 (N_710,N_201,N_209);
and U711 (N_711,In_1927,N_433);
xor U712 (N_712,N_131,In_753);
xnor U713 (N_713,N_117,In_874);
and U714 (N_714,In_1780,N_274);
nand U715 (N_715,In_1264,N_303);
nand U716 (N_716,In_878,N_255);
and U717 (N_717,In_333,In_1527);
nor U718 (N_718,N_377,In_1151);
nand U719 (N_719,In_1233,In_1507);
nand U720 (N_720,N_395,In_1826);
nor U721 (N_721,In_1777,N_438);
or U722 (N_722,In_220,N_289);
or U723 (N_723,In_413,In_1680);
or U724 (N_724,In_760,In_1814);
or U725 (N_725,In_1144,In_765);
and U726 (N_726,In_1208,N_66);
and U727 (N_727,In_779,In_1640);
nand U728 (N_728,N_24,In_398);
or U729 (N_729,In_30,In_796);
xor U730 (N_730,In_1387,N_159);
and U731 (N_731,N_236,In_464);
nand U732 (N_732,In_1394,In_1636);
xnor U733 (N_733,In_1569,In_835);
nand U734 (N_734,N_461,In_1789);
nand U735 (N_735,In_708,In_960);
nor U736 (N_736,In_1794,N_290);
xor U737 (N_737,In_1402,In_1028);
xnor U738 (N_738,N_200,In_280);
nand U739 (N_739,N_121,In_1469);
and U740 (N_740,N_51,N_63);
and U741 (N_741,In_661,In_1652);
nor U742 (N_742,N_129,N_495);
xor U743 (N_743,In_716,N_222);
and U744 (N_744,In_1299,N_301);
and U745 (N_745,N_126,N_293);
xnor U746 (N_746,N_54,In_456);
or U747 (N_747,N_441,In_605);
or U748 (N_748,In_76,N_232);
nor U749 (N_749,In_1189,In_1531);
and U750 (N_750,In_1054,In_530);
nand U751 (N_751,In_1007,In_1118);
and U752 (N_752,N_468,In_1900);
and U753 (N_753,In_365,In_288);
and U754 (N_754,In_1462,In_1805);
or U755 (N_755,In_134,In_1508);
xor U756 (N_756,In_1526,In_1287);
nor U757 (N_757,In_539,In_317);
xor U758 (N_758,In_784,In_614);
and U759 (N_759,In_1162,In_750);
nor U760 (N_760,In_1501,In_232);
or U761 (N_761,In_726,In_1104);
xnor U762 (N_762,In_1160,In_520);
or U763 (N_763,In_1050,In_1506);
nand U764 (N_764,In_1235,N_347);
and U765 (N_765,In_1070,N_288);
nor U766 (N_766,In_811,In_1861);
nor U767 (N_767,N_182,In_519);
xnor U768 (N_768,In_1843,N_439);
xnor U769 (N_769,In_948,In_1896);
or U770 (N_770,N_244,In_908);
xor U771 (N_771,N_34,In_275);
or U772 (N_772,In_442,N_412);
xnor U773 (N_773,In_1365,In_1194);
xnor U774 (N_774,N_499,In_1587);
or U775 (N_775,In_1089,In_458);
or U776 (N_776,In_177,In_483);
or U777 (N_777,In_87,In_1714);
nor U778 (N_778,N_429,In_429);
or U779 (N_779,In_953,N_80);
or U780 (N_780,In_1225,In_1491);
nand U781 (N_781,In_897,N_162);
and U782 (N_782,In_248,In_254);
and U783 (N_783,In_1057,N_465);
or U784 (N_784,N_145,In_869);
xor U785 (N_785,N_186,In_1595);
and U786 (N_786,In_1485,In_816);
and U787 (N_787,In_1660,In_1244);
xnor U788 (N_788,N_220,In_1980);
nor U789 (N_789,N_411,In_1699);
or U790 (N_790,N_278,In_1250);
or U791 (N_791,In_1052,In_1819);
or U792 (N_792,N_144,In_1371);
nor U793 (N_793,N_413,N_497);
and U794 (N_794,In_1685,N_469);
or U795 (N_795,In_945,In_582);
or U796 (N_796,N_124,In_1803);
nand U797 (N_797,In_116,In_1086);
xnor U798 (N_798,N_381,N_254);
and U799 (N_799,N_164,N_489);
or U800 (N_800,N_62,In_443);
nor U801 (N_801,In_1577,In_1955);
and U802 (N_802,N_420,In_97);
nor U803 (N_803,N_304,In_912);
nand U804 (N_804,In_1024,N_43);
or U805 (N_805,N_397,In_1731);
nor U806 (N_806,N_414,N_246);
xnor U807 (N_807,N_205,In_354);
nor U808 (N_808,In_513,In_818);
or U809 (N_809,In_371,In_1366);
nand U810 (N_810,In_1417,In_1073);
nor U811 (N_811,In_1342,In_1319);
or U812 (N_812,In_855,N_243);
and U813 (N_813,In_1957,N_166);
nand U814 (N_814,In_980,In_157);
xnor U815 (N_815,N_373,In_615);
and U816 (N_816,N_329,N_7);
and U817 (N_817,N_38,N_196);
nor U818 (N_818,In_973,In_880);
or U819 (N_819,In_1019,In_363);
or U820 (N_820,N_422,In_1159);
and U821 (N_821,In_284,N_171);
or U822 (N_822,In_1281,In_654);
or U823 (N_823,In_1168,In_1465);
xor U824 (N_824,N_172,In_314);
or U825 (N_825,N_71,N_298);
and U826 (N_826,In_596,In_1209);
xnor U827 (N_827,In_230,In_527);
nor U828 (N_828,In_1199,N_3);
and U829 (N_829,In_1999,In_1364);
xnor U830 (N_830,N_0,In_1061);
nor U831 (N_831,In_1967,In_1701);
and U832 (N_832,In_192,In_255);
or U833 (N_833,In_1370,N_415);
and U834 (N_834,In_1536,N_218);
and U835 (N_835,N_33,In_1998);
xnor U836 (N_836,In_397,N_53);
nand U837 (N_837,In_1338,In_625);
and U838 (N_838,In_1687,In_637);
and U839 (N_839,N_134,In_1498);
nor U840 (N_840,N_118,In_1494);
nor U841 (N_841,N_189,In_793);
nand U842 (N_842,N_317,N_57);
xnor U843 (N_843,N_406,In_1060);
nand U844 (N_844,In_1585,In_696);
nor U845 (N_845,In_71,In_179);
and U846 (N_846,N_157,In_754);
xnor U847 (N_847,N_272,In_10);
xnor U848 (N_848,In_938,N_47);
or U849 (N_849,In_145,In_68);
xor U850 (N_850,In_1588,In_1459);
xor U851 (N_851,N_458,N_360);
and U852 (N_852,In_1785,In_701);
or U853 (N_853,In_546,In_1902);
or U854 (N_854,N_365,In_1612);
xor U855 (N_855,In_979,In_1570);
and U856 (N_856,N_314,In_808);
nor U857 (N_857,In_514,In_642);
or U858 (N_858,In_1987,In_995);
nor U859 (N_859,N_228,N_296);
and U860 (N_860,N_163,N_383);
xnor U861 (N_861,In_53,In_1102);
and U862 (N_862,In_636,N_483);
nand U863 (N_863,In_251,In_1919);
nand U864 (N_864,In_1581,N_78);
or U865 (N_865,In_677,N_340);
or U866 (N_866,In_1174,N_178);
and U867 (N_867,N_443,In_1681);
and U868 (N_868,N_268,In_447);
xor U869 (N_869,In_250,In_787);
or U870 (N_870,In_132,In_1899);
xnor U871 (N_871,In_1767,N_227);
or U872 (N_872,In_94,In_735);
nand U873 (N_873,N_4,In_1127);
and U874 (N_874,N_89,In_1978);
or U875 (N_875,N_486,In_1496);
nor U876 (N_876,N_280,In_342);
and U877 (N_877,N_292,In_1882);
xor U878 (N_878,In_1058,In_273);
or U879 (N_879,N_358,N_285);
or U880 (N_880,N_310,In_1705);
and U881 (N_881,N_146,In_586);
and U882 (N_882,In_825,N_471);
xnor U883 (N_883,N_116,In_1473);
and U884 (N_884,In_826,In_1004);
and U885 (N_885,In_1434,In_1361);
xnor U886 (N_886,N_2,In_410);
or U887 (N_887,N_343,In_579);
nand U888 (N_888,N_212,In_28);
or U889 (N_889,In_246,In_1856);
xor U890 (N_890,In_1659,N_322);
or U891 (N_891,In_176,In_1548);
xor U892 (N_892,N_357,In_1002);
xnor U893 (N_893,N_494,N_279);
or U894 (N_894,In_1147,In_1400);
nor U895 (N_895,In_180,In_1307);
and U896 (N_896,N_307,In_315);
and U897 (N_897,N_17,N_375);
and U898 (N_898,In_1997,N_55);
nor U899 (N_899,In_1039,In_1672);
xor U900 (N_900,N_74,N_136);
nand U901 (N_901,In_190,N_195);
or U902 (N_902,In_864,In_450);
xnor U903 (N_903,In_401,In_470);
or U904 (N_904,In_718,In_409);
nor U905 (N_905,In_1386,N_366);
xor U906 (N_906,N_132,In_129);
nor U907 (N_907,In_1265,N_299);
and U908 (N_908,In_1707,In_849);
xnor U909 (N_909,In_1085,N_39);
nand U910 (N_910,In_1682,N_300);
nand U911 (N_911,In_1959,In_308);
nor U912 (N_912,In_1881,In_1852);
xor U913 (N_913,In_1393,In_83);
nor U914 (N_914,In_1075,In_1864);
xor U915 (N_915,N_463,N_399);
nand U916 (N_916,N_260,In_1128);
nand U917 (N_917,N_437,N_474);
nor U918 (N_918,In_899,In_1108);
and U919 (N_919,N_114,N_419);
and U920 (N_920,In_7,In_649);
or U921 (N_921,In_1426,N_141);
xor U922 (N_922,In_1130,N_106);
or U923 (N_923,In_1615,N_262);
nor U924 (N_924,In_1323,In_1700);
or U925 (N_925,In_841,N_491);
nor U926 (N_926,N_154,In_526);
nand U927 (N_927,In_1661,In_866);
or U928 (N_928,In_522,N_44);
or U929 (N_929,In_1694,In_1854);
nor U930 (N_930,In_924,N_456);
and U931 (N_931,In_1249,In_375);
or U932 (N_932,N_311,In_1693);
nand U933 (N_933,In_261,N_22);
and U934 (N_934,N_332,N_326);
nand U935 (N_935,In_595,N_18);
nand U936 (N_936,N_404,N_165);
or U937 (N_937,In_411,In_1541);
nand U938 (N_938,N_481,N_142);
and U939 (N_939,N_111,N_396);
nand U940 (N_940,In_1928,In_1813);
nor U941 (N_941,In_229,In_815);
nand U942 (N_942,N_318,N_498);
nand U943 (N_943,In_1202,N_472);
nor U944 (N_944,N_151,In_15);
or U945 (N_945,N_398,In_690);
xnor U946 (N_946,N_405,In_1447);
or U947 (N_947,N_371,In_304);
or U948 (N_948,In_128,In_1332);
nor U949 (N_949,In_767,N_418);
or U950 (N_950,In_1610,In_528);
nand U951 (N_951,In_1304,N_423);
nor U952 (N_952,In_1064,N_305);
or U953 (N_953,In_1605,In_58);
nor U954 (N_954,In_999,N_364);
nor U955 (N_955,In_1658,In_1871);
nand U956 (N_956,In_997,In_839);
and U957 (N_957,N_230,N_308);
nor U958 (N_958,N_239,N_161);
nand U959 (N_959,In_807,In_1724);
nand U960 (N_960,In_507,In_1413);
nand U961 (N_961,In_1940,In_146);
nand U962 (N_962,N_231,In_1421);
nand U963 (N_963,In_669,In_1783);
nand U964 (N_964,N_94,N_385);
xnor U965 (N_965,In_687,In_1535);
nand U966 (N_966,In_1416,In_1958);
and U967 (N_967,N_281,In_549);
xnor U968 (N_968,In_1011,In_1214);
nand U969 (N_969,In_1187,N_5);
nor U970 (N_970,N_133,N_61);
nand U971 (N_971,In_1858,In_809);
and U972 (N_972,N_102,N_192);
xnor U973 (N_973,In_171,In_1341);
nor U974 (N_974,In_977,In_63);
nor U975 (N_975,In_717,In_1838);
or U976 (N_976,In_1316,In_290);
and U977 (N_977,In_1692,N_256);
and U978 (N_978,N_394,N_427);
nand U979 (N_979,N_434,N_234);
or U980 (N_980,N_143,In_1106);
nor U981 (N_981,In_1325,In_233);
nor U982 (N_982,N_445,In_1734);
or U983 (N_983,N_112,N_28);
or U984 (N_984,In_505,N_76);
nor U985 (N_985,N_15,In_318);
or U986 (N_986,N_238,N_36);
and U987 (N_987,In_1924,In_904);
or U988 (N_988,In_504,In_1906);
nand U989 (N_989,In_1901,In_1352);
and U990 (N_990,In_1236,In_1676);
nor U991 (N_991,N_149,In_124);
nand U992 (N_992,In_72,In_1476);
or U993 (N_993,In_1378,In_101);
nand U994 (N_994,In_435,In_438);
or U995 (N_995,In_1354,In_311);
xor U996 (N_996,In_1278,In_144);
nand U997 (N_997,N_392,In_1502);
or U998 (N_998,In_1399,N_408);
xnor U999 (N_999,N_69,In_1776);
xnor U1000 (N_1000,In_1949,N_930);
xor U1001 (N_1001,N_818,In_1005);
nand U1002 (N_1002,N_699,In_1243);
xnor U1003 (N_1003,N_737,In_1623);
nor U1004 (N_1004,N_623,N_726);
xnor U1005 (N_1005,N_730,N_49);
xor U1006 (N_1006,N_746,N_783);
nand U1007 (N_1007,N_579,In_581);
xnor U1008 (N_1008,In_1788,N_802);
or U1009 (N_1009,N_945,N_701);
or U1010 (N_1010,N_194,In_476);
nand U1011 (N_1011,In_381,N_552);
or U1012 (N_1012,N_667,N_770);
nand U1013 (N_1013,N_235,In_1137);
nand U1014 (N_1014,In_1995,N_599);
and U1015 (N_1015,N_984,N_857);
nand U1016 (N_1016,N_565,In_8);
and U1017 (N_1017,N_819,In_1484);
or U1018 (N_1018,In_1082,In_14);
nand U1019 (N_1019,In_833,In_1925);
and U1020 (N_1020,N_516,In_1153);
and U1021 (N_1021,N_83,In_968);
nor U1022 (N_1022,N_302,N_331);
and U1023 (N_1023,In_1300,In_1103);
or U1024 (N_1024,N_860,N_710);
nand U1025 (N_1025,In_1574,In_372);
xnor U1026 (N_1026,N_158,N_784);
xor U1027 (N_1027,In_1754,In_1379);
xnor U1028 (N_1028,N_674,In_515);
xnor U1029 (N_1029,In_1878,N_573);
nand U1030 (N_1030,N_859,N_610);
xnor U1031 (N_1031,N_138,N_155);
xnor U1032 (N_1032,N_723,N_30);
and U1033 (N_1033,In_574,N_337);
nor U1034 (N_1034,In_923,N_761);
nand U1035 (N_1035,N_827,In_1372);
xor U1036 (N_1036,N_696,In_1992);
nand U1037 (N_1037,N_722,N_241);
xnor U1038 (N_1038,N_922,N_45);
nand U1039 (N_1039,In_1408,In_1190);
xnor U1040 (N_1040,In_1267,N_872);
nand U1041 (N_1041,N_324,N_742);
or U1042 (N_1042,In_568,N_264);
nand U1043 (N_1043,N_540,In_1991);
xnor U1044 (N_1044,N_828,N_898);
xnor U1045 (N_1045,In_328,In_1247);
nand U1046 (N_1046,In_962,N_496);
and U1047 (N_1047,In_1887,N_936);
and U1048 (N_1048,N_581,N_933);
or U1049 (N_1049,In_889,N_914);
nand U1050 (N_1050,N_250,N_593);
and U1051 (N_1051,N_808,N_541);
or U1052 (N_1052,N_85,In_645);
and U1053 (N_1053,N_609,N_447);
nand U1054 (N_1054,In_1392,In_1559);
xnor U1055 (N_1055,N_992,In_571);
nor U1056 (N_1056,In_1034,In_778);
or U1057 (N_1057,N_35,In_475);
xnor U1058 (N_1058,In_65,N_323);
or U1059 (N_1059,N_969,N_739);
and U1060 (N_1060,N_589,N_334);
or U1061 (N_1061,N_925,N_571);
and U1062 (N_1062,In_1359,N_613);
xnor U1063 (N_1063,N_986,N_807);
xor U1064 (N_1064,N_638,N_856);
nor U1065 (N_1065,N_797,N_961);
nor U1066 (N_1066,N_578,N_775);
or U1067 (N_1067,N_970,In_929);
xnor U1068 (N_1068,N_662,In_1716);
nand U1069 (N_1069,N_139,N_277);
and U1070 (N_1070,N_604,N_353);
nand U1071 (N_1071,In_105,In_558);
and U1072 (N_1072,In_1690,In_325);
xnor U1073 (N_1073,N_630,N_206);
xor U1074 (N_1074,N_904,N_911);
or U1075 (N_1075,N_191,N_833);
nor U1076 (N_1076,In_382,N_873);
nor U1077 (N_1077,N_547,N_316);
and U1078 (N_1078,N_944,N_130);
or U1079 (N_1079,N_608,N_795);
nor U1080 (N_1080,N_724,N_91);
or U1081 (N_1081,N_617,N_233);
xnor U1082 (N_1082,In_781,N_771);
and U1083 (N_1083,N_197,N_772);
or U1084 (N_1084,In_1616,N_920);
xnor U1085 (N_1085,N_641,N_672);
and U1086 (N_1086,In_906,N_490);
or U1087 (N_1087,N_985,N_531);
and U1088 (N_1088,In_725,N_558);
nand U1089 (N_1089,In_890,N_964);
nor U1090 (N_1090,N_9,In_711);
xor U1091 (N_1091,In_41,N_952);
and U1092 (N_1092,N_891,N_957);
or U1093 (N_1093,In_790,N_800);
and U1094 (N_1094,In_106,N_962);
xnor U1095 (N_1095,N_633,N_523);
or U1096 (N_1096,N_816,N_707);
nand U1097 (N_1097,N_46,In_1006);
nand U1098 (N_1098,In_1113,N_963);
xor U1099 (N_1099,In_1431,N_216);
nor U1100 (N_1100,In_624,N_432);
and U1101 (N_1101,N_530,N_452);
nand U1102 (N_1102,N_56,In_1611);
xnor U1103 (N_1103,In_1726,N_907);
and U1104 (N_1104,N_878,N_32);
xnor U1105 (N_1105,N_982,N_661);
or U1106 (N_1106,In_1093,N_152);
xor U1107 (N_1107,N_673,In_1219);
nor U1108 (N_1108,N_572,In_1256);
xor U1109 (N_1109,N_947,In_1081);
or U1110 (N_1110,N_556,N_503);
xor U1111 (N_1111,In_544,N_923);
nand U1112 (N_1112,In_1324,N_98);
or U1113 (N_1113,N_226,In_1533);
xor U1114 (N_1114,N_207,N_595);
or U1115 (N_1115,In_903,N_967);
or U1116 (N_1116,N_528,In_1453);
or U1117 (N_1117,N_518,N_714);
and U1118 (N_1118,N_537,N_847);
and U1119 (N_1119,N_792,N_615);
nor U1120 (N_1120,In_749,N_612);
xor U1121 (N_1121,N_852,N_942);
or U1122 (N_1122,N_690,N_137);
nor U1123 (N_1123,In_1384,In_1708);
nand U1124 (N_1124,N_546,N_321);
xnor U1125 (N_1125,In_1719,N_649);
or U1126 (N_1126,In_536,In_1824);
or U1127 (N_1127,In_834,N_645);
xnor U1128 (N_1128,In_1150,In_1759);
nand U1129 (N_1129,N_763,N_618);
or U1130 (N_1130,N_886,In_1543);
nand U1131 (N_1131,N_168,In_956);
nand U1132 (N_1132,N_596,N_900);
nand U1133 (N_1133,N_948,In_1963);
or U1134 (N_1134,N_505,In_110);
or U1135 (N_1135,N_457,N_670);
and U1136 (N_1136,N_527,N_644);
nor U1137 (N_1137,N_561,N_725);
and U1138 (N_1138,N_586,In_427);
nor U1139 (N_1139,N_939,N_522);
xor U1140 (N_1140,N_539,N_890);
nand U1141 (N_1141,N_950,N_380);
and U1142 (N_1142,N_736,In_845);
nand U1143 (N_1143,In_1969,N_510);
nand U1144 (N_1144,N_888,In_1026);
nand U1145 (N_1145,N_787,N_835);
or U1146 (N_1146,N_682,N_834);
nor U1147 (N_1147,N_862,N_866);
or U1148 (N_1148,In_1481,N_960);
and U1149 (N_1149,In_729,In_907);
nor U1150 (N_1150,In_592,N_753);
xnor U1151 (N_1151,N_449,In_1606);
nor U1152 (N_1152,N_803,N_213);
or U1153 (N_1153,N_829,N_951);
or U1154 (N_1154,In_117,In_1347);
or U1155 (N_1155,N_910,N_16);
nor U1156 (N_1156,In_759,N_467);
or U1157 (N_1157,N_90,In_368);
xor U1158 (N_1158,N_533,N_622);
xor U1159 (N_1159,N_648,In_202);
nand U1160 (N_1160,In_1454,N_335);
nor U1161 (N_1161,In_1613,N_868);
nor U1162 (N_1162,N_431,N_902);
nand U1163 (N_1163,N_758,N_977);
xor U1164 (N_1164,In_1158,N_995);
and U1165 (N_1165,N_273,N_897);
or U1166 (N_1166,N_576,In_1205);
or U1167 (N_1167,N_210,In_532);
nor U1168 (N_1168,N_224,N_253);
or U1169 (N_1169,In_1182,N_875);
or U1170 (N_1170,In_1345,In_1470);
xnor U1171 (N_1171,N_881,In_80);
or U1172 (N_1172,N_177,In_518);
and U1173 (N_1173,N_639,N_750);
nand U1174 (N_1174,N_110,N_70);
or U1175 (N_1175,N_894,In_648);
nand U1176 (N_1176,N_937,In_1781);
or U1177 (N_1177,N_903,In_189);
or U1178 (N_1178,N_257,N_924);
and U1179 (N_1179,N_319,N_480);
nor U1180 (N_1180,N_636,In_222);
nand U1181 (N_1181,N_627,In_612);
nor U1182 (N_1182,N_913,In_1525);
and U1183 (N_1183,N_883,In_1830);
nor U1184 (N_1184,N_42,N_892);
and U1185 (N_1185,In_506,N_631);
nor U1186 (N_1186,N_870,N_837);
nand U1187 (N_1187,N_548,N_584);
nand U1188 (N_1188,N_482,N_974);
or U1189 (N_1189,N_735,N_805);
xor U1190 (N_1190,N_425,N_926);
nor U1191 (N_1191,N_242,In_1248);
nand U1192 (N_1192,N_717,N_801);
xnor U1193 (N_1193,N_777,In_639);
nand U1194 (N_1194,N_603,In_870);
nor U1195 (N_1195,N_685,N_402);
nand U1196 (N_1196,N_748,N_520);
and U1197 (N_1197,N_778,In_1806);
xnor U1198 (N_1198,N_526,In_1550);
nand U1199 (N_1199,N_759,In_35);
or U1200 (N_1200,N_958,In_886);
xnor U1201 (N_1201,In_1609,N_621);
nor U1202 (N_1202,In_550,In_643);
xor U1203 (N_1203,N_731,N_935);
xnor U1204 (N_1204,N_851,In_1772);
nand U1205 (N_1205,N_577,N_743);
nor U1206 (N_1206,In_321,N_677);
xnor U1207 (N_1207,In_1036,N_511);
xor U1208 (N_1208,N_956,In_1675);
nand U1209 (N_1209,N_550,N_884);
xnor U1210 (N_1210,N_104,In_1486);
nor U1211 (N_1211,In_1747,N_477);
nand U1212 (N_1212,N_79,N_651);
and U1213 (N_1213,In_1953,N_506);
nand U1214 (N_1214,In_830,N_738);
xnor U1215 (N_1215,In_460,N_865);
xor U1216 (N_1216,N_602,N_695);
xor U1217 (N_1217,In_1523,In_1231);
or U1218 (N_1218,In_56,In_1572);
nor U1219 (N_1219,N_507,In_1317);
or U1220 (N_1220,N_128,In_523);
nor U1221 (N_1221,N_990,N_700);
xnor U1222 (N_1222,N_713,N_780);
nor U1223 (N_1223,N_683,N_632);
nor U1224 (N_1224,N_694,N_706);
and U1225 (N_1225,N_812,N_766);
and U1226 (N_1226,In_543,N_75);
or U1227 (N_1227,N_607,N_313);
xor U1228 (N_1228,In_1835,N_363);
xnor U1229 (N_1229,In_224,N_728);
and U1230 (N_1230,N_751,In_459);
nand U1231 (N_1231,N_987,In_1649);
xnor U1232 (N_1232,N_679,N_980);
nor U1233 (N_1233,N_867,N_656);
nor U1234 (N_1234,N_989,N_796);
nand U1235 (N_1235,In_353,N_20);
and U1236 (N_1236,N_655,N_830);
nor U1237 (N_1237,In_524,N_665);
or U1238 (N_1238,In_181,In_1903);
xnor U1239 (N_1239,In_1273,In_1291);
nor U1240 (N_1240,In_782,N_916);
and U1241 (N_1241,N_978,N_814);
or U1242 (N_1242,N_949,In_1321);
nor U1243 (N_1243,In_204,N_680);
and U1244 (N_1244,N_806,In_590);
nand U1245 (N_1245,N_844,N_899);
xnor U1246 (N_1246,In_1697,In_156);
and U1247 (N_1247,N_825,N_361);
nand U1248 (N_1248,N_813,N_773);
nor U1249 (N_1249,N_515,In_316);
xor U1250 (N_1250,In_1504,In_1859);
and U1251 (N_1251,In_69,N_749);
nor U1252 (N_1252,N_81,N_646);
nand U1253 (N_1253,In_606,N_588);
nor U1254 (N_1254,In_1730,N_747);
or U1255 (N_1255,N_678,N_614);
nand U1256 (N_1256,N_858,N_534);
and U1257 (N_1257,N_356,N_943);
or U1258 (N_1258,N_619,In_698);
xnor U1259 (N_1259,N_705,In_123);
nor U1260 (N_1260,N_637,In_17);
nor U1261 (N_1261,N_940,N_727);
nor U1262 (N_1262,In_392,N_721);
and U1263 (N_1263,N_583,N_436);
and U1264 (N_1264,N_893,N_601);
and U1265 (N_1265,In_391,N_843);
and U1266 (N_1266,In_704,N_211);
or U1267 (N_1267,N_529,N_663);
xnor U1268 (N_1268,N_379,N_712);
nor U1269 (N_1269,In_989,N_981);
nand U1270 (N_1270,In_1377,In_1404);
xor U1271 (N_1271,N_921,N_459);
or U1272 (N_1272,N_524,In_791);
or U1273 (N_1273,N_513,N_536);
nand U1274 (N_1274,N_740,N_659);
and U1275 (N_1275,In_256,In_1367);
nor U1276 (N_1276,In_563,In_1206);
or U1277 (N_1277,N_817,In_1756);
or U1278 (N_1278,In_240,N_732);
xor U1279 (N_1279,N_776,N_669);
nor U1280 (N_1280,N_876,N_555);
nor U1281 (N_1281,N_823,N_653);
nor U1282 (N_1282,N_369,In_974);
xnor U1283 (N_1283,N_885,In_1195);
and U1284 (N_1284,In_1080,In_1466);
nand U1285 (N_1285,N_764,N_769);
nand U1286 (N_1286,In_942,In_1003);
or U1287 (N_1287,N_850,In_289);
nand U1288 (N_1288,In_1505,N_959);
nand U1289 (N_1289,N_846,N_525);
xor U1290 (N_1290,In_388,In_1204);
or U1291 (N_1291,N_635,N_934);
nor U1292 (N_1292,N_809,N_14);
or U1293 (N_1293,In_1913,N_832);
or U1294 (N_1294,In_77,In_412);
xnor U1295 (N_1295,N_786,In_1276);
or U1296 (N_1296,N_983,N_909);
and U1297 (N_1297,N_824,N_676);
nor U1298 (N_1298,In_223,In_1844);
or U1299 (N_1299,In_1047,N_968);
nand U1300 (N_1300,In_1576,N_996);
nor U1301 (N_1301,N_562,N_202);
or U1302 (N_1302,N_932,In_1079);
nor U1303 (N_1303,N_625,N_927);
and U1304 (N_1304,N_120,N_733);
xor U1305 (N_1305,In_295,N_620);
or U1306 (N_1306,N_785,In_414);
and U1307 (N_1307,N_658,N_598);
or U1308 (N_1308,N_946,N_993);
xor U1309 (N_1309,In_73,In_939);
nor U1310 (N_1310,N_779,N_647);
or U1311 (N_1311,In_451,In_338);
nor U1312 (N_1312,N_841,In_462);
and U1313 (N_1313,In_613,N_587);
xor U1314 (N_1314,In_1985,N_681);
or U1315 (N_1315,N_86,N_869);
or U1316 (N_1316,N_8,In_1041);
and U1317 (N_1317,In_448,In_542);
xor U1318 (N_1318,N_688,N_767);
and U1319 (N_1319,In_689,N_147);
nor U1320 (N_1320,In_1430,N_479);
nor U1321 (N_1321,In_1432,N_811);
or U1322 (N_1322,N_789,In_508);
or U1323 (N_1323,N_991,N_585);
and U1324 (N_1324,N_135,N_693);
and U1325 (N_1325,N_912,N_77);
and U1326 (N_1326,In_1013,N_101);
xor U1327 (N_1327,In_1654,N_788);
or U1328 (N_1328,N_687,N_854);
nor U1329 (N_1329,In_264,In_868);
nor U1330 (N_1330,In_1760,N_838);
and U1331 (N_1331,In_1445,In_355);
xnor U1332 (N_1332,N_831,In_484);
nor U1333 (N_1333,In_1932,N_781);
or U1334 (N_1334,In_153,In_1340);
or U1335 (N_1335,In_1914,N_575);
and U1336 (N_1336,In_1670,In_1738);
xor U1337 (N_1337,In_39,N_27);
nor U1338 (N_1338,In_1732,N_709);
xor U1339 (N_1339,N_861,N_535);
nand U1340 (N_1340,In_1839,N_666);
nor U1341 (N_1341,In_1112,N_590);
nand U1342 (N_1342,In_1968,N_350);
xor U1343 (N_1343,In_1586,N_810);
nor U1344 (N_1344,In_158,N_791);
nand U1345 (N_1345,N_566,N_417);
nand U1346 (N_1346,N_338,N_554);
and U1347 (N_1347,In_1938,N_840);
and U1348 (N_1348,N_569,N_450);
xor U1349 (N_1349,N_58,N_839);
nor U1350 (N_1350,In_1873,In_258);
nor U1351 (N_1351,In_140,N_611);
and U1352 (N_1352,N_19,In_1297);
or U1353 (N_1353,N_689,N_6);
nor U1354 (N_1354,In_1765,In_1020);
and U1355 (N_1355,N_686,N_594);
or U1356 (N_1356,N_570,In_1183);
and U1357 (N_1357,In_1809,N_822);
nor U1358 (N_1358,N_938,N_882);
xnor U1359 (N_1359,N_820,N_826);
and U1360 (N_1360,In_1798,In_1022);
and U1361 (N_1361,N_275,N_794);
nand U1362 (N_1362,In_567,In_1639);
or U1363 (N_1363,N_557,In_1092);
or U1364 (N_1364,N_799,In_276);
nor U1365 (N_1365,In_1910,In_731);
nand U1366 (N_1366,N_845,In_1472);
nor U1367 (N_1367,N_928,N_551);
and U1368 (N_1368,N_634,In_1766);
or U1369 (N_1369,In_681,N_815);
and U1370 (N_1370,In_218,N_698);
nor U1371 (N_1371,In_1309,In_1272);
nor U1372 (N_1372,In_1869,N_716);
or U1373 (N_1373,N_65,N_979);
or U1374 (N_1374,N_650,N_509);
nand U1375 (N_1375,N_756,N_501);
nor U1376 (N_1376,N_328,N_760);
nor U1377 (N_1377,N_512,N_684);
nor U1378 (N_1378,N_874,N_629);
nand U1379 (N_1379,N_173,N_668);
and U1380 (N_1380,N_768,N_798);
or U1381 (N_1381,N_877,N_97);
nor U1382 (N_1382,In_800,N_853);
nand U1383 (N_1383,N_153,N_580);
and U1384 (N_1384,N_263,In_60);
or U1385 (N_1385,N_183,N_582);
xor U1386 (N_1386,In_1911,N_744);
and U1387 (N_1387,In_860,In_1952);
or U1388 (N_1388,N_115,N_745);
xnor U1389 (N_1389,N_757,In_1173);
xnor U1390 (N_1390,In_1909,N_538);
nand U1391 (N_1391,N_351,N_12);
or U1392 (N_1392,N_880,In_901);
xor U1393 (N_1393,In_1044,N_95);
and U1394 (N_1394,In_887,N_368);
and U1395 (N_1395,N_734,In_969);
nand U1396 (N_1396,N_973,In_1232);
nand U1397 (N_1397,In_638,N_521);
xor U1398 (N_1398,N_29,In_1362);
nand U1399 (N_1399,N_821,In_4);
and U1400 (N_1400,N_864,N_345);
and U1401 (N_1401,N_403,N_918);
and U1402 (N_1402,N_718,In_1373);
and U1403 (N_1403,N_972,N_999);
or U1404 (N_1404,N_976,In_1628);
xnor U1405 (N_1405,In_494,In_934);
or U1406 (N_1406,N_592,N_248);
nor U1407 (N_1407,N_691,In_947);
xor U1408 (N_1408,In_1172,N_460);
and U1409 (N_1409,N_466,N_863);
and U1410 (N_1410,N_703,In_819);
and U1411 (N_1411,N_966,In_493);
or U1412 (N_1412,In_1702,N_504);
xnor U1413 (N_1413,N_896,N_628);
xnor U1414 (N_1414,N_391,N_704);
or U1415 (N_1415,In_1774,In_293);
nand U1416 (N_1416,In_1131,N_473);
nor U1417 (N_1417,N_988,In_1863);
or U1418 (N_1418,N_25,N_545);
or U1419 (N_1419,N_532,N_297);
nor U1420 (N_1420,In_43,N_941);
nor U1421 (N_1421,In_1461,N_500);
nor U1422 (N_1422,N_793,N_953);
xnor U1423 (N_1423,N_624,N_919);
nor U1424 (N_1424,In_370,In_1689);
nand U1425 (N_1425,N_560,N_755);
nand U1426 (N_1426,N_836,N_697);
nand U1427 (N_1427,N_428,N_975);
or U1428 (N_1428,In_656,N_568);
nor U1429 (N_1429,N_606,N_998);
nor U1430 (N_1430,N_354,N_198);
or U1431 (N_1431,N_508,N_502);
nor U1432 (N_1432,N_848,In_1315);
nand U1433 (N_1433,N_729,N_188);
or U1434 (N_1434,In_1547,In_710);
and U1435 (N_1435,In_762,N_664);
nand U1436 (N_1436,N_478,N_514);
or U1437 (N_1437,N_543,In_1905);
or U1438 (N_1438,In_1796,N_544);
xnor U1439 (N_1439,N_675,In_434);
and U1440 (N_1440,In_1775,In_1314);
or U1441 (N_1441,In_911,In_1270);
nor U1442 (N_1442,N_917,In_92);
nand U1443 (N_1443,In_1646,N_915);
and U1444 (N_1444,N_597,N_643);
nand U1445 (N_1445,N_549,N_574);
nand U1446 (N_1446,In_159,N_517);
xnor U1447 (N_1447,In_1829,N_563);
and U1448 (N_1448,In_1042,In_47);
nand U1449 (N_1449,In_1401,N_849);
xor U1450 (N_1450,In_182,N_567);
nor U1451 (N_1451,N_50,N_140);
nor U1452 (N_1452,In_403,N_251);
xor U1453 (N_1453,N_542,In_715);
xnor U1454 (N_1454,In_630,N_906);
xnor U1455 (N_1455,N_741,N_270);
nor U1456 (N_1456,In_213,In_1360);
and U1457 (N_1457,In_1832,In_1100);
nor U1458 (N_1458,N_626,N_782);
nor U1459 (N_1459,N_720,In_640);
xnor U1460 (N_1460,N_715,N_889);
or U1461 (N_1461,N_954,N_895);
xnor U1462 (N_1462,N_997,N_711);
and U1463 (N_1463,In_1067,N_72);
or U1464 (N_1464,N_559,In_1695);
or U1465 (N_1465,N_476,In_31);
and U1466 (N_1466,N_184,N_931);
and U1467 (N_1467,In_626,N_519);
nor U1468 (N_1468,N_660,N_905);
nand U1469 (N_1469,N_994,N_719);
nand U1470 (N_1470,In_561,N_855);
or U1471 (N_1471,N_600,N_804);
xor U1472 (N_1472,In_331,N_774);
nand U1473 (N_1473,N_616,In_1091);
and U1474 (N_1474,In_1733,In_810);
and U1475 (N_1475,N_564,N_908);
nand U1476 (N_1476,In_1821,In_1614);
nor U1477 (N_1477,In_1895,N_376);
or U1478 (N_1478,N_692,In_1290);
and U1479 (N_1479,In_112,N_122);
or U1480 (N_1480,N_654,N_605);
nor U1481 (N_1481,N_123,N_708);
and U1482 (N_1482,N_214,In_556);
xnor U1483 (N_1483,N_965,N_929);
and U1484 (N_1484,N_842,N_887);
nor U1485 (N_1485,In_490,N_879);
or U1486 (N_1486,N_871,N_901);
and U1487 (N_1487,In_277,N_485);
or U1488 (N_1488,In_1115,N_442);
xor U1489 (N_1489,N_657,N_702);
xnor U1490 (N_1490,N_754,N_671);
xnor U1491 (N_1491,N_553,N_790);
or U1492 (N_1492,N_765,N_591);
or U1493 (N_1493,In_1188,N_642);
nor U1494 (N_1494,In_1418,N_237);
or U1495 (N_1495,N_762,N_752);
xnor U1496 (N_1496,N_125,N_175);
and U1497 (N_1497,N_971,N_955);
xnor U1498 (N_1498,N_640,N_82);
nor U1499 (N_1499,N_652,N_349);
nand U1500 (N_1500,N_1402,N_1417);
nand U1501 (N_1501,N_1201,N_1346);
nor U1502 (N_1502,N_1207,N_1266);
nand U1503 (N_1503,N_1015,N_1149);
or U1504 (N_1504,N_1358,N_1058);
or U1505 (N_1505,N_1364,N_1180);
and U1506 (N_1506,N_1320,N_1272);
or U1507 (N_1507,N_1369,N_1191);
and U1508 (N_1508,N_1345,N_1000);
and U1509 (N_1509,N_1436,N_1195);
and U1510 (N_1510,N_1498,N_1390);
nand U1511 (N_1511,N_1188,N_1227);
and U1512 (N_1512,N_1018,N_1024);
xnor U1513 (N_1513,N_1156,N_1353);
xnor U1514 (N_1514,N_1397,N_1106);
or U1515 (N_1515,N_1029,N_1268);
and U1516 (N_1516,N_1438,N_1141);
xor U1517 (N_1517,N_1143,N_1261);
and U1518 (N_1518,N_1181,N_1072);
nand U1519 (N_1519,N_1486,N_1271);
and U1520 (N_1520,N_1456,N_1043);
xnor U1521 (N_1521,N_1416,N_1133);
nand U1522 (N_1522,N_1477,N_1145);
xor U1523 (N_1523,N_1273,N_1357);
xor U1524 (N_1524,N_1009,N_1165);
nor U1525 (N_1525,N_1077,N_1304);
nor U1526 (N_1526,N_1326,N_1122);
xnor U1527 (N_1527,N_1105,N_1011);
or U1528 (N_1528,N_1166,N_1295);
or U1529 (N_1529,N_1062,N_1437);
xor U1530 (N_1530,N_1136,N_1359);
and U1531 (N_1531,N_1123,N_1240);
nand U1532 (N_1532,N_1292,N_1441);
or U1533 (N_1533,N_1217,N_1399);
nor U1534 (N_1534,N_1160,N_1265);
and U1535 (N_1535,N_1178,N_1184);
and U1536 (N_1536,N_1244,N_1342);
nor U1537 (N_1537,N_1098,N_1007);
nand U1538 (N_1538,N_1041,N_1443);
nor U1539 (N_1539,N_1352,N_1091);
xor U1540 (N_1540,N_1175,N_1373);
nand U1541 (N_1541,N_1279,N_1107);
nand U1542 (N_1542,N_1259,N_1013);
nand U1543 (N_1543,N_1348,N_1488);
and U1544 (N_1544,N_1117,N_1404);
or U1545 (N_1545,N_1350,N_1118);
or U1546 (N_1546,N_1237,N_1391);
nand U1547 (N_1547,N_1252,N_1487);
and U1548 (N_1548,N_1253,N_1276);
xor U1549 (N_1549,N_1316,N_1021);
and U1550 (N_1550,N_1419,N_1289);
nor U1551 (N_1551,N_1204,N_1473);
and U1552 (N_1552,N_1343,N_1274);
nand U1553 (N_1553,N_1220,N_1039);
xnor U1554 (N_1554,N_1186,N_1340);
xor U1555 (N_1555,N_1079,N_1383);
xor U1556 (N_1556,N_1001,N_1066);
nand U1557 (N_1557,N_1338,N_1494);
xor U1558 (N_1558,N_1499,N_1169);
nand U1559 (N_1559,N_1046,N_1476);
nor U1560 (N_1560,N_1291,N_1398);
xnor U1561 (N_1561,N_1028,N_1228);
xnor U1562 (N_1562,N_1331,N_1019);
nor U1563 (N_1563,N_1005,N_1194);
nand U1564 (N_1564,N_1395,N_1442);
or U1565 (N_1565,N_1170,N_1251);
nor U1566 (N_1566,N_1100,N_1162);
nor U1567 (N_1567,N_1367,N_1474);
or U1568 (N_1568,N_1382,N_1255);
or U1569 (N_1569,N_1017,N_1471);
or U1570 (N_1570,N_1238,N_1030);
xor U1571 (N_1571,N_1366,N_1299);
xnor U1572 (N_1572,N_1294,N_1014);
or U1573 (N_1573,N_1362,N_1139);
and U1574 (N_1574,N_1192,N_1457);
xor U1575 (N_1575,N_1374,N_1298);
nor U1576 (N_1576,N_1097,N_1137);
nor U1577 (N_1577,N_1464,N_1452);
xor U1578 (N_1578,N_1260,N_1067);
xor U1579 (N_1579,N_1293,N_1214);
nand U1580 (N_1580,N_1129,N_1386);
nand U1581 (N_1581,N_1300,N_1212);
and U1582 (N_1582,N_1490,N_1344);
nor U1583 (N_1583,N_1037,N_1224);
or U1584 (N_1584,N_1094,N_1275);
xnor U1585 (N_1585,N_1092,N_1082);
xnor U1586 (N_1586,N_1425,N_1110);
nand U1587 (N_1587,N_1093,N_1329);
or U1588 (N_1588,N_1151,N_1108);
or U1589 (N_1589,N_1065,N_1258);
and U1590 (N_1590,N_1182,N_1307);
nand U1591 (N_1591,N_1284,N_1447);
or U1592 (N_1592,N_1347,N_1269);
nand U1593 (N_1593,N_1341,N_1115);
nand U1594 (N_1594,N_1031,N_1462);
or U1595 (N_1595,N_1140,N_1006);
nor U1596 (N_1596,N_1485,N_1433);
or U1597 (N_1597,N_1286,N_1424);
nor U1598 (N_1598,N_1008,N_1384);
nor U1599 (N_1599,N_1283,N_1247);
and U1600 (N_1600,N_1174,N_1408);
xnor U1601 (N_1601,N_1423,N_1095);
nor U1602 (N_1602,N_1389,N_1309);
nand U1603 (N_1603,N_1057,N_1431);
xnor U1604 (N_1604,N_1125,N_1157);
nor U1605 (N_1605,N_1270,N_1446);
nand U1606 (N_1606,N_1434,N_1463);
xnor U1607 (N_1607,N_1033,N_1250);
nor U1608 (N_1608,N_1484,N_1163);
or U1609 (N_1609,N_1096,N_1303);
nand U1610 (N_1610,N_1004,N_1168);
xor U1611 (N_1611,N_1306,N_1313);
or U1612 (N_1612,N_1056,N_1475);
nand U1613 (N_1613,N_1172,N_1491);
xnor U1614 (N_1614,N_1103,N_1109);
nand U1615 (N_1615,N_1365,N_1439);
and U1616 (N_1616,N_1047,N_1392);
nor U1617 (N_1617,N_1090,N_1128);
and U1618 (N_1618,N_1049,N_1076);
and U1619 (N_1619,N_1314,N_1328);
or U1620 (N_1620,N_1405,N_1327);
nand U1621 (N_1621,N_1460,N_1155);
and U1622 (N_1622,N_1003,N_1311);
and U1623 (N_1623,N_1010,N_1246);
or U1624 (N_1624,N_1078,N_1415);
nor U1625 (N_1625,N_1497,N_1002);
xor U1626 (N_1626,N_1267,N_1130);
nor U1627 (N_1627,N_1429,N_1216);
nand U1628 (N_1628,N_1189,N_1027);
nor U1629 (N_1629,N_1124,N_1150);
xor U1630 (N_1630,N_1281,N_1241);
or U1631 (N_1631,N_1278,N_1127);
xnor U1632 (N_1632,N_1210,N_1202);
and U1633 (N_1633,N_1114,N_1074);
or U1634 (N_1634,N_1104,N_1154);
and U1635 (N_1635,N_1197,N_1226);
and U1636 (N_1636,N_1211,N_1230);
and U1637 (N_1637,N_1467,N_1025);
xnor U1638 (N_1638,N_1396,N_1022);
xor U1639 (N_1639,N_1221,N_1101);
xnor U1640 (N_1640,N_1310,N_1236);
or U1641 (N_1641,N_1451,N_1167);
or U1642 (N_1642,N_1198,N_1054);
or U1643 (N_1643,N_1459,N_1470);
or U1644 (N_1644,N_1371,N_1040);
and U1645 (N_1645,N_1385,N_1083);
nand U1646 (N_1646,N_1445,N_1234);
nor U1647 (N_1647,N_1282,N_1409);
nor U1648 (N_1648,N_1086,N_1052);
nor U1649 (N_1649,N_1361,N_1042);
or U1650 (N_1650,N_1060,N_1356);
and U1651 (N_1651,N_1351,N_1073);
nand U1652 (N_1652,N_1349,N_1063);
nand U1653 (N_1653,N_1323,N_1159);
xor U1654 (N_1654,N_1332,N_1393);
nor U1655 (N_1655,N_1480,N_1089);
or U1656 (N_1656,N_1435,N_1048);
or U1657 (N_1657,N_1355,N_1087);
nor U1658 (N_1658,N_1147,N_1388);
nand U1659 (N_1659,N_1233,N_1161);
xor U1660 (N_1660,N_1449,N_1171);
nand U1661 (N_1661,N_1026,N_1257);
or U1662 (N_1662,N_1229,N_1080);
xor U1663 (N_1663,N_1132,N_1223);
or U1664 (N_1664,N_1177,N_1495);
xor U1665 (N_1665,N_1381,N_1312);
xnor U1666 (N_1666,N_1068,N_1302);
and U1667 (N_1667,N_1187,N_1363);
nor U1668 (N_1668,N_1245,N_1239);
nor U1669 (N_1669,N_1020,N_1318);
or U1670 (N_1670,N_1148,N_1243);
nor U1671 (N_1671,N_1263,N_1315);
xnor U1672 (N_1672,N_1111,N_1413);
nor U1673 (N_1673,N_1297,N_1481);
nor U1674 (N_1674,N_1410,N_1053);
nor U1675 (N_1675,N_1420,N_1036);
nor U1676 (N_1676,N_1045,N_1213);
or U1677 (N_1677,N_1370,N_1375);
or U1678 (N_1678,N_1200,N_1050);
nor U1679 (N_1679,N_1061,N_1102);
nor U1680 (N_1680,N_1085,N_1231);
nor U1681 (N_1681,N_1138,N_1305);
or U1682 (N_1682,N_1038,N_1064);
nor U1683 (N_1683,N_1321,N_1377);
xor U1684 (N_1684,N_1319,N_1450);
and U1685 (N_1685,N_1121,N_1461);
nand U1686 (N_1686,N_1206,N_1354);
xnor U1687 (N_1687,N_1422,N_1120);
or U1688 (N_1688,N_1466,N_1453);
nor U1689 (N_1689,N_1242,N_1492);
nand U1690 (N_1690,N_1472,N_1158);
or U1691 (N_1691,N_1055,N_1478);
nor U1692 (N_1692,N_1360,N_1322);
or U1693 (N_1693,N_1387,N_1209);
or U1694 (N_1694,N_1146,N_1380);
and U1695 (N_1695,N_1482,N_1368);
and U1696 (N_1696,N_1113,N_1222);
xor U1697 (N_1697,N_1135,N_1468);
xor U1698 (N_1698,N_1287,N_1317);
and U1699 (N_1699,N_1185,N_1428);
nor U1700 (N_1700,N_1337,N_1084);
and U1701 (N_1701,N_1333,N_1335);
nand U1702 (N_1702,N_1219,N_1203);
xor U1703 (N_1703,N_1496,N_1248);
nand U1704 (N_1704,N_1112,N_1330);
and U1705 (N_1705,N_1059,N_1406);
and U1706 (N_1706,N_1012,N_1407);
or U1707 (N_1707,N_1465,N_1479);
and U1708 (N_1708,N_1277,N_1264);
nand U1709 (N_1709,N_1193,N_1334);
xnor U1710 (N_1710,N_1215,N_1290);
and U1711 (N_1711,N_1411,N_1099);
nand U1712 (N_1712,N_1430,N_1134);
and U1713 (N_1713,N_1285,N_1131);
xnor U1714 (N_1714,N_1153,N_1454);
nor U1715 (N_1715,N_1262,N_1493);
nor U1716 (N_1716,N_1296,N_1032);
nor U1717 (N_1717,N_1403,N_1249);
nand U1718 (N_1718,N_1235,N_1088);
and U1719 (N_1719,N_1444,N_1034);
nand U1720 (N_1720,N_1075,N_1199);
or U1721 (N_1721,N_1071,N_1288);
nor U1722 (N_1722,N_1218,N_1069);
nand U1723 (N_1723,N_1301,N_1225);
nor U1724 (N_1724,N_1173,N_1081);
and U1725 (N_1725,N_1183,N_1044);
xor U1726 (N_1726,N_1412,N_1394);
nand U1727 (N_1727,N_1376,N_1483);
or U1728 (N_1728,N_1070,N_1256);
nor U1729 (N_1729,N_1280,N_1144);
or U1730 (N_1730,N_1448,N_1116);
nand U1731 (N_1731,N_1336,N_1378);
or U1732 (N_1732,N_1339,N_1489);
nor U1733 (N_1733,N_1372,N_1308);
nor U1734 (N_1734,N_1418,N_1432);
nor U1735 (N_1735,N_1427,N_1440);
or U1736 (N_1736,N_1205,N_1208);
nor U1737 (N_1737,N_1325,N_1179);
and U1738 (N_1738,N_1421,N_1016);
nand U1739 (N_1739,N_1324,N_1379);
and U1740 (N_1740,N_1023,N_1152);
xnor U1741 (N_1741,N_1126,N_1458);
nand U1742 (N_1742,N_1190,N_1455);
xnor U1743 (N_1743,N_1196,N_1119);
nand U1744 (N_1744,N_1426,N_1051);
or U1745 (N_1745,N_1469,N_1176);
xnor U1746 (N_1746,N_1414,N_1142);
xor U1747 (N_1747,N_1400,N_1232);
nor U1748 (N_1748,N_1164,N_1254);
nor U1749 (N_1749,N_1401,N_1035);
and U1750 (N_1750,N_1031,N_1257);
xor U1751 (N_1751,N_1118,N_1412);
nor U1752 (N_1752,N_1477,N_1029);
and U1753 (N_1753,N_1077,N_1386);
nand U1754 (N_1754,N_1074,N_1041);
and U1755 (N_1755,N_1323,N_1115);
or U1756 (N_1756,N_1451,N_1401);
xnor U1757 (N_1757,N_1066,N_1184);
nor U1758 (N_1758,N_1362,N_1103);
nor U1759 (N_1759,N_1054,N_1410);
xnor U1760 (N_1760,N_1276,N_1415);
nand U1761 (N_1761,N_1058,N_1309);
and U1762 (N_1762,N_1376,N_1002);
or U1763 (N_1763,N_1487,N_1297);
and U1764 (N_1764,N_1453,N_1393);
xnor U1765 (N_1765,N_1314,N_1261);
and U1766 (N_1766,N_1049,N_1287);
and U1767 (N_1767,N_1301,N_1366);
and U1768 (N_1768,N_1232,N_1013);
nand U1769 (N_1769,N_1472,N_1270);
and U1770 (N_1770,N_1306,N_1467);
and U1771 (N_1771,N_1297,N_1307);
xor U1772 (N_1772,N_1340,N_1090);
nand U1773 (N_1773,N_1063,N_1069);
or U1774 (N_1774,N_1282,N_1494);
and U1775 (N_1775,N_1171,N_1139);
xor U1776 (N_1776,N_1373,N_1186);
xor U1777 (N_1777,N_1237,N_1042);
nor U1778 (N_1778,N_1315,N_1162);
nand U1779 (N_1779,N_1096,N_1143);
xnor U1780 (N_1780,N_1341,N_1400);
and U1781 (N_1781,N_1125,N_1244);
and U1782 (N_1782,N_1246,N_1151);
or U1783 (N_1783,N_1105,N_1397);
nand U1784 (N_1784,N_1019,N_1310);
and U1785 (N_1785,N_1353,N_1133);
and U1786 (N_1786,N_1118,N_1260);
or U1787 (N_1787,N_1426,N_1215);
nand U1788 (N_1788,N_1066,N_1252);
nor U1789 (N_1789,N_1107,N_1470);
nand U1790 (N_1790,N_1170,N_1016);
xor U1791 (N_1791,N_1261,N_1123);
nor U1792 (N_1792,N_1102,N_1335);
or U1793 (N_1793,N_1128,N_1094);
nor U1794 (N_1794,N_1465,N_1188);
nor U1795 (N_1795,N_1310,N_1165);
nor U1796 (N_1796,N_1162,N_1067);
and U1797 (N_1797,N_1025,N_1212);
nor U1798 (N_1798,N_1026,N_1099);
and U1799 (N_1799,N_1208,N_1100);
nor U1800 (N_1800,N_1045,N_1422);
or U1801 (N_1801,N_1114,N_1069);
xnor U1802 (N_1802,N_1373,N_1131);
nand U1803 (N_1803,N_1410,N_1341);
nand U1804 (N_1804,N_1235,N_1433);
xnor U1805 (N_1805,N_1457,N_1093);
and U1806 (N_1806,N_1258,N_1404);
nand U1807 (N_1807,N_1347,N_1280);
xor U1808 (N_1808,N_1462,N_1434);
xnor U1809 (N_1809,N_1391,N_1499);
and U1810 (N_1810,N_1301,N_1055);
nor U1811 (N_1811,N_1285,N_1494);
xnor U1812 (N_1812,N_1398,N_1200);
or U1813 (N_1813,N_1040,N_1159);
and U1814 (N_1814,N_1187,N_1209);
or U1815 (N_1815,N_1286,N_1194);
and U1816 (N_1816,N_1420,N_1251);
xor U1817 (N_1817,N_1333,N_1325);
or U1818 (N_1818,N_1401,N_1434);
nor U1819 (N_1819,N_1217,N_1471);
nor U1820 (N_1820,N_1135,N_1234);
or U1821 (N_1821,N_1052,N_1178);
or U1822 (N_1822,N_1255,N_1065);
and U1823 (N_1823,N_1280,N_1266);
nand U1824 (N_1824,N_1468,N_1368);
or U1825 (N_1825,N_1219,N_1478);
or U1826 (N_1826,N_1348,N_1260);
xor U1827 (N_1827,N_1462,N_1282);
nand U1828 (N_1828,N_1398,N_1107);
xor U1829 (N_1829,N_1378,N_1476);
and U1830 (N_1830,N_1005,N_1216);
or U1831 (N_1831,N_1001,N_1002);
or U1832 (N_1832,N_1403,N_1113);
nor U1833 (N_1833,N_1478,N_1400);
nor U1834 (N_1834,N_1328,N_1286);
nand U1835 (N_1835,N_1212,N_1224);
or U1836 (N_1836,N_1230,N_1150);
or U1837 (N_1837,N_1243,N_1434);
or U1838 (N_1838,N_1263,N_1296);
nand U1839 (N_1839,N_1338,N_1300);
and U1840 (N_1840,N_1291,N_1223);
xnor U1841 (N_1841,N_1140,N_1354);
and U1842 (N_1842,N_1499,N_1472);
nand U1843 (N_1843,N_1079,N_1334);
or U1844 (N_1844,N_1038,N_1489);
or U1845 (N_1845,N_1419,N_1281);
xnor U1846 (N_1846,N_1490,N_1165);
and U1847 (N_1847,N_1272,N_1335);
nand U1848 (N_1848,N_1227,N_1255);
and U1849 (N_1849,N_1035,N_1141);
nor U1850 (N_1850,N_1054,N_1374);
and U1851 (N_1851,N_1269,N_1451);
xnor U1852 (N_1852,N_1457,N_1039);
xnor U1853 (N_1853,N_1265,N_1068);
or U1854 (N_1854,N_1390,N_1259);
nor U1855 (N_1855,N_1220,N_1138);
nor U1856 (N_1856,N_1174,N_1162);
nor U1857 (N_1857,N_1434,N_1464);
nor U1858 (N_1858,N_1062,N_1069);
nor U1859 (N_1859,N_1060,N_1021);
or U1860 (N_1860,N_1264,N_1340);
xnor U1861 (N_1861,N_1456,N_1204);
and U1862 (N_1862,N_1418,N_1382);
nand U1863 (N_1863,N_1349,N_1366);
or U1864 (N_1864,N_1443,N_1196);
nor U1865 (N_1865,N_1485,N_1070);
and U1866 (N_1866,N_1496,N_1399);
or U1867 (N_1867,N_1396,N_1438);
and U1868 (N_1868,N_1384,N_1028);
nand U1869 (N_1869,N_1073,N_1391);
nor U1870 (N_1870,N_1271,N_1157);
nand U1871 (N_1871,N_1127,N_1266);
xor U1872 (N_1872,N_1146,N_1317);
nand U1873 (N_1873,N_1226,N_1203);
or U1874 (N_1874,N_1078,N_1260);
nand U1875 (N_1875,N_1460,N_1493);
xnor U1876 (N_1876,N_1384,N_1341);
or U1877 (N_1877,N_1056,N_1001);
nand U1878 (N_1878,N_1432,N_1388);
nand U1879 (N_1879,N_1449,N_1185);
nand U1880 (N_1880,N_1087,N_1316);
or U1881 (N_1881,N_1011,N_1376);
nand U1882 (N_1882,N_1008,N_1130);
or U1883 (N_1883,N_1357,N_1183);
xnor U1884 (N_1884,N_1167,N_1175);
xnor U1885 (N_1885,N_1215,N_1253);
or U1886 (N_1886,N_1448,N_1176);
and U1887 (N_1887,N_1167,N_1185);
and U1888 (N_1888,N_1401,N_1333);
nand U1889 (N_1889,N_1358,N_1094);
nor U1890 (N_1890,N_1008,N_1489);
nand U1891 (N_1891,N_1146,N_1178);
nor U1892 (N_1892,N_1302,N_1349);
and U1893 (N_1893,N_1438,N_1246);
nor U1894 (N_1894,N_1488,N_1327);
or U1895 (N_1895,N_1401,N_1429);
and U1896 (N_1896,N_1192,N_1089);
and U1897 (N_1897,N_1388,N_1210);
nand U1898 (N_1898,N_1359,N_1301);
or U1899 (N_1899,N_1125,N_1456);
nor U1900 (N_1900,N_1109,N_1081);
nor U1901 (N_1901,N_1245,N_1177);
nand U1902 (N_1902,N_1030,N_1262);
xnor U1903 (N_1903,N_1371,N_1002);
xnor U1904 (N_1904,N_1131,N_1081);
nand U1905 (N_1905,N_1321,N_1156);
and U1906 (N_1906,N_1325,N_1414);
and U1907 (N_1907,N_1416,N_1149);
nand U1908 (N_1908,N_1472,N_1290);
and U1909 (N_1909,N_1258,N_1485);
or U1910 (N_1910,N_1409,N_1201);
nor U1911 (N_1911,N_1281,N_1295);
xor U1912 (N_1912,N_1285,N_1149);
xor U1913 (N_1913,N_1155,N_1279);
and U1914 (N_1914,N_1380,N_1319);
nand U1915 (N_1915,N_1146,N_1245);
nor U1916 (N_1916,N_1017,N_1413);
xor U1917 (N_1917,N_1048,N_1340);
nand U1918 (N_1918,N_1010,N_1184);
and U1919 (N_1919,N_1381,N_1438);
xor U1920 (N_1920,N_1296,N_1437);
nand U1921 (N_1921,N_1318,N_1334);
nor U1922 (N_1922,N_1190,N_1351);
nand U1923 (N_1923,N_1207,N_1297);
nor U1924 (N_1924,N_1053,N_1232);
or U1925 (N_1925,N_1240,N_1310);
nor U1926 (N_1926,N_1192,N_1415);
xor U1927 (N_1927,N_1399,N_1041);
or U1928 (N_1928,N_1124,N_1037);
nand U1929 (N_1929,N_1002,N_1447);
or U1930 (N_1930,N_1428,N_1378);
and U1931 (N_1931,N_1304,N_1486);
and U1932 (N_1932,N_1077,N_1349);
or U1933 (N_1933,N_1378,N_1273);
or U1934 (N_1934,N_1455,N_1047);
xnor U1935 (N_1935,N_1143,N_1010);
nor U1936 (N_1936,N_1287,N_1318);
and U1937 (N_1937,N_1016,N_1240);
xor U1938 (N_1938,N_1129,N_1068);
and U1939 (N_1939,N_1168,N_1138);
nor U1940 (N_1940,N_1145,N_1476);
or U1941 (N_1941,N_1030,N_1052);
xor U1942 (N_1942,N_1316,N_1282);
nand U1943 (N_1943,N_1474,N_1171);
and U1944 (N_1944,N_1432,N_1004);
nand U1945 (N_1945,N_1429,N_1371);
and U1946 (N_1946,N_1095,N_1474);
nand U1947 (N_1947,N_1358,N_1328);
or U1948 (N_1948,N_1254,N_1168);
nand U1949 (N_1949,N_1238,N_1096);
and U1950 (N_1950,N_1261,N_1427);
xor U1951 (N_1951,N_1130,N_1300);
or U1952 (N_1952,N_1185,N_1145);
and U1953 (N_1953,N_1306,N_1096);
xnor U1954 (N_1954,N_1132,N_1146);
nor U1955 (N_1955,N_1428,N_1417);
and U1956 (N_1956,N_1094,N_1205);
nand U1957 (N_1957,N_1453,N_1424);
nand U1958 (N_1958,N_1376,N_1359);
or U1959 (N_1959,N_1204,N_1388);
nand U1960 (N_1960,N_1056,N_1351);
xnor U1961 (N_1961,N_1379,N_1471);
nand U1962 (N_1962,N_1185,N_1408);
xnor U1963 (N_1963,N_1491,N_1049);
nor U1964 (N_1964,N_1213,N_1220);
xor U1965 (N_1965,N_1214,N_1290);
nor U1966 (N_1966,N_1396,N_1422);
xnor U1967 (N_1967,N_1360,N_1236);
xor U1968 (N_1968,N_1103,N_1039);
nand U1969 (N_1969,N_1042,N_1133);
or U1970 (N_1970,N_1271,N_1427);
xnor U1971 (N_1971,N_1389,N_1344);
and U1972 (N_1972,N_1078,N_1051);
nor U1973 (N_1973,N_1243,N_1435);
or U1974 (N_1974,N_1026,N_1448);
and U1975 (N_1975,N_1093,N_1304);
xnor U1976 (N_1976,N_1096,N_1109);
and U1977 (N_1977,N_1074,N_1153);
xor U1978 (N_1978,N_1181,N_1122);
nor U1979 (N_1979,N_1158,N_1260);
or U1980 (N_1980,N_1437,N_1002);
and U1981 (N_1981,N_1180,N_1379);
or U1982 (N_1982,N_1290,N_1124);
nor U1983 (N_1983,N_1260,N_1466);
xnor U1984 (N_1984,N_1124,N_1239);
nor U1985 (N_1985,N_1123,N_1321);
nor U1986 (N_1986,N_1078,N_1163);
and U1987 (N_1987,N_1056,N_1227);
and U1988 (N_1988,N_1056,N_1113);
nand U1989 (N_1989,N_1265,N_1212);
and U1990 (N_1990,N_1201,N_1476);
and U1991 (N_1991,N_1050,N_1175);
nand U1992 (N_1992,N_1391,N_1384);
xor U1993 (N_1993,N_1031,N_1186);
or U1994 (N_1994,N_1353,N_1260);
or U1995 (N_1995,N_1480,N_1196);
and U1996 (N_1996,N_1283,N_1358);
nor U1997 (N_1997,N_1238,N_1264);
or U1998 (N_1998,N_1402,N_1415);
xor U1999 (N_1999,N_1071,N_1226);
xnor U2000 (N_2000,N_1730,N_1574);
or U2001 (N_2001,N_1595,N_1839);
or U2002 (N_2002,N_1738,N_1723);
or U2003 (N_2003,N_1911,N_1653);
xnor U2004 (N_2004,N_1664,N_1817);
xnor U2005 (N_2005,N_1695,N_1756);
nor U2006 (N_2006,N_1554,N_1724);
nor U2007 (N_2007,N_1780,N_1994);
nor U2008 (N_2008,N_1900,N_1607);
nand U2009 (N_2009,N_1622,N_1733);
nand U2010 (N_2010,N_1890,N_1744);
or U2011 (N_2011,N_1950,N_1689);
nand U2012 (N_2012,N_1975,N_1552);
and U2013 (N_2013,N_1959,N_1840);
and U2014 (N_2014,N_1663,N_1625);
nor U2015 (N_2015,N_1675,N_1518);
and U2016 (N_2016,N_1617,N_1812);
and U2017 (N_2017,N_1714,N_1726);
and U2018 (N_2018,N_1854,N_1636);
nand U2019 (N_2019,N_1877,N_1510);
or U2020 (N_2020,N_1935,N_1519);
nor U2021 (N_2021,N_1741,N_1556);
xnor U2022 (N_2022,N_1543,N_1796);
nand U2023 (N_2023,N_1633,N_1502);
nor U2024 (N_2024,N_1860,N_1951);
and U2025 (N_2025,N_1932,N_1881);
xor U2026 (N_2026,N_1713,N_1962);
xor U2027 (N_2027,N_1568,N_1739);
or U2028 (N_2028,N_1609,N_1642);
nor U2029 (N_2029,N_1922,N_1832);
xnor U2030 (N_2030,N_1838,N_1761);
nor U2031 (N_2031,N_1864,N_1934);
and U2032 (N_2032,N_1997,N_1500);
nor U2033 (N_2033,N_1572,N_1637);
nand U2034 (N_2034,N_1711,N_1649);
nor U2035 (N_2035,N_1770,N_1575);
nor U2036 (N_2036,N_1912,N_1774);
nand U2037 (N_2037,N_1972,N_1512);
and U2038 (N_2038,N_1577,N_1676);
nand U2039 (N_2039,N_1810,N_1555);
nor U2040 (N_2040,N_1866,N_1528);
nor U2041 (N_2041,N_1674,N_1752);
nand U2042 (N_2042,N_1801,N_1677);
nand U2043 (N_2043,N_1580,N_1786);
nor U2044 (N_2044,N_1635,N_1837);
nor U2045 (N_2045,N_1542,N_1769);
xnor U2046 (N_2046,N_1843,N_1847);
and U2047 (N_2047,N_1954,N_1710);
nor U2048 (N_2048,N_1728,N_1971);
or U2049 (N_2049,N_1692,N_1930);
nand U2050 (N_2050,N_1524,N_1772);
or U2051 (N_2051,N_1589,N_1938);
nand U2052 (N_2052,N_1640,N_1682);
nor U2053 (N_2053,N_1665,N_1593);
and U2054 (N_2054,N_1899,N_1605);
nand U2055 (N_2055,N_1888,N_1883);
xor U2056 (N_2056,N_1787,N_1503);
xnor U2057 (N_2057,N_1944,N_1745);
nor U2058 (N_2058,N_1680,N_1978);
xor U2059 (N_2059,N_1852,N_1749);
nor U2060 (N_2060,N_1652,N_1616);
and U2061 (N_2061,N_1983,N_1757);
and U2062 (N_2062,N_1648,N_1981);
xnor U2063 (N_2063,N_1654,N_1816);
xor U2064 (N_2064,N_1514,N_1585);
and U2065 (N_2065,N_1594,N_1600);
and U2066 (N_2066,N_1529,N_1827);
nand U2067 (N_2067,N_1721,N_1579);
nand U2068 (N_2068,N_1910,N_1553);
xor U2069 (N_2069,N_1948,N_1725);
and U2070 (N_2070,N_1707,N_1992);
or U2071 (N_2071,N_1627,N_1591);
nand U2072 (N_2072,N_1976,N_1557);
nor U2073 (N_2073,N_1691,N_1586);
xor U2074 (N_2074,N_1919,N_1802);
xnor U2075 (N_2075,N_1768,N_1679);
nand U2076 (N_2076,N_1969,N_1766);
nor U2077 (N_2077,N_1647,N_1509);
or U2078 (N_2078,N_1566,N_1650);
or U2079 (N_2079,N_1779,N_1988);
and U2080 (N_2080,N_1957,N_1763);
or U2081 (N_2081,N_1611,N_1601);
xnor U2082 (N_2082,N_1578,N_1947);
nor U2083 (N_2083,N_1856,N_1753);
or U2084 (N_2084,N_1781,N_1771);
or U2085 (N_2085,N_1527,N_1719);
and U2086 (N_2086,N_1822,N_1598);
xor U2087 (N_2087,N_1828,N_1638);
nand U2088 (N_2088,N_1927,N_1630);
nor U2089 (N_2089,N_1920,N_1522);
nand U2090 (N_2090,N_1985,N_1987);
nand U2091 (N_2091,N_1865,N_1685);
nand U2092 (N_2092,N_1634,N_1823);
nand U2093 (N_2093,N_1966,N_1955);
nor U2094 (N_2094,N_1884,N_1909);
xor U2095 (N_2095,N_1708,N_1914);
xnor U2096 (N_2096,N_1731,N_1621);
nand U2097 (N_2097,N_1546,N_1850);
and U2098 (N_2098,N_1597,N_1690);
nand U2099 (N_2099,N_1808,N_1937);
nor U2100 (N_2100,N_1820,N_1945);
nand U2101 (N_2101,N_1933,N_1882);
nand U2102 (N_2102,N_1742,N_1619);
nand U2103 (N_2103,N_1946,N_1809);
and U2104 (N_2104,N_1803,N_1508);
xor U2105 (N_2105,N_1861,N_1513);
nor U2106 (N_2106,N_1655,N_1525);
nand U2107 (N_2107,N_1869,N_1658);
nor U2108 (N_2108,N_1748,N_1788);
or U2109 (N_2109,N_1902,N_1567);
nor U2110 (N_2110,N_1558,N_1942);
xnor U2111 (N_2111,N_1806,N_1657);
or U2112 (N_2112,N_1949,N_1547);
xor U2113 (N_2113,N_1829,N_1903);
nor U2114 (N_2114,N_1516,N_1582);
or U2115 (N_2115,N_1639,N_1693);
nand U2116 (N_2116,N_1700,N_1551);
nand U2117 (N_2117,N_1530,N_1610);
and U2118 (N_2118,N_1686,N_1926);
or U2119 (N_2119,N_1506,N_1683);
nand U2120 (N_2120,N_1576,N_1734);
nor U2121 (N_2121,N_1751,N_1931);
and U2122 (N_2122,N_1991,N_1620);
nor U2123 (N_2123,N_1868,N_1520);
nor U2124 (N_2124,N_1684,N_1952);
and U2125 (N_2125,N_1924,N_1886);
and U2126 (N_2126,N_1818,N_1821);
xnor U2127 (N_2127,N_1778,N_1505);
xnor U2128 (N_2128,N_1631,N_1662);
nor U2129 (N_2129,N_1897,N_1916);
and U2130 (N_2130,N_1697,N_1858);
and U2131 (N_2131,N_1590,N_1974);
xor U2132 (N_2132,N_1602,N_1592);
nor U2133 (N_2133,N_1727,N_1996);
xnor U2134 (N_2134,N_1973,N_1666);
nor U2135 (N_2135,N_1583,N_1917);
nor U2136 (N_2136,N_1549,N_1878);
xor U2137 (N_2137,N_1867,N_1737);
nand U2138 (N_2138,N_1792,N_1815);
or U2139 (N_2139,N_1504,N_1669);
xnor U2140 (N_2140,N_1716,N_1501);
or U2141 (N_2141,N_1797,N_1782);
xor U2142 (N_2142,N_1699,N_1898);
xnor U2143 (N_2143,N_1961,N_1805);
xor U2144 (N_2144,N_1963,N_1628);
nand U2145 (N_2145,N_1862,N_1750);
and U2146 (N_2146,N_1703,N_1535);
xor U2147 (N_2147,N_1783,N_1776);
xor U2148 (N_2148,N_1613,N_1706);
xnor U2149 (N_2149,N_1773,N_1587);
nor U2150 (N_2150,N_1672,N_1893);
nor U2151 (N_2151,N_1717,N_1561);
nor U2152 (N_2152,N_1800,N_1863);
nor U2153 (N_2153,N_1762,N_1841);
or U2154 (N_2154,N_1618,N_1901);
xnor U2155 (N_2155,N_1507,N_1671);
xnor U2156 (N_2156,N_1784,N_1967);
or U2157 (N_2157,N_1887,N_1876);
nor U2158 (N_2158,N_1785,N_1874);
xnor U2159 (N_2159,N_1807,N_1831);
xnor U2160 (N_2160,N_1645,N_1571);
and U2161 (N_2161,N_1569,N_1775);
nand U2162 (N_2162,N_1581,N_1906);
or U2163 (N_2163,N_1764,N_1533);
nand U2164 (N_2164,N_1895,N_1790);
nor U2165 (N_2165,N_1688,N_1641);
and U2166 (N_2166,N_1767,N_1646);
and U2167 (N_2167,N_1588,N_1999);
nand U2168 (N_2168,N_1718,N_1870);
nor U2169 (N_2169,N_1941,N_1848);
or U2170 (N_2170,N_1825,N_1824);
nand U2171 (N_2171,N_1842,N_1704);
nand U2172 (N_2172,N_1758,N_1956);
xnor U2173 (N_2173,N_1939,N_1844);
and U2174 (N_2174,N_1880,N_1584);
nand U2175 (N_2175,N_1537,N_1965);
or U2176 (N_2176,N_1830,N_1702);
or U2177 (N_2177,N_1564,N_1875);
xor U2178 (N_2178,N_1980,N_1521);
nand U2179 (N_2179,N_1921,N_1722);
nor U2180 (N_2180,N_1755,N_1612);
or U2181 (N_2181,N_1857,N_1923);
and U2182 (N_2182,N_1615,N_1929);
and U2183 (N_2183,N_1536,N_1604);
and U2184 (N_2184,N_1913,N_1885);
nor U2185 (N_2185,N_1562,N_1896);
or U2186 (N_2186,N_1735,N_1979);
or U2187 (N_2187,N_1759,N_1517);
nor U2188 (N_2188,N_1565,N_1940);
nand U2189 (N_2189,N_1908,N_1993);
and U2190 (N_2190,N_1813,N_1643);
or U2191 (N_2191,N_1541,N_1970);
nor U2192 (N_2192,N_1990,N_1599);
or U2193 (N_2193,N_1960,N_1608);
and U2194 (N_2194,N_1836,N_1743);
nor U2195 (N_2195,N_1667,N_1539);
nand U2196 (N_2196,N_1661,N_1523);
nor U2197 (N_2197,N_1540,N_1977);
and U2198 (N_2198,N_1747,N_1698);
and U2199 (N_2199,N_1964,N_1907);
nor U2200 (N_2200,N_1936,N_1563);
nor U2201 (N_2201,N_1729,N_1573);
nor U2202 (N_2202,N_1559,N_1915);
xnor U2203 (N_2203,N_1548,N_1789);
nand U2204 (N_2204,N_1705,N_1891);
or U2205 (N_2205,N_1835,N_1894);
or U2206 (N_2206,N_1968,N_1793);
or U2207 (N_2207,N_1720,N_1853);
nand U2208 (N_2208,N_1732,N_1550);
nor U2209 (N_2209,N_1928,N_1632);
nand U2210 (N_2210,N_1681,N_1760);
nor U2211 (N_2211,N_1531,N_1791);
xor U2212 (N_2212,N_1626,N_1943);
xnor U2213 (N_2213,N_1795,N_1998);
nor U2214 (N_2214,N_1614,N_1532);
nor U2215 (N_2215,N_1656,N_1765);
xor U2216 (N_2216,N_1958,N_1740);
nand U2217 (N_2217,N_1694,N_1570);
or U2218 (N_2218,N_1709,N_1660);
or U2219 (N_2219,N_1982,N_1814);
xnor U2220 (N_2220,N_1603,N_1855);
or U2221 (N_2221,N_1644,N_1871);
nor U2222 (N_2222,N_1892,N_1873);
xnor U2223 (N_2223,N_1606,N_1798);
or U2224 (N_2224,N_1925,N_1715);
or U2225 (N_2225,N_1986,N_1526);
or U2226 (N_2226,N_1712,N_1624);
nand U2227 (N_2227,N_1995,N_1984);
nand U2228 (N_2228,N_1538,N_1696);
and U2229 (N_2229,N_1754,N_1670);
xor U2230 (N_2230,N_1879,N_1777);
and U2231 (N_2231,N_1651,N_1687);
and U2232 (N_2232,N_1668,N_1544);
and U2233 (N_2233,N_1746,N_1819);
or U2234 (N_2234,N_1534,N_1799);
and U2235 (N_2235,N_1833,N_1659);
nand U2236 (N_2236,N_1678,N_1904);
and U2237 (N_2237,N_1596,N_1845);
nand U2238 (N_2238,N_1511,N_1889);
nor U2239 (N_2239,N_1629,N_1736);
or U2240 (N_2240,N_1851,N_1859);
nor U2241 (N_2241,N_1515,N_1701);
nor U2242 (N_2242,N_1989,N_1872);
xnor U2243 (N_2243,N_1834,N_1623);
and U2244 (N_2244,N_1811,N_1846);
or U2245 (N_2245,N_1953,N_1804);
nand U2246 (N_2246,N_1673,N_1905);
or U2247 (N_2247,N_1826,N_1849);
and U2248 (N_2248,N_1560,N_1918);
or U2249 (N_2249,N_1794,N_1545);
or U2250 (N_2250,N_1612,N_1730);
nor U2251 (N_2251,N_1910,N_1843);
and U2252 (N_2252,N_1858,N_1931);
nor U2253 (N_2253,N_1808,N_1944);
xnor U2254 (N_2254,N_1860,N_1838);
xor U2255 (N_2255,N_1601,N_1842);
xnor U2256 (N_2256,N_1525,N_1605);
or U2257 (N_2257,N_1537,N_1637);
or U2258 (N_2258,N_1771,N_1782);
nor U2259 (N_2259,N_1832,N_1556);
nor U2260 (N_2260,N_1601,N_1976);
xnor U2261 (N_2261,N_1802,N_1510);
and U2262 (N_2262,N_1864,N_1542);
and U2263 (N_2263,N_1846,N_1840);
and U2264 (N_2264,N_1656,N_1516);
xnor U2265 (N_2265,N_1983,N_1824);
or U2266 (N_2266,N_1774,N_1809);
or U2267 (N_2267,N_1892,N_1871);
and U2268 (N_2268,N_1935,N_1508);
nor U2269 (N_2269,N_1961,N_1550);
nor U2270 (N_2270,N_1786,N_1569);
or U2271 (N_2271,N_1626,N_1796);
or U2272 (N_2272,N_1501,N_1611);
nand U2273 (N_2273,N_1589,N_1728);
and U2274 (N_2274,N_1507,N_1643);
xor U2275 (N_2275,N_1736,N_1936);
nand U2276 (N_2276,N_1632,N_1747);
and U2277 (N_2277,N_1875,N_1511);
or U2278 (N_2278,N_1779,N_1976);
or U2279 (N_2279,N_1705,N_1964);
or U2280 (N_2280,N_1956,N_1749);
and U2281 (N_2281,N_1606,N_1976);
or U2282 (N_2282,N_1774,N_1800);
nor U2283 (N_2283,N_1730,N_1848);
nand U2284 (N_2284,N_1598,N_1865);
nand U2285 (N_2285,N_1997,N_1792);
and U2286 (N_2286,N_1531,N_1559);
nand U2287 (N_2287,N_1970,N_1664);
and U2288 (N_2288,N_1561,N_1923);
xor U2289 (N_2289,N_1942,N_1888);
and U2290 (N_2290,N_1990,N_1687);
or U2291 (N_2291,N_1778,N_1834);
xor U2292 (N_2292,N_1825,N_1817);
nand U2293 (N_2293,N_1505,N_1624);
xor U2294 (N_2294,N_1827,N_1601);
or U2295 (N_2295,N_1644,N_1949);
nor U2296 (N_2296,N_1743,N_1872);
nor U2297 (N_2297,N_1526,N_1528);
xor U2298 (N_2298,N_1633,N_1878);
or U2299 (N_2299,N_1833,N_1732);
nor U2300 (N_2300,N_1508,N_1550);
nand U2301 (N_2301,N_1682,N_1689);
nand U2302 (N_2302,N_1558,N_1577);
nor U2303 (N_2303,N_1529,N_1818);
and U2304 (N_2304,N_1938,N_1966);
nor U2305 (N_2305,N_1552,N_1795);
and U2306 (N_2306,N_1839,N_1981);
nand U2307 (N_2307,N_1726,N_1597);
xor U2308 (N_2308,N_1905,N_1963);
nor U2309 (N_2309,N_1859,N_1897);
or U2310 (N_2310,N_1908,N_1728);
or U2311 (N_2311,N_1641,N_1814);
and U2312 (N_2312,N_1793,N_1501);
or U2313 (N_2313,N_1782,N_1566);
nor U2314 (N_2314,N_1886,N_1721);
xnor U2315 (N_2315,N_1947,N_1507);
or U2316 (N_2316,N_1881,N_1948);
nor U2317 (N_2317,N_1755,N_1809);
nand U2318 (N_2318,N_1940,N_1784);
and U2319 (N_2319,N_1585,N_1866);
nand U2320 (N_2320,N_1633,N_1813);
or U2321 (N_2321,N_1829,N_1597);
nor U2322 (N_2322,N_1876,N_1632);
and U2323 (N_2323,N_1613,N_1930);
and U2324 (N_2324,N_1543,N_1999);
nor U2325 (N_2325,N_1826,N_1998);
and U2326 (N_2326,N_1749,N_1837);
nor U2327 (N_2327,N_1927,N_1857);
and U2328 (N_2328,N_1683,N_1637);
nor U2329 (N_2329,N_1723,N_1534);
and U2330 (N_2330,N_1746,N_1937);
nand U2331 (N_2331,N_1687,N_1824);
xnor U2332 (N_2332,N_1723,N_1907);
nor U2333 (N_2333,N_1526,N_1954);
xor U2334 (N_2334,N_1762,N_1579);
xnor U2335 (N_2335,N_1965,N_1764);
and U2336 (N_2336,N_1646,N_1937);
nor U2337 (N_2337,N_1930,N_1720);
nand U2338 (N_2338,N_1639,N_1949);
and U2339 (N_2339,N_1585,N_1503);
xor U2340 (N_2340,N_1713,N_1772);
xnor U2341 (N_2341,N_1759,N_1657);
or U2342 (N_2342,N_1885,N_1896);
and U2343 (N_2343,N_1792,N_1605);
or U2344 (N_2344,N_1980,N_1559);
and U2345 (N_2345,N_1559,N_1583);
and U2346 (N_2346,N_1562,N_1973);
and U2347 (N_2347,N_1734,N_1589);
and U2348 (N_2348,N_1874,N_1695);
and U2349 (N_2349,N_1798,N_1978);
xor U2350 (N_2350,N_1640,N_1750);
or U2351 (N_2351,N_1524,N_1849);
xor U2352 (N_2352,N_1574,N_1759);
nor U2353 (N_2353,N_1910,N_1745);
xor U2354 (N_2354,N_1882,N_1810);
nor U2355 (N_2355,N_1891,N_1877);
and U2356 (N_2356,N_1884,N_1851);
nand U2357 (N_2357,N_1652,N_1687);
nor U2358 (N_2358,N_1605,N_1548);
nor U2359 (N_2359,N_1540,N_1523);
nand U2360 (N_2360,N_1788,N_1607);
or U2361 (N_2361,N_1940,N_1597);
nand U2362 (N_2362,N_1844,N_1702);
nor U2363 (N_2363,N_1696,N_1996);
nor U2364 (N_2364,N_1974,N_1738);
nand U2365 (N_2365,N_1533,N_1723);
or U2366 (N_2366,N_1713,N_1847);
or U2367 (N_2367,N_1711,N_1729);
nor U2368 (N_2368,N_1577,N_1615);
xor U2369 (N_2369,N_1606,N_1861);
nand U2370 (N_2370,N_1690,N_1914);
or U2371 (N_2371,N_1997,N_1607);
nand U2372 (N_2372,N_1646,N_1934);
nor U2373 (N_2373,N_1792,N_1678);
or U2374 (N_2374,N_1819,N_1832);
nor U2375 (N_2375,N_1604,N_1778);
nor U2376 (N_2376,N_1790,N_1548);
and U2377 (N_2377,N_1717,N_1671);
nand U2378 (N_2378,N_1866,N_1764);
or U2379 (N_2379,N_1950,N_1773);
xnor U2380 (N_2380,N_1713,N_1915);
nand U2381 (N_2381,N_1872,N_1754);
xnor U2382 (N_2382,N_1824,N_1904);
nand U2383 (N_2383,N_1841,N_1815);
xnor U2384 (N_2384,N_1500,N_1560);
nor U2385 (N_2385,N_1995,N_1799);
nor U2386 (N_2386,N_1621,N_1637);
nor U2387 (N_2387,N_1616,N_1584);
xor U2388 (N_2388,N_1529,N_1924);
or U2389 (N_2389,N_1842,N_1847);
nor U2390 (N_2390,N_1564,N_1939);
nand U2391 (N_2391,N_1503,N_1704);
or U2392 (N_2392,N_1602,N_1816);
xor U2393 (N_2393,N_1598,N_1765);
or U2394 (N_2394,N_1849,N_1595);
xor U2395 (N_2395,N_1743,N_1711);
or U2396 (N_2396,N_1524,N_1971);
nand U2397 (N_2397,N_1789,N_1980);
xnor U2398 (N_2398,N_1767,N_1671);
or U2399 (N_2399,N_1534,N_1631);
nand U2400 (N_2400,N_1663,N_1878);
nor U2401 (N_2401,N_1666,N_1840);
nor U2402 (N_2402,N_1574,N_1724);
nor U2403 (N_2403,N_1939,N_1676);
and U2404 (N_2404,N_1636,N_1507);
or U2405 (N_2405,N_1518,N_1834);
nand U2406 (N_2406,N_1942,N_1770);
nor U2407 (N_2407,N_1622,N_1958);
nand U2408 (N_2408,N_1947,N_1573);
nor U2409 (N_2409,N_1819,N_1703);
or U2410 (N_2410,N_1822,N_1893);
xnor U2411 (N_2411,N_1886,N_1836);
nor U2412 (N_2412,N_1918,N_1880);
and U2413 (N_2413,N_1665,N_1922);
nor U2414 (N_2414,N_1771,N_1918);
nor U2415 (N_2415,N_1805,N_1556);
and U2416 (N_2416,N_1599,N_1606);
or U2417 (N_2417,N_1772,N_1799);
xnor U2418 (N_2418,N_1525,N_1902);
or U2419 (N_2419,N_1760,N_1713);
or U2420 (N_2420,N_1546,N_1814);
nor U2421 (N_2421,N_1981,N_1751);
xnor U2422 (N_2422,N_1792,N_1735);
or U2423 (N_2423,N_1622,N_1837);
nor U2424 (N_2424,N_1932,N_1576);
and U2425 (N_2425,N_1867,N_1747);
or U2426 (N_2426,N_1646,N_1790);
nor U2427 (N_2427,N_1863,N_1782);
nand U2428 (N_2428,N_1833,N_1964);
nor U2429 (N_2429,N_1994,N_1611);
and U2430 (N_2430,N_1910,N_1740);
nand U2431 (N_2431,N_1859,N_1964);
or U2432 (N_2432,N_1628,N_1713);
xor U2433 (N_2433,N_1916,N_1710);
xnor U2434 (N_2434,N_1783,N_1579);
nor U2435 (N_2435,N_1927,N_1838);
nor U2436 (N_2436,N_1683,N_1897);
nor U2437 (N_2437,N_1692,N_1821);
nor U2438 (N_2438,N_1829,N_1591);
or U2439 (N_2439,N_1581,N_1739);
or U2440 (N_2440,N_1535,N_1618);
xnor U2441 (N_2441,N_1687,N_1696);
xnor U2442 (N_2442,N_1916,N_1701);
nand U2443 (N_2443,N_1610,N_1733);
xor U2444 (N_2444,N_1954,N_1893);
nand U2445 (N_2445,N_1877,N_1951);
nor U2446 (N_2446,N_1872,N_1799);
or U2447 (N_2447,N_1853,N_1877);
and U2448 (N_2448,N_1928,N_1917);
xnor U2449 (N_2449,N_1753,N_1783);
or U2450 (N_2450,N_1978,N_1892);
and U2451 (N_2451,N_1745,N_1767);
nand U2452 (N_2452,N_1777,N_1530);
xnor U2453 (N_2453,N_1884,N_1659);
nand U2454 (N_2454,N_1782,N_1820);
xnor U2455 (N_2455,N_1733,N_1638);
xor U2456 (N_2456,N_1986,N_1749);
or U2457 (N_2457,N_1945,N_1763);
or U2458 (N_2458,N_1859,N_1658);
or U2459 (N_2459,N_1909,N_1936);
xnor U2460 (N_2460,N_1680,N_1990);
nor U2461 (N_2461,N_1774,N_1760);
or U2462 (N_2462,N_1619,N_1850);
nand U2463 (N_2463,N_1819,N_1616);
xnor U2464 (N_2464,N_1617,N_1794);
or U2465 (N_2465,N_1593,N_1922);
nor U2466 (N_2466,N_1559,N_1513);
and U2467 (N_2467,N_1707,N_1854);
nor U2468 (N_2468,N_1986,N_1995);
or U2469 (N_2469,N_1643,N_1731);
nand U2470 (N_2470,N_1960,N_1746);
or U2471 (N_2471,N_1930,N_1825);
or U2472 (N_2472,N_1568,N_1689);
and U2473 (N_2473,N_1697,N_1987);
nor U2474 (N_2474,N_1910,N_1668);
xnor U2475 (N_2475,N_1994,N_1928);
and U2476 (N_2476,N_1692,N_1618);
or U2477 (N_2477,N_1899,N_1920);
or U2478 (N_2478,N_1975,N_1576);
nand U2479 (N_2479,N_1952,N_1907);
xor U2480 (N_2480,N_1917,N_1867);
or U2481 (N_2481,N_1841,N_1931);
and U2482 (N_2482,N_1850,N_1509);
nand U2483 (N_2483,N_1553,N_1971);
or U2484 (N_2484,N_1738,N_1683);
and U2485 (N_2485,N_1964,N_1527);
nor U2486 (N_2486,N_1686,N_1883);
nand U2487 (N_2487,N_1684,N_1946);
or U2488 (N_2488,N_1602,N_1815);
nand U2489 (N_2489,N_1842,N_1873);
or U2490 (N_2490,N_1716,N_1773);
or U2491 (N_2491,N_1502,N_1800);
and U2492 (N_2492,N_1750,N_1532);
nand U2493 (N_2493,N_1705,N_1812);
nor U2494 (N_2494,N_1669,N_1536);
and U2495 (N_2495,N_1527,N_1596);
nor U2496 (N_2496,N_1513,N_1975);
and U2497 (N_2497,N_1804,N_1583);
xor U2498 (N_2498,N_1830,N_1520);
xnor U2499 (N_2499,N_1958,N_1585);
nor U2500 (N_2500,N_2459,N_2424);
nand U2501 (N_2501,N_2045,N_2161);
nor U2502 (N_2502,N_2368,N_2071);
or U2503 (N_2503,N_2474,N_2443);
xor U2504 (N_2504,N_2198,N_2061);
xnor U2505 (N_2505,N_2421,N_2313);
nor U2506 (N_2506,N_2435,N_2302);
and U2507 (N_2507,N_2453,N_2070);
xnor U2508 (N_2508,N_2034,N_2401);
or U2509 (N_2509,N_2239,N_2100);
or U2510 (N_2510,N_2094,N_2301);
xnor U2511 (N_2511,N_2022,N_2457);
xor U2512 (N_2512,N_2321,N_2021);
xor U2513 (N_2513,N_2107,N_2308);
and U2514 (N_2514,N_2402,N_2063);
or U2515 (N_2515,N_2012,N_2188);
xnor U2516 (N_2516,N_2290,N_2440);
and U2517 (N_2517,N_2004,N_2108);
nor U2518 (N_2518,N_2231,N_2236);
nor U2519 (N_2519,N_2078,N_2307);
xor U2520 (N_2520,N_2158,N_2297);
or U2521 (N_2521,N_2284,N_2164);
nor U2522 (N_2522,N_2476,N_2417);
xor U2523 (N_2523,N_2344,N_2254);
xor U2524 (N_2524,N_2466,N_2408);
or U2525 (N_2525,N_2163,N_2358);
or U2526 (N_2526,N_2056,N_2388);
or U2527 (N_2527,N_2391,N_2212);
nand U2528 (N_2528,N_2199,N_2362);
nand U2529 (N_2529,N_2088,N_2327);
xor U2530 (N_2530,N_2248,N_2084);
xnor U2531 (N_2531,N_2037,N_2393);
and U2532 (N_2532,N_2287,N_2291);
or U2533 (N_2533,N_2383,N_2354);
nor U2534 (N_2534,N_2186,N_2222);
nor U2535 (N_2535,N_2109,N_2335);
or U2536 (N_2536,N_2376,N_2489);
nand U2537 (N_2537,N_2110,N_2444);
xnor U2538 (N_2538,N_2389,N_2085);
xor U2539 (N_2539,N_2104,N_2170);
and U2540 (N_2540,N_2140,N_2083);
nor U2541 (N_2541,N_2058,N_2385);
and U2542 (N_2542,N_2018,N_2378);
and U2543 (N_2543,N_2067,N_2487);
xnor U2544 (N_2544,N_2000,N_2255);
nor U2545 (N_2545,N_2230,N_2452);
nand U2546 (N_2546,N_2431,N_2132);
nand U2547 (N_2547,N_2266,N_2166);
xnor U2548 (N_2548,N_2304,N_2364);
and U2549 (N_2549,N_2324,N_2180);
nand U2550 (N_2550,N_2412,N_2332);
nand U2551 (N_2551,N_2423,N_2075);
or U2552 (N_2552,N_2325,N_2374);
nand U2553 (N_2553,N_2322,N_2151);
nand U2554 (N_2554,N_2283,N_2130);
or U2555 (N_2555,N_2319,N_2008);
nand U2556 (N_2556,N_2282,N_2146);
nand U2557 (N_2557,N_2079,N_2098);
or U2558 (N_2558,N_2205,N_2041);
or U2559 (N_2559,N_2211,N_2272);
and U2560 (N_2560,N_2442,N_2315);
nand U2561 (N_2561,N_2365,N_2405);
and U2562 (N_2562,N_2187,N_2481);
or U2563 (N_2563,N_2305,N_2139);
nand U2564 (N_2564,N_2455,N_2360);
or U2565 (N_2565,N_2395,N_2114);
or U2566 (N_2566,N_2415,N_2044);
or U2567 (N_2567,N_2448,N_2386);
and U2568 (N_2568,N_2330,N_2010);
and U2569 (N_2569,N_2251,N_2135);
nor U2570 (N_2570,N_2207,N_2080);
and U2571 (N_2571,N_2495,N_2156);
nor U2572 (N_2572,N_2019,N_2128);
or U2573 (N_2573,N_2030,N_2095);
nor U2574 (N_2574,N_2296,N_2203);
and U2575 (N_2575,N_2329,N_2249);
and U2576 (N_2576,N_2215,N_2064);
or U2577 (N_2577,N_2072,N_2043);
or U2578 (N_2578,N_2150,N_2181);
or U2579 (N_2579,N_2125,N_2160);
nor U2580 (N_2580,N_2377,N_2261);
and U2581 (N_2581,N_2191,N_2102);
or U2582 (N_2582,N_2285,N_2055);
xnor U2583 (N_2583,N_2122,N_2176);
or U2584 (N_2584,N_2407,N_2042);
nor U2585 (N_2585,N_2007,N_2038);
xor U2586 (N_2586,N_2026,N_2464);
nor U2587 (N_2587,N_2023,N_2482);
nand U2588 (N_2588,N_2472,N_2220);
nand U2589 (N_2589,N_2143,N_2197);
and U2590 (N_2590,N_2338,N_2372);
or U2591 (N_2591,N_2468,N_2480);
and U2592 (N_2592,N_2001,N_2003);
nor U2593 (N_2593,N_2097,N_2300);
and U2594 (N_2594,N_2387,N_2185);
nor U2595 (N_2595,N_2265,N_2089);
nand U2596 (N_2596,N_2036,N_2101);
and U2597 (N_2597,N_2491,N_2214);
nand U2598 (N_2598,N_2024,N_2062);
nand U2599 (N_2599,N_2183,N_2414);
nand U2600 (N_2600,N_2317,N_2367);
nor U2601 (N_2601,N_2292,N_2429);
and U2602 (N_2602,N_2328,N_2121);
or U2603 (N_2603,N_2069,N_2277);
or U2604 (N_2604,N_2134,N_2171);
or U2605 (N_2605,N_2047,N_2194);
and U2606 (N_2606,N_2303,N_2493);
nor U2607 (N_2607,N_2339,N_2438);
nor U2608 (N_2608,N_2390,N_2233);
nand U2609 (N_2609,N_2015,N_2473);
nand U2610 (N_2610,N_2373,N_2051);
or U2611 (N_2611,N_2294,N_2419);
or U2612 (N_2612,N_2425,N_2040);
nor U2613 (N_2613,N_2485,N_2127);
nor U2614 (N_2614,N_2342,N_2092);
xor U2615 (N_2615,N_2250,N_2357);
and U2616 (N_2616,N_2426,N_2142);
or U2617 (N_2617,N_2208,N_2123);
xor U2618 (N_2618,N_2093,N_2352);
and U2619 (N_2619,N_2053,N_2269);
nand U2620 (N_2620,N_2168,N_2420);
and U2621 (N_2621,N_2394,N_2178);
nor U2622 (N_2622,N_2226,N_2375);
nor U2623 (N_2623,N_2437,N_2106);
nand U2624 (N_2624,N_2234,N_2157);
xor U2625 (N_2625,N_2016,N_2117);
or U2626 (N_2626,N_2068,N_2065);
nand U2627 (N_2627,N_2293,N_2210);
or U2628 (N_2628,N_2011,N_2082);
or U2629 (N_2629,N_2309,N_2049);
nor U2630 (N_2630,N_2032,N_2430);
and U2631 (N_2631,N_2346,N_2103);
and U2632 (N_2632,N_2242,N_2411);
or U2633 (N_2633,N_2155,N_2190);
or U2634 (N_2634,N_2380,N_2073);
and U2635 (N_2635,N_2091,N_2033);
and U2636 (N_2636,N_2116,N_2439);
xor U2637 (N_2637,N_2275,N_2488);
or U2638 (N_2638,N_2099,N_2148);
nand U2639 (N_2639,N_2252,N_2247);
xor U2640 (N_2640,N_2175,N_2462);
xor U2641 (N_2641,N_2316,N_2235);
and U2642 (N_2642,N_2490,N_2138);
nor U2643 (N_2643,N_2396,N_2471);
nor U2644 (N_2644,N_2469,N_2418);
nor U2645 (N_2645,N_2258,N_2461);
nand U2646 (N_2646,N_2081,N_2113);
nor U2647 (N_2647,N_2406,N_2066);
nand U2648 (N_2648,N_2299,N_2144);
nand U2649 (N_2649,N_2147,N_2312);
or U2650 (N_2650,N_2281,N_2483);
or U2651 (N_2651,N_2031,N_2499);
or U2652 (N_2652,N_2286,N_2154);
nor U2653 (N_2653,N_2165,N_2223);
nor U2654 (N_2654,N_2382,N_2460);
xor U2655 (N_2655,N_2363,N_2172);
xnor U2656 (N_2656,N_2416,N_2274);
and U2657 (N_2657,N_2337,N_2475);
xnor U2658 (N_2658,N_2264,N_2028);
nor U2659 (N_2659,N_2341,N_2177);
nor U2660 (N_2660,N_2369,N_2349);
xnor U2661 (N_2661,N_2027,N_2257);
xor U2662 (N_2662,N_2167,N_2355);
or U2663 (N_2663,N_2436,N_2351);
or U2664 (N_2664,N_2450,N_2217);
nand U2665 (N_2665,N_2115,N_2074);
xor U2666 (N_2666,N_2298,N_2020);
nand U2667 (N_2667,N_2280,N_2174);
or U2668 (N_2668,N_2263,N_2314);
nand U2669 (N_2669,N_2209,N_2306);
and U2670 (N_2670,N_2105,N_2054);
xor U2671 (N_2671,N_2278,N_2048);
nand U2672 (N_2672,N_2271,N_2124);
or U2673 (N_2673,N_2240,N_2111);
and U2674 (N_2674,N_2359,N_2323);
nand U2675 (N_2675,N_2189,N_2295);
and U2676 (N_2676,N_2361,N_2433);
xor U2677 (N_2677,N_2318,N_2410);
xnor U2678 (N_2678,N_2087,N_2029);
nand U2679 (N_2679,N_2467,N_2447);
nand U2680 (N_2680,N_2289,N_2398);
nand U2681 (N_2681,N_2403,N_2347);
and U2682 (N_2682,N_2225,N_2077);
nor U2683 (N_2683,N_2159,N_2486);
nand U2684 (N_2684,N_2076,N_2152);
nand U2685 (N_2685,N_2141,N_2434);
nor U2686 (N_2686,N_2484,N_2201);
nand U2687 (N_2687,N_2131,N_2002);
xnor U2688 (N_2688,N_2463,N_2136);
nor U2689 (N_2689,N_2013,N_2149);
nor U2690 (N_2690,N_2413,N_2126);
nor U2691 (N_2691,N_2059,N_2422);
nand U2692 (N_2692,N_2392,N_2381);
and U2693 (N_2693,N_2279,N_2245);
xor U2694 (N_2694,N_2244,N_2006);
xnor U2695 (N_2695,N_2118,N_2454);
and U2696 (N_2696,N_2005,N_2432);
nand U2697 (N_2697,N_2017,N_2227);
xor U2698 (N_2698,N_2397,N_2276);
or U2699 (N_2699,N_2228,N_2046);
and U2700 (N_2700,N_2238,N_2273);
nor U2701 (N_2701,N_2345,N_2311);
nand U2702 (N_2702,N_2267,N_2241);
or U2703 (N_2703,N_2404,N_2458);
xor U2704 (N_2704,N_2137,N_2182);
nor U2705 (N_2705,N_2206,N_2162);
nor U2706 (N_2706,N_2129,N_2343);
xor U2707 (N_2707,N_2451,N_2259);
or U2708 (N_2708,N_2334,N_2173);
nand U2709 (N_2709,N_2014,N_2492);
xor U2710 (N_2710,N_2246,N_2213);
or U2711 (N_2711,N_2195,N_2052);
nand U2712 (N_2712,N_2370,N_2192);
nor U2713 (N_2713,N_2153,N_2193);
nand U2714 (N_2714,N_2356,N_2243);
xnor U2715 (N_2715,N_2200,N_2253);
nand U2716 (N_2716,N_2112,N_2310);
and U2717 (N_2717,N_2477,N_2456);
or U2718 (N_2718,N_2090,N_2145);
nand U2719 (N_2719,N_2384,N_2409);
nor U2720 (N_2720,N_2256,N_2202);
and U2721 (N_2721,N_2379,N_2035);
nand U2722 (N_2722,N_2366,N_2498);
or U2723 (N_2723,N_2009,N_2270);
and U2724 (N_2724,N_2441,N_2260);
nor U2725 (N_2725,N_2096,N_2216);
nor U2726 (N_2726,N_2086,N_2494);
nor U2727 (N_2727,N_2399,N_2219);
nand U2728 (N_2728,N_2336,N_2169);
nand U2729 (N_2729,N_2446,N_2039);
xnor U2730 (N_2730,N_2427,N_2371);
nor U2731 (N_2731,N_2050,N_2465);
and U2732 (N_2732,N_2470,N_2326);
nor U2733 (N_2733,N_2428,N_2445);
nand U2734 (N_2734,N_2133,N_2262);
and U2735 (N_2735,N_2340,N_2353);
or U2736 (N_2736,N_2479,N_2057);
and U2737 (N_2737,N_2497,N_2400);
nor U2738 (N_2738,N_2232,N_2348);
nand U2739 (N_2739,N_2119,N_2229);
xor U2740 (N_2740,N_2288,N_2204);
nand U2741 (N_2741,N_2179,N_2478);
xnor U2742 (N_2742,N_2333,N_2268);
nand U2743 (N_2743,N_2120,N_2184);
xor U2744 (N_2744,N_2196,N_2331);
nand U2745 (N_2745,N_2496,N_2221);
nand U2746 (N_2746,N_2025,N_2449);
or U2747 (N_2747,N_2218,N_2237);
xnor U2748 (N_2748,N_2320,N_2060);
nand U2749 (N_2749,N_2350,N_2224);
and U2750 (N_2750,N_2308,N_2143);
nand U2751 (N_2751,N_2320,N_2471);
and U2752 (N_2752,N_2239,N_2136);
and U2753 (N_2753,N_2082,N_2330);
nor U2754 (N_2754,N_2041,N_2158);
and U2755 (N_2755,N_2487,N_2335);
xnor U2756 (N_2756,N_2241,N_2124);
and U2757 (N_2757,N_2152,N_2060);
and U2758 (N_2758,N_2392,N_2317);
and U2759 (N_2759,N_2306,N_2421);
nor U2760 (N_2760,N_2144,N_2352);
nor U2761 (N_2761,N_2123,N_2298);
and U2762 (N_2762,N_2223,N_2236);
or U2763 (N_2763,N_2254,N_2034);
or U2764 (N_2764,N_2090,N_2247);
or U2765 (N_2765,N_2014,N_2292);
nor U2766 (N_2766,N_2232,N_2373);
nor U2767 (N_2767,N_2286,N_2395);
nor U2768 (N_2768,N_2489,N_2246);
and U2769 (N_2769,N_2250,N_2499);
and U2770 (N_2770,N_2372,N_2174);
or U2771 (N_2771,N_2209,N_2218);
or U2772 (N_2772,N_2131,N_2364);
nand U2773 (N_2773,N_2240,N_2315);
nand U2774 (N_2774,N_2336,N_2255);
or U2775 (N_2775,N_2147,N_2347);
and U2776 (N_2776,N_2162,N_2367);
nand U2777 (N_2777,N_2357,N_2319);
nor U2778 (N_2778,N_2079,N_2362);
nor U2779 (N_2779,N_2425,N_2430);
nand U2780 (N_2780,N_2065,N_2406);
nor U2781 (N_2781,N_2121,N_2082);
nand U2782 (N_2782,N_2341,N_2049);
nand U2783 (N_2783,N_2236,N_2187);
nand U2784 (N_2784,N_2084,N_2069);
or U2785 (N_2785,N_2381,N_2313);
and U2786 (N_2786,N_2449,N_2186);
nor U2787 (N_2787,N_2053,N_2219);
or U2788 (N_2788,N_2090,N_2434);
or U2789 (N_2789,N_2182,N_2329);
xnor U2790 (N_2790,N_2236,N_2498);
xnor U2791 (N_2791,N_2273,N_2306);
nor U2792 (N_2792,N_2468,N_2013);
and U2793 (N_2793,N_2090,N_2103);
xnor U2794 (N_2794,N_2109,N_2283);
xor U2795 (N_2795,N_2427,N_2313);
xnor U2796 (N_2796,N_2109,N_2482);
or U2797 (N_2797,N_2042,N_2465);
and U2798 (N_2798,N_2362,N_2459);
nand U2799 (N_2799,N_2008,N_2376);
and U2800 (N_2800,N_2041,N_2033);
nand U2801 (N_2801,N_2410,N_2134);
and U2802 (N_2802,N_2435,N_2204);
or U2803 (N_2803,N_2064,N_2204);
nand U2804 (N_2804,N_2490,N_2333);
nor U2805 (N_2805,N_2138,N_2106);
or U2806 (N_2806,N_2259,N_2234);
and U2807 (N_2807,N_2034,N_2369);
or U2808 (N_2808,N_2007,N_2018);
nand U2809 (N_2809,N_2140,N_2223);
and U2810 (N_2810,N_2328,N_2172);
nand U2811 (N_2811,N_2175,N_2067);
xor U2812 (N_2812,N_2157,N_2266);
nand U2813 (N_2813,N_2209,N_2308);
nor U2814 (N_2814,N_2193,N_2322);
xnor U2815 (N_2815,N_2257,N_2031);
xnor U2816 (N_2816,N_2235,N_2031);
xor U2817 (N_2817,N_2071,N_2017);
nand U2818 (N_2818,N_2029,N_2206);
nand U2819 (N_2819,N_2299,N_2192);
nand U2820 (N_2820,N_2259,N_2326);
xor U2821 (N_2821,N_2253,N_2185);
or U2822 (N_2822,N_2102,N_2295);
xor U2823 (N_2823,N_2260,N_2361);
xnor U2824 (N_2824,N_2405,N_2279);
xnor U2825 (N_2825,N_2325,N_2332);
and U2826 (N_2826,N_2417,N_2198);
and U2827 (N_2827,N_2176,N_2132);
or U2828 (N_2828,N_2065,N_2121);
xor U2829 (N_2829,N_2380,N_2476);
and U2830 (N_2830,N_2298,N_2051);
and U2831 (N_2831,N_2237,N_2415);
xor U2832 (N_2832,N_2376,N_2329);
nand U2833 (N_2833,N_2232,N_2237);
and U2834 (N_2834,N_2180,N_2447);
nor U2835 (N_2835,N_2049,N_2170);
nand U2836 (N_2836,N_2034,N_2232);
or U2837 (N_2837,N_2365,N_2488);
or U2838 (N_2838,N_2124,N_2447);
and U2839 (N_2839,N_2090,N_2352);
or U2840 (N_2840,N_2473,N_2320);
and U2841 (N_2841,N_2270,N_2152);
nor U2842 (N_2842,N_2341,N_2153);
nor U2843 (N_2843,N_2204,N_2334);
and U2844 (N_2844,N_2379,N_2411);
nand U2845 (N_2845,N_2372,N_2084);
or U2846 (N_2846,N_2254,N_2193);
and U2847 (N_2847,N_2456,N_2185);
and U2848 (N_2848,N_2004,N_2245);
nand U2849 (N_2849,N_2109,N_2455);
nand U2850 (N_2850,N_2409,N_2012);
and U2851 (N_2851,N_2086,N_2087);
or U2852 (N_2852,N_2482,N_2177);
nand U2853 (N_2853,N_2298,N_2272);
nor U2854 (N_2854,N_2111,N_2257);
nand U2855 (N_2855,N_2034,N_2231);
and U2856 (N_2856,N_2294,N_2015);
xnor U2857 (N_2857,N_2147,N_2443);
or U2858 (N_2858,N_2340,N_2397);
nor U2859 (N_2859,N_2051,N_2413);
xor U2860 (N_2860,N_2439,N_2251);
xnor U2861 (N_2861,N_2443,N_2353);
nor U2862 (N_2862,N_2252,N_2477);
or U2863 (N_2863,N_2436,N_2073);
or U2864 (N_2864,N_2463,N_2236);
or U2865 (N_2865,N_2051,N_2350);
nand U2866 (N_2866,N_2397,N_2109);
and U2867 (N_2867,N_2356,N_2314);
xnor U2868 (N_2868,N_2255,N_2340);
or U2869 (N_2869,N_2222,N_2020);
and U2870 (N_2870,N_2181,N_2053);
or U2871 (N_2871,N_2384,N_2074);
xor U2872 (N_2872,N_2024,N_2416);
nand U2873 (N_2873,N_2172,N_2451);
or U2874 (N_2874,N_2302,N_2199);
and U2875 (N_2875,N_2137,N_2065);
xnor U2876 (N_2876,N_2108,N_2496);
or U2877 (N_2877,N_2301,N_2136);
xnor U2878 (N_2878,N_2093,N_2190);
xnor U2879 (N_2879,N_2307,N_2447);
or U2880 (N_2880,N_2392,N_2072);
and U2881 (N_2881,N_2196,N_2470);
nor U2882 (N_2882,N_2052,N_2305);
and U2883 (N_2883,N_2423,N_2018);
nand U2884 (N_2884,N_2475,N_2062);
nor U2885 (N_2885,N_2493,N_2229);
xor U2886 (N_2886,N_2392,N_2398);
xor U2887 (N_2887,N_2147,N_2144);
nor U2888 (N_2888,N_2296,N_2044);
nor U2889 (N_2889,N_2325,N_2133);
xnor U2890 (N_2890,N_2136,N_2407);
and U2891 (N_2891,N_2360,N_2484);
xnor U2892 (N_2892,N_2466,N_2143);
nor U2893 (N_2893,N_2128,N_2154);
and U2894 (N_2894,N_2476,N_2332);
nor U2895 (N_2895,N_2124,N_2438);
nand U2896 (N_2896,N_2262,N_2051);
xor U2897 (N_2897,N_2370,N_2477);
and U2898 (N_2898,N_2158,N_2191);
and U2899 (N_2899,N_2038,N_2227);
xnor U2900 (N_2900,N_2275,N_2000);
nand U2901 (N_2901,N_2429,N_2490);
and U2902 (N_2902,N_2259,N_2319);
and U2903 (N_2903,N_2321,N_2110);
nor U2904 (N_2904,N_2157,N_2386);
nand U2905 (N_2905,N_2244,N_2316);
or U2906 (N_2906,N_2235,N_2410);
nor U2907 (N_2907,N_2186,N_2387);
nor U2908 (N_2908,N_2458,N_2043);
xor U2909 (N_2909,N_2173,N_2459);
or U2910 (N_2910,N_2404,N_2159);
or U2911 (N_2911,N_2009,N_2385);
nand U2912 (N_2912,N_2440,N_2410);
nand U2913 (N_2913,N_2444,N_2448);
and U2914 (N_2914,N_2021,N_2430);
or U2915 (N_2915,N_2102,N_2112);
nand U2916 (N_2916,N_2200,N_2347);
nand U2917 (N_2917,N_2172,N_2281);
and U2918 (N_2918,N_2469,N_2364);
xor U2919 (N_2919,N_2455,N_2428);
nand U2920 (N_2920,N_2097,N_2298);
and U2921 (N_2921,N_2485,N_2394);
nand U2922 (N_2922,N_2075,N_2047);
or U2923 (N_2923,N_2212,N_2202);
nand U2924 (N_2924,N_2324,N_2283);
or U2925 (N_2925,N_2474,N_2050);
xor U2926 (N_2926,N_2261,N_2203);
and U2927 (N_2927,N_2059,N_2447);
xnor U2928 (N_2928,N_2046,N_2214);
nor U2929 (N_2929,N_2036,N_2326);
nand U2930 (N_2930,N_2170,N_2191);
or U2931 (N_2931,N_2250,N_2446);
nor U2932 (N_2932,N_2087,N_2262);
and U2933 (N_2933,N_2242,N_2334);
xor U2934 (N_2934,N_2165,N_2173);
nand U2935 (N_2935,N_2267,N_2422);
and U2936 (N_2936,N_2433,N_2331);
xor U2937 (N_2937,N_2316,N_2348);
and U2938 (N_2938,N_2159,N_2331);
xor U2939 (N_2939,N_2104,N_2423);
nand U2940 (N_2940,N_2190,N_2158);
xnor U2941 (N_2941,N_2093,N_2098);
xnor U2942 (N_2942,N_2360,N_2217);
nor U2943 (N_2943,N_2421,N_2448);
or U2944 (N_2944,N_2380,N_2002);
and U2945 (N_2945,N_2257,N_2107);
or U2946 (N_2946,N_2247,N_2433);
and U2947 (N_2947,N_2412,N_2489);
xnor U2948 (N_2948,N_2029,N_2002);
xor U2949 (N_2949,N_2497,N_2298);
xnor U2950 (N_2950,N_2436,N_2008);
nor U2951 (N_2951,N_2012,N_2411);
xor U2952 (N_2952,N_2274,N_2290);
nor U2953 (N_2953,N_2323,N_2157);
nor U2954 (N_2954,N_2010,N_2158);
nand U2955 (N_2955,N_2162,N_2305);
and U2956 (N_2956,N_2008,N_2428);
xnor U2957 (N_2957,N_2085,N_2447);
and U2958 (N_2958,N_2168,N_2450);
nor U2959 (N_2959,N_2427,N_2137);
or U2960 (N_2960,N_2175,N_2090);
and U2961 (N_2961,N_2401,N_2205);
nor U2962 (N_2962,N_2171,N_2236);
and U2963 (N_2963,N_2112,N_2029);
nand U2964 (N_2964,N_2193,N_2082);
or U2965 (N_2965,N_2026,N_2041);
nand U2966 (N_2966,N_2140,N_2420);
nor U2967 (N_2967,N_2085,N_2259);
nor U2968 (N_2968,N_2070,N_2144);
nand U2969 (N_2969,N_2289,N_2226);
nor U2970 (N_2970,N_2101,N_2060);
and U2971 (N_2971,N_2128,N_2392);
nor U2972 (N_2972,N_2466,N_2005);
nand U2973 (N_2973,N_2449,N_2448);
nand U2974 (N_2974,N_2302,N_2032);
and U2975 (N_2975,N_2247,N_2220);
xnor U2976 (N_2976,N_2249,N_2327);
and U2977 (N_2977,N_2414,N_2338);
nand U2978 (N_2978,N_2168,N_2369);
or U2979 (N_2979,N_2018,N_2070);
and U2980 (N_2980,N_2421,N_2018);
nor U2981 (N_2981,N_2374,N_2116);
and U2982 (N_2982,N_2458,N_2475);
and U2983 (N_2983,N_2221,N_2342);
or U2984 (N_2984,N_2198,N_2378);
nand U2985 (N_2985,N_2400,N_2485);
and U2986 (N_2986,N_2422,N_2085);
nand U2987 (N_2987,N_2286,N_2057);
and U2988 (N_2988,N_2372,N_2134);
nand U2989 (N_2989,N_2395,N_2026);
nand U2990 (N_2990,N_2205,N_2054);
xnor U2991 (N_2991,N_2372,N_2126);
xnor U2992 (N_2992,N_2019,N_2051);
and U2993 (N_2993,N_2014,N_2377);
or U2994 (N_2994,N_2017,N_2292);
nand U2995 (N_2995,N_2223,N_2379);
nand U2996 (N_2996,N_2440,N_2004);
nor U2997 (N_2997,N_2496,N_2245);
and U2998 (N_2998,N_2445,N_2397);
or U2999 (N_2999,N_2020,N_2292);
nor U3000 (N_3000,N_2544,N_2951);
xor U3001 (N_3001,N_2608,N_2871);
and U3002 (N_3002,N_2561,N_2946);
and U3003 (N_3003,N_2784,N_2598);
nor U3004 (N_3004,N_2707,N_2625);
nor U3005 (N_3005,N_2766,N_2829);
xor U3006 (N_3006,N_2510,N_2635);
and U3007 (N_3007,N_2760,N_2547);
or U3008 (N_3008,N_2789,N_2527);
and U3009 (N_3009,N_2671,N_2588);
or U3010 (N_3010,N_2810,N_2848);
xnor U3011 (N_3011,N_2888,N_2662);
xor U3012 (N_3012,N_2513,N_2713);
and U3013 (N_3013,N_2890,N_2866);
or U3014 (N_3014,N_2920,N_2870);
xnor U3015 (N_3015,N_2819,N_2834);
xnor U3016 (N_3016,N_2833,N_2661);
and U3017 (N_3017,N_2763,N_2668);
nor U3018 (N_3018,N_2591,N_2728);
or U3019 (N_3019,N_2666,N_2585);
or U3020 (N_3020,N_2553,N_2744);
nor U3021 (N_3021,N_2967,N_2646);
or U3022 (N_3022,N_2693,N_2746);
nand U3023 (N_3023,N_2658,N_2874);
xnor U3024 (N_3024,N_2803,N_2759);
or U3025 (N_3025,N_2648,N_2616);
and U3026 (N_3026,N_2783,N_2929);
nand U3027 (N_3027,N_2932,N_2719);
and U3028 (N_3028,N_2786,N_2768);
and U3029 (N_3029,N_2584,N_2808);
and U3030 (N_3030,N_2734,N_2572);
nor U3031 (N_3031,N_2762,N_2990);
nand U3032 (N_3032,N_2704,N_2835);
nand U3033 (N_3033,N_2889,N_2710);
nor U3034 (N_3034,N_2738,N_2700);
or U3035 (N_3035,N_2924,N_2897);
and U3036 (N_3036,N_2577,N_2531);
nor U3037 (N_3037,N_2907,N_2624);
nor U3038 (N_3038,N_2984,N_2583);
and U3039 (N_3039,N_2849,N_2526);
xor U3040 (N_3040,N_2747,N_2593);
nor U3041 (N_3041,N_2902,N_2670);
xor U3042 (N_3042,N_2732,N_2769);
nand U3043 (N_3043,N_2843,N_2823);
nor U3044 (N_3044,N_2511,N_2586);
and U3045 (N_3045,N_2859,N_2726);
or U3046 (N_3046,N_2963,N_2580);
or U3047 (N_3047,N_2539,N_2995);
or U3048 (N_3048,N_2607,N_2838);
xor U3049 (N_3049,N_2743,N_2611);
nand U3050 (N_3050,N_2537,N_2737);
nand U3051 (N_3051,N_2831,N_2817);
nand U3052 (N_3052,N_2623,N_2564);
xor U3053 (N_3053,N_2943,N_2718);
or U3054 (N_3054,N_2745,N_2649);
and U3055 (N_3055,N_2642,N_2968);
or U3056 (N_3056,N_2589,N_2679);
or U3057 (N_3057,N_2617,N_2676);
or U3058 (N_3058,N_2560,N_2566);
xor U3059 (N_3059,N_2742,N_2647);
nand U3060 (N_3060,N_2702,N_2581);
and U3061 (N_3061,N_2785,N_2660);
or U3062 (N_3062,N_2881,N_2931);
nand U3063 (N_3063,N_2797,N_2650);
or U3064 (N_3064,N_2520,N_2555);
nor U3065 (N_3065,N_2590,N_2796);
and U3066 (N_3066,N_2896,N_2621);
nand U3067 (N_3067,N_2892,N_2721);
or U3068 (N_3068,N_2692,N_2651);
or U3069 (N_3069,N_2592,N_2986);
or U3070 (N_3070,N_2543,N_2514);
nor U3071 (N_3071,N_2872,N_2684);
and U3072 (N_3072,N_2916,N_2836);
nand U3073 (N_3073,N_2614,N_2893);
and U3074 (N_3074,N_2842,N_2901);
xnor U3075 (N_3075,N_2534,N_2776);
nand U3076 (N_3076,N_2716,N_2518);
xor U3077 (N_3077,N_2756,N_2998);
xor U3078 (N_3078,N_2636,N_2554);
nand U3079 (N_3079,N_2765,N_2965);
or U3080 (N_3080,N_2500,N_2694);
or U3081 (N_3081,N_2864,N_2612);
nand U3082 (N_3082,N_2613,N_2550);
and U3083 (N_3083,N_2825,N_2939);
and U3084 (N_3084,N_2813,N_2996);
nor U3085 (N_3085,N_2805,N_2643);
xor U3086 (N_3086,N_2877,N_2695);
nor U3087 (N_3087,N_2599,N_2926);
xnor U3088 (N_3088,N_2685,N_2578);
nand U3089 (N_3089,N_2771,N_2711);
and U3090 (N_3090,N_2895,N_2894);
nand U3091 (N_3091,N_2565,N_2787);
and U3092 (N_3092,N_2962,N_2712);
xor U3093 (N_3093,N_2778,N_2818);
xnor U3094 (N_3094,N_2683,N_2837);
nand U3095 (N_3095,N_2677,N_2610);
and U3096 (N_3096,N_2626,N_2714);
or U3097 (N_3097,N_2654,N_2521);
nand U3098 (N_3098,N_2910,N_2921);
nand U3099 (N_3099,N_2930,N_2958);
and U3100 (N_3100,N_2873,N_2727);
nor U3101 (N_3101,N_2657,N_2854);
nor U3102 (N_3102,N_2972,N_2964);
and U3103 (N_3103,N_2826,N_2976);
or U3104 (N_3104,N_2594,N_2655);
nor U3105 (N_3105,N_2780,N_2731);
nor U3106 (N_3106,N_2729,N_2563);
xnor U3107 (N_3107,N_2876,N_2529);
nand U3108 (N_3108,N_2980,N_2767);
or U3109 (N_3109,N_2629,N_2507);
xnor U3110 (N_3110,N_2945,N_2820);
nand U3111 (N_3111,N_2503,N_2758);
nand U3112 (N_3112,N_2698,N_2772);
or U3113 (N_3113,N_2755,N_2687);
or U3114 (N_3114,N_2740,N_2750);
or U3115 (N_3115,N_2664,N_2573);
or U3116 (N_3116,N_2937,N_2627);
or U3117 (N_3117,N_2991,N_2858);
nor U3118 (N_3118,N_2891,N_2523);
nor U3119 (N_3119,N_2541,N_2706);
and U3120 (N_3120,N_2900,N_2882);
nor U3121 (N_3121,N_2999,N_2663);
nand U3122 (N_3122,N_2824,N_2802);
nor U3123 (N_3123,N_2639,N_2909);
nand U3124 (N_3124,N_2691,N_2528);
nor U3125 (N_3125,N_2569,N_2556);
and U3126 (N_3126,N_2770,N_2791);
and U3127 (N_3127,N_2987,N_2512);
and U3128 (N_3128,N_2798,N_2733);
or U3129 (N_3129,N_2782,N_2839);
or U3130 (N_3130,N_2505,N_2886);
or U3131 (N_3131,N_2928,N_2799);
nand U3132 (N_3132,N_2730,N_2530);
nor U3133 (N_3133,N_2884,N_2705);
xor U3134 (N_3134,N_2978,N_2868);
nor U3135 (N_3135,N_2801,N_2804);
or U3136 (N_3136,N_2501,N_2525);
xnor U3137 (N_3137,N_2832,N_2757);
nor U3138 (N_3138,N_2552,N_2508);
or U3139 (N_3139,N_2741,N_2788);
xor U3140 (N_3140,N_2988,N_2997);
or U3141 (N_3141,N_2950,N_2955);
nand U3142 (N_3142,N_2828,N_2830);
and U3143 (N_3143,N_2630,N_2725);
xor U3144 (N_3144,N_2615,N_2689);
nand U3145 (N_3145,N_2722,N_2792);
and U3146 (N_3146,N_2618,N_2956);
nand U3147 (N_3147,N_2574,N_2779);
and U3148 (N_3148,N_2532,N_2923);
nand U3149 (N_3149,N_2863,N_2622);
nor U3150 (N_3150,N_2867,N_2596);
or U3151 (N_3151,N_2811,N_2781);
nand U3152 (N_3152,N_2977,N_2715);
or U3153 (N_3153,N_2952,N_2665);
or U3154 (N_3154,N_2517,N_2678);
nor U3155 (N_3155,N_2961,N_2903);
or U3156 (N_3156,N_2800,N_2860);
or U3157 (N_3157,N_2632,N_2761);
or U3158 (N_3158,N_2869,N_2675);
or U3159 (N_3159,N_2949,N_2970);
xor U3160 (N_3160,N_2673,N_2680);
xor U3161 (N_3161,N_2724,N_2948);
and U3162 (N_3162,N_2773,N_2681);
or U3163 (N_3163,N_2709,N_2807);
nor U3164 (N_3164,N_2855,N_2793);
or U3165 (N_3165,N_2703,N_2570);
or U3166 (N_3166,N_2653,N_2736);
or U3167 (N_3167,N_2915,N_2857);
or U3168 (N_3168,N_2620,N_2571);
xor U3169 (N_3169,N_2749,N_2506);
and U3170 (N_3170,N_2812,N_2919);
xnor U3171 (N_3171,N_2887,N_2899);
nand U3172 (N_3172,N_2845,N_2821);
or U3173 (N_3173,N_2602,N_2953);
xor U3174 (N_3174,N_2861,N_2925);
or U3175 (N_3175,N_2682,N_2753);
and U3176 (N_3176,N_2519,N_2809);
nor U3177 (N_3177,N_2669,N_2908);
nor U3178 (N_3178,N_2633,N_2790);
and U3179 (N_3179,N_2595,N_2806);
nand U3180 (N_3180,N_2548,N_2981);
nor U3181 (N_3181,N_2672,N_2739);
xor U3182 (N_3182,N_2558,N_2989);
xor U3183 (N_3183,N_2912,N_2960);
or U3184 (N_3184,N_2542,N_2880);
nor U3185 (N_3185,N_2841,N_2827);
and U3186 (N_3186,N_2536,N_2904);
and U3187 (N_3187,N_2852,N_2674);
or U3188 (N_3188,N_2582,N_2540);
or U3189 (N_3189,N_2862,N_2559);
nor U3190 (N_3190,N_2774,N_2814);
and U3191 (N_3191,N_2688,N_2992);
nand U3192 (N_3192,N_2579,N_2856);
and U3193 (N_3193,N_2878,N_2644);
nand U3194 (N_3194,N_2522,N_2993);
and U3195 (N_3195,N_2640,N_2546);
or U3196 (N_3196,N_2538,N_2516);
xnor U3197 (N_3197,N_2701,N_2597);
and U3198 (N_3198,N_2603,N_2969);
or U3199 (N_3199,N_2557,N_2922);
or U3200 (N_3200,N_2562,N_2697);
nand U3201 (N_3201,N_2606,N_2935);
xor U3202 (N_3202,N_2587,N_2605);
and U3203 (N_3203,N_2905,N_2634);
nor U3204 (N_3204,N_2975,N_2652);
xor U3205 (N_3205,N_2944,N_2794);
and U3206 (N_3206,N_2940,N_2656);
or U3207 (N_3207,N_2934,N_2567);
nor U3208 (N_3208,N_2840,N_2917);
xnor U3209 (N_3209,N_2690,N_2515);
and U3210 (N_3210,N_2979,N_2601);
nand U3211 (N_3211,N_2954,N_2875);
nor U3212 (N_3212,N_2883,N_2748);
or U3213 (N_3213,N_2957,N_2509);
or U3214 (N_3214,N_2846,N_2966);
xor U3215 (N_3215,N_2898,N_2973);
nor U3216 (N_3216,N_2913,N_2775);
and U3217 (N_3217,N_2502,N_2631);
and U3218 (N_3218,N_2822,N_2600);
nor U3219 (N_3219,N_2764,N_2942);
nand U3220 (N_3220,N_2777,N_2959);
xor U3221 (N_3221,N_2645,N_2974);
and U3222 (N_3222,N_2851,N_2971);
nand U3223 (N_3223,N_2752,N_2568);
nor U3224 (N_3224,N_2815,N_2847);
xor U3225 (N_3225,N_2850,N_2735);
nand U3226 (N_3226,N_2816,N_2885);
nand U3227 (N_3227,N_2696,N_2938);
nand U3228 (N_3228,N_2933,N_2524);
xnor U3229 (N_3229,N_2754,N_2911);
nor U3230 (N_3230,N_2637,N_2985);
or U3231 (N_3231,N_2879,N_2699);
xnor U3232 (N_3232,N_2906,N_2504);
or U3233 (N_3233,N_2723,N_2641);
and U3234 (N_3234,N_2918,N_2576);
xor U3235 (N_3235,N_2983,N_2609);
xnor U3236 (N_3236,N_2720,N_2936);
nor U3237 (N_3237,N_2751,N_2853);
nand U3238 (N_3238,N_2686,N_2994);
and U3239 (N_3239,N_2551,N_2575);
and U3240 (N_3240,N_2604,N_2982);
or U3241 (N_3241,N_2535,N_2533);
nor U3242 (N_3242,N_2708,N_2865);
nor U3243 (N_3243,N_2941,N_2545);
and U3244 (N_3244,N_2667,N_2914);
and U3245 (N_3245,N_2638,N_2927);
nor U3246 (N_3246,N_2844,N_2628);
and U3247 (N_3247,N_2659,N_2947);
xor U3248 (N_3248,N_2717,N_2549);
and U3249 (N_3249,N_2619,N_2795);
nand U3250 (N_3250,N_2758,N_2863);
xnor U3251 (N_3251,N_2752,N_2956);
nor U3252 (N_3252,N_2766,N_2945);
or U3253 (N_3253,N_2520,N_2885);
xnor U3254 (N_3254,N_2794,N_2687);
or U3255 (N_3255,N_2816,N_2845);
nand U3256 (N_3256,N_2817,N_2999);
nand U3257 (N_3257,N_2957,N_2976);
xor U3258 (N_3258,N_2905,N_2577);
or U3259 (N_3259,N_2942,N_2795);
or U3260 (N_3260,N_2975,N_2519);
or U3261 (N_3261,N_2799,N_2511);
nand U3262 (N_3262,N_2783,N_2508);
or U3263 (N_3263,N_2892,N_2641);
nor U3264 (N_3264,N_2761,N_2857);
nor U3265 (N_3265,N_2822,N_2536);
xor U3266 (N_3266,N_2936,N_2517);
nor U3267 (N_3267,N_2871,N_2629);
or U3268 (N_3268,N_2532,N_2571);
and U3269 (N_3269,N_2634,N_2778);
or U3270 (N_3270,N_2575,N_2838);
nand U3271 (N_3271,N_2933,N_2993);
nor U3272 (N_3272,N_2558,N_2797);
and U3273 (N_3273,N_2827,N_2646);
or U3274 (N_3274,N_2681,N_2882);
nand U3275 (N_3275,N_2835,N_2511);
and U3276 (N_3276,N_2731,N_2665);
nor U3277 (N_3277,N_2648,N_2842);
nor U3278 (N_3278,N_2672,N_2654);
xnor U3279 (N_3279,N_2747,N_2862);
xnor U3280 (N_3280,N_2911,N_2631);
or U3281 (N_3281,N_2521,N_2804);
nand U3282 (N_3282,N_2985,N_2524);
nand U3283 (N_3283,N_2731,N_2603);
nand U3284 (N_3284,N_2821,N_2689);
nand U3285 (N_3285,N_2639,N_2728);
nor U3286 (N_3286,N_2837,N_2786);
xor U3287 (N_3287,N_2780,N_2509);
xnor U3288 (N_3288,N_2540,N_2939);
xor U3289 (N_3289,N_2925,N_2505);
nand U3290 (N_3290,N_2657,N_2946);
nor U3291 (N_3291,N_2539,N_2602);
nor U3292 (N_3292,N_2809,N_2985);
xor U3293 (N_3293,N_2541,N_2639);
and U3294 (N_3294,N_2986,N_2674);
or U3295 (N_3295,N_2606,N_2841);
or U3296 (N_3296,N_2814,N_2955);
nand U3297 (N_3297,N_2500,N_2606);
nor U3298 (N_3298,N_2873,N_2868);
or U3299 (N_3299,N_2806,N_2884);
nand U3300 (N_3300,N_2854,N_2947);
and U3301 (N_3301,N_2716,N_2757);
xnor U3302 (N_3302,N_2676,N_2662);
and U3303 (N_3303,N_2898,N_2760);
or U3304 (N_3304,N_2603,N_2932);
and U3305 (N_3305,N_2738,N_2525);
or U3306 (N_3306,N_2520,N_2625);
xnor U3307 (N_3307,N_2843,N_2732);
nand U3308 (N_3308,N_2583,N_2987);
xnor U3309 (N_3309,N_2948,N_2646);
nand U3310 (N_3310,N_2506,N_2958);
nor U3311 (N_3311,N_2790,N_2974);
and U3312 (N_3312,N_2877,N_2999);
and U3313 (N_3313,N_2511,N_2839);
or U3314 (N_3314,N_2761,N_2594);
nor U3315 (N_3315,N_2660,N_2898);
xor U3316 (N_3316,N_2750,N_2927);
or U3317 (N_3317,N_2668,N_2823);
xnor U3318 (N_3318,N_2664,N_2524);
and U3319 (N_3319,N_2738,N_2982);
nand U3320 (N_3320,N_2942,N_2558);
nor U3321 (N_3321,N_2819,N_2896);
or U3322 (N_3322,N_2567,N_2748);
or U3323 (N_3323,N_2621,N_2893);
or U3324 (N_3324,N_2775,N_2694);
nor U3325 (N_3325,N_2797,N_2774);
and U3326 (N_3326,N_2832,N_2581);
nand U3327 (N_3327,N_2580,N_2623);
nor U3328 (N_3328,N_2979,N_2999);
xnor U3329 (N_3329,N_2774,N_2744);
or U3330 (N_3330,N_2909,N_2823);
xnor U3331 (N_3331,N_2603,N_2951);
nor U3332 (N_3332,N_2545,N_2886);
and U3333 (N_3333,N_2980,N_2862);
nand U3334 (N_3334,N_2586,N_2767);
nand U3335 (N_3335,N_2755,N_2838);
and U3336 (N_3336,N_2898,N_2810);
or U3337 (N_3337,N_2529,N_2541);
xor U3338 (N_3338,N_2892,N_2624);
xor U3339 (N_3339,N_2811,N_2759);
nor U3340 (N_3340,N_2647,N_2864);
nand U3341 (N_3341,N_2509,N_2854);
or U3342 (N_3342,N_2531,N_2511);
and U3343 (N_3343,N_2554,N_2632);
nor U3344 (N_3344,N_2541,N_2596);
nand U3345 (N_3345,N_2553,N_2752);
nand U3346 (N_3346,N_2675,N_2764);
and U3347 (N_3347,N_2517,N_2731);
nor U3348 (N_3348,N_2627,N_2906);
and U3349 (N_3349,N_2549,N_2612);
nand U3350 (N_3350,N_2666,N_2795);
xor U3351 (N_3351,N_2964,N_2955);
and U3352 (N_3352,N_2840,N_2906);
nand U3353 (N_3353,N_2596,N_2986);
nor U3354 (N_3354,N_2891,N_2619);
nor U3355 (N_3355,N_2890,N_2901);
nor U3356 (N_3356,N_2617,N_2587);
nor U3357 (N_3357,N_2704,N_2681);
or U3358 (N_3358,N_2701,N_2818);
nor U3359 (N_3359,N_2602,N_2771);
xor U3360 (N_3360,N_2823,N_2875);
and U3361 (N_3361,N_2715,N_2609);
or U3362 (N_3362,N_2977,N_2973);
xnor U3363 (N_3363,N_2638,N_2659);
or U3364 (N_3364,N_2764,N_2548);
xor U3365 (N_3365,N_2771,N_2605);
nor U3366 (N_3366,N_2901,N_2597);
nand U3367 (N_3367,N_2801,N_2844);
xor U3368 (N_3368,N_2726,N_2614);
nand U3369 (N_3369,N_2711,N_2560);
nand U3370 (N_3370,N_2878,N_2653);
nand U3371 (N_3371,N_2669,N_2873);
nor U3372 (N_3372,N_2718,N_2555);
nor U3373 (N_3373,N_2887,N_2650);
or U3374 (N_3374,N_2672,N_2952);
and U3375 (N_3375,N_2540,N_2885);
and U3376 (N_3376,N_2627,N_2616);
xor U3377 (N_3377,N_2796,N_2720);
xor U3378 (N_3378,N_2742,N_2555);
nand U3379 (N_3379,N_2525,N_2636);
nor U3380 (N_3380,N_2632,N_2572);
nand U3381 (N_3381,N_2701,N_2879);
nand U3382 (N_3382,N_2554,N_2899);
nor U3383 (N_3383,N_2838,N_2673);
nand U3384 (N_3384,N_2555,N_2777);
xor U3385 (N_3385,N_2905,N_2857);
or U3386 (N_3386,N_2768,N_2763);
nor U3387 (N_3387,N_2918,N_2601);
nand U3388 (N_3388,N_2959,N_2976);
and U3389 (N_3389,N_2538,N_2918);
xnor U3390 (N_3390,N_2880,N_2611);
nand U3391 (N_3391,N_2665,N_2991);
nand U3392 (N_3392,N_2743,N_2577);
or U3393 (N_3393,N_2583,N_2794);
nand U3394 (N_3394,N_2607,N_2956);
xor U3395 (N_3395,N_2918,N_2713);
and U3396 (N_3396,N_2808,N_2514);
and U3397 (N_3397,N_2504,N_2591);
or U3398 (N_3398,N_2822,N_2724);
nand U3399 (N_3399,N_2986,N_2976);
xnor U3400 (N_3400,N_2634,N_2718);
nand U3401 (N_3401,N_2656,N_2631);
or U3402 (N_3402,N_2874,N_2848);
and U3403 (N_3403,N_2982,N_2813);
xnor U3404 (N_3404,N_2655,N_2855);
nand U3405 (N_3405,N_2977,N_2955);
nand U3406 (N_3406,N_2508,N_2737);
nand U3407 (N_3407,N_2653,N_2709);
xnor U3408 (N_3408,N_2745,N_2914);
and U3409 (N_3409,N_2731,N_2921);
and U3410 (N_3410,N_2863,N_2955);
nand U3411 (N_3411,N_2850,N_2941);
xnor U3412 (N_3412,N_2904,N_2663);
xnor U3413 (N_3413,N_2892,N_2608);
xor U3414 (N_3414,N_2948,N_2916);
nor U3415 (N_3415,N_2505,N_2675);
nor U3416 (N_3416,N_2871,N_2978);
and U3417 (N_3417,N_2816,N_2767);
nand U3418 (N_3418,N_2782,N_2716);
nand U3419 (N_3419,N_2563,N_2516);
nor U3420 (N_3420,N_2752,N_2740);
xnor U3421 (N_3421,N_2914,N_2861);
and U3422 (N_3422,N_2550,N_2532);
nor U3423 (N_3423,N_2757,N_2635);
nand U3424 (N_3424,N_2930,N_2935);
nand U3425 (N_3425,N_2665,N_2928);
and U3426 (N_3426,N_2509,N_2989);
and U3427 (N_3427,N_2734,N_2936);
nand U3428 (N_3428,N_2841,N_2805);
xor U3429 (N_3429,N_2982,N_2767);
and U3430 (N_3430,N_2921,N_2654);
xnor U3431 (N_3431,N_2935,N_2988);
xor U3432 (N_3432,N_2874,N_2732);
and U3433 (N_3433,N_2968,N_2581);
or U3434 (N_3434,N_2974,N_2760);
and U3435 (N_3435,N_2527,N_2893);
nor U3436 (N_3436,N_2753,N_2717);
nor U3437 (N_3437,N_2776,N_2927);
nor U3438 (N_3438,N_2810,N_2501);
nor U3439 (N_3439,N_2900,N_2868);
or U3440 (N_3440,N_2770,N_2912);
xnor U3441 (N_3441,N_2526,N_2965);
xnor U3442 (N_3442,N_2670,N_2775);
nand U3443 (N_3443,N_2741,N_2555);
nand U3444 (N_3444,N_2524,N_2510);
nand U3445 (N_3445,N_2953,N_2874);
nor U3446 (N_3446,N_2885,N_2513);
nand U3447 (N_3447,N_2932,N_2514);
and U3448 (N_3448,N_2653,N_2977);
nand U3449 (N_3449,N_2931,N_2814);
xnor U3450 (N_3450,N_2921,N_2744);
nand U3451 (N_3451,N_2893,N_2926);
or U3452 (N_3452,N_2616,N_2678);
xor U3453 (N_3453,N_2527,N_2961);
xnor U3454 (N_3454,N_2901,N_2504);
or U3455 (N_3455,N_2526,N_2827);
and U3456 (N_3456,N_2997,N_2535);
nor U3457 (N_3457,N_2810,N_2967);
and U3458 (N_3458,N_2783,N_2685);
and U3459 (N_3459,N_2827,N_2623);
nand U3460 (N_3460,N_2768,N_2950);
nor U3461 (N_3461,N_2534,N_2786);
and U3462 (N_3462,N_2649,N_2582);
nor U3463 (N_3463,N_2984,N_2786);
nand U3464 (N_3464,N_2932,N_2702);
or U3465 (N_3465,N_2551,N_2589);
or U3466 (N_3466,N_2934,N_2546);
nand U3467 (N_3467,N_2855,N_2813);
nand U3468 (N_3468,N_2911,N_2860);
nand U3469 (N_3469,N_2831,N_2743);
xnor U3470 (N_3470,N_2750,N_2973);
or U3471 (N_3471,N_2544,N_2518);
and U3472 (N_3472,N_2980,N_2960);
nor U3473 (N_3473,N_2908,N_2574);
nor U3474 (N_3474,N_2831,N_2663);
and U3475 (N_3475,N_2879,N_2963);
nor U3476 (N_3476,N_2765,N_2503);
or U3477 (N_3477,N_2869,N_2682);
nor U3478 (N_3478,N_2936,N_2553);
and U3479 (N_3479,N_2798,N_2806);
or U3480 (N_3480,N_2509,N_2670);
and U3481 (N_3481,N_2753,N_2812);
xnor U3482 (N_3482,N_2944,N_2533);
nand U3483 (N_3483,N_2919,N_2601);
or U3484 (N_3484,N_2512,N_2867);
and U3485 (N_3485,N_2945,N_2869);
nor U3486 (N_3486,N_2989,N_2993);
xor U3487 (N_3487,N_2859,N_2607);
nand U3488 (N_3488,N_2681,N_2727);
and U3489 (N_3489,N_2804,N_2762);
or U3490 (N_3490,N_2500,N_2982);
xor U3491 (N_3491,N_2683,N_2859);
xnor U3492 (N_3492,N_2765,N_2925);
and U3493 (N_3493,N_2891,N_2846);
xnor U3494 (N_3494,N_2522,N_2844);
or U3495 (N_3495,N_2828,N_2988);
xor U3496 (N_3496,N_2503,N_2598);
or U3497 (N_3497,N_2614,N_2730);
and U3498 (N_3498,N_2585,N_2673);
or U3499 (N_3499,N_2501,N_2923);
and U3500 (N_3500,N_3174,N_3097);
nand U3501 (N_3501,N_3326,N_3144);
and U3502 (N_3502,N_3386,N_3225);
and U3503 (N_3503,N_3441,N_3093);
or U3504 (N_3504,N_3087,N_3085);
or U3505 (N_3505,N_3195,N_3179);
and U3506 (N_3506,N_3199,N_3285);
and U3507 (N_3507,N_3076,N_3170);
and U3508 (N_3508,N_3313,N_3283);
nand U3509 (N_3509,N_3395,N_3086);
nor U3510 (N_3510,N_3230,N_3111);
or U3511 (N_3511,N_3425,N_3426);
xnor U3512 (N_3512,N_3487,N_3122);
or U3513 (N_3513,N_3456,N_3279);
nor U3514 (N_3514,N_3020,N_3129);
nor U3515 (N_3515,N_3255,N_3193);
nor U3516 (N_3516,N_3067,N_3183);
and U3517 (N_3517,N_3489,N_3294);
nand U3518 (N_3518,N_3480,N_3379);
xor U3519 (N_3519,N_3246,N_3051);
nor U3520 (N_3520,N_3130,N_3491);
and U3521 (N_3521,N_3013,N_3330);
or U3522 (N_3522,N_3413,N_3100);
or U3523 (N_3523,N_3341,N_3258);
nor U3524 (N_3524,N_3420,N_3103);
xnor U3525 (N_3525,N_3431,N_3479);
nor U3526 (N_3526,N_3264,N_3143);
nor U3527 (N_3527,N_3102,N_3347);
and U3528 (N_3528,N_3339,N_3240);
nor U3529 (N_3529,N_3252,N_3113);
nor U3530 (N_3530,N_3344,N_3437);
xor U3531 (N_3531,N_3007,N_3375);
and U3532 (N_3532,N_3406,N_3371);
and U3533 (N_3533,N_3167,N_3383);
or U3534 (N_3534,N_3254,N_3433);
and U3535 (N_3535,N_3467,N_3042);
or U3536 (N_3536,N_3135,N_3238);
nor U3537 (N_3537,N_3072,N_3354);
nand U3538 (N_3538,N_3182,N_3320);
or U3539 (N_3539,N_3412,N_3319);
or U3540 (N_3540,N_3465,N_3005);
and U3541 (N_3541,N_3378,N_3069);
or U3542 (N_3542,N_3400,N_3328);
nor U3543 (N_3543,N_3058,N_3391);
nand U3544 (N_3544,N_3117,N_3212);
and U3545 (N_3545,N_3178,N_3409);
nand U3546 (N_3546,N_3359,N_3215);
or U3547 (N_3547,N_3162,N_3003);
or U3548 (N_3548,N_3171,N_3098);
or U3549 (N_3549,N_3209,N_3316);
xnor U3550 (N_3550,N_3343,N_3028);
and U3551 (N_3551,N_3234,N_3188);
nand U3552 (N_3552,N_3452,N_3435);
and U3553 (N_3553,N_3457,N_3424);
and U3554 (N_3554,N_3150,N_3271);
xor U3555 (N_3555,N_3082,N_3021);
nor U3556 (N_3556,N_3159,N_3389);
or U3557 (N_3557,N_3318,N_3314);
nand U3558 (N_3558,N_3396,N_3468);
xnor U3559 (N_3559,N_3049,N_3439);
or U3560 (N_3560,N_3398,N_3154);
xor U3561 (N_3561,N_3068,N_3127);
nor U3562 (N_3562,N_3408,N_3251);
nor U3563 (N_3563,N_3044,N_3047);
and U3564 (N_3564,N_3293,N_3486);
nand U3565 (N_3565,N_3229,N_3147);
and U3566 (N_3566,N_3145,N_3104);
or U3567 (N_3567,N_3036,N_3187);
nand U3568 (N_3568,N_3088,N_3181);
nand U3569 (N_3569,N_3261,N_3108);
nor U3570 (N_3570,N_3197,N_3027);
nor U3571 (N_3571,N_3284,N_3393);
xor U3572 (N_3572,N_3454,N_3288);
and U3573 (N_3573,N_3334,N_3474);
or U3574 (N_3574,N_3473,N_3357);
and U3575 (N_3575,N_3053,N_3163);
nor U3576 (N_3576,N_3125,N_3031);
and U3577 (N_3577,N_3185,N_3245);
nand U3578 (N_3578,N_3213,N_3046);
or U3579 (N_3579,N_3311,N_3161);
nand U3580 (N_3580,N_3388,N_3118);
and U3581 (N_3581,N_3340,N_3338);
and U3582 (N_3582,N_3050,N_3410);
nor U3583 (N_3583,N_3430,N_3206);
and U3584 (N_3584,N_3296,N_3180);
or U3585 (N_3585,N_3372,N_3038);
and U3586 (N_3586,N_3352,N_3349);
nor U3587 (N_3587,N_3366,N_3089);
or U3588 (N_3588,N_3052,N_3432);
nand U3589 (N_3589,N_3169,N_3029);
and U3590 (N_3590,N_3418,N_3221);
or U3591 (N_3591,N_3224,N_3061);
nor U3592 (N_3592,N_3115,N_3201);
nand U3593 (N_3593,N_3353,N_3403);
and U3594 (N_3594,N_3011,N_3493);
nor U3595 (N_3595,N_3325,N_3401);
nand U3596 (N_3596,N_3110,N_3070);
and U3597 (N_3597,N_3004,N_3222);
or U3598 (N_3598,N_3034,N_3263);
nor U3599 (N_3599,N_3377,N_3048);
nand U3600 (N_3600,N_3290,N_3278);
or U3601 (N_3601,N_3250,N_3176);
and U3602 (N_3602,N_3131,N_3191);
or U3603 (N_3603,N_3405,N_3152);
or U3604 (N_3604,N_3309,N_3404);
or U3605 (N_3605,N_3270,N_3281);
xor U3606 (N_3606,N_3024,N_3080);
and U3607 (N_3607,N_3422,N_3399);
xor U3608 (N_3608,N_3275,N_3297);
xor U3609 (N_3609,N_3112,N_3464);
and U3610 (N_3610,N_3351,N_3119);
nand U3611 (N_3611,N_3146,N_3350);
or U3612 (N_3612,N_3241,N_3063);
or U3613 (N_3613,N_3466,N_3440);
xnor U3614 (N_3614,N_3387,N_3345);
nand U3615 (N_3615,N_3329,N_3062);
nor U3616 (N_3616,N_3210,N_3177);
nor U3617 (N_3617,N_3227,N_3476);
nand U3618 (N_3618,N_3190,N_3078);
or U3619 (N_3619,N_3358,N_3216);
xor U3620 (N_3620,N_3262,N_3196);
nor U3621 (N_3621,N_3233,N_3189);
and U3622 (N_3622,N_3211,N_3026);
or U3623 (N_3623,N_3172,N_3443);
or U3624 (N_3624,N_3370,N_3120);
and U3625 (N_3625,N_3337,N_3256);
nand U3626 (N_3626,N_3090,N_3018);
or U3627 (N_3627,N_3166,N_3333);
or U3628 (N_3628,N_3360,N_3304);
and U3629 (N_3629,N_3203,N_3324);
or U3630 (N_3630,N_3390,N_3267);
nand U3631 (N_3631,N_3123,N_3362);
nor U3632 (N_3632,N_3280,N_3132);
or U3633 (N_3633,N_3308,N_3105);
xnor U3634 (N_3634,N_3484,N_3242);
or U3635 (N_3635,N_3427,N_3429);
or U3636 (N_3636,N_3461,N_3156);
nor U3637 (N_3637,N_3081,N_3083);
nor U3638 (N_3638,N_3361,N_3015);
nor U3639 (N_3639,N_3434,N_3327);
and U3640 (N_3640,N_3499,N_3355);
nor U3641 (N_3641,N_3009,N_3248);
and U3642 (N_3642,N_3107,N_3019);
xnor U3643 (N_3643,N_3186,N_3202);
nor U3644 (N_3644,N_3016,N_3470);
and U3645 (N_3645,N_3236,N_3217);
xor U3646 (N_3646,N_3367,N_3269);
xor U3647 (N_3647,N_3055,N_3315);
nand U3648 (N_3648,N_3376,N_3247);
or U3649 (N_3649,N_3444,N_3368);
nor U3650 (N_3650,N_3200,N_3272);
nand U3651 (N_3651,N_3471,N_3045);
and U3652 (N_3652,N_3385,N_3092);
or U3653 (N_3653,N_3000,N_3207);
nand U3654 (N_3654,N_3079,N_3266);
nor U3655 (N_3655,N_3475,N_3300);
and U3656 (N_3656,N_3126,N_3498);
or U3657 (N_3657,N_3239,N_3419);
and U3658 (N_3658,N_3134,N_3151);
and U3659 (N_3659,N_3402,N_3459);
or U3660 (N_3660,N_3001,N_3095);
xor U3661 (N_3661,N_3446,N_3023);
or U3662 (N_3662,N_3084,N_3198);
nor U3663 (N_3663,N_3346,N_3482);
xor U3664 (N_3664,N_3056,N_3039);
and U3665 (N_3665,N_3157,N_3160);
or U3666 (N_3666,N_3260,N_3133);
nand U3667 (N_3667,N_3356,N_3164);
or U3668 (N_3668,N_3137,N_3116);
or U3669 (N_3669,N_3175,N_3253);
nor U3670 (N_3670,N_3397,N_3173);
nor U3671 (N_3671,N_3394,N_3244);
nand U3672 (N_3672,N_3421,N_3043);
xor U3673 (N_3673,N_3014,N_3249);
xor U3674 (N_3674,N_3073,N_3373);
xnor U3675 (N_3675,N_3060,N_3041);
and U3676 (N_3676,N_3306,N_3295);
or U3677 (N_3677,N_3381,N_3449);
or U3678 (N_3678,N_3428,N_3292);
and U3679 (N_3679,N_3040,N_3037);
nor U3680 (N_3680,N_3148,N_3149);
nand U3681 (N_3681,N_3231,N_3168);
and U3682 (N_3682,N_3192,N_3074);
or U3683 (N_3683,N_3477,N_3305);
nand U3684 (N_3684,N_3106,N_3139);
xor U3685 (N_3685,N_3226,N_3322);
xnor U3686 (N_3686,N_3423,N_3075);
nor U3687 (N_3687,N_3382,N_3455);
xnor U3688 (N_3688,N_3492,N_3331);
and U3689 (N_3689,N_3463,N_3483);
or U3690 (N_3690,N_3287,N_3298);
nor U3691 (N_3691,N_3059,N_3458);
nand U3692 (N_3692,N_3128,N_3495);
or U3693 (N_3693,N_3485,N_3342);
or U3694 (N_3694,N_3416,N_3008);
nor U3695 (N_3695,N_3140,N_3099);
nor U3696 (N_3696,N_3469,N_3310);
nor U3697 (N_3697,N_3243,N_3235);
or U3698 (N_3698,N_3438,N_3364);
and U3699 (N_3699,N_3096,N_3054);
and U3700 (N_3700,N_3274,N_3017);
nor U3701 (N_3701,N_3276,N_3460);
nand U3702 (N_3702,N_3323,N_3436);
nand U3703 (N_3703,N_3277,N_3445);
or U3704 (N_3704,N_3321,N_3204);
nand U3705 (N_3705,N_3155,N_3035);
nand U3706 (N_3706,N_3265,N_3348);
and U3707 (N_3707,N_3153,N_3442);
xnor U3708 (N_3708,N_3417,N_3286);
xor U3709 (N_3709,N_3257,N_3071);
or U3710 (N_3710,N_3494,N_3374);
or U3711 (N_3711,N_3121,N_3448);
nor U3712 (N_3712,N_3065,N_3335);
xor U3713 (N_3713,N_3138,N_3312);
nand U3714 (N_3714,N_3273,N_3223);
and U3715 (N_3715,N_3488,N_3218);
nand U3716 (N_3716,N_3481,N_3077);
nor U3717 (N_3717,N_3259,N_3317);
nor U3718 (N_3718,N_3025,N_3232);
xnor U3719 (N_3719,N_3064,N_3136);
nand U3720 (N_3720,N_3496,N_3291);
or U3721 (N_3721,N_3141,N_3006);
nor U3722 (N_3722,N_3109,N_3497);
or U3723 (N_3723,N_3332,N_3392);
nor U3724 (N_3724,N_3010,N_3462);
and U3725 (N_3725,N_3237,N_3214);
xor U3726 (N_3726,N_3472,N_3478);
or U3727 (N_3727,N_3384,N_3184);
nand U3728 (N_3728,N_3453,N_3301);
nor U3729 (N_3729,N_3208,N_3032);
nand U3730 (N_3730,N_3158,N_3094);
nand U3731 (N_3731,N_3369,N_3033);
nor U3732 (N_3732,N_3002,N_3407);
nand U3733 (N_3733,N_3091,N_3336);
xnor U3734 (N_3734,N_3268,N_3282);
and U3735 (N_3735,N_3365,N_3414);
or U3736 (N_3736,N_3219,N_3030);
nand U3737 (N_3737,N_3415,N_3165);
nor U3738 (N_3738,N_3022,N_3057);
nor U3739 (N_3739,N_3114,N_3101);
xnor U3740 (N_3740,N_3142,N_3451);
xor U3741 (N_3741,N_3012,N_3490);
nor U3742 (N_3742,N_3299,N_3205);
nand U3743 (N_3743,N_3447,N_3194);
nand U3744 (N_3744,N_3220,N_3289);
and U3745 (N_3745,N_3307,N_3363);
and U3746 (N_3746,N_3450,N_3302);
or U3747 (N_3747,N_3228,N_3303);
xnor U3748 (N_3748,N_3066,N_3411);
nand U3749 (N_3749,N_3380,N_3124);
nor U3750 (N_3750,N_3111,N_3203);
or U3751 (N_3751,N_3132,N_3353);
and U3752 (N_3752,N_3384,N_3370);
nand U3753 (N_3753,N_3368,N_3360);
nor U3754 (N_3754,N_3191,N_3399);
nor U3755 (N_3755,N_3021,N_3109);
xnor U3756 (N_3756,N_3210,N_3478);
xor U3757 (N_3757,N_3295,N_3359);
nor U3758 (N_3758,N_3258,N_3376);
nand U3759 (N_3759,N_3182,N_3043);
and U3760 (N_3760,N_3375,N_3031);
xor U3761 (N_3761,N_3459,N_3416);
or U3762 (N_3762,N_3373,N_3440);
or U3763 (N_3763,N_3002,N_3419);
or U3764 (N_3764,N_3239,N_3258);
xnor U3765 (N_3765,N_3307,N_3483);
nand U3766 (N_3766,N_3452,N_3280);
nor U3767 (N_3767,N_3479,N_3261);
and U3768 (N_3768,N_3035,N_3019);
nor U3769 (N_3769,N_3314,N_3163);
and U3770 (N_3770,N_3124,N_3248);
nor U3771 (N_3771,N_3046,N_3301);
xnor U3772 (N_3772,N_3126,N_3034);
xnor U3773 (N_3773,N_3373,N_3401);
nor U3774 (N_3774,N_3338,N_3109);
or U3775 (N_3775,N_3443,N_3021);
nand U3776 (N_3776,N_3167,N_3219);
xor U3777 (N_3777,N_3449,N_3216);
nand U3778 (N_3778,N_3403,N_3067);
and U3779 (N_3779,N_3190,N_3247);
xor U3780 (N_3780,N_3161,N_3205);
xor U3781 (N_3781,N_3332,N_3144);
xnor U3782 (N_3782,N_3107,N_3044);
xnor U3783 (N_3783,N_3098,N_3046);
nand U3784 (N_3784,N_3092,N_3047);
nand U3785 (N_3785,N_3441,N_3272);
and U3786 (N_3786,N_3101,N_3190);
xor U3787 (N_3787,N_3096,N_3199);
nor U3788 (N_3788,N_3171,N_3487);
and U3789 (N_3789,N_3226,N_3183);
and U3790 (N_3790,N_3096,N_3231);
and U3791 (N_3791,N_3033,N_3065);
or U3792 (N_3792,N_3036,N_3316);
nor U3793 (N_3793,N_3245,N_3046);
or U3794 (N_3794,N_3405,N_3189);
nand U3795 (N_3795,N_3491,N_3467);
xor U3796 (N_3796,N_3288,N_3220);
xnor U3797 (N_3797,N_3454,N_3492);
nor U3798 (N_3798,N_3387,N_3327);
nand U3799 (N_3799,N_3274,N_3046);
nor U3800 (N_3800,N_3235,N_3298);
nand U3801 (N_3801,N_3013,N_3035);
and U3802 (N_3802,N_3107,N_3184);
xor U3803 (N_3803,N_3381,N_3279);
xor U3804 (N_3804,N_3459,N_3109);
or U3805 (N_3805,N_3129,N_3041);
and U3806 (N_3806,N_3199,N_3203);
or U3807 (N_3807,N_3090,N_3349);
and U3808 (N_3808,N_3238,N_3185);
and U3809 (N_3809,N_3290,N_3096);
xor U3810 (N_3810,N_3065,N_3122);
nor U3811 (N_3811,N_3336,N_3391);
and U3812 (N_3812,N_3430,N_3242);
xnor U3813 (N_3813,N_3444,N_3207);
or U3814 (N_3814,N_3300,N_3386);
and U3815 (N_3815,N_3306,N_3369);
nand U3816 (N_3816,N_3462,N_3101);
xnor U3817 (N_3817,N_3247,N_3288);
or U3818 (N_3818,N_3363,N_3425);
or U3819 (N_3819,N_3145,N_3323);
xnor U3820 (N_3820,N_3225,N_3109);
xor U3821 (N_3821,N_3416,N_3152);
and U3822 (N_3822,N_3158,N_3344);
nand U3823 (N_3823,N_3188,N_3214);
xnor U3824 (N_3824,N_3369,N_3070);
nor U3825 (N_3825,N_3172,N_3111);
or U3826 (N_3826,N_3329,N_3379);
xor U3827 (N_3827,N_3118,N_3405);
or U3828 (N_3828,N_3222,N_3295);
xor U3829 (N_3829,N_3461,N_3050);
and U3830 (N_3830,N_3241,N_3216);
xnor U3831 (N_3831,N_3223,N_3002);
nand U3832 (N_3832,N_3084,N_3290);
xor U3833 (N_3833,N_3066,N_3058);
nand U3834 (N_3834,N_3350,N_3089);
nand U3835 (N_3835,N_3278,N_3238);
xor U3836 (N_3836,N_3355,N_3224);
nor U3837 (N_3837,N_3008,N_3156);
or U3838 (N_3838,N_3237,N_3109);
or U3839 (N_3839,N_3268,N_3463);
nor U3840 (N_3840,N_3431,N_3068);
or U3841 (N_3841,N_3172,N_3334);
xnor U3842 (N_3842,N_3184,N_3011);
or U3843 (N_3843,N_3247,N_3029);
xor U3844 (N_3844,N_3245,N_3117);
nand U3845 (N_3845,N_3408,N_3387);
or U3846 (N_3846,N_3133,N_3441);
or U3847 (N_3847,N_3344,N_3209);
nor U3848 (N_3848,N_3481,N_3207);
xor U3849 (N_3849,N_3002,N_3175);
nand U3850 (N_3850,N_3129,N_3392);
nand U3851 (N_3851,N_3162,N_3266);
or U3852 (N_3852,N_3082,N_3269);
or U3853 (N_3853,N_3366,N_3277);
nor U3854 (N_3854,N_3221,N_3303);
nand U3855 (N_3855,N_3305,N_3165);
or U3856 (N_3856,N_3490,N_3392);
and U3857 (N_3857,N_3327,N_3264);
and U3858 (N_3858,N_3054,N_3314);
or U3859 (N_3859,N_3158,N_3475);
nor U3860 (N_3860,N_3370,N_3121);
and U3861 (N_3861,N_3178,N_3227);
or U3862 (N_3862,N_3091,N_3121);
xnor U3863 (N_3863,N_3328,N_3173);
nand U3864 (N_3864,N_3224,N_3414);
nor U3865 (N_3865,N_3175,N_3254);
xor U3866 (N_3866,N_3346,N_3325);
xor U3867 (N_3867,N_3467,N_3167);
xor U3868 (N_3868,N_3011,N_3206);
xnor U3869 (N_3869,N_3178,N_3366);
or U3870 (N_3870,N_3349,N_3386);
and U3871 (N_3871,N_3198,N_3179);
nand U3872 (N_3872,N_3095,N_3307);
or U3873 (N_3873,N_3132,N_3225);
or U3874 (N_3874,N_3416,N_3121);
nor U3875 (N_3875,N_3155,N_3420);
xnor U3876 (N_3876,N_3386,N_3323);
or U3877 (N_3877,N_3137,N_3495);
or U3878 (N_3878,N_3064,N_3033);
or U3879 (N_3879,N_3047,N_3172);
nand U3880 (N_3880,N_3446,N_3140);
or U3881 (N_3881,N_3035,N_3419);
or U3882 (N_3882,N_3243,N_3285);
nand U3883 (N_3883,N_3388,N_3112);
nor U3884 (N_3884,N_3086,N_3379);
nand U3885 (N_3885,N_3424,N_3421);
or U3886 (N_3886,N_3194,N_3176);
nor U3887 (N_3887,N_3071,N_3230);
xnor U3888 (N_3888,N_3219,N_3082);
nor U3889 (N_3889,N_3160,N_3130);
and U3890 (N_3890,N_3013,N_3066);
or U3891 (N_3891,N_3066,N_3417);
xor U3892 (N_3892,N_3176,N_3193);
nand U3893 (N_3893,N_3252,N_3234);
xor U3894 (N_3894,N_3323,N_3118);
xor U3895 (N_3895,N_3447,N_3000);
nor U3896 (N_3896,N_3341,N_3058);
xnor U3897 (N_3897,N_3135,N_3491);
nor U3898 (N_3898,N_3226,N_3283);
and U3899 (N_3899,N_3387,N_3015);
nand U3900 (N_3900,N_3463,N_3228);
xor U3901 (N_3901,N_3338,N_3454);
and U3902 (N_3902,N_3372,N_3199);
or U3903 (N_3903,N_3068,N_3440);
xnor U3904 (N_3904,N_3206,N_3270);
nand U3905 (N_3905,N_3197,N_3061);
and U3906 (N_3906,N_3494,N_3228);
nand U3907 (N_3907,N_3231,N_3084);
or U3908 (N_3908,N_3412,N_3122);
and U3909 (N_3909,N_3084,N_3118);
nor U3910 (N_3910,N_3369,N_3272);
nand U3911 (N_3911,N_3483,N_3281);
nand U3912 (N_3912,N_3113,N_3273);
and U3913 (N_3913,N_3145,N_3298);
nor U3914 (N_3914,N_3431,N_3435);
nand U3915 (N_3915,N_3161,N_3145);
or U3916 (N_3916,N_3339,N_3343);
nand U3917 (N_3917,N_3199,N_3253);
and U3918 (N_3918,N_3101,N_3015);
nor U3919 (N_3919,N_3280,N_3250);
and U3920 (N_3920,N_3175,N_3274);
and U3921 (N_3921,N_3018,N_3114);
and U3922 (N_3922,N_3136,N_3169);
xor U3923 (N_3923,N_3380,N_3481);
xnor U3924 (N_3924,N_3446,N_3327);
or U3925 (N_3925,N_3388,N_3139);
xnor U3926 (N_3926,N_3265,N_3407);
xnor U3927 (N_3927,N_3292,N_3402);
nand U3928 (N_3928,N_3450,N_3342);
nor U3929 (N_3929,N_3197,N_3376);
or U3930 (N_3930,N_3331,N_3084);
nand U3931 (N_3931,N_3167,N_3141);
and U3932 (N_3932,N_3096,N_3075);
xor U3933 (N_3933,N_3388,N_3008);
nand U3934 (N_3934,N_3411,N_3368);
or U3935 (N_3935,N_3392,N_3454);
xor U3936 (N_3936,N_3311,N_3196);
xnor U3937 (N_3937,N_3385,N_3085);
and U3938 (N_3938,N_3315,N_3391);
nor U3939 (N_3939,N_3344,N_3172);
nor U3940 (N_3940,N_3355,N_3345);
or U3941 (N_3941,N_3202,N_3467);
xnor U3942 (N_3942,N_3303,N_3270);
and U3943 (N_3943,N_3178,N_3185);
xnor U3944 (N_3944,N_3071,N_3315);
nor U3945 (N_3945,N_3027,N_3453);
nand U3946 (N_3946,N_3412,N_3458);
and U3947 (N_3947,N_3019,N_3070);
xnor U3948 (N_3948,N_3068,N_3281);
or U3949 (N_3949,N_3081,N_3129);
or U3950 (N_3950,N_3186,N_3118);
or U3951 (N_3951,N_3268,N_3215);
and U3952 (N_3952,N_3447,N_3366);
xnor U3953 (N_3953,N_3426,N_3421);
xor U3954 (N_3954,N_3214,N_3355);
and U3955 (N_3955,N_3090,N_3445);
nor U3956 (N_3956,N_3302,N_3208);
or U3957 (N_3957,N_3145,N_3497);
nor U3958 (N_3958,N_3244,N_3065);
or U3959 (N_3959,N_3395,N_3337);
xnor U3960 (N_3960,N_3045,N_3199);
xnor U3961 (N_3961,N_3071,N_3336);
nand U3962 (N_3962,N_3163,N_3223);
nor U3963 (N_3963,N_3000,N_3127);
xnor U3964 (N_3964,N_3130,N_3047);
nor U3965 (N_3965,N_3479,N_3226);
and U3966 (N_3966,N_3185,N_3216);
nor U3967 (N_3967,N_3442,N_3028);
nand U3968 (N_3968,N_3231,N_3276);
and U3969 (N_3969,N_3127,N_3250);
and U3970 (N_3970,N_3320,N_3307);
nor U3971 (N_3971,N_3296,N_3349);
or U3972 (N_3972,N_3312,N_3475);
and U3973 (N_3973,N_3136,N_3251);
xnor U3974 (N_3974,N_3323,N_3141);
nand U3975 (N_3975,N_3175,N_3359);
nand U3976 (N_3976,N_3208,N_3351);
nor U3977 (N_3977,N_3333,N_3319);
nor U3978 (N_3978,N_3299,N_3062);
xor U3979 (N_3979,N_3485,N_3405);
nand U3980 (N_3980,N_3054,N_3014);
xnor U3981 (N_3981,N_3004,N_3062);
or U3982 (N_3982,N_3051,N_3156);
nor U3983 (N_3983,N_3071,N_3005);
nand U3984 (N_3984,N_3197,N_3152);
xnor U3985 (N_3985,N_3225,N_3323);
xor U3986 (N_3986,N_3469,N_3060);
or U3987 (N_3987,N_3001,N_3109);
xor U3988 (N_3988,N_3024,N_3267);
xnor U3989 (N_3989,N_3274,N_3425);
xnor U3990 (N_3990,N_3028,N_3417);
nor U3991 (N_3991,N_3224,N_3018);
and U3992 (N_3992,N_3118,N_3027);
xor U3993 (N_3993,N_3270,N_3110);
and U3994 (N_3994,N_3186,N_3336);
and U3995 (N_3995,N_3006,N_3045);
nor U3996 (N_3996,N_3201,N_3097);
xor U3997 (N_3997,N_3404,N_3183);
nand U3998 (N_3998,N_3048,N_3121);
and U3999 (N_3999,N_3033,N_3242);
xnor U4000 (N_4000,N_3886,N_3506);
and U4001 (N_4001,N_3968,N_3723);
nand U4002 (N_4002,N_3975,N_3809);
xnor U4003 (N_4003,N_3790,N_3631);
nor U4004 (N_4004,N_3696,N_3837);
and U4005 (N_4005,N_3547,N_3966);
nor U4006 (N_4006,N_3662,N_3930);
nand U4007 (N_4007,N_3819,N_3843);
and U4008 (N_4008,N_3762,N_3946);
and U4009 (N_4009,N_3561,N_3761);
nor U4010 (N_4010,N_3636,N_3539);
xnor U4011 (N_4011,N_3524,N_3647);
xor U4012 (N_4012,N_3667,N_3535);
nand U4013 (N_4013,N_3801,N_3879);
and U4014 (N_4014,N_3604,N_3536);
nand U4015 (N_4015,N_3908,N_3791);
and U4016 (N_4016,N_3534,N_3617);
nor U4017 (N_4017,N_3601,N_3677);
nand U4018 (N_4018,N_3693,N_3513);
nor U4019 (N_4019,N_3951,N_3666);
nor U4020 (N_4020,N_3736,N_3960);
nand U4021 (N_4021,N_3713,N_3896);
or U4022 (N_4022,N_3740,N_3532);
and U4023 (N_4023,N_3518,N_3597);
and U4024 (N_4024,N_3562,N_3977);
xor U4025 (N_4025,N_3575,N_3942);
xnor U4026 (N_4026,N_3796,N_3804);
nand U4027 (N_4027,N_3721,N_3774);
or U4028 (N_4028,N_3555,N_3656);
and U4029 (N_4029,N_3755,N_3730);
nor U4030 (N_4030,N_3607,N_3620);
and U4031 (N_4031,N_3654,N_3888);
and U4032 (N_4032,N_3593,N_3890);
nand U4033 (N_4033,N_3912,N_3688);
nor U4034 (N_4034,N_3906,N_3619);
nand U4035 (N_4035,N_3627,N_3997);
xor U4036 (N_4036,N_3588,N_3559);
nand U4037 (N_4037,N_3797,N_3786);
nand U4038 (N_4038,N_3611,N_3698);
and U4039 (N_4039,N_3687,N_3978);
nor U4040 (N_4040,N_3871,N_3976);
xnor U4041 (N_4041,N_3516,N_3509);
and U4042 (N_4042,N_3515,N_3629);
nor U4043 (N_4043,N_3616,N_3982);
nand U4044 (N_4044,N_3959,N_3807);
xor U4045 (N_4045,N_3727,N_3702);
nor U4046 (N_4046,N_3928,N_3504);
nor U4047 (N_4047,N_3899,N_3738);
xor U4048 (N_4048,N_3981,N_3712);
nand U4049 (N_4049,N_3512,N_3757);
and U4050 (N_4050,N_3766,N_3560);
nor U4051 (N_4051,N_3963,N_3709);
nor U4052 (N_4052,N_3722,N_3889);
nor U4053 (N_4053,N_3686,N_3500);
nand U4054 (N_4054,N_3983,N_3840);
nor U4055 (N_4055,N_3695,N_3805);
nor U4056 (N_4056,N_3557,N_3967);
and U4057 (N_4057,N_3670,N_3910);
nor U4058 (N_4058,N_3567,N_3935);
nand U4059 (N_4059,N_3682,N_3759);
nand U4060 (N_4060,N_3582,N_3577);
nor U4061 (N_4061,N_3718,N_3638);
nor U4062 (N_4062,N_3590,N_3566);
or U4063 (N_4063,N_3626,N_3992);
and U4064 (N_4064,N_3770,N_3583);
nand U4065 (N_4065,N_3692,N_3955);
and U4066 (N_4066,N_3948,N_3668);
nor U4067 (N_4067,N_3584,N_3589);
nor U4068 (N_4068,N_3657,N_3551);
xor U4069 (N_4069,N_3877,N_3831);
nor U4070 (N_4070,N_3537,N_3674);
and U4071 (N_4071,N_3939,N_3909);
and U4072 (N_4072,N_3507,N_3731);
nor U4073 (N_4073,N_3943,N_3733);
nand U4074 (N_4074,N_3962,N_3663);
and U4075 (N_4075,N_3864,N_3618);
nor U4076 (N_4076,N_3749,N_3684);
xor U4077 (N_4077,N_3641,N_3918);
nor U4078 (N_4078,N_3606,N_3933);
nand U4079 (N_4079,N_3503,N_3845);
nand U4080 (N_4080,N_3985,N_3549);
or U4081 (N_4081,N_3869,N_3699);
xor U4082 (N_4082,N_3573,N_3958);
and U4083 (N_4083,N_3758,N_3768);
or U4084 (N_4084,N_3979,N_3865);
nand U4085 (N_4085,N_3907,N_3765);
or U4086 (N_4086,N_3706,N_3818);
nand U4087 (N_4087,N_3803,N_3510);
xor U4088 (N_4088,N_3875,N_3836);
nand U4089 (N_4089,N_3614,N_3707);
and U4090 (N_4090,N_3711,N_3891);
or U4091 (N_4091,N_3940,N_3971);
nand U4092 (N_4092,N_3862,N_3863);
and U4093 (N_4093,N_3756,N_3897);
nand U4094 (N_4094,N_3779,N_3690);
nor U4095 (N_4095,N_3591,N_3576);
and U4096 (N_4096,N_3911,N_3554);
or U4097 (N_4097,N_3822,N_3934);
or U4098 (N_4098,N_3697,N_3676);
nor U4099 (N_4099,N_3915,N_3505);
nand U4100 (N_4100,N_3605,N_3720);
or U4101 (N_4101,N_3926,N_3900);
nor U4102 (N_4102,N_3645,N_3587);
nor U4103 (N_4103,N_3598,N_3988);
nand U4104 (N_4104,N_3530,N_3970);
and U4105 (N_4105,N_3511,N_3672);
and U4106 (N_4106,N_3776,N_3866);
and U4107 (N_4107,N_3525,N_3793);
nand U4108 (N_4108,N_3552,N_3528);
xor U4109 (N_4109,N_3508,N_3944);
nand U4110 (N_4110,N_3887,N_3628);
or U4111 (N_4111,N_3609,N_3777);
and U4112 (N_4112,N_3522,N_3834);
nor U4113 (N_4113,N_3961,N_3594);
or U4114 (N_4114,N_3816,N_3635);
or U4115 (N_4115,N_3991,N_3613);
and U4116 (N_4116,N_3680,N_3823);
xor U4117 (N_4117,N_3853,N_3742);
nand U4118 (N_4118,N_3844,N_3633);
nand U4119 (N_4119,N_3568,N_3773);
and U4120 (N_4120,N_3748,N_3994);
nor U4121 (N_4121,N_3732,N_3519);
and U4122 (N_4122,N_3728,N_3980);
and U4123 (N_4123,N_3655,N_3838);
xor U4124 (N_4124,N_3531,N_3745);
nor U4125 (N_4125,N_3743,N_3719);
and U4126 (N_4126,N_3828,N_3610);
and U4127 (N_4127,N_3529,N_3545);
and U4128 (N_4128,N_3673,N_3872);
nor U4129 (N_4129,N_3927,N_3945);
and U4130 (N_4130,N_3810,N_3581);
xnor U4131 (N_4131,N_3789,N_3726);
nand U4132 (N_4132,N_3920,N_3964);
nand U4133 (N_4133,N_3556,N_3553);
xnor U4134 (N_4134,N_3775,N_3744);
or U4135 (N_4135,N_3894,N_3929);
nor U4136 (N_4136,N_3632,N_3881);
and U4137 (N_4137,N_3901,N_3989);
or U4138 (N_4138,N_3760,N_3919);
nand U4139 (N_4139,N_3754,N_3624);
nor U4140 (N_4140,N_3652,N_3716);
nand U4141 (N_4141,N_3651,N_3665);
and U4142 (N_4142,N_3832,N_3850);
or U4143 (N_4143,N_3788,N_3675);
and U4144 (N_4144,N_3785,N_3705);
nand U4145 (N_4145,N_3847,N_3826);
and U4146 (N_4146,N_3973,N_3800);
and U4147 (N_4147,N_3859,N_3572);
nor U4148 (N_4148,N_3694,N_3579);
and U4149 (N_4149,N_3501,N_3679);
nor U4150 (N_4150,N_3842,N_3903);
and U4151 (N_4151,N_3725,N_3922);
nor U4152 (N_4152,N_3905,N_3867);
nor U4153 (N_4153,N_3569,N_3746);
or U4154 (N_4154,N_3787,N_3650);
xnor U4155 (N_4155,N_3639,N_3841);
and U4156 (N_4156,N_3565,N_3520);
and U4157 (N_4157,N_3729,N_3764);
and U4158 (N_4158,N_3857,N_3714);
or U4159 (N_4159,N_3811,N_3808);
xor U4160 (N_4160,N_3936,N_3703);
nor U4161 (N_4161,N_3681,N_3846);
nor U4162 (N_4162,N_3851,N_3794);
xor U4163 (N_4163,N_3602,N_3526);
nand U4164 (N_4164,N_3778,N_3986);
nor U4165 (N_4165,N_3615,N_3972);
nor U4166 (N_4166,N_3792,N_3683);
xor U4167 (N_4167,N_3678,N_3741);
xnor U4168 (N_4168,N_3739,N_3974);
xnor U4169 (N_4169,N_3839,N_3885);
nand U4170 (N_4170,N_3752,N_3932);
xnor U4171 (N_4171,N_3817,N_3521);
xnor U4172 (N_4172,N_3824,N_3820);
xnor U4173 (N_4173,N_3852,N_3646);
and U4174 (N_4174,N_3541,N_3916);
and U4175 (N_4175,N_3814,N_3987);
nor U4176 (N_4176,N_3671,N_3585);
nand U4177 (N_4177,N_3813,N_3874);
or U4178 (N_4178,N_3659,N_3600);
nand U4179 (N_4179,N_3898,N_3815);
nand U4180 (N_4180,N_3802,N_3751);
xnor U4181 (N_4181,N_3917,N_3795);
nand U4182 (N_4182,N_3873,N_3625);
or U4183 (N_4183,N_3586,N_3855);
nor U4184 (N_4184,N_3644,N_3848);
nand U4185 (N_4185,N_3548,N_3799);
xnor U4186 (N_4186,N_3542,N_3747);
nand U4187 (N_4187,N_3737,N_3514);
nor U4188 (N_4188,N_3941,N_3685);
and U4189 (N_4189,N_3861,N_3984);
nor U4190 (N_4190,N_3999,N_3782);
xnor U4191 (N_4191,N_3781,N_3595);
nor U4192 (N_4192,N_3772,N_3715);
and U4193 (N_4193,N_3517,N_3753);
nand U4194 (N_4194,N_3658,N_3868);
or U4195 (N_4195,N_3876,N_3830);
nor U4196 (N_4196,N_3883,N_3950);
or U4197 (N_4197,N_3637,N_3704);
nand U4198 (N_4198,N_3750,N_3735);
nor U4199 (N_4199,N_3564,N_3767);
xnor U4200 (N_4200,N_3734,N_3550);
xnor U4201 (N_4201,N_3812,N_3546);
xnor U4202 (N_4202,N_3882,N_3701);
xnor U4203 (N_4203,N_3621,N_3931);
nand U4204 (N_4204,N_3806,N_3578);
xor U4205 (N_4205,N_3612,N_3769);
xnor U4206 (N_4206,N_3902,N_3630);
or U4207 (N_4207,N_3763,N_3558);
nor U4208 (N_4208,N_3798,N_3710);
xor U4209 (N_4209,N_3827,N_3821);
or U4210 (N_4210,N_3904,N_3953);
xnor U4211 (N_4211,N_3856,N_3623);
and U4212 (N_4212,N_3527,N_3825);
and U4213 (N_4213,N_3957,N_3523);
or U4214 (N_4214,N_3592,N_3689);
or U4215 (N_4215,N_3533,N_3913);
nor U4216 (N_4216,N_3661,N_3544);
and U4217 (N_4217,N_3640,N_3858);
and U4218 (N_4218,N_3993,N_3771);
or U4219 (N_4219,N_3538,N_3717);
nand U4220 (N_4220,N_3574,N_3780);
or U4221 (N_4221,N_3880,N_3634);
xnor U4222 (N_4222,N_3691,N_3502);
nor U4223 (N_4223,N_3938,N_3829);
xnor U4224 (N_4224,N_3956,N_3700);
xnor U4225 (N_4225,N_3540,N_3599);
nor U4226 (N_4226,N_3870,N_3608);
and U4227 (N_4227,N_3708,N_3893);
xor U4228 (N_4228,N_3664,N_3996);
nor U4229 (N_4229,N_3849,N_3724);
or U4230 (N_4230,N_3603,N_3925);
nor U4231 (N_4231,N_3884,N_3923);
nand U4232 (N_4232,N_3570,N_3669);
xnor U4233 (N_4233,N_3965,N_3835);
and U4234 (N_4234,N_3543,N_3833);
nor U4235 (N_4235,N_3947,N_3914);
or U4236 (N_4236,N_3784,N_3924);
nor U4237 (N_4237,N_3854,N_3921);
or U4238 (N_4238,N_3642,N_3643);
and U4239 (N_4239,N_3648,N_3783);
xor U4240 (N_4240,N_3660,N_3895);
nor U4241 (N_4241,N_3892,N_3998);
or U4242 (N_4242,N_3937,N_3622);
or U4243 (N_4243,N_3653,N_3969);
and U4244 (N_4244,N_3954,N_3580);
nor U4245 (N_4245,N_3990,N_3571);
or U4246 (N_4246,N_3649,N_3563);
or U4247 (N_4247,N_3878,N_3860);
nor U4248 (N_4248,N_3995,N_3949);
or U4249 (N_4249,N_3952,N_3596);
and U4250 (N_4250,N_3688,N_3966);
nand U4251 (N_4251,N_3932,N_3826);
nand U4252 (N_4252,N_3989,N_3571);
xnor U4253 (N_4253,N_3656,N_3896);
and U4254 (N_4254,N_3668,N_3542);
nor U4255 (N_4255,N_3595,N_3757);
nand U4256 (N_4256,N_3702,N_3562);
nor U4257 (N_4257,N_3826,N_3851);
nand U4258 (N_4258,N_3929,N_3611);
nand U4259 (N_4259,N_3717,N_3667);
nor U4260 (N_4260,N_3680,N_3544);
or U4261 (N_4261,N_3693,N_3725);
nand U4262 (N_4262,N_3789,N_3756);
and U4263 (N_4263,N_3804,N_3712);
or U4264 (N_4264,N_3958,N_3914);
nor U4265 (N_4265,N_3973,N_3545);
nor U4266 (N_4266,N_3945,N_3503);
nor U4267 (N_4267,N_3723,N_3667);
and U4268 (N_4268,N_3547,N_3928);
and U4269 (N_4269,N_3964,N_3798);
or U4270 (N_4270,N_3527,N_3982);
or U4271 (N_4271,N_3502,N_3955);
xor U4272 (N_4272,N_3711,N_3967);
and U4273 (N_4273,N_3903,N_3636);
nor U4274 (N_4274,N_3781,N_3510);
nor U4275 (N_4275,N_3587,N_3652);
nor U4276 (N_4276,N_3689,N_3745);
xnor U4277 (N_4277,N_3902,N_3855);
or U4278 (N_4278,N_3575,N_3752);
or U4279 (N_4279,N_3609,N_3922);
nor U4280 (N_4280,N_3802,N_3986);
nand U4281 (N_4281,N_3538,N_3873);
or U4282 (N_4282,N_3781,N_3898);
nor U4283 (N_4283,N_3514,N_3848);
and U4284 (N_4284,N_3530,N_3986);
and U4285 (N_4285,N_3646,N_3672);
nand U4286 (N_4286,N_3617,N_3629);
xor U4287 (N_4287,N_3669,N_3790);
and U4288 (N_4288,N_3593,N_3981);
xnor U4289 (N_4289,N_3807,N_3845);
nor U4290 (N_4290,N_3771,N_3910);
nor U4291 (N_4291,N_3734,N_3773);
nand U4292 (N_4292,N_3834,N_3540);
nand U4293 (N_4293,N_3617,N_3624);
xnor U4294 (N_4294,N_3668,N_3775);
or U4295 (N_4295,N_3578,N_3894);
and U4296 (N_4296,N_3540,N_3857);
nand U4297 (N_4297,N_3555,N_3983);
and U4298 (N_4298,N_3892,N_3767);
or U4299 (N_4299,N_3640,N_3589);
or U4300 (N_4300,N_3998,N_3930);
xnor U4301 (N_4301,N_3628,N_3737);
or U4302 (N_4302,N_3754,N_3836);
and U4303 (N_4303,N_3876,N_3591);
nor U4304 (N_4304,N_3752,N_3767);
and U4305 (N_4305,N_3908,N_3809);
nor U4306 (N_4306,N_3674,N_3535);
nor U4307 (N_4307,N_3531,N_3592);
nor U4308 (N_4308,N_3698,N_3881);
nand U4309 (N_4309,N_3737,N_3808);
and U4310 (N_4310,N_3969,N_3631);
xor U4311 (N_4311,N_3764,N_3748);
or U4312 (N_4312,N_3804,N_3553);
xor U4313 (N_4313,N_3535,N_3759);
or U4314 (N_4314,N_3936,N_3668);
and U4315 (N_4315,N_3781,N_3934);
nand U4316 (N_4316,N_3777,N_3573);
nand U4317 (N_4317,N_3675,N_3549);
or U4318 (N_4318,N_3872,N_3830);
xnor U4319 (N_4319,N_3599,N_3828);
or U4320 (N_4320,N_3614,N_3506);
or U4321 (N_4321,N_3979,N_3685);
and U4322 (N_4322,N_3685,N_3908);
xor U4323 (N_4323,N_3545,N_3882);
nor U4324 (N_4324,N_3641,N_3547);
or U4325 (N_4325,N_3556,N_3502);
or U4326 (N_4326,N_3993,N_3826);
xor U4327 (N_4327,N_3854,N_3678);
nand U4328 (N_4328,N_3968,N_3709);
xor U4329 (N_4329,N_3503,N_3948);
and U4330 (N_4330,N_3819,N_3509);
nor U4331 (N_4331,N_3908,N_3743);
xor U4332 (N_4332,N_3619,N_3813);
nor U4333 (N_4333,N_3992,N_3932);
or U4334 (N_4334,N_3964,N_3780);
nor U4335 (N_4335,N_3888,N_3641);
xnor U4336 (N_4336,N_3584,N_3646);
or U4337 (N_4337,N_3582,N_3764);
or U4338 (N_4338,N_3871,N_3626);
xnor U4339 (N_4339,N_3568,N_3728);
nand U4340 (N_4340,N_3872,N_3773);
nand U4341 (N_4341,N_3599,N_3693);
xor U4342 (N_4342,N_3529,N_3547);
and U4343 (N_4343,N_3902,N_3769);
and U4344 (N_4344,N_3981,N_3581);
nor U4345 (N_4345,N_3535,N_3615);
or U4346 (N_4346,N_3929,N_3778);
or U4347 (N_4347,N_3921,N_3539);
nor U4348 (N_4348,N_3883,N_3584);
nand U4349 (N_4349,N_3957,N_3562);
or U4350 (N_4350,N_3869,N_3899);
nand U4351 (N_4351,N_3903,N_3544);
and U4352 (N_4352,N_3800,N_3688);
nand U4353 (N_4353,N_3818,N_3739);
and U4354 (N_4354,N_3734,N_3767);
nor U4355 (N_4355,N_3980,N_3992);
xor U4356 (N_4356,N_3571,N_3743);
or U4357 (N_4357,N_3780,N_3555);
and U4358 (N_4358,N_3703,N_3945);
nor U4359 (N_4359,N_3913,N_3932);
xor U4360 (N_4360,N_3539,N_3591);
or U4361 (N_4361,N_3734,N_3588);
xor U4362 (N_4362,N_3557,N_3514);
nand U4363 (N_4363,N_3823,N_3721);
xor U4364 (N_4364,N_3546,N_3928);
nor U4365 (N_4365,N_3802,N_3749);
xnor U4366 (N_4366,N_3578,N_3621);
or U4367 (N_4367,N_3674,N_3665);
and U4368 (N_4368,N_3766,N_3915);
and U4369 (N_4369,N_3614,N_3783);
xor U4370 (N_4370,N_3563,N_3545);
xor U4371 (N_4371,N_3792,N_3891);
or U4372 (N_4372,N_3703,N_3524);
nor U4373 (N_4373,N_3684,N_3816);
xnor U4374 (N_4374,N_3500,N_3815);
nand U4375 (N_4375,N_3554,N_3935);
xnor U4376 (N_4376,N_3863,N_3544);
nand U4377 (N_4377,N_3627,N_3631);
nor U4378 (N_4378,N_3974,N_3565);
xnor U4379 (N_4379,N_3942,N_3793);
or U4380 (N_4380,N_3664,N_3677);
xor U4381 (N_4381,N_3755,N_3920);
nor U4382 (N_4382,N_3691,N_3604);
nor U4383 (N_4383,N_3909,N_3731);
nand U4384 (N_4384,N_3833,N_3624);
or U4385 (N_4385,N_3516,N_3700);
xnor U4386 (N_4386,N_3723,N_3644);
or U4387 (N_4387,N_3963,N_3928);
nor U4388 (N_4388,N_3836,N_3559);
or U4389 (N_4389,N_3568,N_3879);
nand U4390 (N_4390,N_3589,N_3558);
xnor U4391 (N_4391,N_3914,N_3500);
or U4392 (N_4392,N_3763,N_3668);
and U4393 (N_4393,N_3808,N_3775);
nand U4394 (N_4394,N_3663,N_3619);
nor U4395 (N_4395,N_3685,N_3981);
nand U4396 (N_4396,N_3921,N_3558);
and U4397 (N_4397,N_3665,N_3626);
nor U4398 (N_4398,N_3511,N_3996);
or U4399 (N_4399,N_3807,N_3960);
nor U4400 (N_4400,N_3749,N_3905);
nor U4401 (N_4401,N_3611,N_3552);
nand U4402 (N_4402,N_3814,N_3591);
or U4403 (N_4403,N_3925,N_3795);
xnor U4404 (N_4404,N_3965,N_3505);
nand U4405 (N_4405,N_3814,N_3706);
xor U4406 (N_4406,N_3637,N_3933);
xnor U4407 (N_4407,N_3860,N_3817);
nor U4408 (N_4408,N_3835,N_3555);
nor U4409 (N_4409,N_3990,N_3623);
xnor U4410 (N_4410,N_3855,N_3898);
xnor U4411 (N_4411,N_3667,N_3674);
xor U4412 (N_4412,N_3836,N_3561);
xor U4413 (N_4413,N_3815,N_3639);
or U4414 (N_4414,N_3635,N_3901);
nand U4415 (N_4415,N_3697,N_3656);
nand U4416 (N_4416,N_3765,N_3938);
xor U4417 (N_4417,N_3835,N_3878);
xnor U4418 (N_4418,N_3695,N_3981);
nand U4419 (N_4419,N_3858,N_3606);
xor U4420 (N_4420,N_3896,N_3916);
or U4421 (N_4421,N_3757,N_3793);
nand U4422 (N_4422,N_3739,N_3856);
nor U4423 (N_4423,N_3738,N_3597);
and U4424 (N_4424,N_3672,N_3892);
or U4425 (N_4425,N_3953,N_3507);
xnor U4426 (N_4426,N_3546,N_3791);
nand U4427 (N_4427,N_3753,N_3722);
xnor U4428 (N_4428,N_3537,N_3806);
nand U4429 (N_4429,N_3980,N_3658);
xor U4430 (N_4430,N_3920,N_3660);
nand U4431 (N_4431,N_3658,N_3729);
xor U4432 (N_4432,N_3858,N_3530);
xnor U4433 (N_4433,N_3836,N_3604);
xnor U4434 (N_4434,N_3828,N_3660);
and U4435 (N_4435,N_3500,N_3834);
and U4436 (N_4436,N_3833,N_3752);
and U4437 (N_4437,N_3781,N_3967);
and U4438 (N_4438,N_3823,N_3708);
xnor U4439 (N_4439,N_3856,N_3899);
and U4440 (N_4440,N_3657,N_3567);
nor U4441 (N_4441,N_3955,N_3865);
or U4442 (N_4442,N_3660,N_3777);
nor U4443 (N_4443,N_3940,N_3885);
nand U4444 (N_4444,N_3528,N_3926);
nand U4445 (N_4445,N_3969,N_3618);
nand U4446 (N_4446,N_3819,N_3712);
nor U4447 (N_4447,N_3969,N_3848);
nand U4448 (N_4448,N_3853,N_3941);
nand U4449 (N_4449,N_3510,N_3993);
nand U4450 (N_4450,N_3512,N_3915);
nor U4451 (N_4451,N_3833,N_3885);
nor U4452 (N_4452,N_3505,N_3638);
xnor U4453 (N_4453,N_3856,N_3846);
or U4454 (N_4454,N_3785,N_3716);
and U4455 (N_4455,N_3700,N_3938);
xor U4456 (N_4456,N_3550,N_3724);
nand U4457 (N_4457,N_3798,N_3671);
nand U4458 (N_4458,N_3768,N_3733);
and U4459 (N_4459,N_3822,N_3753);
xor U4460 (N_4460,N_3549,N_3737);
and U4461 (N_4461,N_3989,N_3663);
nand U4462 (N_4462,N_3610,N_3707);
or U4463 (N_4463,N_3764,N_3591);
and U4464 (N_4464,N_3890,N_3565);
xnor U4465 (N_4465,N_3658,N_3671);
or U4466 (N_4466,N_3753,N_3882);
and U4467 (N_4467,N_3912,N_3606);
xnor U4468 (N_4468,N_3599,N_3842);
nor U4469 (N_4469,N_3988,N_3647);
and U4470 (N_4470,N_3735,N_3747);
xnor U4471 (N_4471,N_3668,N_3675);
xor U4472 (N_4472,N_3799,N_3813);
nor U4473 (N_4473,N_3709,N_3978);
xor U4474 (N_4474,N_3800,N_3524);
nor U4475 (N_4475,N_3793,N_3826);
or U4476 (N_4476,N_3508,N_3896);
nor U4477 (N_4477,N_3505,N_3944);
or U4478 (N_4478,N_3971,N_3658);
or U4479 (N_4479,N_3656,N_3644);
nor U4480 (N_4480,N_3599,N_3759);
nor U4481 (N_4481,N_3644,N_3760);
nand U4482 (N_4482,N_3712,N_3926);
nor U4483 (N_4483,N_3771,N_3840);
or U4484 (N_4484,N_3970,N_3529);
nor U4485 (N_4485,N_3562,N_3645);
nor U4486 (N_4486,N_3972,N_3820);
xnor U4487 (N_4487,N_3513,N_3577);
or U4488 (N_4488,N_3628,N_3876);
or U4489 (N_4489,N_3534,N_3981);
xor U4490 (N_4490,N_3867,N_3535);
xnor U4491 (N_4491,N_3980,N_3720);
and U4492 (N_4492,N_3974,N_3910);
xnor U4493 (N_4493,N_3913,N_3680);
nor U4494 (N_4494,N_3768,N_3702);
or U4495 (N_4495,N_3503,N_3599);
or U4496 (N_4496,N_3947,N_3901);
nand U4497 (N_4497,N_3990,N_3542);
nand U4498 (N_4498,N_3571,N_3789);
nor U4499 (N_4499,N_3943,N_3827);
or U4500 (N_4500,N_4268,N_4345);
nand U4501 (N_4501,N_4449,N_4298);
xor U4502 (N_4502,N_4464,N_4071);
nor U4503 (N_4503,N_4107,N_4208);
or U4504 (N_4504,N_4392,N_4012);
or U4505 (N_4505,N_4431,N_4276);
nor U4506 (N_4506,N_4424,N_4486);
and U4507 (N_4507,N_4415,N_4144);
nand U4508 (N_4508,N_4153,N_4084);
or U4509 (N_4509,N_4381,N_4390);
or U4510 (N_4510,N_4356,N_4172);
or U4511 (N_4511,N_4458,N_4343);
nand U4512 (N_4512,N_4081,N_4294);
and U4513 (N_4513,N_4272,N_4467);
nor U4514 (N_4514,N_4309,N_4470);
nor U4515 (N_4515,N_4443,N_4151);
xnor U4516 (N_4516,N_4375,N_4197);
or U4517 (N_4517,N_4454,N_4473);
xnor U4518 (N_4518,N_4179,N_4279);
and U4519 (N_4519,N_4429,N_4273);
and U4520 (N_4520,N_4036,N_4230);
xor U4521 (N_4521,N_4111,N_4001);
or U4522 (N_4522,N_4237,N_4337);
nor U4523 (N_4523,N_4320,N_4317);
or U4524 (N_4524,N_4070,N_4421);
xor U4525 (N_4525,N_4060,N_4086);
nor U4526 (N_4526,N_4231,N_4117);
nor U4527 (N_4527,N_4485,N_4112);
or U4528 (N_4528,N_4057,N_4394);
nand U4529 (N_4529,N_4247,N_4064);
or U4530 (N_4530,N_4270,N_4336);
xor U4531 (N_4531,N_4203,N_4187);
and U4532 (N_4532,N_4040,N_4284);
and U4533 (N_4533,N_4372,N_4166);
or U4534 (N_4534,N_4063,N_4009);
nand U4535 (N_4535,N_4435,N_4286);
and U4536 (N_4536,N_4366,N_4481);
or U4537 (N_4537,N_4008,N_4432);
or U4538 (N_4538,N_4027,N_4422);
nor U4539 (N_4539,N_4423,N_4271);
nor U4540 (N_4540,N_4174,N_4065);
and U4541 (N_4541,N_4314,N_4163);
or U4542 (N_4542,N_4085,N_4358);
nor U4543 (N_4543,N_4398,N_4183);
nor U4544 (N_4544,N_4258,N_4096);
or U4545 (N_4545,N_4420,N_4411);
nand U4546 (N_4546,N_4000,N_4005);
and U4547 (N_4547,N_4243,N_4408);
nor U4548 (N_4548,N_4266,N_4251);
or U4549 (N_4549,N_4130,N_4329);
and U4550 (N_4550,N_4407,N_4169);
nor U4551 (N_4551,N_4078,N_4410);
nor U4552 (N_4552,N_4457,N_4121);
nor U4553 (N_4553,N_4168,N_4134);
nor U4554 (N_4554,N_4210,N_4461);
nor U4555 (N_4555,N_4010,N_4220);
nand U4556 (N_4556,N_4020,N_4003);
nand U4557 (N_4557,N_4437,N_4412);
nor U4558 (N_4558,N_4325,N_4100);
nand U4559 (N_4559,N_4239,N_4355);
and U4560 (N_4560,N_4048,N_4339);
xor U4561 (N_4561,N_4054,N_4075);
xor U4562 (N_4562,N_4116,N_4438);
nand U4563 (N_4563,N_4155,N_4221);
and U4564 (N_4564,N_4290,N_4182);
nand U4565 (N_4565,N_4259,N_4335);
nor U4566 (N_4566,N_4206,N_4032);
nand U4567 (N_4567,N_4326,N_4088);
and U4568 (N_4568,N_4049,N_4154);
nor U4569 (N_4569,N_4436,N_4159);
and U4570 (N_4570,N_4139,N_4141);
or U4571 (N_4571,N_4022,N_4311);
nand U4572 (N_4572,N_4280,N_4434);
nor U4573 (N_4573,N_4142,N_4489);
xnor U4574 (N_4574,N_4149,N_4226);
or U4575 (N_4575,N_4277,N_4393);
nor U4576 (N_4576,N_4232,N_4330);
nand U4577 (N_4577,N_4108,N_4228);
nor U4578 (N_4578,N_4033,N_4246);
xor U4579 (N_4579,N_4475,N_4338);
or U4580 (N_4580,N_4254,N_4238);
nand U4581 (N_4581,N_4453,N_4030);
nand U4582 (N_4582,N_4171,N_4414);
xnor U4583 (N_4583,N_4176,N_4318);
nor U4584 (N_4584,N_4214,N_4255);
nor U4585 (N_4585,N_4248,N_4133);
or U4586 (N_4586,N_4476,N_4409);
xor U4587 (N_4587,N_4045,N_4161);
xnor U4588 (N_4588,N_4403,N_4496);
nor U4589 (N_4589,N_4162,N_4334);
and U4590 (N_4590,N_4360,N_4310);
nor U4591 (N_4591,N_4354,N_4331);
or U4592 (N_4592,N_4028,N_4397);
and U4593 (N_4593,N_4074,N_4348);
nand U4594 (N_4594,N_4387,N_4384);
nor U4595 (N_4595,N_4031,N_4115);
or U4596 (N_4596,N_4080,N_4050);
and U4597 (N_4597,N_4287,N_4223);
nand U4598 (N_4598,N_4455,N_4011);
nand U4599 (N_4599,N_4077,N_4440);
xnor U4600 (N_4600,N_4105,N_4289);
xnor U4601 (N_4601,N_4364,N_4465);
nand U4602 (N_4602,N_4146,N_4102);
nor U4603 (N_4603,N_4201,N_4477);
nand U4604 (N_4604,N_4383,N_4262);
xnor U4605 (N_4605,N_4138,N_4006);
nand U4606 (N_4606,N_4321,N_4260);
nand U4607 (N_4607,N_4341,N_4079);
nor U4608 (N_4608,N_4216,N_4186);
or U4609 (N_4609,N_4059,N_4180);
and U4610 (N_4610,N_4474,N_4352);
nand U4611 (N_4611,N_4445,N_4382);
nand U4612 (N_4612,N_4098,N_4113);
nand U4613 (N_4613,N_4093,N_4026);
xnor U4614 (N_4614,N_4456,N_4361);
or U4615 (N_4615,N_4488,N_4224);
nand U4616 (N_4616,N_4484,N_4189);
xor U4617 (N_4617,N_4332,N_4209);
xor U4618 (N_4618,N_4158,N_4413);
nand U4619 (N_4619,N_4013,N_4192);
nand U4620 (N_4620,N_4056,N_4150);
nand U4621 (N_4621,N_4215,N_4069);
and U4622 (N_4622,N_4401,N_4388);
nand U4623 (N_4623,N_4344,N_4140);
and U4624 (N_4624,N_4014,N_4068);
and U4625 (N_4625,N_4370,N_4442);
and U4626 (N_4626,N_4114,N_4347);
or U4627 (N_4627,N_4023,N_4213);
nor U4628 (N_4628,N_4425,N_4285);
or U4629 (N_4629,N_4205,N_4073);
nor U4630 (N_4630,N_4312,N_4178);
nand U4631 (N_4631,N_4292,N_4204);
xnor U4632 (N_4632,N_4229,N_4357);
nand U4633 (N_4633,N_4135,N_4333);
xnor U4634 (N_4634,N_4256,N_4097);
nor U4635 (N_4635,N_4015,N_4417);
nand U4636 (N_4636,N_4089,N_4296);
nand U4637 (N_4637,N_4281,N_4095);
or U4638 (N_4638,N_4132,N_4200);
and U4639 (N_4639,N_4127,N_4125);
nand U4640 (N_4640,N_4402,N_4124);
nand U4641 (N_4641,N_4240,N_4173);
and U4642 (N_4642,N_4244,N_4342);
nand U4643 (N_4643,N_4491,N_4055);
and U4644 (N_4644,N_4148,N_4207);
and U4645 (N_4645,N_4051,N_4092);
nand U4646 (N_4646,N_4406,N_4123);
and U4647 (N_4647,N_4136,N_4378);
xor U4648 (N_4648,N_4295,N_4362);
xor U4649 (N_4649,N_4188,N_4042);
xnor U4650 (N_4650,N_4447,N_4018);
or U4651 (N_4651,N_4359,N_4460);
xor U4652 (N_4652,N_4195,N_4119);
xnor U4653 (N_4653,N_4156,N_4034);
xnor U4654 (N_4654,N_4374,N_4264);
or U4655 (N_4655,N_4120,N_4293);
and U4656 (N_4656,N_4469,N_4194);
nand U4657 (N_4657,N_4024,N_4087);
or U4658 (N_4658,N_4450,N_4043);
and U4659 (N_4659,N_4373,N_4419);
nor U4660 (N_4660,N_4396,N_4118);
nor U4661 (N_4661,N_4416,N_4323);
nor U4662 (N_4662,N_4307,N_4041);
xor U4663 (N_4663,N_4494,N_4389);
nand U4664 (N_4664,N_4322,N_4482);
nand U4665 (N_4665,N_4303,N_4368);
nor U4666 (N_4666,N_4044,N_4346);
nand U4667 (N_4667,N_4191,N_4066);
or U4668 (N_4668,N_4170,N_4316);
xor U4669 (N_4669,N_4395,N_4212);
nor U4670 (N_4670,N_4426,N_4035);
nand U4671 (N_4671,N_4380,N_4103);
nand U4672 (N_4672,N_4021,N_4288);
and U4673 (N_4673,N_4131,N_4452);
nor U4674 (N_4674,N_4499,N_4386);
and U4675 (N_4675,N_4106,N_4091);
or U4676 (N_4676,N_4275,N_4218);
or U4677 (N_4677,N_4165,N_4250);
nand U4678 (N_4678,N_4302,N_4269);
nand U4679 (N_4679,N_4283,N_4369);
nor U4680 (N_4680,N_4137,N_4446);
or U4681 (N_4681,N_4492,N_4062);
xor U4682 (N_4682,N_4181,N_4493);
nor U4683 (N_4683,N_4351,N_4016);
xnor U4684 (N_4684,N_4462,N_4400);
and U4685 (N_4685,N_4076,N_4480);
or U4686 (N_4686,N_4451,N_4046);
and U4687 (N_4687,N_4267,N_4448);
or U4688 (N_4688,N_4297,N_4090);
nand U4689 (N_4689,N_4029,N_4004);
or U4690 (N_4690,N_4002,N_4196);
xnor U4691 (N_4691,N_4053,N_4037);
or U4692 (N_4692,N_4164,N_4101);
or U4693 (N_4693,N_4299,N_4157);
nand U4694 (N_4694,N_4058,N_4025);
nor U4695 (N_4695,N_4353,N_4278);
or U4696 (N_4696,N_4099,N_4219);
or U4697 (N_4697,N_4129,N_4007);
xnor U4698 (N_4698,N_4143,N_4211);
nor U4699 (N_4699,N_4495,N_4235);
xnor U4700 (N_4700,N_4038,N_4405);
or U4701 (N_4701,N_4313,N_4167);
xor U4702 (N_4702,N_4072,N_4067);
xnor U4703 (N_4703,N_4291,N_4233);
nor U4704 (N_4704,N_4466,N_4300);
or U4705 (N_4705,N_4225,N_4472);
or U4706 (N_4706,N_4241,N_4441);
or U4707 (N_4707,N_4126,N_4110);
or U4708 (N_4708,N_4253,N_4252);
nor U4709 (N_4709,N_4305,N_4487);
nor U4710 (N_4710,N_4094,N_4202);
nor U4711 (N_4711,N_4047,N_4463);
xnor U4712 (N_4712,N_4483,N_4430);
and U4713 (N_4713,N_4324,N_4152);
xor U4714 (N_4714,N_4190,N_4459);
and U4715 (N_4715,N_4350,N_4319);
xor U4716 (N_4716,N_4471,N_4261);
nor U4717 (N_4717,N_4385,N_4160);
nor U4718 (N_4718,N_4177,N_4306);
or U4719 (N_4719,N_4198,N_4404);
nand U4720 (N_4720,N_4377,N_4104);
xor U4721 (N_4721,N_4308,N_4444);
and U4722 (N_4722,N_4128,N_4391);
or U4723 (N_4723,N_4439,N_4061);
nor U4724 (N_4724,N_4367,N_4418);
and U4725 (N_4725,N_4245,N_4340);
nand U4726 (N_4726,N_4242,N_4109);
xor U4727 (N_4727,N_4249,N_4217);
nor U4728 (N_4728,N_4498,N_4428);
xnor U4729 (N_4729,N_4497,N_4371);
xor U4730 (N_4730,N_4039,N_4052);
nand U4731 (N_4731,N_4227,N_4265);
nor U4732 (N_4732,N_4199,N_4327);
nor U4733 (N_4733,N_4082,N_4363);
or U4734 (N_4734,N_4222,N_4274);
and U4735 (N_4735,N_4427,N_4490);
nand U4736 (N_4736,N_4399,N_4122);
or U4737 (N_4737,N_4282,N_4193);
nand U4738 (N_4738,N_4019,N_4304);
nor U4739 (N_4739,N_4083,N_4478);
and U4740 (N_4740,N_4145,N_4175);
xor U4741 (N_4741,N_4263,N_4017);
xnor U4742 (N_4742,N_4468,N_4365);
nor U4743 (N_4743,N_4433,N_4349);
nor U4744 (N_4744,N_4301,N_4147);
or U4745 (N_4745,N_4184,N_4328);
or U4746 (N_4746,N_4236,N_4257);
xor U4747 (N_4747,N_4479,N_4185);
xor U4748 (N_4748,N_4315,N_4379);
nand U4749 (N_4749,N_4234,N_4376);
and U4750 (N_4750,N_4377,N_4251);
nor U4751 (N_4751,N_4486,N_4378);
xnor U4752 (N_4752,N_4243,N_4474);
or U4753 (N_4753,N_4144,N_4141);
nand U4754 (N_4754,N_4260,N_4401);
xnor U4755 (N_4755,N_4179,N_4194);
nor U4756 (N_4756,N_4183,N_4332);
and U4757 (N_4757,N_4277,N_4292);
and U4758 (N_4758,N_4234,N_4454);
or U4759 (N_4759,N_4329,N_4399);
nand U4760 (N_4760,N_4365,N_4033);
nor U4761 (N_4761,N_4460,N_4394);
and U4762 (N_4762,N_4300,N_4454);
nor U4763 (N_4763,N_4185,N_4335);
nand U4764 (N_4764,N_4286,N_4158);
and U4765 (N_4765,N_4394,N_4436);
and U4766 (N_4766,N_4057,N_4185);
and U4767 (N_4767,N_4222,N_4019);
nor U4768 (N_4768,N_4082,N_4210);
nor U4769 (N_4769,N_4074,N_4350);
and U4770 (N_4770,N_4030,N_4251);
xor U4771 (N_4771,N_4015,N_4411);
nor U4772 (N_4772,N_4034,N_4498);
xor U4773 (N_4773,N_4176,N_4334);
nand U4774 (N_4774,N_4047,N_4245);
and U4775 (N_4775,N_4123,N_4022);
or U4776 (N_4776,N_4377,N_4246);
and U4777 (N_4777,N_4355,N_4476);
xor U4778 (N_4778,N_4183,N_4351);
xor U4779 (N_4779,N_4429,N_4474);
nor U4780 (N_4780,N_4054,N_4015);
and U4781 (N_4781,N_4401,N_4430);
nand U4782 (N_4782,N_4168,N_4380);
or U4783 (N_4783,N_4081,N_4091);
and U4784 (N_4784,N_4109,N_4024);
nand U4785 (N_4785,N_4219,N_4174);
xor U4786 (N_4786,N_4367,N_4332);
and U4787 (N_4787,N_4264,N_4237);
nand U4788 (N_4788,N_4054,N_4451);
xnor U4789 (N_4789,N_4051,N_4141);
or U4790 (N_4790,N_4401,N_4286);
nor U4791 (N_4791,N_4447,N_4122);
and U4792 (N_4792,N_4154,N_4178);
xnor U4793 (N_4793,N_4113,N_4108);
nor U4794 (N_4794,N_4271,N_4153);
nor U4795 (N_4795,N_4357,N_4272);
nor U4796 (N_4796,N_4180,N_4019);
nand U4797 (N_4797,N_4085,N_4000);
nor U4798 (N_4798,N_4175,N_4037);
nand U4799 (N_4799,N_4116,N_4201);
nor U4800 (N_4800,N_4012,N_4291);
nand U4801 (N_4801,N_4001,N_4164);
or U4802 (N_4802,N_4242,N_4049);
and U4803 (N_4803,N_4231,N_4319);
and U4804 (N_4804,N_4241,N_4173);
nand U4805 (N_4805,N_4284,N_4069);
nor U4806 (N_4806,N_4466,N_4028);
nand U4807 (N_4807,N_4217,N_4304);
nand U4808 (N_4808,N_4117,N_4013);
and U4809 (N_4809,N_4027,N_4433);
and U4810 (N_4810,N_4324,N_4414);
xnor U4811 (N_4811,N_4254,N_4210);
xnor U4812 (N_4812,N_4251,N_4186);
or U4813 (N_4813,N_4321,N_4114);
xor U4814 (N_4814,N_4217,N_4380);
nor U4815 (N_4815,N_4188,N_4198);
nand U4816 (N_4816,N_4311,N_4133);
or U4817 (N_4817,N_4421,N_4270);
and U4818 (N_4818,N_4029,N_4226);
nand U4819 (N_4819,N_4490,N_4008);
nor U4820 (N_4820,N_4294,N_4366);
and U4821 (N_4821,N_4246,N_4008);
nand U4822 (N_4822,N_4006,N_4028);
xor U4823 (N_4823,N_4302,N_4225);
nand U4824 (N_4824,N_4250,N_4182);
xnor U4825 (N_4825,N_4403,N_4042);
xnor U4826 (N_4826,N_4332,N_4265);
or U4827 (N_4827,N_4057,N_4110);
nor U4828 (N_4828,N_4151,N_4047);
xnor U4829 (N_4829,N_4221,N_4218);
xor U4830 (N_4830,N_4152,N_4149);
or U4831 (N_4831,N_4172,N_4124);
or U4832 (N_4832,N_4440,N_4460);
xor U4833 (N_4833,N_4307,N_4304);
xor U4834 (N_4834,N_4025,N_4083);
nand U4835 (N_4835,N_4076,N_4149);
nand U4836 (N_4836,N_4021,N_4206);
xnor U4837 (N_4837,N_4101,N_4330);
nor U4838 (N_4838,N_4221,N_4342);
xnor U4839 (N_4839,N_4225,N_4027);
nand U4840 (N_4840,N_4044,N_4479);
or U4841 (N_4841,N_4179,N_4287);
nor U4842 (N_4842,N_4253,N_4181);
nand U4843 (N_4843,N_4253,N_4295);
or U4844 (N_4844,N_4238,N_4366);
nor U4845 (N_4845,N_4242,N_4087);
xnor U4846 (N_4846,N_4472,N_4085);
nor U4847 (N_4847,N_4288,N_4123);
or U4848 (N_4848,N_4133,N_4350);
xnor U4849 (N_4849,N_4495,N_4097);
and U4850 (N_4850,N_4201,N_4356);
and U4851 (N_4851,N_4233,N_4160);
and U4852 (N_4852,N_4127,N_4028);
nor U4853 (N_4853,N_4023,N_4125);
and U4854 (N_4854,N_4307,N_4214);
nand U4855 (N_4855,N_4241,N_4258);
nor U4856 (N_4856,N_4212,N_4249);
or U4857 (N_4857,N_4160,N_4277);
xnor U4858 (N_4858,N_4017,N_4269);
nand U4859 (N_4859,N_4498,N_4432);
and U4860 (N_4860,N_4372,N_4329);
and U4861 (N_4861,N_4258,N_4312);
xnor U4862 (N_4862,N_4416,N_4200);
xnor U4863 (N_4863,N_4442,N_4319);
or U4864 (N_4864,N_4410,N_4255);
and U4865 (N_4865,N_4398,N_4051);
nor U4866 (N_4866,N_4203,N_4220);
or U4867 (N_4867,N_4192,N_4263);
or U4868 (N_4868,N_4463,N_4343);
xnor U4869 (N_4869,N_4185,N_4237);
xor U4870 (N_4870,N_4311,N_4276);
xnor U4871 (N_4871,N_4232,N_4375);
and U4872 (N_4872,N_4225,N_4045);
or U4873 (N_4873,N_4328,N_4360);
nor U4874 (N_4874,N_4499,N_4058);
xor U4875 (N_4875,N_4234,N_4475);
nand U4876 (N_4876,N_4371,N_4490);
nand U4877 (N_4877,N_4134,N_4121);
nand U4878 (N_4878,N_4088,N_4403);
xor U4879 (N_4879,N_4279,N_4385);
nor U4880 (N_4880,N_4068,N_4055);
nor U4881 (N_4881,N_4061,N_4301);
nor U4882 (N_4882,N_4024,N_4186);
xor U4883 (N_4883,N_4211,N_4045);
nor U4884 (N_4884,N_4478,N_4374);
nand U4885 (N_4885,N_4217,N_4079);
nand U4886 (N_4886,N_4237,N_4189);
xnor U4887 (N_4887,N_4211,N_4332);
xnor U4888 (N_4888,N_4211,N_4457);
xor U4889 (N_4889,N_4419,N_4236);
and U4890 (N_4890,N_4162,N_4284);
and U4891 (N_4891,N_4065,N_4467);
or U4892 (N_4892,N_4024,N_4490);
or U4893 (N_4893,N_4143,N_4266);
nand U4894 (N_4894,N_4303,N_4268);
nand U4895 (N_4895,N_4201,N_4154);
nand U4896 (N_4896,N_4255,N_4126);
nand U4897 (N_4897,N_4084,N_4348);
xnor U4898 (N_4898,N_4491,N_4372);
xnor U4899 (N_4899,N_4118,N_4267);
or U4900 (N_4900,N_4250,N_4236);
xnor U4901 (N_4901,N_4439,N_4100);
and U4902 (N_4902,N_4481,N_4000);
or U4903 (N_4903,N_4308,N_4174);
or U4904 (N_4904,N_4442,N_4109);
nand U4905 (N_4905,N_4118,N_4019);
and U4906 (N_4906,N_4348,N_4490);
or U4907 (N_4907,N_4145,N_4030);
and U4908 (N_4908,N_4354,N_4163);
nor U4909 (N_4909,N_4029,N_4016);
or U4910 (N_4910,N_4321,N_4323);
nand U4911 (N_4911,N_4165,N_4403);
or U4912 (N_4912,N_4466,N_4331);
nand U4913 (N_4913,N_4155,N_4014);
and U4914 (N_4914,N_4023,N_4123);
nand U4915 (N_4915,N_4225,N_4217);
nor U4916 (N_4916,N_4062,N_4150);
nor U4917 (N_4917,N_4303,N_4029);
nand U4918 (N_4918,N_4099,N_4124);
nand U4919 (N_4919,N_4013,N_4245);
xor U4920 (N_4920,N_4424,N_4315);
and U4921 (N_4921,N_4424,N_4199);
nand U4922 (N_4922,N_4281,N_4497);
and U4923 (N_4923,N_4336,N_4140);
nand U4924 (N_4924,N_4089,N_4156);
or U4925 (N_4925,N_4330,N_4344);
nand U4926 (N_4926,N_4411,N_4190);
nand U4927 (N_4927,N_4059,N_4161);
nand U4928 (N_4928,N_4394,N_4162);
xor U4929 (N_4929,N_4288,N_4295);
and U4930 (N_4930,N_4064,N_4276);
xor U4931 (N_4931,N_4177,N_4133);
xnor U4932 (N_4932,N_4307,N_4246);
nand U4933 (N_4933,N_4469,N_4375);
and U4934 (N_4934,N_4455,N_4387);
or U4935 (N_4935,N_4305,N_4026);
nor U4936 (N_4936,N_4485,N_4492);
nand U4937 (N_4937,N_4442,N_4378);
and U4938 (N_4938,N_4312,N_4113);
xor U4939 (N_4939,N_4194,N_4175);
nand U4940 (N_4940,N_4010,N_4451);
nor U4941 (N_4941,N_4375,N_4351);
or U4942 (N_4942,N_4265,N_4282);
or U4943 (N_4943,N_4050,N_4147);
nor U4944 (N_4944,N_4081,N_4250);
nand U4945 (N_4945,N_4258,N_4485);
or U4946 (N_4946,N_4053,N_4117);
or U4947 (N_4947,N_4486,N_4155);
xnor U4948 (N_4948,N_4414,N_4378);
xnor U4949 (N_4949,N_4484,N_4032);
nor U4950 (N_4950,N_4374,N_4143);
and U4951 (N_4951,N_4179,N_4056);
xnor U4952 (N_4952,N_4199,N_4090);
nand U4953 (N_4953,N_4426,N_4045);
and U4954 (N_4954,N_4400,N_4123);
xor U4955 (N_4955,N_4044,N_4415);
nand U4956 (N_4956,N_4202,N_4368);
and U4957 (N_4957,N_4034,N_4496);
xnor U4958 (N_4958,N_4410,N_4361);
and U4959 (N_4959,N_4456,N_4215);
nand U4960 (N_4960,N_4164,N_4397);
or U4961 (N_4961,N_4088,N_4200);
or U4962 (N_4962,N_4391,N_4409);
nand U4963 (N_4963,N_4410,N_4127);
nor U4964 (N_4964,N_4153,N_4492);
xor U4965 (N_4965,N_4297,N_4187);
or U4966 (N_4966,N_4247,N_4031);
nand U4967 (N_4967,N_4066,N_4314);
xnor U4968 (N_4968,N_4432,N_4119);
nand U4969 (N_4969,N_4220,N_4130);
nor U4970 (N_4970,N_4244,N_4306);
xnor U4971 (N_4971,N_4138,N_4027);
or U4972 (N_4972,N_4492,N_4357);
nand U4973 (N_4973,N_4010,N_4295);
or U4974 (N_4974,N_4204,N_4269);
nand U4975 (N_4975,N_4106,N_4171);
or U4976 (N_4976,N_4256,N_4488);
or U4977 (N_4977,N_4099,N_4061);
xor U4978 (N_4978,N_4128,N_4057);
and U4979 (N_4979,N_4430,N_4477);
nand U4980 (N_4980,N_4063,N_4317);
nor U4981 (N_4981,N_4057,N_4277);
nand U4982 (N_4982,N_4410,N_4406);
xor U4983 (N_4983,N_4005,N_4271);
or U4984 (N_4984,N_4189,N_4493);
nor U4985 (N_4985,N_4197,N_4175);
nand U4986 (N_4986,N_4209,N_4231);
nand U4987 (N_4987,N_4395,N_4305);
nor U4988 (N_4988,N_4402,N_4198);
nor U4989 (N_4989,N_4265,N_4455);
nor U4990 (N_4990,N_4166,N_4009);
nand U4991 (N_4991,N_4093,N_4180);
xor U4992 (N_4992,N_4244,N_4030);
nand U4993 (N_4993,N_4402,N_4216);
or U4994 (N_4994,N_4119,N_4041);
xnor U4995 (N_4995,N_4174,N_4266);
nor U4996 (N_4996,N_4056,N_4174);
nand U4997 (N_4997,N_4337,N_4077);
or U4998 (N_4998,N_4118,N_4062);
nor U4999 (N_4999,N_4475,N_4210);
xor U5000 (N_5000,N_4621,N_4764);
nor U5001 (N_5001,N_4583,N_4554);
and U5002 (N_5002,N_4885,N_4972);
xor U5003 (N_5003,N_4745,N_4798);
xnor U5004 (N_5004,N_4556,N_4518);
nor U5005 (N_5005,N_4910,N_4855);
nand U5006 (N_5006,N_4647,N_4771);
nand U5007 (N_5007,N_4635,N_4586);
or U5008 (N_5008,N_4801,N_4630);
and U5009 (N_5009,N_4715,N_4723);
or U5010 (N_5010,N_4835,N_4736);
or U5011 (N_5011,N_4534,N_4645);
or U5012 (N_5012,N_4991,N_4914);
or U5013 (N_5013,N_4742,N_4578);
xnor U5014 (N_5014,N_4685,N_4956);
or U5015 (N_5015,N_4865,N_4516);
and U5016 (N_5016,N_4659,N_4670);
nor U5017 (N_5017,N_4967,N_4584);
nand U5018 (N_5018,N_4672,N_4821);
or U5019 (N_5019,N_4653,N_4733);
or U5020 (N_5020,N_4760,N_4531);
xnor U5021 (N_5021,N_4796,N_4544);
nor U5022 (N_5022,N_4523,N_4698);
and U5023 (N_5023,N_4548,N_4982);
or U5024 (N_5024,N_4740,N_4607);
and U5025 (N_5025,N_4935,N_4842);
and U5026 (N_5026,N_4528,N_4961);
xnor U5027 (N_5027,N_4900,N_4755);
and U5028 (N_5028,N_4758,N_4933);
or U5029 (N_5029,N_4674,N_4619);
and U5030 (N_5030,N_4952,N_4839);
nor U5031 (N_5031,N_4538,N_4934);
nand U5032 (N_5032,N_4943,N_4772);
nor U5033 (N_5033,N_4730,N_4996);
and U5034 (N_5034,N_4823,N_4515);
nand U5035 (N_5035,N_4638,N_4894);
nand U5036 (N_5036,N_4882,N_4896);
xor U5037 (N_5037,N_4696,N_4994);
nand U5038 (N_5038,N_4908,N_4721);
nor U5039 (N_5039,N_4564,N_4642);
nand U5040 (N_5040,N_4873,N_4596);
and U5041 (N_5041,N_4686,N_4646);
and U5042 (N_5042,N_4524,N_4840);
nor U5043 (N_5043,N_4716,N_4738);
and U5044 (N_5044,N_4520,N_4631);
xnor U5045 (N_5045,N_4566,N_4727);
nand U5046 (N_5046,N_4678,N_4939);
and U5047 (N_5047,N_4780,N_4773);
xor U5048 (N_5048,N_4907,N_4507);
or U5049 (N_5049,N_4699,N_4902);
or U5050 (N_5050,N_4567,N_4500);
nor U5051 (N_5051,N_4810,N_4866);
or U5052 (N_5052,N_4605,N_4924);
or U5053 (N_5053,N_4775,N_4676);
xnor U5054 (N_5054,N_4973,N_4981);
nor U5055 (N_5055,N_4948,N_4622);
xor U5056 (N_5056,N_4937,N_4750);
and U5057 (N_5057,N_4824,N_4802);
nor U5058 (N_5058,N_4711,N_4841);
or U5059 (N_5059,N_4774,N_4519);
and U5060 (N_5060,N_4641,N_4843);
and U5061 (N_5061,N_4884,N_4929);
and U5062 (N_5062,N_4502,N_4893);
and U5063 (N_5063,N_4787,N_4809);
nor U5064 (N_5064,N_4580,N_4541);
nor U5065 (N_5065,N_4992,N_4714);
xnor U5066 (N_5066,N_4833,N_4980);
and U5067 (N_5067,N_4606,N_4928);
nor U5068 (N_5068,N_4718,N_4664);
or U5069 (N_5069,N_4648,N_4610);
nor U5070 (N_5070,N_4526,N_4739);
and U5071 (N_5071,N_4741,N_4585);
or U5072 (N_5072,N_4511,N_4964);
xor U5073 (N_5073,N_4684,N_4504);
xnor U5074 (N_5074,N_4940,N_4673);
and U5075 (N_5075,N_4953,N_4747);
or U5076 (N_5076,N_4612,N_4765);
xor U5077 (N_5077,N_4633,N_4881);
and U5078 (N_5078,N_4751,N_4997);
and U5079 (N_5079,N_4789,N_4995);
nand U5080 (N_5080,N_4665,N_4555);
and U5081 (N_5081,N_4949,N_4691);
and U5082 (N_5082,N_4923,N_4588);
xnor U5083 (N_5083,N_4912,N_4752);
and U5084 (N_5084,N_4689,N_4532);
xnor U5085 (N_5085,N_4877,N_4743);
or U5086 (N_5086,N_4720,N_4827);
xnor U5087 (N_5087,N_4770,N_4667);
or U5088 (N_5088,N_4844,N_4959);
and U5089 (N_5089,N_4623,N_4592);
and U5090 (N_5090,N_4547,N_4792);
xor U5091 (N_5091,N_4918,N_4830);
nor U5092 (N_5092,N_4966,N_4581);
xor U5093 (N_5093,N_4977,N_4834);
or U5094 (N_5094,N_4620,N_4737);
nand U5095 (N_5095,N_4553,N_4651);
or U5096 (N_5096,N_4860,N_4875);
or U5097 (N_5097,N_4668,N_4955);
and U5098 (N_5098,N_4692,N_4861);
xnor U5099 (N_5099,N_4826,N_4944);
nand U5100 (N_5100,N_4671,N_4722);
xor U5101 (N_5101,N_4859,N_4890);
nand U5102 (N_5102,N_4536,N_4597);
xor U5103 (N_5103,N_4878,N_4962);
and U5104 (N_5104,N_4702,N_4958);
nor U5105 (N_5105,N_4763,N_4628);
or U5106 (N_5106,N_4549,N_4570);
xnor U5107 (N_5107,N_4811,N_4909);
xor U5108 (N_5108,N_4895,N_4899);
nor U5109 (N_5109,N_4617,N_4706);
nand U5110 (N_5110,N_4782,N_4726);
or U5111 (N_5111,N_4975,N_4540);
and U5112 (N_5112,N_4911,N_4946);
or U5113 (N_5113,N_4666,N_4757);
nand U5114 (N_5114,N_4938,N_4627);
and U5115 (N_5115,N_4563,N_4974);
or U5116 (N_5116,N_4998,N_4777);
nor U5117 (N_5117,N_4573,N_4710);
xor U5118 (N_5118,N_4954,N_4759);
nor U5119 (N_5119,N_4892,N_4695);
or U5120 (N_5120,N_4568,N_4779);
and U5121 (N_5121,N_4927,N_4569);
and U5122 (N_5122,N_4816,N_4897);
nor U5123 (N_5123,N_4529,N_4604);
or U5124 (N_5124,N_4626,N_4768);
or U5125 (N_5125,N_4703,N_4876);
or U5126 (N_5126,N_4886,N_4797);
or U5127 (N_5127,N_4986,N_4883);
nor U5128 (N_5128,N_4913,N_4799);
and U5129 (N_5129,N_4976,N_4784);
or U5130 (N_5130,N_4571,N_4945);
or U5131 (N_5131,N_4576,N_4558);
and U5132 (N_5132,N_4969,N_4871);
nor U5133 (N_5133,N_4906,N_4829);
nand U5134 (N_5134,N_4688,N_4679);
and U5135 (N_5135,N_4690,N_4624);
nand U5136 (N_5136,N_4560,N_4748);
nand U5137 (N_5137,N_4735,N_4904);
nor U5138 (N_5138,N_4550,N_4942);
and U5139 (N_5139,N_4815,N_4761);
nand U5140 (N_5140,N_4562,N_4947);
and U5141 (N_5141,N_4662,N_4932);
nor U5142 (N_5142,N_4599,N_4919);
xor U5143 (N_5143,N_4655,N_4926);
nand U5144 (N_5144,N_4514,N_4632);
or U5145 (N_5145,N_4543,N_4629);
xnor U5146 (N_5146,N_4870,N_4682);
xor U5147 (N_5147,N_4704,N_4832);
nand U5148 (N_5148,N_4533,N_4990);
and U5149 (N_5149,N_4616,N_4708);
and U5150 (N_5150,N_4851,N_4879);
or U5151 (N_5151,N_4634,N_4729);
xnor U5152 (N_5152,N_4746,N_4681);
nand U5153 (N_5153,N_4970,N_4791);
xnor U5154 (N_5154,N_4788,N_4577);
and U5155 (N_5155,N_4808,N_4591);
or U5156 (N_5156,N_4936,N_4505);
nand U5157 (N_5157,N_4931,N_4762);
and U5158 (N_5158,N_4978,N_4614);
nor U5159 (N_5159,N_4551,N_4579);
or U5160 (N_5160,N_4989,N_4650);
nor U5161 (N_5161,N_4805,N_4868);
and U5162 (N_5162,N_4968,N_4680);
nand U5163 (N_5163,N_4887,N_4734);
nand U5164 (N_5164,N_4595,N_4517);
or U5165 (N_5165,N_4603,N_4640);
or U5166 (N_5166,N_4687,N_4510);
nand U5167 (N_5167,N_4983,N_4921);
or U5168 (N_5168,N_4693,N_4786);
and U5169 (N_5169,N_4916,N_4888);
xor U5170 (N_5170,N_4863,N_4776);
and U5171 (N_5171,N_4643,N_4769);
and U5172 (N_5172,N_4661,N_4999);
xor U5173 (N_5173,N_4705,N_4660);
nor U5174 (N_5174,N_4766,N_4856);
or U5175 (N_5175,N_4854,N_4793);
and U5176 (N_5176,N_4767,N_4625);
and U5177 (N_5177,N_4867,N_4656);
nor U5178 (N_5178,N_4637,N_4901);
or U5179 (N_5179,N_4971,N_4806);
nor U5180 (N_5180,N_4898,N_4657);
and U5181 (N_5181,N_4542,N_4857);
or U5182 (N_5182,N_4828,N_4663);
xnor U5183 (N_5183,N_4869,N_4905);
xnor U5184 (N_5184,N_4838,N_4522);
nand U5185 (N_5185,N_4852,N_4930);
or U5186 (N_5186,N_4858,N_4535);
and U5187 (N_5187,N_4594,N_4920);
nand U5188 (N_5188,N_4988,N_4575);
xnor U5189 (N_5189,N_4864,N_4749);
nor U5190 (N_5190,N_4880,N_4552);
xnor U5191 (N_5191,N_4836,N_4589);
nand U5192 (N_5192,N_4611,N_4889);
xor U5193 (N_5193,N_4848,N_4963);
xor U5194 (N_5194,N_4506,N_4820);
nor U5195 (N_5195,N_4728,N_4781);
nand U5196 (N_5196,N_4756,N_4559);
xor U5197 (N_5197,N_4587,N_4600);
or U5198 (N_5198,N_4565,N_4818);
and U5199 (N_5199,N_4675,N_4965);
and U5200 (N_5200,N_4922,N_4850);
nand U5201 (N_5201,N_4545,N_4941);
nor U5202 (N_5202,N_4530,N_4778);
xor U5203 (N_5203,N_4669,N_4795);
xor U5204 (N_5204,N_4618,N_4574);
nor U5205 (N_5205,N_4987,N_4649);
nor U5206 (N_5206,N_4874,N_4639);
xor U5207 (N_5207,N_4803,N_4717);
xnor U5208 (N_5208,N_4993,N_4712);
or U5209 (N_5209,N_4754,N_4785);
and U5210 (N_5210,N_4593,N_4509);
nor U5211 (N_5211,N_4845,N_4501);
nor U5212 (N_5212,N_4694,N_4812);
xnor U5213 (N_5213,N_4615,N_4903);
and U5214 (N_5214,N_4512,N_4697);
xnor U5215 (N_5215,N_4725,N_4950);
or U5216 (N_5216,N_4525,N_4713);
nor U5217 (N_5217,N_4825,N_4521);
and U5218 (N_5218,N_4508,N_4794);
nand U5219 (N_5219,N_4783,N_4731);
or U5220 (N_5220,N_4701,N_4837);
xnor U5221 (N_5221,N_4813,N_4546);
nand U5222 (N_5222,N_4537,N_4853);
xor U5223 (N_5223,N_4557,N_4744);
nor U5224 (N_5224,N_4822,N_4819);
xnor U5225 (N_5225,N_4572,N_4644);
or U5226 (N_5226,N_4561,N_4539);
nand U5227 (N_5227,N_4636,N_4917);
and U5228 (N_5228,N_4658,N_4609);
and U5229 (N_5229,N_4915,N_4891);
xor U5230 (N_5230,N_4847,N_4700);
xnor U5231 (N_5231,N_4817,N_4790);
nor U5232 (N_5232,N_4979,N_4503);
xor U5233 (N_5233,N_4707,N_4862);
nor U5234 (N_5234,N_4872,N_4598);
or U5235 (N_5235,N_4652,N_4960);
xnor U5236 (N_5236,N_4601,N_4513);
or U5237 (N_5237,N_4800,N_4719);
or U5238 (N_5238,N_4724,N_4527);
nor U5239 (N_5239,N_4709,N_4677);
or U5240 (N_5240,N_4814,N_4846);
nor U5241 (N_5241,N_4654,N_4849);
nand U5242 (N_5242,N_4613,N_4582);
or U5243 (N_5243,N_4804,N_4925);
xnor U5244 (N_5244,N_4602,N_4753);
or U5245 (N_5245,N_4985,N_4951);
nor U5246 (N_5246,N_4608,N_4957);
nor U5247 (N_5247,N_4590,N_4683);
nand U5248 (N_5248,N_4831,N_4732);
or U5249 (N_5249,N_4984,N_4807);
and U5250 (N_5250,N_4915,N_4693);
or U5251 (N_5251,N_4573,N_4936);
nand U5252 (N_5252,N_4657,N_4578);
nor U5253 (N_5253,N_4972,N_4862);
nor U5254 (N_5254,N_4636,N_4922);
and U5255 (N_5255,N_4640,N_4563);
and U5256 (N_5256,N_4846,N_4832);
and U5257 (N_5257,N_4836,N_4597);
nor U5258 (N_5258,N_4703,N_4860);
nor U5259 (N_5259,N_4965,N_4872);
or U5260 (N_5260,N_4776,N_4567);
or U5261 (N_5261,N_4953,N_4559);
nand U5262 (N_5262,N_4837,N_4514);
xor U5263 (N_5263,N_4600,N_4669);
xnor U5264 (N_5264,N_4687,N_4638);
nand U5265 (N_5265,N_4512,N_4918);
nand U5266 (N_5266,N_4562,N_4976);
and U5267 (N_5267,N_4846,N_4587);
nor U5268 (N_5268,N_4827,N_4620);
nand U5269 (N_5269,N_4603,N_4921);
nor U5270 (N_5270,N_4958,N_4512);
nor U5271 (N_5271,N_4546,N_4541);
xor U5272 (N_5272,N_4544,N_4675);
xor U5273 (N_5273,N_4671,N_4628);
or U5274 (N_5274,N_4789,N_4618);
xor U5275 (N_5275,N_4507,N_4859);
or U5276 (N_5276,N_4808,N_4882);
nand U5277 (N_5277,N_4510,N_4852);
nand U5278 (N_5278,N_4630,N_4875);
and U5279 (N_5279,N_4646,N_4881);
nand U5280 (N_5280,N_4973,N_4752);
or U5281 (N_5281,N_4718,N_4562);
and U5282 (N_5282,N_4585,N_4945);
and U5283 (N_5283,N_4526,N_4768);
or U5284 (N_5284,N_4859,N_4719);
nor U5285 (N_5285,N_4733,N_4851);
nor U5286 (N_5286,N_4864,N_4909);
or U5287 (N_5287,N_4831,N_4763);
or U5288 (N_5288,N_4839,N_4949);
nand U5289 (N_5289,N_4916,N_4852);
and U5290 (N_5290,N_4960,N_4608);
nand U5291 (N_5291,N_4648,N_4708);
nor U5292 (N_5292,N_4527,N_4546);
nand U5293 (N_5293,N_4667,N_4601);
and U5294 (N_5294,N_4980,N_4882);
nand U5295 (N_5295,N_4912,N_4513);
xor U5296 (N_5296,N_4589,N_4850);
nor U5297 (N_5297,N_4980,N_4913);
or U5298 (N_5298,N_4520,N_4800);
xor U5299 (N_5299,N_4560,N_4900);
nor U5300 (N_5300,N_4882,N_4814);
xor U5301 (N_5301,N_4935,N_4703);
nor U5302 (N_5302,N_4762,N_4535);
or U5303 (N_5303,N_4752,N_4823);
nand U5304 (N_5304,N_4884,N_4718);
nand U5305 (N_5305,N_4699,N_4660);
xnor U5306 (N_5306,N_4753,N_4559);
and U5307 (N_5307,N_4528,N_4867);
and U5308 (N_5308,N_4518,N_4917);
xor U5309 (N_5309,N_4777,N_4714);
nand U5310 (N_5310,N_4984,N_4759);
nor U5311 (N_5311,N_4562,N_4641);
xor U5312 (N_5312,N_4697,N_4531);
or U5313 (N_5313,N_4664,N_4667);
and U5314 (N_5314,N_4519,N_4651);
or U5315 (N_5315,N_4733,N_4970);
nor U5316 (N_5316,N_4526,N_4730);
nand U5317 (N_5317,N_4793,N_4680);
or U5318 (N_5318,N_4768,N_4620);
nor U5319 (N_5319,N_4832,N_4617);
nand U5320 (N_5320,N_4679,N_4993);
nand U5321 (N_5321,N_4686,N_4696);
nor U5322 (N_5322,N_4668,N_4799);
nor U5323 (N_5323,N_4840,N_4922);
and U5324 (N_5324,N_4535,N_4803);
and U5325 (N_5325,N_4860,N_4905);
nand U5326 (N_5326,N_4562,N_4689);
and U5327 (N_5327,N_4575,N_4735);
nor U5328 (N_5328,N_4560,N_4599);
or U5329 (N_5329,N_4731,N_4897);
xor U5330 (N_5330,N_4514,N_4650);
xor U5331 (N_5331,N_4903,N_4790);
nor U5332 (N_5332,N_4613,N_4606);
or U5333 (N_5333,N_4723,N_4940);
or U5334 (N_5334,N_4925,N_4881);
or U5335 (N_5335,N_4525,N_4619);
nand U5336 (N_5336,N_4596,N_4799);
or U5337 (N_5337,N_4668,N_4692);
nand U5338 (N_5338,N_4876,N_4571);
nor U5339 (N_5339,N_4960,N_4766);
xor U5340 (N_5340,N_4891,N_4626);
nor U5341 (N_5341,N_4754,N_4643);
nor U5342 (N_5342,N_4748,N_4720);
and U5343 (N_5343,N_4910,N_4622);
and U5344 (N_5344,N_4729,N_4989);
xor U5345 (N_5345,N_4762,N_4794);
and U5346 (N_5346,N_4584,N_4618);
or U5347 (N_5347,N_4522,N_4750);
nor U5348 (N_5348,N_4777,N_4621);
nand U5349 (N_5349,N_4977,N_4710);
nand U5350 (N_5350,N_4665,N_4709);
xor U5351 (N_5351,N_4565,N_4518);
or U5352 (N_5352,N_4598,N_4911);
nor U5353 (N_5353,N_4577,N_4846);
or U5354 (N_5354,N_4955,N_4992);
xnor U5355 (N_5355,N_4943,N_4652);
xor U5356 (N_5356,N_4910,N_4531);
nor U5357 (N_5357,N_4963,N_4968);
nand U5358 (N_5358,N_4738,N_4704);
and U5359 (N_5359,N_4594,N_4527);
nand U5360 (N_5360,N_4689,N_4826);
xor U5361 (N_5361,N_4591,N_4593);
and U5362 (N_5362,N_4540,N_4657);
nor U5363 (N_5363,N_4817,N_4912);
nand U5364 (N_5364,N_4679,N_4666);
nand U5365 (N_5365,N_4643,N_4987);
or U5366 (N_5366,N_4675,N_4543);
or U5367 (N_5367,N_4509,N_4640);
nor U5368 (N_5368,N_4752,N_4697);
nand U5369 (N_5369,N_4756,N_4584);
or U5370 (N_5370,N_4968,N_4694);
xnor U5371 (N_5371,N_4950,N_4745);
or U5372 (N_5372,N_4931,N_4969);
and U5373 (N_5373,N_4747,N_4565);
and U5374 (N_5374,N_4876,N_4934);
and U5375 (N_5375,N_4674,N_4828);
nand U5376 (N_5376,N_4816,N_4887);
and U5377 (N_5377,N_4908,N_4591);
and U5378 (N_5378,N_4578,N_4913);
or U5379 (N_5379,N_4939,N_4587);
and U5380 (N_5380,N_4945,N_4972);
xor U5381 (N_5381,N_4792,N_4700);
xor U5382 (N_5382,N_4887,N_4648);
nor U5383 (N_5383,N_4814,N_4566);
nor U5384 (N_5384,N_4818,N_4705);
xnor U5385 (N_5385,N_4978,N_4814);
nor U5386 (N_5386,N_4815,N_4925);
nor U5387 (N_5387,N_4905,N_4809);
or U5388 (N_5388,N_4644,N_4954);
nor U5389 (N_5389,N_4787,N_4794);
and U5390 (N_5390,N_4944,N_4577);
nor U5391 (N_5391,N_4847,N_4684);
nor U5392 (N_5392,N_4982,N_4701);
nor U5393 (N_5393,N_4636,N_4862);
or U5394 (N_5394,N_4771,N_4906);
and U5395 (N_5395,N_4879,N_4977);
nor U5396 (N_5396,N_4819,N_4554);
or U5397 (N_5397,N_4864,N_4586);
and U5398 (N_5398,N_4642,N_4740);
nand U5399 (N_5399,N_4580,N_4979);
nand U5400 (N_5400,N_4734,N_4500);
and U5401 (N_5401,N_4806,N_4815);
and U5402 (N_5402,N_4514,N_4706);
nor U5403 (N_5403,N_4583,N_4748);
xor U5404 (N_5404,N_4865,N_4980);
or U5405 (N_5405,N_4746,N_4677);
and U5406 (N_5406,N_4657,N_4512);
xnor U5407 (N_5407,N_4925,N_4613);
xnor U5408 (N_5408,N_4533,N_4788);
and U5409 (N_5409,N_4946,N_4784);
or U5410 (N_5410,N_4530,N_4603);
xnor U5411 (N_5411,N_4835,N_4747);
nand U5412 (N_5412,N_4781,N_4777);
nor U5413 (N_5413,N_4729,N_4638);
nor U5414 (N_5414,N_4629,N_4715);
or U5415 (N_5415,N_4791,N_4922);
xnor U5416 (N_5416,N_4630,N_4771);
nor U5417 (N_5417,N_4709,N_4990);
xnor U5418 (N_5418,N_4635,N_4913);
and U5419 (N_5419,N_4709,N_4514);
xnor U5420 (N_5420,N_4619,N_4663);
nor U5421 (N_5421,N_4607,N_4645);
xor U5422 (N_5422,N_4559,N_4629);
or U5423 (N_5423,N_4967,N_4935);
nor U5424 (N_5424,N_4990,N_4969);
nand U5425 (N_5425,N_4781,N_4725);
xor U5426 (N_5426,N_4830,N_4712);
or U5427 (N_5427,N_4715,N_4895);
and U5428 (N_5428,N_4691,N_4761);
nand U5429 (N_5429,N_4727,N_4792);
nand U5430 (N_5430,N_4945,N_4750);
or U5431 (N_5431,N_4848,N_4744);
xnor U5432 (N_5432,N_4605,N_4721);
nand U5433 (N_5433,N_4746,N_4806);
xnor U5434 (N_5434,N_4787,N_4667);
nor U5435 (N_5435,N_4758,N_4584);
and U5436 (N_5436,N_4968,N_4979);
nand U5437 (N_5437,N_4917,N_4655);
and U5438 (N_5438,N_4751,N_4965);
nand U5439 (N_5439,N_4560,N_4920);
nor U5440 (N_5440,N_4730,N_4900);
or U5441 (N_5441,N_4598,N_4720);
and U5442 (N_5442,N_4696,N_4551);
nor U5443 (N_5443,N_4552,N_4625);
xor U5444 (N_5444,N_4553,N_4876);
or U5445 (N_5445,N_4895,N_4615);
and U5446 (N_5446,N_4510,N_4679);
nand U5447 (N_5447,N_4647,N_4684);
nand U5448 (N_5448,N_4632,N_4943);
nor U5449 (N_5449,N_4870,N_4978);
nand U5450 (N_5450,N_4678,N_4876);
and U5451 (N_5451,N_4616,N_4513);
or U5452 (N_5452,N_4993,N_4802);
nand U5453 (N_5453,N_4783,N_4909);
or U5454 (N_5454,N_4624,N_4721);
nor U5455 (N_5455,N_4956,N_4783);
nor U5456 (N_5456,N_4926,N_4607);
and U5457 (N_5457,N_4874,N_4876);
nand U5458 (N_5458,N_4564,N_4569);
xor U5459 (N_5459,N_4761,N_4828);
and U5460 (N_5460,N_4603,N_4887);
and U5461 (N_5461,N_4773,N_4833);
xnor U5462 (N_5462,N_4570,N_4657);
or U5463 (N_5463,N_4909,N_4838);
xor U5464 (N_5464,N_4882,N_4937);
nand U5465 (N_5465,N_4664,N_4700);
nor U5466 (N_5466,N_4727,N_4790);
or U5467 (N_5467,N_4512,N_4682);
xor U5468 (N_5468,N_4964,N_4822);
or U5469 (N_5469,N_4818,N_4860);
and U5470 (N_5470,N_4616,N_4518);
and U5471 (N_5471,N_4993,N_4550);
nor U5472 (N_5472,N_4780,N_4747);
nor U5473 (N_5473,N_4652,N_4621);
xor U5474 (N_5474,N_4647,N_4882);
xor U5475 (N_5475,N_4877,N_4732);
nand U5476 (N_5476,N_4869,N_4671);
or U5477 (N_5477,N_4698,N_4924);
or U5478 (N_5478,N_4611,N_4701);
nor U5479 (N_5479,N_4652,N_4538);
nor U5480 (N_5480,N_4565,N_4585);
and U5481 (N_5481,N_4528,N_4890);
xnor U5482 (N_5482,N_4952,N_4768);
nand U5483 (N_5483,N_4755,N_4983);
or U5484 (N_5484,N_4837,N_4902);
or U5485 (N_5485,N_4660,N_4609);
and U5486 (N_5486,N_4985,N_4509);
and U5487 (N_5487,N_4732,N_4674);
nor U5488 (N_5488,N_4546,N_4701);
and U5489 (N_5489,N_4648,N_4778);
nor U5490 (N_5490,N_4810,N_4695);
nor U5491 (N_5491,N_4807,N_4812);
and U5492 (N_5492,N_4641,N_4850);
xnor U5493 (N_5493,N_4843,N_4816);
xnor U5494 (N_5494,N_4713,N_4995);
and U5495 (N_5495,N_4959,N_4968);
xor U5496 (N_5496,N_4814,N_4994);
or U5497 (N_5497,N_4562,N_4598);
and U5498 (N_5498,N_4972,N_4649);
and U5499 (N_5499,N_4913,N_4961);
nand U5500 (N_5500,N_5238,N_5050);
or U5501 (N_5501,N_5466,N_5119);
xor U5502 (N_5502,N_5024,N_5318);
and U5503 (N_5503,N_5038,N_5243);
or U5504 (N_5504,N_5230,N_5492);
nand U5505 (N_5505,N_5478,N_5116);
nor U5506 (N_5506,N_5097,N_5216);
nand U5507 (N_5507,N_5013,N_5272);
nand U5508 (N_5508,N_5113,N_5017);
and U5509 (N_5509,N_5093,N_5254);
nor U5510 (N_5510,N_5134,N_5086);
xor U5511 (N_5511,N_5154,N_5208);
or U5512 (N_5512,N_5162,N_5486);
or U5513 (N_5513,N_5153,N_5413);
nand U5514 (N_5514,N_5020,N_5346);
and U5515 (N_5515,N_5055,N_5166);
nand U5516 (N_5516,N_5372,N_5213);
xnor U5517 (N_5517,N_5395,N_5256);
nand U5518 (N_5518,N_5267,N_5355);
nand U5519 (N_5519,N_5033,N_5091);
nor U5520 (N_5520,N_5464,N_5306);
nor U5521 (N_5521,N_5049,N_5034);
nor U5522 (N_5522,N_5239,N_5235);
nand U5523 (N_5523,N_5224,N_5269);
nand U5524 (N_5524,N_5392,N_5291);
nand U5525 (N_5525,N_5487,N_5202);
and U5526 (N_5526,N_5427,N_5410);
xor U5527 (N_5527,N_5484,N_5350);
nor U5528 (N_5528,N_5001,N_5477);
or U5529 (N_5529,N_5152,N_5102);
nor U5530 (N_5530,N_5348,N_5449);
nor U5531 (N_5531,N_5402,N_5356);
or U5532 (N_5532,N_5136,N_5359);
or U5533 (N_5533,N_5457,N_5183);
nand U5534 (N_5534,N_5138,N_5388);
or U5535 (N_5535,N_5149,N_5083);
and U5536 (N_5536,N_5416,N_5014);
xor U5537 (N_5537,N_5336,N_5377);
xnor U5538 (N_5538,N_5035,N_5100);
and U5539 (N_5539,N_5178,N_5022);
or U5540 (N_5540,N_5491,N_5191);
nand U5541 (N_5541,N_5173,N_5098);
nor U5542 (N_5542,N_5005,N_5171);
or U5543 (N_5543,N_5276,N_5419);
and U5544 (N_5544,N_5205,N_5160);
nor U5545 (N_5545,N_5234,N_5462);
nor U5546 (N_5546,N_5112,N_5441);
and U5547 (N_5547,N_5360,N_5385);
and U5548 (N_5548,N_5233,N_5000);
and U5549 (N_5549,N_5253,N_5414);
or U5550 (N_5550,N_5303,N_5424);
nand U5551 (N_5551,N_5222,N_5431);
or U5552 (N_5552,N_5244,N_5417);
nor U5553 (N_5553,N_5320,N_5255);
nor U5554 (N_5554,N_5494,N_5274);
and U5555 (N_5555,N_5258,N_5029);
or U5556 (N_5556,N_5064,N_5271);
nor U5557 (N_5557,N_5193,N_5241);
xor U5558 (N_5558,N_5296,N_5032);
and U5559 (N_5559,N_5023,N_5314);
and U5560 (N_5560,N_5015,N_5174);
and U5561 (N_5561,N_5011,N_5293);
or U5562 (N_5562,N_5054,N_5135);
and U5563 (N_5563,N_5219,N_5435);
nand U5564 (N_5564,N_5245,N_5057);
and U5565 (N_5565,N_5075,N_5073);
xnor U5566 (N_5566,N_5027,N_5079);
and U5567 (N_5567,N_5378,N_5109);
or U5568 (N_5568,N_5483,N_5123);
xor U5569 (N_5569,N_5374,N_5268);
or U5570 (N_5570,N_5406,N_5009);
xor U5571 (N_5571,N_5010,N_5369);
nand U5572 (N_5572,N_5430,N_5217);
and U5573 (N_5573,N_5184,N_5480);
nor U5574 (N_5574,N_5115,N_5396);
or U5575 (N_5575,N_5329,N_5006);
and U5576 (N_5576,N_5150,N_5042);
nand U5577 (N_5577,N_5158,N_5052);
and U5578 (N_5578,N_5056,N_5349);
nor U5579 (N_5579,N_5315,N_5401);
nand U5580 (N_5580,N_5190,N_5141);
nand U5581 (N_5581,N_5436,N_5283);
nand U5582 (N_5582,N_5422,N_5469);
and U5583 (N_5583,N_5428,N_5311);
xnor U5584 (N_5584,N_5447,N_5188);
or U5585 (N_5585,N_5408,N_5361);
or U5586 (N_5586,N_5096,N_5232);
and U5587 (N_5587,N_5442,N_5351);
or U5588 (N_5588,N_5357,N_5316);
and U5589 (N_5589,N_5493,N_5117);
and U5590 (N_5590,N_5026,N_5110);
xor U5591 (N_5591,N_5310,N_5328);
and U5592 (N_5592,N_5265,N_5111);
xor U5593 (N_5593,N_5227,N_5437);
nor U5594 (N_5594,N_5454,N_5037);
nor U5595 (N_5595,N_5168,N_5161);
or U5596 (N_5596,N_5394,N_5334);
nand U5597 (N_5597,N_5330,N_5308);
nor U5598 (N_5598,N_5352,N_5434);
nand U5599 (N_5599,N_5312,N_5445);
nor U5600 (N_5600,N_5105,N_5016);
and U5601 (N_5601,N_5278,N_5209);
nor U5602 (N_5602,N_5400,N_5423);
or U5603 (N_5603,N_5313,N_5081);
nand U5604 (N_5604,N_5249,N_5072);
nor U5605 (N_5605,N_5210,N_5327);
xnor U5606 (N_5606,N_5365,N_5326);
xor U5607 (N_5607,N_5182,N_5008);
xnor U5608 (N_5608,N_5192,N_5467);
nor U5609 (N_5609,N_5286,N_5139);
and U5610 (N_5610,N_5066,N_5455);
or U5611 (N_5611,N_5087,N_5175);
nand U5612 (N_5612,N_5304,N_5155);
xor U5613 (N_5613,N_5387,N_5472);
and U5614 (N_5614,N_5067,N_5197);
nand U5615 (N_5615,N_5187,N_5439);
or U5616 (N_5616,N_5137,N_5379);
xor U5617 (N_5617,N_5498,N_5172);
nand U5618 (N_5618,N_5131,N_5220);
xor U5619 (N_5619,N_5363,N_5186);
nor U5620 (N_5620,N_5089,N_5475);
nand U5621 (N_5621,N_5405,N_5198);
xor U5622 (N_5622,N_5065,N_5176);
or U5623 (N_5623,N_5163,N_5383);
or U5624 (N_5624,N_5384,N_5031);
xnor U5625 (N_5625,N_5353,N_5450);
xnor U5626 (N_5626,N_5221,N_5021);
nand U5627 (N_5627,N_5456,N_5451);
or U5628 (N_5628,N_5063,N_5339);
and U5629 (N_5629,N_5389,N_5459);
and U5630 (N_5630,N_5252,N_5370);
nand U5631 (N_5631,N_5332,N_5180);
and U5632 (N_5632,N_5298,N_5092);
and U5633 (N_5633,N_5277,N_5046);
nor U5634 (N_5634,N_5465,N_5266);
or U5635 (N_5635,N_5068,N_5479);
nor U5636 (N_5636,N_5040,N_5094);
and U5637 (N_5637,N_5047,N_5200);
nand U5638 (N_5638,N_5151,N_5347);
nand U5639 (N_5639,N_5364,N_5362);
and U5640 (N_5640,N_5130,N_5251);
xnor U5641 (N_5641,N_5125,N_5126);
xor U5642 (N_5642,N_5028,N_5390);
or U5643 (N_5643,N_5421,N_5319);
xor U5644 (N_5644,N_5212,N_5165);
or U5645 (N_5645,N_5043,N_5289);
nor U5646 (N_5646,N_5107,N_5474);
xnor U5647 (N_5647,N_5211,N_5382);
xnor U5648 (N_5648,N_5425,N_5167);
and U5649 (N_5649,N_5106,N_5061);
or U5650 (N_5650,N_5337,N_5203);
or U5651 (N_5651,N_5146,N_5003);
xnor U5652 (N_5652,N_5285,N_5367);
nor U5653 (N_5653,N_5380,N_5452);
or U5654 (N_5654,N_5129,N_5341);
nor U5655 (N_5655,N_5403,N_5460);
or U5656 (N_5656,N_5263,N_5275);
and U5657 (N_5657,N_5489,N_5124);
and U5658 (N_5658,N_5012,N_5189);
nand U5659 (N_5659,N_5307,N_5019);
nor U5660 (N_5660,N_5261,N_5273);
and U5661 (N_5661,N_5411,N_5103);
nand U5662 (N_5662,N_5331,N_5397);
nand U5663 (N_5663,N_5077,N_5280);
nand U5664 (N_5664,N_5438,N_5342);
nand U5665 (N_5665,N_5407,N_5053);
and U5666 (N_5666,N_5426,N_5458);
xnor U5667 (N_5667,N_5170,N_5247);
or U5668 (N_5668,N_5481,N_5444);
xor U5669 (N_5669,N_5488,N_5287);
xor U5670 (N_5670,N_5470,N_5440);
nand U5671 (N_5671,N_5371,N_5099);
nor U5672 (N_5672,N_5322,N_5195);
or U5673 (N_5673,N_5071,N_5448);
nand U5674 (N_5674,N_5340,N_5108);
nor U5675 (N_5675,N_5299,N_5157);
nand U5676 (N_5676,N_5386,N_5433);
or U5677 (N_5677,N_5338,N_5218);
nand U5678 (N_5678,N_5294,N_5080);
nor U5679 (N_5679,N_5366,N_5499);
xnor U5680 (N_5680,N_5250,N_5122);
nor U5681 (N_5681,N_5084,N_5468);
and U5682 (N_5682,N_5301,N_5144);
or U5683 (N_5683,N_5104,N_5282);
or U5684 (N_5684,N_5143,N_5264);
nand U5685 (N_5685,N_5226,N_5240);
and U5686 (N_5686,N_5132,N_5398);
or U5687 (N_5687,N_5044,N_5323);
or U5688 (N_5688,N_5194,N_5058);
or U5689 (N_5689,N_5145,N_5295);
xnor U5690 (N_5690,N_5185,N_5085);
or U5691 (N_5691,N_5300,N_5181);
or U5692 (N_5692,N_5030,N_5215);
nand U5693 (N_5693,N_5207,N_5078);
nand U5694 (N_5694,N_5476,N_5048);
nand U5695 (N_5695,N_5127,N_5159);
and U5696 (N_5696,N_5090,N_5461);
and U5697 (N_5697,N_5399,N_5169);
nor U5698 (N_5698,N_5305,N_5004);
or U5699 (N_5699,N_5120,N_5018);
xor U5700 (N_5700,N_5497,N_5281);
nand U5701 (N_5701,N_5196,N_5375);
nand U5702 (N_5702,N_5335,N_5074);
and U5703 (N_5703,N_5242,N_5237);
and U5704 (N_5704,N_5095,N_5333);
xnor U5705 (N_5705,N_5420,N_5373);
nand U5706 (N_5706,N_5325,N_5345);
nand U5707 (N_5707,N_5446,N_5025);
xnor U5708 (N_5708,N_5412,N_5344);
nand U5709 (N_5709,N_5060,N_5236);
nor U5710 (N_5710,N_5453,N_5041);
nor U5711 (N_5711,N_5381,N_5393);
nor U5712 (N_5712,N_5292,N_5270);
nor U5713 (N_5713,N_5404,N_5432);
nand U5714 (N_5714,N_5260,N_5229);
or U5715 (N_5715,N_5045,N_5101);
nor U5716 (N_5716,N_5070,N_5463);
and U5717 (N_5717,N_5214,N_5206);
xnor U5718 (N_5718,N_5290,N_5496);
and U5719 (N_5719,N_5199,N_5223);
and U5720 (N_5720,N_5490,N_5302);
nand U5721 (N_5721,N_5179,N_5391);
or U5722 (N_5722,N_5059,N_5088);
nor U5723 (N_5723,N_5177,N_5118);
xor U5724 (N_5724,N_5482,N_5443);
and U5725 (N_5725,N_5204,N_5262);
nand U5726 (N_5726,N_5036,N_5354);
nand U5727 (N_5727,N_5473,N_5002);
or U5728 (N_5728,N_5164,N_5259);
xor U5729 (N_5729,N_5309,N_5121);
and U5730 (N_5730,N_5257,N_5429);
nand U5731 (N_5731,N_5082,N_5343);
or U5732 (N_5732,N_5368,N_5114);
nor U5733 (N_5733,N_5228,N_5076);
or U5734 (N_5734,N_5133,N_5051);
and U5735 (N_5735,N_5485,N_5495);
xor U5736 (N_5736,N_5288,N_5358);
or U5737 (N_5737,N_5324,N_5248);
nor U5738 (N_5738,N_5471,N_5297);
and U5739 (N_5739,N_5279,N_5140);
xor U5740 (N_5740,N_5321,N_5156);
nor U5741 (N_5741,N_5376,N_5201);
nand U5742 (N_5742,N_5225,N_5409);
nand U5743 (N_5743,N_5317,N_5246);
or U5744 (N_5744,N_5231,N_5142);
and U5745 (N_5745,N_5039,N_5148);
nand U5746 (N_5746,N_5415,N_5062);
nand U5747 (N_5747,N_5069,N_5418);
nor U5748 (N_5748,N_5007,N_5284);
nor U5749 (N_5749,N_5128,N_5147);
xor U5750 (N_5750,N_5432,N_5176);
and U5751 (N_5751,N_5466,N_5098);
and U5752 (N_5752,N_5024,N_5415);
and U5753 (N_5753,N_5017,N_5046);
and U5754 (N_5754,N_5104,N_5142);
or U5755 (N_5755,N_5229,N_5487);
or U5756 (N_5756,N_5214,N_5035);
xnor U5757 (N_5757,N_5047,N_5382);
nand U5758 (N_5758,N_5045,N_5084);
nand U5759 (N_5759,N_5070,N_5377);
and U5760 (N_5760,N_5012,N_5218);
or U5761 (N_5761,N_5140,N_5346);
nor U5762 (N_5762,N_5371,N_5205);
nand U5763 (N_5763,N_5441,N_5005);
and U5764 (N_5764,N_5008,N_5223);
xor U5765 (N_5765,N_5007,N_5088);
or U5766 (N_5766,N_5370,N_5016);
xor U5767 (N_5767,N_5194,N_5112);
and U5768 (N_5768,N_5424,N_5127);
nor U5769 (N_5769,N_5003,N_5414);
nor U5770 (N_5770,N_5113,N_5491);
and U5771 (N_5771,N_5315,N_5198);
nand U5772 (N_5772,N_5194,N_5254);
or U5773 (N_5773,N_5450,N_5453);
nor U5774 (N_5774,N_5381,N_5330);
xor U5775 (N_5775,N_5331,N_5361);
and U5776 (N_5776,N_5095,N_5190);
or U5777 (N_5777,N_5374,N_5326);
xor U5778 (N_5778,N_5135,N_5410);
or U5779 (N_5779,N_5196,N_5109);
and U5780 (N_5780,N_5191,N_5082);
xnor U5781 (N_5781,N_5180,N_5428);
nor U5782 (N_5782,N_5357,N_5414);
and U5783 (N_5783,N_5167,N_5031);
and U5784 (N_5784,N_5171,N_5413);
nand U5785 (N_5785,N_5181,N_5049);
and U5786 (N_5786,N_5484,N_5430);
and U5787 (N_5787,N_5182,N_5215);
xnor U5788 (N_5788,N_5255,N_5092);
and U5789 (N_5789,N_5022,N_5369);
xor U5790 (N_5790,N_5295,N_5256);
or U5791 (N_5791,N_5257,N_5112);
or U5792 (N_5792,N_5342,N_5287);
nand U5793 (N_5793,N_5434,N_5067);
and U5794 (N_5794,N_5165,N_5155);
or U5795 (N_5795,N_5233,N_5066);
nor U5796 (N_5796,N_5156,N_5282);
nor U5797 (N_5797,N_5017,N_5188);
xnor U5798 (N_5798,N_5337,N_5232);
nor U5799 (N_5799,N_5286,N_5492);
nand U5800 (N_5800,N_5147,N_5432);
and U5801 (N_5801,N_5441,N_5438);
xnor U5802 (N_5802,N_5219,N_5171);
xnor U5803 (N_5803,N_5157,N_5166);
xor U5804 (N_5804,N_5025,N_5011);
nand U5805 (N_5805,N_5131,N_5122);
or U5806 (N_5806,N_5344,N_5013);
nor U5807 (N_5807,N_5232,N_5117);
nand U5808 (N_5808,N_5002,N_5332);
nor U5809 (N_5809,N_5365,N_5255);
and U5810 (N_5810,N_5132,N_5074);
nor U5811 (N_5811,N_5350,N_5326);
nand U5812 (N_5812,N_5044,N_5455);
xnor U5813 (N_5813,N_5359,N_5385);
and U5814 (N_5814,N_5053,N_5017);
nor U5815 (N_5815,N_5208,N_5145);
or U5816 (N_5816,N_5399,N_5203);
nand U5817 (N_5817,N_5448,N_5311);
xnor U5818 (N_5818,N_5211,N_5006);
nand U5819 (N_5819,N_5332,N_5418);
xnor U5820 (N_5820,N_5212,N_5381);
nor U5821 (N_5821,N_5026,N_5377);
and U5822 (N_5822,N_5120,N_5089);
nand U5823 (N_5823,N_5376,N_5151);
and U5824 (N_5824,N_5435,N_5109);
and U5825 (N_5825,N_5463,N_5146);
or U5826 (N_5826,N_5126,N_5476);
xor U5827 (N_5827,N_5402,N_5315);
nand U5828 (N_5828,N_5214,N_5191);
and U5829 (N_5829,N_5266,N_5191);
nor U5830 (N_5830,N_5182,N_5108);
or U5831 (N_5831,N_5174,N_5060);
and U5832 (N_5832,N_5255,N_5237);
xnor U5833 (N_5833,N_5328,N_5199);
nand U5834 (N_5834,N_5400,N_5277);
nor U5835 (N_5835,N_5301,N_5260);
nand U5836 (N_5836,N_5123,N_5304);
nor U5837 (N_5837,N_5356,N_5410);
nand U5838 (N_5838,N_5118,N_5035);
nor U5839 (N_5839,N_5274,N_5280);
and U5840 (N_5840,N_5364,N_5116);
or U5841 (N_5841,N_5175,N_5165);
nand U5842 (N_5842,N_5246,N_5382);
xor U5843 (N_5843,N_5031,N_5350);
and U5844 (N_5844,N_5047,N_5022);
nor U5845 (N_5845,N_5444,N_5330);
nor U5846 (N_5846,N_5357,N_5269);
nor U5847 (N_5847,N_5424,N_5356);
xor U5848 (N_5848,N_5285,N_5132);
xnor U5849 (N_5849,N_5003,N_5080);
or U5850 (N_5850,N_5383,N_5386);
xnor U5851 (N_5851,N_5318,N_5433);
or U5852 (N_5852,N_5476,N_5070);
nor U5853 (N_5853,N_5495,N_5108);
nor U5854 (N_5854,N_5155,N_5347);
nor U5855 (N_5855,N_5142,N_5030);
nand U5856 (N_5856,N_5025,N_5498);
or U5857 (N_5857,N_5270,N_5472);
xnor U5858 (N_5858,N_5153,N_5243);
xnor U5859 (N_5859,N_5348,N_5124);
nor U5860 (N_5860,N_5440,N_5022);
or U5861 (N_5861,N_5209,N_5087);
xnor U5862 (N_5862,N_5320,N_5094);
and U5863 (N_5863,N_5349,N_5126);
nand U5864 (N_5864,N_5469,N_5382);
or U5865 (N_5865,N_5141,N_5101);
and U5866 (N_5866,N_5452,N_5168);
and U5867 (N_5867,N_5441,N_5478);
xnor U5868 (N_5868,N_5151,N_5277);
or U5869 (N_5869,N_5241,N_5218);
xor U5870 (N_5870,N_5013,N_5270);
or U5871 (N_5871,N_5109,N_5190);
nor U5872 (N_5872,N_5164,N_5160);
nand U5873 (N_5873,N_5167,N_5396);
and U5874 (N_5874,N_5021,N_5288);
nor U5875 (N_5875,N_5043,N_5353);
and U5876 (N_5876,N_5278,N_5160);
xnor U5877 (N_5877,N_5412,N_5050);
nor U5878 (N_5878,N_5098,N_5096);
xor U5879 (N_5879,N_5134,N_5078);
xnor U5880 (N_5880,N_5375,N_5420);
nor U5881 (N_5881,N_5374,N_5203);
xor U5882 (N_5882,N_5481,N_5416);
and U5883 (N_5883,N_5169,N_5442);
and U5884 (N_5884,N_5217,N_5318);
xor U5885 (N_5885,N_5269,N_5100);
or U5886 (N_5886,N_5004,N_5450);
xnor U5887 (N_5887,N_5191,N_5035);
nor U5888 (N_5888,N_5305,N_5484);
and U5889 (N_5889,N_5377,N_5031);
or U5890 (N_5890,N_5317,N_5260);
or U5891 (N_5891,N_5389,N_5029);
and U5892 (N_5892,N_5389,N_5101);
nand U5893 (N_5893,N_5348,N_5499);
nor U5894 (N_5894,N_5009,N_5031);
and U5895 (N_5895,N_5490,N_5140);
or U5896 (N_5896,N_5328,N_5213);
xor U5897 (N_5897,N_5162,N_5434);
nand U5898 (N_5898,N_5186,N_5145);
nand U5899 (N_5899,N_5402,N_5433);
or U5900 (N_5900,N_5453,N_5076);
xor U5901 (N_5901,N_5337,N_5390);
and U5902 (N_5902,N_5295,N_5023);
nand U5903 (N_5903,N_5098,N_5003);
and U5904 (N_5904,N_5298,N_5111);
and U5905 (N_5905,N_5340,N_5464);
xnor U5906 (N_5906,N_5236,N_5076);
xor U5907 (N_5907,N_5273,N_5310);
nand U5908 (N_5908,N_5357,N_5454);
nand U5909 (N_5909,N_5414,N_5463);
or U5910 (N_5910,N_5322,N_5237);
or U5911 (N_5911,N_5481,N_5147);
nor U5912 (N_5912,N_5208,N_5134);
nand U5913 (N_5913,N_5073,N_5030);
or U5914 (N_5914,N_5268,N_5390);
xor U5915 (N_5915,N_5398,N_5055);
xor U5916 (N_5916,N_5246,N_5482);
nor U5917 (N_5917,N_5122,N_5006);
nand U5918 (N_5918,N_5323,N_5319);
and U5919 (N_5919,N_5393,N_5152);
xor U5920 (N_5920,N_5263,N_5397);
nand U5921 (N_5921,N_5443,N_5228);
or U5922 (N_5922,N_5423,N_5316);
nand U5923 (N_5923,N_5124,N_5179);
or U5924 (N_5924,N_5235,N_5267);
or U5925 (N_5925,N_5458,N_5372);
nor U5926 (N_5926,N_5435,N_5112);
nand U5927 (N_5927,N_5041,N_5299);
nor U5928 (N_5928,N_5110,N_5424);
or U5929 (N_5929,N_5358,N_5173);
nor U5930 (N_5930,N_5311,N_5055);
nand U5931 (N_5931,N_5030,N_5184);
or U5932 (N_5932,N_5359,N_5197);
or U5933 (N_5933,N_5490,N_5308);
xor U5934 (N_5934,N_5326,N_5309);
nand U5935 (N_5935,N_5421,N_5177);
nor U5936 (N_5936,N_5109,N_5065);
nor U5937 (N_5937,N_5449,N_5275);
and U5938 (N_5938,N_5007,N_5077);
or U5939 (N_5939,N_5048,N_5014);
nand U5940 (N_5940,N_5056,N_5430);
nor U5941 (N_5941,N_5347,N_5174);
or U5942 (N_5942,N_5478,N_5470);
or U5943 (N_5943,N_5465,N_5109);
or U5944 (N_5944,N_5257,N_5215);
nor U5945 (N_5945,N_5033,N_5060);
and U5946 (N_5946,N_5306,N_5093);
nor U5947 (N_5947,N_5000,N_5307);
or U5948 (N_5948,N_5254,N_5079);
nor U5949 (N_5949,N_5142,N_5112);
xor U5950 (N_5950,N_5166,N_5253);
and U5951 (N_5951,N_5413,N_5161);
or U5952 (N_5952,N_5246,N_5022);
nand U5953 (N_5953,N_5420,N_5096);
nor U5954 (N_5954,N_5414,N_5170);
nor U5955 (N_5955,N_5197,N_5391);
or U5956 (N_5956,N_5158,N_5113);
and U5957 (N_5957,N_5107,N_5102);
or U5958 (N_5958,N_5398,N_5114);
and U5959 (N_5959,N_5120,N_5410);
and U5960 (N_5960,N_5190,N_5352);
nor U5961 (N_5961,N_5077,N_5011);
nand U5962 (N_5962,N_5027,N_5116);
or U5963 (N_5963,N_5059,N_5324);
xor U5964 (N_5964,N_5362,N_5245);
nor U5965 (N_5965,N_5283,N_5098);
and U5966 (N_5966,N_5331,N_5477);
or U5967 (N_5967,N_5468,N_5051);
nor U5968 (N_5968,N_5040,N_5280);
nand U5969 (N_5969,N_5132,N_5077);
nor U5970 (N_5970,N_5381,N_5179);
or U5971 (N_5971,N_5237,N_5311);
xor U5972 (N_5972,N_5073,N_5322);
xnor U5973 (N_5973,N_5176,N_5397);
nor U5974 (N_5974,N_5033,N_5202);
xnor U5975 (N_5975,N_5354,N_5116);
or U5976 (N_5976,N_5105,N_5045);
xnor U5977 (N_5977,N_5387,N_5353);
nor U5978 (N_5978,N_5116,N_5172);
nand U5979 (N_5979,N_5450,N_5103);
or U5980 (N_5980,N_5273,N_5103);
xor U5981 (N_5981,N_5424,N_5385);
xor U5982 (N_5982,N_5244,N_5319);
nand U5983 (N_5983,N_5418,N_5058);
nand U5984 (N_5984,N_5092,N_5076);
or U5985 (N_5985,N_5478,N_5122);
xor U5986 (N_5986,N_5063,N_5418);
nor U5987 (N_5987,N_5424,N_5050);
or U5988 (N_5988,N_5101,N_5032);
nand U5989 (N_5989,N_5093,N_5449);
nand U5990 (N_5990,N_5210,N_5425);
or U5991 (N_5991,N_5156,N_5486);
or U5992 (N_5992,N_5075,N_5223);
or U5993 (N_5993,N_5336,N_5434);
and U5994 (N_5994,N_5071,N_5488);
or U5995 (N_5995,N_5324,N_5035);
nor U5996 (N_5996,N_5438,N_5325);
nand U5997 (N_5997,N_5011,N_5369);
nor U5998 (N_5998,N_5457,N_5170);
or U5999 (N_5999,N_5088,N_5430);
nand U6000 (N_6000,N_5767,N_5893);
nand U6001 (N_6001,N_5680,N_5827);
nor U6002 (N_6002,N_5528,N_5540);
or U6003 (N_6003,N_5689,N_5803);
nand U6004 (N_6004,N_5994,N_5949);
and U6005 (N_6005,N_5718,N_5860);
nand U6006 (N_6006,N_5802,N_5877);
nand U6007 (N_6007,N_5886,N_5721);
nand U6008 (N_6008,N_5610,N_5837);
and U6009 (N_6009,N_5789,N_5587);
nor U6010 (N_6010,N_5525,N_5653);
nor U6011 (N_6011,N_5894,N_5513);
nor U6012 (N_6012,N_5874,N_5751);
nand U6013 (N_6013,N_5698,N_5656);
nor U6014 (N_6014,N_5942,N_5547);
and U6015 (N_6015,N_5965,N_5558);
or U6016 (N_6016,N_5768,N_5934);
and U6017 (N_6017,N_5628,N_5992);
nand U6018 (N_6018,N_5616,N_5676);
nor U6019 (N_6019,N_5695,N_5622);
or U6020 (N_6020,N_5574,N_5601);
nor U6021 (N_6021,N_5604,N_5771);
or U6022 (N_6022,N_5760,N_5909);
nor U6023 (N_6023,N_5902,N_5754);
xnor U6024 (N_6024,N_5922,N_5642);
nand U6025 (N_6025,N_5801,N_5815);
and U6026 (N_6026,N_5570,N_5581);
nor U6027 (N_6027,N_5609,N_5649);
and U6028 (N_6028,N_5555,N_5692);
xnor U6029 (N_6029,N_5707,N_5770);
or U6030 (N_6030,N_5843,N_5944);
xnor U6031 (N_6031,N_5667,N_5685);
xnor U6032 (N_6032,N_5614,N_5853);
xnor U6033 (N_6033,N_5966,N_5811);
xnor U6034 (N_6034,N_5535,N_5539);
and U6035 (N_6035,N_5793,N_5746);
xor U6036 (N_6036,N_5903,N_5573);
nand U6037 (N_6037,N_5638,N_5559);
nor U6038 (N_6038,N_5560,N_5504);
xnor U6039 (N_6039,N_5820,N_5505);
or U6040 (N_6040,N_5727,N_5995);
and U6041 (N_6041,N_5659,N_5910);
or U6042 (N_6042,N_5654,N_5800);
xnor U6043 (N_6043,N_5948,N_5591);
nor U6044 (N_6044,N_5683,N_5854);
nor U6045 (N_6045,N_5631,N_5589);
and U6046 (N_6046,N_5921,N_5621);
nand U6047 (N_6047,N_5788,N_5963);
nand U6048 (N_6048,N_5749,N_5930);
and U6049 (N_6049,N_5700,N_5779);
nand U6050 (N_6050,N_5943,N_5594);
nand U6051 (N_6051,N_5812,N_5915);
and U6052 (N_6052,N_5896,N_5805);
nor U6053 (N_6053,N_5858,N_5791);
xor U6054 (N_6054,N_5567,N_5534);
and U6055 (N_6055,N_5947,N_5565);
or U6056 (N_6056,N_5536,N_5872);
nor U6057 (N_6057,N_5512,N_5806);
and U6058 (N_6058,N_5748,N_5813);
or U6059 (N_6059,N_5730,N_5905);
xnor U6060 (N_6060,N_5875,N_5797);
nor U6061 (N_6061,N_5762,N_5712);
nand U6062 (N_6062,N_5979,N_5816);
nand U6063 (N_6063,N_5550,N_5696);
or U6064 (N_6064,N_5546,N_5742);
nor U6065 (N_6065,N_5529,N_5744);
nand U6066 (N_6066,N_5969,N_5509);
nor U6067 (N_6067,N_5941,N_5929);
or U6068 (N_6068,N_5832,N_5599);
nor U6069 (N_6069,N_5703,N_5554);
and U6070 (N_6070,N_5898,N_5849);
xor U6071 (N_6071,N_5835,N_5527);
or U6072 (N_6072,N_5850,N_5545);
nor U6073 (N_6073,N_5734,N_5597);
xor U6074 (N_6074,N_5920,N_5794);
nor U6075 (N_6075,N_5764,N_5900);
or U6076 (N_6076,N_5838,N_5919);
nand U6077 (N_6077,N_5911,N_5724);
nand U6078 (N_6078,N_5510,N_5772);
and U6079 (N_6079,N_5731,N_5785);
nor U6080 (N_6080,N_5758,N_5636);
nand U6081 (N_6081,N_5757,N_5799);
and U6082 (N_6082,N_5926,N_5964);
xnor U6083 (N_6083,N_5501,N_5627);
nand U6084 (N_6084,N_5989,N_5766);
nor U6085 (N_6085,N_5928,N_5603);
nand U6086 (N_6086,N_5795,N_5723);
nand U6087 (N_6087,N_5836,N_5739);
or U6088 (N_6088,N_5821,N_5613);
xnor U6089 (N_6089,N_5857,N_5950);
nand U6090 (N_6090,N_5952,N_5852);
and U6091 (N_6091,N_5842,N_5881);
and U6092 (N_6092,N_5940,N_5787);
or U6093 (N_6093,N_5830,N_5693);
xnor U6094 (N_6094,N_5755,N_5522);
xor U6095 (N_6095,N_5887,N_5959);
xnor U6096 (N_6096,N_5737,N_5732);
nand U6097 (N_6097,N_5652,N_5885);
xnor U6098 (N_6098,N_5583,N_5983);
or U6099 (N_6099,N_5974,N_5745);
nor U6100 (N_6100,N_5569,N_5880);
xnor U6101 (N_6101,N_5508,N_5516);
and U6102 (N_6102,N_5579,N_5765);
or U6103 (N_6103,N_5935,N_5968);
nand U6104 (N_6104,N_5862,N_5517);
nor U6105 (N_6105,N_5895,N_5997);
nor U6106 (N_6106,N_5503,N_5980);
xor U6107 (N_6107,N_5936,N_5780);
nand U6108 (N_6108,N_5932,N_5595);
and U6109 (N_6109,N_5551,N_5564);
nor U6110 (N_6110,N_5592,N_5677);
xnor U6111 (N_6111,N_5848,N_5580);
nand U6112 (N_6112,N_5702,N_5533);
nand U6113 (N_6113,N_5688,N_5657);
nor U6114 (N_6114,N_5866,N_5856);
and U6115 (N_6115,N_5519,N_5892);
nand U6116 (N_6116,N_5699,N_5648);
and U6117 (N_6117,N_5725,N_5623);
or U6118 (N_6118,N_5669,N_5863);
xnor U6119 (N_6119,N_5781,N_5984);
xor U6120 (N_6120,N_5641,N_5982);
or U6121 (N_6121,N_5690,N_5810);
nand U6122 (N_6122,N_5606,N_5809);
or U6123 (N_6123,N_5607,N_5675);
or U6124 (N_6124,N_5951,N_5988);
nor U6125 (N_6125,N_5655,N_5883);
xor U6126 (N_6126,N_5532,N_5553);
and U6127 (N_6127,N_5956,N_5868);
nor U6128 (N_6128,N_5520,N_5914);
or U6129 (N_6129,N_5987,N_5684);
or U6130 (N_6130,N_5720,N_5640);
nand U6131 (N_6131,N_5687,N_5998);
or U6132 (N_6132,N_5518,N_5598);
nor U6133 (N_6133,N_5918,N_5960);
nor U6134 (N_6134,N_5869,N_5679);
and U6135 (N_6135,N_5973,N_5955);
nand U6136 (N_6136,N_5888,N_5643);
nand U6137 (N_6137,N_5753,N_5818);
or U6138 (N_6138,N_5879,N_5639);
nand U6139 (N_6139,N_5741,N_5511);
and U6140 (N_6140,N_5701,N_5904);
nand U6141 (N_6141,N_5912,N_5939);
or U6142 (N_6142,N_5870,N_5549);
nor U6143 (N_6143,N_5637,N_5826);
nand U6144 (N_6144,N_5530,N_5543);
nand U6145 (N_6145,N_5844,N_5867);
nor U6146 (N_6146,N_5552,N_5713);
or U6147 (N_6147,N_5538,N_5600);
or U6148 (N_6148,N_5889,N_5661);
xnor U6149 (N_6149,N_5673,N_5873);
nor U6150 (N_6150,N_5861,N_5711);
nor U6151 (N_6151,N_5761,N_5938);
nand U6152 (N_6152,N_5747,N_5927);
xor U6153 (N_6153,N_5976,N_5996);
or U6154 (N_6154,N_5561,N_5807);
and U6155 (N_6155,N_5937,N_5515);
xor U6156 (N_6156,N_5882,N_5953);
nor U6157 (N_6157,N_5773,N_5786);
xnor U6158 (N_6158,N_5541,N_5735);
nor U6159 (N_6159,N_5878,N_5967);
xnor U6160 (N_6160,N_5908,N_5819);
and U6161 (N_6161,N_5664,N_5563);
nor U6162 (N_6162,N_5716,N_5526);
or U6163 (N_6163,N_5733,N_5993);
xnor U6164 (N_6164,N_5681,N_5593);
or U6165 (N_6165,N_5740,N_5970);
nand U6166 (N_6166,N_5962,N_5670);
xor U6167 (N_6167,N_5682,N_5602);
or U6168 (N_6168,N_5626,N_5986);
or U6169 (N_6169,N_5708,N_5778);
or U6170 (N_6170,N_5822,N_5808);
xnor U6171 (N_6171,N_5899,N_5829);
and U6172 (N_6172,N_5999,N_5769);
and U6173 (N_6173,N_5705,N_5542);
and U6174 (N_6174,N_5906,N_5584);
nor U6175 (N_6175,N_5840,N_5972);
xnor U6176 (N_6176,N_5715,N_5500);
and U6177 (N_6177,N_5971,N_5804);
and U6178 (N_6178,N_5650,N_5834);
xor U6179 (N_6179,N_5884,N_5586);
nand U6180 (N_6180,N_5923,N_5665);
xor U6181 (N_6181,N_5714,N_5946);
and U6182 (N_6182,N_5756,N_5671);
xor U6183 (N_6183,N_5577,N_5644);
nand U6184 (N_6184,N_5890,N_5502);
or U6185 (N_6185,N_5719,N_5846);
xnor U6186 (N_6186,N_5945,N_5825);
xor U6187 (N_6187,N_5859,N_5871);
or U6188 (N_6188,N_5991,N_5845);
nand U6189 (N_6189,N_5612,N_5537);
and U6190 (N_6190,N_5833,N_5824);
or U6191 (N_6191,N_5514,N_5691);
nand U6192 (N_6192,N_5978,N_5814);
and U6193 (N_6193,N_5647,N_5726);
and U6194 (N_6194,N_5568,N_5663);
and U6195 (N_6195,N_5524,N_5575);
xnor U6196 (N_6196,N_5585,N_5752);
xnor U6197 (N_6197,N_5672,N_5706);
nor U6198 (N_6198,N_5710,N_5775);
or U6199 (N_6199,N_5562,N_5704);
or U6200 (N_6200,N_5617,N_5728);
nand U6201 (N_6201,N_5578,N_5783);
xor U6202 (N_6202,N_5544,N_5777);
xnor U6203 (N_6203,N_5658,N_5957);
nor U6204 (N_6204,N_5763,N_5847);
and U6205 (N_6205,N_5615,N_5774);
and U6206 (N_6206,N_5851,N_5865);
xnor U6207 (N_6207,N_5556,N_5784);
nor U6208 (N_6208,N_5990,N_5931);
xnor U6209 (N_6209,N_5660,N_5817);
nor U6210 (N_6210,N_5736,N_5611);
or U6211 (N_6211,N_5782,N_5662);
and U6212 (N_6212,N_5828,N_5645);
xnor U6213 (N_6213,N_5855,N_5605);
or U6214 (N_6214,N_5633,N_5717);
nand U6215 (N_6215,N_5531,N_5632);
and U6216 (N_6216,N_5975,N_5548);
nor U6217 (N_6217,N_5722,N_5743);
and U6218 (N_6218,N_5954,N_5521);
and U6219 (N_6219,N_5933,N_5619);
and U6220 (N_6220,N_5738,N_5566);
and U6221 (N_6221,N_5917,N_5796);
nand U6222 (N_6222,N_5588,N_5913);
nand U6223 (N_6223,N_5582,N_5666);
and U6224 (N_6224,N_5646,N_5925);
nor U6225 (N_6225,N_5864,N_5590);
nor U6226 (N_6226,N_5823,N_5958);
and U6227 (N_6227,N_5694,N_5596);
and U6228 (N_6228,N_5651,N_5608);
and U6229 (N_6229,N_5897,N_5759);
nand U6230 (N_6230,N_5841,N_5798);
or U6231 (N_6231,N_5924,N_5624);
nand U6232 (N_6232,N_5790,N_5674);
and U6233 (N_6233,N_5776,N_5839);
and U6234 (N_6234,N_5686,N_5916);
and U6235 (N_6235,N_5876,N_5620);
and U6236 (N_6236,N_5961,N_5635);
nand U6237 (N_6237,N_5697,N_5985);
nor U6238 (N_6238,N_5792,N_5634);
xnor U6239 (N_6239,N_5977,N_5618);
nand U6240 (N_6240,N_5709,N_5576);
and U6241 (N_6241,N_5629,N_5891);
and U6242 (N_6242,N_5750,N_5630);
nor U6243 (N_6243,N_5572,N_5907);
nand U6244 (N_6244,N_5901,N_5729);
xor U6245 (N_6245,N_5557,N_5981);
xnor U6246 (N_6246,N_5668,N_5678);
nand U6247 (N_6247,N_5571,N_5523);
nand U6248 (N_6248,N_5831,N_5507);
nor U6249 (N_6249,N_5506,N_5625);
or U6250 (N_6250,N_5904,N_5823);
nor U6251 (N_6251,N_5889,N_5963);
nor U6252 (N_6252,N_5534,N_5895);
nand U6253 (N_6253,N_5528,N_5753);
xor U6254 (N_6254,N_5756,N_5635);
xnor U6255 (N_6255,N_5809,N_5916);
nand U6256 (N_6256,N_5516,N_5973);
nand U6257 (N_6257,N_5670,N_5650);
nor U6258 (N_6258,N_5790,N_5562);
xor U6259 (N_6259,N_5628,N_5639);
and U6260 (N_6260,N_5505,N_5972);
and U6261 (N_6261,N_5729,N_5760);
and U6262 (N_6262,N_5805,N_5661);
nand U6263 (N_6263,N_5642,N_5610);
or U6264 (N_6264,N_5701,N_5950);
and U6265 (N_6265,N_5511,N_5717);
and U6266 (N_6266,N_5876,N_5545);
xnor U6267 (N_6267,N_5545,N_5793);
or U6268 (N_6268,N_5728,N_5654);
and U6269 (N_6269,N_5745,N_5805);
nor U6270 (N_6270,N_5660,N_5996);
xor U6271 (N_6271,N_5673,N_5753);
xnor U6272 (N_6272,N_5561,N_5655);
nand U6273 (N_6273,N_5579,N_5607);
or U6274 (N_6274,N_5504,N_5941);
nand U6275 (N_6275,N_5879,N_5671);
nand U6276 (N_6276,N_5580,N_5875);
nand U6277 (N_6277,N_5982,N_5992);
xnor U6278 (N_6278,N_5707,N_5983);
nor U6279 (N_6279,N_5688,N_5953);
xnor U6280 (N_6280,N_5715,N_5723);
nor U6281 (N_6281,N_5535,N_5905);
xnor U6282 (N_6282,N_5898,N_5762);
or U6283 (N_6283,N_5848,N_5934);
and U6284 (N_6284,N_5865,N_5882);
xnor U6285 (N_6285,N_5996,N_5655);
nor U6286 (N_6286,N_5810,N_5507);
and U6287 (N_6287,N_5756,N_5893);
or U6288 (N_6288,N_5682,N_5996);
nor U6289 (N_6289,N_5953,N_5846);
nand U6290 (N_6290,N_5723,N_5755);
nand U6291 (N_6291,N_5623,N_5818);
and U6292 (N_6292,N_5976,N_5966);
or U6293 (N_6293,N_5949,N_5951);
nor U6294 (N_6294,N_5721,N_5972);
or U6295 (N_6295,N_5563,N_5672);
nor U6296 (N_6296,N_5610,N_5822);
xor U6297 (N_6297,N_5785,N_5950);
nor U6298 (N_6298,N_5786,N_5886);
xor U6299 (N_6299,N_5587,N_5726);
nand U6300 (N_6300,N_5689,N_5665);
nor U6301 (N_6301,N_5843,N_5846);
nor U6302 (N_6302,N_5734,N_5731);
or U6303 (N_6303,N_5916,N_5579);
nor U6304 (N_6304,N_5972,N_5658);
nand U6305 (N_6305,N_5798,N_5852);
nand U6306 (N_6306,N_5771,N_5778);
nor U6307 (N_6307,N_5837,N_5984);
and U6308 (N_6308,N_5641,N_5904);
nand U6309 (N_6309,N_5854,N_5829);
xnor U6310 (N_6310,N_5990,N_5557);
nand U6311 (N_6311,N_5857,N_5769);
nor U6312 (N_6312,N_5576,N_5942);
nor U6313 (N_6313,N_5907,N_5594);
xor U6314 (N_6314,N_5981,N_5700);
xor U6315 (N_6315,N_5786,N_5718);
xnor U6316 (N_6316,N_5768,N_5558);
and U6317 (N_6317,N_5922,N_5937);
xor U6318 (N_6318,N_5888,N_5605);
or U6319 (N_6319,N_5979,N_5746);
nand U6320 (N_6320,N_5727,N_5641);
or U6321 (N_6321,N_5944,N_5542);
xor U6322 (N_6322,N_5643,N_5646);
nand U6323 (N_6323,N_5999,N_5762);
xnor U6324 (N_6324,N_5908,N_5739);
or U6325 (N_6325,N_5967,N_5555);
nand U6326 (N_6326,N_5763,N_5764);
nand U6327 (N_6327,N_5760,N_5569);
nor U6328 (N_6328,N_5979,N_5594);
nor U6329 (N_6329,N_5512,N_5980);
and U6330 (N_6330,N_5727,N_5559);
xor U6331 (N_6331,N_5692,N_5973);
or U6332 (N_6332,N_5642,N_5673);
nand U6333 (N_6333,N_5788,N_5810);
nor U6334 (N_6334,N_5792,N_5811);
nor U6335 (N_6335,N_5580,N_5568);
or U6336 (N_6336,N_5649,N_5711);
xnor U6337 (N_6337,N_5976,N_5954);
and U6338 (N_6338,N_5609,N_5681);
or U6339 (N_6339,N_5782,N_5626);
or U6340 (N_6340,N_5562,N_5911);
xor U6341 (N_6341,N_5546,N_5542);
and U6342 (N_6342,N_5839,N_5816);
nor U6343 (N_6343,N_5966,N_5958);
nor U6344 (N_6344,N_5994,N_5540);
nand U6345 (N_6345,N_5536,N_5770);
xor U6346 (N_6346,N_5665,N_5610);
nor U6347 (N_6347,N_5723,N_5564);
nand U6348 (N_6348,N_5882,N_5916);
xnor U6349 (N_6349,N_5965,N_5707);
or U6350 (N_6350,N_5982,N_5888);
and U6351 (N_6351,N_5705,N_5632);
and U6352 (N_6352,N_5678,N_5729);
and U6353 (N_6353,N_5674,N_5913);
nand U6354 (N_6354,N_5991,N_5526);
or U6355 (N_6355,N_5561,N_5993);
and U6356 (N_6356,N_5773,N_5972);
and U6357 (N_6357,N_5950,N_5613);
nand U6358 (N_6358,N_5614,N_5663);
or U6359 (N_6359,N_5508,N_5835);
xnor U6360 (N_6360,N_5624,N_5799);
nor U6361 (N_6361,N_5661,N_5834);
and U6362 (N_6362,N_5875,N_5741);
or U6363 (N_6363,N_5830,N_5861);
nand U6364 (N_6364,N_5601,N_5733);
and U6365 (N_6365,N_5757,N_5696);
or U6366 (N_6366,N_5582,N_5888);
nand U6367 (N_6367,N_5517,N_5974);
and U6368 (N_6368,N_5560,N_5932);
nor U6369 (N_6369,N_5598,N_5781);
or U6370 (N_6370,N_5623,N_5988);
nand U6371 (N_6371,N_5552,N_5859);
nor U6372 (N_6372,N_5551,N_5672);
and U6373 (N_6373,N_5738,N_5864);
xor U6374 (N_6374,N_5635,N_5676);
xnor U6375 (N_6375,N_5980,N_5500);
nor U6376 (N_6376,N_5545,N_5739);
and U6377 (N_6377,N_5682,N_5591);
nand U6378 (N_6378,N_5704,N_5816);
and U6379 (N_6379,N_5615,N_5757);
nor U6380 (N_6380,N_5984,N_5557);
nand U6381 (N_6381,N_5600,N_5894);
nand U6382 (N_6382,N_5862,N_5557);
and U6383 (N_6383,N_5584,N_5561);
or U6384 (N_6384,N_5656,N_5563);
xnor U6385 (N_6385,N_5667,N_5720);
or U6386 (N_6386,N_5739,N_5822);
nor U6387 (N_6387,N_5925,N_5801);
nand U6388 (N_6388,N_5933,N_5612);
nor U6389 (N_6389,N_5701,N_5672);
or U6390 (N_6390,N_5573,N_5703);
nand U6391 (N_6391,N_5915,N_5521);
nand U6392 (N_6392,N_5753,N_5703);
xnor U6393 (N_6393,N_5564,N_5752);
nor U6394 (N_6394,N_5780,N_5808);
nor U6395 (N_6395,N_5999,N_5626);
or U6396 (N_6396,N_5648,N_5757);
xor U6397 (N_6397,N_5658,N_5771);
or U6398 (N_6398,N_5864,N_5913);
nand U6399 (N_6399,N_5956,N_5890);
or U6400 (N_6400,N_5587,N_5937);
or U6401 (N_6401,N_5950,N_5723);
xor U6402 (N_6402,N_5831,N_5715);
and U6403 (N_6403,N_5623,N_5999);
or U6404 (N_6404,N_5725,N_5708);
or U6405 (N_6405,N_5734,N_5867);
nor U6406 (N_6406,N_5629,N_5538);
nand U6407 (N_6407,N_5618,N_5507);
nand U6408 (N_6408,N_5659,N_5897);
or U6409 (N_6409,N_5597,N_5884);
nor U6410 (N_6410,N_5877,N_5770);
nor U6411 (N_6411,N_5586,N_5807);
and U6412 (N_6412,N_5876,N_5972);
nand U6413 (N_6413,N_5593,N_5684);
and U6414 (N_6414,N_5927,N_5857);
nand U6415 (N_6415,N_5550,N_5598);
or U6416 (N_6416,N_5709,N_5521);
xnor U6417 (N_6417,N_5911,N_5656);
or U6418 (N_6418,N_5675,N_5960);
nor U6419 (N_6419,N_5659,N_5900);
nand U6420 (N_6420,N_5872,N_5740);
or U6421 (N_6421,N_5923,N_5816);
or U6422 (N_6422,N_5811,N_5894);
or U6423 (N_6423,N_5922,N_5608);
or U6424 (N_6424,N_5946,N_5764);
nand U6425 (N_6425,N_5992,N_5655);
nand U6426 (N_6426,N_5664,N_5680);
or U6427 (N_6427,N_5658,N_5644);
and U6428 (N_6428,N_5965,N_5826);
or U6429 (N_6429,N_5870,N_5696);
or U6430 (N_6430,N_5746,N_5973);
xnor U6431 (N_6431,N_5867,N_5859);
or U6432 (N_6432,N_5606,N_5548);
nand U6433 (N_6433,N_5961,N_5773);
and U6434 (N_6434,N_5731,N_5910);
xor U6435 (N_6435,N_5882,N_5987);
and U6436 (N_6436,N_5885,N_5958);
nor U6437 (N_6437,N_5922,N_5738);
nor U6438 (N_6438,N_5792,N_5779);
xnor U6439 (N_6439,N_5818,N_5981);
or U6440 (N_6440,N_5500,N_5673);
or U6441 (N_6441,N_5904,N_5882);
and U6442 (N_6442,N_5695,N_5786);
nand U6443 (N_6443,N_5820,N_5641);
nor U6444 (N_6444,N_5738,N_5640);
and U6445 (N_6445,N_5567,N_5729);
and U6446 (N_6446,N_5840,N_5606);
nand U6447 (N_6447,N_5638,N_5685);
nand U6448 (N_6448,N_5971,N_5597);
xor U6449 (N_6449,N_5989,N_5571);
nor U6450 (N_6450,N_5808,N_5994);
or U6451 (N_6451,N_5984,N_5614);
nor U6452 (N_6452,N_5876,N_5634);
xnor U6453 (N_6453,N_5866,N_5557);
nor U6454 (N_6454,N_5727,N_5749);
xnor U6455 (N_6455,N_5798,N_5598);
and U6456 (N_6456,N_5539,N_5725);
nand U6457 (N_6457,N_5625,N_5593);
or U6458 (N_6458,N_5662,N_5515);
or U6459 (N_6459,N_5816,N_5615);
xnor U6460 (N_6460,N_5789,N_5666);
nor U6461 (N_6461,N_5946,N_5624);
nand U6462 (N_6462,N_5934,N_5942);
xnor U6463 (N_6463,N_5500,N_5564);
or U6464 (N_6464,N_5792,N_5586);
nand U6465 (N_6465,N_5800,N_5510);
xnor U6466 (N_6466,N_5732,N_5577);
nand U6467 (N_6467,N_5553,N_5976);
nor U6468 (N_6468,N_5567,N_5924);
and U6469 (N_6469,N_5551,N_5646);
xor U6470 (N_6470,N_5790,N_5571);
or U6471 (N_6471,N_5950,N_5915);
xor U6472 (N_6472,N_5877,N_5815);
and U6473 (N_6473,N_5774,N_5543);
or U6474 (N_6474,N_5701,N_5740);
nand U6475 (N_6475,N_5880,N_5596);
nor U6476 (N_6476,N_5794,N_5869);
and U6477 (N_6477,N_5621,N_5728);
nand U6478 (N_6478,N_5689,N_5768);
nand U6479 (N_6479,N_5992,N_5563);
nand U6480 (N_6480,N_5872,N_5634);
nand U6481 (N_6481,N_5706,N_5897);
or U6482 (N_6482,N_5897,N_5788);
nand U6483 (N_6483,N_5974,N_5695);
xor U6484 (N_6484,N_5927,N_5529);
and U6485 (N_6485,N_5607,N_5656);
and U6486 (N_6486,N_5649,N_5562);
nand U6487 (N_6487,N_5956,N_5839);
and U6488 (N_6488,N_5803,N_5542);
nor U6489 (N_6489,N_5653,N_5644);
xnor U6490 (N_6490,N_5632,N_5861);
nand U6491 (N_6491,N_5974,N_5734);
xnor U6492 (N_6492,N_5617,N_5931);
or U6493 (N_6493,N_5563,N_5849);
nor U6494 (N_6494,N_5774,N_5560);
nor U6495 (N_6495,N_5792,N_5960);
nand U6496 (N_6496,N_5967,N_5974);
nand U6497 (N_6497,N_5683,N_5710);
or U6498 (N_6498,N_5798,N_5959);
nor U6499 (N_6499,N_5946,N_5532);
nand U6500 (N_6500,N_6223,N_6001);
nand U6501 (N_6501,N_6067,N_6043);
nor U6502 (N_6502,N_6019,N_6193);
and U6503 (N_6503,N_6023,N_6374);
xnor U6504 (N_6504,N_6215,N_6300);
xnor U6505 (N_6505,N_6158,N_6259);
nor U6506 (N_6506,N_6005,N_6137);
or U6507 (N_6507,N_6159,N_6454);
nand U6508 (N_6508,N_6060,N_6085);
nand U6509 (N_6509,N_6165,N_6465);
nand U6510 (N_6510,N_6065,N_6253);
or U6511 (N_6511,N_6007,N_6452);
nand U6512 (N_6512,N_6451,N_6036);
and U6513 (N_6513,N_6309,N_6236);
and U6514 (N_6514,N_6275,N_6395);
and U6515 (N_6515,N_6360,N_6419);
and U6516 (N_6516,N_6366,N_6473);
and U6517 (N_6517,N_6108,N_6328);
and U6518 (N_6518,N_6289,N_6111);
nand U6519 (N_6519,N_6181,N_6341);
xor U6520 (N_6520,N_6481,N_6029);
and U6521 (N_6521,N_6082,N_6324);
nand U6522 (N_6522,N_6078,N_6327);
and U6523 (N_6523,N_6089,N_6378);
nand U6524 (N_6524,N_6225,N_6350);
xor U6525 (N_6525,N_6017,N_6206);
nor U6526 (N_6526,N_6457,N_6381);
and U6527 (N_6527,N_6006,N_6117);
and U6528 (N_6528,N_6427,N_6315);
xor U6529 (N_6529,N_6485,N_6428);
nand U6530 (N_6530,N_6266,N_6425);
and U6531 (N_6531,N_6140,N_6476);
nand U6532 (N_6532,N_6415,N_6359);
and U6533 (N_6533,N_6035,N_6471);
and U6534 (N_6534,N_6299,N_6077);
and U6535 (N_6535,N_6002,N_6346);
nor U6536 (N_6536,N_6279,N_6308);
or U6537 (N_6537,N_6151,N_6333);
and U6538 (N_6538,N_6087,N_6373);
nor U6539 (N_6539,N_6458,N_6405);
nand U6540 (N_6540,N_6478,N_6335);
and U6541 (N_6541,N_6355,N_6139);
and U6542 (N_6542,N_6201,N_6310);
or U6543 (N_6543,N_6363,N_6008);
nor U6544 (N_6544,N_6039,N_6463);
and U6545 (N_6545,N_6109,N_6073);
xor U6546 (N_6546,N_6276,N_6311);
or U6547 (N_6547,N_6442,N_6093);
or U6548 (N_6548,N_6025,N_6216);
or U6549 (N_6549,N_6095,N_6453);
nand U6550 (N_6550,N_6084,N_6022);
and U6551 (N_6551,N_6116,N_6396);
and U6552 (N_6552,N_6479,N_6297);
xor U6553 (N_6553,N_6034,N_6021);
or U6554 (N_6554,N_6145,N_6123);
nand U6555 (N_6555,N_6287,N_6343);
or U6556 (N_6556,N_6278,N_6371);
nand U6557 (N_6557,N_6440,N_6293);
nand U6558 (N_6558,N_6254,N_6393);
nor U6559 (N_6559,N_6238,N_6198);
or U6560 (N_6560,N_6285,N_6450);
nand U6561 (N_6561,N_6199,N_6301);
nor U6562 (N_6562,N_6464,N_6026);
nand U6563 (N_6563,N_6132,N_6334);
or U6564 (N_6564,N_6076,N_6369);
and U6565 (N_6565,N_6409,N_6296);
and U6566 (N_6566,N_6177,N_6098);
nor U6567 (N_6567,N_6414,N_6200);
and U6568 (N_6568,N_6348,N_6243);
nand U6569 (N_6569,N_6188,N_6171);
nor U6570 (N_6570,N_6056,N_6179);
or U6571 (N_6571,N_6062,N_6375);
xor U6572 (N_6572,N_6252,N_6050);
xor U6573 (N_6573,N_6417,N_6340);
or U6574 (N_6574,N_6048,N_6064);
and U6575 (N_6575,N_6434,N_6175);
and U6576 (N_6576,N_6474,N_6424);
and U6577 (N_6577,N_6319,N_6103);
and U6578 (N_6578,N_6086,N_6125);
and U6579 (N_6579,N_6420,N_6379);
and U6580 (N_6580,N_6102,N_6245);
nor U6581 (N_6581,N_6160,N_6352);
nand U6582 (N_6582,N_6012,N_6263);
xnor U6583 (N_6583,N_6129,N_6045);
nand U6584 (N_6584,N_6155,N_6498);
nand U6585 (N_6585,N_6030,N_6456);
xnor U6586 (N_6586,N_6314,N_6257);
nor U6587 (N_6587,N_6380,N_6219);
or U6588 (N_6588,N_6217,N_6265);
nand U6589 (N_6589,N_6090,N_6063);
or U6590 (N_6590,N_6182,N_6234);
and U6591 (N_6591,N_6467,N_6264);
nor U6592 (N_6592,N_6221,N_6397);
nand U6593 (N_6593,N_6488,N_6432);
nor U6594 (N_6594,N_6059,N_6307);
xnor U6595 (N_6595,N_6429,N_6241);
and U6596 (N_6596,N_6148,N_6183);
xor U6597 (N_6597,N_6180,N_6291);
or U6598 (N_6598,N_6016,N_6038);
xnor U6599 (N_6599,N_6455,N_6196);
nand U6600 (N_6600,N_6051,N_6430);
and U6601 (N_6601,N_6439,N_6357);
xnor U6602 (N_6602,N_6230,N_6482);
nand U6603 (N_6603,N_6469,N_6233);
and U6604 (N_6604,N_6143,N_6411);
xor U6605 (N_6605,N_6449,N_6492);
nand U6606 (N_6606,N_6274,N_6162);
xor U6607 (N_6607,N_6068,N_6150);
nor U6608 (N_6608,N_6049,N_6489);
xor U6609 (N_6609,N_6448,N_6403);
xnor U6610 (N_6610,N_6486,N_6094);
xor U6611 (N_6611,N_6009,N_6401);
nor U6612 (N_6612,N_6041,N_6295);
nor U6613 (N_6613,N_6462,N_6244);
and U6614 (N_6614,N_6246,N_6337);
and U6615 (N_6615,N_6214,N_6120);
or U6616 (N_6616,N_6024,N_6205);
nor U6617 (N_6617,N_6433,N_6326);
nand U6618 (N_6618,N_6010,N_6100);
xor U6619 (N_6619,N_6031,N_6446);
and U6620 (N_6620,N_6203,N_6262);
and U6621 (N_6621,N_6218,N_6437);
nand U6622 (N_6622,N_6280,N_6362);
nor U6623 (N_6623,N_6410,N_6057);
or U6624 (N_6624,N_6174,N_6475);
nor U6625 (N_6625,N_6080,N_6130);
nor U6626 (N_6626,N_6018,N_6407);
nand U6627 (N_6627,N_6075,N_6466);
or U6628 (N_6628,N_6000,N_6261);
nand U6629 (N_6629,N_6081,N_6367);
nand U6630 (N_6630,N_6389,N_6282);
nor U6631 (N_6631,N_6222,N_6040);
nor U6632 (N_6632,N_6232,N_6114);
nand U6633 (N_6633,N_6110,N_6304);
nand U6634 (N_6634,N_6496,N_6406);
and U6635 (N_6635,N_6322,N_6185);
and U6636 (N_6636,N_6088,N_6320);
and U6637 (N_6637,N_6186,N_6163);
xnor U6638 (N_6638,N_6204,N_6107);
nand U6639 (N_6639,N_6248,N_6497);
nor U6640 (N_6640,N_6164,N_6286);
or U6641 (N_6641,N_6388,N_6484);
nand U6642 (N_6642,N_6493,N_6166);
or U6643 (N_6643,N_6436,N_6161);
nor U6644 (N_6644,N_6459,N_6172);
or U6645 (N_6645,N_6237,N_6312);
nand U6646 (N_6646,N_6046,N_6447);
nor U6647 (N_6647,N_6313,N_6037);
or U6648 (N_6648,N_6384,N_6468);
nand U6649 (N_6649,N_6404,N_6231);
xnor U6650 (N_6650,N_6272,N_6480);
nand U6651 (N_6651,N_6047,N_6271);
xor U6652 (N_6652,N_6494,N_6247);
nand U6653 (N_6653,N_6118,N_6028);
nand U6654 (N_6654,N_6273,N_6268);
nor U6655 (N_6655,N_6240,N_6044);
nor U6656 (N_6656,N_6113,N_6444);
xnor U6657 (N_6657,N_6441,N_6070);
xnor U6658 (N_6658,N_6336,N_6292);
and U6659 (N_6659,N_6147,N_6499);
nand U6660 (N_6660,N_6156,N_6170);
or U6661 (N_6661,N_6235,N_6144);
or U6662 (N_6662,N_6472,N_6119);
and U6663 (N_6663,N_6364,N_6052);
or U6664 (N_6664,N_6211,N_6220);
or U6665 (N_6665,N_6255,N_6491);
xnor U6666 (N_6666,N_6288,N_6423);
or U6667 (N_6667,N_6399,N_6391);
or U6668 (N_6668,N_6256,N_6318);
xnor U6669 (N_6669,N_6408,N_6135);
nand U6670 (N_6670,N_6074,N_6011);
nor U6671 (N_6671,N_6412,N_6226);
nor U6672 (N_6672,N_6136,N_6126);
nor U6673 (N_6673,N_6416,N_6099);
and U6674 (N_6674,N_6014,N_6385);
or U6675 (N_6675,N_6338,N_6382);
xnor U6676 (N_6676,N_6013,N_6305);
or U6677 (N_6677,N_6197,N_6202);
or U6678 (N_6678,N_6210,N_6277);
nor U6679 (N_6679,N_6176,N_6072);
or U6680 (N_6680,N_6258,N_6242);
and U6681 (N_6681,N_6394,N_6386);
or U6682 (N_6682,N_6392,N_6435);
and U6683 (N_6683,N_6191,N_6091);
and U6684 (N_6684,N_6490,N_6368);
or U6685 (N_6685,N_6267,N_6418);
or U6686 (N_6686,N_6227,N_6122);
nand U6687 (N_6687,N_6269,N_6330);
nand U6688 (N_6688,N_6487,N_6224);
nor U6689 (N_6689,N_6194,N_6195);
and U6690 (N_6690,N_6347,N_6290);
nor U6691 (N_6691,N_6317,N_6303);
nor U6692 (N_6692,N_6323,N_6331);
and U6693 (N_6693,N_6079,N_6146);
nand U6694 (N_6694,N_6376,N_6101);
xor U6695 (N_6695,N_6104,N_6192);
and U6696 (N_6696,N_6281,N_6115);
xnor U6697 (N_6697,N_6069,N_6157);
or U6698 (N_6698,N_6128,N_6460);
and U6699 (N_6699,N_6345,N_6053);
xor U6700 (N_6700,N_6402,N_6298);
xor U6701 (N_6701,N_6431,N_6426);
or U6702 (N_6702,N_6054,N_6342);
or U6703 (N_6703,N_6332,N_6004);
or U6704 (N_6704,N_6131,N_6339);
xor U6705 (N_6705,N_6027,N_6377);
nand U6706 (N_6706,N_6189,N_6461);
and U6707 (N_6707,N_6066,N_6260);
xnor U6708 (N_6708,N_6096,N_6400);
xnor U6709 (N_6709,N_6354,N_6284);
xnor U6710 (N_6710,N_6344,N_6212);
or U6711 (N_6711,N_6083,N_6370);
and U6712 (N_6712,N_6365,N_6351);
nand U6713 (N_6713,N_6142,N_6356);
and U6714 (N_6714,N_6124,N_6187);
or U6715 (N_6715,N_6495,N_6390);
or U6716 (N_6716,N_6239,N_6121);
xor U6717 (N_6717,N_6294,N_6190);
xnor U6718 (N_6718,N_6209,N_6106);
and U6719 (N_6719,N_6207,N_6283);
nand U6720 (N_6720,N_6015,N_6020);
nor U6721 (N_6721,N_6306,N_6168);
and U6722 (N_6722,N_6152,N_6316);
nor U6723 (N_6723,N_6438,N_6184);
xor U6724 (N_6724,N_6361,N_6228);
or U6725 (N_6725,N_6092,N_6445);
or U6726 (N_6726,N_6033,N_6229);
nand U6727 (N_6727,N_6134,N_6270);
nand U6728 (N_6728,N_6138,N_6213);
and U6729 (N_6729,N_6398,N_6071);
nor U6730 (N_6730,N_6169,N_6154);
and U6731 (N_6731,N_6112,N_6042);
or U6732 (N_6732,N_6329,N_6422);
nand U6733 (N_6733,N_6208,N_6105);
and U6734 (N_6734,N_6032,N_6383);
or U6735 (N_6735,N_6353,N_6127);
and U6736 (N_6736,N_6058,N_6178);
or U6737 (N_6737,N_6302,N_6421);
or U6738 (N_6738,N_6251,N_6443);
nor U6739 (N_6739,N_6153,N_6173);
nand U6740 (N_6740,N_6387,N_6061);
and U6741 (N_6741,N_6483,N_6133);
and U6742 (N_6742,N_6167,N_6413);
nand U6743 (N_6743,N_6470,N_6372);
xor U6744 (N_6744,N_6325,N_6097);
nand U6745 (N_6745,N_6003,N_6055);
nand U6746 (N_6746,N_6141,N_6249);
nand U6747 (N_6747,N_6149,N_6250);
or U6748 (N_6748,N_6477,N_6349);
or U6749 (N_6749,N_6358,N_6321);
xnor U6750 (N_6750,N_6083,N_6071);
nor U6751 (N_6751,N_6186,N_6489);
or U6752 (N_6752,N_6000,N_6127);
and U6753 (N_6753,N_6007,N_6281);
nand U6754 (N_6754,N_6110,N_6129);
nor U6755 (N_6755,N_6427,N_6060);
or U6756 (N_6756,N_6002,N_6315);
or U6757 (N_6757,N_6448,N_6178);
nor U6758 (N_6758,N_6163,N_6251);
nor U6759 (N_6759,N_6420,N_6192);
or U6760 (N_6760,N_6289,N_6355);
nand U6761 (N_6761,N_6175,N_6346);
xnor U6762 (N_6762,N_6075,N_6045);
and U6763 (N_6763,N_6110,N_6256);
and U6764 (N_6764,N_6221,N_6071);
and U6765 (N_6765,N_6163,N_6348);
xnor U6766 (N_6766,N_6188,N_6010);
and U6767 (N_6767,N_6438,N_6318);
and U6768 (N_6768,N_6249,N_6454);
nor U6769 (N_6769,N_6211,N_6379);
or U6770 (N_6770,N_6238,N_6214);
nor U6771 (N_6771,N_6014,N_6134);
nor U6772 (N_6772,N_6141,N_6046);
nor U6773 (N_6773,N_6141,N_6422);
or U6774 (N_6774,N_6210,N_6370);
and U6775 (N_6775,N_6452,N_6149);
nand U6776 (N_6776,N_6456,N_6336);
nand U6777 (N_6777,N_6196,N_6229);
or U6778 (N_6778,N_6033,N_6460);
xor U6779 (N_6779,N_6430,N_6250);
nand U6780 (N_6780,N_6325,N_6457);
nand U6781 (N_6781,N_6379,N_6297);
nor U6782 (N_6782,N_6455,N_6274);
nor U6783 (N_6783,N_6141,N_6070);
nand U6784 (N_6784,N_6356,N_6179);
nand U6785 (N_6785,N_6131,N_6184);
nor U6786 (N_6786,N_6389,N_6145);
nand U6787 (N_6787,N_6206,N_6093);
xor U6788 (N_6788,N_6023,N_6220);
nor U6789 (N_6789,N_6272,N_6101);
xnor U6790 (N_6790,N_6367,N_6460);
nand U6791 (N_6791,N_6096,N_6298);
nand U6792 (N_6792,N_6215,N_6419);
nor U6793 (N_6793,N_6231,N_6478);
nand U6794 (N_6794,N_6204,N_6379);
nor U6795 (N_6795,N_6476,N_6200);
nand U6796 (N_6796,N_6406,N_6129);
nand U6797 (N_6797,N_6483,N_6344);
nor U6798 (N_6798,N_6250,N_6133);
and U6799 (N_6799,N_6430,N_6167);
or U6800 (N_6800,N_6323,N_6384);
and U6801 (N_6801,N_6476,N_6395);
nand U6802 (N_6802,N_6447,N_6028);
nand U6803 (N_6803,N_6234,N_6162);
nand U6804 (N_6804,N_6338,N_6372);
or U6805 (N_6805,N_6060,N_6200);
or U6806 (N_6806,N_6272,N_6214);
or U6807 (N_6807,N_6399,N_6356);
or U6808 (N_6808,N_6230,N_6196);
nand U6809 (N_6809,N_6257,N_6406);
nand U6810 (N_6810,N_6146,N_6439);
or U6811 (N_6811,N_6053,N_6042);
nor U6812 (N_6812,N_6370,N_6473);
nand U6813 (N_6813,N_6320,N_6344);
nand U6814 (N_6814,N_6304,N_6302);
nand U6815 (N_6815,N_6397,N_6083);
or U6816 (N_6816,N_6127,N_6329);
nor U6817 (N_6817,N_6482,N_6367);
nor U6818 (N_6818,N_6394,N_6408);
or U6819 (N_6819,N_6345,N_6132);
nand U6820 (N_6820,N_6189,N_6425);
nand U6821 (N_6821,N_6116,N_6181);
xnor U6822 (N_6822,N_6328,N_6373);
or U6823 (N_6823,N_6454,N_6482);
nor U6824 (N_6824,N_6199,N_6469);
nor U6825 (N_6825,N_6149,N_6119);
or U6826 (N_6826,N_6375,N_6453);
nor U6827 (N_6827,N_6025,N_6367);
xor U6828 (N_6828,N_6302,N_6379);
xnor U6829 (N_6829,N_6216,N_6427);
and U6830 (N_6830,N_6083,N_6482);
xor U6831 (N_6831,N_6167,N_6185);
and U6832 (N_6832,N_6232,N_6220);
xor U6833 (N_6833,N_6036,N_6034);
and U6834 (N_6834,N_6347,N_6140);
nand U6835 (N_6835,N_6021,N_6474);
nand U6836 (N_6836,N_6382,N_6333);
and U6837 (N_6837,N_6003,N_6157);
xnor U6838 (N_6838,N_6205,N_6268);
xor U6839 (N_6839,N_6167,N_6173);
xor U6840 (N_6840,N_6290,N_6274);
nand U6841 (N_6841,N_6410,N_6004);
xnor U6842 (N_6842,N_6473,N_6263);
nand U6843 (N_6843,N_6383,N_6401);
nand U6844 (N_6844,N_6089,N_6449);
or U6845 (N_6845,N_6225,N_6307);
and U6846 (N_6846,N_6086,N_6037);
nor U6847 (N_6847,N_6189,N_6109);
nand U6848 (N_6848,N_6210,N_6264);
nand U6849 (N_6849,N_6468,N_6322);
and U6850 (N_6850,N_6054,N_6337);
or U6851 (N_6851,N_6341,N_6083);
nor U6852 (N_6852,N_6244,N_6149);
xor U6853 (N_6853,N_6406,N_6389);
or U6854 (N_6854,N_6233,N_6428);
and U6855 (N_6855,N_6331,N_6443);
and U6856 (N_6856,N_6379,N_6270);
and U6857 (N_6857,N_6233,N_6119);
and U6858 (N_6858,N_6244,N_6264);
nor U6859 (N_6859,N_6013,N_6402);
nand U6860 (N_6860,N_6453,N_6261);
nand U6861 (N_6861,N_6492,N_6487);
or U6862 (N_6862,N_6077,N_6437);
or U6863 (N_6863,N_6463,N_6499);
nand U6864 (N_6864,N_6137,N_6312);
xnor U6865 (N_6865,N_6232,N_6359);
and U6866 (N_6866,N_6352,N_6002);
nor U6867 (N_6867,N_6181,N_6003);
nor U6868 (N_6868,N_6345,N_6272);
or U6869 (N_6869,N_6118,N_6492);
or U6870 (N_6870,N_6179,N_6297);
xnor U6871 (N_6871,N_6277,N_6092);
xnor U6872 (N_6872,N_6224,N_6246);
xor U6873 (N_6873,N_6133,N_6205);
nand U6874 (N_6874,N_6029,N_6431);
xnor U6875 (N_6875,N_6154,N_6489);
or U6876 (N_6876,N_6070,N_6363);
nand U6877 (N_6877,N_6050,N_6281);
and U6878 (N_6878,N_6470,N_6085);
or U6879 (N_6879,N_6255,N_6450);
and U6880 (N_6880,N_6273,N_6301);
nand U6881 (N_6881,N_6103,N_6195);
and U6882 (N_6882,N_6065,N_6100);
nor U6883 (N_6883,N_6344,N_6284);
nand U6884 (N_6884,N_6199,N_6461);
and U6885 (N_6885,N_6057,N_6391);
and U6886 (N_6886,N_6114,N_6394);
nand U6887 (N_6887,N_6151,N_6210);
xnor U6888 (N_6888,N_6077,N_6022);
or U6889 (N_6889,N_6189,N_6284);
and U6890 (N_6890,N_6080,N_6280);
nor U6891 (N_6891,N_6496,N_6355);
and U6892 (N_6892,N_6496,N_6415);
or U6893 (N_6893,N_6491,N_6250);
and U6894 (N_6894,N_6198,N_6125);
nand U6895 (N_6895,N_6213,N_6461);
and U6896 (N_6896,N_6460,N_6489);
xor U6897 (N_6897,N_6306,N_6474);
nand U6898 (N_6898,N_6248,N_6112);
xor U6899 (N_6899,N_6111,N_6215);
nor U6900 (N_6900,N_6417,N_6358);
or U6901 (N_6901,N_6302,N_6189);
and U6902 (N_6902,N_6187,N_6110);
nor U6903 (N_6903,N_6459,N_6242);
xor U6904 (N_6904,N_6377,N_6492);
xnor U6905 (N_6905,N_6223,N_6244);
xor U6906 (N_6906,N_6040,N_6457);
xor U6907 (N_6907,N_6498,N_6227);
xor U6908 (N_6908,N_6043,N_6251);
and U6909 (N_6909,N_6182,N_6465);
or U6910 (N_6910,N_6496,N_6267);
xor U6911 (N_6911,N_6237,N_6005);
xnor U6912 (N_6912,N_6249,N_6066);
and U6913 (N_6913,N_6168,N_6149);
or U6914 (N_6914,N_6380,N_6386);
and U6915 (N_6915,N_6273,N_6316);
nor U6916 (N_6916,N_6472,N_6399);
xor U6917 (N_6917,N_6382,N_6346);
and U6918 (N_6918,N_6070,N_6324);
nor U6919 (N_6919,N_6223,N_6402);
nand U6920 (N_6920,N_6400,N_6143);
nand U6921 (N_6921,N_6331,N_6234);
nand U6922 (N_6922,N_6357,N_6442);
and U6923 (N_6923,N_6110,N_6128);
nor U6924 (N_6924,N_6046,N_6301);
nand U6925 (N_6925,N_6107,N_6223);
and U6926 (N_6926,N_6453,N_6268);
nand U6927 (N_6927,N_6272,N_6252);
xor U6928 (N_6928,N_6059,N_6414);
or U6929 (N_6929,N_6109,N_6126);
nor U6930 (N_6930,N_6369,N_6420);
or U6931 (N_6931,N_6091,N_6352);
and U6932 (N_6932,N_6382,N_6491);
nor U6933 (N_6933,N_6114,N_6081);
nor U6934 (N_6934,N_6301,N_6070);
xor U6935 (N_6935,N_6290,N_6394);
xnor U6936 (N_6936,N_6239,N_6305);
xnor U6937 (N_6937,N_6129,N_6049);
and U6938 (N_6938,N_6145,N_6264);
nor U6939 (N_6939,N_6416,N_6037);
and U6940 (N_6940,N_6259,N_6453);
and U6941 (N_6941,N_6159,N_6458);
nand U6942 (N_6942,N_6192,N_6081);
xnor U6943 (N_6943,N_6406,N_6310);
xor U6944 (N_6944,N_6416,N_6403);
xnor U6945 (N_6945,N_6108,N_6354);
and U6946 (N_6946,N_6269,N_6146);
xnor U6947 (N_6947,N_6134,N_6078);
and U6948 (N_6948,N_6107,N_6093);
nand U6949 (N_6949,N_6259,N_6391);
nand U6950 (N_6950,N_6423,N_6221);
or U6951 (N_6951,N_6468,N_6389);
nand U6952 (N_6952,N_6241,N_6125);
xnor U6953 (N_6953,N_6324,N_6388);
nand U6954 (N_6954,N_6386,N_6370);
or U6955 (N_6955,N_6290,N_6325);
nor U6956 (N_6956,N_6438,N_6202);
nand U6957 (N_6957,N_6477,N_6206);
nor U6958 (N_6958,N_6314,N_6062);
nand U6959 (N_6959,N_6424,N_6159);
or U6960 (N_6960,N_6493,N_6205);
nand U6961 (N_6961,N_6310,N_6279);
xor U6962 (N_6962,N_6049,N_6467);
nand U6963 (N_6963,N_6171,N_6361);
or U6964 (N_6964,N_6237,N_6426);
nand U6965 (N_6965,N_6337,N_6207);
nand U6966 (N_6966,N_6210,N_6434);
nand U6967 (N_6967,N_6490,N_6474);
nand U6968 (N_6968,N_6433,N_6135);
nand U6969 (N_6969,N_6404,N_6495);
nor U6970 (N_6970,N_6244,N_6040);
xor U6971 (N_6971,N_6102,N_6220);
or U6972 (N_6972,N_6227,N_6454);
xnor U6973 (N_6973,N_6046,N_6357);
and U6974 (N_6974,N_6045,N_6385);
xor U6975 (N_6975,N_6334,N_6434);
nor U6976 (N_6976,N_6340,N_6356);
xor U6977 (N_6977,N_6036,N_6395);
nor U6978 (N_6978,N_6442,N_6068);
nor U6979 (N_6979,N_6308,N_6322);
nand U6980 (N_6980,N_6154,N_6313);
xor U6981 (N_6981,N_6251,N_6489);
or U6982 (N_6982,N_6455,N_6023);
nand U6983 (N_6983,N_6437,N_6337);
xnor U6984 (N_6984,N_6168,N_6185);
nand U6985 (N_6985,N_6007,N_6224);
nand U6986 (N_6986,N_6185,N_6323);
xor U6987 (N_6987,N_6272,N_6484);
xnor U6988 (N_6988,N_6097,N_6035);
or U6989 (N_6989,N_6061,N_6242);
nor U6990 (N_6990,N_6108,N_6090);
and U6991 (N_6991,N_6491,N_6283);
and U6992 (N_6992,N_6436,N_6044);
nand U6993 (N_6993,N_6001,N_6068);
or U6994 (N_6994,N_6092,N_6062);
nand U6995 (N_6995,N_6128,N_6218);
or U6996 (N_6996,N_6099,N_6329);
or U6997 (N_6997,N_6254,N_6450);
or U6998 (N_6998,N_6001,N_6451);
and U6999 (N_6999,N_6222,N_6275);
nand U7000 (N_7000,N_6979,N_6732);
nand U7001 (N_7001,N_6548,N_6850);
nand U7002 (N_7002,N_6805,N_6720);
or U7003 (N_7003,N_6676,N_6827);
and U7004 (N_7004,N_6917,N_6881);
or U7005 (N_7005,N_6928,N_6655);
nand U7006 (N_7006,N_6714,N_6648);
and U7007 (N_7007,N_6656,N_6746);
nor U7008 (N_7008,N_6927,N_6970);
nand U7009 (N_7009,N_6954,N_6911);
nand U7010 (N_7010,N_6856,N_6697);
xnor U7011 (N_7011,N_6510,N_6978);
and U7012 (N_7012,N_6859,N_6992);
or U7013 (N_7013,N_6711,N_6902);
nand U7014 (N_7014,N_6782,N_6769);
xnor U7015 (N_7015,N_6799,N_6562);
nand U7016 (N_7016,N_6605,N_6767);
or U7017 (N_7017,N_6557,N_6907);
or U7018 (N_7018,N_6612,N_6895);
nand U7019 (N_7019,N_6649,N_6729);
nor U7020 (N_7020,N_6749,N_6646);
or U7021 (N_7021,N_6584,N_6855);
or U7022 (N_7022,N_6873,N_6880);
nand U7023 (N_7023,N_6781,N_6694);
nor U7024 (N_7024,N_6900,N_6857);
nand U7025 (N_7025,N_6804,N_6922);
nand U7026 (N_7026,N_6773,N_6607);
xnor U7027 (N_7027,N_6645,N_6643);
nand U7028 (N_7028,N_6709,N_6872);
nand U7029 (N_7029,N_6555,N_6915);
nor U7030 (N_7030,N_6823,N_6606);
nor U7031 (N_7031,N_6620,N_6705);
nor U7032 (N_7032,N_6968,N_6544);
or U7033 (N_7033,N_6817,N_6719);
xnor U7034 (N_7034,N_6835,N_6683);
nor U7035 (N_7035,N_6977,N_6766);
nand U7036 (N_7036,N_6721,N_6563);
nand U7037 (N_7037,N_6520,N_6863);
and U7038 (N_7038,N_6508,N_6809);
and U7039 (N_7039,N_6901,N_6972);
xor U7040 (N_7040,N_6813,N_6945);
or U7041 (N_7041,N_6851,N_6765);
nand U7042 (N_7042,N_6808,N_6586);
nand U7043 (N_7043,N_6757,N_6576);
and U7044 (N_7044,N_6879,N_6830);
and U7045 (N_7045,N_6688,N_6819);
or U7046 (N_7046,N_6654,N_6681);
and U7047 (N_7047,N_6780,N_6628);
xnor U7048 (N_7048,N_6989,N_6678);
xnor U7049 (N_7049,N_6957,N_6952);
and U7050 (N_7050,N_6843,N_6999);
nand U7051 (N_7051,N_6869,N_6938);
or U7052 (N_7052,N_6906,N_6867);
or U7053 (N_7053,N_6501,N_6741);
or U7054 (N_7054,N_6725,N_6824);
and U7055 (N_7055,N_6959,N_6583);
xor U7056 (N_7056,N_6702,N_6998);
and U7057 (N_7057,N_6600,N_6523);
and U7058 (N_7058,N_6975,N_6937);
nand U7059 (N_7059,N_6886,N_6580);
or U7060 (N_7060,N_6524,N_6762);
nand U7061 (N_7061,N_6662,N_6770);
and U7062 (N_7062,N_6955,N_6953);
nor U7063 (N_7063,N_6944,N_6517);
xnor U7064 (N_7064,N_6986,N_6512);
nand U7065 (N_7065,N_6667,N_6644);
or U7066 (N_7066,N_6818,N_6784);
or U7067 (N_7067,N_6558,N_6540);
or U7068 (N_7068,N_6533,N_6883);
nor U7069 (N_7069,N_6587,N_6786);
and U7070 (N_7070,N_6526,N_6931);
xnor U7071 (N_7071,N_6845,N_6939);
or U7072 (N_7072,N_6897,N_6949);
and U7073 (N_7073,N_6751,N_6595);
nor U7074 (N_7074,N_6511,N_6619);
nand U7075 (N_7075,N_6575,N_6987);
and U7076 (N_7076,N_6599,N_6613);
or U7077 (N_7077,N_6803,N_6704);
or U7078 (N_7078,N_6635,N_6829);
and U7079 (N_7079,N_6858,N_6918);
and U7080 (N_7080,N_6534,N_6618);
xor U7081 (N_7081,N_6842,N_6878);
xnor U7082 (N_7082,N_6754,N_6973);
nor U7083 (N_7083,N_6984,N_6592);
nand U7084 (N_7084,N_6737,N_6726);
and U7085 (N_7085,N_6779,N_6525);
xnor U7086 (N_7086,N_6701,N_6797);
or U7087 (N_7087,N_6788,N_6854);
and U7088 (N_7088,N_6904,N_6868);
and U7089 (N_7089,N_6752,N_6825);
xor U7090 (N_7090,N_6846,N_6509);
or U7091 (N_7091,N_6703,N_6602);
nor U7092 (N_7092,N_6964,N_6798);
xor U7093 (N_7093,N_6995,N_6545);
nor U7094 (N_7094,N_6996,N_6764);
nor U7095 (N_7095,N_6727,N_6930);
xnor U7096 (N_7096,N_6932,N_6514);
or U7097 (N_7097,N_6549,N_6621);
and U7098 (N_7098,N_6682,N_6617);
xnor U7099 (N_7099,N_6743,N_6696);
and U7100 (N_7100,N_6724,N_6777);
nor U7101 (N_7101,N_6862,N_6861);
nor U7102 (N_7102,N_6903,N_6899);
nor U7103 (N_7103,N_6666,N_6958);
nor U7104 (N_7104,N_6734,N_6527);
xnor U7105 (N_7105,N_6971,N_6876);
or U7106 (N_7106,N_6691,N_6756);
nor U7107 (N_7107,N_6626,N_6513);
xor U7108 (N_7108,N_6594,N_6636);
nand U7109 (N_7109,N_6565,N_6951);
or U7110 (N_7110,N_6875,N_6969);
or U7111 (N_7111,N_6559,N_6547);
nor U7112 (N_7112,N_6651,N_6844);
xnor U7113 (N_7113,N_6864,N_6577);
and U7114 (N_7114,N_6976,N_6556);
nand U7115 (N_7115,N_6624,N_6736);
nand U7116 (N_7116,N_6776,N_6553);
nand U7117 (N_7117,N_6874,N_6647);
or U7118 (N_7118,N_6745,N_6740);
and U7119 (N_7119,N_6625,N_6710);
and U7120 (N_7120,N_6708,N_6733);
xor U7121 (N_7121,N_6763,N_6689);
or U7122 (N_7122,N_6622,N_6965);
nor U7123 (N_7123,N_6564,N_6921);
and U7124 (N_7124,N_6674,N_6759);
or U7125 (N_7125,N_6695,N_6811);
nor U7126 (N_7126,N_6632,N_6603);
and U7127 (N_7127,N_6578,N_6812);
xnor U7128 (N_7128,N_6891,N_6518);
or U7129 (N_7129,N_6985,N_6761);
xnor U7130 (N_7130,N_6896,N_6833);
xnor U7131 (N_7131,N_6742,N_6551);
or U7132 (N_7132,N_6980,N_6807);
or U7133 (N_7133,N_6659,N_6841);
xnor U7134 (N_7134,N_6794,N_6774);
or U7135 (N_7135,N_6848,N_6601);
or U7136 (N_7136,N_6739,N_6672);
nor U7137 (N_7137,N_6700,N_6828);
nand U7138 (N_7138,N_6680,N_6693);
and U7139 (N_7139,N_6669,N_6806);
nor U7140 (N_7140,N_6816,N_6870);
and U7141 (N_7141,N_6546,N_6639);
or U7142 (N_7142,N_6832,N_6660);
nand U7143 (N_7143,N_6983,N_6608);
nand U7144 (N_7144,N_6566,N_6963);
nor U7145 (N_7145,N_6554,N_6597);
xor U7146 (N_7146,N_6994,N_6919);
and U7147 (N_7147,N_6790,N_6589);
or U7148 (N_7148,N_6570,N_6820);
nand U7149 (N_7149,N_6860,N_6650);
xor U7150 (N_7150,N_6528,N_6991);
and U7151 (N_7151,N_6853,N_6627);
nand U7152 (N_7152,N_6529,N_6609);
xnor U7153 (N_7153,N_6793,N_6671);
nand U7154 (N_7154,N_6502,N_6849);
nand U7155 (N_7155,N_6661,N_6738);
nand U7156 (N_7156,N_6747,N_6950);
or U7157 (N_7157,N_6568,N_6506);
and U7158 (N_7158,N_6685,N_6715);
nand U7159 (N_7159,N_6722,N_6658);
nand U7160 (N_7160,N_6614,N_6538);
and U7161 (N_7161,N_6503,N_6634);
or U7162 (N_7162,N_6912,N_6591);
and U7163 (N_7163,N_6935,N_6974);
or U7164 (N_7164,N_6686,N_6598);
or U7165 (N_7165,N_6967,N_6698);
xnor U7166 (N_7166,N_6800,N_6673);
and U7167 (N_7167,N_6934,N_6877);
and U7168 (N_7168,N_6560,N_6760);
or U7169 (N_7169,N_6638,N_6585);
xor U7170 (N_7170,N_6888,N_6615);
nand U7171 (N_7171,N_6839,N_6926);
and U7172 (N_7172,N_6679,N_6961);
or U7173 (N_7173,N_6909,N_6611);
xnor U7174 (N_7174,N_6982,N_6692);
and U7175 (N_7175,N_6730,N_6519);
xor U7176 (N_7176,N_6796,N_6535);
and U7177 (N_7177,N_6834,N_6567);
xor U7178 (N_7178,N_6943,N_6997);
or U7179 (N_7179,N_6706,N_6596);
nor U7180 (N_7180,N_6956,N_6947);
or U7181 (N_7181,N_6775,N_6581);
nand U7182 (N_7182,N_6604,N_6731);
xor U7183 (N_7183,N_6795,N_6684);
xnor U7184 (N_7184,N_6532,N_6801);
and U7185 (N_7185,N_6552,N_6791);
nor U7186 (N_7186,N_6936,N_6582);
or U7187 (N_7187,N_6981,N_6753);
xnor U7188 (N_7188,N_6542,N_6574);
or U7189 (N_7189,N_6838,N_6713);
or U7190 (N_7190,N_6718,N_6537);
nor U7191 (N_7191,N_6665,N_6758);
nor U7192 (N_7192,N_6561,N_6633);
xnor U7193 (N_7193,N_6707,N_6593);
and U7194 (N_7194,N_6924,N_6892);
nor U7195 (N_7195,N_6573,N_6810);
xor U7196 (N_7196,N_6815,N_6925);
xnor U7197 (N_7197,N_6623,N_6664);
or U7198 (N_7198,N_6933,N_6687);
xor U7199 (N_7199,N_6590,N_6908);
nor U7200 (N_7200,N_6630,N_6550);
nor U7201 (N_7201,N_6913,N_6588);
nand U7202 (N_7202,N_6675,N_6629);
nor U7203 (N_7203,N_6822,N_6530);
nand U7204 (N_7204,N_6768,N_6852);
nor U7205 (N_7205,N_6993,N_6500);
xor U7206 (N_7206,N_6882,N_6914);
or U7207 (N_7207,N_6699,N_6962);
xor U7208 (N_7208,N_6516,N_6960);
nor U7209 (N_7209,N_6946,N_6889);
nor U7210 (N_7210,N_6748,N_6966);
and U7211 (N_7211,N_6531,N_6717);
and U7212 (N_7212,N_6657,N_6865);
xnor U7213 (N_7213,N_6836,N_6920);
nand U7214 (N_7214,N_6887,N_6785);
or U7215 (N_7215,N_6543,N_6579);
nor U7216 (N_7216,N_6610,N_6988);
and U7217 (N_7217,N_6894,N_6572);
nand U7218 (N_7218,N_6755,N_6885);
and U7219 (N_7219,N_6942,N_6821);
nor U7220 (N_7220,N_6505,N_6783);
xnor U7221 (N_7221,N_6890,N_6668);
and U7222 (N_7222,N_6652,N_6663);
or U7223 (N_7223,N_6670,N_6884);
and U7224 (N_7224,N_6814,N_6792);
nor U7225 (N_7225,N_6789,N_6637);
nor U7226 (N_7226,N_6735,N_6941);
nor U7227 (N_7227,N_6772,N_6916);
or U7228 (N_7228,N_6515,N_6522);
and U7229 (N_7229,N_6840,N_6948);
xor U7230 (N_7230,N_6905,N_6893);
nor U7231 (N_7231,N_6541,N_6571);
and U7232 (N_7232,N_6871,N_6866);
nor U7233 (N_7233,N_6750,N_6504);
and U7234 (N_7234,N_6712,N_6539);
nor U7235 (N_7235,N_6847,N_6787);
nor U7236 (N_7236,N_6744,N_6723);
nand U7237 (N_7237,N_6569,N_6929);
nand U7238 (N_7238,N_6990,N_6940);
nand U7239 (N_7239,N_6728,N_6831);
or U7240 (N_7240,N_6716,N_6641);
and U7241 (N_7241,N_6837,N_6690);
and U7242 (N_7242,N_6910,N_6507);
nand U7243 (N_7243,N_6631,N_6771);
nor U7244 (N_7244,N_6536,N_6640);
and U7245 (N_7245,N_6826,N_6616);
nand U7246 (N_7246,N_6521,N_6802);
and U7247 (N_7247,N_6642,N_6923);
nor U7248 (N_7248,N_6898,N_6677);
xor U7249 (N_7249,N_6653,N_6778);
and U7250 (N_7250,N_6991,N_6965);
nor U7251 (N_7251,N_6504,N_6561);
or U7252 (N_7252,N_6765,N_6897);
nor U7253 (N_7253,N_6639,N_6891);
nand U7254 (N_7254,N_6598,N_6984);
xor U7255 (N_7255,N_6903,N_6516);
nor U7256 (N_7256,N_6939,N_6549);
and U7257 (N_7257,N_6646,N_6904);
nand U7258 (N_7258,N_6526,N_6837);
and U7259 (N_7259,N_6862,N_6850);
and U7260 (N_7260,N_6537,N_6972);
xor U7261 (N_7261,N_6619,N_6647);
xnor U7262 (N_7262,N_6608,N_6682);
nor U7263 (N_7263,N_6908,N_6846);
nor U7264 (N_7264,N_6657,N_6882);
xnor U7265 (N_7265,N_6546,N_6796);
nand U7266 (N_7266,N_6821,N_6666);
nor U7267 (N_7267,N_6577,N_6819);
nor U7268 (N_7268,N_6581,N_6582);
nor U7269 (N_7269,N_6501,N_6937);
nand U7270 (N_7270,N_6895,N_6997);
or U7271 (N_7271,N_6643,N_6544);
or U7272 (N_7272,N_6832,N_6927);
nand U7273 (N_7273,N_6736,N_6597);
xor U7274 (N_7274,N_6815,N_6616);
or U7275 (N_7275,N_6781,N_6621);
nor U7276 (N_7276,N_6569,N_6651);
and U7277 (N_7277,N_6775,N_6854);
nor U7278 (N_7278,N_6722,N_6515);
or U7279 (N_7279,N_6663,N_6502);
nand U7280 (N_7280,N_6794,N_6573);
nand U7281 (N_7281,N_6913,N_6992);
nor U7282 (N_7282,N_6856,N_6733);
nor U7283 (N_7283,N_6594,N_6819);
or U7284 (N_7284,N_6880,N_6945);
and U7285 (N_7285,N_6603,N_6718);
nand U7286 (N_7286,N_6937,N_6952);
nand U7287 (N_7287,N_6796,N_6977);
and U7288 (N_7288,N_6890,N_6781);
and U7289 (N_7289,N_6706,N_6503);
and U7290 (N_7290,N_6586,N_6819);
and U7291 (N_7291,N_6841,N_6988);
or U7292 (N_7292,N_6986,N_6955);
nor U7293 (N_7293,N_6635,N_6905);
and U7294 (N_7294,N_6571,N_6779);
xor U7295 (N_7295,N_6791,N_6625);
xnor U7296 (N_7296,N_6789,N_6783);
nor U7297 (N_7297,N_6965,N_6736);
or U7298 (N_7298,N_6621,N_6991);
and U7299 (N_7299,N_6645,N_6852);
nor U7300 (N_7300,N_6733,N_6979);
and U7301 (N_7301,N_6561,N_6551);
xnor U7302 (N_7302,N_6584,N_6907);
and U7303 (N_7303,N_6807,N_6530);
nor U7304 (N_7304,N_6741,N_6837);
and U7305 (N_7305,N_6585,N_6782);
xnor U7306 (N_7306,N_6987,N_6759);
nor U7307 (N_7307,N_6579,N_6599);
nand U7308 (N_7308,N_6697,N_6897);
nand U7309 (N_7309,N_6722,N_6729);
and U7310 (N_7310,N_6645,N_6956);
xnor U7311 (N_7311,N_6932,N_6792);
nor U7312 (N_7312,N_6583,N_6600);
nand U7313 (N_7313,N_6910,N_6839);
or U7314 (N_7314,N_6607,N_6870);
nand U7315 (N_7315,N_6517,N_6697);
nand U7316 (N_7316,N_6580,N_6653);
xor U7317 (N_7317,N_6602,N_6847);
nand U7318 (N_7318,N_6803,N_6715);
nor U7319 (N_7319,N_6989,N_6572);
or U7320 (N_7320,N_6687,N_6751);
and U7321 (N_7321,N_6509,N_6937);
or U7322 (N_7322,N_6503,N_6964);
and U7323 (N_7323,N_6870,N_6508);
nand U7324 (N_7324,N_6556,N_6954);
xnor U7325 (N_7325,N_6706,N_6703);
and U7326 (N_7326,N_6869,N_6711);
or U7327 (N_7327,N_6699,N_6523);
nor U7328 (N_7328,N_6921,N_6605);
xnor U7329 (N_7329,N_6681,N_6694);
nand U7330 (N_7330,N_6521,N_6788);
nor U7331 (N_7331,N_6629,N_6589);
xor U7332 (N_7332,N_6699,N_6745);
nor U7333 (N_7333,N_6973,N_6638);
or U7334 (N_7334,N_6913,N_6677);
and U7335 (N_7335,N_6825,N_6638);
nand U7336 (N_7336,N_6901,N_6756);
or U7337 (N_7337,N_6904,N_6892);
or U7338 (N_7338,N_6667,N_6740);
and U7339 (N_7339,N_6862,N_6598);
nor U7340 (N_7340,N_6641,N_6664);
nand U7341 (N_7341,N_6767,N_6529);
nor U7342 (N_7342,N_6846,N_6768);
xnor U7343 (N_7343,N_6629,N_6905);
nand U7344 (N_7344,N_6803,N_6565);
nor U7345 (N_7345,N_6603,N_6726);
nor U7346 (N_7346,N_6505,N_6731);
nand U7347 (N_7347,N_6647,N_6834);
nand U7348 (N_7348,N_6976,N_6578);
or U7349 (N_7349,N_6625,N_6891);
nand U7350 (N_7350,N_6949,N_6755);
nand U7351 (N_7351,N_6700,N_6644);
or U7352 (N_7352,N_6759,N_6680);
xor U7353 (N_7353,N_6768,N_6788);
and U7354 (N_7354,N_6976,N_6642);
or U7355 (N_7355,N_6935,N_6504);
or U7356 (N_7356,N_6739,N_6891);
nor U7357 (N_7357,N_6927,N_6929);
nand U7358 (N_7358,N_6626,N_6549);
and U7359 (N_7359,N_6638,N_6806);
or U7360 (N_7360,N_6573,N_6657);
or U7361 (N_7361,N_6592,N_6773);
or U7362 (N_7362,N_6641,N_6818);
or U7363 (N_7363,N_6794,N_6931);
nand U7364 (N_7364,N_6734,N_6836);
or U7365 (N_7365,N_6988,N_6866);
xnor U7366 (N_7366,N_6843,N_6751);
or U7367 (N_7367,N_6978,N_6838);
nand U7368 (N_7368,N_6506,N_6648);
xnor U7369 (N_7369,N_6935,N_6508);
nand U7370 (N_7370,N_6584,N_6970);
nand U7371 (N_7371,N_6557,N_6588);
nor U7372 (N_7372,N_6720,N_6734);
nand U7373 (N_7373,N_6937,N_6604);
nor U7374 (N_7374,N_6848,N_6743);
nand U7375 (N_7375,N_6645,N_6928);
nor U7376 (N_7376,N_6593,N_6558);
or U7377 (N_7377,N_6569,N_6817);
nor U7378 (N_7378,N_6794,N_6831);
nor U7379 (N_7379,N_6605,N_6717);
nor U7380 (N_7380,N_6636,N_6516);
nor U7381 (N_7381,N_6874,N_6841);
xor U7382 (N_7382,N_6965,N_6958);
and U7383 (N_7383,N_6886,N_6756);
xnor U7384 (N_7384,N_6552,N_6643);
and U7385 (N_7385,N_6640,N_6603);
or U7386 (N_7386,N_6644,N_6934);
or U7387 (N_7387,N_6524,N_6988);
nand U7388 (N_7388,N_6744,N_6658);
or U7389 (N_7389,N_6627,N_6742);
nor U7390 (N_7390,N_6922,N_6552);
xnor U7391 (N_7391,N_6656,N_6916);
and U7392 (N_7392,N_6895,N_6790);
and U7393 (N_7393,N_6587,N_6701);
or U7394 (N_7394,N_6787,N_6758);
nand U7395 (N_7395,N_6787,N_6991);
or U7396 (N_7396,N_6913,N_6917);
nor U7397 (N_7397,N_6638,N_6969);
xnor U7398 (N_7398,N_6982,N_6578);
nor U7399 (N_7399,N_6527,N_6627);
nand U7400 (N_7400,N_6600,N_6929);
xor U7401 (N_7401,N_6975,N_6904);
or U7402 (N_7402,N_6639,N_6784);
or U7403 (N_7403,N_6570,N_6569);
nand U7404 (N_7404,N_6959,N_6933);
and U7405 (N_7405,N_6945,N_6971);
nand U7406 (N_7406,N_6927,N_6671);
and U7407 (N_7407,N_6813,N_6720);
and U7408 (N_7408,N_6574,N_6615);
or U7409 (N_7409,N_6912,N_6630);
or U7410 (N_7410,N_6966,N_6676);
xnor U7411 (N_7411,N_6859,N_6555);
or U7412 (N_7412,N_6975,N_6842);
nor U7413 (N_7413,N_6776,N_6880);
nor U7414 (N_7414,N_6587,N_6808);
xnor U7415 (N_7415,N_6640,N_6591);
and U7416 (N_7416,N_6562,N_6590);
or U7417 (N_7417,N_6642,N_6796);
nand U7418 (N_7418,N_6533,N_6557);
or U7419 (N_7419,N_6655,N_6962);
nand U7420 (N_7420,N_6889,N_6938);
xor U7421 (N_7421,N_6961,N_6695);
xor U7422 (N_7422,N_6592,N_6963);
or U7423 (N_7423,N_6964,N_6937);
nand U7424 (N_7424,N_6774,N_6775);
or U7425 (N_7425,N_6992,N_6609);
and U7426 (N_7426,N_6924,N_6554);
and U7427 (N_7427,N_6556,N_6922);
nor U7428 (N_7428,N_6875,N_6849);
xor U7429 (N_7429,N_6888,N_6936);
nor U7430 (N_7430,N_6913,N_6770);
nor U7431 (N_7431,N_6988,N_6808);
and U7432 (N_7432,N_6682,N_6526);
or U7433 (N_7433,N_6843,N_6774);
xor U7434 (N_7434,N_6862,N_6809);
or U7435 (N_7435,N_6856,N_6698);
or U7436 (N_7436,N_6953,N_6945);
nand U7437 (N_7437,N_6520,N_6594);
or U7438 (N_7438,N_6586,N_6674);
or U7439 (N_7439,N_6620,N_6894);
nand U7440 (N_7440,N_6888,N_6520);
nand U7441 (N_7441,N_6543,N_6818);
xnor U7442 (N_7442,N_6584,N_6788);
and U7443 (N_7443,N_6690,N_6650);
nor U7444 (N_7444,N_6877,N_6500);
and U7445 (N_7445,N_6541,N_6895);
xor U7446 (N_7446,N_6951,N_6788);
or U7447 (N_7447,N_6684,N_6859);
or U7448 (N_7448,N_6690,N_6551);
nor U7449 (N_7449,N_6881,N_6714);
nand U7450 (N_7450,N_6589,N_6707);
xor U7451 (N_7451,N_6800,N_6652);
nor U7452 (N_7452,N_6901,N_6596);
nor U7453 (N_7453,N_6715,N_6827);
and U7454 (N_7454,N_6713,N_6612);
or U7455 (N_7455,N_6958,N_6662);
or U7456 (N_7456,N_6504,N_6696);
nor U7457 (N_7457,N_6662,N_6631);
or U7458 (N_7458,N_6777,N_6518);
nor U7459 (N_7459,N_6719,N_6957);
or U7460 (N_7460,N_6897,N_6805);
xnor U7461 (N_7461,N_6813,N_6944);
nand U7462 (N_7462,N_6678,N_6760);
and U7463 (N_7463,N_6692,N_6620);
nand U7464 (N_7464,N_6855,N_6909);
nand U7465 (N_7465,N_6866,N_6857);
nand U7466 (N_7466,N_6762,N_6713);
and U7467 (N_7467,N_6940,N_6659);
or U7468 (N_7468,N_6880,N_6519);
nor U7469 (N_7469,N_6825,N_6503);
or U7470 (N_7470,N_6795,N_6759);
xnor U7471 (N_7471,N_6532,N_6565);
or U7472 (N_7472,N_6652,N_6700);
nand U7473 (N_7473,N_6717,N_6895);
and U7474 (N_7474,N_6518,N_6699);
or U7475 (N_7475,N_6680,N_6794);
nor U7476 (N_7476,N_6905,N_6784);
xor U7477 (N_7477,N_6573,N_6506);
xnor U7478 (N_7478,N_6971,N_6532);
and U7479 (N_7479,N_6515,N_6731);
or U7480 (N_7480,N_6630,N_6553);
nor U7481 (N_7481,N_6608,N_6606);
xor U7482 (N_7482,N_6806,N_6595);
xor U7483 (N_7483,N_6617,N_6551);
xnor U7484 (N_7484,N_6811,N_6600);
nor U7485 (N_7485,N_6669,N_6847);
or U7486 (N_7486,N_6653,N_6721);
nand U7487 (N_7487,N_6530,N_6681);
nand U7488 (N_7488,N_6865,N_6661);
or U7489 (N_7489,N_6997,N_6719);
nand U7490 (N_7490,N_6565,N_6783);
nor U7491 (N_7491,N_6979,N_6540);
or U7492 (N_7492,N_6960,N_6812);
nor U7493 (N_7493,N_6629,N_6844);
nor U7494 (N_7494,N_6838,N_6920);
xnor U7495 (N_7495,N_6743,N_6552);
or U7496 (N_7496,N_6804,N_6862);
and U7497 (N_7497,N_6590,N_6621);
nor U7498 (N_7498,N_6565,N_6595);
xor U7499 (N_7499,N_6656,N_6987);
nor U7500 (N_7500,N_7086,N_7367);
nand U7501 (N_7501,N_7435,N_7446);
nand U7502 (N_7502,N_7464,N_7234);
or U7503 (N_7503,N_7498,N_7315);
and U7504 (N_7504,N_7073,N_7459);
nor U7505 (N_7505,N_7474,N_7243);
and U7506 (N_7506,N_7433,N_7164);
and U7507 (N_7507,N_7001,N_7242);
nand U7508 (N_7508,N_7463,N_7019);
nor U7509 (N_7509,N_7153,N_7372);
xor U7510 (N_7510,N_7487,N_7137);
nand U7511 (N_7511,N_7323,N_7353);
and U7512 (N_7512,N_7223,N_7340);
or U7513 (N_7513,N_7026,N_7413);
or U7514 (N_7514,N_7484,N_7378);
nor U7515 (N_7515,N_7215,N_7241);
nand U7516 (N_7516,N_7300,N_7059);
nor U7517 (N_7517,N_7229,N_7496);
xnor U7518 (N_7518,N_7062,N_7076);
and U7519 (N_7519,N_7111,N_7365);
or U7520 (N_7520,N_7453,N_7410);
xor U7521 (N_7521,N_7382,N_7097);
nand U7522 (N_7522,N_7003,N_7047);
nand U7523 (N_7523,N_7472,N_7267);
nor U7524 (N_7524,N_7452,N_7371);
and U7525 (N_7525,N_7170,N_7202);
xnor U7526 (N_7526,N_7254,N_7424);
or U7527 (N_7527,N_7263,N_7205);
and U7528 (N_7528,N_7327,N_7402);
nor U7529 (N_7529,N_7189,N_7320);
or U7530 (N_7530,N_7416,N_7412);
or U7531 (N_7531,N_7099,N_7444);
nand U7532 (N_7532,N_7030,N_7049);
and U7533 (N_7533,N_7125,N_7058);
nor U7534 (N_7534,N_7477,N_7143);
nand U7535 (N_7535,N_7417,N_7129);
nor U7536 (N_7536,N_7376,N_7489);
nand U7537 (N_7537,N_7262,N_7311);
and U7538 (N_7538,N_7273,N_7008);
nand U7539 (N_7539,N_7406,N_7092);
xnor U7540 (N_7540,N_7492,N_7466);
and U7541 (N_7541,N_7405,N_7377);
or U7542 (N_7542,N_7113,N_7203);
nand U7543 (N_7543,N_7185,N_7115);
nand U7544 (N_7544,N_7269,N_7044);
or U7545 (N_7545,N_7209,N_7430);
or U7546 (N_7546,N_7290,N_7291);
nand U7547 (N_7547,N_7048,N_7027);
and U7548 (N_7548,N_7038,N_7407);
or U7549 (N_7549,N_7355,N_7260);
or U7550 (N_7550,N_7102,N_7158);
xor U7551 (N_7551,N_7188,N_7257);
nor U7552 (N_7552,N_7018,N_7043);
nor U7553 (N_7553,N_7427,N_7411);
nor U7554 (N_7554,N_7429,N_7422);
or U7555 (N_7555,N_7303,N_7014);
xor U7556 (N_7556,N_7392,N_7383);
nand U7557 (N_7557,N_7431,N_7419);
and U7558 (N_7558,N_7272,N_7293);
and U7559 (N_7559,N_7436,N_7179);
and U7560 (N_7560,N_7332,N_7298);
xnor U7561 (N_7561,N_7056,N_7445);
nor U7562 (N_7562,N_7404,N_7398);
or U7563 (N_7563,N_7385,N_7114);
xor U7564 (N_7564,N_7232,N_7283);
nor U7565 (N_7565,N_7105,N_7220);
nand U7566 (N_7566,N_7089,N_7231);
nand U7567 (N_7567,N_7370,N_7035);
nand U7568 (N_7568,N_7213,N_7434);
or U7569 (N_7569,N_7138,N_7186);
or U7570 (N_7570,N_7493,N_7235);
or U7571 (N_7571,N_7447,N_7344);
nor U7572 (N_7572,N_7473,N_7324);
and U7573 (N_7573,N_7308,N_7451);
nand U7574 (N_7574,N_7418,N_7022);
nand U7575 (N_7575,N_7469,N_7460);
nand U7576 (N_7576,N_7187,N_7321);
nand U7577 (N_7577,N_7266,N_7210);
nand U7578 (N_7578,N_7237,N_7072);
nor U7579 (N_7579,N_7197,N_7031);
nor U7580 (N_7580,N_7211,N_7393);
nor U7581 (N_7581,N_7346,N_7196);
or U7582 (N_7582,N_7178,N_7024);
xor U7583 (N_7583,N_7248,N_7455);
nor U7584 (N_7584,N_7177,N_7401);
nor U7585 (N_7585,N_7415,N_7336);
and U7586 (N_7586,N_7318,N_7119);
and U7587 (N_7587,N_7329,N_7139);
nand U7588 (N_7588,N_7294,N_7161);
nand U7589 (N_7589,N_7396,N_7354);
and U7590 (N_7590,N_7159,N_7199);
nand U7591 (N_7591,N_7258,N_7441);
and U7592 (N_7592,N_7091,N_7352);
nand U7593 (N_7593,N_7238,N_7479);
xnor U7594 (N_7594,N_7075,N_7157);
xnor U7595 (N_7595,N_7442,N_7369);
xor U7596 (N_7596,N_7192,N_7067);
and U7597 (N_7597,N_7065,N_7397);
nor U7598 (N_7598,N_7270,N_7309);
nand U7599 (N_7599,N_7148,N_7005);
or U7600 (N_7600,N_7100,N_7359);
or U7601 (N_7601,N_7122,N_7165);
and U7602 (N_7602,N_7313,N_7182);
or U7603 (N_7603,N_7448,N_7218);
nor U7604 (N_7604,N_7335,N_7098);
or U7605 (N_7605,N_7130,N_7384);
nand U7606 (N_7606,N_7387,N_7020);
and U7607 (N_7607,N_7316,N_7212);
and U7608 (N_7608,N_7015,N_7465);
or U7609 (N_7609,N_7361,N_7146);
or U7610 (N_7610,N_7214,N_7297);
nand U7611 (N_7611,N_7126,N_7201);
and U7612 (N_7612,N_7358,N_7456);
or U7613 (N_7613,N_7247,N_7368);
nand U7614 (N_7614,N_7039,N_7204);
nand U7615 (N_7615,N_7071,N_7360);
or U7616 (N_7616,N_7307,N_7194);
and U7617 (N_7617,N_7000,N_7118);
xor U7618 (N_7618,N_7305,N_7389);
nand U7619 (N_7619,N_7082,N_7362);
or U7620 (N_7620,N_7068,N_7162);
nor U7621 (N_7621,N_7364,N_7347);
nor U7622 (N_7622,N_7061,N_7490);
and U7623 (N_7623,N_7083,N_7032);
xor U7624 (N_7624,N_7328,N_7481);
xnor U7625 (N_7625,N_7227,N_7478);
nand U7626 (N_7626,N_7066,N_7259);
xor U7627 (N_7627,N_7495,N_7317);
nand U7628 (N_7628,N_7380,N_7004);
xnor U7629 (N_7629,N_7333,N_7342);
nor U7630 (N_7630,N_7304,N_7280);
or U7631 (N_7631,N_7124,N_7168);
or U7632 (N_7632,N_7440,N_7034);
or U7633 (N_7633,N_7322,N_7017);
nand U7634 (N_7634,N_7131,N_7467);
nand U7635 (N_7635,N_7287,N_7443);
nand U7636 (N_7636,N_7136,N_7261);
xor U7637 (N_7637,N_7302,N_7295);
nor U7638 (N_7638,N_7045,N_7449);
and U7639 (N_7639,N_7133,N_7399);
and U7640 (N_7640,N_7264,N_7357);
and U7641 (N_7641,N_7421,N_7348);
and U7642 (N_7642,N_7052,N_7491);
nand U7643 (N_7643,N_7007,N_7079);
nand U7644 (N_7644,N_7334,N_7011);
or U7645 (N_7645,N_7037,N_7426);
and U7646 (N_7646,N_7036,N_7166);
nor U7647 (N_7647,N_7256,N_7296);
and U7648 (N_7648,N_7468,N_7246);
xor U7649 (N_7649,N_7458,N_7470);
nor U7650 (N_7650,N_7391,N_7379);
nand U7651 (N_7651,N_7163,N_7425);
nor U7652 (N_7652,N_7351,N_7239);
nor U7653 (N_7653,N_7276,N_7169);
xor U7654 (N_7654,N_7106,N_7128);
nor U7655 (N_7655,N_7480,N_7116);
and U7656 (N_7656,N_7135,N_7233);
and U7657 (N_7657,N_7174,N_7085);
or U7658 (N_7658,N_7012,N_7471);
or U7659 (N_7659,N_7255,N_7292);
or U7660 (N_7660,N_7181,N_7054);
and U7661 (N_7661,N_7094,N_7077);
nand U7662 (N_7662,N_7141,N_7151);
nor U7663 (N_7663,N_7438,N_7288);
nand U7664 (N_7664,N_7142,N_7228);
xnor U7665 (N_7665,N_7310,N_7225);
nor U7666 (N_7666,N_7494,N_7070);
nand U7667 (N_7667,N_7193,N_7366);
or U7668 (N_7668,N_7450,N_7482);
nand U7669 (N_7669,N_7084,N_7023);
xnor U7670 (N_7670,N_7284,N_7095);
xnor U7671 (N_7671,N_7109,N_7488);
nand U7672 (N_7672,N_7394,N_7108);
nand U7673 (N_7673,N_7274,N_7282);
and U7674 (N_7674,N_7499,N_7016);
and U7675 (N_7675,N_7190,N_7338);
nor U7676 (N_7676,N_7326,N_7285);
nor U7677 (N_7677,N_7152,N_7224);
xnor U7678 (N_7678,N_7090,N_7053);
nor U7679 (N_7679,N_7078,N_7439);
nor U7680 (N_7680,N_7176,N_7183);
or U7681 (N_7681,N_7330,N_7400);
nand U7682 (N_7682,N_7010,N_7356);
and U7683 (N_7683,N_7437,N_7110);
nand U7684 (N_7684,N_7155,N_7454);
nor U7685 (N_7685,N_7497,N_7373);
nor U7686 (N_7686,N_7341,N_7041);
and U7687 (N_7687,N_7486,N_7457);
nand U7688 (N_7688,N_7221,N_7149);
nor U7689 (N_7689,N_7200,N_7132);
nor U7690 (N_7690,N_7171,N_7206);
nand U7691 (N_7691,N_7277,N_7042);
and U7692 (N_7692,N_7409,N_7060);
or U7693 (N_7693,N_7345,N_7281);
or U7694 (N_7694,N_7306,N_7278);
xor U7695 (N_7695,N_7160,N_7156);
nor U7696 (N_7696,N_7408,N_7101);
xnor U7697 (N_7697,N_7390,N_7051);
xnor U7698 (N_7698,N_7216,N_7428);
nor U7699 (N_7699,N_7134,N_7167);
xnor U7700 (N_7700,N_7096,N_7271);
nor U7701 (N_7701,N_7299,N_7103);
or U7702 (N_7702,N_7029,N_7063);
nor U7703 (N_7703,N_7325,N_7475);
xor U7704 (N_7704,N_7374,N_7144);
or U7705 (N_7705,N_7198,N_7127);
nand U7706 (N_7706,N_7363,N_7207);
and U7707 (N_7707,N_7033,N_7222);
nand U7708 (N_7708,N_7217,N_7080);
or U7709 (N_7709,N_7253,N_7343);
nor U7710 (N_7710,N_7240,N_7172);
xnor U7711 (N_7711,N_7025,N_7175);
and U7712 (N_7712,N_7485,N_7002);
or U7713 (N_7713,N_7319,N_7230);
xor U7714 (N_7714,N_7462,N_7286);
nor U7715 (N_7715,N_7057,N_7013);
nor U7716 (N_7716,N_7249,N_7147);
and U7717 (N_7717,N_7432,N_7104);
nor U7718 (N_7718,N_7381,N_7021);
and U7719 (N_7719,N_7173,N_7386);
or U7720 (N_7720,N_7423,N_7150);
or U7721 (N_7721,N_7250,N_7009);
xor U7722 (N_7722,N_7117,N_7403);
xor U7723 (N_7723,N_7195,N_7265);
nand U7724 (N_7724,N_7145,N_7244);
xnor U7725 (N_7725,N_7081,N_7121);
nand U7726 (N_7726,N_7180,N_7046);
nor U7727 (N_7727,N_7331,N_7339);
nor U7728 (N_7728,N_7040,N_7251);
nand U7729 (N_7729,N_7088,N_7483);
xor U7730 (N_7730,N_7093,N_7208);
xor U7731 (N_7731,N_7476,N_7120);
nor U7732 (N_7732,N_7461,N_7289);
nor U7733 (N_7733,N_7006,N_7395);
and U7734 (N_7734,N_7245,N_7268);
nor U7735 (N_7735,N_7349,N_7087);
xnor U7736 (N_7736,N_7069,N_7184);
or U7737 (N_7737,N_7350,N_7301);
xnor U7738 (N_7738,N_7055,N_7191);
or U7739 (N_7739,N_7074,N_7388);
nand U7740 (N_7740,N_7219,N_7028);
and U7741 (N_7741,N_7123,N_7337);
nand U7742 (N_7742,N_7154,N_7236);
nand U7743 (N_7743,N_7064,N_7312);
and U7744 (N_7744,N_7275,N_7414);
nor U7745 (N_7745,N_7140,N_7420);
or U7746 (N_7746,N_7314,N_7050);
or U7747 (N_7747,N_7252,N_7375);
nand U7748 (N_7748,N_7112,N_7279);
or U7749 (N_7749,N_7107,N_7226);
or U7750 (N_7750,N_7089,N_7422);
nand U7751 (N_7751,N_7216,N_7288);
xnor U7752 (N_7752,N_7453,N_7217);
xnor U7753 (N_7753,N_7409,N_7043);
or U7754 (N_7754,N_7144,N_7181);
and U7755 (N_7755,N_7280,N_7496);
nor U7756 (N_7756,N_7343,N_7319);
and U7757 (N_7757,N_7218,N_7098);
nand U7758 (N_7758,N_7395,N_7271);
xnor U7759 (N_7759,N_7017,N_7076);
and U7760 (N_7760,N_7340,N_7156);
or U7761 (N_7761,N_7457,N_7253);
xnor U7762 (N_7762,N_7216,N_7411);
nor U7763 (N_7763,N_7177,N_7118);
and U7764 (N_7764,N_7448,N_7128);
or U7765 (N_7765,N_7459,N_7383);
nand U7766 (N_7766,N_7225,N_7042);
and U7767 (N_7767,N_7099,N_7426);
xnor U7768 (N_7768,N_7162,N_7091);
and U7769 (N_7769,N_7401,N_7199);
and U7770 (N_7770,N_7292,N_7303);
or U7771 (N_7771,N_7380,N_7175);
nor U7772 (N_7772,N_7234,N_7098);
nor U7773 (N_7773,N_7333,N_7451);
xor U7774 (N_7774,N_7494,N_7427);
xnor U7775 (N_7775,N_7048,N_7432);
nor U7776 (N_7776,N_7234,N_7022);
and U7777 (N_7777,N_7234,N_7246);
or U7778 (N_7778,N_7192,N_7158);
and U7779 (N_7779,N_7460,N_7394);
xor U7780 (N_7780,N_7335,N_7466);
and U7781 (N_7781,N_7240,N_7104);
xnor U7782 (N_7782,N_7427,N_7227);
or U7783 (N_7783,N_7261,N_7092);
nor U7784 (N_7784,N_7201,N_7009);
xor U7785 (N_7785,N_7150,N_7383);
nor U7786 (N_7786,N_7290,N_7487);
nand U7787 (N_7787,N_7353,N_7013);
or U7788 (N_7788,N_7334,N_7070);
or U7789 (N_7789,N_7368,N_7401);
xor U7790 (N_7790,N_7352,N_7013);
and U7791 (N_7791,N_7350,N_7006);
or U7792 (N_7792,N_7356,N_7498);
and U7793 (N_7793,N_7042,N_7457);
xnor U7794 (N_7794,N_7214,N_7463);
xor U7795 (N_7795,N_7087,N_7117);
nor U7796 (N_7796,N_7247,N_7002);
xnor U7797 (N_7797,N_7445,N_7220);
xor U7798 (N_7798,N_7336,N_7376);
nand U7799 (N_7799,N_7356,N_7102);
nor U7800 (N_7800,N_7211,N_7292);
nor U7801 (N_7801,N_7413,N_7363);
xor U7802 (N_7802,N_7477,N_7369);
nand U7803 (N_7803,N_7469,N_7431);
or U7804 (N_7804,N_7423,N_7075);
nand U7805 (N_7805,N_7097,N_7230);
or U7806 (N_7806,N_7031,N_7051);
nor U7807 (N_7807,N_7116,N_7297);
nand U7808 (N_7808,N_7080,N_7362);
and U7809 (N_7809,N_7068,N_7346);
xnor U7810 (N_7810,N_7093,N_7450);
nor U7811 (N_7811,N_7275,N_7171);
nor U7812 (N_7812,N_7228,N_7347);
nor U7813 (N_7813,N_7268,N_7324);
nand U7814 (N_7814,N_7050,N_7217);
nand U7815 (N_7815,N_7300,N_7471);
nand U7816 (N_7816,N_7145,N_7196);
nor U7817 (N_7817,N_7309,N_7145);
xnor U7818 (N_7818,N_7245,N_7427);
xnor U7819 (N_7819,N_7302,N_7043);
nand U7820 (N_7820,N_7366,N_7178);
and U7821 (N_7821,N_7125,N_7176);
or U7822 (N_7822,N_7321,N_7075);
xor U7823 (N_7823,N_7095,N_7256);
and U7824 (N_7824,N_7379,N_7083);
and U7825 (N_7825,N_7230,N_7134);
and U7826 (N_7826,N_7339,N_7342);
nand U7827 (N_7827,N_7075,N_7498);
nand U7828 (N_7828,N_7078,N_7024);
nand U7829 (N_7829,N_7382,N_7178);
and U7830 (N_7830,N_7142,N_7273);
xnor U7831 (N_7831,N_7265,N_7080);
nor U7832 (N_7832,N_7464,N_7427);
nand U7833 (N_7833,N_7136,N_7245);
or U7834 (N_7834,N_7102,N_7338);
nor U7835 (N_7835,N_7014,N_7363);
nand U7836 (N_7836,N_7169,N_7244);
nand U7837 (N_7837,N_7362,N_7497);
and U7838 (N_7838,N_7097,N_7104);
or U7839 (N_7839,N_7158,N_7027);
nor U7840 (N_7840,N_7004,N_7471);
xnor U7841 (N_7841,N_7062,N_7110);
nor U7842 (N_7842,N_7398,N_7454);
nand U7843 (N_7843,N_7367,N_7319);
nand U7844 (N_7844,N_7028,N_7187);
nor U7845 (N_7845,N_7042,N_7184);
nor U7846 (N_7846,N_7073,N_7355);
and U7847 (N_7847,N_7324,N_7239);
or U7848 (N_7848,N_7068,N_7454);
or U7849 (N_7849,N_7352,N_7331);
xor U7850 (N_7850,N_7235,N_7471);
nand U7851 (N_7851,N_7227,N_7076);
or U7852 (N_7852,N_7349,N_7004);
xnor U7853 (N_7853,N_7338,N_7065);
xor U7854 (N_7854,N_7263,N_7460);
and U7855 (N_7855,N_7391,N_7344);
xor U7856 (N_7856,N_7082,N_7153);
xor U7857 (N_7857,N_7436,N_7460);
xnor U7858 (N_7858,N_7437,N_7223);
nand U7859 (N_7859,N_7104,N_7100);
nand U7860 (N_7860,N_7299,N_7187);
xor U7861 (N_7861,N_7485,N_7156);
or U7862 (N_7862,N_7313,N_7068);
and U7863 (N_7863,N_7456,N_7248);
or U7864 (N_7864,N_7110,N_7122);
nor U7865 (N_7865,N_7187,N_7015);
or U7866 (N_7866,N_7480,N_7205);
xor U7867 (N_7867,N_7430,N_7127);
or U7868 (N_7868,N_7385,N_7376);
xor U7869 (N_7869,N_7303,N_7129);
nand U7870 (N_7870,N_7288,N_7342);
nor U7871 (N_7871,N_7029,N_7261);
xnor U7872 (N_7872,N_7378,N_7444);
nor U7873 (N_7873,N_7423,N_7466);
nand U7874 (N_7874,N_7450,N_7060);
nand U7875 (N_7875,N_7495,N_7445);
nor U7876 (N_7876,N_7409,N_7465);
xnor U7877 (N_7877,N_7025,N_7015);
and U7878 (N_7878,N_7439,N_7322);
xnor U7879 (N_7879,N_7268,N_7156);
nor U7880 (N_7880,N_7283,N_7446);
xnor U7881 (N_7881,N_7007,N_7417);
nand U7882 (N_7882,N_7011,N_7418);
nor U7883 (N_7883,N_7164,N_7197);
xnor U7884 (N_7884,N_7361,N_7338);
xnor U7885 (N_7885,N_7107,N_7048);
and U7886 (N_7886,N_7139,N_7471);
nor U7887 (N_7887,N_7356,N_7405);
or U7888 (N_7888,N_7060,N_7100);
and U7889 (N_7889,N_7333,N_7032);
and U7890 (N_7890,N_7229,N_7189);
xor U7891 (N_7891,N_7440,N_7157);
xnor U7892 (N_7892,N_7035,N_7038);
and U7893 (N_7893,N_7111,N_7125);
nand U7894 (N_7894,N_7204,N_7135);
or U7895 (N_7895,N_7034,N_7290);
or U7896 (N_7896,N_7100,N_7149);
nor U7897 (N_7897,N_7055,N_7075);
nor U7898 (N_7898,N_7156,N_7280);
nor U7899 (N_7899,N_7031,N_7235);
or U7900 (N_7900,N_7166,N_7432);
nor U7901 (N_7901,N_7334,N_7091);
nand U7902 (N_7902,N_7177,N_7077);
nand U7903 (N_7903,N_7415,N_7132);
nand U7904 (N_7904,N_7266,N_7272);
and U7905 (N_7905,N_7438,N_7072);
and U7906 (N_7906,N_7057,N_7002);
nor U7907 (N_7907,N_7424,N_7238);
nor U7908 (N_7908,N_7038,N_7144);
and U7909 (N_7909,N_7073,N_7096);
nand U7910 (N_7910,N_7200,N_7334);
and U7911 (N_7911,N_7160,N_7028);
xor U7912 (N_7912,N_7127,N_7467);
and U7913 (N_7913,N_7398,N_7395);
xor U7914 (N_7914,N_7179,N_7224);
and U7915 (N_7915,N_7346,N_7168);
or U7916 (N_7916,N_7196,N_7445);
or U7917 (N_7917,N_7322,N_7498);
and U7918 (N_7918,N_7097,N_7375);
nand U7919 (N_7919,N_7297,N_7273);
or U7920 (N_7920,N_7314,N_7198);
nor U7921 (N_7921,N_7032,N_7220);
nor U7922 (N_7922,N_7088,N_7464);
and U7923 (N_7923,N_7366,N_7257);
xor U7924 (N_7924,N_7321,N_7481);
and U7925 (N_7925,N_7308,N_7341);
nor U7926 (N_7926,N_7094,N_7153);
nand U7927 (N_7927,N_7183,N_7309);
nand U7928 (N_7928,N_7495,N_7385);
nor U7929 (N_7929,N_7021,N_7017);
nand U7930 (N_7930,N_7231,N_7251);
or U7931 (N_7931,N_7286,N_7193);
or U7932 (N_7932,N_7154,N_7194);
xor U7933 (N_7933,N_7026,N_7315);
or U7934 (N_7934,N_7264,N_7299);
nand U7935 (N_7935,N_7373,N_7348);
or U7936 (N_7936,N_7230,N_7086);
xor U7937 (N_7937,N_7168,N_7209);
and U7938 (N_7938,N_7056,N_7126);
xor U7939 (N_7939,N_7360,N_7431);
nand U7940 (N_7940,N_7007,N_7185);
nand U7941 (N_7941,N_7038,N_7016);
or U7942 (N_7942,N_7433,N_7228);
nor U7943 (N_7943,N_7433,N_7040);
and U7944 (N_7944,N_7143,N_7192);
xnor U7945 (N_7945,N_7010,N_7125);
xnor U7946 (N_7946,N_7437,N_7153);
nand U7947 (N_7947,N_7061,N_7013);
nor U7948 (N_7948,N_7213,N_7077);
nand U7949 (N_7949,N_7086,N_7066);
xnor U7950 (N_7950,N_7280,N_7044);
or U7951 (N_7951,N_7475,N_7409);
nor U7952 (N_7952,N_7144,N_7016);
nor U7953 (N_7953,N_7127,N_7025);
xor U7954 (N_7954,N_7025,N_7106);
nor U7955 (N_7955,N_7097,N_7071);
or U7956 (N_7956,N_7269,N_7478);
xor U7957 (N_7957,N_7286,N_7031);
nor U7958 (N_7958,N_7131,N_7314);
and U7959 (N_7959,N_7008,N_7352);
nand U7960 (N_7960,N_7430,N_7329);
nand U7961 (N_7961,N_7171,N_7423);
or U7962 (N_7962,N_7199,N_7392);
or U7963 (N_7963,N_7467,N_7136);
or U7964 (N_7964,N_7334,N_7492);
or U7965 (N_7965,N_7228,N_7023);
xor U7966 (N_7966,N_7164,N_7264);
nand U7967 (N_7967,N_7349,N_7040);
and U7968 (N_7968,N_7053,N_7073);
or U7969 (N_7969,N_7100,N_7366);
xnor U7970 (N_7970,N_7271,N_7194);
nor U7971 (N_7971,N_7102,N_7448);
or U7972 (N_7972,N_7445,N_7133);
nor U7973 (N_7973,N_7082,N_7336);
and U7974 (N_7974,N_7444,N_7454);
nand U7975 (N_7975,N_7184,N_7180);
and U7976 (N_7976,N_7143,N_7285);
nand U7977 (N_7977,N_7244,N_7270);
nor U7978 (N_7978,N_7352,N_7450);
and U7979 (N_7979,N_7467,N_7044);
xnor U7980 (N_7980,N_7350,N_7356);
nand U7981 (N_7981,N_7003,N_7065);
nand U7982 (N_7982,N_7337,N_7367);
or U7983 (N_7983,N_7297,N_7007);
xor U7984 (N_7984,N_7415,N_7218);
xor U7985 (N_7985,N_7099,N_7093);
nor U7986 (N_7986,N_7054,N_7400);
or U7987 (N_7987,N_7014,N_7216);
and U7988 (N_7988,N_7151,N_7030);
nor U7989 (N_7989,N_7063,N_7259);
xnor U7990 (N_7990,N_7223,N_7447);
or U7991 (N_7991,N_7451,N_7358);
nor U7992 (N_7992,N_7082,N_7469);
or U7993 (N_7993,N_7216,N_7325);
or U7994 (N_7994,N_7447,N_7310);
and U7995 (N_7995,N_7252,N_7100);
nor U7996 (N_7996,N_7415,N_7174);
and U7997 (N_7997,N_7095,N_7043);
nor U7998 (N_7998,N_7186,N_7293);
nand U7999 (N_7999,N_7449,N_7257);
nor U8000 (N_8000,N_7756,N_7507);
or U8001 (N_8001,N_7557,N_7747);
nor U8002 (N_8002,N_7834,N_7519);
nor U8003 (N_8003,N_7993,N_7816);
or U8004 (N_8004,N_7535,N_7994);
nand U8005 (N_8005,N_7788,N_7828);
or U8006 (N_8006,N_7934,N_7527);
and U8007 (N_8007,N_7639,N_7784);
and U8008 (N_8008,N_7667,N_7549);
or U8009 (N_8009,N_7746,N_7678);
xnor U8010 (N_8010,N_7524,N_7745);
and U8011 (N_8011,N_7712,N_7805);
and U8012 (N_8012,N_7655,N_7677);
or U8013 (N_8013,N_7670,N_7932);
and U8014 (N_8014,N_7744,N_7986);
nor U8015 (N_8015,N_7806,N_7763);
and U8016 (N_8016,N_7701,N_7915);
and U8017 (N_8017,N_7928,N_7841);
xor U8018 (N_8018,N_7778,N_7869);
xnor U8019 (N_8019,N_7888,N_7774);
nor U8020 (N_8020,N_7919,N_7975);
nand U8021 (N_8021,N_7553,N_7521);
and U8022 (N_8022,N_7573,N_7815);
nand U8023 (N_8023,N_7617,N_7679);
or U8024 (N_8024,N_7540,N_7939);
and U8025 (N_8025,N_7562,N_7983);
and U8026 (N_8026,N_7623,N_7558);
nand U8027 (N_8027,N_7689,N_7593);
nor U8028 (N_8028,N_7675,N_7742);
xor U8029 (N_8029,N_7965,N_7637);
or U8030 (N_8030,N_7785,N_7950);
xnor U8031 (N_8031,N_7614,N_7587);
or U8032 (N_8032,N_7613,N_7804);
and U8033 (N_8033,N_7879,N_7810);
nor U8034 (N_8034,N_7567,N_7578);
xnor U8035 (N_8035,N_7631,N_7911);
nor U8036 (N_8036,N_7596,N_7657);
nor U8037 (N_8037,N_7964,N_7510);
nor U8038 (N_8038,N_7793,N_7990);
and U8039 (N_8039,N_7846,N_7699);
nand U8040 (N_8040,N_7982,N_7594);
nand U8041 (N_8041,N_7548,N_7731);
and U8042 (N_8042,N_7538,N_7737);
xnor U8043 (N_8043,N_7904,N_7545);
nand U8044 (N_8044,N_7800,N_7999);
or U8045 (N_8045,N_7766,N_7839);
and U8046 (N_8046,N_7760,N_7612);
nor U8047 (N_8047,N_7901,N_7768);
nor U8048 (N_8048,N_7843,N_7781);
or U8049 (N_8049,N_7948,N_7798);
or U8050 (N_8050,N_7516,N_7571);
nand U8051 (N_8051,N_7925,N_7807);
xor U8052 (N_8052,N_7970,N_7917);
nand U8053 (N_8053,N_7875,N_7977);
or U8054 (N_8054,N_7650,N_7971);
and U8055 (N_8055,N_7876,N_7542);
nand U8056 (N_8056,N_7674,N_7634);
or U8057 (N_8057,N_7811,N_7642);
or U8058 (N_8058,N_7752,N_7695);
and U8059 (N_8059,N_7974,N_7830);
nor U8060 (N_8060,N_7987,N_7600);
nor U8061 (N_8061,N_7802,N_7561);
or U8062 (N_8062,N_7621,N_7660);
xnor U8063 (N_8063,N_7889,N_7525);
and U8064 (N_8064,N_7543,N_7606);
nor U8065 (N_8065,N_7855,N_7690);
nor U8066 (N_8066,N_7880,N_7622);
or U8067 (N_8067,N_7503,N_7592);
nor U8068 (N_8068,N_7933,N_7653);
nor U8069 (N_8069,N_7887,N_7582);
or U8070 (N_8070,N_7603,N_7685);
nand U8071 (N_8071,N_7898,N_7743);
nor U8072 (N_8072,N_7936,N_7908);
xor U8073 (N_8073,N_7814,N_7619);
nor U8074 (N_8074,N_7905,N_7555);
xor U8075 (N_8075,N_7691,N_7513);
and U8076 (N_8076,N_7852,N_7820);
nor U8077 (N_8077,N_7803,N_7520);
and U8078 (N_8078,N_7626,N_7570);
or U8079 (N_8079,N_7597,N_7709);
or U8080 (N_8080,N_7514,N_7770);
nand U8081 (N_8081,N_7552,N_7539);
nand U8082 (N_8082,N_7884,N_7668);
and U8083 (N_8083,N_7515,N_7713);
nor U8084 (N_8084,N_7837,N_7794);
and U8085 (N_8085,N_7604,N_7892);
or U8086 (N_8086,N_7676,N_7844);
or U8087 (N_8087,N_7651,N_7707);
and U8088 (N_8088,N_7568,N_7808);
nand U8089 (N_8089,N_7824,N_7862);
or U8090 (N_8090,N_7534,N_7981);
and U8091 (N_8091,N_7995,N_7696);
nor U8092 (N_8092,N_7686,N_7681);
or U8093 (N_8093,N_7938,N_7704);
or U8094 (N_8094,N_7969,N_7511);
xnor U8095 (N_8095,N_7636,N_7792);
nand U8096 (N_8096,N_7789,N_7740);
nand U8097 (N_8097,N_7702,N_7959);
or U8098 (N_8098,N_7847,N_7845);
xnor U8099 (N_8099,N_7705,N_7903);
xor U8100 (N_8100,N_7818,N_7758);
nor U8101 (N_8101,N_7899,N_7790);
nor U8102 (N_8102,N_7656,N_7868);
nand U8103 (N_8103,N_7663,N_7733);
and U8104 (N_8104,N_7501,N_7652);
and U8105 (N_8105,N_7937,N_7698);
nand U8106 (N_8106,N_7963,N_7585);
xnor U8107 (N_8107,N_7550,N_7978);
nor U8108 (N_8108,N_7502,N_7536);
nor U8109 (N_8109,N_7867,N_7769);
xor U8110 (N_8110,N_7836,N_7997);
nand U8111 (N_8111,N_7627,N_7608);
nand U8112 (N_8112,N_7533,N_7941);
and U8113 (N_8113,N_7711,N_7863);
nand U8114 (N_8114,N_7755,N_7838);
or U8115 (N_8115,N_7649,N_7753);
xor U8116 (N_8116,N_7882,N_7878);
nand U8117 (N_8117,N_7710,N_7894);
and U8118 (N_8118,N_7916,N_7574);
and U8119 (N_8119,N_7735,N_7902);
or U8120 (N_8120,N_7881,N_7706);
or U8121 (N_8121,N_7508,N_7909);
and U8122 (N_8122,N_7598,N_7942);
nor U8123 (N_8123,N_7773,N_7833);
or U8124 (N_8124,N_7559,N_7835);
xnor U8125 (N_8125,N_7547,N_7541);
or U8126 (N_8126,N_7730,N_7727);
and U8127 (N_8127,N_7641,N_7854);
or U8128 (N_8128,N_7813,N_7715);
or U8129 (N_8129,N_7998,N_7732);
nor U8130 (N_8130,N_7584,N_7777);
and U8131 (N_8131,N_7840,N_7851);
or U8132 (N_8132,N_7849,N_7958);
nor U8133 (N_8133,N_7703,N_7683);
xor U8134 (N_8134,N_7771,N_7762);
or U8135 (N_8135,N_7967,N_7864);
xnor U8136 (N_8136,N_7848,N_7962);
nand U8137 (N_8137,N_7628,N_7692);
or U8138 (N_8138,N_7616,N_7826);
nor U8139 (N_8139,N_7748,N_7946);
nor U8140 (N_8140,N_7923,N_7522);
nor U8141 (N_8141,N_7662,N_7754);
nor U8142 (N_8142,N_7858,N_7544);
or U8143 (N_8143,N_7504,N_7554);
nor U8144 (N_8144,N_7989,N_7687);
and U8145 (N_8145,N_7643,N_7607);
or U8146 (N_8146,N_7796,N_7575);
nor U8147 (N_8147,N_7896,N_7609);
xor U8148 (N_8148,N_7821,N_7883);
nor U8149 (N_8149,N_7610,N_7947);
nor U8150 (N_8150,N_7688,N_7960);
nand U8151 (N_8151,N_7801,N_7684);
nand U8152 (N_8152,N_7890,N_7629);
and U8153 (N_8153,N_7996,N_7611);
nor U8154 (N_8154,N_7531,N_7669);
nor U8155 (N_8155,N_7556,N_7640);
nor U8156 (N_8156,N_7759,N_7595);
nor U8157 (N_8157,N_7586,N_7924);
and U8158 (N_8158,N_7772,N_7625);
and U8159 (N_8159,N_7935,N_7783);
or U8160 (N_8160,N_7955,N_7832);
nand U8161 (N_8161,N_7865,N_7500);
xor U8162 (N_8162,N_7786,N_7659);
or U8163 (N_8163,N_7647,N_7985);
xor U8164 (N_8164,N_7871,N_7900);
nand U8165 (N_8165,N_7966,N_7723);
and U8166 (N_8166,N_7749,N_7661);
and U8167 (N_8167,N_7700,N_7589);
or U8168 (N_8168,N_7529,N_7856);
nand U8169 (N_8169,N_7714,N_7968);
nor U8170 (N_8170,N_7927,N_7718);
nand U8171 (N_8171,N_7775,N_7873);
nand U8172 (N_8172,N_7734,N_7633);
nor U8173 (N_8173,N_7954,N_7601);
nor U8174 (N_8174,N_7819,N_7726);
nor U8175 (N_8175,N_7877,N_7644);
xor U8176 (N_8176,N_7861,N_7591);
and U8177 (N_8177,N_7931,N_7918);
nor U8178 (N_8178,N_7929,N_7823);
nor U8179 (N_8179,N_7646,N_7664);
nand U8180 (N_8180,N_7635,N_7886);
and U8181 (N_8181,N_7817,N_7782);
or U8182 (N_8182,N_7630,N_7870);
nor U8183 (N_8183,N_7741,N_7913);
or U8184 (N_8184,N_7827,N_7665);
or U8185 (N_8185,N_7728,N_7729);
xnor U8186 (N_8186,N_7523,N_7588);
or U8187 (N_8187,N_7565,N_7648);
or U8188 (N_8188,N_7615,N_7885);
xnor U8189 (N_8189,N_7654,N_7984);
or U8190 (N_8190,N_7551,N_7672);
or U8191 (N_8191,N_7682,N_7632);
xnor U8192 (N_8192,N_7859,N_7512);
nor U8193 (N_8193,N_7724,N_7618);
nand U8194 (N_8194,N_7895,N_7951);
nand U8195 (N_8195,N_7509,N_7751);
nand U8196 (N_8196,N_7893,N_7949);
nor U8197 (N_8197,N_7767,N_7776);
and U8198 (N_8198,N_7590,N_7853);
and U8199 (N_8199,N_7973,N_7576);
nor U8200 (N_8200,N_7795,N_7972);
nor U8201 (N_8201,N_7638,N_7693);
and U8202 (N_8202,N_7906,N_7528);
xnor U8203 (N_8203,N_7765,N_7812);
and U8204 (N_8204,N_7722,N_7566);
and U8205 (N_8205,N_7779,N_7572);
or U8206 (N_8206,N_7857,N_7988);
and U8207 (N_8207,N_7721,N_7897);
and U8208 (N_8208,N_7944,N_7658);
or U8209 (N_8209,N_7530,N_7526);
nor U8210 (N_8210,N_7992,N_7860);
or U8211 (N_8211,N_7563,N_7505);
and U8212 (N_8212,N_7953,N_7922);
and U8213 (N_8213,N_7940,N_7952);
or U8214 (N_8214,N_7738,N_7930);
nand U8215 (N_8215,N_7716,N_7506);
nor U8216 (N_8216,N_7797,N_7787);
nor U8217 (N_8217,N_7957,N_7912);
nand U8218 (N_8218,N_7825,N_7891);
or U8219 (N_8219,N_7680,N_7874);
nor U8220 (N_8220,N_7569,N_7581);
nor U8221 (N_8221,N_7809,N_7914);
and U8222 (N_8222,N_7850,N_7872);
or U8223 (N_8223,N_7920,N_7829);
and U8224 (N_8224,N_7673,N_7945);
nand U8225 (N_8225,N_7697,N_7991);
nand U8226 (N_8226,N_7910,N_7750);
nor U8227 (N_8227,N_7671,N_7645);
and U8228 (N_8228,N_7943,N_7518);
or U8229 (N_8229,N_7799,N_7620);
nor U8230 (N_8230,N_7546,N_7907);
xor U8231 (N_8231,N_7757,N_7532);
xor U8232 (N_8232,N_7822,N_7580);
and U8233 (N_8233,N_7842,N_7761);
and U8234 (N_8234,N_7831,N_7708);
or U8235 (N_8235,N_7564,N_7739);
xor U8236 (N_8236,N_7720,N_7921);
nor U8237 (N_8237,N_7624,N_7926);
nor U8238 (N_8238,N_7717,N_7666);
xor U8239 (N_8239,N_7780,N_7605);
xor U8240 (N_8240,N_7599,N_7517);
nand U8241 (N_8241,N_7694,N_7980);
nand U8242 (N_8242,N_7976,N_7736);
xnor U8243 (N_8243,N_7961,N_7956);
or U8244 (N_8244,N_7719,N_7979);
xor U8245 (N_8245,N_7866,N_7725);
and U8246 (N_8246,N_7560,N_7764);
xor U8247 (N_8247,N_7602,N_7577);
nand U8248 (N_8248,N_7537,N_7791);
or U8249 (N_8249,N_7583,N_7579);
or U8250 (N_8250,N_7842,N_7610);
nand U8251 (N_8251,N_7527,N_7567);
xor U8252 (N_8252,N_7665,N_7876);
or U8253 (N_8253,N_7896,N_7562);
and U8254 (N_8254,N_7952,N_7908);
nand U8255 (N_8255,N_7921,N_7582);
xor U8256 (N_8256,N_7720,N_7761);
xor U8257 (N_8257,N_7821,N_7558);
nor U8258 (N_8258,N_7709,N_7860);
xor U8259 (N_8259,N_7855,N_7546);
xnor U8260 (N_8260,N_7997,N_7904);
or U8261 (N_8261,N_7500,N_7862);
xnor U8262 (N_8262,N_7843,N_7729);
and U8263 (N_8263,N_7553,N_7838);
or U8264 (N_8264,N_7672,N_7987);
nor U8265 (N_8265,N_7800,N_7998);
and U8266 (N_8266,N_7832,N_7810);
xnor U8267 (N_8267,N_7716,N_7992);
nor U8268 (N_8268,N_7852,N_7613);
xnor U8269 (N_8269,N_7837,N_7683);
nor U8270 (N_8270,N_7808,N_7690);
xor U8271 (N_8271,N_7559,N_7787);
nand U8272 (N_8272,N_7734,N_7951);
xnor U8273 (N_8273,N_7951,N_7749);
nor U8274 (N_8274,N_7975,N_7961);
nor U8275 (N_8275,N_7711,N_7621);
xnor U8276 (N_8276,N_7649,N_7987);
nand U8277 (N_8277,N_7900,N_7848);
nor U8278 (N_8278,N_7881,N_7900);
nor U8279 (N_8279,N_7955,N_7506);
xor U8280 (N_8280,N_7920,N_7854);
or U8281 (N_8281,N_7882,N_7976);
nor U8282 (N_8282,N_7981,N_7781);
xor U8283 (N_8283,N_7711,N_7527);
or U8284 (N_8284,N_7948,N_7819);
or U8285 (N_8285,N_7721,N_7772);
nor U8286 (N_8286,N_7920,N_7706);
nor U8287 (N_8287,N_7781,N_7865);
or U8288 (N_8288,N_7606,N_7615);
nor U8289 (N_8289,N_7605,N_7760);
nand U8290 (N_8290,N_7890,N_7990);
or U8291 (N_8291,N_7775,N_7909);
or U8292 (N_8292,N_7860,N_7786);
or U8293 (N_8293,N_7878,N_7573);
nor U8294 (N_8294,N_7606,N_7854);
xnor U8295 (N_8295,N_7597,N_7551);
and U8296 (N_8296,N_7599,N_7740);
and U8297 (N_8297,N_7718,N_7903);
or U8298 (N_8298,N_7996,N_7766);
xor U8299 (N_8299,N_7672,N_7601);
or U8300 (N_8300,N_7943,N_7650);
and U8301 (N_8301,N_7725,N_7854);
and U8302 (N_8302,N_7635,N_7715);
or U8303 (N_8303,N_7599,N_7967);
and U8304 (N_8304,N_7985,N_7610);
nand U8305 (N_8305,N_7954,N_7668);
nor U8306 (N_8306,N_7723,N_7631);
or U8307 (N_8307,N_7602,N_7777);
or U8308 (N_8308,N_7535,N_7884);
nand U8309 (N_8309,N_7756,N_7792);
nand U8310 (N_8310,N_7597,N_7994);
nand U8311 (N_8311,N_7955,N_7522);
xor U8312 (N_8312,N_7671,N_7786);
or U8313 (N_8313,N_7794,N_7559);
nor U8314 (N_8314,N_7532,N_7662);
and U8315 (N_8315,N_7766,N_7908);
nand U8316 (N_8316,N_7666,N_7677);
xor U8317 (N_8317,N_7720,N_7597);
or U8318 (N_8318,N_7922,N_7504);
and U8319 (N_8319,N_7758,N_7919);
xnor U8320 (N_8320,N_7593,N_7909);
and U8321 (N_8321,N_7688,N_7959);
and U8322 (N_8322,N_7897,N_7681);
xnor U8323 (N_8323,N_7939,N_7815);
nor U8324 (N_8324,N_7890,N_7680);
and U8325 (N_8325,N_7636,N_7586);
nor U8326 (N_8326,N_7614,N_7928);
or U8327 (N_8327,N_7965,N_7565);
nand U8328 (N_8328,N_7595,N_7643);
or U8329 (N_8329,N_7527,N_7820);
nor U8330 (N_8330,N_7629,N_7924);
and U8331 (N_8331,N_7935,N_7535);
xor U8332 (N_8332,N_7633,N_7590);
xor U8333 (N_8333,N_7931,N_7900);
nor U8334 (N_8334,N_7637,N_7906);
or U8335 (N_8335,N_7591,N_7533);
nor U8336 (N_8336,N_7912,N_7703);
nand U8337 (N_8337,N_7625,N_7650);
or U8338 (N_8338,N_7555,N_7919);
and U8339 (N_8339,N_7569,N_7757);
and U8340 (N_8340,N_7870,N_7813);
or U8341 (N_8341,N_7502,N_7682);
nor U8342 (N_8342,N_7546,N_7961);
or U8343 (N_8343,N_7666,N_7563);
nand U8344 (N_8344,N_7997,N_7527);
and U8345 (N_8345,N_7937,N_7837);
or U8346 (N_8346,N_7686,N_7633);
xnor U8347 (N_8347,N_7569,N_7658);
nor U8348 (N_8348,N_7761,N_7789);
xnor U8349 (N_8349,N_7771,N_7538);
nor U8350 (N_8350,N_7614,N_7541);
nand U8351 (N_8351,N_7554,N_7807);
nor U8352 (N_8352,N_7962,N_7521);
xor U8353 (N_8353,N_7866,N_7975);
nor U8354 (N_8354,N_7981,N_7921);
xor U8355 (N_8355,N_7826,N_7892);
nor U8356 (N_8356,N_7971,N_7968);
nor U8357 (N_8357,N_7807,N_7687);
or U8358 (N_8358,N_7528,N_7691);
nor U8359 (N_8359,N_7904,N_7890);
nor U8360 (N_8360,N_7529,N_7590);
nor U8361 (N_8361,N_7798,N_7739);
xnor U8362 (N_8362,N_7699,N_7509);
and U8363 (N_8363,N_7619,N_7502);
xor U8364 (N_8364,N_7662,N_7833);
and U8365 (N_8365,N_7518,N_7662);
xnor U8366 (N_8366,N_7736,N_7969);
xor U8367 (N_8367,N_7856,N_7760);
nor U8368 (N_8368,N_7899,N_7771);
nor U8369 (N_8369,N_7623,N_7572);
and U8370 (N_8370,N_7743,N_7983);
xnor U8371 (N_8371,N_7874,N_7904);
xor U8372 (N_8372,N_7859,N_7544);
xnor U8373 (N_8373,N_7965,N_7906);
and U8374 (N_8374,N_7791,N_7629);
or U8375 (N_8375,N_7706,N_7786);
or U8376 (N_8376,N_7506,N_7824);
and U8377 (N_8377,N_7676,N_7930);
xor U8378 (N_8378,N_7773,N_7614);
nor U8379 (N_8379,N_7521,N_7855);
nand U8380 (N_8380,N_7692,N_7620);
and U8381 (N_8381,N_7947,N_7970);
nand U8382 (N_8382,N_7535,N_7745);
or U8383 (N_8383,N_7580,N_7984);
and U8384 (N_8384,N_7626,N_7530);
nor U8385 (N_8385,N_7892,N_7580);
or U8386 (N_8386,N_7889,N_7621);
nand U8387 (N_8387,N_7743,N_7904);
or U8388 (N_8388,N_7831,N_7775);
nand U8389 (N_8389,N_7978,N_7990);
xnor U8390 (N_8390,N_7638,N_7842);
and U8391 (N_8391,N_7575,N_7809);
or U8392 (N_8392,N_7919,N_7677);
xnor U8393 (N_8393,N_7594,N_7510);
or U8394 (N_8394,N_7530,N_7519);
nand U8395 (N_8395,N_7706,N_7503);
or U8396 (N_8396,N_7737,N_7536);
xnor U8397 (N_8397,N_7799,N_7717);
xnor U8398 (N_8398,N_7770,N_7685);
nor U8399 (N_8399,N_7591,N_7914);
xor U8400 (N_8400,N_7532,N_7673);
or U8401 (N_8401,N_7558,N_7537);
xnor U8402 (N_8402,N_7709,N_7621);
and U8403 (N_8403,N_7652,N_7963);
xor U8404 (N_8404,N_7851,N_7573);
nand U8405 (N_8405,N_7944,N_7592);
or U8406 (N_8406,N_7851,N_7710);
nand U8407 (N_8407,N_7584,N_7969);
or U8408 (N_8408,N_7762,N_7642);
nand U8409 (N_8409,N_7505,N_7922);
xor U8410 (N_8410,N_7869,N_7689);
xnor U8411 (N_8411,N_7817,N_7952);
or U8412 (N_8412,N_7572,N_7787);
and U8413 (N_8413,N_7765,N_7731);
nor U8414 (N_8414,N_7581,N_7735);
nand U8415 (N_8415,N_7798,N_7869);
nor U8416 (N_8416,N_7974,N_7949);
nand U8417 (N_8417,N_7725,N_7699);
or U8418 (N_8418,N_7963,N_7561);
and U8419 (N_8419,N_7540,N_7970);
xnor U8420 (N_8420,N_7760,N_7708);
or U8421 (N_8421,N_7535,N_7870);
or U8422 (N_8422,N_7714,N_7983);
nor U8423 (N_8423,N_7606,N_7995);
nor U8424 (N_8424,N_7758,N_7634);
nor U8425 (N_8425,N_7832,N_7807);
and U8426 (N_8426,N_7585,N_7650);
or U8427 (N_8427,N_7653,N_7947);
nand U8428 (N_8428,N_7540,N_7749);
nor U8429 (N_8429,N_7601,N_7526);
nand U8430 (N_8430,N_7575,N_7623);
nor U8431 (N_8431,N_7916,N_7585);
and U8432 (N_8432,N_7624,N_7985);
or U8433 (N_8433,N_7936,N_7505);
xnor U8434 (N_8434,N_7729,N_7702);
and U8435 (N_8435,N_7797,N_7984);
and U8436 (N_8436,N_7752,N_7970);
or U8437 (N_8437,N_7581,N_7854);
and U8438 (N_8438,N_7728,N_7504);
or U8439 (N_8439,N_7884,N_7630);
or U8440 (N_8440,N_7763,N_7577);
nor U8441 (N_8441,N_7806,N_7988);
nor U8442 (N_8442,N_7864,N_7602);
and U8443 (N_8443,N_7654,N_7825);
nor U8444 (N_8444,N_7924,N_7891);
nand U8445 (N_8445,N_7911,N_7727);
xor U8446 (N_8446,N_7541,N_7654);
nand U8447 (N_8447,N_7827,N_7957);
nand U8448 (N_8448,N_7559,N_7764);
and U8449 (N_8449,N_7968,N_7532);
nor U8450 (N_8450,N_7632,N_7516);
nand U8451 (N_8451,N_7852,N_7623);
nor U8452 (N_8452,N_7983,N_7803);
nand U8453 (N_8453,N_7611,N_7699);
or U8454 (N_8454,N_7548,N_7691);
or U8455 (N_8455,N_7923,N_7857);
xnor U8456 (N_8456,N_7617,N_7707);
nand U8457 (N_8457,N_7855,N_7649);
or U8458 (N_8458,N_7546,N_7899);
nor U8459 (N_8459,N_7637,N_7602);
and U8460 (N_8460,N_7845,N_7890);
or U8461 (N_8461,N_7950,N_7775);
or U8462 (N_8462,N_7888,N_7703);
and U8463 (N_8463,N_7799,N_7760);
nor U8464 (N_8464,N_7620,N_7682);
and U8465 (N_8465,N_7647,N_7794);
xor U8466 (N_8466,N_7634,N_7867);
xor U8467 (N_8467,N_7749,N_7739);
and U8468 (N_8468,N_7954,N_7901);
nor U8469 (N_8469,N_7500,N_7889);
and U8470 (N_8470,N_7863,N_7924);
nor U8471 (N_8471,N_7523,N_7632);
nand U8472 (N_8472,N_7791,N_7825);
or U8473 (N_8473,N_7930,N_7928);
nor U8474 (N_8474,N_7744,N_7592);
nand U8475 (N_8475,N_7619,N_7909);
xnor U8476 (N_8476,N_7576,N_7838);
or U8477 (N_8477,N_7981,N_7644);
and U8478 (N_8478,N_7642,N_7904);
or U8479 (N_8479,N_7979,N_7696);
nor U8480 (N_8480,N_7809,N_7762);
nand U8481 (N_8481,N_7805,N_7547);
xor U8482 (N_8482,N_7838,N_7794);
or U8483 (N_8483,N_7769,N_7845);
nand U8484 (N_8484,N_7985,N_7644);
xnor U8485 (N_8485,N_7501,N_7556);
and U8486 (N_8486,N_7865,N_7550);
xnor U8487 (N_8487,N_7837,N_7553);
and U8488 (N_8488,N_7719,N_7677);
nor U8489 (N_8489,N_7931,N_7994);
xor U8490 (N_8490,N_7768,N_7762);
or U8491 (N_8491,N_7867,N_7640);
nand U8492 (N_8492,N_7709,N_7538);
and U8493 (N_8493,N_7878,N_7783);
and U8494 (N_8494,N_7733,N_7834);
and U8495 (N_8495,N_7523,N_7972);
xnor U8496 (N_8496,N_7527,N_7550);
xnor U8497 (N_8497,N_7557,N_7739);
or U8498 (N_8498,N_7842,N_7501);
or U8499 (N_8499,N_7969,N_7760);
nand U8500 (N_8500,N_8013,N_8147);
xnor U8501 (N_8501,N_8202,N_8314);
or U8502 (N_8502,N_8040,N_8459);
and U8503 (N_8503,N_8135,N_8364);
nor U8504 (N_8504,N_8282,N_8145);
nand U8505 (N_8505,N_8144,N_8227);
nor U8506 (N_8506,N_8468,N_8067);
or U8507 (N_8507,N_8212,N_8425);
xor U8508 (N_8508,N_8204,N_8396);
and U8509 (N_8509,N_8035,N_8229);
nand U8510 (N_8510,N_8262,N_8061);
nand U8511 (N_8511,N_8426,N_8276);
and U8512 (N_8512,N_8255,N_8194);
and U8513 (N_8513,N_8087,N_8449);
or U8514 (N_8514,N_8153,N_8011);
and U8515 (N_8515,N_8402,N_8301);
and U8516 (N_8516,N_8384,N_8029);
or U8517 (N_8517,N_8018,N_8234);
nor U8518 (N_8518,N_8043,N_8116);
and U8519 (N_8519,N_8217,N_8454);
xor U8520 (N_8520,N_8092,N_8272);
xor U8521 (N_8521,N_8333,N_8342);
nor U8522 (N_8522,N_8407,N_8466);
and U8523 (N_8523,N_8334,N_8039);
xor U8524 (N_8524,N_8437,N_8486);
nor U8525 (N_8525,N_8123,N_8027);
or U8526 (N_8526,N_8286,N_8237);
nor U8527 (N_8527,N_8455,N_8481);
and U8528 (N_8528,N_8440,N_8177);
xnor U8529 (N_8529,N_8496,N_8274);
xnor U8530 (N_8530,N_8424,N_8076);
nor U8531 (N_8531,N_8347,N_8370);
nand U8532 (N_8532,N_8383,N_8081);
or U8533 (N_8533,N_8290,N_8288);
or U8534 (N_8534,N_8253,N_8193);
nand U8535 (N_8535,N_8242,N_8281);
or U8536 (N_8536,N_8054,N_8287);
nand U8537 (N_8537,N_8125,N_8256);
and U8538 (N_8538,N_8138,N_8353);
nand U8539 (N_8539,N_8430,N_8474);
nand U8540 (N_8540,N_8360,N_8317);
and U8541 (N_8541,N_8016,N_8167);
nor U8542 (N_8542,N_8012,N_8351);
nor U8543 (N_8543,N_8379,N_8192);
nand U8544 (N_8544,N_8032,N_8085);
xnor U8545 (N_8545,N_8302,N_8431);
xor U8546 (N_8546,N_8448,N_8289);
and U8547 (N_8547,N_8278,N_8174);
and U8548 (N_8548,N_8355,N_8093);
xor U8549 (N_8549,N_8099,N_8291);
or U8550 (N_8550,N_8005,N_8017);
nor U8551 (N_8551,N_8419,N_8120);
nand U8552 (N_8552,N_8443,N_8000);
nor U8553 (N_8553,N_8015,N_8221);
and U8554 (N_8554,N_8470,N_8042);
and U8555 (N_8555,N_8456,N_8298);
and U8556 (N_8556,N_8075,N_8141);
nor U8557 (N_8557,N_8423,N_8339);
or U8558 (N_8558,N_8079,N_8063);
nor U8559 (N_8559,N_8416,N_8247);
and U8560 (N_8560,N_8445,N_8241);
or U8561 (N_8561,N_8306,N_8166);
nor U8562 (N_8562,N_8300,N_8332);
or U8563 (N_8563,N_8315,N_8258);
or U8564 (N_8564,N_8374,N_8422);
xor U8565 (N_8565,N_8393,N_8146);
xnor U8566 (N_8566,N_8435,N_8080);
nand U8567 (N_8567,N_8411,N_8223);
xnor U8568 (N_8568,N_8238,N_8205);
and U8569 (N_8569,N_8464,N_8140);
or U8570 (N_8570,N_8324,N_8378);
and U8571 (N_8571,N_8284,N_8121);
nor U8572 (N_8572,N_8127,N_8451);
or U8573 (N_8573,N_8312,N_8458);
xnor U8574 (N_8574,N_8152,N_8463);
nor U8575 (N_8575,N_8235,N_8338);
xor U8576 (N_8576,N_8248,N_8206);
or U8577 (N_8577,N_8006,N_8348);
nand U8578 (N_8578,N_8483,N_8354);
and U8579 (N_8579,N_8077,N_8465);
nor U8580 (N_8580,N_8260,N_8283);
xor U8581 (N_8581,N_8294,N_8047);
or U8582 (N_8582,N_8088,N_8444);
nor U8583 (N_8583,N_8219,N_8335);
xor U8584 (N_8584,N_8429,N_8110);
xnor U8585 (N_8585,N_8002,N_8408);
xnor U8586 (N_8586,N_8400,N_8263);
nor U8587 (N_8587,N_8178,N_8210);
or U8588 (N_8588,N_8213,N_8363);
xor U8589 (N_8589,N_8420,N_8494);
and U8590 (N_8590,N_8475,N_8112);
or U8591 (N_8591,N_8367,N_8139);
nand U8592 (N_8592,N_8115,N_8478);
xor U8593 (N_8593,N_8059,N_8498);
and U8594 (N_8594,N_8190,N_8183);
and U8595 (N_8595,N_8296,N_8074);
or U8596 (N_8596,N_8195,N_8180);
nand U8597 (N_8597,N_8409,N_8009);
and U8598 (N_8598,N_8482,N_8182);
nand U8599 (N_8599,N_8095,N_8410);
xnor U8600 (N_8600,N_8479,N_8169);
xnor U8601 (N_8601,N_8053,N_8428);
nand U8602 (N_8602,N_8391,N_8057);
nor U8603 (N_8603,N_8490,N_8421);
nor U8604 (N_8604,N_8239,N_8215);
xnor U8605 (N_8605,N_8472,N_8022);
nor U8606 (N_8606,N_8325,N_8297);
nand U8607 (N_8607,N_8129,N_8196);
or U8608 (N_8608,N_8028,N_8280);
nor U8609 (N_8609,N_8025,N_8091);
xnor U8610 (N_8610,N_8222,N_8181);
nand U8611 (N_8611,N_8102,N_8062);
or U8612 (N_8612,N_8014,N_8020);
and U8613 (N_8613,N_8154,N_8151);
or U8614 (N_8614,N_8341,N_8362);
nand U8615 (N_8615,N_8089,N_8251);
and U8616 (N_8616,N_8436,N_8148);
xnor U8617 (N_8617,N_8450,N_8390);
and U8618 (N_8618,N_8292,N_8208);
or U8619 (N_8619,N_8403,N_8070);
nand U8620 (N_8620,N_8230,N_8111);
or U8621 (N_8621,N_8173,N_8082);
and U8622 (N_8622,N_8398,N_8031);
xor U8623 (N_8623,N_8069,N_8316);
nor U8624 (N_8624,N_8279,N_8249);
or U8625 (N_8625,N_8343,N_8244);
xnor U8626 (N_8626,N_8228,N_8160);
xor U8627 (N_8627,N_8149,N_8476);
and U8628 (N_8628,N_8240,N_8376);
nor U8629 (N_8629,N_8264,N_8285);
and U8630 (N_8630,N_8184,N_8245);
nand U8631 (N_8631,N_8049,N_8023);
xnor U8632 (N_8632,N_8096,N_8224);
nand U8633 (N_8633,N_8107,N_8392);
and U8634 (N_8634,N_8377,N_8344);
xnor U8635 (N_8635,N_8488,N_8331);
and U8636 (N_8636,N_8055,N_8101);
and U8637 (N_8637,N_8133,N_8467);
and U8638 (N_8638,N_8188,N_8433);
or U8639 (N_8639,N_8446,N_8124);
xor U8640 (N_8640,N_8083,N_8480);
or U8641 (N_8641,N_8381,N_8243);
nand U8642 (N_8642,N_8405,N_8322);
and U8643 (N_8643,N_8484,N_8220);
or U8644 (N_8644,N_8457,N_8113);
nand U8645 (N_8645,N_8037,N_8293);
xor U8646 (N_8646,N_8257,N_8350);
and U8647 (N_8647,N_8492,N_8261);
or U8648 (N_8648,N_8368,N_8313);
nor U8649 (N_8649,N_8214,N_8216);
nand U8650 (N_8650,N_8303,N_8375);
and U8651 (N_8651,N_8162,N_8345);
xor U8652 (N_8652,N_8318,N_8019);
nor U8653 (N_8653,N_8386,N_8199);
xnor U8654 (N_8654,N_8186,N_8265);
nor U8655 (N_8655,N_8060,N_8106);
nand U8656 (N_8656,N_8485,N_8136);
nor U8657 (N_8657,N_8010,N_8109);
nor U8658 (N_8658,N_8191,N_8084);
or U8659 (N_8659,N_8389,N_8358);
nand U8660 (N_8660,N_8197,N_8462);
and U8661 (N_8661,N_8030,N_8471);
nand U8662 (N_8662,N_8372,N_8225);
nor U8663 (N_8663,N_8078,N_8026);
and U8664 (N_8664,N_8118,N_8327);
or U8665 (N_8665,N_8439,N_8130);
xor U8666 (N_8666,N_8491,N_8226);
nand U8667 (N_8667,N_8034,N_8388);
xor U8668 (N_8668,N_8114,N_8356);
nor U8669 (N_8669,N_8236,N_8307);
xnor U8670 (N_8670,N_8487,N_8326);
nand U8671 (N_8671,N_8414,N_8404);
and U8672 (N_8672,N_8366,N_8399);
or U8673 (N_8673,N_8051,N_8117);
xor U8674 (N_8674,N_8477,N_8359);
and U8675 (N_8675,N_8072,N_8495);
or U8676 (N_8676,N_8328,N_8352);
or U8677 (N_8677,N_8371,N_8295);
and U8678 (N_8678,N_8365,N_8176);
nor U8679 (N_8679,N_8277,N_8021);
nand U8680 (N_8680,N_8086,N_8126);
and U8681 (N_8681,N_8171,N_8382);
nor U8682 (N_8682,N_8311,N_8385);
and U8683 (N_8683,N_8321,N_8142);
or U8684 (N_8684,N_8268,N_8337);
nor U8685 (N_8685,N_8170,N_8461);
and U8686 (N_8686,N_8175,N_8453);
nor U8687 (N_8687,N_8050,N_8068);
nand U8688 (N_8688,N_8203,N_8273);
and U8689 (N_8689,N_8150,N_8187);
and U8690 (N_8690,N_8189,N_8447);
and U8691 (N_8691,N_8158,N_8232);
nor U8692 (N_8692,N_8269,N_8233);
xnor U8693 (N_8693,N_8064,N_8323);
or U8694 (N_8694,N_8340,N_8033);
nor U8695 (N_8695,N_8380,N_8052);
xnor U8696 (N_8696,N_8460,N_8165);
xnor U8697 (N_8697,N_8131,N_8156);
and U8698 (N_8698,N_8103,N_8469);
and U8699 (N_8699,N_8441,N_8038);
or U8700 (N_8700,N_8308,N_8209);
nor U8701 (N_8701,N_8098,N_8003);
xor U8702 (N_8702,N_8309,N_8442);
xnor U8703 (N_8703,N_8045,N_8252);
and U8704 (N_8704,N_8406,N_8172);
and U8705 (N_8705,N_8250,N_8304);
nor U8706 (N_8706,N_8427,N_8200);
nand U8707 (N_8707,N_8434,N_8090);
xor U8708 (N_8708,N_8157,N_8394);
nand U8709 (N_8709,N_8361,N_8155);
nand U8710 (N_8710,N_8305,N_8259);
xor U8711 (N_8711,N_8132,N_8413);
nand U8712 (N_8712,N_8143,N_8369);
nor U8713 (N_8713,N_8105,N_8489);
nand U8714 (N_8714,N_8211,N_8266);
xnor U8715 (N_8715,N_8024,N_8271);
xor U8716 (N_8716,N_8048,N_8104);
xor U8717 (N_8717,N_8134,N_8218);
or U8718 (N_8718,N_8119,N_8056);
nand U8719 (N_8719,N_8036,N_8357);
nand U8720 (N_8720,N_8066,N_8071);
or U8721 (N_8721,N_8310,N_8044);
and U8722 (N_8722,N_8415,N_8207);
xor U8723 (N_8723,N_8073,N_8397);
nor U8724 (N_8724,N_8185,N_8001);
nor U8725 (N_8725,N_8065,N_8159);
xor U8726 (N_8726,N_8254,N_8137);
nand U8727 (N_8727,N_8179,N_8097);
and U8728 (N_8728,N_8246,N_8417);
or U8729 (N_8729,N_8163,N_8164);
nor U8730 (N_8730,N_8108,N_8497);
nand U8731 (N_8731,N_8094,N_8122);
xor U8732 (N_8732,N_8046,N_8418);
or U8733 (N_8733,N_8401,N_8395);
xnor U8734 (N_8734,N_8452,N_8198);
nor U8735 (N_8735,N_8346,N_8387);
xnor U8736 (N_8736,N_8330,N_8412);
nand U8737 (N_8737,N_8499,N_8100);
nor U8738 (N_8738,N_8319,N_8336);
or U8739 (N_8739,N_8008,N_8329);
nor U8740 (N_8740,N_8349,N_8299);
and U8741 (N_8741,N_8320,N_8161);
xnor U8742 (N_8742,N_8493,N_8128);
or U8743 (N_8743,N_8473,N_8373);
xnor U8744 (N_8744,N_8201,N_8432);
xor U8745 (N_8745,N_8058,N_8168);
or U8746 (N_8746,N_8004,N_8267);
and U8747 (N_8747,N_8041,N_8270);
or U8748 (N_8748,N_8007,N_8231);
nor U8749 (N_8749,N_8275,N_8438);
xor U8750 (N_8750,N_8365,N_8256);
nand U8751 (N_8751,N_8228,N_8274);
xnor U8752 (N_8752,N_8100,N_8408);
nand U8753 (N_8753,N_8317,N_8204);
xnor U8754 (N_8754,N_8120,N_8332);
nor U8755 (N_8755,N_8239,N_8080);
and U8756 (N_8756,N_8460,N_8440);
nor U8757 (N_8757,N_8463,N_8242);
or U8758 (N_8758,N_8323,N_8000);
nor U8759 (N_8759,N_8106,N_8153);
or U8760 (N_8760,N_8397,N_8242);
nor U8761 (N_8761,N_8318,N_8092);
or U8762 (N_8762,N_8186,N_8426);
nor U8763 (N_8763,N_8489,N_8267);
xnor U8764 (N_8764,N_8304,N_8266);
and U8765 (N_8765,N_8082,N_8415);
or U8766 (N_8766,N_8319,N_8220);
xnor U8767 (N_8767,N_8213,N_8105);
or U8768 (N_8768,N_8449,N_8371);
nor U8769 (N_8769,N_8074,N_8443);
xnor U8770 (N_8770,N_8226,N_8331);
nor U8771 (N_8771,N_8006,N_8116);
and U8772 (N_8772,N_8006,N_8133);
nor U8773 (N_8773,N_8156,N_8327);
or U8774 (N_8774,N_8184,N_8170);
or U8775 (N_8775,N_8292,N_8287);
nand U8776 (N_8776,N_8439,N_8020);
xor U8777 (N_8777,N_8245,N_8481);
nand U8778 (N_8778,N_8401,N_8176);
and U8779 (N_8779,N_8356,N_8495);
nor U8780 (N_8780,N_8034,N_8370);
and U8781 (N_8781,N_8052,N_8140);
or U8782 (N_8782,N_8039,N_8289);
nand U8783 (N_8783,N_8342,N_8441);
or U8784 (N_8784,N_8013,N_8390);
nand U8785 (N_8785,N_8420,N_8434);
nor U8786 (N_8786,N_8269,N_8461);
xnor U8787 (N_8787,N_8457,N_8433);
nor U8788 (N_8788,N_8028,N_8115);
nand U8789 (N_8789,N_8227,N_8392);
or U8790 (N_8790,N_8257,N_8388);
or U8791 (N_8791,N_8461,N_8029);
nor U8792 (N_8792,N_8175,N_8419);
and U8793 (N_8793,N_8353,N_8081);
or U8794 (N_8794,N_8252,N_8371);
or U8795 (N_8795,N_8497,N_8361);
or U8796 (N_8796,N_8114,N_8321);
xor U8797 (N_8797,N_8429,N_8069);
or U8798 (N_8798,N_8235,N_8045);
nand U8799 (N_8799,N_8458,N_8331);
or U8800 (N_8800,N_8094,N_8411);
nand U8801 (N_8801,N_8465,N_8156);
or U8802 (N_8802,N_8068,N_8010);
and U8803 (N_8803,N_8378,N_8365);
nor U8804 (N_8804,N_8093,N_8016);
and U8805 (N_8805,N_8301,N_8186);
nand U8806 (N_8806,N_8421,N_8401);
nor U8807 (N_8807,N_8307,N_8178);
nand U8808 (N_8808,N_8325,N_8289);
nor U8809 (N_8809,N_8459,N_8175);
nor U8810 (N_8810,N_8378,N_8054);
nor U8811 (N_8811,N_8474,N_8481);
nand U8812 (N_8812,N_8370,N_8109);
or U8813 (N_8813,N_8326,N_8192);
nor U8814 (N_8814,N_8064,N_8359);
or U8815 (N_8815,N_8098,N_8472);
nor U8816 (N_8816,N_8177,N_8262);
nor U8817 (N_8817,N_8403,N_8444);
nor U8818 (N_8818,N_8055,N_8468);
nor U8819 (N_8819,N_8495,N_8354);
and U8820 (N_8820,N_8278,N_8087);
nor U8821 (N_8821,N_8315,N_8451);
or U8822 (N_8822,N_8408,N_8183);
and U8823 (N_8823,N_8454,N_8306);
xor U8824 (N_8824,N_8421,N_8245);
xor U8825 (N_8825,N_8428,N_8091);
nor U8826 (N_8826,N_8019,N_8066);
nand U8827 (N_8827,N_8165,N_8120);
nor U8828 (N_8828,N_8143,N_8265);
nand U8829 (N_8829,N_8231,N_8334);
nor U8830 (N_8830,N_8208,N_8381);
nand U8831 (N_8831,N_8213,N_8443);
nand U8832 (N_8832,N_8136,N_8371);
or U8833 (N_8833,N_8372,N_8307);
or U8834 (N_8834,N_8098,N_8206);
xor U8835 (N_8835,N_8098,N_8028);
xor U8836 (N_8836,N_8403,N_8077);
and U8837 (N_8837,N_8277,N_8294);
or U8838 (N_8838,N_8457,N_8477);
nor U8839 (N_8839,N_8170,N_8041);
xnor U8840 (N_8840,N_8259,N_8058);
xnor U8841 (N_8841,N_8010,N_8463);
nor U8842 (N_8842,N_8001,N_8089);
or U8843 (N_8843,N_8115,N_8440);
or U8844 (N_8844,N_8406,N_8452);
nand U8845 (N_8845,N_8499,N_8440);
xnor U8846 (N_8846,N_8334,N_8148);
or U8847 (N_8847,N_8203,N_8450);
or U8848 (N_8848,N_8101,N_8428);
nor U8849 (N_8849,N_8478,N_8381);
xnor U8850 (N_8850,N_8018,N_8092);
xnor U8851 (N_8851,N_8200,N_8335);
xor U8852 (N_8852,N_8115,N_8083);
nand U8853 (N_8853,N_8239,N_8034);
nor U8854 (N_8854,N_8409,N_8053);
nor U8855 (N_8855,N_8145,N_8028);
or U8856 (N_8856,N_8438,N_8185);
and U8857 (N_8857,N_8479,N_8137);
and U8858 (N_8858,N_8122,N_8034);
xor U8859 (N_8859,N_8280,N_8158);
nor U8860 (N_8860,N_8274,N_8259);
or U8861 (N_8861,N_8381,N_8197);
and U8862 (N_8862,N_8253,N_8204);
xor U8863 (N_8863,N_8499,N_8126);
nor U8864 (N_8864,N_8325,N_8208);
nand U8865 (N_8865,N_8130,N_8179);
and U8866 (N_8866,N_8221,N_8145);
and U8867 (N_8867,N_8090,N_8330);
nor U8868 (N_8868,N_8293,N_8421);
or U8869 (N_8869,N_8419,N_8324);
nor U8870 (N_8870,N_8329,N_8086);
and U8871 (N_8871,N_8206,N_8221);
or U8872 (N_8872,N_8056,N_8037);
and U8873 (N_8873,N_8164,N_8137);
xnor U8874 (N_8874,N_8035,N_8133);
and U8875 (N_8875,N_8465,N_8049);
or U8876 (N_8876,N_8265,N_8179);
or U8877 (N_8877,N_8421,N_8220);
nor U8878 (N_8878,N_8495,N_8093);
nor U8879 (N_8879,N_8053,N_8283);
or U8880 (N_8880,N_8350,N_8034);
and U8881 (N_8881,N_8230,N_8008);
nand U8882 (N_8882,N_8374,N_8403);
xnor U8883 (N_8883,N_8142,N_8087);
nor U8884 (N_8884,N_8068,N_8231);
or U8885 (N_8885,N_8315,N_8264);
xor U8886 (N_8886,N_8433,N_8327);
xor U8887 (N_8887,N_8056,N_8060);
nor U8888 (N_8888,N_8345,N_8252);
nor U8889 (N_8889,N_8129,N_8339);
and U8890 (N_8890,N_8058,N_8183);
or U8891 (N_8891,N_8109,N_8326);
or U8892 (N_8892,N_8220,N_8022);
nor U8893 (N_8893,N_8047,N_8476);
and U8894 (N_8894,N_8057,N_8417);
xor U8895 (N_8895,N_8373,N_8494);
xnor U8896 (N_8896,N_8032,N_8101);
and U8897 (N_8897,N_8295,N_8465);
xor U8898 (N_8898,N_8121,N_8325);
and U8899 (N_8899,N_8143,N_8181);
nand U8900 (N_8900,N_8400,N_8453);
or U8901 (N_8901,N_8283,N_8087);
or U8902 (N_8902,N_8331,N_8375);
and U8903 (N_8903,N_8184,N_8210);
xnor U8904 (N_8904,N_8487,N_8149);
or U8905 (N_8905,N_8371,N_8058);
or U8906 (N_8906,N_8355,N_8459);
nand U8907 (N_8907,N_8496,N_8443);
nor U8908 (N_8908,N_8172,N_8350);
or U8909 (N_8909,N_8216,N_8279);
xnor U8910 (N_8910,N_8039,N_8498);
or U8911 (N_8911,N_8247,N_8308);
and U8912 (N_8912,N_8270,N_8014);
or U8913 (N_8913,N_8346,N_8239);
and U8914 (N_8914,N_8015,N_8354);
and U8915 (N_8915,N_8183,N_8351);
or U8916 (N_8916,N_8308,N_8168);
or U8917 (N_8917,N_8217,N_8028);
xnor U8918 (N_8918,N_8087,N_8377);
nand U8919 (N_8919,N_8132,N_8220);
xor U8920 (N_8920,N_8014,N_8291);
nor U8921 (N_8921,N_8255,N_8152);
xnor U8922 (N_8922,N_8164,N_8035);
nand U8923 (N_8923,N_8340,N_8071);
nand U8924 (N_8924,N_8367,N_8460);
xnor U8925 (N_8925,N_8111,N_8004);
xnor U8926 (N_8926,N_8463,N_8266);
xor U8927 (N_8927,N_8039,N_8329);
and U8928 (N_8928,N_8038,N_8054);
and U8929 (N_8929,N_8214,N_8478);
or U8930 (N_8930,N_8036,N_8463);
xor U8931 (N_8931,N_8276,N_8082);
nor U8932 (N_8932,N_8320,N_8378);
xnor U8933 (N_8933,N_8243,N_8052);
nor U8934 (N_8934,N_8240,N_8118);
or U8935 (N_8935,N_8285,N_8092);
nand U8936 (N_8936,N_8423,N_8072);
or U8937 (N_8937,N_8096,N_8110);
nor U8938 (N_8938,N_8452,N_8263);
nor U8939 (N_8939,N_8006,N_8299);
nor U8940 (N_8940,N_8465,N_8087);
nand U8941 (N_8941,N_8458,N_8182);
nand U8942 (N_8942,N_8378,N_8219);
nor U8943 (N_8943,N_8087,N_8170);
nand U8944 (N_8944,N_8383,N_8013);
nor U8945 (N_8945,N_8266,N_8323);
nand U8946 (N_8946,N_8215,N_8307);
and U8947 (N_8947,N_8337,N_8161);
nand U8948 (N_8948,N_8423,N_8457);
and U8949 (N_8949,N_8054,N_8383);
nand U8950 (N_8950,N_8177,N_8277);
nor U8951 (N_8951,N_8244,N_8105);
xnor U8952 (N_8952,N_8042,N_8153);
xnor U8953 (N_8953,N_8180,N_8108);
or U8954 (N_8954,N_8357,N_8291);
xor U8955 (N_8955,N_8162,N_8229);
nor U8956 (N_8956,N_8496,N_8453);
nand U8957 (N_8957,N_8144,N_8021);
nand U8958 (N_8958,N_8046,N_8209);
and U8959 (N_8959,N_8144,N_8337);
nand U8960 (N_8960,N_8231,N_8109);
or U8961 (N_8961,N_8084,N_8107);
nand U8962 (N_8962,N_8090,N_8246);
or U8963 (N_8963,N_8256,N_8426);
and U8964 (N_8964,N_8275,N_8440);
or U8965 (N_8965,N_8381,N_8031);
and U8966 (N_8966,N_8138,N_8054);
nor U8967 (N_8967,N_8048,N_8302);
and U8968 (N_8968,N_8198,N_8394);
nand U8969 (N_8969,N_8386,N_8463);
nor U8970 (N_8970,N_8238,N_8413);
or U8971 (N_8971,N_8057,N_8360);
and U8972 (N_8972,N_8335,N_8401);
or U8973 (N_8973,N_8492,N_8198);
and U8974 (N_8974,N_8050,N_8490);
or U8975 (N_8975,N_8280,N_8291);
xor U8976 (N_8976,N_8328,N_8244);
and U8977 (N_8977,N_8354,N_8410);
and U8978 (N_8978,N_8477,N_8399);
or U8979 (N_8979,N_8121,N_8313);
nand U8980 (N_8980,N_8358,N_8235);
nor U8981 (N_8981,N_8128,N_8319);
and U8982 (N_8982,N_8080,N_8155);
or U8983 (N_8983,N_8119,N_8363);
nand U8984 (N_8984,N_8200,N_8314);
nand U8985 (N_8985,N_8402,N_8134);
or U8986 (N_8986,N_8383,N_8274);
and U8987 (N_8987,N_8019,N_8190);
nor U8988 (N_8988,N_8126,N_8072);
nor U8989 (N_8989,N_8216,N_8348);
nor U8990 (N_8990,N_8417,N_8427);
xor U8991 (N_8991,N_8133,N_8451);
or U8992 (N_8992,N_8352,N_8070);
nand U8993 (N_8993,N_8079,N_8027);
or U8994 (N_8994,N_8142,N_8420);
xnor U8995 (N_8995,N_8445,N_8272);
nand U8996 (N_8996,N_8416,N_8395);
nor U8997 (N_8997,N_8122,N_8181);
and U8998 (N_8998,N_8012,N_8353);
and U8999 (N_8999,N_8319,N_8391);
and U9000 (N_9000,N_8885,N_8998);
or U9001 (N_9001,N_8595,N_8586);
and U9002 (N_9002,N_8684,N_8833);
nor U9003 (N_9003,N_8515,N_8717);
or U9004 (N_9004,N_8901,N_8800);
xnor U9005 (N_9005,N_8808,N_8894);
and U9006 (N_9006,N_8792,N_8990);
and U9007 (N_9007,N_8993,N_8771);
or U9008 (N_9008,N_8567,N_8528);
nand U9009 (N_9009,N_8588,N_8610);
nand U9010 (N_9010,N_8682,N_8531);
nand U9011 (N_9011,N_8738,N_8557);
xnor U9012 (N_9012,N_8571,N_8881);
xnor U9013 (N_9013,N_8855,N_8604);
nor U9014 (N_9014,N_8675,N_8561);
or U9015 (N_9015,N_8629,N_8893);
or U9016 (N_9016,N_8699,N_8826);
or U9017 (N_9017,N_8917,N_8525);
nand U9018 (N_9018,N_8667,N_8841);
nor U9019 (N_9019,N_8552,N_8678);
nor U9020 (N_9020,N_8820,N_8697);
nor U9021 (N_9021,N_8908,N_8563);
nor U9022 (N_9022,N_8829,N_8932);
nor U9023 (N_9023,N_8972,N_8980);
nor U9024 (N_9024,N_8910,N_8871);
and U9025 (N_9025,N_8711,N_8831);
nor U9026 (N_9026,N_8774,N_8956);
and U9027 (N_9027,N_8553,N_8679);
xnor U9028 (N_9028,N_8676,N_8746);
or U9029 (N_9029,N_8537,N_8749);
and U9030 (N_9030,N_8937,N_8695);
nand U9031 (N_9031,N_8704,N_8876);
and U9032 (N_9032,N_8880,N_8989);
nor U9033 (N_9033,N_8607,N_8896);
nand U9034 (N_9034,N_8756,N_8776);
and U9035 (N_9035,N_8565,N_8779);
xor U9036 (N_9036,N_8665,N_8784);
nor U9037 (N_9037,N_8971,N_8743);
and U9038 (N_9038,N_8560,N_8637);
xor U9039 (N_9039,N_8509,N_8873);
xnor U9040 (N_9040,N_8582,N_8838);
nor U9041 (N_9041,N_8631,N_8857);
or U9042 (N_9042,N_8986,N_8705);
and U9043 (N_9043,N_8544,N_8798);
nand U9044 (N_9044,N_8849,N_8801);
nor U9045 (N_9045,N_8897,N_8538);
nand U9046 (N_9046,N_8813,N_8994);
nand U9047 (N_9047,N_8527,N_8625);
or U9048 (N_9048,N_8739,N_8612);
nand U9049 (N_9049,N_8765,N_8673);
nor U9050 (N_9050,N_8715,N_8650);
nor U9051 (N_9051,N_8951,N_8783);
nand U9052 (N_9052,N_8955,N_8760);
xnor U9053 (N_9053,N_8891,N_8981);
nor U9054 (N_9054,N_8840,N_8593);
or U9055 (N_9055,N_8969,N_8599);
and U9056 (N_9056,N_8940,N_8983);
xor U9057 (N_9057,N_8888,N_8758);
and U9058 (N_9058,N_8514,N_8764);
nand U9059 (N_9059,N_8848,N_8968);
nor U9060 (N_9060,N_8733,N_8680);
nand U9061 (N_9061,N_8523,N_8519);
and U9062 (N_9062,N_8920,N_8741);
and U9063 (N_9063,N_8978,N_8953);
or U9064 (N_9064,N_8787,N_8858);
nand U9065 (N_9065,N_8874,N_8555);
or U9066 (N_9066,N_8830,N_8558);
nand U9067 (N_9067,N_8618,N_8533);
xnor U9068 (N_9068,N_8559,N_8921);
xnor U9069 (N_9069,N_8626,N_8662);
nor U9070 (N_9070,N_8622,N_8782);
or U9071 (N_9071,N_8817,N_8729);
and U9072 (N_9072,N_8750,N_8892);
nand U9073 (N_9073,N_8652,N_8959);
and U9074 (N_9074,N_8938,N_8814);
or U9075 (N_9075,N_8686,N_8661);
and U9076 (N_9076,N_8580,N_8827);
or U9077 (N_9077,N_8770,N_8534);
xor U9078 (N_9078,N_8668,N_8924);
nor U9079 (N_9079,N_8694,N_8708);
nor U9080 (N_9080,N_8658,N_8524);
and U9081 (N_9081,N_8608,N_8630);
nand U9082 (N_9082,N_8719,N_8616);
nor U9083 (N_9083,N_8825,N_8796);
nor U9084 (N_9084,N_8913,N_8882);
or U9085 (N_9085,N_8666,N_8898);
xor U9086 (N_9086,N_8850,N_8532);
nand U9087 (N_9087,N_8907,N_8832);
or U9088 (N_9088,N_8736,N_8816);
nor U9089 (N_9089,N_8887,N_8574);
nor U9090 (N_9090,N_8957,N_8721);
xor U9091 (N_9091,N_8962,N_8950);
xor U9092 (N_9092,N_8812,N_8999);
nor U9093 (N_9093,N_8778,N_8585);
nand U9094 (N_9094,N_8510,N_8573);
or U9095 (N_9095,N_8594,N_8797);
nand U9096 (N_9096,N_8728,N_8766);
nor U9097 (N_9097,N_8546,N_8867);
xor U9098 (N_9098,N_8720,N_8554);
and U9099 (N_9099,N_8562,N_8791);
xnor U9100 (N_9100,N_8692,N_8852);
nand U9101 (N_9101,N_8603,N_8579);
nor U9102 (N_9102,N_8621,N_8761);
xor U9103 (N_9103,N_8731,N_8570);
or U9104 (N_9104,N_8501,N_8638);
and U9105 (N_9105,N_8646,N_8768);
nand U9106 (N_9106,N_8949,N_8714);
and U9107 (N_9107,N_8641,N_8656);
nor U9108 (N_9108,N_8918,N_8550);
and U9109 (N_9109,N_8974,N_8987);
nor U9110 (N_9110,N_8506,N_8644);
nand U9111 (N_9111,N_8965,N_8824);
nor U9112 (N_9112,N_8961,N_8909);
xor U9113 (N_9113,N_8916,N_8627);
xor U9114 (N_9114,N_8681,N_8706);
or U9115 (N_9115,N_8500,N_8810);
and U9116 (N_9116,N_8605,N_8919);
or U9117 (N_9117,N_8591,N_8723);
or U9118 (N_9118,N_8520,N_8879);
xnor U9119 (N_9119,N_8996,N_8763);
and U9120 (N_9120,N_8698,N_8549);
nand U9121 (N_9121,N_8772,N_8773);
nand U9122 (N_9122,N_8602,N_8799);
xor U9123 (N_9123,N_8564,N_8914);
xnor U9124 (N_9124,N_8922,N_8903);
nand U9125 (N_9125,N_8870,N_8828);
xnor U9126 (N_9126,N_8865,N_8823);
or U9127 (N_9127,N_8842,N_8700);
xor U9128 (N_9128,N_8615,N_8929);
nand U9129 (N_9129,N_8657,N_8889);
or U9130 (N_9130,N_8516,N_8740);
xor U9131 (N_9131,N_8997,N_8687);
nor U9132 (N_9132,N_8732,N_8780);
nor U9133 (N_9133,N_8503,N_8596);
xnor U9134 (N_9134,N_8521,N_8718);
nor U9135 (N_9135,N_8716,N_8789);
xnor U9136 (N_9136,N_8781,N_8566);
nor U9137 (N_9137,N_8674,N_8624);
xor U9138 (N_9138,N_8755,N_8727);
nor U9139 (N_9139,N_8642,N_8734);
nand U9140 (N_9140,N_8691,N_8647);
nand U9141 (N_9141,N_8522,N_8786);
nor U9142 (N_9142,N_8899,N_8737);
nor U9143 (N_9143,N_8979,N_8707);
nand U9144 (N_9144,N_8725,N_8912);
and U9145 (N_9145,N_8539,N_8693);
nor U9146 (N_9146,N_8854,N_8685);
xnor U9147 (N_9147,N_8948,N_8722);
nand U9148 (N_9148,N_8540,N_8609);
nor U9149 (N_9149,N_8548,N_8655);
nor U9150 (N_9150,N_8536,N_8505);
and U9151 (N_9151,N_8902,N_8572);
or U9152 (N_9152,N_8995,N_8724);
xor U9153 (N_9153,N_8613,N_8973);
nor U9154 (N_9154,N_8590,N_8883);
xor U9155 (N_9155,N_8793,N_8877);
nand U9156 (N_9156,N_8688,N_8712);
nand U9157 (N_9157,N_8504,N_8811);
nand U9158 (N_9158,N_8703,N_8943);
xor U9159 (N_9159,N_8664,N_8795);
or U9160 (N_9160,N_8933,N_8958);
nor U9161 (N_9161,N_8587,N_8847);
or U9162 (N_9162,N_8767,N_8982);
nand U9163 (N_9163,N_8803,N_8518);
nor U9164 (N_9164,N_8752,N_8915);
and U9165 (N_9165,N_8878,N_8690);
and U9166 (N_9166,N_8569,N_8836);
nand U9167 (N_9167,N_8818,N_8512);
xor U9168 (N_9168,N_8805,N_8581);
and U9169 (N_9169,N_8611,N_8551);
and U9170 (N_9170,N_8985,N_8785);
or U9171 (N_9171,N_8906,N_8702);
xor U9172 (N_9172,N_8821,N_8640);
xor U9173 (N_9173,N_8804,N_8744);
or U9174 (N_9174,N_8508,N_8806);
nand U9175 (N_9175,N_8672,N_8872);
nand U9176 (N_9176,N_8670,N_8984);
nand U9177 (N_9177,N_8577,N_8934);
or U9178 (N_9178,N_8967,N_8936);
and U9179 (N_9179,N_8935,N_8730);
xor U9180 (N_9180,N_8890,N_8851);
xor U9181 (N_9181,N_8930,N_8619);
nor U9182 (N_9182,N_8923,N_8807);
xnor U9183 (N_9183,N_8643,N_8663);
or U9184 (N_9184,N_8925,N_8511);
nor U9185 (N_9185,N_8617,N_8946);
xnor U9186 (N_9186,N_8839,N_8545);
nand U9187 (N_9187,N_8726,N_8895);
nor U9188 (N_9188,N_8904,N_8844);
xnor U9189 (N_9189,N_8677,N_8775);
and U9190 (N_9190,N_8600,N_8794);
and U9191 (N_9191,N_8556,N_8926);
nor U9192 (N_9192,N_8835,N_8753);
nor U9193 (N_9193,N_8623,N_8576);
nand U9194 (N_9194,N_8660,N_8942);
nor U9195 (N_9195,N_8866,N_8952);
nor U9196 (N_9196,N_8671,N_8751);
or U9197 (N_9197,N_8975,N_8601);
nand U9198 (N_9198,N_8659,N_8701);
or U9199 (N_9199,N_8541,N_8529);
xor U9200 (N_9200,N_8762,N_8822);
and U9201 (N_9201,N_8769,N_8598);
nand U9202 (N_9202,N_8941,N_8815);
or U9203 (N_9203,N_8649,N_8592);
nand U9204 (N_9204,N_8911,N_8991);
nand U9205 (N_9205,N_8620,N_8502);
nor U9206 (N_9206,N_8614,N_8584);
and U9207 (N_9207,N_8589,N_8868);
and U9208 (N_9208,N_8683,N_8964);
nor U9209 (N_9209,N_8819,N_8834);
or U9210 (N_9210,N_8526,N_8954);
or U9211 (N_9211,N_8837,N_8861);
and U9212 (N_9212,N_8530,N_8859);
or U9213 (N_9213,N_8875,N_8869);
nor U9214 (N_9214,N_8742,N_8568);
and U9215 (N_9215,N_8754,N_8628);
and U9216 (N_9216,N_8633,N_8713);
xnor U9217 (N_9217,N_8966,N_8710);
nand U9218 (N_9218,N_8864,N_8517);
nand U9219 (N_9219,N_8689,N_8944);
nor U9220 (N_9220,N_8960,N_8759);
or U9221 (N_9221,N_8853,N_8777);
nor U9222 (N_9222,N_8970,N_8977);
xor U9223 (N_9223,N_8632,N_8735);
or U9224 (N_9224,N_8634,N_8597);
xor U9225 (N_9225,N_8575,N_8535);
xnor U9226 (N_9226,N_8843,N_8884);
or U9227 (N_9227,N_8583,N_8860);
or U9228 (N_9228,N_8809,N_8748);
xor U9229 (N_9229,N_8976,N_8745);
or U9230 (N_9230,N_8757,N_8947);
xor U9231 (N_9231,N_8963,N_8863);
or U9232 (N_9232,N_8606,N_8578);
nand U9233 (N_9233,N_8645,N_8845);
and U9234 (N_9234,N_8856,N_8507);
and U9235 (N_9235,N_8542,N_8928);
or U9236 (N_9236,N_8696,N_8988);
and U9237 (N_9237,N_8648,N_8513);
nor U9238 (N_9238,N_8905,N_8992);
nor U9239 (N_9239,N_8939,N_8747);
and U9240 (N_9240,N_8653,N_8802);
and U9241 (N_9241,N_8927,N_8945);
and U9242 (N_9242,N_8900,N_8931);
or U9243 (N_9243,N_8790,N_8636);
nor U9244 (N_9244,N_8654,N_8635);
xor U9245 (N_9245,N_8709,N_8788);
xor U9246 (N_9246,N_8846,N_8639);
and U9247 (N_9247,N_8886,N_8547);
xor U9248 (N_9248,N_8669,N_8651);
or U9249 (N_9249,N_8862,N_8543);
xnor U9250 (N_9250,N_8651,N_8845);
or U9251 (N_9251,N_8882,N_8853);
and U9252 (N_9252,N_8609,N_8804);
nand U9253 (N_9253,N_8644,N_8807);
or U9254 (N_9254,N_8825,N_8769);
or U9255 (N_9255,N_8511,N_8860);
and U9256 (N_9256,N_8804,N_8835);
nand U9257 (N_9257,N_8626,N_8711);
nand U9258 (N_9258,N_8741,N_8905);
or U9259 (N_9259,N_8527,N_8578);
and U9260 (N_9260,N_8839,N_8689);
or U9261 (N_9261,N_8612,N_8720);
nand U9262 (N_9262,N_8693,N_8888);
xnor U9263 (N_9263,N_8876,N_8850);
xor U9264 (N_9264,N_8652,N_8827);
and U9265 (N_9265,N_8828,N_8626);
nor U9266 (N_9266,N_8967,N_8969);
xnor U9267 (N_9267,N_8869,N_8708);
xnor U9268 (N_9268,N_8974,N_8928);
nand U9269 (N_9269,N_8718,N_8837);
nor U9270 (N_9270,N_8987,N_8837);
xnor U9271 (N_9271,N_8932,N_8605);
nand U9272 (N_9272,N_8966,N_8584);
and U9273 (N_9273,N_8846,N_8823);
nand U9274 (N_9274,N_8956,N_8873);
xnor U9275 (N_9275,N_8589,N_8804);
nor U9276 (N_9276,N_8644,N_8751);
or U9277 (N_9277,N_8913,N_8821);
xor U9278 (N_9278,N_8798,N_8929);
nand U9279 (N_9279,N_8753,N_8783);
and U9280 (N_9280,N_8728,N_8909);
nand U9281 (N_9281,N_8919,N_8984);
nand U9282 (N_9282,N_8864,N_8998);
nor U9283 (N_9283,N_8505,N_8769);
nor U9284 (N_9284,N_8921,N_8632);
xor U9285 (N_9285,N_8613,N_8692);
nor U9286 (N_9286,N_8687,N_8791);
xor U9287 (N_9287,N_8798,N_8900);
nand U9288 (N_9288,N_8872,N_8948);
xor U9289 (N_9289,N_8615,N_8588);
or U9290 (N_9290,N_8881,N_8931);
xor U9291 (N_9291,N_8530,N_8734);
or U9292 (N_9292,N_8854,N_8937);
and U9293 (N_9293,N_8707,N_8983);
and U9294 (N_9294,N_8728,N_8887);
nor U9295 (N_9295,N_8642,N_8982);
xnor U9296 (N_9296,N_8856,N_8972);
nor U9297 (N_9297,N_8786,N_8941);
or U9298 (N_9298,N_8997,N_8634);
or U9299 (N_9299,N_8817,N_8611);
nand U9300 (N_9300,N_8633,N_8670);
nand U9301 (N_9301,N_8912,N_8792);
nor U9302 (N_9302,N_8581,N_8855);
nor U9303 (N_9303,N_8656,N_8539);
nor U9304 (N_9304,N_8835,N_8690);
and U9305 (N_9305,N_8747,N_8737);
nor U9306 (N_9306,N_8884,N_8950);
nand U9307 (N_9307,N_8885,N_8891);
and U9308 (N_9308,N_8994,N_8765);
nor U9309 (N_9309,N_8864,N_8829);
and U9310 (N_9310,N_8667,N_8704);
and U9311 (N_9311,N_8646,N_8755);
nor U9312 (N_9312,N_8753,N_8897);
nor U9313 (N_9313,N_8608,N_8564);
or U9314 (N_9314,N_8701,N_8948);
xnor U9315 (N_9315,N_8636,N_8925);
and U9316 (N_9316,N_8503,N_8727);
and U9317 (N_9317,N_8995,N_8844);
nor U9318 (N_9318,N_8939,N_8925);
and U9319 (N_9319,N_8599,N_8602);
xnor U9320 (N_9320,N_8527,N_8941);
nand U9321 (N_9321,N_8788,N_8653);
or U9322 (N_9322,N_8672,N_8630);
xnor U9323 (N_9323,N_8884,N_8658);
nand U9324 (N_9324,N_8602,N_8660);
nor U9325 (N_9325,N_8782,N_8637);
and U9326 (N_9326,N_8821,N_8963);
nor U9327 (N_9327,N_8504,N_8764);
and U9328 (N_9328,N_8753,N_8703);
or U9329 (N_9329,N_8566,N_8674);
and U9330 (N_9330,N_8652,N_8728);
xor U9331 (N_9331,N_8523,N_8569);
nand U9332 (N_9332,N_8975,N_8588);
nand U9333 (N_9333,N_8574,N_8608);
xor U9334 (N_9334,N_8811,N_8642);
nand U9335 (N_9335,N_8589,N_8980);
or U9336 (N_9336,N_8882,N_8827);
xor U9337 (N_9337,N_8681,N_8599);
xnor U9338 (N_9338,N_8532,N_8540);
and U9339 (N_9339,N_8948,N_8559);
or U9340 (N_9340,N_8629,N_8604);
nor U9341 (N_9341,N_8643,N_8670);
nor U9342 (N_9342,N_8696,N_8761);
or U9343 (N_9343,N_8852,N_8581);
nand U9344 (N_9344,N_8974,N_8668);
nand U9345 (N_9345,N_8532,N_8687);
nand U9346 (N_9346,N_8852,N_8661);
nor U9347 (N_9347,N_8693,N_8893);
and U9348 (N_9348,N_8822,N_8957);
or U9349 (N_9349,N_8957,N_8537);
nand U9350 (N_9350,N_8631,N_8981);
nand U9351 (N_9351,N_8913,N_8530);
nor U9352 (N_9352,N_8733,N_8763);
nor U9353 (N_9353,N_8548,N_8695);
and U9354 (N_9354,N_8784,N_8811);
and U9355 (N_9355,N_8821,N_8920);
xor U9356 (N_9356,N_8821,N_8709);
and U9357 (N_9357,N_8820,N_8559);
xnor U9358 (N_9358,N_8826,N_8863);
nand U9359 (N_9359,N_8617,N_8818);
xnor U9360 (N_9360,N_8637,N_8544);
or U9361 (N_9361,N_8785,N_8633);
and U9362 (N_9362,N_8924,N_8951);
or U9363 (N_9363,N_8525,N_8680);
xor U9364 (N_9364,N_8562,N_8660);
xor U9365 (N_9365,N_8612,N_8804);
xor U9366 (N_9366,N_8721,N_8822);
or U9367 (N_9367,N_8945,N_8589);
or U9368 (N_9368,N_8670,N_8535);
nand U9369 (N_9369,N_8617,N_8656);
and U9370 (N_9370,N_8870,N_8664);
nor U9371 (N_9371,N_8973,N_8644);
xor U9372 (N_9372,N_8530,N_8523);
and U9373 (N_9373,N_8576,N_8524);
and U9374 (N_9374,N_8707,N_8999);
nor U9375 (N_9375,N_8979,N_8616);
nor U9376 (N_9376,N_8929,N_8621);
and U9377 (N_9377,N_8554,N_8674);
nand U9378 (N_9378,N_8687,N_8771);
xnor U9379 (N_9379,N_8544,N_8532);
and U9380 (N_9380,N_8897,N_8532);
or U9381 (N_9381,N_8795,N_8515);
and U9382 (N_9382,N_8850,N_8527);
and U9383 (N_9383,N_8938,N_8676);
xnor U9384 (N_9384,N_8768,N_8703);
xor U9385 (N_9385,N_8538,N_8561);
or U9386 (N_9386,N_8942,N_8676);
xor U9387 (N_9387,N_8770,N_8765);
nand U9388 (N_9388,N_8980,N_8995);
xnor U9389 (N_9389,N_8755,N_8639);
xor U9390 (N_9390,N_8641,N_8735);
nor U9391 (N_9391,N_8670,N_8530);
or U9392 (N_9392,N_8843,N_8805);
or U9393 (N_9393,N_8897,N_8979);
nand U9394 (N_9394,N_8739,N_8587);
nor U9395 (N_9395,N_8622,N_8501);
nand U9396 (N_9396,N_8867,N_8687);
or U9397 (N_9397,N_8687,N_8615);
nand U9398 (N_9398,N_8774,N_8701);
xor U9399 (N_9399,N_8836,N_8894);
nand U9400 (N_9400,N_8549,N_8796);
and U9401 (N_9401,N_8608,N_8968);
or U9402 (N_9402,N_8552,N_8715);
xnor U9403 (N_9403,N_8860,N_8870);
nand U9404 (N_9404,N_8999,N_8577);
or U9405 (N_9405,N_8786,N_8727);
and U9406 (N_9406,N_8580,N_8618);
nor U9407 (N_9407,N_8840,N_8773);
or U9408 (N_9408,N_8559,N_8696);
and U9409 (N_9409,N_8964,N_8653);
xnor U9410 (N_9410,N_8620,N_8752);
and U9411 (N_9411,N_8892,N_8751);
and U9412 (N_9412,N_8796,N_8643);
nand U9413 (N_9413,N_8657,N_8867);
or U9414 (N_9414,N_8632,N_8765);
or U9415 (N_9415,N_8637,N_8839);
or U9416 (N_9416,N_8737,N_8785);
xor U9417 (N_9417,N_8780,N_8518);
nor U9418 (N_9418,N_8668,N_8915);
nand U9419 (N_9419,N_8543,N_8541);
nand U9420 (N_9420,N_8984,N_8715);
xor U9421 (N_9421,N_8725,N_8917);
nand U9422 (N_9422,N_8863,N_8717);
xnor U9423 (N_9423,N_8804,N_8885);
or U9424 (N_9424,N_8898,N_8966);
and U9425 (N_9425,N_8540,N_8779);
xnor U9426 (N_9426,N_8609,N_8524);
nor U9427 (N_9427,N_8804,N_8696);
or U9428 (N_9428,N_8583,N_8597);
and U9429 (N_9429,N_8561,N_8772);
and U9430 (N_9430,N_8520,N_8758);
xnor U9431 (N_9431,N_8524,N_8558);
nor U9432 (N_9432,N_8720,N_8645);
nand U9433 (N_9433,N_8588,N_8904);
nand U9434 (N_9434,N_8804,N_8747);
xnor U9435 (N_9435,N_8898,N_8883);
nand U9436 (N_9436,N_8838,N_8553);
nand U9437 (N_9437,N_8533,N_8582);
and U9438 (N_9438,N_8802,N_8751);
and U9439 (N_9439,N_8623,N_8675);
nor U9440 (N_9440,N_8672,N_8878);
and U9441 (N_9441,N_8925,N_8725);
or U9442 (N_9442,N_8559,N_8623);
nand U9443 (N_9443,N_8554,N_8558);
and U9444 (N_9444,N_8575,N_8572);
nor U9445 (N_9445,N_8511,N_8777);
and U9446 (N_9446,N_8812,N_8551);
or U9447 (N_9447,N_8769,N_8815);
or U9448 (N_9448,N_8598,N_8533);
xor U9449 (N_9449,N_8849,N_8745);
xor U9450 (N_9450,N_8590,N_8940);
xnor U9451 (N_9451,N_8875,N_8685);
nor U9452 (N_9452,N_8520,N_8686);
and U9453 (N_9453,N_8830,N_8808);
xnor U9454 (N_9454,N_8652,N_8717);
or U9455 (N_9455,N_8833,N_8696);
and U9456 (N_9456,N_8678,N_8760);
or U9457 (N_9457,N_8550,N_8926);
nand U9458 (N_9458,N_8607,N_8869);
nand U9459 (N_9459,N_8700,N_8627);
xor U9460 (N_9460,N_8730,N_8994);
nand U9461 (N_9461,N_8615,N_8949);
nor U9462 (N_9462,N_8953,N_8951);
nand U9463 (N_9463,N_8792,N_8504);
and U9464 (N_9464,N_8994,N_8634);
or U9465 (N_9465,N_8729,N_8944);
nor U9466 (N_9466,N_8890,N_8964);
xnor U9467 (N_9467,N_8950,N_8519);
nor U9468 (N_9468,N_8773,N_8713);
nand U9469 (N_9469,N_8886,N_8564);
and U9470 (N_9470,N_8632,N_8904);
and U9471 (N_9471,N_8842,N_8844);
and U9472 (N_9472,N_8500,N_8766);
or U9473 (N_9473,N_8637,N_8989);
and U9474 (N_9474,N_8622,N_8644);
nand U9475 (N_9475,N_8821,N_8931);
nor U9476 (N_9476,N_8514,N_8628);
and U9477 (N_9477,N_8684,N_8779);
or U9478 (N_9478,N_8764,N_8602);
and U9479 (N_9479,N_8615,N_8651);
xnor U9480 (N_9480,N_8647,N_8630);
and U9481 (N_9481,N_8848,N_8761);
nor U9482 (N_9482,N_8978,N_8889);
and U9483 (N_9483,N_8995,N_8673);
or U9484 (N_9484,N_8954,N_8628);
xor U9485 (N_9485,N_8676,N_8629);
nor U9486 (N_9486,N_8715,N_8604);
and U9487 (N_9487,N_8548,N_8723);
or U9488 (N_9488,N_8965,N_8789);
or U9489 (N_9489,N_8785,N_8830);
and U9490 (N_9490,N_8604,N_8996);
nor U9491 (N_9491,N_8513,N_8766);
nor U9492 (N_9492,N_8870,N_8963);
xor U9493 (N_9493,N_8886,N_8740);
and U9494 (N_9494,N_8833,N_8736);
nor U9495 (N_9495,N_8706,N_8957);
or U9496 (N_9496,N_8794,N_8741);
or U9497 (N_9497,N_8735,N_8649);
nand U9498 (N_9498,N_8860,N_8737);
nor U9499 (N_9499,N_8894,N_8677);
xor U9500 (N_9500,N_9464,N_9232);
or U9501 (N_9501,N_9276,N_9009);
xnor U9502 (N_9502,N_9081,N_9296);
and U9503 (N_9503,N_9165,N_9173);
nand U9504 (N_9504,N_9431,N_9086);
xor U9505 (N_9505,N_9472,N_9361);
nand U9506 (N_9506,N_9167,N_9060);
nor U9507 (N_9507,N_9380,N_9351);
nor U9508 (N_9508,N_9368,N_9181);
or U9509 (N_9509,N_9451,N_9034);
nor U9510 (N_9510,N_9303,N_9427);
nor U9511 (N_9511,N_9308,N_9184);
or U9512 (N_9512,N_9172,N_9033);
xor U9513 (N_9513,N_9058,N_9051);
or U9514 (N_9514,N_9062,N_9254);
xnor U9515 (N_9515,N_9367,N_9126);
or U9516 (N_9516,N_9100,N_9493);
nor U9517 (N_9517,N_9372,N_9204);
xnor U9518 (N_9518,N_9483,N_9435);
or U9519 (N_9519,N_9484,N_9320);
xnor U9520 (N_9520,N_9155,N_9392);
xor U9521 (N_9521,N_9359,N_9331);
nand U9522 (N_9522,N_9156,N_9273);
and U9523 (N_9523,N_9246,N_9010);
or U9524 (N_9524,N_9417,N_9411);
nor U9525 (N_9525,N_9142,N_9406);
nor U9526 (N_9526,N_9404,N_9026);
nand U9527 (N_9527,N_9257,N_9337);
nor U9528 (N_9528,N_9133,N_9301);
or U9529 (N_9529,N_9350,N_9007);
nor U9530 (N_9530,N_9251,N_9466);
or U9531 (N_9531,N_9347,N_9469);
or U9532 (N_9532,N_9087,N_9252);
nor U9533 (N_9533,N_9475,N_9462);
nand U9534 (N_9534,N_9290,N_9478);
xor U9535 (N_9535,N_9023,N_9274);
nor U9536 (N_9536,N_9281,N_9410);
nor U9537 (N_9537,N_9069,N_9446);
nand U9538 (N_9538,N_9066,N_9068);
nor U9539 (N_9539,N_9434,N_9024);
xor U9540 (N_9540,N_9113,N_9208);
and U9541 (N_9541,N_9219,N_9352);
or U9542 (N_9542,N_9234,N_9382);
nor U9543 (N_9543,N_9111,N_9452);
nor U9544 (N_9544,N_9095,N_9283);
and U9545 (N_9545,N_9178,N_9148);
xor U9546 (N_9546,N_9362,N_9166);
xnor U9547 (N_9547,N_9210,N_9025);
nand U9548 (N_9548,N_9363,N_9358);
xnor U9549 (N_9549,N_9237,N_9398);
xor U9550 (N_9550,N_9371,N_9098);
nand U9551 (N_9551,N_9271,N_9152);
and U9552 (N_9552,N_9220,N_9312);
or U9553 (N_9553,N_9415,N_9272);
nand U9554 (N_9554,N_9035,N_9116);
nand U9555 (N_9555,N_9141,N_9473);
or U9556 (N_9556,N_9340,N_9366);
nand U9557 (N_9557,N_9265,N_9109);
nand U9558 (N_9558,N_9316,N_9117);
nand U9559 (N_9559,N_9393,N_9425);
and U9560 (N_9560,N_9499,N_9082);
and U9561 (N_9561,N_9479,N_9342);
or U9562 (N_9562,N_9319,N_9092);
or U9563 (N_9563,N_9416,N_9032);
and U9564 (N_9564,N_9375,N_9294);
xnor U9565 (N_9565,N_9130,N_9430);
nor U9566 (N_9566,N_9145,N_9465);
nand U9567 (N_9567,N_9075,N_9106);
nor U9568 (N_9568,N_9201,N_9162);
nor U9569 (N_9569,N_9150,N_9074);
nor U9570 (N_9570,N_9004,N_9450);
xor U9571 (N_9571,N_9467,N_9238);
nand U9572 (N_9572,N_9346,N_9055);
nand U9573 (N_9573,N_9151,N_9215);
nand U9574 (N_9574,N_9453,N_9225);
nor U9575 (N_9575,N_9063,N_9182);
xor U9576 (N_9576,N_9481,N_9037);
and U9577 (N_9577,N_9241,N_9029);
and U9578 (N_9578,N_9212,N_9408);
xor U9579 (N_9579,N_9344,N_9268);
nand U9580 (N_9580,N_9080,N_9441);
xnor U9581 (N_9581,N_9053,N_9138);
nor U9582 (N_9582,N_9048,N_9176);
nor U9583 (N_9583,N_9461,N_9269);
nand U9584 (N_9584,N_9123,N_9059);
or U9585 (N_9585,N_9031,N_9146);
nor U9586 (N_9586,N_9468,N_9270);
and U9587 (N_9587,N_9258,N_9044);
nand U9588 (N_9588,N_9209,N_9492);
and U9589 (N_9589,N_9012,N_9399);
xnor U9590 (N_9590,N_9437,N_9459);
and U9591 (N_9591,N_9047,N_9327);
nand U9592 (N_9592,N_9125,N_9355);
or U9593 (N_9593,N_9057,N_9214);
nor U9594 (N_9594,N_9174,N_9199);
and U9595 (N_9595,N_9083,N_9288);
nand U9596 (N_9596,N_9292,N_9315);
or U9597 (N_9597,N_9096,N_9188);
nand U9598 (N_9598,N_9022,N_9402);
and U9599 (N_9599,N_9448,N_9042);
or U9600 (N_9600,N_9357,N_9134);
nand U9601 (N_9601,N_9256,N_9231);
xnor U9602 (N_9602,N_9305,N_9159);
and U9603 (N_9603,N_9262,N_9020);
xnor U9604 (N_9604,N_9287,N_9282);
and U9605 (N_9605,N_9221,N_9127);
and U9606 (N_9606,N_9115,N_9110);
nor U9607 (N_9607,N_9299,N_9235);
or U9608 (N_9608,N_9414,N_9045);
xnor U9609 (N_9609,N_9280,N_9300);
xnor U9610 (N_9610,N_9005,N_9236);
xnor U9611 (N_9611,N_9409,N_9379);
nor U9612 (N_9612,N_9496,N_9318);
and U9613 (N_9613,N_9071,N_9217);
xnor U9614 (N_9614,N_9384,N_9284);
xnor U9615 (N_9615,N_9264,N_9003);
and U9616 (N_9616,N_9480,N_9482);
xor U9617 (N_9617,N_9444,N_9070);
and U9618 (N_9618,N_9144,N_9193);
xor U9619 (N_9619,N_9438,N_9291);
nand U9620 (N_9620,N_9476,N_9163);
xnor U9621 (N_9621,N_9385,N_9027);
or U9622 (N_9622,N_9107,N_9226);
xnor U9623 (N_9623,N_9240,N_9149);
nor U9624 (N_9624,N_9397,N_9378);
nor U9625 (N_9625,N_9317,N_9248);
nor U9626 (N_9626,N_9157,N_9454);
xnor U9627 (N_9627,N_9136,N_9353);
or U9628 (N_9628,N_9383,N_9046);
or U9629 (N_9629,N_9495,N_9354);
or U9630 (N_9630,N_9065,N_9374);
xor U9631 (N_9631,N_9213,N_9021);
nand U9632 (N_9632,N_9423,N_9341);
or U9633 (N_9633,N_9131,N_9094);
or U9634 (N_9634,N_9436,N_9485);
xnor U9635 (N_9635,N_9442,N_9191);
nand U9636 (N_9636,N_9449,N_9293);
xnor U9637 (N_9637,N_9322,N_9477);
and U9638 (N_9638,N_9064,N_9386);
and U9639 (N_9639,N_9323,N_9028);
or U9640 (N_9640,N_9348,N_9297);
nand U9641 (N_9641,N_9286,N_9013);
or U9642 (N_9642,N_9329,N_9334);
or U9643 (N_9643,N_9049,N_9185);
nor U9644 (N_9644,N_9019,N_9298);
and U9645 (N_9645,N_9067,N_9158);
and U9646 (N_9646,N_9389,N_9443);
xnor U9647 (N_9647,N_9360,N_9186);
or U9648 (N_9648,N_9494,N_9242);
nor U9649 (N_9649,N_9326,N_9207);
xnor U9650 (N_9650,N_9008,N_9061);
and U9651 (N_9651,N_9405,N_9486);
nor U9652 (N_9652,N_9222,N_9330);
and U9653 (N_9653,N_9135,N_9306);
nor U9654 (N_9654,N_9164,N_9439);
xor U9655 (N_9655,N_9089,N_9054);
or U9656 (N_9656,N_9377,N_9364);
xor U9657 (N_9657,N_9309,N_9119);
or U9658 (N_9658,N_9088,N_9120);
nand U9659 (N_9659,N_9161,N_9000);
nand U9660 (N_9660,N_9030,N_9394);
nand U9661 (N_9661,N_9369,N_9233);
nor U9662 (N_9662,N_9097,N_9421);
and U9663 (N_9663,N_9140,N_9224);
xnor U9664 (N_9664,N_9103,N_9079);
xor U9665 (N_9665,N_9339,N_9203);
or U9666 (N_9666,N_9139,N_9200);
and U9667 (N_9667,N_9244,N_9267);
xnor U9668 (N_9668,N_9104,N_9147);
xnor U9669 (N_9669,N_9228,N_9419);
or U9670 (N_9670,N_9324,N_9036);
and U9671 (N_9671,N_9403,N_9078);
xor U9672 (N_9672,N_9381,N_9422);
nor U9673 (N_9673,N_9400,N_9278);
or U9674 (N_9674,N_9018,N_9457);
nand U9675 (N_9675,N_9407,N_9420);
nor U9676 (N_9676,N_9460,N_9170);
xnor U9677 (N_9677,N_9491,N_9335);
nand U9678 (N_9678,N_9310,N_9455);
xnor U9679 (N_9679,N_9277,N_9202);
nor U9680 (N_9680,N_9255,N_9040);
nor U9681 (N_9681,N_9311,N_9043);
nor U9682 (N_9682,N_9333,N_9218);
nand U9683 (N_9683,N_9194,N_9445);
and U9684 (N_9684,N_9216,N_9413);
nor U9685 (N_9685,N_9121,N_9307);
xnor U9686 (N_9686,N_9249,N_9471);
nor U9687 (N_9687,N_9247,N_9160);
nor U9688 (N_9688,N_9412,N_9429);
nor U9689 (N_9689,N_9015,N_9002);
xor U9690 (N_9690,N_9370,N_9050);
nor U9691 (N_9691,N_9108,N_9304);
or U9692 (N_9692,N_9401,N_9498);
nor U9693 (N_9693,N_9243,N_9175);
and U9694 (N_9694,N_9205,N_9314);
xnor U9695 (N_9695,N_9376,N_9321);
or U9696 (N_9696,N_9017,N_9014);
nand U9697 (N_9697,N_9090,N_9391);
or U9698 (N_9698,N_9390,N_9489);
or U9699 (N_9699,N_9470,N_9189);
nand U9700 (N_9700,N_9313,N_9458);
nor U9701 (N_9701,N_9105,N_9190);
or U9702 (N_9702,N_9227,N_9154);
nand U9703 (N_9703,N_9076,N_9102);
nor U9704 (N_9704,N_9196,N_9072);
or U9705 (N_9705,N_9129,N_9356);
and U9706 (N_9706,N_9245,N_9132);
nand U9707 (N_9707,N_9016,N_9295);
or U9708 (N_9708,N_9038,N_9349);
or U9709 (N_9709,N_9259,N_9285);
xnor U9710 (N_9710,N_9039,N_9230);
or U9711 (N_9711,N_9183,N_9260);
nor U9712 (N_9712,N_9153,N_9328);
nor U9713 (N_9713,N_9488,N_9085);
xor U9714 (N_9714,N_9056,N_9041);
or U9715 (N_9715,N_9474,N_9229);
or U9716 (N_9716,N_9396,N_9497);
or U9717 (N_9717,N_9192,N_9179);
or U9718 (N_9718,N_9338,N_9387);
or U9719 (N_9719,N_9101,N_9302);
or U9720 (N_9720,N_9325,N_9118);
xnor U9721 (N_9721,N_9093,N_9052);
nor U9722 (N_9722,N_9084,N_9266);
xor U9723 (N_9723,N_9487,N_9490);
and U9724 (N_9724,N_9279,N_9128);
or U9725 (N_9725,N_9169,N_9345);
or U9726 (N_9726,N_9187,N_9011);
nor U9727 (N_9727,N_9426,N_9332);
nand U9728 (N_9728,N_9418,N_9261);
and U9729 (N_9729,N_9177,N_9171);
and U9730 (N_9730,N_9343,N_9073);
nand U9731 (N_9731,N_9137,N_9001);
and U9732 (N_9732,N_9206,N_9250);
and U9733 (N_9733,N_9424,N_9432);
nor U9734 (N_9734,N_9223,N_9253);
and U9735 (N_9735,N_9428,N_9143);
and U9736 (N_9736,N_9263,N_9112);
and U9737 (N_9737,N_9239,N_9168);
and U9738 (N_9738,N_9124,N_9195);
xor U9739 (N_9739,N_9091,N_9456);
nor U9740 (N_9740,N_9388,N_9275);
and U9741 (N_9741,N_9122,N_9211);
and U9742 (N_9742,N_9365,N_9077);
nand U9743 (N_9743,N_9114,N_9006);
xor U9744 (N_9744,N_9336,N_9463);
nand U9745 (N_9745,N_9395,N_9447);
nor U9746 (N_9746,N_9289,N_9198);
nand U9747 (N_9747,N_9180,N_9433);
and U9748 (N_9748,N_9197,N_9440);
or U9749 (N_9749,N_9373,N_9099);
and U9750 (N_9750,N_9162,N_9226);
or U9751 (N_9751,N_9207,N_9482);
and U9752 (N_9752,N_9463,N_9158);
and U9753 (N_9753,N_9063,N_9084);
and U9754 (N_9754,N_9147,N_9436);
xnor U9755 (N_9755,N_9271,N_9138);
nand U9756 (N_9756,N_9056,N_9389);
nand U9757 (N_9757,N_9020,N_9067);
and U9758 (N_9758,N_9389,N_9020);
or U9759 (N_9759,N_9465,N_9278);
xor U9760 (N_9760,N_9182,N_9421);
and U9761 (N_9761,N_9322,N_9393);
or U9762 (N_9762,N_9481,N_9424);
nor U9763 (N_9763,N_9066,N_9498);
nand U9764 (N_9764,N_9263,N_9198);
nor U9765 (N_9765,N_9176,N_9349);
and U9766 (N_9766,N_9106,N_9136);
nand U9767 (N_9767,N_9135,N_9208);
nand U9768 (N_9768,N_9236,N_9207);
nor U9769 (N_9769,N_9467,N_9340);
and U9770 (N_9770,N_9272,N_9165);
and U9771 (N_9771,N_9260,N_9139);
nand U9772 (N_9772,N_9429,N_9328);
xor U9773 (N_9773,N_9170,N_9367);
xnor U9774 (N_9774,N_9042,N_9249);
nand U9775 (N_9775,N_9219,N_9480);
or U9776 (N_9776,N_9154,N_9490);
nand U9777 (N_9777,N_9281,N_9143);
and U9778 (N_9778,N_9130,N_9434);
or U9779 (N_9779,N_9137,N_9124);
or U9780 (N_9780,N_9237,N_9153);
nand U9781 (N_9781,N_9291,N_9095);
nand U9782 (N_9782,N_9208,N_9058);
nor U9783 (N_9783,N_9340,N_9343);
and U9784 (N_9784,N_9229,N_9181);
nand U9785 (N_9785,N_9014,N_9259);
xor U9786 (N_9786,N_9324,N_9144);
nor U9787 (N_9787,N_9499,N_9052);
nor U9788 (N_9788,N_9333,N_9457);
xor U9789 (N_9789,N_9330,N_9390);
nor U9790 (N_9790,N_9114,N_9001);
nand U9791 (N_9791,N_9073,N_9203);
nor U9792 (N_9792,N_9016,N_9276);
and U9793 (N_9793,N_9410,N_9441);
and U9794 (N_9794,N_9412,N_9249);
or U9795 (N_9795,N_9095,N_9155);
nand U9796 (N_9796,N_9167,N_9341);
nand U9797 (N_9797,N_9141,N_9070);
and U9798 (N_9798,N_9147,N_9017);
and U9799 (N_9799,N_9009,N_9242);
nor U9800 (N_9800,N_9063,N_9164);
nor U9801 (N_9801,N_9463,N_9421);
or U9802 (N_9802,N_9444,N_9028);
nand U9803 (N_9803,N_9017,N_9381);
or U9804 (N_9804,N_9172,N_9419);
nor U9805 (N_9805,N_9067,N_9151);
nand U9806 (N_9806,N_9471,N_9200);
and U9807 (N_9807,N_9018,N_9212);
xnor U9808 (N_9808,N_9198,N_9272);
xnor U9809 (N_9809,N_9177,N_9212);
nor U9810 (N_9810,N_9414,N_9344);
or U9811 (N_9811,N_9062,N_9123);
and U9812 (N_9812,N_9035,N_9413);
and U9813 (N_9813,N_9370,N_9382);
nor U9814 (N_9814,N_9025,N_9379);
nor U9815 (N_9815,N_9047,N_9281);
nand U9816 (N_9816,N_9472,N_9465);
or U9817 (N_9817,N_9190,N_9354);
xor U9818 (N_9818,N_9118,N_9299);
nor U9819 (N_9819,N_9284,N_9412);
nand U9820 (N_9820,N_9064,N_9180);
nor U9821 (N_9821,N_9373,N_9006);
nor U9822 (N_9822,N_9049,N_9101);
or U9823 (N_9823,N_9438,N_9393);
xnor U9824 (N_9824,N_9271,N_9136);
and U9825 (N_9825,N_9005,N_9357);
and U9826 (N_9826,N_9376,N_9227);
and U9827 (N_9827,N_9141,N_9037);
and U9828 (N_9828,N_9411,N_9007);
and U9829 (N_9829,N_9234,N_9375);
and U9830 (N_9830,N_9113,N_9383);
xnor U9831 (N_9831,N_9098,N_9157);
or U9832 (N_9832,N_9370,N_9399);
and U9833 (N_9833,N_9214,N_9497);
nor U9834 (N_9834,N_9351,N_9498);
nor U9835 (N_9835,N_9495,N_9075);
nor U9836 (N_9836,N_9126,N_9060);
and U9837 (N_9837,N_9044,N_9082);
and U9838 (N_9838,N_9307,N_9393);
xor U9839 (N_9839,N_9376,N_9487);
or U9840 (N_9840,N_9452,N_9442);
and U9841 (N_9841,N_9357,N_9194);
nor U9842 (N_9842,N_9250,N_9388);
nor U9843 (N_9843,N_9483,N_9026);
or U9844 (N_9844,N_9225,N_9019);
nor U9845 (N_9845,N_9197,N_9366);
nor U9846 (N_9846,N_9482,N_9137);
and U9847 (N_9847,N_9322,N_9305);
or U9848 (N_9848,N_9124,N_9353);
xnor U9849 (N_9849,N_9455,N_9385);
nor U9850 (N_9850,N_9281,N_9381);
nor U9851 (N_9851,N_9335,N_9025);
and U9852 (N_9852,N_9066,N_9013);
nor U9853 (N_9853,N_9455,N_9107);
nand U9854 (N_9854,N_9028,N_9273);
nand U9855 (N_9855,N_9135,N_9404);
xor U9856 (N_9856,N_9359,N_9019);
and U9857 (N_9857,N_9330,N_9449);
nand U9858 (N_9858,N_9083,N_9400);
and U9859 (N_9859,N_9397,N_9415);
and U9860 (N_9860,N_9025,N_9172);
nand U9861 (N_9861,N_9442,N_9310);
and U9862 (N_9862,N_9073,N_9495);
xor U9863 (N_9863,N_9090,N_9214);
nor U9864 (N_9864,N_9332,N_9126);
and U9865 (N_9865,N_9429,N_9050);
nor U9866 (N_9866,N_9325,N_9458);
nand U9867 (N_9867,N_9068,N_9098);
nor U9868 (N_9868,N_9481,N_9071);
and U9869 (N_9869,N_9018,N_9427);
and U9870 (N_9870,N_9062,N_9198);
xnor U9871 (N_9871,N_9046,N_9254);
and U9872 (N_9872,N_9294,N_9006);
and U9873 (N_9873,N_9018,N_9046);
and U9874 (N_9874,N_9122,N_9373);
or U9875 (N_9875,N_9388,N_9274);
and U9876 (N_9876,N_9177,N_9048);
xnor U9877 (N_9877,N_9104,N_9134);
and U9878 (N_9878,N_9043,N_9307);
or U9879 (N_9879,N_9055,N_9017);
xnor U9880 (N_9880,N_9078,N_9190);
xor U9881 (N_9881,N_9086,N_9009);
or U9882 (N_9882,N_9308,N_9438);
nor U9883 (N_9883,N_9439,N_9368);
xnor U9884 (N_9884,N_9294,N_9387);
and U9885 (N_9885,N_9315,N_9433);
nor U9886 (N_9886,N_9175,N_9354);
nand U9887 (N_9887,N_9453,N_9233);
and U9888 (N_9888,N_9042,N_9489);
and U9889 (N_9889,N_9027,N_9021);
xor U9890 (N_9890,N_9010,N_9400);
nand U9891 (N_9891,N_9396,N_9215);
and U9892 (N_9892,N_9069,N_9352);
nand U9893 (N_9893,N_9335,N_9058);
xnor U9894 (N_9894,N_9361,N_9225);
nor U9895 (N_9895,N_9307,N_9407);
or U9896 (N_9896,N_9331,N_9074);
xor U9897 (N_9897,N_9150,N_9212);
nor U9898 (N_9898,N_9269,N_9076);
xor U9899 (N_9899,N_9410,N_9139);
xor U9900 (N_9900,N_9181,N_9424);
nand U9901 (N_9901,N_9490,N_9409);
and U9902 (N_9902,N_9263,N_9290);
xor U9903 (N_9903,N_9317,N_9185);
and U9904 (N_9904,N_9017,N_9331);
xor U9905 (N_9905,N_9094,N_9065);
xnor U9906 (N_9906,N_9336,N_9400);
and U9907 (N_9907,N_9107,N_9138);
xor U9908 (N_9908,N_9449,N_9073);
xnor U9909 (N_9909,N_9469,N_9453);
and U9910 (N_9910,N_9048,N_9495);
and U9911 (N_9911,N_9121,N_9190);
xnor U9912 (N_9912,N_9330,N_9120);
nor U9913 (N_9913,N_9249,N_9009);
nand U9914 (N_9914,N_9345,N_9401);
xor U9915 (N_9915,N_9127,N_9041);
nand U9916 (N_9916,N_9002,N_9359);
nor U9917 (N_9917,N_9377,N_9000);
or U9918 (N_9918,N_9471,N_9175);
nor U9919 (N_9919,N_9164,N_9445);
and U9920 (N_9920,N_9185,N_9294);
nor U9921 (N_9921,N_9313,N_9085);
nand U9922 (N_9922,N_9281,N_9319);
and U9923 (N_9923,N_9161,N_9291);
or U9924 (N_9924,N_9151,N_9236);
and U9925 (N_9925,N_9373,N_9138);
and U9926 (N_9926,N_9244,N_9094);
or U9927 (N_9927,N_9045,N_9307);
xor U9928 (N_9928,N_9008,N_9195);
nand U9929 (N_9929,N_9248,N_9314);
nor U9930 (N_9930,N_9263,N_9081);
xor U9931 (N_9931,N_9422,N_9100);
nor U9932 (N_9932,N_9106,N_9145);
or U9933 (N_9933,N_9216,N_9439);
or U9934 (N_9934,N_9137,N_9351);
nand U9935 (N_9935,N_9191,N_9342);
nor U9936 (N_9936,N_9273,N_9220);
xnor U9937 (N_9937,N_9240,N_9336);
xnor U9938 (N_9938,N_9122,N_9462);
nand U9939 (N_9939,N_9463,N_9187);
xnor U9940 (N_9940,N_9309,N_9389);
nor U9941 (N_9941,N_9417,N_9389);
xor U9942 (N_9942,N_9376,N_9369);
and U9943 (N_9943,N_9096,N_9489);
nand U9944 (N_9944,N_9258,N_9389);
nand U9945 (N_9945,N_9249,N_9055);
or U9946 (N_9946,N_9088,N_9245);
xnor U9947 (N_9947,N_9254,N_9084);
or U9948 (N_9948,N_9293,N_9137);
xnor U9949 (N_9949,N_9267,N_9315);
and U9950 (N_9950,N_9350,N_9117);
and U9951 (N_9951,N_9461,N_9009);
xnor U9952 (N_9952,N_9121,N_9020);
nor U9953 (N_9953,N_9088,N_9177);
and U9954 (N_9954,N_9099,N_9279);
nor U9955 (N_9955,N_9145,N_9185);
and U9956 (N_9956,N_9038,N_9169);
and U9957 (N_9957,N_9497,N_9371);
and U9958 (N_9958,N_9108,N_9063);
or U9959 (N_9959,N_9181,N_9427);
and U9960 (N_9960,N_9270,N_9261);
xnor U9961 (N_9961,N_9105,N_9077);
nor U9962 (N_9962,N_9492,N_9006);
nand U9963 (N_9963,N_9036,N_9372);
nand U9964 (N_9964,N_9150,N_9080);
or U9965 (N_9965,N_9069,N_9172);
and U9966 (N_9966,N_9204,N_9236);
nor U9967 (N_9967,N_9030,N_9361);
and U9968 (N_9968,N_9260,N_9129);
nand U9969 (N_9969,N_9197,N_9218);
nand U9970 (N_9970,N_9138,N_9156);
nand U9971 (N_9971,N_9051,N_9241);
xor U9972 (N_9972,N_9255,N_9178);
nor U9973 (N_9973,N_9097,N_9381);
or U9974 (N_9974,N_9361,N_9187);
and U9975 (N_9975,N_9333,N_9029);
nor U9976 (N_9976,N_9315,N_9029);
or U9977 (N_9977,N_9167,N_9063);
nand U9978 (N_9978,N_9470,N_9122);
or U9979 (N_9979,N_9125,N_9338);
and U9980 (N_9980,N_9452,N_9478);
xnor U9981 (N_9981,N_9185,N_9490);
or U9982 (N_9982,N_9308,N_9010);
nand U9983 (N_9983,N_9368,N_9158);
and U9984 (N_9984,N_9428,N_9177);
or U9985 (N_9985,N_9091,N_9432);
or U9986 (N_9986,N_9099,N_9408);
and U9987 (N_9987,N_9476,N_9272);
and U9988 (N_9988,N_9288,N_9345);
nor U9989 (N_9989,N_9109,N_9489);
nor U9990 (N_9990,N_9272,N_9040);
nand U9991 (N_9991,N_9444,N_9320);
or U9992 (N_9992,N_9335,N_9007);
or U9993 (N_9993,N_9290,N_9479);
or U9994 (N_9994,N_9183,N_9396);
nand U9995 (N_9995,N_9292,N_9332);
nor U9996 (N_9996,N_9129,N_9391);
or U9997 (N_9997,N_9310,N_9419);
or U9998 (N_9998,N_9290,N_9007);
nand U9999 (N_9999,N_9059,N_9171);
and U10000 (N_10000,N_9690,N_9777);
or U10001 (N_10001,N_9618,N_9974);
nor U10002 (N_10002,N_9887,N_9709);
nand U10003 (N_10003,N_9877,N_9570);
nor U10004 (N_10004,N_9504,N_9822);
nand U10005 (N_10005,N_9846,N_9872);
nand U10006 (N_10006,N_9585,N_9999);
nand U10007 (N_10007,N_9672,N_9766);
and U10008 (N_10008,N_9749,N_9513);
and U10009 (N_10009,N_9988,N_9686);
and U10010 (N_10010,N_9806,N_9623);
nand U10011 (N_10011,N_9732,N_9918);
xnor U10012 (N_10012,N_9910,N_9971);
nor U10013 (N_10013,N_9949,N_9747);
xor U10014 (N_10014,N_9557,N_9642);
nor U10015 (N_10015,N_9700,N_9738);
nand U10016 (N_10016,N_9679,N_9631);
or U10017 (N_10017,N_9848,N_9780);
or U10018 (N_10018,N_9650,N_9677);
or U10019 (N_10019,N_9647,N_9879);
nand U10020 (N_10020,N_9892,N_9836);
and U10021 (N_10021,N_9621,N_9997);
or U10022 (N_10022,N_9832,N_9627);
or U10023 (N_10023,N_9763,N_9838);
nand U10024 (N_10024,N_9519,N_9615);
xor U10025 (N_10025,N_9691,N_9626);
nand U10026 (N_10026,N_9609,N_9937);
nand U10027 (N_10027,N_9592,N_9904);
xor U10028 (N_10028,N_9710,N_9753);
xor U10029 (N_10029,N_9678,N_9707);
or U10030 (N_10030,N_9829,N_9587);
and U10031 (N_10031,N_9956,N_9975);
xnor U10032 (N_10032,N_9617,N_9771);
nand U10033 (N_10033,N_9600,N_9545);
nor U10034 (N_10034,N_9919,N_9880);
and U10035 (N_10035,N_9718,N_9554);
xor U10036 (N_10036,N_9522,N_9851);
or U10037 (N_10037,N_9509,N_9696);
nand U10038 (N_10038,N_9952,N_9885);
nor U10039 (N_10039,N_9957,N_9648);
and U10040 (N_10040,N_9932,N_9850);
xnor U10041 (N_10041,N_9538,N_9940);
and U10042 (N_10042,N_9576,N_9756);
nor U10043 (N_10043,N_9767,N_9722);
xor U10044 (N_10044,N_9544,N_9794);
or U10045 (N_10045,N_9665,N_9673);
xor U10046 (N_10046,N_9982,N_9843);
nor U10047 (N_10047,N_9841,N_9898);
xnor U10048 (N_10048,N_9531,N_9693);
nand U10049 (N_10049,N_9876,N_9955);
xor U10050 (N_10050,N_9998,N_9800);
and U10051 (N_10051,N_9614,N_9827);
xnor U10052 (N_10052,N_9658,N_9757);
nand U10053 (N_10053,N_9933,N_9962);
xor U10054 (N_10054,N_9640,N_9868);
xor U10055 (N_10055,N_9731,N_9994);
nand U10056 (N_10056,N_9584,N_9636);
nand U10057 (N_10057,N_9938,N_9697);
and U10058 (N_10058,N_9859,N_9858);
nor U10059 (N_10059,N_9951,N_9840);
xor U10060 (N_10060,N_9849,N_9842);
nor U10061 (N_10061,N_9863,N_9525);
and U10062 (N_10062,N_9801,N_9810);
or U10063 (N_10063,N_9629,N_9993);
or U10064 (N_10064,N_9534,N_9628);
xor U10065 (N_10065,N_9856,N_9635);
and U10066 (N_10066,N_9946,N_9907);
or U10067 (N_10067,N_9903,N_9987);
xnor U10068 (N_10068,N_9921,N_9797);
nor U10069 (N_10069,N_9733,N_9581);
and U10070 (N_10070,N_9969,N_9637);
xnor U10071 (N_10071,N_9713,N_9524);
and U10072 (N_10072,N_9689,N_9549);
nor U10073 (N_10073,N_9813,N_9820);
or U10074 (N_10074,N_9518,N_9819);
or U10075 (N_10075,N_9839,N_9764);
or U10076 (N_10076,N_9541,N_9878);
nor U10077 (N_10077,N_9873,N_9726);
or U10078 (N_10078,N_9865,N_9936);
or U10079 (N_10079,N_9579,N_9977);
and U10080 (N_10080,N_9651,N_9608);
or U10081 (N_10081,N_9695,N_9663);
nor U10082 (N_10082,N_9681,N_9888);
nand U10083 (N_10083,N_9620,N_9536);
and U10084 (N_10084,N_9565,N_9785);
nand U10085 (N_10085,N_9929,N_9564);
xnor U10086 (N_10086,N_9506,N_9744);
or U10087 (N_10087,N_9824,N_9791);
and U10088 (N_10088,N_9669,N_9743);
or U10089 (N_10089,N_9594,N_9721);
nor U10090 (N_10090,N_9643,N_9563);
nand U10091 (N_10091,N_9502,N_9899);
nor U10092 (N_10092,N_9566,N_9884);
nor U10093 (N_10093,N_9543,N_9928);
nor U10094 (N_10094,N_9772,N_9769);
or U10095 (N_10095,N_9908,N_9860);
or U10096 (N_10096,N_9688,N_9912);
and U10097 (N_10097,N_9817,N_9597);
nor U10098 (N_10098,N_9990,N_9625);
nor U10099 (N_10099,N_9553,N_9740);
xnor U10100 (N_10100,N_9529,N_9533);
or U10101 (N_10101,N_9501,N_9857);
xnor U10102 (N_10102,N_9653,N_9532);
xor U10103 (N_10103,N_9925,N_9634);
nand U10104 (N_10104,N_9583,N_9755);
nand U10105 (N_10105,N_9901,N_9917);
or U10106 (N_10106,N_9909,N_9891);
nand U10107 (N_10107,N_9889,N_9963);
xor U10108 (N_10108,N_9598,N_9516);
xnor U10109 (N_10109,N_9805,N_9811);
xor U10110 (N_10110,N_9599,N_9630);
nand U10111 (N_10111,N_9922,N_9708);
xor U10112 (N_10112,N_9652,N_9881);
nand U10113 (N_10113,N_9604,N_9567);
xor U10114 (N_10114,N_9790,N_9862);
or U10115 (N_10115,N_9793,N_9715);
or U10116 (N_10116,N_9735,N_9638);
or U10117 (N_10117,N_9900,N_9573);
xnor U10118 (N_10118,N_9542,N_9560);
nand U10119 (N_10119,N_9844,N_9588);
and U10120 (N_10120,N_9702,N_9894);
nand U10121 (N_10121,N_9816,N_9762);
nor U10122 (N_10122,N_9507,N_9537);
nor U10123 (N_10123,N_9751,N_9510);
and U10124 (N_10124,N_9748,N_9720);
nor U10125 (N_10125,N_9883,N_9935);
nand U10126 (N_10126,N_9986,N_9562);
and U10127 (N_10127,N_9976,N_9633);
or U10128 (N_10128,N_9812,N_9984);
nor U10129 (N_10129,N_9779,N_9947);
nand U10130 (N_10130,N_9815,N_9979);
xor U10131 (N_10131,N_9703,N_9953);
and U10132 (N_10132,N_9520,N_9568);
nand U10133 (N_10133,N_9970,N_9692);
or U10134 (N_10134,N_9895,N_9613);
nand U10135 (N_10135,N_9991,N_9833);
and U10136 (N_10136,N_9578,N_9978);
xor U10137 (N_10137,N_9742,N_9835);
nor U10138 (N_10138,N_9734,N_9814);
xnor U10139 (N_10139,N_9804,N_9716);
or U10140 (N_10140,N_9964,N_9589);
and U10141 (N_10141,N_9717,N_9959);
nand U10142 (N_10142,N_9622,N_9577);
or U10143 (N_10143,N_9983,N_9965);
or U10144 (N_10144,N_9701,N_9792);
xnor U10145 (N_10145,N_9818,N_9927);
and U10146 (N_10146,N_9931,N_9985);
and U10147 (N_10147,N_9641,N_9923);
or U10148 (N_10148,N_9809,N_9656);
nand U10149 (N_10149,N_9612,N_9556);
or U10150 (N_10150,N_9788,N_9661);
or U10151 (N_10151,N_9645,N_9761);
and U10152 (N_10152,N_9593,N_9550);
nor U10153 (N_10153,N_9992,N_9837);
nand U10154 (N_10154,N_9765,N_9760);
and U10155 (N_10155,N_9803,N_9770);
nand U10156 (N_10156,N_9714,N_9505);
nor U10157 (N_10157,N_9853,N_9607);
nor U10158 (N_10158,N_9754,N_9911);
nand U10159 (N_10159,N_9528,N_9741);
and U10160 (N_10160,N_9610,N_9914);
xor U10161 (N_10161,N_9941,N_9575);
and U10162 (N_10162,N_9540,N_9930);
xnor U10163 (N_10163,N_9739,N_9569);
nand U10164 (N_10164,N_9896,N_9954);
nor U10165 (N_10165,N_9616,N_9727);
and U10166 (N_10166,N_9920,N_9905);
or U10167 (N_10167,N_9611,N_9552);
xor U10168 (N_10168,N_9605,N_9867);
xor U10169 (N_10169,N_9527,N_9834);
xor U10170 (N_10170,N_9778,N_9723);
and U10171 (N_10171,N_9596,N_9795);
nand U10172 (N_10172,N_9752,N_9632);
xor U10173 (N_10173,N_9773,N_9666);
nor U10174 (N_10174,N_9644,N_9826);
or U10175 (N_10175,N_9646,N_9870);
or U10176 (N_10176,N_9852,N_9893);
xor U10177 (N_10177,N_9730,N_9559);
and U10178 (N_10178,N_9847,N_9775);
or U10179 (N_10179,N_9861,N_9728);
and U10180 (N_10180,N_9874,N_9875);
or U10181 (N_10181,N_9967,N_9758);
nor U10182 (N_10182,N_9948,N_9668);
and U10183 (N_10183,N_9698,N_9624);
and U10184 (N_10184,N_9704,N_9582);
or U10185 (N_10185,N_9574,N_9591);
nor U10186 (N_10186,N_9706,N_9966);
or U10187 (N_10187,N_9670,N_9750);
and U10188 (N_10188,N_9886,N_9864);
nor U10189 (N_10189,N_9547,N_9786);
nand U10190 (N_10190,N_9561,N_9699);
and U10191 (N_10191,N_9590,N_9572);
and U10192 (N_10192,N_9551,N_9807);
nand U10193 (N_10193,N_9828,N_9960);
or U10194 (N_10194,N_9659,N_9711);
or U10195 (N_10195,N_9737,N_9958);
xor U10196 (N_10196,N_9783,N_9725);
and U10197 (N_10197,N_9890,N_9664);
nor U10198 (N_10198,N_9657,N_9687);
nor U10199 (N_10199,N_9897,N_9784);
and U10200 (N_10200,N_9526,N_9802);
or U10201 (N_10201,N_9662,N_9705);
nand U10202 (N_10202,N_9972,N_9586);
xor U10203 (N_10203,N_9759,N_9831);
xor U10204 (N_10204,N_9535,N_9667);
nor U10205 (N_10205,N_9676,N_9654);
nor U10206 (N_10206,N_9546,N_9845);
nor U10207 (N_10207,N_9508,N_9639);
and U10208 (N_10208,N_9973,N_9798);
nor U10209 (N_10209,N_9511,N_9674);
xnor U10210 (N_10210,N_9712,N_9796);
nor U10211 (N_10211,N_9980,N_9736);
xor U10212 (N_10212,N_9683,N_9950);
or U10213 (N_10213,N_9512,N_9830);
nor U10214 (N_10214,N_9916,N_9961);
nor U10215 (N_10215,N_9924,N_9671);
xor U10216 (N_10216,N_9781,N_9968);
xnor U10217 (N_10217,N_9539,N_9854);
and U10218 (N_10218,N_9774,N_9571);
nand U10219 (N_10219,N_9869,N_9823);
or U10220 (N_10220,N_9649,N_9787);
xnor U10221 (N_10221,N_9724,N_9619);
xnor U10222 (N_10222,N_9580,N_9768);
and U10223 (N_10223,N_9995,N_9521);
or U10224 (N_10224,N_9926,N_9746);
nand U10225 (N_10225,N_9808,N_9981);
or U10226 (N_10226,N_9660,N_9530);
nor U10227 (N_10227,N_9555,N_9943);
nand U10228 (N_10228,N_9799,N_9944);
nand U10229 (N_10229,N_9934,N_9548);
and U10230 (N_10230,N_9680,N_9601);
and U10231 (N_10231,N_9595,N_9866);
xnor U10232 (N_10232,N_9685,N_9821);
nor U10233 (N_10233,N_9655,N_9915);
nor U10234 (N_10234,N_9558,N_9789);
or U10235 (N_10235,N_9515,N_9500);
and U10236 (N_10236,N_9902,N_9945);
and U10237 (N_10237,N_9719,N_9606);
and U10238 (N_10238,N_9523,N_9745);
and U10239 (N_10239,N_9871,N_9989);
nand U10240 (N_10240,N_9694,N_9503);
nand U10241 (N_10241,N_9913,N_9882);
and U10242 (N_10242,N_9514,N_9906);
xor U10243 (N_10243,N_9825,N_9776);
nand U10244 (N_10244,N_9603,N_9729);
nor U10245 (N_10245,N_9942,N_9684);
and U10246 (N_10246,N_9996,N_9675);
and U10247 (N_10247,N_9517,N_9855);
nor U10248 (N_10248,N_9782,N_9939);
nand U10249 (N_10249,N_9602,N_9682);
xor U10250 (N_10250,N_9873,N_9770);
nand U10251 (N_10251,N_9878,N_9943);
nor U10252 (N_10252,N_9647,N_9589);
or U10253 (N_10253,N_9651,N_9733);
nor U10254 (N_10254,N_9869,N_9892);
xnor U10255 (N_10255,N_9808,N_9583);
and U10256 (N_10256,N_9621,N_9528);
nor U10257 (N_10257,N_9564,N_9600);
nand U10258 (N_10258,N_9841,N_9586);
nor U10259 (N_10259,N_9717,N_9549);
nor U10260 (N_10260,N_9636,N_9696);
nor U10261 (N_10261,N_9980,N_9681);
and U10262 (N_10262,N_9955,N_9622);
or U10263 (N_10263,N_9900,N_9619);
nand U10264 (N_10264,N_9848,N_9845);
or U10265 (N_10265,N_9761,N_9609);
xor U10266 (N_10266,N_9647,N_9688);
xor U10267 (N_10267,N_9577,N_9811);
or U10268 (N_10268,N_9638,N_9639);
nor U10269 (N_10269,N_9758,N_9818);
nor U10270 (N_10270,N_9695,N_9783);
nor U10271 (N_10271,N_9712,N_9746);
nand U10272 (N_10272,N_9962,N_9623);
or U10273 (N_10273,N_9985,N_9917);
and U10274 (N_10274,N_9535,N_9838);
nand U10275 (N_10275,N_9797,N_9567);
xor U10276 (N_10276,N_9723,N_9981);
or U10277 (N_10277,N_9769,N_9554);
and U10278 (N_10278,N_9862,N_9694);
and U10279 (N_10279,N_9974,N_9985);
nor U10280 (N_10280,N_9739,N_9600);
nand U10281 (N_10281,N_9696,N_9684);
xor U10282 (N_10282,N_9848,N_9560);
or U10283 (N_10283,N_9973,N_9524);
nand U10284 (N_10284,N_9914,N_9828);
and U10285 (N_10285,N_9807,N_9857);
or U10286 (N_10286,N_9552,N_9963);
nand U10287 (N_10287,N_9506,N_9927);
nand U10288 (N_10288,N_9556,N_9744);
xor U10289 (N_10289,N_9837,N_9766);
and U10290 (N_10290,N_9800,N_9708);
xor U10291 (N_10291,N_9926,N_9939);
xnor U10292 (N_10292,N_9555,N_9906);
or U10293 (N_10293,N_9987,N_9847);
or U10294 (N_10294,N_9534,N_9708);
and U10295 (N_10295,N_9977,N_9834);
or U10296 (N_10296,N_9893,N_9559);
nor U10297 (N_10297,N_9795,N_9771);
or U10298 (N_10298,N_9625,N_9912);
and U10299 (N_10299,N_9592,N_9789);
nand U10300 (N_10300,N_9972,N_9627);
xnor U10301 (N_10301,N_9939,N_9593);
nand U10302 (N_10302,N_9541,N_9751);
xor U10303 (N_10303,N_9591,N_9828);
or U10304 (N_10304,N_9794,N_9904);
or U10305 (N_10305,N_9878,N_9738);
nor U10306 (N_10306,N_9531,N_9976);
nor U10307 (N_10307,N_9652,N_9736);
or U10308 (N_10308,N_9690,N_9921);
nand U10309 (N_10309,N_9637,N_9886);
or U10310 (N_10310,N_9622,N_9760);
nor U10311 (N_10311,N_9832,N_9833);
xor U10312 (N_10312,N_9878,N_9539);
nor U10313 (N_10313,N_9888,N_9857);
nor U10314 (N_10314,N_9898,N_9768);
xnor U10315 (N_10315,N_9682,N_9516);
or U10316 (N_10316,N_9907,N_9621);
or U10317 (N_10317,N_9551,N_9503);
and U10318 (N_10318,N_9824,N_9745);
or U10319 (N_10319,N_9889,N_9561);
nand U10320 (N_10320,N_9712,N_9965);
xnor U10321 (N_10321,N_9659,N_9691);
and U10322 (N_10322,N_9988,N_9802);
and U10323 (N_10323,N_9634,N_9827);
nor U10324 (N_10324,N_9663,N_9960);
xnor U10325 (N_10325,N_9971,N_9560);
xnor U10326 (N_10326,N_9981,N_9617);
or U10327 (N_10327,N_9974,N_9611);
and U10328 (N_10328,N_9923,N_9632);
and U10329 (N_10329,N_9766,N_9783);
and U10330 (N_10330,N_9700,N_9584);
and U10331 (N_10331,N_9838,N_9549);
and U10332 (N_10332,N_9712,N_9592);
nand U10333 (N_10333,N_9967,N_9638);
xnor U10334 (N_10334,N_9767,N_9803);
nor U10335 (N_10335,N_9518,N_9680);
or U10336 (N_10336,N_9605,N_9858);
and U10337 (N_10337,N_9666,N_9646);
nand U10338 (N_10338,N_9664,N_9603);
and U10339 (N_10339,N_9623,N_9621);
xnor U10340 (N_10340,N_9513,N_9879);
nor U10341 (N_10341,N_9918,N_9742);
or U10342 (N_10342,N_9607,N_9527);
nand U10343 (N_10343,N_9806,N_9878);
nand U10344 (N_10344,N_9578,N_9796);
or U10345 (N_10345,N_9666,N_9714);
nor U10346 (N_10346,N_9847,N_9734);
and U10347 (N_10347,N_9572,N_9978);
and U10348 (N_10348,N_9831,N_9685);
or U10349 (N_10349,N_9902,N_9711);
or U10350 (N_10350,N_9733,N_9649);
and U10351 (N_10351,N_9630,N_9570);
nand U10352 (N_10352,N_9925,N_9685);
and U10353 (N_10353,N_9749,N_9695);
nor U10354 (N_10354,N_9506,N_9610);
and U10355 (N_10355,N_9584,N_9856);
and U10356 (N_10356,N_9678,N_9792);
xnor U10357 (N_10357,N_9870,N_9510);
or U10358 (N_10358,N_9559,N_9580);
xor U10359 (N_10359,N_9975,N_9660);
nand U10360 (N_10360,N_9540,N_9793);
or U10361 (N_10361,N_9758,N_9688);
xor U10362 (N_10362,N_9936,N_9963);
or U10363 (N_10363,N_9996,N_9691);
nand U10364 (N_10364,N_9868,N_9992);
nand U10365 (N_10365,N_9618,N_9972);
xnor U10366 (N_10366,N_9571,N_9533);
or U10367 (N_10367,N_9580,N_9798);
and U10368 (N_10368,N_9607,N_9665);
nand U10369 (N_10369,N_9582,N_9975);
xnor U10370 (N_10370,N_9523,N_9586);
and U10371 (N_10371,N_9808,N_9964);
nand U10372 (N_10372,N_9879,N_9627);
nor U10373 (N_10373,N_9624,N_9595);
nor U10374 (N_10374,N_9794,N_9723);
nor U10375 (N_10375,N_9680,N_9919);
or U10376 (N_10376,N_9980,N_9504);
xor U10377 (N_10377,N_9764,N_9815);
or U10378 (N_10378,N_9976,N_9644);
nand U10379 (N_10379,N_9720,N_9713);
or U10380 (N_10380,N_9681,N_9782);
or U10381 (N_10381,N_9707,N_9952);
nor U10382 (N_10382,N_9986,N_9549);
or U10383 (N_10383,N_9580,N_9720);
xnor U10384 (N_10384,N_9722,N_9801);
or U10385 (N_10385,N_9726,N_9923);
nand U10386 (N_10386,N_9929,N_9811);
nor U10387 (N_10387,N_9676,N_9735);
xor U10388 (N_10388,N_9551,N_9657);
nor U10389 (N_10389,N_9519,N_9924);
nand U10390 (N_10390,N_9610,N_9724);
or U10391 (N_10391,N_9947,N_9971);
and U10392 (N_10392,N_9953,N_9811);
or U10393 (N_10393,N_9633,N_9530);
and U10394 (N_10394,N_9798,N_9839);
and U10395 (N_10395,N_9993,N_9977);
xor U10396 (N_10396,N_9512,N_9858);
or U10397 (N_10397,N_9859,N_9813);
nand U10398 (N_10398,N_9928,N_9690);
xnor U10399 (N_10399,N_9595,N_9728);
and U10400 (N_10400,N_9618,N_9559);
and U10401 (N_10401,N_9959,N_9810);
or U10402 (N_10402,N_9576,N_9585);
nand U10403 (N_10403,N_9669,N_9595);
nor U10404 (N_10404,N_9651,N_9787);
and U10405 (N_10405,N_9828,N_9844);
xor U10406 (N_10406,N_9694,N_9769);
nor U10407 (N_10407,N_9957,N_9916);
and U10408 (N_10408,N_9698,N_9725);
xnor U10409 (N_10409,N_9806,N_9817);
nor U10410 (N_10410,N_9798,N_9657);
nand U10411 (N_10411,N_9692,N_9671);
nor U10412 (N_10412,N_9859,N_9688);
nand U10413 (N_10413,N_9683,N_9589);
and U10414 (N_10414,N_9864,N_9941);
and U10415 (N_10415,N_9898,N_9954);
or U10416 (N_10416,N_9601,N_9903);
nand U10417 (N_10417,N_9620,N_9924);
xor U10418 (N_10418,N_9545,N_9936);
or U10419 (N_10419,N_9548,N_9831);
nor U10420 (N_10420,N_9902,N_9562);
xnor U10421 (N_10421,N_9721,N_9954);
and U10422 (N_10422,N_9932,N_9893);
or U10423 (N_10423,N_9582,N_9815);
and U10424 (N_10424,N_9889,N_9580);
nor U10425 (N_10425,N_9526,N_9833);
and U10426 (N_10426,N_9777,N_9609);
xor U10427 (N_10427,N_9900,N_9979);
xnor U10428 (N_10428,N_9998,N_9879);
nor U10429 (N_10429,N_9744,N_9976);
nor U10430 (N_10430,N_9575,N_9757);
xnor U10431 (N_10431,N_9808,N_9613);
or U10432 (N_10432,N_9564,N_9755);
nor U10433 (N_10433,N_9979,N_9818);
nor U10434 (N_10434,N_9871,N_9927);
and U10435 (N_10435,N_9568,N_9709);
nor U10436 (N_10436,N_9784,N_9837);
or U10437 (N_10437,N_9754,N_9930);
xor U10438 (N_10438,N_9589,N_9992);
or U10439 (N_10439,N_9575,N_9843);
xnor U10440 (N_10440,N_9952,N_9881);
or U10441 (N_10441,N_9523,N_9676);
or U10442 (N_10442,N_9818,N_9911);
and U10443 (N_10443,N_9786,N_9815);
nor U10444 (N_10444,N_9911,N_9836);
xnor U10445 (N_10445,N_9950,N_9946);
nand U10446 (N_10446,N_9953,N_9534);
and U10447 (N_10447,N_9971,N_9891);
or U10448 (N_10448,N_9578,N_9613);
xnor U10449 (N_10449,N_9962,N_9830);
nand U10450 (N_10450,N_9977,N_9955);
nor U10451 (N_10451,N_9964,N_9968);
nand U10452 (N_10452,N_9927,N_9868);
xor U10453 (N_10453,N_9603,N_9977);
or U10454 (N_10454,N_9635,N_9644);
or U10455 (N_10455,N_9962,N_9573);
xor U10456 (N_10456,N_9529,N_9566);
nor U10457 (N_10457,N_9805,N_9899);
nand U10458 (N_10458,N_9943,N_9797);
nand U10459 (N_10459,N_9954,N_9673);
and U10460 (N_10460,N_9535,N_9612);
xor U10461 (N_10461,N_9975,N_9678);
nand U10462 (N_10462,N_9929,N_9606);
nor U10463 (N_10463,N_9946,N_9510);
xor U10464 (N_10464,N_9739,N_9781);
xnor U10465 (N_10465,N_9582,N_9663);
and U10466 (N_10466,N_9571,N_9620);
nand U10467 (N_10467,N_9667,N_9500);
nor U10468 (N_10468,N_9561,N_9722);
and U10469 (N_10469,N_9698,N_9821);
xor U10470 (N_10470,N_9660,N_9789);
nor U10471 (N_10471,N_9528,N_9558);
and U10472 (N_10472,N_9746,N_9945);
and U10473 (N_10473,N_9971,N_9501);
and U10474 (N_10474,N_9667,N_9815);
or U10475 (N_10475,N_9500,N_9600);
xor U10476 (N_10476,N_9981,N_9855);
xor U10477 (N_10477,N_9723,N_9865);
or U10478 (N_10478,N_9643,N_9797);
and U10479 (N_10479,N_9951,N_9565);
and U10480 (N_10480,N_9668,N_9672);
nor U10481 (N_10481,N_9636,N_9703);
nand U10482 (N_10482,N_9654,N_9819);
and U10483 (N_10483,N_9993,N_9541);
nor U10484 (N_10484,N_9834,N_9599);
or U10485 (N_10485,N_9572,N_9551);
and U10486 (N_10486,N_9674,N_9545);
nand U10487 (N_10487,N_9661,N_9800);
xnor U10488 (N_10488,N_9617,N_9689);
nand U10489 (N_10489,N_9655,N_9934);
nor U10490 (N_10490,N_9686,N_9508);
nand U10491 (N_10491,N_9818,N_9625);
nand U10492 (N_10492,N_9914,N_9660);
xor U10493 (N_10493,N_9548,N_9725);
and U10494 (N_10494,N_9857,N_9552);
nor U10495 (N_10495,N_9977,N_9879);
and U10496 (N_10496,N_9770,N_9514);
or U10497 (N_10497,N_9773,N_9966);
nand U10498 (N_10498,N_9733,N_9671);
and U10499 (N_10499,N_9863,N_9868);
and U10500 (N_10500,N_10408,N_10057);
nor U10501 (N_10501,N_10104,N_10005);
nor U10502 (N_10502,N_10031,N_10073);
nor U10503 (N_10503,N_10422,N_10130);
or U10504 (N_10504,N_10294,N_10330);
nor U10505 (N_10505,N_10495,N_10204);
or U10506 (N_10506,N_10424,N_10065);
and U10507 (N_10507,N_10351,N_10440);
xnor U10508 (N_10508,N_10215,N_10076);
or U10509 (N_10509,N_10323,N_10121);
nor U10510 (N_10510,N_10273,N_10433);
xor U10511 (N_10511,N_10372,N_10193);
nand U10512 (N_10512,N_10167,N_10345);
nor U10513 (N_10513,N_10151,N_10080);
and U10514 (N_10514,N_10385,N_10418);
nor U10515 (N_10515,N_10075,N_10211);
or U10516 (N_10516,N_10149,N_10302);
nor U10517 (N_10517,N_10056,N_10441);
xnor U10518 (N_10518,N_10474,N_10340);
or U10519 (N_10519,N_10050,N_10079);
or U10520 (N_10520,N_10451,N_10335);
and U10521 (N_10521,N_10048,N_10216);
xnor U10522 (N_10522,N_10404,N_10152);
or U10523 (N_10523,N_10009,N_10192);
xor U10524 (N_10524,N_10012,N_10169);
xor U10525 (N_10525,N_10450,N_10489);
xor U10526 (N_10526,N_10324,N_10061);
nand U10527 (N_10527,N_10431,N_10163);
xor U10528 (N_10528,N_10157,N_10174);
and U10529 (N_10529,N_10446,N_10242);
xor U10530 (N_10530,N_10485,N_10358);
and U10531 (N_10531,N_10382,N_10329);
and U10532 (N_10532,N_10363,N_10069);
or U10533 (N_10533,N_10352,N_10046);
nand U10534 (N_10534,N_10305,N_10331);
or U10535 (N_10535,N_10209,N_10112);
or U10536 (N_10536,N_10154,N_10334);
nand U10537 (N_10537,N_10300,N_10098);
nor U10538 (N_10538,N_10254,N_10405);
or U10539 (N_10539,N_10459,N_10371);
nor U10540 (N_10540,N_10359,N_10093);
and U10541 (N_10541,N_10191,N_10203);
nor U10542 (N_10542,N_10237,N_10486);
xor U10543 (N_10543,N_10150,N_10473);
nand U10544 (N_10544,N_10052,N_10325);
nand U10545 (N_10545,N_10219,N_10103);
nor U10546 (N_10546,N_10399,N_10230);
or U10547 (N_10547,N_10132,N_10176);
or U10548 (N_10548,N_10004,N_10170);
nand U10549 (N_10549,N_10053,N_10465);
nand U10550 (N_10550,N_10249,N_10160);
and U10551 (N_10551,N_10311,N_10417);
xnor U10552 (N_10552,N_10018,N_10309);
xor U10553 (N_10553,N_10042,N_10397);
xnor U10554 (N_10554,N_10247,N_10088);
nand U10555 (N_10555,N_10288,N_10128);
nor U10556 (N_10556,N_10124,N_10402);
xor U10557 (N_10557,N_10196,N_10341);
nor U10558 (N_10558,N_10387,N_10299);
and U10559 (N_10559,N_10458,N_10062);
nand U10560 (N_10560,N_10117,N_10162);
nor U10561 (N_10561,N_10036,N_10392);
xor U10562 (N_10562,N_10228,N_10333);
and U10563 (N_10563,N_10074,N_10161);
nor U10564 (N_10564,N_10183,N_10051);
nor U10565 (N_10565,N_10089,N_10493);
xor U10566 (N_10566,N_10155,N_10409);
nand U10567 (N_10567,N_10456,N_10339);
nor U10568 (N_10568,N_10308,N_10401);
and U10569 (N_10569,N_10058,N_10281);
nor U10570 (N_10570,N_10238,N_10202);
nor U10571 (N_10571,N_10264,N_10270);
nor U10572 (N_10572,N_10159,N_10426);
and U10573 (N_10573,N_10208,N_10258);
xnor U10574 (N_10574,N_10095,N_10147);
or U10575 (N_10575,N_10452,N_10472);
xor U10576 (N_10576,N_10410,N_10269);
nand U10577 (N_10577,N_10438,N_10086);
xnor U10578 (N_10578,N_10421,N_10097);
or U10579 (N_10579,N_10355,N_10184);
and U10580 (N_10580,N_10102,N_10129);
and U10581 (N_10581,N_10322,N_10388);
and U10582 (N_10582,N_10142,N_10415);
nand U10583 (N_10583,N_10252,N_10085);
and U10584 (N_10584,N_10034,N_10468);
xnor U10585 (N_10585,N_10108,N_10146);
nor U10586 (N_10586,N_10092,N_10127);
or U10587 (N_10587,N_10497,N_10317);
or U10588 (N_10588,N_10181,N_10318);
and U10589 (N_10589,N_10251,N_10448);
xnor U10590 (N_10590,N_10343,N_10398);
nand U10591 (N_10591,N_10266,N_10032);
nor U10592 (N_10592,N_10241,N_10059);
nand U10593 (N_10593,N_10122,N_10187);
or U10594 (N_10594,N_10475,N_10006);
or U10595 (N_10595,N_10442,N_10349);
nand U10596 (N_10596,N_10244,N_10153);
and U10597 (N_10597,N_10115,N_10416);
and U10598 (N_10598,N_10367,N_10419);
and U10599 (N_10599,N_10078,N_10413);
nand U10600 (N_10600,N_10235,N_10429);
nor U10601 (N_10601,N_10243,N_10297);
and U10602 (N_10602,N_10188,N_10360);
or U10603 (N_10603,N_10082,N_10227);
nor U10604 (N_10604,N_10123,N_10290);
or U10605 (N_10605,N_10453,N_10487);
nor U10606 (N_10606,N_10137,N_10282);
and U10607 (N_10607,N_10091,N_10172);
nor U10608 (N_10608,N_10384,N_10289);
xnor U10609 (N_10609,N_10220,N_10178);
xnor U10610 (N_10610,N_10250,N_10041);
nor U10611 (N_10611,N_10236,N_10490);
or U10612 (N_10612,N_10262,N_10284);
nor U10613 (N_10613,N_10411,N_10319);
or U10614 (N_10614,N_10260,N_10233);
and U10615 (N_10615,N_10276,N_10499);
or U10616 (N_10616,N_10435,N_10466);
nand U10617 (N_10617,N_10023,N_10222);
or U10618 (N_10618,N_10186,N_10423);
and U10619 (N_10619,N_10044,N_10301);
or U10620 (N_10620,N_10140,N_10210);
nand U10621 (N_10621,N_10463,N_10332);
or U10622 (N_10622,N_10027,N_10087);
or U10623 (N_10623,N_10481,N_10001);
xor U10624 (N_10624,N_10175,N_10179);
xor U10625 (N_10625,N_10439,N_10221);
and U10626 (N_10626,N_10229,N_10496);
or U10627 (N_10627,N_10190,N_10425);
nor U10628 (N_10628,N_10028,N_10370);
nand U10629 (N_10629,N_10195,N_10164);
and U10630 (N_10630,N_10099,N_10457);
and U10631 (N_10631,N_10267,N_10286);
nand U10632 (N_10632,N_10125,N_10047);
and U10633 (N_10633,N_10476,N_10200);
and U10634 (N_10634,N_10263,N_10107);
or U10635 (N_10635,N_10067,N_10436);
nor U10636 (N_10636,N_10198,N_10376);
and U10637 (N_10637,N_10096,N_10136);
and U10638 (N_10638,N_10428,N_10165);
and U10639 (N_10639,N_10315,N_10239);
nand U10640 (N_10640,N_10071,N_10390);
or U10641 (N_10641,N_10434,N_10158);
nor U10642 (N_10642,N_10105,N_10464);
or U10643 (N_10643,N_10484,N_10454);
xnor U10644 (N_10644,N_10396,N_10328);
nor U10645 (N_10645,N_10245,N_10437);
xor U10646 (N_10646,N_10101,N_10182);
or U10647 (N_10647,N_10498,N_10477);
and U10648 (N_10648,N_10491,N_10072);
xnor U10649 (N_10649,N_10467,N_10257);
or U10650 (N_10650,N_10407,N_10283);
or U10651 (N_10651,N_10060,N_10037);
and U10652 (N_10652,N_10010,N_10040);
or U10653 (N_10653,N_10391,N_10213);
nand U10654 (N_10654,N_10406,N_10038);
or U10655 (N_10655,N_10427,N_10455);
and U10656 (N_10656,N_10314,N_10015);
nand U10657 (N_10657,N_10145,N_10460);
and U10658 (N_10658,N_10109,N_10444);
or U10659 (N_10659,N_10357,N_10274);
or U10660 (N_10660,N_10177,N_10114);
xor U10661 (N_10661,N_10312,N_10008);
or U10662 (N_10662,N_10120,N_10106);
and U10663 (N_10663,N_10365,N_10225);
nor U10664 (N_10664,N_10166,N_10373);
or U10665 (N_10665,N_10389,N_10386);
or U10666 (N_10666,N_10253,N_10445);
or U10667 (N_10667,N_10492,N_10189);
nor U10668 (N_10668,N_10261,N_10256);
nand U10669 (N_10669,N_10346,N_10279);
nand U10670 (N_10670,N_10338,N_10400);
xor U10671 (N_10671,N_10070,N_10226);
or U10672 (N_10672,N_10347,N_10321);
or U10673 (N_10673,N_10064,N_10234);
or U10674 (N_10674,N_10030,N_10206);
or U10675 (N_10675,N_10138,N_10374);
and U10676 (N_10676,N_10483,N_10194);
nand U10677 (N_10677,N_10268,N_10039);
nand U10678 (N_10678,N_10197,N_10461);
and U10679 (N_10679,N_10063,N_10081);
nand U10680 (N_10680,N_10271,N_10224);
nor U10681 (N_10681,N_10135,N_10113);
xor U10682 (N_10682,N_10139,N_10231);
xor U10683 (N_10683,N_10207,N_10369);
or U10684 (N_10684,N_10443,N_10381);
nand U10685 (N_10685,N_10310,N_10021);
xnor U10686 (N_10686,N_10110,N_10144);
or U10687 (N_10687,N_10043,N_10470);
nand U10688 (N_10688,N_10316,N_10205);
or U10689 (N_10689,N_10143,N_10111);
nand U10690 (N_10690,N_10077,N_10116);
nor U10691 (N_10691,N_10180,N_10275);
xnor U10692 (N_10692,N_10218,N_10118);
or U10693 (N_10693,N_10296,N_10024);
nand U10694 (N_10694,N_10049,N_10248);
xor U10695 (N_10695,N_10094,N_10214);
xnor U10696 (N_10696,N_10432,N_10232);
or U10697 (N_10697,N_10011,N_10126);
nor U10698 (N_10698,N_10326,N_10393);
and U10699 (N_10699,N_10033,N_10482);
xnor U10700 (N_10700,N_10320,N_10488);
nand U10701 (N_10701,N_10016,N_10020);
or U10702 (N_10702,N_10019,N_10265);
or U10703 (N_10703,N_10000,N_10494);
nand U10704 (N_10704,N_10272,N_10469);
nand U10705 (N_10705,N_10480,N_10378);
or U10706 (N_10706,N_10055,N_10199);
and U10707 (N_10707,N_10141,N_10100);
nand U10708 (N_10708,N_10292,N_10479);
and U10709 (N_10709,N_10291,N_10156);
nor U10710 (N_10710,N_10134,N_10403);
nand U10711 (N_10711,N_10361,N_10313);
nor U10712 (N_10712,N_10344,N_10342);
xnor U10713 (N_10713,N_10395,N_10394);
nand U10714 (N_10714,N_10045,N_10277);
and U10715 (N_10715,N_10350,N_10304);
nor U10716 (N_10716,N_10298,N_10287);
nand U10717 (N_10717,N_10295,N_10337);
xnor U10718 (N_10718,N_10414,N_10131);
nand U10719 (N_10719,N_10364,N_10471);
nor U10720 (N_10720,N_10447,N_10375);
xnor U10721 (N_10721,N_10246,N_10449);
nand U10722 (N_10722,N_10379,N_10336);
and U10723 (N_10723,N_10383,N_10380);
nand U10724 (N_10724,N_10462,N_10306);
nor U10725 (N_10725,N_10054,N_10084);
nand U10726 (N_10726,N_10066,N_10083);
and U10727 (N_10727,N_10293,N_10017);
or U10728 (N_10728,N_10173,N_10168);
xnor U10729 (N_10729,N_10259,N_10133);
and U10730 (N_10730,N_10029,N_10223);
and U10731 (N_10731,N_10022,N_10478);
nand U10732 (N_10732,N_10212,N_10377);
or U10733 (N_10733,N_10307,N_10217);
nand U10734 (N_10734,N_10368,N_10420);
or U10735 (N_10735,N_10354,N_10348);
and U10736 (N_10736,N_10285,N_10362);
or U10737 (N_10737,N_10171,N_10148);
nor U10738 (N_10738,N_10014,N_10353);
or U10739 (N_10739,N_10026,N_10201);
or U10740 (N_10740,N_10007,N_10090);
or U10741 (N_10741,N_10068,N_10303);
xor U10742 (N_10742,N_10013,N_10185);
nor U10743 (N_10743,N_10003,N_10366);
and U10744 (N_10744,N_10280,N_10240);
and U10745 (N_10745,N_10327,N_10255);
and U10746 (N_10746,N_10278,N_10412);
nor U10747 (N_10747,N_10119,N_10430);
xnor U10748 (N_10748,N_10035,N_10002);
nand U10749 (N_10749,N_10025,N_10356);
or U10750 (N_10750,N_10241,N_10391);
or U10751 (N_10751,N_10280,N_10387);
and U10752 (N_10752,N_10000,N_10401);
or U10753 (N_10753,N_10034,N_10079);
xor U10754 (N_10754,N_10318,N_10132);
nand U10755 (N_10755,N_10277,N_10445);
xnor U10756 (N_10756,N_10205,N_10297);
xor U10757 (N_10757,N_10278,N_10492);
nand U10758 (N_10758,N_10411,N_10323);
and U10759 (N_10759,N_10468,N_10080);
or U10760 (N_10760,N_10161,N_10038);
or U10761 (N_10761,N_10252,N_10366);
xnor U10762 (N_10762,N_10484,N_10026);
and U10763 (N_10763,N_10347,N_10132);
nand U10764 (N_10764,N_10169,N_10386);
nor U10765 (N_10765,N_10213,N_10431);
nand U10766 (N_10766,N_10433,N_10030);
nand U10767 (N_10767,N_10292,N_10362);
and U10768 (N_10768,N_10093,N_10173);
nand U10769 (N_10769,N_10225,N_10471);
or U10770 (N_10770,N_10142,N_10147);
or U10771 (N_10771,N_10318,N_10273);
and U10772 (N_10772,N_10223,N_10325);
nand U10773 (N_10773,N_10428,N_10349);
or U10774 (N_10774,N_10181,N_10253);
nand U10775 (N_10775,N_10397,N_10141);
nand U10776 (N_10776,N_10237,N_10265);
nor U10777 (N_10777,N_10077,N_10466);
xnor U10778 (N_10778,N_10385,N_10122);
and U10779 (N_10779,N_10050,N_10404);
or U10780 (N_10780,N_10297,N_10324);
nand U10781 (N_10781,N_10080,N_10130);
or U10782 (N_10782,N_10473,N_10460);
and U10783 (N_10783,N_10148,N_10143);
and U10784 (N_10784,N_10392,N_10329);
or U10785 (N_10785,N_10221,N_10048);
or U10786 (N_10786,N_10411,N_10252);
nor U10787 (N_10787,N_10387,N_10492);
and U10788 (N_10788,N_10227,N_10349);
xnor U10789 (N_10789,N_10410,N_10121);
nand U10790 (N_10790,N_10133,N_10454);
nor U10791 (N_10791,N_10233,N_10196);
xnor U10792 (N_10792,N_10386,N_10499);
or U10793 (N_10793,N_10085,N_10008);
nand U10794 (N_10794,N_10244,N_10321);
xor U10795 (N_10795,N_10272,N_10003);
and U10796 (N_10796,N_10473,N_10112);
and U10797 (N_10797,N_10273,N_10310);
xor U10798 (N_10798,N_10018,N_10257);
nor U10799 (N_10799,N_10403,N_10398);
nor U10800 (N_10800,N_10014,N_10347);
and U10801 (N_10801,N_10233,N_10032);
and U10802 (N_10802,N_10091,N_10330);
nand U10803 (N_10803,N_10070,N_10377);
nand U10804 (N_10804,N_10279,N_10404);
and U10805 (N_10805,N_10277,N_10407);
and U10806 (N_10806,N_10041,N_10113);
or U10807 (N_10807,N_10306,N_10131);
or U10808 (N_10808,N_10445,N_10212);
or U10809 (N_10809,N_10163,N_10276);
nand U10810 (N_10810,N_10185,N_10232);
and U10811 (N_10811,N_10344,N_10120);
xor U10812 (N_10812,N_10279,N_10498);
nand U10813 (N_10813,N_10216,N_10124);
xnor U10814 (N_10814,N_10077,N_10049);
nand U10815 (N_10815,N_10406,N_10121);
and U10816 (N_10816,N_10195,N_10484);
xnor U10817 (N_10817,N_10030,N_10251);
and U10818 (N_10818,N_10212,N_10297);
or U10819 (N_10819,N_10430,N_10421);
and U10820 (N_10820,N_10303,N_10207);
and U10821 (N_10821,N_10396,N_10211);
and U10822 (N_10822,N_10029,N_10095);
nand U10823 (N_10823,N_10456,N_10432);
nand U10824 (N_10824,N_10124,N_10403);
or U10825 (N_10825,N_10324,N_10475);
nand U10826 (N_10826,N_10358,N_10431);
and U10827 (N_10827,N_10260,N_10068);
xnor U10828 (N_10828,N_10112,N_10251);
and U10829 (N_10829,N_10177,N_10326);
or U10830 (N_10830,N_10428,N_10464);
nor U10831 (N_10831,N_10004,N_10017);
nand U10832 (N_10832,N_10465,N_10343);
nor U10833 (N_10833,N_10017,N_10355);
or U10834 (N_10834,N_10186,N_10146);
nand U10835 (N_10835,N_10428,N_10083);
or U10836 (N_10836,N_10192,N_10026);
and U10837 (N_10837,N_10032,N_10119);
nand U10838 (N_10838,N_10336,N_10305);
or U10839 (N_10839,N_10456,N_10213);
xor U10840 (N_10840,N_10195,N_10107);
and U10841 (N_10841,N_10433,N_10406);
nand U10842 (N_10842,N_10045,N_10251);
nand U10843 (N_10843,N_10044,N_10485);
and U10844 (N_10844,N_10262,N_10310);
nand U10845 (N_10845,N_10012,N_10152);
xnor U10846 (N_10846,N_10041,N_10278);
or U10847 (N_10847,N_10412,N_10306);
or U10848 (N_10848,N_10122,N_10400);
xor U10849 (N_10849,N_10022,N_10311);
or U10850 (N_10850,N_10147,N_10402);
or U10851 (N_10851,N_10358,N_10094);
or U10852 (N_10852,N_10351,N_10170);
xnor U10853 (N_10853,N_10490,N_10166);
or U10854 (N_10854,N_10244,N_10458);
nand U10855 (N_10855,N_10350,N_10280);
or U10856 (N_10856,N_10045,N_10477);
nand U10857 (N_10857,N_10281,N_10068);
or U10858 (N_10858,N_10163,N_10471);
or U10859 (N_10859,N_10086,N_10182);
or U10860 (N_10860,N_10282,N_10461);
nor U10861 (N_10861,N_10409,N_10112);
and U10862 (N_10862,N_10054,N_10274);
nor U10863 (N_10863,N_10148,N_10445);
and U10864 (N_10864,N_10220,N_10320);
nand U10865 (N_10865,N_10456,N_10105);
xor U10866 (N_10866,N_10330,N_10325);
xor U10867 (N_10867,N_10344,N_10484);
and U10868 (N_10868,N_10406,N_10204);
or U10869 (N_10869,N_10394,N_10134);
xor U10870 (N_10870,N_10224,N_10154);
nor U10871 (N_10871,N_10446,N_10389);
xnor U10872 (N_10872,N_10437,N_10313);
xnor U10873 (N_10873,N_10195,N_10379);
or U10874 (N_10874,N_10201,N_10368);
or U10875 (N_10875,N_10008,N_10473);
nand U10876 (N_10876,N_10069,N_10072);
nor U10877 (N_10877,N_10322,N_10195);
nand U10878 (N_10878,N_10291,N_10029);
or U10879 (N_10879,N_10413,N_10145);
nand U10880 (N_10880,N_10149,N_10412);
xnor U10881 (N_10881,N_10275,N_10392);
nor U10882 (N_10882,N_10302,N_10169);
and U10883 (N_10883,N_10416,N_10270);
xnor U10884 (N_10884,N_10235,N_10314);
nor U10885 (N_10885,N_10359,N_10486);
and U10886 (N_10886,N_10082,N_10352);
nand U10887 (N_10887,N_10084,N_10010);
and U10888 (N_10888,N_10296,N_10018);
xor U10889 (N_10889,N_10411,N_10448);
nor U10890 (N_10890,N_10005,N_10027);
nand U10891 (N_10891,N_10372,N_10427);
xnor U10892 (N_10892,N_10372,N_10277);
xnor U10893 (N_10893,N_10380,N_10488);
and U10894 (N_10894,N_10430,N_10051);
xor U10895 (N_10895,N_10459,N_10051);
nand U10896 (N_10896,N_10413,N_10221);
or U10897 (N_10897,N_10178,N_10211);
and U10898 (N_10898,N_10103,N_10047);
nor U10899 (N_10899,N_10439,N_10061);
xor U10900 (N_10900,N_10190,N_10458);
xor U10901 (N_10901,N_10427,N_10088);
nor U10902 (N_10902,N_10428,N_10046);
and U10903 (N_10903,N_10340,N_10281);
and U10904 (N_10904,N_10020,N_10194);
and U10905 (N_10905,N_10187,N_10334);
or U10906 (N_10906,N_10497,N_10116);
or U10907 (N_10907,N_10207,N_10048);
nand U10908 (N_10908,N_10093,N_10269);
or U10909 (N_10909,N_10071,N_10315);
or U10910 (N_10910,N_10133,N_10088);
nand U10911 (N_10911,N_10480,N_10251);
xor U10912 (N_10912,N_10252,N_10056);
or U10913 (N_10913,N_10382,N_10385);
nand U10914 (N_10914,N_10302,N_10207);
nand U10915 (N_10915,N_10456,N_10424);
or U10916 (N_10916,N_10421,N_10259);
nor U10917 (N_10917,N_10174,N_10108);
xor U10918 (N_10918,N_10090,N_10284);
or U10919 (N_10919,N_10157,N_10430);
nand U10920 (N_10920,N_10429,N_10463);
and U10921 (N_10921,N_10399,N_10121);
nor U10922 (N_10922,N_10414,N_10209);
and U10923 (N_10923,N_10497,N_10351);
and U10924 (N_10924,N_10164,N_10125);
or U10925 (N_10925,N_10213,N_10361);
or U10926 (N_10926,N_10424,N_10048);
nand U10927 (N_10927,N_10357,N_10193);
and U10928 (N_10928,N_10196,N_10439);
nand U10929 (N_10929,N_10203,N_10267);
nor U10930 (N_10930,N_10140,N_10378);
nand U10931 (N_10931,N_10362,N_10051);
nor U10932 (N_10932,N_10264,N_10361);
or U10933 (N_10933,N_10379,N_10057);
xnor U10934 (N_10934,N_10153,N_10170);
nand U10935 (N_10935,N_10444,N_10058);
xnor U10936 (N_10936,N_10152,N_10341);
or U10937 (N_10937,N_10141,N_10425);
nand U10938 (N_10938,N_10114,N_10049);
and U10939 (N_10939,N_10246,N_10152);
or U10940 (N_10940,N_10010,N_10082);
and U10941 (N_10941,N_10073,N_10177);
or U10942 (N_10942,N_10295,N_10417);
or U10943 (N_10943,N_10447,N_10094);
nor U10944 (N_10944,N_10445,N_10210);
and U10945 (N_10945,N_10097,N_10071);
and U10946 (N_10946,N_10171,N_10264);
xor U10947 (N_10947,N_10143,N_10018);
nand U10948 (N_10948,N_10275,N_10404);
xor U10949 (N_10949,N_10147,N_10308);
nor U10950 (N_10950,N_10354,N_10411);
nor U10951 (N_10951,N_10042,N_10295);
xnor U10952 (N_10952,N_10228,N_10428);
xor U10953 (N_10953,N_10405,N_10122);
nand U10954 (N_10954,N_10406,N_10087);
and U10955 (N_10955,N_10472,N_10375);
and U10956 (N_10956,N_10305,N_10006);
nor U10957 (N_10957,N_10115,N_10363);
and U10958 (N_10958,N_10294,N_10182);
xor U10959 (N_10959,N_10454,N_10230);
xor U10960 (N_10960,N_10043,N_10269);
nor U10961 (N_10961,N_10228,N_10414);
nand U10962 (N_10962,N_10477,N_10025);
nand U10963 (N_10963,N_10231,N_10232);
and U10964 (N_10964,N_10113,N_10496);
nand U10965 (N_10965,N_10333,N_10099);
or U10966 (N_10966,N_10403,N_10143);
nor U10967 (N_10967,N_10193,N_10201);
nor U10968 (N_10968,N_10087,N_10183);
nand U10969 (N_10969,N_10480,N_10488);
and U10970 (N_10970,N_10073,N_10484);
and U10971 (N_10971,N_10323,N_10276);
xnor U10972 (N_10972,N_10070,N_10321);
nor U10973 (N_10973,N_10463,N_10210);
nor U10974 (N_10974,N_10268,N_10224);
xnor U10975 (N_10975,N_10101,N_10081);
xor U10976 (N_10976,N_10269,N_10231);
and U10977 (N_10977,N_10095,N_10323);
or U10978 (N_10978,N_10075,N_10201);
nand U10979 (N_10979,N_10220,N_10140);
nand U10980 (N_10980,N_10096,N_10267);
xnor U10981 (N_10981,N_10347,N_10164);
xor U10982 (N_10982,N_10084,N_10183);
nor U10983 (N_10983,N_10083,N_10458);
nand U10984 (N_10984,N_10138,N_10455);
xor U10985 (N_10985,N_10459,N_10291);
or U10986 (N_10986,N_10314,N_10101);
nand U10987 (N_10987,N_10461,N_10189);
nor U10988 (N_10988,N_10456,N_10379);
and U10989 (N_10989,N_10374,N_10282);
xor U10990 (N_10990,N_10320,N_10365);
nor U10991 (N_10991,N_10358,N_10040);
xnor U10992 (N_10992,N_10465,N_10047);
nand U10993 (N_10993,N_10407,N_10462);
and U10994 (N_10994,N_10071,N_10343);
nand U10995 (N_10995,N_10109,N_10353);
nand U10996 (N_10996,N_10221,N_10070);
xor U10997 (N_10997,N_10326,N_10033);
nand U10998 (N_10998,N_10053,N_10110);
and U10999 (N_10999,N_10482,N_10139);
nand U11000 (N_11000,N_10528,N_10585);
or U11001 (N_11001,N_10930,N_10726);
xor U11002 (N_11002,N_10614,N_10977);
nor U11003 (N_11003,N_10625,N_10583);
and U11004 (N_11004,N_10667,N_10699);
nor U11005 (N_11005,N_10959,N_10693);
xnor U11006 (N_11006,N_10775,N_10786);
or U11007 (N_11007,N_10730,N_10993);
or U11008 (N_11008,N_10743,N_10516);
xnor U11009 (N_11009,N_10764,N_10579);
and U11010 (N_11010,N_10745,N_10759);
and U11011 (N_11011,N_10879,N_10575);
and U11012 (N_11012,N_10713,N_10893);
xnor U11013 (N_11013,N_10891,N_10783);
nand U11014 (N_11014,N_10750,N_10762);
nand U11015 (N_11015,N_10828,N_10763);
and U11016 (N_11016,N_10551,N_10690);
xor U11017 (N_11017,N_10607,N_10902);
nor U11018 (N_11018,N_10541,N_10578);
nand U11019 (N_11019,N_10535,N_10527);
or U11020 (N_11020,N_10935,N_10809);
or U11021 (N_11021,N_10950,N_10524);
or U11022 (N_11022,N_10905,N_10587);
or U11023 (N_11023,N_10807,N_10518);
and U11024 (N_11024,N_10938,N_10994);
nor U11025 (N_11025,N_10790,N_10644);
nand U11026 (N_11026,N_10571,N_10632);
nand U11027 (N_11027,N_10586,N_10623);
xor U11028 (N_11028,N_10920,N_10820);
and U11029 (N_11029,N_10642,N_10936);
xnor U11030 (N_11030,N_10620,N_10666);
nor U11031 (N_11031,N_10789,N_10765);
xor U11032 (N_11032,N_10982,N_10537);
xor U11033 (N_11033,N_10684,N_10749);
and U11034 (N_11034,N_10716,N_10829);
or U11035 (N_11035,N_10768,N_10856);
or U11036 (N_11036,N_10988,N_10594);
nor U11037 (N_11037,N_10530,N_10853);
and U11038 (N_11038,N_10798,N_10843);
nand U11039 (N_11039,N_10507,N_10830);
nor U11040 (N_11040,N_10539,N_10646);
xor U11041 (N_11041,N_10515,N_10990);
or U11042 (N_11042,N_10903,N_10967);
nor U11043 (N_11043,N_10796,N_10728);
nor U11044 (N_11044,N_10540,N_10593);
nand U11045 (N_11045,N_10552,N_10532);
nand U11046 (N_11046,N_10549,N_10928);
xor U11047 (N_11047,N_10673,N_10776);
nor U11048 (N_11048,N_10504,N_10640);
xor U11049 (N_11049,N_10948,N_10956);
or U11050 (N_11050,N_10940,N_10659);
xor U11051 (N_11051,N_10562,N_10556);
xnor U11052 (N_11052,N_10704,N_10616);
nand U11053 (N_11053,N_10714,N_10734);
xor U11054 (N_11054,N_10870,N_10800);
and U11055 (N_11055,N_10611,N_10894);
or U11056 (N_11056,N_10845,N_10933);
and U11057 (N_11057,N_10769,N_10958);
and U11058 (N_11058,N_10603,N_10941);
and U11059 (N_11059,N_10598,N_10580);
nand U11060 (N_11060,N_10564,N_10841);
nor U11061 (N_11061,N_10984,N_10559);
nand U11062 (N_11062,N_10808,N_10858);
nor U11063 (N_11063,N_10873,N_10817);
or U11064 (N_11064,N_10525,N_10760);
nor U11065 (N_11065,N_10857,N_10918);
or U11066 (N_11066,N_10900,N_10850);
xor U11067 (N_11067,N_10505,N_10874);
and U11068 (N_11068,N_10634,N_10823);
nor U11069 (N_11069,N_10937,N_10797);
or U11070 (N_11070,N_10927,N_10706);
and U11071 (N_11071,N_10710,N_10741);
and U11072 (N_11072,N_10631,N_10814);
and U11073 (N_11073,N_10742,N_10782);
or U11074 (N_11074,N_10919,N_10682);
and U11075 (N_11075,N_10980,N_10847);
xor U11076 (N_11076,N_10952,N_10672);
and U11077 (N_11077,N_10628,N_10998);
or U11078 (N_11078,N_10915,N_10723);
xnor U11079 (N_11079,N_10863,N_10914);
nand U11080 (N_11080,N_10793,N_10653);
xnor U11081 (N_11081,N_10944,N_10819);
xnor U11082 (N_11082,N_10751,N_10788);
xor U11083 (N_11083,N_10503,N_10971);
nor U11084 (N_11084,N_10735,N_10953);
and U11085 (N_11085,N_10691,N_10925);
nor U11086 (N_11086,N_10636,N_10983);
and U11087 (N_11087,N_10577,N_10865);
xnor U11088 (N_11088,N_10717,N_10707);
or U11089 (N_11089,N_10923,N_10754);
nand U11090 (N_11090,N_10589,N_10558);
and U11091 (N_11091,N_10621,N_10599);
and U11092 (N_11092,N_10746,N_10912);
xnor U11093 (N_11093,N_10926,N_10889);
nor U11094 (N_11094,N_10785,N_10722);
and U11095 (N_11095,N_10791,N_10637);
xnor U11096 (N_11096,N_10604,N_10834);
xnor U11097 (N_11097,N_10547,N_10802);
nor U11098 (N_11098,N_10694,N_10804);
xnor U11099 (N_11099,N_10908,N_10622);
nand U11100 (N_11100,N_10757,N_10657);
or U11101 (N_11101,N_10844,N_10934);
or U11102 (N_11102,N_10679,N_10605);
and U11103 (N_11103,N_10766,N_10668);
nand U11104 (N_11104,N_10612,N_10655);
or U11105 (N_11105,N_10981,N_10794);
and U11106 (N_11106,N_10961,N_10861);
xor U11107 (N_11107,N_10995,N_10945);
nor U11108 (N_11108,N_10999,N_10574);
and U11109 (N_11109,N_10805,N_10855);
and U11110 (N_11110,N_10572,N_10949);
xnor U11111 (N_11111,N_10985,N_10965);
or U11112 (N_11112,N_10779,N_10678);
nand U11113 (N_11113,N_10955,N_10618);
and U11114 (N_11114,N_10639,N_10600);
nand U11115 (N_11115,N_10866,N_10692);
and U11116 (N_11116,N_10840,N_10836);
nand U11117 (N_11117,N_10588,N_10546);
nand U11118 (N_11118,N_10772,N_10663);
or U11119 (N_11119,N_10748,N_10991);
xor U11120 (N_11120,N_10522,N_10851);
xor U11121 (N_11121,N_10810,N_10560);
xor U11122 (N_11122,N_10773,N_10831);
nand U11123 (N_11123,N_10881,N_10521);
and U11124 (N_11124,N_10806,N_10997);
nand U11125 (N_11125,N_10536,N_10992);
nand U11126 (N_11126,N_10633,N_10615);
and U11127 (N_11127,N_10630,N_10500);
and U11128 (N_11128,N_10904,N_10610);
and U11129 (N_11129,N_10712,N_10921);
and U11130 (N_11130,N_10709,N_10916);
and U11131 (N_11131,N_10774,N_10681);
nand U11132 (N_11132,N_10761,N_10677);
and U11133 (N_11133,N_10606,N_10570);
or U11134 (N_11134,N_10732,N_10553);
and U11135 (N_11135,N_10898,N_10601);
or U11136 (N_11136,N_10947,N_10512);
xnor U11137 (N_11137,N_10520,N_10895);
xor U11138 (N_11138,N_10647,N_10838);
nand U11139 (N_11139,N_10534,N_10839);
nor U11140 (N_11140,N_10591,N_10872);
and U11141 (N_11141,N_10877,N_10526);
xor U11142 (N_11142,N_10784,N_10543);
or U11143 (N_11143,N_10884,N_10602);
or U11144 (N_11144,N_10563,N_10654);
or U11145 (N_11145,N_10738,N_10868);
nand U11146 (N_11146,N_10922,N_10523);
or U11147 (N_11147,N_10883,N_10544);
xor U11148 (N_11148,N_10711,N_10917);
xnor U11149 (N_11149,N_10899,N_10932);
nand U11150 (N_11150,N_10687,N_10510);
nor U11151 (N_11151,N_10892,N_10701);
nand U11152 (N_11152,N_10733,N_10986);
and U11153 (N_11153,N_10860,N_10582);
and U11154 (N_11154,N_10533,N_10652);
nand U11155 (N_11155,N_10573,N_10987);
nand U11156 (N_11156,N_10826,N_10758);
and U11157 (N_11157,N_10566,N_10929);
xnor U11158 (N_11158,N_10729,N_10882);
and U11159 (N_11159,N_10705,N_10897);
and U11160 (N_11160,N_10676,N_10662);
nor U11161 (N_11161,N_10816,N_10565);
or U11162 (N_11162,N_10906,N_10799);
and U11163 (N_11163,N_10561,N_10969);
xnor U11164 (N_11164,N_10590,N_10671);
nor U11165 (N_11165,N_10939,N_10852);
and U11166 (N_11166,N_10624,N_10670);
nand U11167 (N_11167,N_10686,N_10837);
nand U11168 (N_11168,N_10548,N_10629);
and U11169 (N_11169,N_10910,N_10627);
and U11170 (N_11170,N_10951,N_10744);
xnor U11171 (N_11171,N_10660,N_10954);
xnor U11172 (N_11172,N_10645,N_10824);
nand U11173 (N_11173,N_10755,N_10978);
or U11174 (N_11174,N_10854,N_10555);
xnor U11175 (N_11175,N_10907,N_10812);
nand U11176 (N_11176,N_10825,N_10698);
or U11177 (N_11177,N_10656,N_10833);
and U11178 (N_11178,N_10752,N_10635);
xor U11179 (N_11179,N_10875,N_10513);
or U11180 (N_11180,N_10596,N_10975);
nand U11181 (N_11181,N_10508,N_10901);
nor U11182 (N_11182,N_10649,N_10996);
or U11183 (N_11183,N_10970,N_10979);
nor U11184 (N_11184,N_10962,N_10966);
and U11185 (N_11185,N_10887,N_10648);
xnor U11186 (N_11186,N_10680,N_10931);
nand U11187 (N_11187,N_10674,N_10864);
nand U11188 (N_11188,N_10724,N_10803);
xnor U11189 (N_11189,N_10664,N_10641);
xor U11190 (N_11190,N_10832,N_10911);
and U11191 (N_11191,N_10613,N_10584);
and U11192 (N_11192,N_10688,N_10675);
and U11193 (N_11193,N_10801,N_10792);
xor U11194 (N_11194,N_10683,N_10725);
and U11195 (N_11195,N_10943,N_10721);
and U11196 (N_11196,N_10545,N_10718);
or U11197 (N_11197,N_10708,N_10859);
nand U11198 (N_11198,N_10976,N_10715);
and U11199 (N_11199,N_10942,N_10538);
nor U11200 (N_11200,N_10963,N_10576);
nand U11201 (N_11201,N_10502,N_10777);
xnor U11202 (N_11202,N_10913,N_10542);
xnor U11203 (N_11203,N_10509,N_10695);
and U11204 (N_11204,N_10568,N_10795);
nor U11205 (N_11205,N_10880,N_10703);
xor U11206 (N_11206,N_10862,N_10696);
nor U11207 (N_11207,N_10946,N_10554);
nor U11208 (N_11208,N_10835,N_10960);
xnor U11209 (N_11209,N_10501,N_10909);
nor U11210 (N_11210,N_10739,N_10661);
or U11211 (N_11211,N_10506,N_10778);
and U11212 (N_11212,N_10876,N_10517);
nand U11213 (N_11213,N_10964,N_10973);
xor U11214 (N_11214,N_10731,N_10815);
or U11215 (N_11215,N_10651,N_10848);
or U11216 (N_11216,N_10719,N_10813);
xnor U11217 (N_11217,N_10753,N_10702);
nor U11218 (N_11218,N_10569,N_10867);
nor U11219 (N_11219,N_10770,N_10989);
or U11220 (N_11220,N_10972,N_10818);
nand U11221 (N_11221,N_10685,N_10780);
xnor U11222 (N_11222,N_10617,N_10638);
nand U11223 (N_11223,N_10740,N_10581);
or U11224 (N_11224,N_10519,N_10811);
xnor U11225 (N_11225,N_10821,N_10514);
xor U11226 (N_11226,N_10720,N_10869);
or U11227 (N_11227,N_10609,N_10665);
and U11228 (N_11228,N_10849,N_10595);
nand U11229 (N_11229,N_10747,N_10787);
or U11230 (N_11230,N_10531,N_10567);
and U11231 (N_11231,N_10697,N_10626);
or U11232 (N_11232,N_10885,N_10781);
and U11233 (N_11233,N_10767,N_10827);
nand U11234 (N_11234,N_10737,N_10727);
nand U11235 (N_11235,N_10890,N_10529);
nor U11236 (N_11236,N_10888,N_10550);
nor U11237 (N_11237,N_10592,N_10643);
nor U11238 (N_11238,N_10557,N_10822);
and U11239 (N_11239,N_10650,N_10771);
xnor U11240 (N_11240,N_10511,N_10924);
and U11241 (N_11241,N_10846,N_10597);
nand U11242 (N_11242,N_10886,N_10756);
and U11243 (N_11243,N_10974,N_10689);
xnor U11244 (N_11244,N_10658,N_10842);
or U11245 (N_11245,N_10608,N_10957);
or U11246 (N_11246,N_10700,N_10878);
and U11247 (N_11247,N_10871,N_10968);
xor U11248 (N_11248,N_10736,N_10896);
xor U11249 (N_11249,N_10669,N_10619);
or U11250 (N_11250,N_10605,N_10507);
and U11251 (N_11251,N_10778,N_10835);
xnor U11252 (N_11252,N_10876,N_10524);
xor U11253 (N_11253,N_10947,N_10934);
and U11254 (N_11254,N_10857,N_10637);
and U11255 (N_11255,N_10618,N_10986);
and U11256 (N_11256,N_10572,N_10899);
and U11257 (N_11257,N_10998,N_10786);
or U11258 (N_11258,N_10932,N_10964);
xnor U11259 (N_11259,N_10964,N_10718);
xnor U11260 (N_11260,N_10747,N_10702);
xnor U11261 (N_11261,N_10694,N_10568);
nand U11262 (N_11262,N_10915,N_10822);
nor U11263 (N_11263,N_10746,N_10551);
and U11264 (N_11264,N_10749,N_10562);
and U11265 (N_11265,N_10622,N_10939);
nor U11266 (N_11266,N_10882,N_10668);
nor U11267 (N_11267,N_10804,N_10875);
nor U11268 (N_11268,N_10990,N_10701);
nand U11269 (N_11269,N_10586,N_10643);
or U11270 (N_11270,N_10706,N_10757);
xor U11271 (N_11271,N_10851,N_10954);
xnor U11272 (N_11272,N_10732,N_10846);
or U11273 (N_11273,N_10721,N_10625);
nand U11274 (N_11274,N_10862,N_10893);
nand U11275 (N_11275,N_10984,N_10953);
or U11276 (N_11276,N_10772,N_10752);
xor U11277 (N_11277,N_10560,N_10505);
nand U11278 (N_11278,N_10798,N_10574);
and U11279 (N_11279,N_10538,N_10998);
and U11280 (N_11280,N_10683,N_10592);
or U11281 (N_11281,N_10558,N_10603);
nand U11282 (N_11282,N_10675,N_10588);
xnor U11283 (N_11283,N_10981,N_10879);
nor U11284 (N_11284,N_10810,N_10537);
nand U11285 (N_11285,N_10960,N_10742);
nor U11286 (N_11286,N_10809,N_10926);
nand U11287 (N_11287,N_10835,N_10567);
nor U11288 (N_11288,N_10643,N_10973);
and U11289 (N_11289,N_10763,N_10933);
and U11290 (N_11290,N_10603,N_10991);
nor U11291 (N_11291,N_10578,N_10990);
and U11292 (N_11292,N_10783,N_10930);
and U11293 (N_11293,N_10770,N_10548);
nand U11294 (N_11294,N_10650,N_10519);
nand U11295 (N_11295,N_10882,N_10617);
nand U11296 (N_11296,N_10680,N_10551);
or U11297 (N_11297,N_10698,N_10856);
xor U11298 (N_11298,N_10598,N_10517);
or U11299 (N_11299,N_10879,N_10794);
and U11300 (N_11300,N_10913,N_10848);
nor U11301 (N_11301,N_10952,N_10889);
nor U11302 (N_11302,N_10737,N_10634);
nor U11303 (N_11303,N_10631,N_10615);
xor U11304 (N_11304,N_10930,N_10953);
or U11305 (N_11305,N_10822,N_10754);
nor U11306 (N_11306,N_10560,N_10593);
nor U11307 (N_11307,N_10996,N_10803);
or U11308 (N_11308,N_10976,N_10636);
or U11309 (N_11309,N_10543,N_10985);
and U11310 (N_11310,N_10769,N_10801);
or U11311 (N_11311,N_10707,N_10822);
nor U11312 (N_11312,N_10619,N_10645);
nand U11313 (N_11313,N_10933,N_10913);
and U11314 (N_11314,N_10885,N_10592);
and U11315 (N_11315,N_10927,N_10728);
nor U11316 (N_11316,N_10834,N_10521);
and U11317 (N_11317,N_10793,N_10690);
nor U11318 (N_11318,N_10925,N_10725);
and U11319 (N_11319,N_10840,N_10721);
nand U11320 (N_11320,N_10526,N_10624);
nand U11321 (N_11321,N_10922,N_10649);
nand U11322 (N_11322,N_10697,N_10993);
xor U11323 (N_11323,N_10595,N_10653);
xnor U11324 (N_11324,N_10838,N_10784);
or U11325 (N_11325,N_10589,N_10564);
xnor U11326 (N_11326,N_10810,N_10703);
nand U11327 (N_11327,N_10897,N_10935);
or U11328 (N_11328,N_10613,N_10500);
nand U11329 (N_11329,N_10841,N_10900);
nor U11330 (N_11330,N_10754,N_10878);
or U11331 (N_11331,N_10818,N_10673);
or U11332 (N_11332,N_10585,N_10836);
or U11333 (N_11333,N_10980,N_10874);
nor U11334 (N_11334,N_10957,N_10846);
nor U11335 (N_11335,N_10820,N_10712);
nor U11336 (N_11336,N_10973,N_10929);
or U11337 (N_11337,N_10876,N_10592);
xnor U11338 (N_11338,N_10651,N_10522);
or U11339 (N_11339,N_10835,N_10703);
nor U11340 (N_11340,N_10578,N_10542);
nand U11341 (N_11341,N_10760,N_10841);
nor U11342 (N_11342,N_10733,N_10754);
or U11343 (N_11343,N_10761,N_10983);
and U11344 (N_11344,N_10579,N_10983);
and U11345 (N_11345,N_10771,N_10903);
and U11346 (N_11346,N_10952,N_10692);
or U11347 (N_11347,N_10633,N_10930);
and U11348 (N_11348,N_10802,N_10734);
and U11349 (N_11349,N_10537,N_10590);
xnor U11350 (N_11350,N_10942,N_10996);
nand U11351 (N_11351,N_10939,N_10686);
nand U11352 (N_11352,N_10732,N_10771);
nor U11353 (N_11353,N_10770,N_10668);
xor U11354 (N_11354,N_10982,N_10800);
or U11355 (N_11355,N_10911,N_10880);
and U11356 (N_11356,N_10715,N_10927);
or U11357 (N_11357,N_10527,N_10724);
nor U11358 (N_11358,N_10978,N_10806);
nand U11359 (N_11359,N_10755,N_10964);
nand U11360 (N_11360,N_10657,N_10768);
and U11361 (N_11361,N_10587,N_10881);
nand U11362 (N_11362,N_10666,N_10552);
and U11363 (N_11363,N_10877,N_10764);
or U11364 (N_11364,N_10523,N_10692);
nor U11365 (N_11365,N_10745,N_10894);
or U11366 (N_11366,N_10735,N_10575);
xnor U11367 (N_11367,N_10895,N_10630);
xnor U11368 (N_11368,N_10667,N_10937);
and U11369 (N_11369,N_10880,N_10640);
or U11370 (N_11370,N_10710,N_10774);
or U11371 (N_11371,N_10571,N_10943);
nor U11372 (N_11372,N_10770,N_10962);
xor U11373 (N_11373,N_10798,N_10989);
or U11374 (N_11374,N_10696,N_10507);
nand U11375 (N_11375,N_10570,N_10687);
xnor U11376 (N_11376,N_10686,N_10846);
nor U11377 (N_11377,N_10889,N_10865);
nand U11378 (N_11378,N_10887,N_10884);
nor U11379 (N_11379,N_10763,N_10953);
or U11380 (N_11380,N_10684,N_10907);
xnor U11381 (N_11381,N_10834,N_10629);
or U11382 (N_11382,N_10764,N_10782);
or U11383 (N_11383,N_10637,N_10558);
or U11384 (N_11384,N_10980,N_10502);
nand U11385 (N_11385,N_10885,N_10939);
or U11386 (N_11386,N_10579,N_10934);
xor U11387 (N_11387,N_10571,N_10587);
nor U11388 (N_11388,N_10802,N_10577);
or U11389 (N_11389,N_10655,N_10585);
nor U11390 (N_11390,N_10788,N_10994);
xor U11391 (N_11391,N_10959,N_10762);
nand U11392 (N_11392,N_10856,N_10753);
and U11393 (N_11393,N_10603,N_10986);
and U11394 (N_11394,N_10645,N_10715);
or U11395 (N_11395,N_10641,N_10723);
and U11396 (N_11396,N_10976,N_10640);
nand U11397 (N_11397,N_10698,N_10751);
or U11398 (N_11398,N_10823,N_10659);
nor U11399 (N_11399,N_10601,N_10683);
or U11400 (N_11400,N_10880,N_10772);
xor U11401 (N_11401,N_10619,N_10881);
or U11402 (N_11402,N_10955,N_10832);
xnor U11403 (N_11403,N_10515,N_10564);
or U11404 (N_11404,N_10523,N_10920);
or U11405 (N_11405,N_10725,N_10678);
xor U11406 (N_11406,N_10901,N_10753);
nor U11407 (N_11407,N_10647,N_10697);
nor U11408 (N_11408,N_10924,N_10521);
and U11409 (N_11409,N_10662,N_10749);
xnor U11410 (N_11410,N_10938,N_10921);
xnor U11411 (N_11411,N_10735,N_10636);
nor U11412 (N_11412,N_10521,N_10882);
or U11413 (N_11413,N_10513,N_10695);
nand U11414 (N_11414,N_10767,N_10521);
and U11415 (N_11415,N_10748,N_10696);
xnor U11416 (N_11416,N_10744,N_10953);
nor U11417 (N_11417,N_10966,N_10595);
and U11418 (N_11418,N_10892,N_10755);
or U11419 (N_11419,N_10589,N_10904);
nand U11420 (N_11420,N_10999,N_10728);
nor U11421 (N_11421,N_10555,N_10938);
or U11422 (N_11422,N_10531,N_10721);
or U11423 (N_11423,N_10536,N_10601);
or U11424 (N_11424,N_10921,N_10795);
nor U11425 (N_11425,N_10998,N_10745);
or U11426 (N_11426,N_10512,N_10685);
or U11427 (N_11427,N_10552,N_10891);
nand U11428 (N_11428,N_10741,N_10718);
and U11429 (N_11429,N_10856,N_10760);
or U11430 (N_11430,N_10774,N_10717);
nand U11431 (N_11431,N_10689,N_10688);
nor U11432 (N_11432,N_10997,N_10807);
nor U11433 (N_11433,N_10668,N_10777);
and U11434 (N_11434,N_10980,N_10786);
nand U11435 (N_11435,N_10679,N_10766);
nor U11436 (N_11436,N_10598,N_10676);
or U11437 (N_11437,N_10650,N_10837);
nor U11438 (N_11438,N_10907,N_10808);
xor U11439 (N_11439,N_10745,N_10935);
xor U11440 (N_11440,N_10573,N_10661);
xor U11441 (N_11441,N_10634,N_10540);
xnor U11442 (N_11442,N_10795,N_10787);
xnor U11443 (N_11443,N_10676,N_10901);
and U11444 (N_11444,N_10558,N_10615);
and U11445 (N_11445,N_10727,N_10924);
nand U11446 (N_11446,N_10989,N_10634);
nor U11447 (N_11447,N_10902,N_10928);
nor U11448 (N_11448,N_10852,N_10968);
nor U11449 (N_11449,N_10942,N_10919);
xnor U11450 (N_11450,N_10993,N_10658);
and U11451 (N_11451,N_10903,N_10666);
xnor U11452 (N_11452,N_10724,N_10717);
nor U11453 (N_11453,N_10869,N_10660);
or U11454 (N_11454,N_10823,N_10774);
nand U11455 (N_11455,N_10703,N_10886);
nor U11456 (N_11456,N_10620,N_10713);
and U11457 (N_11457,N_10550,N_10871);
nor U11458 (N_11458,N_10998,N_10607);
nor U11459 (N_11459,N_10991,N_10814);
xnor U11460 (N_11460,N_10844,N_10991);
xor U11461 (N_11461,N_10981,N_10855);
or U11462 (N_11462,N_10904,N_10958);
nor U11463 (N_11463,N_10886,N_10983);
and U11464 (N_11464,N_10568,N_10847);
and U11465 (N_11465,N_10983,N_10911);
xnor U11466 (N_11466,N_10901,N_10523);
or U11467 (N_11467,N_10879,N_10819);
nand U11468 (N_11468,N_10793,N_10640);
nand U11469 (N_11469,N_10673,N_10681);
or U11470 (N_11470,N_10601,N_10976);
nand U11471 (N_11471,N_10764,N_10742);
nand U11472 (N_11472,N_10749,N_10948);
and U11473 (N_11473,N_10896,N_10755);
or U11474 (N_11474,N_10680,N_10615);
or U11475 (N_11475,N_10672,N_10594);
or U11476 (N_11476,N_10856,N_10715);
or U11477 (N_11477,N_10681,N_10588);
nand U11478 (N_11478,N_10676,N_10692);
nand U11479 (N_11479,N_10741,N_10632);
and U11480 (N_11480,N_10645,N_10566);
xnor U11481 (N_11481,N_10942,N_10643);
nor U11482 (N_11482,N_10971,N_10882);
or U11483 (N_11483,N_10660,N_10826);
and U11484 (N_11484,N_10808,N_10834);
nor U11485 (N_11485,N_10682,N_10691);
nor U11486 (N_11486,N_10869,N_10893);
and U11487 (N_11487,N_10663,N_10868);
or U11488 (N_11488,N_10646,N_10590);
and U11489 (N_11489,N_10697,N_10527);
and U11490 (N_11490,N_10890,N_10536);
and U11491 (N_11491,N_10648,N_10810);
or U11492 (N_11492,N_10721,N_10540);
and U11493 (N_11493,N_10996,N_10955);
nand U11494 (N_11494,N_10870,N_10689);
nor U11495 (N_11495,N_10515,N_10625);
xnor U11496 (N_11496,N_10768,N_10759);
and U11497 (N_11497,N_10853,N_10991);
and U11498 (N_11498,N_10573,N_10552);
xnor U11499 (N_11499,N_10865,N_10930);
xnor U11500 (N_11500,N_11001,N_11288);
and U11501 (N_11501,N_11477,N_11424);
and U11502 (N_11502,N_11365,N_11071);
nand U11503 (N_11503,N_11276,N_11274);
xnor U11504 (N_11504,N_11454,N_11403);
nand U11505 (N_11505,N_11136,N_11229);
and U11506 (N_11506,N_11332,N_11449);
xor U11507 (N_11507,N_11357,N_11193);
and U11508 (N_11508,N_11455,N_11283);
nor U11509 (N_11509,N_11298,N_11101);
xor U11510 (N_11510,N_11231,N_11361);
or U11511 (N_11511,N_11255,N_11210);
xnor U11512 (N_11512,N_11351,N_11490);
or U11513 (N_11513,N_11063,N_11095);
nand U11514 (N_11514,N_11385,N_11056);
or U11515 (N_11515,N_11014,N_11368);
xnor U11516 (N_11516,N_11486,N_11147);
xnor U11517 (N_11517,N_11083,N_11328);
xor U11518 (N_11518,N_11460,N_11320);
and U11519 (N_11519,N_11119,N_11051);
nand U11520 (N_11520,N_11026,N_11059);
nand U11521 (N_11521,N_11176,N_11387);
and U11522 (N_11522,N_11090,N_11036);
nor U11523 (N_11523,N_11470,N_11240);
nand U11524 (N_11524,N_11248,N_11114);
or U11525 (N_11525,N_11463,N_11293);
or U11526 (N_11526,N_11411,N_11238);
nor U11527 (N_11527,N_11271,N_11377);
xnor U11528 (N_11528,N_11444,N_11348);
or U11529 (N_11529,N_11367,N_11372);
or U11530 (N_11530,N_11042,N_11220);
nand U11531 (N_11531,N_11419,N_11228);
or U11532 (N_11532,N_11296,N_11185);
xnor U11533 (N_11533,N_11405,N_11408);
xor U11534 (N_11534,N_11047,N_11282);
and U11535 (N_11535,N_11128,N_11010);
xnor U11536 (N_11536,N_11032,N_11187);
and U11537 (N_11537,N_11390,N_11378);
or U11538 (N_11538,N_11321,N_11339);
xor U11539 (N_11539,N_11438,N_11275);
nor U11540 (N_11540,N_11015,N_11191);
nand U11541 (N_11541,N_11386,N_11013);
nand U11542 (N_11542,N_11172,N_11107);
or U11543 (N_11543,N_11395,N_11466);
or U11544 (N_11544,N_11149,N_11195);
or U11545 (N_11545,N_11098,N_11439);
or U11546 (N_11546,N_11121,N_11201);
nand U11547 (N_11547,N_11103,N_11425);
or U11548 (N_11548,N_11144,N_11409);
xnor U11549 (N_11549,N_11197,N_11171);
or U11550 (N_11550,N_11011,N_11491);
or U11551 (N_11551,N_11402,N_11338);
nor U11552 (N_11552,N_11480,N_11140);
or U11553 (N_11553,N_11018,N_11102);
xnor U11554 (N_11554,N_11141,N_11483);
xnor U11555 (N_11555,N_11353,N_11041);
xnor U11556 (N_11556,N_11113,N_11315);
nor U11557 (N_11557,N_11007,N_11418);
or U11558 (N_11558,N_11162,N_11268);
and U11559 (N_11559,N_11199,N_11284);
nand U11560 (N_11560,N_11239,N_11091);
xor U11561 (N_11561,N_11330,N_11062);
nand U11562 (N_11562,N_11421,N_11342);
or U11563 (N_11563,N_11299,N_11226);
and U11564 (N_11564,N_11383,N_11326);
nand U11565 (N_11565,N_11325,N_11203);
xnor U11566 (N_11566,N_11314,N_11027);
and U11567 (N_11567,N_11401,N_11459);
nor U11568 (N_11568,N_11252,N_11394);
xnor U11569 (N_11569,N_11300,N_11287);
nor U11570 (N_11570,N_11082,N_11153);
nor U11571 (N_11571,N_11442,N_11078);
and U11572 (N_11572,N_11392,N_11165);
nor U11573 (N_11573,N_11108,N_11178);
nor U11574 (N_11574,N_11020,N_11498);
and U11575 (N_11575,N_11017,N_11106);
or U11576 (N_11576,N_11475,N_11242);
nor U11577 (N_11577,N_11137,N_11363);
nand U11578 (N_11578,N_11168,N_11495);
nor U11579 (N_11579,N_11125,N_11478);
and U11580 (N_11580,N_11150,N_11039);
and U11581 (N_11581,N_11012,N_11089);
xnor U11582 (N_11582,N_11190,N_11142);
nor U11583 (N_11583,N_11004,N_11318);
nor U11584 (N_11584,N_11170,N_11290);
and U11585 (N_11585,N_11343,N_11451);
or U11586 (N_11586,N_11110,N_11092);
nor U11587 (N_11587,N_11370,N_11236);
xor U11588 (N_11588,N_11474,N_11327);
or U11589 (N_11589,N_11499,N_11436);
xnor U11590 (N_11590,N_11182,N_11204);
xnor U11591 (N_11591,N_11253,N_11345);
xor U11592 (N_11592,N_11251,N_11373);
and U11593 (N_11593,N_11127,N_11235);
nor U11594 (N_11594,N_11305,N_11006);
nand U11595 (N_11595,N_11067,N_11316);
or U11596 (N_11596,N_11245,N_11008);
nor U11597 (N_11597,N_11494,N_11400);
xor U11598 (N_11598,N_11064,N_11434);
nand U11599 (N_11599,N_11329,N_11260);
xor U11600 (N_11600,N_11484,N_11181);
nor U11601 (N_11601,N_11159,N_11234);
nand U11602 (N_11602,N_11212,N_11265);
xnor U11603 (N_11603,N_11133,N_11446);
and U11604 (N_11604,N_11350,N_11324);
or U11605 (N_11605,N_11111,N_11489);
or U11606 (N_11606,N_11122,N_11105);
xor U11607 (N_11607,N_11382,N_11109);
and U11608 (N_11608,N_11087,N_11081);
nor U11609 (N_11609,N_11344,N_11280);
xor U11610 (N_11610,N_11286,N_11479);
or U11611 (N_11611,N_11038,N_11346);
nor U11612 (N_11612,N_11323,N_11319);
nor U11613 (N_11613,N_11033,N_11227);
nor U11614 (N_11614,N_11048,N_11224);
nand U11615 (N_11615,N_11311,N_11313);
and U11616 (N_11616,N_11154,N_11115);
nand U11617 (N_11617,N_11233,N_11487);
or U11618 (N_11618,N_11453,N_11369);
xor U11619 (N_11619,N_11295,N_11429);
nor U11620 (N_11620,N_11029,N_11285);
nand U11621 (N_11621,N_11093,N_11347);
xor U11622 (N_11622,N_11473,N_11232);
nand U11623 (N_11623,N_11189,N_11497);
and U11624 (N_11624,N_11132,N_11481);
and U11625 (N_11625,N_11023,N_11075);
xnor U11626 (N_11626,N_11270,N_11471);
nand U11627 (N_11627,N_11356,N_11289);
xnor U11628 (N_11628,N_11221,N_11374);
and U11629 (N_11629,N_11393,N_11021);
or U11630 (N_11630,N_11179,N_11217);
nor U11631 (N_11631,N_11052,N_11423);
nor U11632 (N_11632,N_11492,N_11244);
nor U11633 (N_11633,N_11375,N_11143);
xnor U11634 (N_11634,N_11123,N_11246);
nor U11635 (N_11635,N_11138,N_11045);
nor U11636 (N_11636,N_11493,N_11292);
or U11637 (N_11637,N_11126,N_11073);
and U11638 (N_11638,N_11404,N_11218);
and U11639 (N_11639,N_11198,N_11397);
and U11640 (N_11640,N_11371,N_11219);
and U11641 (N_11641,N_11044,N_11389);
xor U11642 (N_11642,N_11037,N_11183);
nand U11643 (N_11643,N_11333,N_11146);
xor U11644 (N_11644,N_11476,N_11254);
or U11645 (N_11645,N_11175,N_11452);
or U11646 (N_11646,N_11396,N_11427);
nor U11647 (N_11647,N_11448,N_11349);
or U11648 (N_11648,N_11428,N_11065);
or U11649 (N_11649,N_11117,N_11272);
xnor U11650 (N_11650,N_11049,N_11202);
or U11651 (N_11651,N_11118,N_11264);
and U11652 (N_11652,N_11364,N_11031);
or U11653 (N_11653,N_11024,N_11307);
xnor U11654 (N_11654,N_11208,N_11009);
xnor U11655 (N_11655,N_11261,N_11173);
and U11656 (N_11656,N_11359,N_11407);
xnor U11657 (N_11657,N_11310,N_11070);
nor U11658 (N_11658,N_11099,N_11080);
and U11659 (N_11659,N_11104,N_11053);
or U11660 (N_11660,N_11291,N_11100);
or U11661 (N_11661,N_11069,N_11222);
nand U11662 (N_11662,N_11209,N_11376);
nor U11663 (N_11663,N_11417,N_11112);
nor U11664 (N_11664,N_11464,N_11277);
and U11665 (N_11665,N_11163,N_11458);
nor U11666 (N_11666,N_11462,N_11243);
or U11667 (N_11667,N_11269,N_11158);
nand U11668 (N_11668,N_11360,N_11258);
nand U11669 (N_11669,N_11177,N_11225);
and U11670 (N_11670,N_11304,N_11312);
or U11671 (N_11671,N_11211,N_11336);
and U11672 (N_11672,N_11482,N_11076);
nand U11673 (N_11673,N_11040,N_11431);
nor U11674 (N_11674,N_11384,N_11461);
and U11675 (N_11675,N_11335,N_11030);
or U11676 (N_11676,N_11050,N_11362);
nor U11677 (N_11677,N_11447,N_11379);
xor U11678 (N_11678,N_11263,N_11194);
or U11679 (N_11679,N_11381,N_11437);
nor U11680 (N_11680,N_11161,N_11456);
and U11681 (N_11681,N_11022,N_11034);
or U11682 (N_11682,N_11160,N_11278);
xnor U11683 (N_11683,N_11096,N_11388);
nor U11684 (N_11684,N_11317,N_11398);
nand U11685 (N_11685,N_11213,N_11035);
and U11686 (N_11686,N_11139,N_11309);
nor U11687 (N_11687,N_11188,N_11457);
and U11688 (N_11688,N_11416,N_11019);
xnor U11689 (N_11689,N_11061,N_11167);
and U11690 (N_11690,N_11028,N_11354);
or U11691 (N_11691,N_11145,N_11247);
xnor U11692 (N_11692,N_11430,N_11174);
and U11693 (N_11693,N_11303,N_11422);
xnor U11694 (N_11694,N_11441,N_11334);
xor U11695 (N_11695,N_11249,N_11124);
nor U11696 (N_11696,N_11426,N_11155);
or U11697 (N_11697,N_11433,N_11164);
nand U11698 (N_11698,N_11206,N_11000);
nor U11699 (N_11699,N_11223,N_11281);
nand U11700 (N_11700,N_11025,N_11072);
and U11701 (N_11701,N_11169,N_11337);
nand U11702 (N_11702,N_11131,N_11079);
or U11703 (N_11703,N_11432,N_11440);
and U11704 (N_11704,N_11465,N_11306);
nand U11705 (N_11705,N_11380,N_11086);
and U11706 (N_11706,N_11266,N_11420);
xor U11707 (N_11707,N_11273,N_11472);
and U11708 (N_11708,N_11331,N_11412);
nor U11709 (N_11709,N_11066,N_11443);
nand U11710 (N_11710,N_11406,N_11414);
nor U11711 (N_11711,N_11267,N_11468);
nand U11712 (N_11712,N_11060,N_11279);
xnor U11713 (N_11713,N_11186,N_11074);
nand U11714 (N_11714,N_11413,N_11120);
xnor U11715 (N_11715,N_11077,N_11415);
or U11716 (N_11716,N_11341,N_11205);
nor U11717 (N_11717,N_11485,N_11301);
or U11718 (N_11718,N_11046,N_11322);
nor U11719 (N_11719,N_11085,N_11184);
nand U11720 (N_11720,N_11157,N_11302);
or U11721 (N_11721,N_11496,N_11399);
nand U11722 (N_11722,N_11084,N_11241);
and U11723 (N_11723,N_11488,N_11002);
or U11724 (N_11724,N_11097,N_11294);
nand U11725 (N_11725,N_11237,N_11391);
or U11726 (N_11726,N_11215,N_11148);
xnor U11727 (N_11727,N_11057,N_11308);
nand U11728 (N_11728,N_11088,N_11467);
xnor U11729 (N_11729,N_11340,N_11216);
nor U11730 (N_11730,N_11192,N_11166);
nor U11731 (N_11731,N_11003,N_11410);
nand U11732 (N_11732,N_11445,N_11358);
nor U11733 (N_11733,N_11016,N_11156);
nand U11734 (N_11734,N_11043,N_11151);
and U11735 (N_11735,N_11180,N_11435);
xor U11736 (N_11736,N_11116,N_11256);
or U11737 (N_11737,N_11297,N_11469);
or U11738 (N_11738,N_11055,N_11355);
xnor U11739 (N_11739,N_11058,N_11054);
nor U11740 (N_11740,N_11196,N_11207);
nand U11741 (N_11741,N_11257,N_11130);
and U11742 (N_11742,N_11094,N_11134);
nor U11743 (N_11743,N_11450,N_11262);
and U11744 (N_11744,N_11129,N_11152);
and U11745 (N_11745,N_11135,N_11200);
or U11746 (N_11746,N_11214,N_11230);
nor U11747 (N_11747,N_11005,N_11352);
nor U11748 (N_11748,N_11250,N_11259);
and U11749 (N_11749,N_11068,N_11366);
nor U11750 (N_11750,N_11174,N_11026);
nand U11751 (N_11751,N_11183,N_11306);
nor U11752 (N_11752,N_11487,N_11071);
or U11753 (N_11753,N_11416,N_11029);
nand U11754 (N_11754,N_11486,N_11490);
or U11755 (N_11755,N_11402,N_11016);
nand U11756 (N_11756,N_11328,N_11299);
and U11757 (N_11757,N_11096,N_11470);
xor U11758 (N_11758,N_11136,N_11401);
nor U11759 (N_11759,N_11312,N_11400);
and U11760 (N_11760,N_11071,N_11083);
and U11761 (N_11761,N_11125,N_11362);
nand U11762 (N_11762,N_11132,N_11303);
or U11763 (N_11763,N_11137,N_11288);
xor U11764 (N_11764,N_11249,N_11271);
xor U11765 (N_11765,N_11089,N_11312);
and U11766 (N_11766,N_11341,N_11497);
nand U11767 (N_11767,N_11293,N_11381);
nand U11768 (N_11768,N_11040,N_11398);
or U11769 (N_11769,N_11061,N_11301);
nor U11770 (N_11770,N_11103,N_11343);
or U11771 (N_11771,N_11278,N_11287);
and U11772 (N_11772,N_11145,N_11281);
xnor U11773 (N_11773,N_11445,N_11239);
or U11774 (N_11774,N_11223,N_11014);
and U11775 (N_11775,N_11073,N_11422);
or U11776 (N_11776,N_11037,N_11234);
and U11777 (N_11777,N_11128,N_11214);
nand U11778 (N_11778,N_11211,N_11108);
xnor U11779 (N_11779,N_11425,N_11040);
nor U11780 (N_11780,N_11245,N_11388);
xnor U11781 (N_11781,N_11330,N_11179);
nand U11782 (N_11782,N_11261,N_11283);
nand U11783 (N_11783,N_11112,N_11371);
nand U11784 (N_11784,N_11452,N_11135);
nor U11785 (N_11785,N_11014,N_11397);
nand U11786 (N_11786,N_11408,N_11107);
nor U11787 (N_11787,N_11419,N_11023);
and U11788 (N_11788,N_11008,N_11494);
and U11789 (N_11789,N_11485,N_11344);
or U11790 (N_11790,N_11442,N_11297);
or U11791 (N_11791,N_11267,N_11304);
nor U11792 (N_11792,N_11023,N_11072);
nor U11793 (N_11793,N_11410,N_11377);
nand U11794 (N_11794,N_11422,N_11389);
nor U11795 (N_11795,N_11308,N_11424);
and U11796 (N_11796,N_11157,N_11392);
or U11797 (N_11797,N_11457,N_11311);
xor U11798 (N_11798,N_11168,N_11346);
xnor U11799 (N_11799,N_11444,N_11295);
or U11800 (N_11800,N_11092,N_11087);
nand U11801 (N_11801,N_11376,N_11473);
nor U11802 (N_11802,N_11066,N_11309);
nor U11803 (N_11803,N_11496,N_11120);
and U11804 (N_11804,N_11329,N_11124);
nand U11805 (N_11805,N_11418,N_11362);
nand U11806 (N_11806,N_11423,N_11258);
and U11807 (N_11807,N_11089,N_11355);
or U11808 (N_11808,N_11497,N_11137);
xnor U11809 (N_11809,N_11079,N_11416);
or U11810 (N_11810,N_11007,N_11397);
xnor U11811 (N_11811,N_11134,N_11449);
or U11812 (N_11812,N_11274,N_11323);
nor U11813 (N_11813,N_11113,N_11415);
and U11814 (N_11814,N_11375,N_11117);
and U11815 (N_11815,N_11496,N_11412);
or U11816 (N_11816,N_11285,N_11472);
xor U11817 (N_11817,N_11438,N_11053);
nand U11818 (N_11818,N_11265,N_11295);
or U11819 (N_11819,N_11411,N_11216);
nor U11820 (N_11820,N_11371,N_11318);
or U11821 (N_11821,N_11435,N_11118);
or U11822 (N_11822,N_11347,N_11126);
nand U11823 (N_11823,N_11173,N_11123);
xor U11824 (N_11824,N_11217,N_11017);
nor U11825 (N_11825,N_11463,N_11426);
or U11826 (N_11826,N_11472,N_11038);
or U11827 (N_11827,N_11083,N_11183);
or U11828 (N_11828,N_11376,N_11407);
xor U11829 (N_11829,N_11266,N_11192);
nand U11830 (N_11830,N_11023,N_11298);
and U11831 (N_11831,N_11143,N_11429);
nand U11832 (N_11832,N_11005,N_11453);
and U11833 (N_11833,N_11166,N_11220);
or U11834 (N_11834,N_11490,N_11109);
nand U11835 (N_11835,N_11487,N_11428);
xnor U11836 (N_11836,N_11304,N_11023);
nand U11837 (N_11837,N_11044,N_11476);
or U11838 (N_11838,N_11449,N_11169);
nand U11839 (N_11839,N_11089,N_11493);
xor U11840 (N_11840,N_11246,N_11420);
nor U11841 (N_11841,N_11151,N_11238);
nor U11842 (N_11842,N_11037,N_11355);
nand U11843 (N_11843,N_11466,N_11438);
nor U11844 (N_11844,N_11282,N_11002);
or U11845 (N_11845,N_11114,N_11383);
nor U11846 (N_11846,N_11097,N_11255);
nor U11847 (N_11847,N_11224,N_11171);
and U11848 (N_11848,N_11278,N_11162);
or U11849 (N_11849,N_11097,N_11009);
nor U11850 (N_11850,N_11380,N_11400);
xor U11851 (N_11851,N_11474,N_11344);
or U11852 (N_11852,N_11223,N_11318);
nor U11853 (N_11853,N_11365,N_11277);
xor U11854 (N_11854,N_11065,N_11445);
nor U11855 (N_11855,N_11408,N_11201);
and U11856 (N_11856,N_11288,N_11197);
xnor U11857 (N_11857,N_11359,N_11290);
and U11858 (N_11858,N_11087,N_11252);
nor U11859 (N_11859,N_11007,N_11124);
or U11860 (N_11860,N_11494,N_11169);
or U11861 (N_11861,N_11233,N_11438);
and U11862 (N_11862,N_11065,N_11150);
nor U11863 (N_11863,N_11457,N_11279);
nand U11864 (N_11864,N_11437,N_11339);
or U11865 (N_11865,N_11176,N_11057);
nor U11866 (N_11866,N_11387,N_11043);
nor U11867 (N_11867,N_11239,N_11298);
nand U11868 (N_11868,N_11246,N_11105);
xor U11869 (N_11869,N_11456,N_11471);
nor U11870 (N_11870,N_11423,N_11032);
nor U11871 (N_11871,N_11188,N_11179);
and U11872 (N_11872,N_11194,N_11362);
nand U11873 (N_11873,N_11053,N_11071);
nor U11874 (N_11874,N_11379,N_11086);
or U11875 (N_11875,N_11103,N_11474);
or U11876 (N_11876,N_11165,N_11237);
nor U11877 (N_11877,N_11335,N_11139);
and U11878 (N_11878,N_11305,N_11442);
nor U11879 (N_11879,N_11374,N_11174);
or U11880 (N_11880,N_11142,N_11085);
xnor U11881 (N_11881,N_11310,N_11493);
xor U11882 (N_11882,N_11049,N_11228);
xor U11883 (N_11883,N_11053,N_11036);
and U11884 (N_11884,N_11036,N_11466);
or U11885 (N_11885,N_11354,N_11301);
or U11886 (N_11886,N_11153,N_11418);
nand U11887 (N_11887,N_11341,N_11036);
nand U11888 (N_11888,N_11400,N_11191);
xor U11889 (N_11889,N_11070,N_11286);
or U11890 (N_11890,N_11415,N_11424);
and U11891 (N_11891,N_11368,N_11026);
nand U11892 (N_11892,N_11162,N_11109);
xnor U11893 (N_11893,N_11280,N_11056);
and U11894 (N_11894,N_11434,N_11298);
nand U11895 (N_11895,N_11476,N_11366);
nand U11896 (N_11896,N_11392,N_11021);
and U11897 (N_11897,N_11310,N_11043);
or U11898 (N_11898,N_11249,N_11462);
xor U11899 (N_11899,N_11088,N_11251);
and U11900 (N_11900,N_11160,N_11019);
xor U11901 (N_11901,N_11333,N_11277);
and U11902 (N_11902,N_11335,N_11360);
or U11903 (N_11903,N_11238,N_11356);
or U11904 (N_11904,N_11091,N_11260);
and U11905 (N_11905,N_11496,N_11264);
and U11906 (N_11906,N_11305,N_11206);
or U11907 (N_11907,N_11332,N_11256);
nand U11908 (N_11908,N_11130,N_11189);
nor U11909 (N_11909,N_11017,N_11114);
nand U11910 (N_11910,N_11301,N_11399);
and U11911 (N_11911,N_11141,N_11025);
xor U11912 (N_11912,N_11478,N_11318);
nand U11913 (N_11913,N_11386,N_11023);
nand U11914 (N_11914,N_11128,N_11057);
and U11915 (N_11915,N_11225,N_11321);
xor U11916 (N_11916,N_11275,N_11258);
and U11917 (N_11917,N_11326,N_11402);
or U11918 (N_11918,N_11436,N_11082);
nand U11919 (N_11919,N_11042,N_11126);
and U11920 (N_11920,N_11108,N_11498);
and U11921 (N_11921,N_11315,N_11267);
xnor U11922 (N_11922,N_11368,N_11113);
nor U11923 (N_11923,N_11230,N_11395);
xor U11924 (N_11924,N_11176,N_11076);
and U11925 (N_11925,N_11228,N_11207);
nor U11926 (N_11926,N_11411,N_11009);
nand U11927 (N_11927,N_11461,N_11365);
and U11928 (N_11928,N_11179,N_11106);
nor U11929 (N_11929,N_11120,N_11444);
xnor U11930 (N_11930,N_11459,N_11049);
and U11931 (N_11931,N_11193,N_11109);
and U11932 (N_11932,N_11219,N_11186);
xor U11933 (N_11933,N_11284,N_11499);
nor U11934 (N_11934,N_11422,N_11008);
nor U11935 (N_11935,N_11144,N_11380);
nand U11936 (N_11936,N_11264,N_11013);
nor U11937 (N_11937,N_11099,N_11139);
xor U11938 (N_11938,N_11303,N_11202);
nand U11939 (N_11939,N_11334,N_11349);
xor U11940 (N_11940,N_11175,N_11075);
nand U11941 (N_11941,N_11095,N_11256);
or U11942 (N_11942,N_11162,N_11375);
nand U11943 (N_11943,N_11388,N_11068);
nand U11944 (N_11944,N_11491,N_11277);
nor U11945 (N_11945,N_11445,N_11208);
xnor U11946 (N_11946,N_11339,N_11202);
and U11947 (N_11947,N_11074,N_11035);
and U11948 (N_11948,N_11176,N_11106);
nand U11949 (N_11949,N_11427,N_11178);
and U11950 (N_11950,N_11263,N_11289);
nand U11951 (N_11951,N_11471,N_11149);
xnor U11952 (N_11952,N_11183,N_11049);
xor U11953 (N_11953,N_11447,N_11046);
nor U11954 (N_11954,N_11322,N_11011);
nor U11955 (N_11955,N_11484,N_11167);
xor U11956 (N_11956,N_11485,N_11103);
xnor U11957 (N_11957,N_11228,N_11100);
or U11958 (N_11958,N_11368,N_11446);
and U11959 (N_11959,N_11359,N_11360);
and U11960 (N_11960,N_11317,N_11196);
and U11961 (N_11961,N_11336,N_11026);
xnor U11962 (N_11962,N_11187,N_11483);
xnor U11963 (N_11963,N_11084,N_11382);
and U11964 (N_11964,N_11044,N_11370);
or U11965 (N_11965,N_11090,N_11475);
or U11966 (N_11966,N_11202,N_11361);
nor U11967 (N_11967,N_11434,N_11363);
xnor U11968 (N_11968,N_11197,N_11349);
nor U11969 (N_11969,N_11216,N_11237);
or U11970 (N_11970,N_11316,N_11174);
nor U11971 (N_11971,N_11471,N_11231);
nor U11972 (N_11972,N_11468,N_11454);
or U11973 (N_11973,N_11087,N_11117);
nand U11974 (N_11974,N_11380,N_11053);
and U11975 (N_11975,N_11381,N_11422);
nor U11976 (N_11976,N_11176,N_11109);
nor U11977 (N_11977,N_11007,N_11380);
nand U11978 (N_11978,N_11395,N_11197);
and U11979 (N_11979,N_11075,N_11072);
or U11980 (N_11980,N_11056,N_11156);
and U11981 (N_11981,N_11437,N_11266);
and U11982 (N_11982,N_11349,N_11061);
and U11983 (N_11983,N_11060,N_11368);
and U11984 (N_11984,N_11002,N_11011);
nor U11985 (N_11985,N_11088,N_11469);
nor U11986 (N_11986,N_11482,N_11364);
nand U11987 (N_11987,N_11015,N_11078);
xor U11988 (N_11988,N_11342,N_11250);
xnor U11989 (N_11989,N_11160,N_11022);
and U11990 (N_11990,N_11221,N_11187);
or U11991 (N_11991,N_11109,N_11303);
xor U11992 (N_11992,N_11227,N_11383);
or U11993 (N_11993,N_11177,N_11152);
or U11994 (N_11994,N_11458,N_11314);
and U11995 (N_11995,N_11128,N_11262);
and U11996 (N_11996,N_11383,N_11107);
and U11997 (N_11997,N_11154,N_11293);
and U11998 (N_11998,N_11339,N_11132);
and U11999 (N_11999,N_11133,N_11250);
xor U12000 (N_12000,N_11504,N_11583);
xor U12001 (N_12001,N_11888,N_11813);
and U12002 (N_12002,N_11856,N_11996);
nor U12003 (N_12003,N_11749,N_11681);
nor U12004 (N_12004,N_11928,N_11848);
nor U12005 (N_12005,N_11724,N_11574);
xor U12006 (N_12006,N_11839,N_11559);
and U12007 (N_12007,N_11897,N_11834);
nor U12008 (N_12008,N_11604,N_11692);
nor U12009 (N_12009,N_11793,N_11977);
or U12010 (N_12010,N_11893,N_11846);
nand U12011 (N_12011,N_11614,N_11657);
nor U12012 (N_12012,N_11830,N_11648);
and U12013 (N_12013,N_11968,N_11932);
xnor U12014 (N_12014,N_11627,N_11655);
xnor U12015 (N_12015,N_11649,N_11855);
and U12016 (N_12016,N_11898,N_11904);
and U12017 (N_12017,N_11506,N_11701);
or U12018 (N_12018,N_11779,N_11538);
and U12019 (N_12019,N_11659,N_11700);
and U12020 (N_12020,N_11915,N_11640);
and U12021 (N_12021,N_11948,N_11656);
or U12022 (N_12022,N_11611,N_11533);
or U12023 (N_12023,N_11597,N_11573);
nor U12024 (N_12024,N_11929,N_11894);
xor U12025 (N_12025,N_11757,N_11868);
nor U12026 (N_12026,N_11952,N_11716);
and U12027 (N_12027,N_11866,N_11963);
and U12028 (N_12028,N_11748,N_11861);
xor U12029 (N_12029,N_11661,N_11828);
xnor U12030 (N_12030,N_11651,N_11989);
xnor U12031 (N_12031,N_11671,N_11742);
or U12032 (N_12032,N_11763,N_11688);
nand U12033 (N_12033,N_11557,N_11726);
xnor U12034 (N_12034,N_11721,N_11605);
nand U12035 (N_12035,N_11728,N_11523);
xnor U12036 (N_12036,N_11809,N_11775);
or U12037 (N_12037,N_11542,N_11590);
or U12038 (N_12038,N_11550,N_11566);
and U12039 (N_12039,N_11630,N_11667);
xnor U12040 (N_12040,N_11707,N_11907);
xor U12041 (N_12041,N_11632,N_11927);
nor U12042 (N_12042,N_11791,N_11825);
or U12043 (N_12043,N_11801,N_11954);
or U12044 (N_12044,N_11680,N_11704);
nand U12045 (N_12045,N_11911,N_11575);
nor U12046 (N_12046,N_11754,N_11781);
and U12047 (N_12047,N_11608,N_11685);
nand U12048 (N_12048,N_11979,N_11703);
and U12049 (N_12049,N_11556,N_11511);
or U12050 (N_12050,N_11658,N_11978);
or U12051 (N_12051,N_11746,N_11755);
or U12052 (N_12052,N_11699,N_11788);
or U12053 (N_12053,N_11878,N_11772);
and U12054 (N_12054,N_11870,N_11546);
nand U12055 (N_12055,N_11509,N_11578);
and U12056 (N_12056,N_11949,N_11529);
and U12057 (N_12057,N_11924,N_11872);
nor U12058 (N_12058,N_11747,N_11956);
nand U12059 (N_12059,N_11545,N_11994);
xor U12060 (N_12060,N_11946,N_11923);
or U12061 (N_12061,N_11774,N_11508);
nor U12062 (N_12062,N_11899,N_11702);
nand U12063 (N_12063,N_11633,N_11690);
xor U12064 (N_12064,N_11715,N_11739);
nor U12065 (N_12065,N_11891,N_11693);
xnor U12066 (N_12066,N_11816,N_11879);
nor U12067 (N_12067,N_11618,N_11803);
xnor U12068 (N_12068,N_11760,N_11769);
xor U12069 (N_12069,N_11615,N_11564);
nand U12070 (N_12070,N_11887,N_11727);
and U12071 (N_12071,N_11500,N_11600);
and U12072 (N_12072,N_11764,N_11524);
and U12073 (N_12073,N_11964,N_11877);
nand U12074 (N_12074,N_11598,N_11939);
and U12075 (N_12075,N_11859,N_11507);
nand U12076 (N_12076,N_11531,N_11718);
or U12077 (N_12077,N_11806,N_11503);
xor U12078 (N_12078,N_11517,N_11944);
nand U12079 (N_12079,N_11722,N_11595);
nand U12080 (N_12080,N_11672,N_11743);
nand U12081 (N_12081,N_11885,N_11822);
or U12082 (N_12082,N_11596,N_11565);
nor U12083 (N_12083,N_11577,N_11636);
nor U12084 (N_12084,N_11663,N_11833);
nor U12085 (N_12085,N_11841,N_11543);
or U12086 (N_12086,N_11960,N_11937);
nor U12087 (N_12087,N_11972,N_11621);
and U12088 (N_12088,N_11799,N_11850);
nor U12089 (N_12089,N_11892,N_11555);
or U12090 (N_12090,N_11991,N_11941);
and U12091 (N_12091,N_11647,N_11761);
nor U12092 (N_12092,N_11992,N_11539);
and U12093 (N_12093,N_11646,N_11852);
nor U12094 (N_12094,N_11936,N_11567);
nor U12095 (N_12095,N_11687,N_11705);
or U12096 (N_12096,N_11515,N_11957);
nand U12097 (N_12097,N_11725,N_11925);
or U12098 (N_12098,N_11862,N_11522);
and U12099 (N_12099,N_11969,N_11798);
and U12100 (N_12100,N_11625,N_11778);
nor U12101 (N_12101,N_11712,N_11934);
and U12102 (N_12102,N_11942,N_11631);
and U12103 (N_12103,N_11562,N_11812);
or U12104 (N_12104,N_11909,N_11512);
xnor U12105 (N_12105,N_11532,N_11931);
nand U12106 (N_12106,N_11759,N_11623);
and U12107 (N_12107,N_11820,N_11734);
xor U12108 (N_12108,N_11860,N_11970);
and U12109 (N_12109,N_11612,N_11794);
or U12110 (N_12110,N_11973,N_11917);
nand U12111 (N_12111,N_11738,N_11582);
nand U12112 (N_12112,N_11854,N_11635);
and U12113 (N_12113,N_11766,N_11980);
xnor U12114 (N_12114,N_11518,N_11995);
xnor U12115 (N_12115,N_11851,N_11535);
and U12116 (N_12116,N_11650,N_11731);
and U12117 (N_12117,N_11634,N_11609);
and U12118 (N_12118,N_11843,N_11768);
and U12119 (N_12119,N_11818,N_11686);
nand U12120 (N_12120,N_11638,N_11570);
or U12121 (N_12121,N_11717,N_11584);
xor U12122 (N_12122,N_11714,N_11784);
or U12123 (N_12123,N_11514,N_11758);
or U12124 (N_12124,N_11698,N_11984);
xnor U12125 (N_12125,N_11875,N_11720);
nor U12126 (N_12126,N_11881,N_11594);
or U12127 (N_12127,N_11771,N_11913);
xnor U12128 (N_12128,N_11643,N_11876);
xor U12129 (N_12129,N_11628,N_11900);
and U12130 (N_12130,N_11938,N_11677);
nand U12131 (N_12131,N_11541,N_11551);
and U12132 (N_12132,N_11607,N_11958);
and U12133 (N_12133,N_11780,N_11886);
xnor U12134 (N_12134,N_11997,N_11800);
nor U12135 (N_12135,N_11817,N_11889);
and U12136 (N_12136,N_11732,N_11619);
nor U12137 (N_12137,N_11563,N_11940);
nand U12138 (N_12138,N_11521,N_11639);
or U12139 (N_12139,N_11926,N_11988);
nand U12140 (N_12140,N_11593,N_11976);
nand U12141 (N_12141,N_11914,N_11827);
nand U12142 (N_12142,N_11697,N_11883);
xor U12143 (N_12143,N_11815,N_11767);
xnor U12144 (N_12144,N_11975,N_11537);
nor U12145 (N_12145,N_11986,N_11528);
nand U12146 (N_12146,N_11987,N_11581);
and U12147 (N_12147,N_11708,N_11867);
or U12148 (N_12148,N_11829,N_11795);
nand U12149 (N_12149,N_11982,N_11603);
and U12150 (N_12150,N_11840,N_11930);
or U12151 (N_12151,N_11790,N_11560);
xor U12152 (N_12152,N_11525,N_11985);
xor U12153 (N_12153,N_11579,N_11933);
or U12154 (N_12154,N_11906,N_11510);
and U12155 (N_12155,N_11955,N_11971);
nand U12156 (N_12156,N_11540,N_11552);
nand U12157 (N_12157,N_11673,N_11804);
and U12158 (N_12158,N_11787,N_11601);
xor U12159 (N_12159,N_11990,N_11961);
or U12160 (N_12160,N_11950,N_11873);
and U12161 (N_12161,N_11620,N_11536);
and U12162 (N_12162,N_11684,N_11824);
xnor U12163 (N_12163,N_11910,N_11967);
and U12164 (N_12164,N_11864,N_11918);
or U12165 (N_12165,N_11805,N_11723);
nor U12166 (N_12166,N_11641,N_11905);
and U12167 (N_12167,N_11849,N_11965);
and U12168 (N_12168,N_11586,N_11665);
nand U12169 (N_12169,N_11808,N_11762);
or U12170 (N_12170,N_11660,N_11580);
xor U12171 (N_12171,N_11902,N_11674);
or U12172 (N_12172,N_11526,N_11617);
nor U12173 (N_12173,N_11951,N_11544);
and U12174 (N_12174,N_11576,N_11519);
nor U12175 (N_12175,N_11777,N_11896);
or U12176 (N_12176,N_11880,N_11884);
nor U12177 (N_12177,N_11821,N_11842);
or U12178 (N_12178,N_11783,N_11653);
nand U12179 (N_12179,N_11682,N_11568);
nor U12180 (N_12180,N_11935,N_11502);
xnor U12181 (N_12181,N_11706,N_11895);
nor U12182 (N_12182,N_11890,N_11814);
nor U12183 (N_12183,N_11826,N_11610);
nand U12184 (N_12184,N_11752,N_11776);
nor U12185 (N_12185,N_11669,N_11652);
and U12186 (N_12186,N_11737,N_11616);
and U12187 (N_12187,N_11865,N_11750);
xnor U12188 (N_12188,N_11505,N_11516);
or U12189 (N_12189,N_11863,N_11844);
nor U12190 (N_12190,N_11689,N_11624);
nand U12191 (N_12191,N_11554,N_11945);
nor U12192 (N_12192,N_11530,N_11974);
nand U12193 (N_12193,N_11810,N_11901);
nor U12194 (N_12194,N_11709,N_11733);
or U12195 (N_12195,N_11959,N_11785);
nand U12196 (N_12196,N_11558,N_11588);
nand U12197 (N_12197,N_11741,N_11591);
xor U12198 (N_12198,N_11819,N_11548);
xnor U12199 (N_12199,N_11694,N_11999);
or U12200 (N_12200,N_11679,N_11920);
nand U12201 (N_12201,N_11683,N_11908);
and U12202 (N_12202,N_11912,N_11592);
or U12203 (N_12203,N_11549,N_11802);
and U12204 (N_12204,N_11606,N_11943);
and U12205 (N_12205,N_11637,N_11642);
or U12206 (N_12206,N_11613,N_11947);
and U12207 (N_12207,N_11773,N_11501);
nor U12208 (N_12208,N_11644,N_11666);
and U12209 (N_12209,N_11730,N_11670);
or U12210 (N_12210,N_11869,N_11792);
nor U12211 (N_12211,N_11664,N_11599);
and U12212 (N_12212,N_11962,N_11527);
nor U12213 (N_12213,N_11654,N_11691);
nor U12214 (N_12214,N_11711,N_11903);
nand U12215 (N_12215,N_11589,N_11857);
and U12216 (N_12216,N_11729,N_11534);
nand U12217 (N_12217,N_11547,N_11837);
xnor U12218 (N_12218,N_11753,N_11953);
and U12219 (N_12219,N_11585,N_11838);
nand U12220 (N_12220,N_11858,N_11983);
xnor U12221 (N_12221,N_11735,N_11796);
or U12222 (N_12222,N_11695,N_11847);
nor U12223 (N_12223,N_11981,N_11645);
and U12224 (N_12224,N_11569,N_11629);
nand U12225 (N_12225,N_11553,N_11710);
or U12226 (N_12226,N_11719,N_11993);
nor U12227 (N_12227,N_11882,N_11921);
nand U12228 (N_12228,N_11736,N_11668);
xor U12229 (N_12229,N_11853,N_11572);
nor U12230 (N_12230,N_11998,N_11916);
or U12231 (N_12231,N_11765,N_11845);
nand U12232 (N_12232,N_11786,N_11874);
or U12233 (N_12233,N_11807,N_11751);
xor U12234 (N_12234,N_11744,N_11676);
nand U12235 (N_12235,N_11966,N_11782);
nand U12236 (N_12236,N_11662,N_11770);
xor U12237 (N_12237,N_11622,N_11626);
xnor U12238 (N_12238,N_11675,N_11745);
xnor U12239 (N_12239,N_11571,N_11756);
nand U12240 (N_12240,N_11836,N_11871);
or U12241 (N_12241,N_11520,N_11831);
or U12242 (N_12242,N_11561,N_11832);
nor U12243 (N_12243,N_11740,N_11811);
xor U12244 (N_12244,N_11678,N_11922);
nor U12245 (N_12245,N_11835,N_11513);
xnor U12246 (N_12246,N_11696,N_11823);
and U12247 (N_12247,N_11602,N_11713);
xor U12248 (N_12248,N_11919,N_11797);
nor U12249 (N_12249,N_11587,N_11789);
or U12250 (N_12250,N_11851,N_11794);
nand U12251 (N_12251,N_11576,N_11534);
xnor U12252 (N_12252,N_11717,N_11879);
or U12253 (N_12253,N_11963,N_11833);
nand U12254 (N_12254,N_11516,N_11774);
nand U12255 (N_12255,N_11732,N_11640);
and U12256 (N_12256,N_11746,N_11665);
or U12257 (N_12257,N_11972,N_11893);
and U12258 (N_12258,N_11791,N_11827);
nand U12259 (N_12259,N_11927,N_11625);
and U12260 (N_12260,N_11609,N_11671);
nand U12261 (N_12261,N_11674,N_11873);
and U12262 (N_12262,N_11517,N_11986);
and U12263 (N_12263,N_11717,N_11931);
nand U12264 (N_12264,N_11643,N_11533);
nand U12265 (N_12265,N_11553,N_11918);
and U12266 (N_12266,N_11575,N_11576);
xnor U12267 (N_12267,N_11711,N_11984);
nand U12268 (N_12268,N_11929,N_11763);
nand U12269 (N_12269,N_11513,N_11956);
xnor U12270 (N_12270,N_11552,N_11913);
nor U12271 (N_12271,N_11783,N_11905);
and U12272 (N_12272,N_11599,N_11918);
and U12273 (N_12273,N_11927,N_11999);
nor U12274 (N_12274,N_11611,N_11543);
nand U12275 (N_12275,N_11552,N_11875);
nand U12276 (N_12276,N_11822,N_11991);
nand U12277 (N_12277,N_11839,N_11556);
nor U12278 (N_12278,N_11654,N_11926);
nor U12279 (N_12279,N_11901,N_11504);
xnor U12280 (N_12280,N_11821,N_11958);
or U12281 (N_12281,N_11527,N_11695);
nor U12282 (N_12282,N_11713,N_11531);
nand U12283 (N_12283,N_11991,N_11883);
or U12284 (N_12284,N_11901,N_11786);
xor U12285 (N_12285,N_11608,N_11900);
and U12286 (N_12286,N_11521,N_11501);
or U12287 (N_12287,N_11932,N_11639);
or U12288 (N_12288,N_11608,N_11975);
xnor U12289 (N_12289,N_11576,N_11558);
xnor U12290 (N_12290,N_11779,N_11908);
or U12291 (N_12291,N_11939,N_11935);
nor U12292 (N_12292,N_11970,N_11846);
nor U12293 (N_12293,N_11958,N_11718);
xnor U12294 (N_12294,N_11538,N_11612);
and U12295 (N_12295,N_11618,N_11676);
nor U12296 (N_12296,N_11930,N_11916);
nor U12297 (N_12297,N_11621,N_11976);
xor U12298 (N_12298,N_11770,N_11554);
or U12299 (N_12299,N_11533,N_11997);
nor U12300 (N_12300,N_11960,N_11575);
or U12301 (N_12301,N_11904,N_11681);
and U12302 (N_12302,N_11525,N_11578);
xnor U12303 (N_12303,N_11698,N_11783);
nand U12304 (N_12304,N_11928,N_11708);
xor U12305 (N_12305,N_11900,N_11713);
and U12306 (N_12306,N_11721,N_11958);
xnor U12307 (N_12307,N_11661,N_11974);
nand U12308 (N_12308,N_11549,N_11812);
nand U12309 (N_12309,N_11679,N_11999);
xor U12310 (N_12310,N_11889,N_11945);
nand U12311 (N_12311,N_11638,N_11640);
xnor U12312 (N_12312,N_11919,N_11680);
and U12313 (N_12313,N_11844,N_11712);
and U12314 (N_12314,N_11871,N_11663);
xor U12315 (N_12315,N_11798,N_11948);
and U12316 (N_12316,N_11668,N_11532);
or U12317 (N_12317,N_11533,N_11979);
and U12318 (N_12318,N_11525,N_11909);
and U12319 (N_12319,N_11656,N_11944);
nand U12320 (N_12320,N_11613,N_11643);
nand U12321 (N_12321,N_11713,N_11606);
nor U12322 (N_12322,N_11997,N_11507);
nor U12323 (N_12323,N_11927,N_11627);
nor U12324 (N_12324,N_11888,N_11715);
or U12325 (N_12325,N_11611,N_11616);
and U12326 (N_12326,N_11849,N_11604);
and U12327 (N_12327,N_11600,N_11849);
and U12328 (N_12328,N_11722,N_11904);
or U12329 (N_12329,N_11569,N_11671);
and U12330 (N_12330,N_11715,N_11846);
nand U12331 (N_12331,N_11752,N_11757);
and U12332 (N_12332,N_11572,N_11767);
nand U12333 (N_12333,N_11993,N_11723);
nand U12334 (N_12334,N_11671,N_11655);
and U12335 (N_12335,N_11937,N_11834);
nor U12336 (N_12336,N_11794,N_11898);
nor U12337 (N_12337,N_11962,N_11687);
xor U12338 (N_12338,N_11613,N_11620);
or U12339 (N_12339,N_11585,N_11911);
nor U12340 (N_12340,N_11934,N_11871);
nand U12341 (N_12341,N_11967,N_11987);
nand U12342 (N_12342,N_11942,N_11797);
or U12343 (N_12343,N_11981,N_11541);
and U12344 (N_12344,N_11755,N_11843);
and U12345 (N_12345,N_11979,N_11777);
nor U12346 (N_12346,N_11674,N_11640);
or U12347 (N_12347,N_11746,N_11978);
xor U12348 (N_12348,N_11574,N_11757);
and U12349 (N_12349,N_11589,N_11963);
nor U12350 (N_12350,N_11554,N_11758);
nor U12351 (N_12351,N_11653,N_11522);
xor U12352 (N_12352,N_11573,N_11792);
or U12353 (N_12353,N_11978,N_11518);
nand U12354 (N_12354,N_11821,N_11876);
xor U12355 (N_12355,N_11736,N_11554);
and U12356 (N_12356,N_11803,N_11678);
nand U12357 (N_12357,N_11704,N_11742);
nand U12358 (N_12358,N_11989,N_11609);
or U12359 (N_12359,N_11956,N_11603);
or U12360 (N_12360,N_11816,N_11888);
or U12361 (N_12361,N_11850,N_11568);
or U12362 (N_12362,N_11623,N_11635);
xnor U12363 (N_12363,N_11731,N_11991);
nand U12364 (N_12364,N_11734,N_11577);
nor U12365 (N_12365,N_11866,N_11607);
nor U12366 (N_12366,N_11559,N_11954);
and U12367 (N_12367,N_11782,N_11885);
and U12368 (N_12368,N_11836,N_11706);
and U12369 (N_12369,N_11602,N_11593);
and U12370 (N_12370,N_11528,N_11857);
or U12371 (N_12371,N_11981,N_11729);
nand U12372 (N_12372,N_11561,N_11503);
xnor U12373 (N_12373,N_11931,N_11905);
nand U12374 (N_12374,N_11901,N_11668);
or U12375 (N_12375,N_11985,N_11518);
nor U12376 (N_12376,N_11506,N_11771);
nor U12377 (N_12377,N_11522,N_11767);
and U12378 (N_12378,N_11770,N_11524);
and U12379 (N_12379,N_11789,N_11632);
or U12380 (N_12380,N_11519,N_11784);
nor U12381 (N_12381,N_11506,N_11606);
or U12382 (N_12382,N_11965,N_11562);
nand U12383 (N_12383,N_11849,N_11697);
and U12384 (N_12384,N_11535,N_11835);
nor U12385 (N_12385,N_11867,N_11728);
nand U12386 (N_12386,N_11712,N_11611);
nor U12387 (N_12387,N_11580,N_11602);
or U12388 (N_12388,N_11822,N_11949);
or U12389 (N_12389,N_11636,N_11757);
nand U12390 (N_12390,N_11777,N_11663);
and U12391 (N_12391,N_11899,N_11826);
nor U12392 (N_12392,N_11702,N_11990);
nor U12393 (N_12393,N_11995,N_11832);
and U12394 (N_12394,N_11794,N_11761);
xor U12395 (N_12395,N_11933,N_11904);
nor U12396 (N_12396,N_11948,N_11848);
nand U12397 (N_12397,N_11806,N_11902);
xnor U12398 (N_12398,N_11520,N_11638);
nand U12399 (N_12399,N_11667,N_11841);
xnor U12400 (N_12400,N_11621,N_11940);
nor U12401 (N_12401,N_11929,N_11674);
nand U12402 (N_12402,N_11692,N_11945);
nor U12403 (N_12403,N_11900,N_11771);
or U12404 (N_12404,N_11758,N_11564);
or U12405 (N_12405,N_11568,N_11984);
xor U12406 (N_12406,N_11854,N_11595);
nor U12407 (N_12407,N_11761,N_11615);
nor U12408 (N_12408,N_11845,N_11949);
xor U12409 (N_12409,N_11975,N_11669);
nand U12410 (N_12410,N_11838,N_11524);
and U12411 (N_12411,N_11552,N_11795);
nor U12412 (N_12412,N_11932,N_11518);
xnor U12413 (N_12413,N_11607,N_11875);
nand U12414 (N_12414,N_11900,N_11907);
or U12415 (N_12415,N_11686,N_11840);
nor U12416 (N_12416,N_11575,N_11685);
and U12417 (N_12417,N_11926,N_11842);
and U12418 (N_12418,N_11770,N_11898);
nand U12419 (N_12419,N_11701,N_11997);
nor U12420 (N_12420,N_11799,N_11536);
nand U12421 (N_12421,N_11962,N_11909);
or U12422 (N_12422,N_11737,N_11757);
and U12423 (N_12423,N_11503,N_11593);
nand U12424 (N_12424,N_11818,N_11615);
and U12425 (N_12425,N_11706,N_11700);
nor U12426 (N_12426,N_11704,N_11611);
or U12427 (N_12427,N_11706,N_11663);
and U12428 (N_12428,N_11513,N_11543);
and U12429 (N_12429,N_11979,N_11960);
and U12430 (N_12430,N_11931,N_11629);
and U12431 (N_12431,N_11626,N_11914);
nor U12432 (N_12432,N_11913,N_11572);
nand U12433 (N_12433,N_11752,N_11824);
nand U12434 (N_12434,N_11746,N_11640);
nand U12435 (N_12435,N_11504,N_11704);
nor U12436 (N_12436,N_11945,N_11732);
nand U12437 (N_12437,N_11772,N_11530);
xor U12438 (N_12438,N_11682,N_11811);
and U12439 (N_12439,N_11942,N_11964);
nor U12440 (N_12440,N_11758,N_11805);
and U12441 (N_12441,N_11792,N_11864);
or U12442 (N_12442,N_11825,N_11912);
or U12443 (N_12443,N_11610,N_11761);
nor U12444 (N_12444,N_11530,N_11802);
and U12445 (N_12445,N_11575,N_11567);
nand U12446 (N_12446,N_11873,N_11855);
nand U12447 (N_12447,N_11849,N_11531);
xor U12448 (N_12448,N_11706,N_11619);
nand U12449 (N_12449,N_11966,N_11600);
nor U12450 (N_12450,N_11720,N_11546);
nor U12451 (N_12451,N_11903,N_11934);
xnor U12452 (N_12452,N_11515,N_11651);
nor U12453 (N_12453,N_11882,N_11919);
or U12454 (N_12454,N_11631,N_11725);
nor U12455 (N_12455,N_11885,N_11929);
xnor U12456 (N_12456,N_11557,N_11650);
xor U12457 (N_12457,N_11852,N_11621);
xor U12458 (N_12458,N_11844,N_11715);
xnor U12459 (N_12459,N_11733,N_11686);
nand U12460 (N_12460,N_11632,N_11503);
or U12461 (N_12461,N_11544,N_11918);
and U12462 (N_12462,N_11623,N_11505);
nand U12463 (N_12463,N_11988,N_11690);
nor U12464 (N_12464,N_11937,N_11975);
nand U12465 (N_12465,N_11517,N_11696);
and U12466 (N_12466,N_11511,N_11780);
or U12467 (N_12467,N_11511,N_11707);
or U12468 (N_12468,N_11928,N_11664);
nand U12469 (N_12469,N_11619,N_11852);
nor U12470 (N_12470,N_11588,N_11745);
nand U12471 (N_12471,N_11542,N_11600);
xor U12472 (N_12472,N_11783,N_11716);
and U12473 (N_12473,N_11771,N_11537);
xnor U12474 (N_12474,N_11982,N_11718);
nand U12475 (N_12475,N_11685,N_11910);
and U12476 (N_12476,N_11918,N_11761);
nor U12477 (N_12477,N_11520,N_11802);
or U12478 (N_12478,N_11742,N_11796);
or U12479 (N_12479,N_11830,N_11738);
nand U12480 (N_12480,N_11819,N_11534);
nand U12481 (N_12481,N_11799,N_11907);
nor U12482 (N_12482,N_11899,N_11808);
nand U12483 (N_12483,N_11893,N_11823);
xnor U12484 (N_12484,N_11576,N_11510);
nor U12485 (N_12485,N_11692,N_11612);
xnor U12486 (N_12486,N_11611,N_11532);
nand U12487 (N_12487,N_11683,N_11898);
nand U12488 (N_12488,N_11516,N_11674);
or U12489 (N_12489,N_11608,N_11776);
xnor U12490 (N_12490,N_11892,N_11604);
or U12491 (N_12491,N_11834,N_11957);
or U12492 (N_12492,N_11866,N_11616);
nor U12493 (N_12493,N_11684,N_11603);
or U12494 (N_12494,N_11606,N_11631);
xnor U12495 (N_12495,N_11839,N_11652);
nand U12496 (N_12496,N_11687,N_11996);
nand U12497 (N_12497,N_11550,N_11613);
nor U12498 (N_12498,N_11677,N_11703);
and U12499 (N_12499,N_11673,N_11617);
nand U12500 (N_12500,N_12192,N_12109);
xor U12501 (N_12501,N_12257,N_12449);
and U12502 (N_12502,N_12350,N_12322);
or U12503 (N_12503,N_12336,N_12218);
xor U12504 (N_12504,N_12389,N_12465);
nand U12505 (N_12505,N_12393,N_12460);
nor U12506 (N_12506,N_12497,N_12209);
xor U12507 (N_12507,N_12335,N_12021);
nor U12508 (N_12508,N_12440,N_12373);
and U12509 (N_12509,N_12341,N_12199);
or U12510 (N_12510,N_12281,N_12365);
nor U12511 (N_12511,N_12427,N_12187);
xor U12512 (N_12512,N_12263,N_12489);
and U12513 (N_12513,N_12158,N_12385);
or U12514 (N_12514,N_12374,N_12207);
and U12515 (N_12515,N_12115,N_12044);
nor U12516 (N_12516,N_12047,N_12306);
nand U12517 (N_12517,N_12215,N_12434);
nand U12518 (N_12518,N_12052,N_12086);
and U12519 (N_12519,N_12185,N_12136);
nand U12520 (N_12520,N_12252,N_12233);
nand U12521 (N_12521,N_12048,N_12349);
nor U12522 (N_12522,N_12193,N_12019);
or U12523 (N_12523,N_12283,N_12162);
nor U12524 (N_12524,N_12334,N_12168);
nor U12525 (N_12525,N_12386,N_12205);
or U12526 (N_12526,N_12108,N_12305);
nand U12527 (N_12527,N_12074,N_12183);
nand U12528 (N_12528,N_12290,N_12255);
and U12529 (N_12529,N_12447,N_12130);
or U12530 (N_12530,N_12325,N_12494);
or U12531 (N_12531,N_12147,N_12362);
and U12532 (N_12532,N_12396,N_12188);
nand U12533 (N_12533,N_12309,N_12190);
and U12534 (N_12534,N_12286,N_12211);
or U12535 (N_12535,N_12467,N_12295);
xor U12536 (N_12536,N_12073,N_12229);
nand U12537 (N_12537,N_12480,N_12101);
nand U12538 (N_12538,N_12079,N_12296);
and U12539 (N_12539,N_12022,N_12264);
nand U12540 (N_12540,N_12144,N_12143);
nor U12541 (N_12541,N_12405,N_12164);
xnor U12542 (N_12542,N_12453,N_12438);
xor U12543 (N_12543,N_12124,N_12107);
nor U12544 (N_12544,N_12236,N_12129);
or U12545 (N_12545,N_12063,N_12093);
xnor U12546 (N_12546,N_12135,N_12031);
and U12547 (N_12547,N_12046,N_12384);
or U12548 (N_12548,N_12251,N_12118);
nor U12549 (N_12549,N_12452,N_12308);
nand U12550 (N_12550,N_12399,N_12456);
nand U12551 (N_12551,N_12020,N_12410);
or U12552 (N_12552,N_12112,N_12003);
nand U12553 (N_12553,N_12298,N_12470);
xor U12554 (N_12554,N_12213,N_12037);
xor U12555 (N_12555,N_12080,N_12420);
and U12556 (N_12556,N_12104,N_12352);
nor U12557 (N_12557,N_12432,N_12398);
or U12558 (N_12558,N_12087,N_12189);
xor U12559 (N_12559,N_12234,N_12089);
xor U12560 (N_12560,N_12176,N_12378);
nor U12561 (N_12561,N_12311,N_12139);
or U12562 (N_12562,N_12149,N_12499);
and U12563 (N_12563,N_12217,N_12276);
or U12564 (N_12564,N_12040,N_12239);
or U12565 (N_12565,N_12237,N_12071);
nand U12566 (N_12566,N_12007,N_12284);
xor U12567 (N_12567,N_12125,N_12201);
nand U12568 (N_12568,N_12408,N_12429);
xnor U12569 (N_12569,N_12267,N_12464);
or U12570 (N_12570,N_12485,N_12203);
or U12571 (N_12571,N_12491,N_12002);
nand U12572 (N_12572,N_12412,N_12307);
xnor U12573 (N_12573,N_12382,N_12430);
and U12574 (N_12574,N_12156,N_12026);
nand U12575 (N_12575,N_12053,N_12262);
nand U12576 (N_12576,N_12253,N_12197);
nor U12577 (N_12577,N_12417,N_12045);
nand U12578 (N_12578,N_12355,N_12072);
xor U12579 (N_12579,N_12221,N_12419);
and U12580 (N_12580,N_12445,N_12466);
nand U12581 (N_12581,N_12312,N_12220);
nand U12582 (N_12582,N_12064,N_12208);
or U12583 (N_12583,N_12292,N_12323);
and U12584 (N_12584,N_12401,N_12161);
nor U12585 (N_12585,N_12145,N_12383);
nand U12586 (N_12586,N_12018,N_12120);
and U12587 (N_12587,N_12038,N_12122);
xor U12588 (N_12588,N_12461,N_12273);
xnor U12589 (N_12589,N_12214,N_12011);
and U12590 (N_12590,N_12414,N_12171);
nand U12591 (N_12591,N_12090,N_12059);
or U12592 (N_12592,N_12486,N_12110);
and U12593 (N_12593,N_12299,N_12354);
and U12594 (N_12594,N_12403,N_12196);
nor U12595 (N_12595,N_12226,N_12084);
nor U12596 (N_12596,N_12289,N_12075);
nor U12597 (N_12597,N_12318,N_12463);
and U12598 (N_12598,N_12132,N_12462);
and U12599 (N_12599,N_12042,N_12395);
nor U12600 (N_12600,N_12015,N_12177);
and U12601 (N_12601,N_12016,N_12367);
xnor U12602 (N_12602,N_12065,N_12433);
or U12603 (N_12603,N_12036,N_12260);
or U12604 (N_12604,N_12076,N_12024);
xnor U12605 (N_12605,N_12448,N_12259);
nand U12606 (N_12606,N_12297,N_12165);
xnor U12607 (N_12607,N_12202,N_12223);
nand U12608 (N_12608,N_12310,N_12092);
xor U12609 (N_12609,N_12041,N_12428);
nor U12610 (N_12610,N_12418,N_12392);
and U12611 (N_12611,N_12319,N_12070);
nand U12612 (N_12612,N_12478,N_12191);
and U12613 (N_12613,N_12128,N_12353);
xor U12614 (N_12614,N_12359,N_12066);
and U12615 (N_12615,N_12397,N_12210);
and U12616 (N_12616,N_12194,N_12009);
xnor U12617 (N_12617,N_12238,N_12057);
xnor U12618 (N_12618,N_12150,N_12415);
or U12619 (N_12619,N_12379,N_12155);
and U12620 (N_12620,N_12081,N_12186);
nor U12621 (N_12621,N_12138,N_12232);
nor U12622 (N_12622,N_12265,N_12443);
xor U12623 (N_12623,N_12316,N_12339);
nor U12624 (N_12624,N_12457,N_12247);
or U12625 (N_12625,N_12056,N_12082);
nor U12626 (N_12626,N_12416,N_12097);
nor U12627 (N_12627,N_12206,N_12370);
or U12628 (N_12628,N_12200,N_12285);
xnor U12629 (N_12629,N_12431,N_12030);
nor U12630 (N_12630,N_12248,N_12357);
nand U12631 (N_12631,N_12400,N_12008);
xor U12632 (N_12632,N_12182,N_12250);
and U12633 (N_12633,N_12424,N_12142);
nand U12634 (N_12634,N_12175,N_12106);
or U12635 (N_12635,N_12490,N_12148);
or U12636 (N_12636,N_12437,N_12146);
nand U12637 (N_12637,N_12083,N_12402);
or U12638 (N_12638,N_12058,N_12288);
nand U12639 (N_12639,N_12013,N_12458);
and U12640 (N_12640,N_12102,N_12291);
nand U12641 (N_12641,N_12167,N_12356);
or U12642 (N_12642,N_12174,N_12421);
xor U12643 (N_12643,N_12231,N_12039);
nand U12644 (N_12644,N_12344,N_12028);
and U12645 (N_12645,N_12303,N_12368);
xor U12646 (N_12646,N_12409,N_12111);
nor U12647 (N_12647,N_12219,N_12241);
nand U12648 (N_12648,N_12023,N_12278);
nor U12649 (N_12649,N_12375,N_12377);
or U12650 (N_12650,N_12178,N_12034);
or U12651 (N_12651,N_12371,N_12387);
xnor U12652 (N_12652,N_12001,N_12269);
nand U12653 (N_12653,N_12321,N_12282);
or U12654 (N_12654,N_12204,N_12360);
nor U12655 (N_12655,N_12159,N_12179);
and U12656 (N_12656,N_12484,N_12180);
nand U12657 (N_12657,N_12266,N_12498);
nand U12658 (N_12658,N_12361,N_12004);
or U12659 (N_12659,N_12450,N_12348);
xnor U12660 (N_12660,N_12436,N_12181);
nand U12661 (N_12661,N_12088,N_12258);
nor U12662 (N_12662,N_12105,N_12469);
and U12663 (N_12663,N_12243,N_12198);
xnor U12664 (N_12664,N_12329,N_12479);
xor U12665 (N_12665,N_12473,N_12471);
nor U12666 (N_12666,N_12027,N_12294);
or U12667 (N_12667,N_12277,N_12212);
or U12668 (N_12668,N_12422,N_12006);
nor U12669 (N_12669,N_12025,N_12423);
nand U12670 (N_12670,N_12119,N_12482);
and U12671 (N_12671,N_12117,N_12315);
nor U12672 (N_12672,N_12035,N_12406);
or U12673 (N_12673,N_12372,N_12351);
nor U12674 (N_12674,N_12363,N_12496);
or U12675 (N_12675,N_12331,N_12012);
xor U12676 (N_12676,N_12451,N_12326);
xor U12677 (N_12677,N_12345,N_12426);
xor U12678 (N_12678,N_12261,N_12195);
nor U12679 (N_12679,N_12272,N_12166);
nand U12680 (N_12680,N_12327,N_12304);
and U12681 (N_12681,N_12133,N_12358);
and U12682 (N_12682,N_12131,N_12293);
or U12683 (N_12683,N_12330,N_12225);
and U12684 (N_12684,N_12390,N_12274);
nor U12685 (N_12685,N_12301,N_12230);
nor U12686 (N_12686,N_12246,N_12366);
or U12687 (N_12687,N_12320,N_12151);
nand U12688 (N_12688,N_12280,N_12442);
nand U12689 (N_12689,N_12407,N_12160);
nor U12690 (N_12690,N_12227,N_12380);
or U12691 (N_12691,N_12488,N_12113);
nand U12692 (N_12692,N_12342,N_12444);
and U12693 (N_12693,N_12094,N_12346);
or U12694 (N_12694,N_12474,N_12347);
nand U12695 (N_12695,N_12340,N_12224);
or U12696 (N_12696,N_12275,N_12014);
nor U12697 (N_12697,N_12069,N_12376);
xnor U12698 (N_12698,N_12245,N_12099);
and U12699 (N_12699,N_12459,N_12369);
xor U12700 (N_12700,N_12439,N_12029);
nor U12701 (N_12701,N_12077,N_12477);
and U12702 (N_12702,N_12121,N_12153);
and U12703 (N_12703,N_12184,N_12157);
nor U12704 (N_12704,N_12085,N_12054);
nor U12705 (N_12705,N_12043,N_12222);
xnor U12706 (N_12706,N_12140,N_12017);
nand U12707 (N_12707,N_12240,N_12333);
nor U12708 (N_12708,N_12061,N_12287);
or U12709 (N_12709,N_12249,N_12254);
and U12710 (N_12710,N_12425,N_12091);
nor U12711 (N_12711,N_12068,N_12067);
nor U12712 (N_12712,N_12126,N_12095);
xor U12713 (N_12713,N_12271,N_12314);
and U12714 (N_12714,N_12476,N_12435);
and U12715 (N_12715,N_12098,N_12242);
or U12716 (N_12716,N_12313,N_12413);
xnor U12717 (N_12717,N_12051,N_12338);
nand U12718 (N_12718,N_12388,N_12337);
or U12719 (N_12719,N_12235,N_12100);
and U12720 (N_12720,N_12343,N_12487);
or U12721 (N_12721,N_12134,N_12170);
and U12722 (N_12722,N_12137,N_12172);
and U12723 (N_12723,N_12127,N_12332);
nor U12724 (N_12724,N_12062,N_12493);
nand U12725 (N_12725,N_12010,N_12078);
and U12726 (N_12726,N_12300,N_12060);
nor U12727 (N_12727,N_12154,N_12324);
nor U12728 (N_12728,N_12317,N_12483);
xnor U12729 (N_12729,N_12163,N_12441);
and U12730 (N_12730,N_12472,N_12270);
or U12731 (N_12731,N_12446,N_12495);
nor U12732 (N_12732,N_12404,N_12103);
and U12733 (N_12733,N_12391,N_12050);
and U12734 (N_12734,N_12481,N_12328);
or U12735 (N_12735,N_12141,N_12244);
nand U12736 (N_12736,N_12268,N_12228);
xor U12737 (N_12737,N_12411,N_12455);
or U12738 (N_12738,N_12256,N_12492);
xor U12739 (N_12739,N_12123,N_12049);
and U12740 (N_12740,N_12096,N_12116);
and U12741 (N_12741,N_12364,N_12173);
or U12742 (N_12742,N_12468,N_12152);
nor U12743 (N_12743,N_12302,N_12005);
nor U12744 (N_12744,N_12000,N_12114);
or U12745 (N_12745,N_12033,N_12279);
and U12746 (N_12746,N_12475,N_12169);
or U12747 (N_12747,N_12216,N_12055);
and U12748 (N_12748,N_12394,N_12032);
nand U12749 (N_12749,N_12381,N_12454);
nand U12750 (N_12750,N_12308,N_12164);
and U12751 (N_12751,N_12470,N_12417);
nand U12752 (N_12752,N_12075,N_12417);
and U12753 (N_12753,N_12253,N_12240);
nor U12754 (N_12754,N_12060,N_12229);
nand U12755 (N_12755,N_12178,N_12376);
nor U12756 (N_12756,N_12356,N_12191);
nand U12757 (N_12757,N_12044,N_12356);
or U12758 (N_12758,N_12312,N_12176);
nand U12759 (N_12759,N_12384,N_12489);
or U12760 (N_12760,N_12477,N_12472);
and U12761 (N_12761,N_12114,N_12072);
and U12762 (N_12762,N_12031,N_12016);
xnor U12763 (N_12763,N_12362,N_12314);
xor U12764 (N_12764,N_12126,N_12428);
xnor U12765 (N_12765,N_12195,N_12391);
and U12766 (N_12766,N_12460,N_12232);
nand U12767 (N_12767,N_12420,N_12463);
nand U12768 (N_12768,N_12069,N_12170);
nand U12769 (N_12769,N_12191,N_12258);
nor U12770 (N_12770,N_12019,N_12214);
and U12771 (N_12771,N_12197,N_12455);
nand U12772 (N_12772,N_12374,N_12343);
nand U12773 (N_12773,N_12215,N_12451);
xor U12774 (N_12774,N_12311,N_12455);
nand U12775 (N_12775,N_12177,N_12139);
nand U12776 (N_12776,N_12084,N_12197);
or U12777 (N_12777,N_12112,N_12345);
and U12778 (N_12778,N_12445,N_12106);
and U12779 (N_12779,N_12364,N_12460);
nand U12780 (N_12780,N_12424,N_12014);
nand U12781 (N_12781,N_12494,N_12267);
nand U12782 (N_12782,N_12365,N_12179);
xor U12783 (N_12783,N_12453,N_12392);
and U12784 (N_12784,N_12044,N_12459);
nor U12785 (N_12785,N_12205,N_12421);
nand U12786 (N_12786,N_12220,N_12113);
or U12787 (N_12787,N_12347,N_12209);
or U12788 (N_12788,N_12083,N_12337);
and U12789 (N_12789,N_12333,N_12180);
nand U12790 (N_12790,N_12186,N_12454);
xnor U12791 (N_12791,N_12356,N_12251);
nand U12792 (N_12792,N_12224,N_12421);
nand U12793 (N_12793,N_12061,N_12410);
and U12794 (N_12794,N_12128,N_12426);
nor U12795 (N_12795,N_12151,N_12242);
xor U12796 (N_12796,N_12056,N_12249);
xor U12797 (N_12797,N_12385,N_12263);
or U12798 (N_12798,N_12135,N_12421);
nand U12799 (N_12799,N_12378,N_12073);
and U12800 (N_12800,N_12286,N_12306);
nand U12801 (N_12801,N_12476,N_12369);
or U12802 (N_12802,N_12263,N_12153);
nor U12803 (N_12803,N_12312,N_12271);
nand U12804 (N_12804,N_12410,N_12473);
and U12805 (N_12805,N_12164,N_12229);
nand U12806 (N_12806,N_12131,N_12274);
nand U12807 (N_12807,N_12316,N_12376);
or U12808 (N_12808,N_12386,N_12259);
nor U12809 (N_12809,N_12245,N_12260);
nor U12810 (N_12810,N_12361,N_12044);
nand U12811 (N_12811,N_12060,N_12033);
xnor U12812 (N_12812,N_12171,N_12364);
nand U12813 (N_12813,N_12387,N_12058);
nand U12814 (N_12814,N_12336,N_12131);
xnor U12815 (N_12815,N_12495,N_12087);
nand U12816 (N_12816,N_12465,N_12382);
nor U12817 (N_12817,N_12481,N_12380);
nand U12818 (N_12818,N_12300,N_12164);
and U12819 (N_12819,N_12399,N_12428);
and U12820 (N_12820,N_12347,N_12283);
and U12821 (N_12821,N_12452,N_12270);
and U12822 (N_12822,N_12174,N_12350);
nor U12823 (N_12823,N_12278,N_12385);
xnor U12824 (N_12824,N_12176,N_12059);
nand U12825 (N_12825,N_12175,N_12305);
and U12826 (N_12826,N_12171,N_12259);
or U12827 (N_12827,N_12020,N_12158);
or U12828 (N_12828,N_12199,N_12042);
nand U12829 (N_12829,N_12385,N_12200);
nand U12830 (N_12830,N_12457,N_12373);
and U12831 (N_12831,N_12274,N_12092);
and U12832 (N_12832,N_12375,N_12379);
xnor U12833 (N_12833,N_12421,N_12223);
nand U12834 (N_12834,N_12065,N_12223);
or U12835 (N_12835,N_12349,N_12277);
nor U12836 (N_12836,N_12385,N_12186);
or U12837 (N_12837,N_12138,N_12270);
nor U12838 (N_12838,N_12025,N_12253);
or U12839 (N_12839,N_12101,N_12286);
or U12840 (N_12840,N_12238,N_12051);
xnor U12841 (N_12841,N_12470,N_12456);
xnor U12842 (N_12842,N_12069,N_12125);
or U12843 (N_12843,N_12169,N_12073);
nor U12844 (N_12844,N_12018,N_12399);
and U12845 (N_12845,N_12348,N_12014);
xnor U12846 (N_12846,N_12172,N_12102);
xor U12847 (N_12847,N_12463,N_12350);
xnor U12848 (N_12848,N_12278,N_12244);
xor U12849 (N_12849,N_12034,N_12221);
and U12850 (N_12850,N_12289,N_12375);
and U12851 (N_12851,N_12400,N_12160);
nand U12852 (N_12852,N_12488,N_12084);
xor U12853 (N_12853,N_12125,N_12056);
or U12854 (N_12854,N_12402,N_12264);
nand U12855 (N_12855,N_12153,N_12056);
xnor U12856 (N_12856,N_12078,N_12352);
and U12857 (N_12857,N_12342,N_12459);
nand U12858 (N_12858,N_12302,N_12388);
and U12859 (N_12859,N_12284,N_12017);
xor U12860 (N_12860,N_12348,N_12436);
or U12861 (N_12861,N_12224,N_12260);
and U12862 (N_12862,N_12370,N_12266);
nand U12863 (N_12863,N_12375,N_12440);
or U12864 (N_12864,N_12319,N_12121);
xor U12865 (N_12865,N_12014,N_12449);
nand U12866 (N_12866,N_12345,N_12479);
xnor U12867 (N_12867,N_12085,N_12148);
nand U12868 (N_12868,N_12493,N_12321);
xor U12869 (N_12869,N_12241,N_12210);
xor U12870 (N_12870,N_12025,N_12382);
and U12871 (N_12871,N_12005,N_12142);
and U12872 (N_12872,N_12049,N_12041);
nor U12873 (N_12873,N_12262,N_12034);
xor U12874 (N_12874,N_12069,N_12402);
xor U12875 (N_12875,N_12307,N_12191);
nand U12876 (N_12876,N_12371,N_12049);
nor U12877 (N_12877,N_12430,N_12440);
xnor U12878 (N_12878,N_12461,N_12328);
nor U12879 (N_12879,N_12306,N_12130);
xor U12880 (N_12880,N_12077,N_12007);
xor U12881 (N_12881,N_12211,N_12107);
xor U12882 (N_12882,N_12365,N_12481);
or U12883 (N_12883,N_12217,N_12014);
or U12884 (N_12884,N_12043,N_12060);
or U12885 (N_12885,N_12003,N_12172);
nor U12886 (N_12886,N_12212,N_12102);
nor U12887 (N_12887,N_12482,N_12108);
nand U12888 (N_12888,N_12115,N_12476);
nand U12889 (N_12889,N_12267,N_12250);
nor U12890 (N_12890,N_12053,N_12488);
nand U12891 (N_12891,N_12305,N_12086);
xor U12892 (N_12892,N_12025,N_12144);
and U12893 (N_12893,N_12248,N_12026);
nand U12894 (N_12894,N_12309,N_12250);
and U12895 (N_12895,N_12088,N_12181);
and U12896 (N_12896,N_12413,N_12415);
nor U12897 (N_12897,N_12127,N_12318);
nand U12898 (N_12898,N_12436,N_12112);
nand U12899 (N_12899,N_12399,N_12136);
and U12900 (N_12900,N_12194,N_12193);
nand U12901 (N_12901,N_12110,N_12231);
nor U12902 (N_12902,N_12179,N_12149);
nand U12903 (N_12903,N_12013,N_12356);
nand U12904 (N_12904,N_12385,N_12321);
xnor U12905 (N_12905,N_12153,N_12321);
and U12906 (N_12906,N_12003,N_12313);
nor U12907 (N_12907,N_12311,N_12291);
or U12908 (N_12908,N_12222,N_12247);
or U12909 (N_12909,N_12040,N_12380);
xor U12910 (N_12910,N_12002,N_12401);
nor U12911 (N_12911,N_12104,N_12457);
xnor U12912 (N_12912,N_12127,N_12006);
nor U12913 (N_12913,N_12252,N_12323);
and U12914 (N_12914,N_12372,N_12473);
xor U12915 (N_12915,N_12231,N_12017);
nor U12916 (N_12916,N_12137,N_12343);
xor U12917 (N_12917,N_12429,N_12315);
and U12918 (N_12918,N_12301,N_12140);
nor U12919 (N_12919,N_12112,N_12091);
and U12920 (N_12920,N_12280,N_12070);
and U12921 (N_12921,N_12364,N_12465);
nand U12922 (N_12922,N_12289,N_12141);
nand U12923 (N_12923,N_12425,N_12418);
nand U12924 (N_12924,N_12163,N_12316);
nand U12925 (N_12925,N_12234,N_12424);
nor U12926 (N_12926,N_12078,N_12365);
xnor U12927 (N_12927,N_12419,N_12218);
and U12928 (N_12928,N_12166,N_12453);
or U12929 (N_12929,N_12357,N_12176);
and U12930 (N_12930,N_12491,N_12389);
or U12931 (N_12931,N_12147,N_12378);
and U12932 (N_12932,N_12409,N_12354);
nand U12933 (N_12933,N_12411,N_12498);
nand U12934 (N_12934,N_12394,N_12196);
or U12935 (N_12935,N_12156,N_12320);
xnor U12936 (N_12936,N_12436,N_12024);
or U12937 (N_12937,N_12067,N_12102);
xnor U12938 (N_12938,N_12429,N_12005);
and U12939 (N_12939,N_12039,N_12344);
and U12940 (N_12940,N_12421,N_12145);
nor U12941 (N_12941,N_12311,N_12398);
xor U12942 (N_12942,N_12485,N_12250);
and U12943 (N_12943,N_12162,N_12449);
or U12944 (N_12944,N_12299,N_12403);
xnor U12945 (N_12945,N_12119,N_12080);
nand U12946 (N_12946,N_12441,N_12326);
xnor U12947 (N_12947,N_12439,N_12192);
and U12948 (N_12948,N_12191,N_12210);
xor U12949 (N_12949,N_12199,N_12417);
xor U12950 (N_12950,N_12378,N_12253);
xor U12951 (N_12951,N_12477,N_12111);
or U12952 (N_12952,N_12409,N_12079);
nand U12953 (N_12953,N_12063,N_12102);
nor U12954 (N_12954,N_12212,N_12258);
and U12955 (N_12955,N_12379,N_12130);
or U12956 (N_12956,N_12337,N_12050);
xor U12957 (N_12957,N_12314,N_12088);
and U12958 (N_12958,N_12017,N_12362);
nand U12959 (N_12959,N_12459,N_12349);
nor U12960 (N_12960,N_12271,N_12238);
and U12961 (N_12961,N_12210,N_12330);
and U12962 (N_12962,N_12030,N_12464);
and U12963 (N_12963,N_12063,N_12469);
or U12964 (N_12964,N_12089,N_12242);
or U12965 (N_12965,N_12039,N_12170);
nor U12966 (N_12966,N_12156,N_12384);
xnor U12967 (N_12967,N_12467,N_12021);
or U12968 (N_12968,N_12453,N_12391);
nor U12969 (N_12969,N_12016,N_12242);
nor U12970 (N_12970,N_12155,N_12478);
nand U12971 (N_12971,N_12441,N_12175);
nand U12972 (N_12972,N_12254,N_12456);
nand U12973 (N_12973,N_12259,N_12074);
nand U12974 (N_12974,N_12102,N_12370);
nor U12975 (N_12975,N_12141,N_12452);
nand U12976 (N_12976,N_12272,N_12157);
and U12977 (N_12977,N_12467,N_12071);
xor U12978 (N_12978,N_12166,N_12307);
or U12979 (N_12979,N_12038,N_12260);
or U12980 (N_12980,N_12360,N_12183);
nor U12981 (N_12981,N_12200,N_12154);
nand U12982 (N_12982,N_12492,N_12431);
and U12983 (N_12983,N_12060,N_12365);
xnor U12984 (N_12984,N_12318,N_12362);
and U12985 (N_12985,N_12274,N_12470);
and U12986 (N_12986,N_12196,N_12275);
nor U12987 (N_12987,N_12364,N_12445);
nand U12988 (N_12988,N_12368,N_12476);
nor U12989 (N_12989,N_12279,N_12120);
nor U12990 (N_12990,N_12270,N_12054);
or U12991 (N_12991,N_12076,N_12399);
nand U12992 (N_12992,N_12167,N_12026);
and U12993 (N_12993,N_12051,N_12469);
and U12994 (N_12994,N_12354,N_12289);
nor U12995 (N_12995,N_12433,N_12031);
and U12996 (N_12996,N_12141,N_12268);
and U12997 (N_12997,N_12012,N_12264);
or U12998 (N_12998,N_12382,N_12298);
or U12999 (N_12999,N_12327,N_12223);
and U13000 (N_13000,N_12540,N_12718);
or U13001 (N_13001,N_12731,N_12987);
xor U13002 (N_13002,N_12904,N_12711);
nor U13003 (N_13003,N_12631,N_12984);
nand U13004 (N_13004,N_12698,N_12957);
nand U13005 (N_13005,N_12894,N_12520);
and U13006 (N_13006,N_12703,N_12535);
and U13007 (N_13007,N_12830,N_12612);
and U13008 (N_13008,N_12893,N_12760);
or U13009 (N_13009,N_12958,N_12614);
and U13010 (N_13010,N_12586,N_12873);
and U13011 (N_13011,N_12645,N_12521);
or U13012 (N_13012,N_12677,N_12647);
or U13013 (N_13013,N_12638,N_12616);
or U13014 (N_13014,N_12835,N_12658);
or U13015 (N_13015,N_12902,N_12544);
and U13016 (N_13016,N_12571,N_12562);
nand U13017 (N_13017,N_12591,N_12945);
nor U13018 (N_13018,N_12793,N_12692);
or U13019 (N_13019,N_12869,N_12615);
nand U13020 (N_13020,N_12595,N_12964);
nand U13021 (N_13021,N_12757,N_12817);
nor U13022 (N_13022,N_12821,N_12702);
nor U13023 (N_13023,N_12989,N_12791);
xor U13024 (N_13024,N_12978,N_12685);
xnor U13025 (N_13025,N_12525,N_12834);
and U13026 (N_13026,N_12510,N_12802);
nand U13027 (N_13027,N_12708,N_12657);
nand U13028 (N_13028,N_12778,N_12988);
nand U13029 (N_13029,N_12626,N_12582);
xor U13030 (N_13030,N_12787,N_12678);
xnor U13031 (N_13031,N_12857,N_12624);
nor U13032 (N_13032,N_12801,N_12738);
or U13033 (N_13033,N_12829,N_12949);
nand U13034 (N_13034,N_12963,N_12734);
and U13035 (N_13035,N_12906,N_12909);
and U13036 (N_13036,N_12669,N_12747);
xor U13037 (N_13037,N_12532,N_12663);
nand U13038 (N_13038,N_12765,N_12683);
and U13039 (N_13039,N_12795,N_12995);
or U13040 (N_13040,N_12719,N_12974);
and U13041 (N_13041,N_12975,N_12985);
xnor U13042 (N_13042,N_12961,N_12870);
nor U13043 (N_13043,N_12642,N_12650);
xor U13044 (N_13044,N_12789,N_12596);
nor U13045 (N_13045,N_12608,N_12790);
xnor U13046 (N_13046,N_12861,N_12932);
xor U13047 (N_13047,N_12737,N_12558);
xnor U13048 (N_13048,N_12664,N_12509);
nor U13049 (N_13049,N_12753,N_12848);
xor U13050 (N_13050,N_12823,N_12607);
and U13051 (N_13051,N_12888,N_12892);
and U13052 (N_13052,N_12813,N_12547);
and U13053 (N_13053,N_12864,N_12621);
or U13054 (N_13054,N_12567,N_12947);
xor U13055 (N_13055,N_12666,N_12751);
xor U13056 (N_13056,N_12966,N_12794);
xor U13057 (N_13057,N_12598,N_12710);
xnor U13058 (N_13058,N_12517,N_12929);
nor U13059 (N_13059,N_12648,N_12889);
nor U13060 (N_13060,N_12552,N_12972);
nor U13061 (N_13061,N_12604,N_12541);
xor U13062 (N_13062,N_12836,N_12976);
or U13063 (N_13063,N_12516,N_12686);
nand U13064 (N_13064,N_12956,N_12943);
nor U13065 (N_13065,N_12706,N_12763);
xnor U13066 (N_13066,N_12611,N_12629);
nor U13067 (N_13067,N_12898,N_12806);
or U13068 (N_13068,N_12785,N_12724);
nand U13069 (N_13069,N_12699,N_12653);
nand U13070 (N_13070,N_12977,N_12917);
nand U13071 (N_13071,N_12996,N_12646);
and U13072 (N_13072,N_12695,N_12837);
and U13073 (N_13073,N_12529,N_12636);
xnor U13074 (N_13074,N_12742,N_12903);
and U13075 (N_13075,N_12878,N_12508);
nand U13076 (N_13076,N_12655,N_12774);
nand U13077 (N_13077,N_12758,N_12736);
nand U13078 (N_13078,N_12761,N_12661);
or U13079 (N_13079,N_12730,N_12746);
nand U13080 (N_13080,N_12969,N_12576);
xnor U13081 (N_13081,N_12735,N_12849);
or U13082 (N_13082,N_12905,N_12784);
nor U13083 (N_13083,N_12716,N_12992);
or U13084 (N_13084,N_12707,N_12752);
nor U13085 (N_13085,N_12759,N_12748);
nand U13086 (N_13086,N_12727,N_12845);
and U13087 (N_13087,N_12769,N_12512);
and U13088 (N_13088,N_12578,N_12715);
or U13089 (N_13089,N_12553,N_12662);
nand U13090 (N_13090,N_12939,N_12628);
or U13091 (N_13091,N_12907,N_12526);
nor U13092 (N_13092,N_12536,N_12643);
and U13093 (N_13093,N_12915,N_12729);
xor U13094 (N_13094,N_12871,N_12862);
nand U13095 (N_13095,N_12965,N_12779);
xnor U13096 (N_13096,N_12998,N_12931);
nand U13097 (N_13097,N_12649,N_12705);
or U13098 (N_13098,N_12739,N_12809);
or U13099 (N_13099,N_12660,N_12533);
nor U13100 (N_13100,N_12798,N_12606);
xnor U13101 (N_13101,N_12808,N_12887);
or U13102 (N_13102,N_12786,N_12524);
nor U13103 (N_13103,N_12539,N_12816);
and U13104 (N_13104,N_12620,N_12986);
and U13105 (N_13105,N_12556,N_12843);
or U13106 (N_13106,N_12781,N_12542);
and U13107 (N_13107,N_12518,N_12818);
xor U13108 (N_13108,N_12537,N_12637);
xnor U13109 (N_13109,N_12920,N_12704);
xor U13110 (N_13110,N_12523,N_12897);
xor U13111 (N_13111,N_12687,N_12910);
xor U13112 (N_13112,N_12555,N_12850);
nand U13113 (N_13113,N_12565,N_12619);
nor U13114 (N_13114,N_12581,N_12713);
nand U13115 (N_13115,N_12842,N_12652);
xnor U13116 (N_13116,N_12772,N_12866);
nand U13117 (N_13117,N_12639,N_12783);
nand U13118 (N_13118,N_12538,N_12709);
or U13119 (N_13119,N_12840,N_12951);
xor U13120 (N_13120,N_12580,N_12827);
nand U13121 (N_13121,N_12914,N_12851);
xnor U13122 (N_13122,N_12665,N_12531);
or U13123 (N_13123,N_12796,N_12979);
xor U13124 (N_13124,N_12853,N_12993);
and U13125 (N_13125,N_12560,N_12839);
and U13126 (N_13126,N_12955,N_12749);
or U13127 (N_13127,N_12792,N_12859);
xnor U13128 (N_13128,N_12880,N_12812);
and U13129 (N_13129,N_12575,N_12923);
nand U13130 (N_13130,N_12755,N_12745);
and U13131 (N_13131,N_12550,N_12981);
nand U13132 (N_13132,N_12673,N_12997);
nor U13133 (N_13133,N_12999,N_12912);
nor U13134 (N_13134,N_12824,N_12674);
nand U13135 (N_13135,N_12603,N_12900);
xnor U13136 (N_13136,N_12971,N_12500);
or U13137 (N_13137,N_12640,N_12811);
and U13138 (N_13138,N_12896,N_12968);
xnor U13139 (N_13139,N_12950,N_12941);
nor U13140 (N_13140,N_12882,N_12916);
xor U13141 (N_13141,N_12501,N_12651);
nor U13142 (N_13142,N_12919,N_12743);
xor U13143 (N_13143,N_12505,N_12933);
or U13144 (N_13144,N_12881,N_12630);
xnor U13145 (N_13145,N_12583,N_12800);
or U13146 (N_13146,N_12574,N_12566);
and U13147 (N_13147,N_12515,N_12854);
nand U13148 (N_13148,N_12828,N_12723);
xnor U13149 (N_13149,N_12768,N_12938);
or U13150 (N_13150,N_12623,N_12921);
nor U13151 (N_13151,N_12918,N_12573);
nor U13152 (N_13152,N_12617,N_12762);
xor U13153 (N_13153,N_12569,N_12886);
and U13154 (N_13154,N_12770,N_12925);
or U13155 (N_13155,N_12502,N_12568);
nand U13156 (N_13156,N_12590,N_12973);
nor U13157 (N_13157,N_12883,N_12668);
nor U13158 (N_13158,N_12884,N_12775);
or U13159 (N_13159,N_12940,N_12740);
xnor U13160 (N_13160,N_12970,N_12530);
xor U13161 (N_13161,N_12507,N_12534);
or U13162 (N_13162,N_12874,N_12506);
nor U13163 (N_13163,N_12585,N_12641);
and U13164 (N_13164,N_12511,N_12503);
xnor U13165 (N_13165,N_12927,N_12960);
xnor U13166 (N_13166,N_12814,N_12557);
or U13167 (N_13167,N_12670,N_12924);
and U13168 (N_13168,N_12764,N_12911);
or U13169 (N_13169,N_12721,N_12600);
and U13170 (N_13170,N_12601,N_12717);
and U13171 (N_13171,N_12519,N_12691);
xnor U13172 (N_13172,N_12936,N_12788);
xor U13173 (N_13173,N_12618,N_12667);
xor U13174 (N_13174,N_12934,N_12797);
and U13175 (N_13175,N_12644,N_12587);
nor U13176 (N_13176,N_12528,N_12863);
and U13177 (N_13177,N_12782,N_12820);
or U13178 (N_13178,N_12563,N_12991);
xor U13179 (N_13179,N_12690,N_12688);
xor U13180 (N_13180,N_12609,N_12545);
xnor U13181 (N_13181,N_12953,N_12588);
and U13182 (N_13182,N_12926,N_12865);
xor U13183 (N_13183,N_12773,N_12899);
and U13184 (N_13184,N_12799,N_12895);
xor U13185 (N_13185,N_12944,N_12728);
or U13186 (N_13186,N_12838,N_12803);
xor U13187 (N_13187,N_12634,N_12659);
and U13188 (N_13188,N_12771,N_12689);
or U13189 (N_13189,N_12831,N_12879);
nor U13190 (N_13190,N_12697,N_12846);
and U13191 (N_13191,N_12696,N_12513);
or U13192 (N_13192,N_12844,N_12858);
xor U13193 (N_13193,N_12543,N_12935);
or U13194 (N_13194,N_12684,N_12891);
nand U13195 (N_13195,N_12613,N_12875);
or U13196 (N_13196,N_12867,N_12610);
and U13197 (N_13197,N_12832,N_12942);
and U13198 (N_13198,N_12671,N_12672);
nor U13199 (N_13199,N_12675,N_12514);
xnor U13200 (N_13200,N_12913,N_12805);
xor U13201 (N_13201,N_12732,N_12930);
nand U13202 (N_13202,N_12990,N_12983);
nand U13203 (N_13203,N_12627,N_12744);
nor U13204 (N_13204,N_12527,N_12777);
or U13205 (N_13205,N_12701,N_12780);
and U13206 (N_13206,N_12712,N_12890);
nor U13207 (N_13207,N_12833,N_12682);
and U13208 (N_13208,N_12577,N_12554);
or U13209 (N_13209,N_12852,N_12570);
or U13210 (N_13210,N_12522,N_12579);
xor U13211 (N_13211,N_12714,N_12726);
nand U13212 (N_13212,N_12559,N_12605);
xnor U13213 (N_13213,N_12922,N_12632);
xnor U13214 (N_13214,N_12810,N_12948);
nand U13215 (N_13215,N_12928,N_12901);
nand U13216 (N_13216,N_12872,N_12720);
nor U13217 (N_13217,N_12967,N_12756);
xnor U13218 (N_13218,N_12593,N_12959);
or U13219 (N_13219,N_12681,N_12819);
nand U13220 (N_13220,N_12847,N_12725);
xor U13221 (N_13221,N_12548,N_12822);
or U13222 (N_13222,N_12954,N_12622);
nand U13223 (N_13223,N_12980,N_12767);
or U13224 (N_13224,N_12592,N_12572);
nor U13225 (N_13225,N_12722,N_12680);
and U13226 (N_13226,N_12885,N_12504);
xor U13227 (N_13227,N_12856,N_12676);
nor U13228 (N_13228,N_12860,N_12584);
nand U13229 (N_13229,N_12750,N_12602);
nor U13230 (N_13230,N_12654,N_12633);
nor U13231 (N_13231,N_12804,N_12855);
nand U13232 (N_13232,N_12825,N_12994);
and U13233 (N_13233,N_12807,N_12868);
xor U13234 (N_13234,N_12546,N_12733);
and U13235 (N_13235,N_12754,N_12815);
nand U13236 (N_13236,N_12952,N_12594);
and U13237 (N_13237,N_12700,N_12876);
or U13238 (N_13238,N_12656,N_12693);
and U13239 (N_13239,N_12561,N_12766);
xor U13240 (N_13240,N_12776,N_12589);
and U13241 (N_13241,N_12946,N_12937);
nor U13242 (N_13242,N_12741,N_12841);
or U13243 (N_13243,N_12826,N_12635);
xnor U13244 (N_13244,N_12625,N_12908);
and U13245 (N_13245,N_12679,N_12551);
or U13246 (N_13246,N_12597,N_12599);
or U13247 (N_13247,N_12564,N_12694);
nor U13248 (N_13248,N_12877,N_12549);
nor U13249 (N_13249,N_12962,N_12982);
nand U13250 (N_13250,N_12977,N_12559);
xnor U13251 (N_13251,N_12529,N_12702);
nor U13252 (N_13252,N_12750,N_12716);
xnor U13253 (N_13253,N_12718,N_12583);
and U13254 (N_13254,N_12755,N_12881);
and U13255 (N_13255,N_12762,N_12828);
xnor U13256 (N_13256,N_12674,N_12571);
nand U13257 (N_13257,N_12552,N_12798);
nand U13258 (N_13258,N_12743,N_12573);
or U13259 (N_13259,N_12899,N_12808);
nand U13260 (N_13260,N_12910,N_12553);
xor U13261 (N_13261,N_12864,N_12721);
and U13262 (N_13262,N_12637,N_12858);
and U13263 (N_13263,N_12930,N_12643);
nor U13264 (N_13264,N_12533,N_12904);
or U13265 (N_13265,N_12604,N_12606);
nand U13266 (N_13266,N_12501,N_12826);
xnor U13267 (N_13267,N_12954,N_12542);
nand U13268 (N_13268,N_12645,N_12811);
or U13269 (N_13269,N_12978,N_12640);
and U13270 (N_13270,N_12515,N_12846);
and U13271 (N_13271,N_12549,N_12931);
nor U13272 (N_13272,N_12682,N_12584);
or U13273 (N_13273,N_12855,N_12522);
nor U13274 (N_13274,N_12768,N_12661);
or U13275 (N_13275,N_12657,N_12694);
xnor U13276 (N_13276,N_12532,N_12827);
xnor U13277 (N_13277,N_12557,N_12652);
xor U13278 (N_13278,N_12641,N_12557);
and U13279 (N_13279,N_12683,N_12519);
nand U13280 (N_13280,N_12856,N_12532);
nor U13281 (N_13281,N_12973,N_12900);
nand U13282 (N_13282,N_12743,N_12629);
or U13283 (N_13283,N_12763,N_12652);
xnor U13284 (N_13284,N_12510,N_12702);
or U13285 (N_13285,N_12831,N_12797);
xnor U13286 (N_13286,N_12937,N_12721);
xor U13287 (N_13287,N_12632,N_12527);
nand U13288 (N_13288,N_12618,N_12971);
and U13289 (N_13289,N_12509,N_12686);
nand U13290 (N_13290,N_12946,N_12547);
nand U13291 (N_13291,N_12558,N_12579);
nor U13292 (N_13292,N_12762,N_12712);
or U13293 (N_13293,N_12809,N_12773);
and U13294 (N_13294,N_12757,N_12682);
or U13295 (N_13295,N_12827,N_12930);
and U13296 (N_13296,N_12922,N_12743);
xor U13297 (N_13297,N_12849,N_12995);
and U13298 (N_13298,N_12761,N_12926);
or U13299 (N_13299,N_12690,N_12950);
nand U13300 (N_13300,N_12645,N_12926);
and U13301 (N_13301,N_12750,N_12507);
or U13302 (N_13302,N_12628,N_12775);
or U13303 (N_13303,N_12542,N_12867);
xor U13304 (N_13304,N_12753,N_12811);
or U13305 (N_13305,N_12531,N_12833);
nor U13306 (N_13306,N_12761,N_12975);
or U13307 (N_13307,N_12885,N_12512);
nand U13308 (N_13308,N_12553,N_12933);
nand U13309 (N_13309,N_12652,N_12653);
and U13310 (N_13310,N_12547,N_12631);
and U13311 (N_13311,N_12875,N_12597);
xor U13312 (N_13312,N_12909,N_12667);
xnor U13313 (N_13313,N_12558,N_12960);
nor U13314 (N_13314,N_12838,N_12699);
or U13315 (N_13315,N_12778,N_12591);
or U13316 (N_13316,N_12963,N_12897);
and U13317 (N_13317,N_12992,N_12699);
and U13318 (N_13318,N_12513,N_12521);
nor U13319 (N_13319,N_12522,N_12573);
and U13320 (N_13320,N_12779,N_12676);
or U13321 (N_13321,N_12774,N_12630);
or U13322 (N_13322,N_12818,N_12744);
nor U13323 (N_13323,N_12710,N_12587);
and U13324 (N_13324,N_12670,N_12538);
nor U13325 (N_13325,N_12896,N_12798);
nor U13326 (N_13326,N_12730,N_12551);
and U13327 (N_13327,N_12647,N_12987);
or U13328 (N_13328,N_12652,N_12761);
nand U13329 (N_13329,N_12700,N_12871);
or U13330 (N_13330,N_12791,N_12878);
nand U13331 (N_13331,N_12932,N_12906);
or U13332 (N_13332,N_12541,N_12832);
xnor U13333 (N_13333,N_12662,N_12752);
or U13334 (N_13334,N_12769,N_12639);
nor U13335 (N_13335,N_12784,N_12686);
or U13336 (N_13336,N_12892,N_12845);
nor U13337 (N_13337,N_12899,N_12836);
or U13338 (N_13338,N_12809,N_12778);
and U13339 (N_13339,N_12953,N_12848);
and U13340 (N_13340,N_12698,N_12862);
nand U13341 (N_13341,N_12822,N_12562);
xnor U13342 (N_13342,N_12713,N_12721);
nor U13343 (N_13343,N_12746,N_12818);
and U13344 (N_13344,N_12966,N_12855);
xnor U13345 (N_13345,N_12547,N_12656);
nand U13346 (N_13346,N_12872,N_12643);
nand U13347 (N_13347,N_12680,N_12578);
xor U13348 (N_13348,N_12771,N_12918);
xnor U13349 (N_13349,N_12523,N_12874);
nand U13350 (N_13350,N_12901,N_12770);
nand U13351 (N_13351,N_12924,N_12643);
nand U13352 (N_13352,N_12855,N_12667);
xnor U13353 (N_13353,N_12822,N_12526);
nor U13354 (N_13354,N_12840,N_12890);
or U13355 (N_13355,N_12924,N_12631);
and U13356 (N_13356,N_12799,N_12772);
and U13357 (N_13357,N_12983,N_12738);
or U13358 (N_13358,N_12711,N_12572);
nand U13359 (N_13359,N_12737,N_12704);
and U13360 (N_13360,N_12953,N_12716);
and U13361 (N_13361,N_12664,N_12563);
xnor U13362 (N_13362,N_12808,N_12909);
or U13363 (N_13363,N_12634,N_12783);
nor U13364 (N_13364,N_12701,N_12869);
xnor U13365 (N_13365,N_12754,N_12700);
nor U13366 (N_13366,N_12979,N_12565);
nand U13367 (N_13367,N_12615,N_12878);
and U13368 (N_13368,N_12966,N_12751);
and U13369 (N_13369,N_12596,N_12660);
xor U13370 (N_13370,N_12644,N_12706);
nand U13371 (N_13371,N_12683,N_12700);
nand U13372 (N_13372,N_12796,N_12977);
nand U13373 (N_13373,N_12654,N_12921);
nand U13374 (N_13374,N_12555,N_12501);
nand U13375 (N_13375,N_12990,N_12971);
xor U13376 (N_13376,N_12994,N_12624);
nand U13377 (N_13377,N_12898,N_12867);
or U13378 (N_13378,N_12824,N_12734);
nand U13379 (N_13379,N_12886,N_12596);
and U13380 (N_13380,N_12979,N_12855);
and U13381 (N_13381,N_12701,N_12516);
nand U13382 (N_13382,N_12987,N_12777);
and U13383 (N_13383,N_12718,N_12533);
nand U13384 (N_13384,N_12516,N_12784);
xor U13385 (N_13385,N_12765,N_12969);
nor U13386 (N_13386,N_12851,N_12963);
or U13387 (N_13387,N_12929,N_12742);
nor U13388 (N_13388,N_12637,N_12526);
nand U13389 (N_13389,N_12669,N_12592);
xor U13390 (N_13390,N_12701,N_12893);
or U13391 (N_13391,N_12718,N_12508);
and U13392 (N_13392,N_12520,N_12506);
and U13393 (N_13393,N_12835,N_12552);
xnor U13394 (N_13394,N_12647,N_12759);
nor U13395 (N_13395,N_12751,N_12675);
nand U13396 (N_13396,N_12910,N_12895);
nand U13397 (N_13397,N_12769,N_12809);
xnor U13398 (N_13398,N_12716,N_12526);
nor U13399 (N_13399,N_12972,N_12903);
nand U13400 (N_13400,N_12899,N_12859);
or U13401 (N_13401,N_12612,N_12807);
nor U13402 (N_13402,N_12957,N_12829);
nand U13403 (N_13403,N_12897,N_12823);
nand U13404 (N_13404,N_12525,N_12801);
xnor U13405 (N_13405,N_12733,N_12690);
nor U13406 (N_13406,N_12513,N_12502);
and U13407 (N_13407,N_12933,N_12527);
and U13408 (N_13408,N_12754,N_12705);
xor U13409 (N_13409,N_12862,N_12857);
xnor U13410 (N_13410,N_12526,N_12665);
xor U13411 (N_13411,N_12971,N_12548);
nor U13412 (N_13412,N_12938,N_12585);
nand U13413 (N_13413,N_12678,N_12598);
or U13414 (N_13414,N_12893,N_12957);
nand U13415 (N_13415,N_12908,N_12691);
nor U13416 (N_13416,N_12758,N_12936);
xor U13417 (N_13417,N_12887,N_12991);
and U13418 (N_13418,N_12992,N_12782);
or U13419 (N_13419,N_12696,N_12846);
or U13420 (N_13420,N_12511,N_12767);
nor U13421 (N_13421,N_12995,N_12617);
nor U13422 (N_13422,N_12642,N_12959);
nor U13423 (N_13423,N_12708,N_12629);
xnor U13424 (N_13424,N_12947,N_12568);
and U13425 (N_13425,N_12908,N_12893);
or U13426 (N_13426,N_12505,N_12937);
xor U13427 (N_13427,N_12964,N_12977);
and U13428 (N_13428,N_12944,N_12576);
nor U13429 (N_13429,N_12553,N_12552);
or U13430 (N_13430,N_12937,N_12631);
nor U13431 (N_13431,N_12707,N_12888);
and U13432 (N_13432,N_12748,N_12736);
nand U13433 (N_13433,N_12708,N_12572);
and U13434 (N_13434,N_12562,N_12512);
and U13435 (N_13435,N_12662,N_12854);
nand U13436 (N_13436,N_12640,N_12896);
or U13437 (N_13437,N_12935,N_12501);
nor U13438 (N_13438,N_12789,N_12699);
nand U13439 (N_13439,N_12797,N_12612);
or U13440 (N_13440,N_12985,N_12692);
nor U13441 (N_13441,N_12751,N_12747);
nor U13442 (N_13442,N_12702,N_12862);
nand U13443 (N_13443,N_12857,N_12884);
and U13444 (N_13444,N_12705,N_12914);
xor U13445 (N_13445,N_12620,N_12735);
nor U13446 (N_13446,N_12779,N_12653);
xnor U13447 (N_13447,N_12621,N_12707);
xnor U13448 (N_13448,N_12593,N_12777);
or U13449 (N_13449,N_12552,N_12717);
or U13450 (N_13450,N_12748,N_12888);
xor U13451 (N_13451,N_12714,N_12838);
and U13452 (N_13452,N_12700,N_12706);
nand U13453 (N_13453,N_12724,N_12973);
xnor U13454 (N_13454,N_12543,N_12971);
nor U13455 (N_13455,N_12818,N_12856);
xnor U13456 (N_13456,N_12664,N_12669);
xor U13457 (N_13457,N_12794,N_12597);
nand U13458 (N_13458,N_12886,N_12721);
xor U13459 (N_13459,N_12548,N_12927);
nor U13460 (N_13460,N_12882,N_12863);
and U13461 (N_13461,N_12983,N_12534);
or U13462 (N_13462,N_12594,N_12603);
nor U13463 (N_13463,N_12696,N_12529);
nor U13464 (N_13464,N_12824,N_12709);
nor U13465 (N_13465,N_12972,N_12543);
or U13466 (N_13466,N_12784,N_12533);
or U13467 (N_13467,N_12583,N_12586);
nand U13468 (N_13468,N_12688,N_12502);
nand U13469 (N_13469,N_12658,N_12877);
or U13470 (N_13470,N_12917,N_12585);
nor U13471 (N_13471,N_12792,N_12664);
nand U13472 (N_13472,N_12538,N_12698);
nand U13473 (N_13473,N_12931,N_12674);
xor U13474 (N_13474,N_12976,N_12686);
nor U13475 (N_13475,N_12622,N_12708);
xor U13476 (N_13476,N_12655,N_12838);
xnor U13477 (N_13477,N_12533,N_12735);
or U13478 (N_13478,N_12602,N_12645);
xnor U13479 (N_13479,N_12509,N_12828);
and U13480 (N_13480,N_12593,N_12744);
or U13481 (N_13481,N_12985,N_12551);
and U13482 (N_13482,N_12587,N_12887);
or U13483 (N_13483,N_12837,N_12547);
and U13484 (N_13484,N_12912,N_12602);
or U13485 (N_13485,N_12804,N_12918);
nand U13486 (N_13486,N_12934,N_12833);
nand U13487 (N_13487,N_12646,N_12637);
or U13488 (N_13488,N_12531,N_12579);
nand U13489 (N_13489,N_12981,N_12908);
or U13490 (N_13490,N_12581,N_12652);
nand U13491 (N_13491,N_12944,N_12839);
and U13492 (N_13492,N_12904,N_12610);
nand U13493 (N_13493,N_12928,N_12755);
nand U13494 (N_13494,N_12623,N_12677);
or U13495 (N_13495,N_12913,N_12662);
and U13496 (N_13496,N_12771,N_12851);
xnor U13497 (N_13497,N_12644,N_12841);
xnor U13498 (N_13498,N_12713,N_12527);
nand U13499 (N_13499,N_12590,N_12998);
nand U13500 (N_13500,N_13009,N_13192);
and U13501 (N_13501,N_13314,N_13019);
xor U13502 (N_13502,N_13116,N_13073);
nor U13503 (N_13503,N_13223,N_13341);
or U13504 (N_13504,N_13124,N_13328);
and U13505 (N_13505,N_13117,N_13059);
xnor U13506 (N_13506,N_13312,N_13180);
or U13507 (N_13507,N_13078,N_13371);
nor U13508 (N_13508,N_13159,N_13228);
nand U13509 (N_13509,N_13160,N_13275);
or U13510 (N_13510,N_13149,N_13102);
nor U13511 (N_13511,N_13225,N_13268);
nand U13512 (N_13512,N_13274,N_13114);
nor U13513 (N_13513,N_13375,N_13016);
xnor U13514 (N_13514,N_13435,N_13253);
or U13515 (N_13515,N_13144,N_13076);
nand U13516 (N_13516,N_13337,N_13445);
or U13517 (N_13517,N_13134,N_13476);
xor U13518 (N_13518,N_13470,N_13377);
or U13519 (N_13519,N_13405,N_13446);
and U13520 (N_13520,N_13096,N_13421);
nor U13521 (N_13521,N_13174,N_13282);
or U13522 (N_13522,N_13012,N_13250);
nand U13523 (N_13523,N_13081,N_13220);
and U13524 (N_13524,N_13013,N_13015);
nand U13525 (N_13525,N_13480,N_13256);
nor U13526 (N_13526,N_13479,N_13370);
and U13527 (N_13527,N_13289,N_13473);
nor U13528 (N_13528,N_13153,N_13173);
nand U13529 (N_13529,N_13464,N_13146);
xor U13530 (N_13530,N_13133,N_13041);
or U13531 (N_13531,N_13376,N_13419);
nor U13532 (N_13532,N_13257,N_13478);
nor U13533 (N_13533,N_13205,N_13097);
xor U13534 (N_13534,N_13202,N_13093);
and U13535 (N_13535,N_13339,N_13482);
nor U13536 (N_13536,N_13054,N_13237);
xnor U13537 (N_13537,N_13235,N_13293);
nand U13538 (N_13538,N_13443,N_13322);
and U13539 (N_13539,N_13332,N_13335);
or U13540 (N_13540,N_13474,N_13025);
or U13541 (N_13541,N_13121,N_13462);
nand U13542 (N_13542,N_13347,N_13083);
nor U13543 (N_13543,N_13033,N_13366);
or U13544 (N_13544,N_13037,N_13069);
nand U13545 (N_13545,N_13457,N_13388);
and U13546 (N_13546,N_13089,N_13086);
nand U13547 (N_13547,N_13058,N_13447);
or U13548 (N_13548,N_13271,N_13494);
xnor U13549 (N_13549,N_13175,N_13362);
xor U13550 (N_13550,N_13100,N_13245);
nor U13551 (N_13551,N_13183,N_13196);
nor U13552 (N_13552,N_13369,N_13358);
nor U13553 (N_13553,N_13468,N_13024);
nor U13554 (N_13554,N_13346,N_13353);
nand U13555 (N_13555,N_13357,N_13152);
xnor U13556 (N_13556,N_13374,N_13492);
and U13557 (N_13557,N_13137,N_13291);
nand U13558 (N_13558,N_13394,N_13184);
nor U13559 (N_13559,N_13434,N_13057);
nand U13560 (N_13560,N_13000,N_13002);
or U13561 (N_13561,N_13484,N_13277);
and U13562 (N_13562,N_13384,N_13359);
nand U13563 (N_13563,N_13049,N_13380);
xor U13564 (N_13564,N_13030,N_13109);
xor U13565 (N_13565,N_13046,N_13390);
nand U13566 (N_13566,N_13182,N_13067);
and U13567 (N_13567,N_13488,N_13317);
or U13568 (N_13568,N_13234,N_13211);
xor U13569 (N_13569,N_13396,N_13308);
and U13570 (N_13570,N_13307,N_13261);
xnor U13571 (N_13571,N_13349,N_13393);
nor U13572 (N_13572,N_13055,N_13352);
nor U13573 (N_13573,N_13471,N_13284);
xnor U13574 (N_13574,N_13378,N_13456);
or U13575 (N_13575,N_13368,N_13411);
and U13576 (N_13576,N_13401,N_13201);
nand U13577 (N_13577,N_13227,N_13392);
and U13578 (N_13578,N_13112,N_13415);
nand U13579 (N_13579,N_13195,N_13306);
xor U13580 (N_13580,N_13423,N_13383);
and U13581 (N_13581,N_13316,N_13188);
nand U13582 (N_13582,N_13404,N_13338);
and U13583 (N_13583,N_13321,N_13451);
or U13584 (N_13584,N_13226,N_13336);
nand U13585 (N_13585,N_13218,N_13241);
nand U13586 (N_13586,N_13424,N_13491);
and U13587 (N_13587,N_13136,N_13425);
xor U13588 (N_13588,N_13351,N_13130);
or U13589 (N_13589,N_13417,N_13242);
nor U13590 (N_13590,N_13035,N_13427);
and U13591 (N_13591,N_13219,N_13053);
xnor U13592 (N_13592,N_13348,N_13098);
nand U13593 (N_13593,N_13119,N_13062);
or U13594 (N_13594,N_13023,N_13483);
nor U13595 (N_13595,N_13051,N_13458);
and U13596 (N_13596,N_13315,N_13397);
and U13597 (N_13597,N_13481,N_13255);
and U13598 (N_13598,N_13444,N_13150);
xor U13599 (N_13599,N_13386,N_13356);
or U13600 (N_13600,N_13466,N_13420);
and U13601 (N_13601,N_13038,N_13005);
or U13602 (N_13602,N_13467,N_13333);
or U13603 (N_13603,N_13001,N_13068);
and U13604 (N_13604,N_13320,N_13283);
nor U13605 (N_13605,N_13224,N_13441);
xor U13606 (N_13606,N_13095,N_13265);
nor U13607 (N_13607,N_13400,N_13155);
xnor U13608 (N_13608,N_13216,N_13285);
and U13609 (N_13609,N_13452,N_13309);
or U13610 (N_13610,N_13270,N_13170);
and U13611 (N_13611,N_13497,N_13298);
or U13612 (N_13612,N_13197,N_13151);
or U13613 (N_13613,N_13360,N_13442);
nand U13614 (N_13614,N_13344,N_13387);
nor U13615 (N_13615,N_13279,N_13403);
nand U13616 (N_13616,N_13052,N_13409);
or U13617 (N_13617,N_13171,N_13495);
nor U13618 (N_13618,N_13413,N_13026);
nor U13619 (N_13619,N_13094,N_13310);
nand U13620 (N_13620,N_13436,N_13493);
nor U13621 (N_13621,N_13258,N_13162);
xnor U13622 (N_13622,N_13191,N_13263);
and U13623 (N_13623,N_13007,N_13115);
or U13624 (N_13624,N_13430,N_13004);
and U13625 (N_13625,N_13172,N_13131);
nor U13626 (N_13626,N_13440,N_13465);
and U13627 (N_13627,N_13103,N_13463);
and U13628 (N_13628,N_13166,N_13181);
or U13629 (N_13629,N_13450,N_13290);
xor U13630 (N_13630,N_13060,N_13003);
nor U13631 (N_13631,N_13039,N_13240);
nor U13632 (N_13632,N_13105,N_13084);
or U13633 (N_13633,N_13248,N_13247);
nand U13634 (N_13634,N_13295,N_13199);
or U13635 (N_13635,N_13303,N_13043);
and U13636 (N_13636,N_13350,N_13072);
xnor U13637 (N_13637,N_13204,N_13319);
and U13638 (N_13638,N_13264,N_13085);
and U13639 (N_13639,N_13373,N_13048);
or U13640 (N_13640,N_13074,N_13432);
nor U13641 (N_13641,N_13176,N_13126);
and U13642 (N_13642,N_13212,N_13200);
and U13643 (N_13643,N_13262,N_13203);
or U13644 (N_13644,N_13066,N_13042);
xnor U13645 (N_13645,N_13148,N_13207);
or U13646 (N_13646,N_13499,N_13489);
nor U13647 (N_13647,N_13382,N_13008);
or U13648 (N_13648,N_13429,N_13395);
and U13649 (N_13649,N_13461,N_13208);
nor U13650 (N_13650,N_13077,N_13402);
and U13651 (N_13651,N_13281,N_13300);
xnor U13652 (N_13652,N_13034,N_13260);
nand U13653 (N_13653,N_13127,N_13334);
nor U13654 (N_13654,N_13006,N_13305);
or U13655 (N_13655,N_13323,N_13361);
nand U13656 (N_13656,N_13111,N_13331);
xor U13657 (N_13657,N_13414,N_13090);
and U13658 (N_13658,N_13138,N_13193);
and U13659 (N_13659,N_13454,N_13324);
nor U13660 (N_13660,N_13355,N_13177);
and U13661 (N_13661,N_13179,N_13278);
xnor U13662 (N_13662,N_13189,N_13406);
nand U13663 (N_13663,N_13070,N_13367);
nor U13664 (N_13664,N_13311,N_13244);
nand U13665 (N_13665,N_13106,N_13017);
nand U13666 (N_13666,N_13294,N_13164);
and U13667 (N_13667,N_13287,N_13433);
or U13668 (N_13668,N_13063,N_13222);
nand U13669 (N_13669,N_13010,N_13029);
or U13670 (N_13670,N_13439,N_13141);
nor U13671 (N_13671,N_13455,N_13104);
nor U13672 (N_13672,N_13232,N_13139);
or U13673 (N_13673,N_13286,N_13142);
xor U13674 (N_13674,N_13496,N_13354);
xor U13675 (N_13675,N_13485,N_13243);
and U13676 (N_13676,N_13221,N_13469);
or U13677 (N_13677,N_13296,N_13194);
or U13678 (N_13678,N_13259,N_13459);
nor U13679 (N_13679,N_13249,N_13190);
nor U13680 (N_13680,N_13113,N_13299);
or U13681 (N_13681,N_13011,N_13431);
nand U13682 (N_13682,N_13318,N_13163);
or U13683 (N_13683,N_13178,N_13246);
and U13684 (N_13684,N_13428,N_13056);
xor U13685 (N_13685,N_13036,N_13028);
or U13686 (N_13686,N_13280,N_13448);
and U13687 (N_13687,N_13107,N_13267);
xnor U13688 (N_13688,N_13158,N_13426);
and U13689 (N_13689,N_13022,N_13301);
nand U13690 (N_13690,N_13018,N_13110);
nand U13691 (N_13691,N_13140,N_13065);
nand U13692 (N_13692,N_13120,N_13381);
and U13693 (N_13693,N_13418,N_13343);
or U13694 (N_13694,N_13214,N_13327);
xor U13695 (N_13695,N_13449,N_13101);
or U13696 (N_13696,N_13125,N_13385);
nor U13697 (N_13697,N_13391,N_13330);
and U13698 (N_13698,N_13132,N_13365);
or U13699 (N_13699,N_13157,N_13313);
nand U13700 (N_13700,N_13147,N_13088);
xor U13701 (N_13701,N_13292,N_13297);
nor U13702 (N_13702,N_13198,N_13422);
and U13703 (N_13703,N_13486,N_13020);
and U13704 (N_13704,N_13014,N_13075);
nor U13705 (N_13705,N_13438,N_13082);
nand U13706 (N_13706,N_13071,N_13206);
or U13707 (N_13707,N_13122,N_13040);
or U13708 (N_13708,N_13210,N_13399);
and U13709 (N_13709,N_13475,N_13302);
nor U13710 (N_13710,N_13252,N_13407);
xnor U13711 (N_13711,N_13326,N_13498);
nor U13712 (N_13712,N_13437,N_13118);
or U13713 (N_13713,N_13364,N_13080);
nor U13714 (N_13714,N_13161,N_13304);
xor U13715 (N_13715,N_13389,N_13031);
and U13716 (N_13716,N_13398,N_13143);
or U13717 (N_13717,N_13276,N_13236);
nor U13718 (N_13718,N_13050,N_13169);
xnor U13719 (N_13719,N_13213,N_13032);
nand U13720 (N_13720,N_13329,N_13156);
xor U13721 (N_13721,N_13123,N_13363);
nand U13722 (N_13722,N_13273,N_13325);
nor U13723 (N_13723,N_13231,N_13091);
nand U13724 (N_13724,N_13129,N_13145);
xnor U13725 (N_13725,N_13099,N_13408);
nand U13726 (N_13726,N_13154,N_13230);
or U13727 (N_13727,N_13272,N_13079);
and U13728 (N_13728,N_13047,N_13379);
or U13729 (N_13729,N_13345,N_13168);
xnor U13730 (N_13730,N_13044,N_13266);
and U13731 (N_13731,N_13187,N_13108);
xor U13732 (N_13732,N_13128,N_13472);
or U13733 (N_13733,N_13416,N_13238);
nor U13734 (N_13734,N_13412,N_13165);
nor U13735 (N_13735,N_13215,N_13251);
nor U13736 (N_13736,N_13410,N_13487);
and U13737 (N_13737,N_13490,N_13027);
nand U13738 (N_13738,N_13229,N_13021);
or U13739 (N_13739,N_13045,N_13217);
nand U13740 (N_13740,N_13167,N_13233);
and U13741 (N_13741,N_13061,N_13185);
nand U13742 (N_13742,N_13135,N_13092);
nor U13743 (N_13743,N_13340,N_13477);
nand U13744 (N_13744,N_13269,N_13372);
or U13745 (N_13745,N_13186,N_13087);
and U13746 (N_13746,N_13288,N_13460);
or U13747 (N_13747,N_13453,N_13064);
nand U13748 (N_13748,N_13342,N_13239);
and U13749 (N_13749,N_13254,N_13209);
xor U13750 (N_13750,N_13353,N_13485);
and U13751 (N_13751,N_13199,N_13420);
nand U13752 (N_13752,N_13219,N_13144);
and U13753 (N_13753,N_13344,N_13154);
nand U13754 (N_13754,N_13307,N_13259);
or U13755 (N_13755,N_13484,N_13003);
nor U13756 (N_13756,N_13003,N_13357);
xor U13757 (N_13757,N_13261,N_13013);
nand U13758 (N_13758,N_13384,N_13389);
nor U13759 (N_13759,N_13239,N_13233);
xor U13760 (N_13760,N_13417,N_13239);
xor U13761 (N_13761,N_13132,N_13340);
xor U13762 (N_13762,N_13196,N_13423);
or U13763 (N_13763,N_13067,N_13043);
nor U13764 (N_13764,N_13173,N_13074);
and U13765 (N_13765,N_13413,N_13469);
or U13766 (N_13766,N_13345,N_13450);
or U13767 (N_13767,N_13315,N_13477);
nand U13768 (N_13768,N_13486,N_13174);
or U13769 (N_13769,N_13392,N_13345);
xnor U13770 (N_13770,N_13290,N_13370);
xnor U13771 (N_13771,N_13363,N_13035);
or U13772 (N_13772,N_13126,N_13408);
and U13773 (N_13773,N_13027,N_13154);
xnor U13774 (N_13774,N_13403,N_13113);
or U13775 (N_13775,N_13181,N_13232);
xor U13776 (N_13776,N_13147,N_13356);
nand U13777 (N_13777,N_13210,N_13176);
xor U13778 (N_13778,N_13357,N_13403);
or U13779 (N_13779,N_13430,N_13097);
and U13780 (N_13780,N_13465,N_13191);
xor U13781 (N_13781,N_13275,N_13119);
nor U13782 (N_13782,N_13238,N_13363);
nor U13783 (N_13783,N_13150,N_13248);
nor U13784 (N_13784,N_13479,N_13249);
xor U13785 (N_13785,N_13103,N_13472);
and U13786 (N_13786,N_13339,N_13055);
xnor U13787 (N_13787,N_13412,N_13006);
or U13788 (N_13788,N_13008,N_13115);
and U13789 (N_13789,N_13441,N_13129);
xor U13790 (N_13790,N_13139,N_13328);
xnor U13791 (N_13791,N_13400,N_13030);
and U13792 (N_13792,N_13477,N_13015);
or U13793 (N_13793,N_13479,N_13050);
nor U13794 (N_13794,N_13017,N_13078);
nor U13795 (N_13795,N_13012,N_13276);
nand U13796 (N_13796,N_13498,N_13368);
nand U13797 (N_13797,N_13070,N_13425);
or U13798 (N_13798,N_13293,N_13349);
nor U13799 (N_13799,N_13179,N_13236);
xor U13800 (N_13800,N_13100,N_13087);
or U13801 (N_13801,N_13012,N_13051);
nand U13802 (N_13802,N_13431,N_13006);
nand U13803 (N_13803,N_13168,N_13190);
nand U13804 (N_13804,N_13034,N_13318);
nor U13805 (N_13805,N_13424,N_13111);
or U13806 (N_13806,N_13381,N_13475);
and U13807 (N_13807,N_13032,N_13327);
xnor U13808 (N_13808,N_13046,N_13463);
nor U13809 (N_13809,N_13322,N_13345);
nor U13810 (N_13810,N_13269,N_13010);
nor U13811 (N_13811,N_13286,N_13053);
nand U13812 (N_13812,N_13253,N_13052);
nand U13813 (N_13813,N_13209,N_13479);
xor U13814 (N_13814,N_13067,N_13084);
nor U13815 (N_13815,N_13188,N_13470);
and U13816 (N_13816,N_13414,N_13486);
nand U13817 (N_13817,N_13446,N_13236);
nor U13818 (N_13818,N_13096,N_13276);
nor U13819 (N_13819,N_13081,N_13176);
nor U13820 (N_13820,N_13048,N_13460);
nor U13821 (N_13821,N_13409,N_13252);
and U13822 (N_13822,N_13071,N_13402);
nor U13823 (N_13823,N_13164,N_13367);
or U13824 (N_13824,N_13426,N_13486);
nor U13825 (N_13825,N_13310,N_13355);
or U13826 (N_13826,N_13138,N_13221);
and U13827 (N_13827,N_13165,N_13292);
nand U13828 (N_13828,N_13151,N_13380);
nor U13829 (N_13829,N_13070,N_13019);
nand U13830 (N_13830,N_13363,N_13386);
nand U13831 (N_13831,N_13121,N_13325);
nor U13832 (N_13832,N_13337,N_13130);
nand U13833 (N_13833,N_13480,N_13421);
nor U13834 (N_13834,N_13353,N_13330);
xor U13835 (N_13835,N_13465,N_13368);
or U13836 (N_13836,N_13493,N_13245);
and U13837 (N_13837,N_13343,N_13297);
or U13838 (N_13838,N_13157,N_13499);
or U13839 (N_13839,N_13439,N_13222);
xnor U13840 (N_13840,N_13334,N_13146);
nand U13841 (N_13841,N_13165,N_13136);
or U13842 (N_13842,N_13319,N_13294);
nand U13843 (N_13843,N_13314,N_13292);
or U13844 (N_13844,N_13024,N_13128);
or U13845 (N_13845,N_13461,N_13025);
or U13846 (N_13846,N_13226,N_13169);
nand U13847 (N_13847,N_13235,N_13238);
nor U13848 (N_13848,N_13042,N_13299);
nor U13849 (N_13849,N_13414,N_13028);
xor U13850 (N_13850,N_13259,N_13302);
or U13851 (N_13851,N_13385,N_13293);
or U13852 (N_13852,N_13376,N_13221);
nand U13853 (N_13853,N_13386,N_13261);
or U13854 (N_13854,N_13253,N_13197);
nand U13855 (N_13855,N_13105,N_13109);
nor U13856 (N_13856,N_13301,N_13104);
and U13857 (N_13857,N_13047,N_13475);
nor U13858 (N_13858,N_13019,N_13426);
nand U13859 (N_13859,N_13208,N_13169);
or U13860 (N_13860,N_13291,N_13251);
nor U13861 (N_13861,N_13311,N_13404);
nand U13862 (N_13862,N_13091,N_13057);
or U13863 (N_13863,N_13168,N_13489);
or U13864 (N_13864,N_13154,N_13454);
and U13865 (N_13865,N_13114,N_13306);
xnor U13866 (N_13866,N_13432,N_13291);
nand U13867 (N_13867,N_13041,N_13476);
or U13868 (N_13868,N_13434,N_13234);
xnor U13869 (N_13869,N_13402,N_13057);
nand U13870 (N_13870,N_13273,N_13135);
xnor U13871 (N_13871,N_13458,N_13334);
or U13872 (N_13872,N_13305,N_13348);
xnor U13873 (N_13873,N_13134,N_13264);
and U13874 (N_13874,N_13278,N_13265);
xnor U13875 (N_13875,N_13289,N_13232);
and U13876 (N_13876,N_13142,N_13221);
xnor U13877 (N_13877,N_13457,N_13264);
and U13878 (N_13878,N_13357,N_13296);
xnor U13879 (N_13879,N_13397,N_13495);
nor U13880 (N_13880,N_13256,N_13083);
nand U13881 (N_13881,N_13218,N_13087);
nor U13882 (N_13882,N_13219,N_13174);
and U13883 (N_13883,N_13471,N_13385);
nor U13884 (N_13884,N_13294,N_13351);
nand U13885 (N_13885,N_13106,N_13071);
or U13886 (N_13886,N_13174,N_13329);
and U13887 (N_13887,N_13303,N_13186);
nand U13888 (N_13888,N_13349,N_13221);
and U13889 (N_13889,N_13396,N_13242);
nand U13890 (N_13890,N_13347,N_13297);
nand U13891 (N_13891,N_13245,N_13462);
xor U13892 (N_13892,N_13038,N_13096);
nor U13893 (N_13893,N_13367,N_13051);
nand U13894 (N_13894,N_13453,N_13122);
nand U13895 (N_13895,N_13481,N_13254);
and U13896 (N_13896,N_13374,N_13007);
xnor U13897 (N_13897,N_13098,N_13489);
and U13898 (N_13898,N_13456,N_13140);
xor U13899 (N_13899,N_13225,N_13463);
nor U13900 (N_13900,N_13119,N_13189);
or U13901 (N_13901,N_13271,N_13261);
xnor U13902 (N_13902,N_13132,N_13304);
nand U13903 (N_13903,N_13177,N_13343);
nand U13904 (N_13904,N_13318,N_13255);
nand U13905 (N_13905,N_13134,N_13413);
nand U13906 (N_13906,N_13359,N_13270);
or U13907 (N_13907,N_13420,N_13092);
nor U13908 (N_13908,N_13092,N_13238);
nand U13909 (N_13909,N_13237,N_13440);
xnor U13910 (N_13910,N_13494,N_13249);
xor U13911 (N_13911,N_13299,N_13456);
and U13912 (N_13912,N_13466,N_13323);
or U13913 (N_13913,N_13389,N_13051);
nor U13914 (N_13914,N_13026,N_13222);
or U13915 (N_13915,N_13145,N_13003);
xor U13916 (N_13916,N_13361,N_13098);
xor U13917 (N_13917,N_13033,N_13442);
nor U13918 (N_13918,N_13482,N_13046);
xor U13919 (N_13919,N_13261,N_13017);
nand U13920 (N_13920,N_13228,N_13285);
xor U13921 (N_13921,N_13390,N_13300);
nor U13922 (N_13922,N_13437,N_13029);
and U13923 (N_13923,N_13014,N_13324);
and U13924 (N_13924,N_13191,N_13366);
xnor U13925 (N_13925,N_13408,N_13245);
nand U13926 (N_13926,N_13248,N_13282);
and U13927 (N_13927,N_13157,N_13483);
xnor U13928 (N_13928,N_13016,N_13120);
xnor U13929 (N_13929,N_13148,N_13012);
nand U13930 (N_13930,N_13305,N_13382);
or U13931 (N_13931,N_13115,N_13298);
and U13932 (N_13932,N_13008,N_13271);
nor U13933 (N_13933,N_13355,N_13416);
nor U13934 (N_13934,N_13471,N_13041);
or U13935 (N_13935,N_13442,N_13356);
or U13936 (N_13936,N_13266,N_13371);
nand U13937 (N_13937,N_13366,N_13379);
and U13938 (N_13938,N_13363,N_13432);
nand U13939 (N_13939,N_13413,N_13327);
nor U13940 (N_13940,N_13452,N_13184);
xor U13941 (N_13941,N_13225,N_13145);
or U13942 (N_13942,N_13040,N_13444);
and U13943 (N_13943,N_13237,N_13408);
and U13944 (N_13944,N_13461,N_13289);
xnor U13945 (N_13945,N_13096,N_13418);
nand U13946 (N_13946,N_13184,N_13432);
nand U13947 (N_13947,N_13023,N_13228);
or U13948 (N_13948,N_13185,N_13408);
or U13949 (N_13949,N_13042,N_13136);
or U13950 (N_13950,N_13124,N_13418);
or U13951 (N_13951,N_13231,N_13152);
nor U13952 (N_13952,N_13387,N_13445);
or U13953 (N_13953,N_13303,N_13019);
nor U13954 (N_13954,N_13036,N_13202);
xnor U13955 (N_13955,N_13132,N_13237);
or U13956 (N_13956,N_13351,N_13406);
xor U13957 (N_13957,N_13043,N_13209);
xnor U13958 (N_13958,N_13103,N_13280);
and U13959 (N_13959,N_13434,N_13135);
and U13960 (N_13960,N_13014,N_13242);
and U13961 (N_13961,N_13046,N_13296);
xor U13962 (N_13962,N_13050,N_13312);
xnor U13963 (N_13963,N_13030,N_13234);
nor U13964 (N_13964,N_13167,N_13315);
nor U13965 (N_13965,N_13486,N_13234);
or U13966 (N_13966,N_13109,N_13251);
nor U13967 (N_13967,N_13252,N_13204);
xor U13968 (N_13968,N_13458,N_13310);
nand U13969 (N_13969,N_13246,N_13217);
xnor U13970 (N_13970,N_13157,N_13198);
or U13971 (N_13971,N_13308,N_13440);
nand U13972 (N_13972,N_13045,N_13061);
or U13973 (N_13973,N_13188,N_13198);
xor U13974 (N_13974,N_13107,N_13264);
nor U13975 (N_13975,N_13005,N_13477);
nand U13976 (N_13976,N_13244,N_13236);
or U13977 (N_13977,N_13466,N_13369);
or U13978 (N_13978,N_13165,N_13366);
and U13979 (N_13979,N_13256,N_13396);
nor U13980 (N_13980,N_13384,N_13020);
nor U13981 (N_13981,N_13074,N_13028);
xnor U13982 (N_13982,N_13187,N_13454);
nor U13983 (N_13983,N_13148,N_13310);
nand U13984 (N_13984,N_13337,N_13334);
nand U13985 (N_13985,N_13216,N_13336);
xnor U13986 (N_13986,N_13085,N_13435);
and U13987 (N_13987,N_13283,N_13241);
and U13988 (N_13988,N_13173,N_13001);
xor U13989 (N_13989,N_13074,N_13083);
xor U13990 (N_13990,N_13196,N_13043);
and U13991 (N_13991,N_13346,N_13284);
or U13992 (N_13992,N_13290,N_13323);
xor U13993 (N_13993,N_13044,N_13474);
xor U13994 (N_13994,N_13201,N_13048);
xnor U13995 (N_13995,N_13452,N_13256);
nand U13996 (N_13996,N_13207,N_13085);
xnor U13997 (N_13997,N_13099,N_13084);
nand U13998 (N_13998,N_13409,N_13174);
nand U13999 (N_13999,N_13453,N_13098);
nand U14000 (N_14000,N_13897,N_13537);
and U14001 (N_14001,N_13981,N_13994);
nor U14002 (N_14002,N_13977,N_13590);
and U14003 (N_14003,N_13786,N_13561);
or U14004 (N_14004,N_13796,N_13920);
or U14005 (N_14005,N_13598,N_13885);
nand U14006 (N_14006,N_13696,N_13926);
or U14007 (N_14007,N_13705,N_13925);
xor U14008 (N_14008,N_13556,N_13616);
or U14009 (N_14009,N_13749,N_13686);
and U14010 (N_14010,N_13575,N_13778);
xnor U14011 (N_14011,N_13916,N_13985);
and U14012 (N_14012,N_13924,N_13941);
nor U14013 (N_14013,N_13738,N_13852);
nand U14014 (N_14014,N_13634,N_13784);
xor U14015 (N_14015,N_13624,N_13583);
nand U14016 (N_14016,N_13503,N_13798);
and U14017 (N_14017,N_13806,N_13727);
xnor U14018 (N_14018,N_13544,N_13639);
and U14019 (N_14019,N_13965,N_13815);
or U14020 (N_14020,N_13578,N_13695);
and U14021 (N_14021,N_13528,N_13619);
and U14022 (N_14022,N_13701,N_13501);
nand U14023 (N_14023,N_13819,N_13911);
or U14024 (N_14024,N_13551,N_13703);
nand U14025 (N_14025,N_13874,N_13827);
xor U14026 (N_14026,N_13771,N_13859);
or U14027 (N_14027,N_13998,N_13972);
or U14028 (N_14028,N_13567,N_13524);
xnor U14029 (N_14029,N_13765,N_13564);
nand U14030 (N_14030,N_13900,N_13987);
nand U14031 (N_14031,N_13950,N_13902);
nand U14032 (N_14032,N_13877,N_13582);
or U14033 (N_14033,N_13767,N_13881);
or U14034 (N_14034,N_13893,N_13631);
nor U14035 (N_14035,N_13657,N_13795);
nor U14036 (N_14036,N_13706,N_13645);
or U14037 (N_14037,N_13870,N_13535);
nor U14038 (N_14038,N_13814,N_13579);
nor U14039 (N_14039,N_13646,N_13605);
nand U14040 (N_14040,N_13527,N_13975);
or U14041 (N_14041,N_13770,N_13895);
xnor U14042 (N_14042,N_13500,N_13937);
xnor U14043 (N_14043,N_13680,N_13983);
or U14044 (N_14044,N_13662,N_13620);
nor U14045 (N_14045,N_13709,N_13607);
or U14046 (N_14046,N_13737,N_13540);
nor U14047 (N_14047,N_13943,N_13871);
and U14048 (N_14048,N_13628,N_13692);
and U14049 (N_14049,N_13946,N_13808);
and U14050 (N_14050,N_13775,N_13515);
or U14051 (N_14051,N_13860,N_13802);
or U14052 (N_14052,N_13614,N_13728);
nand U14053 (N_14053,N_13674,N_13685);
or U14054 (N_14054,N_13514,N_13650);
and U14055 (N_14055,N_13894,N_13682);
xor U14056 (N_14056,N_13595,N_13876);
or U14057 (N_14057,N_13826,N_13840);
nand U14058 (N_14058,N_13714,N_13967);
nor U14059 (N_14059,N_13785,N_13707);
xnor U14060 (N_14060,N_13831,N_13512);
nand U14061 (N_14061,N_13821,N_13875);
nand U14062 (N_14062,N_13841,N_13764);
or U14063 (N_14063,N_13508,N_13603);
xnor U14064 (N_14064,N_13675,N_13918);
and U14065 (N_14065,N_13612,N_13606);
nand U14066 (N_14066,N_13930,N_13807);
or U14067 (N_14067,N_13577,N_13873);
nand U14068 (N_14068,N_13995,N_13823);
nor U14069 (N_14069,N_13659,N_13847);
nor U14070 (N_14070,N_13539,N_13947);
or U14071 (N_14071,N_13790,N_13687);
or U14072 (N_14072,N_13792,N_13836);
xor U14073 (N_14073,N_13519,N_13812);
xnor U14074 (N_14074,N_13867,N_13759);
xnor U14075 (N_14075,N_13825,N_13751);
xor U14076 (N_14076,N_13776,N_13622);
nand U14077 (N_14077,N_13664,N_13934);
or U14078 (N_14078,N_13923,N_13525);
xnor U14079 (N_14079,N_13509,N_13518);
or U14080 (N_14080,N_13691,N_13677);
nand U14081 (N_14081,N_13810,N_13978);
or U14082 (N_14082,N_13948,N_13780);
xnor U14083 (N_14083,N_13991,N_13699);
or U14084 (N_14084,N_13627,N_13963);
nand U14085 (N_14085,N_13853,N_13794);
or U14086 (N_14086,N_13681,N_13846);
and U14087 (N_14087,N_13960,N_13640);
nor U14088 (N_14088,N_13604,N_13654);
or U14089 (N_14089,N_13732,N_13625);
or U14090 (N_14090,N_13623,N_13666);
or U14091 (N_14091,N_13953,N_13610);
nand U14092 (N_14092,N_13572,N_13964);
nor U14093 (N_14093,N_13955,N_13736);
xnor U14094 (N_14094,N_13858,N_13855);
and U14095 (N_14095,N_13854,N_13717);
xnor U14096 (N_14096,N_13884,N_13660);
or U14097 (N_14097,N_13891,N_13915);
nand U14098 (N_14098,N_13734,N_13904);
or U14099 (N_14099,N_13754,N_13626);
xor U14100 (N_14100,N_13928,N_13538);
and U14101 (N_14101,N_13559,N_13907);
or U14102 (N_14102,N_13718,N_13988);
or U14103 (N_14103,N_13601,N_13574);
nand U14104 (N_14104,N_13615,N_13944);
nor U14105 (N_14105,N_13850,N_13550);
nand U14106 (N_14106,N_13589,N_13993);
nand U14107 (N_14107,N_13848,N_13952);
or U14108 (N_14108,N_13642,N_13849);
nand U14109 (N_14109,N_13880,N_13912);
xor U14110 (N_14110,N_13684,N_13688);
nand U14111 (N_14111,N_13762,N_13839);
xnor U14112 (N_14112,N_13745,N_13800);
or U14113 (N_14113,N_13581,N_13708);
nand U14114 (N_14114,N_13989,N_13868);
xor U14115 (N_14115,N_13635,N_13648);
and U14116 (N_14116,N_13571,N_13979);
nor U14117 (N_14117,N_13511,N_13788);
and U14118 (N_14118,N_13502,N_13750);
and U14119 (N_14119,N_13643,N_13939);
nand U14120 (N_14120,N_13742,N_13676);
nand U14121 (N_14121,N_13609,N_13747);
or U14122 (N_14122,N_13730,N_13986);
and U14123 (N_14123,N_13921,N_13898);
nand U14124 (N_14124,N_13824,N_13663);
and U14125 (N_14125,N_13956,N_13722);
nor U14126 (N_14126,N_13938,N_13633);
xnor U14127 (N_14127,N_13629,N_13689);
xnor U14128 (N_14128,N_13534,N_13698);
or U14129 (N_14129,N_13553,N_13670);
or U14130 (N_14130,N_13565,N_13573);
or U14131 (N_14131,N_13748,N_13593);
xnor U14132 (N_14132,N_13996,N_13818);
nand U14133 (N_14133,N_13910,N_13618);
nor U14134 (N_14134,N_13720,N_13638);
nand U14135 (N_14135,N_13513,N_13545);
nand U14136 (N_14136,N_13673,N_13845);
and U14137 (N_14137,N_13542,N_13892);
or U14138 (N_14138,N_13617,N_13526);
nor U14139 (N_14139,N_13562,N_13782);
nor U14140 (N_14140,N_13984,N_13769);
xnor U14141 (N_14141,N_13655,N_13768);
and U14142 (N_14142,N_13822,N_13594);
or U14143 (N_14143,N_13585,N_13844);
and U14144 (N_14144,N_13935,N_13777);
and U14145 (N_14145,N_13863,N_13940);
nor U14146 (N_14146,N_13861,N_13725);
or U14147 (N_14147,N_13766,N_13611);
nor U14148 (N_14148,N_13908,N_13668);
xor U14149 (N_14149,N_13731,N_13715);
and U14150 (N_14150,N_13733,N_13922);
and U14151 (N_14151,N_13557,N_13890);
nand U14152 (N_14152,N_13584,N_13679);
nand U14153 (N_14153,N_13596,N_13957);
and U14154 (N_14154,N_13805,N_13905);
nor U14155 (N_14155,N_13530,N_13971);
xnor U14156 (N_14156,N_13746,N_13903);
and U14157 (N_14157,N_13803,N_13813);
nand U14158 (N_14158,N_13866,N_13969);
and U14159 (N_14159,N_13569,N_13997);
or U14160 (N_14160,N_13931,N_13644);
xor U14161 (N_14161,N_13529,N_13586);
nand U14162 (N_14162,N_13774,N_13832);
xnor U14163 (N_14163,N_13543,N_13933);
nor U14164 (N_14164,N_13828,N_13563);
or U14165 (N_14165,N_13758,N_13879);
and U14166 (N_14166,N_13756,N_13830);
nand U14167 (N_14167,N_13882,N_13787);
xnor U14168 (N_14168,N_13917,N_13761);
and U14169 (N_14169,N_13906,N_13547);
nor U14170 (N_14170,N_13864,N_13962);
nor U14171 (N_14171,N_13945,N_13667);
nor U14172 (N_14172,N_13773,N_13954);
or U14173 (N_14173,N_13752,N_13653);
or U14174 (N_14174,N_13541,N_13697);
and U14175 (N_14175,N_13783,N_13506);
or U14176 (N_14176,N_13741,N_13932);
or U14177 (N_14177,N_13560,N_13702);
xor U14178 (N_14178,N_13704,N_13942);
nand U14179 (N_14179,N_13713,N_13743);
and U14180 (N_14180,N_13936,N_13723);
xor U14181 (N_14181,N_13763,N_13592);
xnor U14182 (N_14182,N_13729,N_13558);
nand U14183 (N_14183,N_13816,N_13966);
nor U14184 (N_14184,N_13716,N_13973);
and U14185 (N_14185,N_13672,N_13974);
nor U14186 (N_14186,N_13833,N_13656);
and U14187 (N_14187,N_13929,N_13883);
nand U14188 (N_14188,N_13522,N_13982);
or U14189 (N_14189,N_13834,N_13505);
and U14190 (N_14190,N_13869,N_13789);
or U14191 (N_14191,N_13533,N_13641);
nand U14192 (N_14192,N_13878,N_13914);
nand U14193 (N_14193,N_13711,N_13548);
xor U14194 (N_14194,N_13842,N_13817);
nor U14195 (N_14195,N_13901,N_13968);
xor U14196 (N_14196,N_13896,N_13552);
nor U14197 (N_14197,N_13630,N_13600);
xnor U14198 (N_14198,N_13566,N_13724);
nor U14199 (N_14199,N_13909,N_13531);
xor U14200 (N_14200,N_13652,N_13857);
and U14201 (N_14201,N_13793,N_13632);
xnor U14202 (N_14202,N_13521,N_13886);
xnor U14203 (N_14203,N_13719,N_13959);
nand U14204 (N_14204,N_13507,N_13591);
nand U14205 (N_14205,N_13700,N_13951);
and U14206 (N_14206,N_13851,N_13580);
nand U14207 (N_14207,N_13837,N_13888);
nor U14208 (N_14208,N_13608,N_13549);
or U14209 (N_14209,N_13576,N_13781);
and U14210 (N_14210,N_13669,N_13791);
nor U14211 (N_14211,N_13637,N_13694);
nor U14212 (N_14212,N_13970,N_13801);
nand U14213 (N_14213,N_13913,N_13690);
nand U14214 (N_14214,N_13990,N_13961);
nor U14215 (N_14215,N_13510,N_13865);
xor U14216 (N_14216,N_13744,N_13532);
nor U14217 (N_14217,N_13602,N_13712);
xor U14218 (N_14218,N_13889,N_13799);
and U14219 (N_14219,N_13710,N_13651);
nor U14220 (N_14220,N_13887,N_13588);
xnor U14221 (N_14221,N_13862,N_13980);
xor U14222 (N_14222,N_13999,N_13992);
nor U14223 (N_14223,N_13809,N_13899);
and U14224 (N_14224,N_13504,N_13658);
nand U14225 (N_14225,N_13678,N_13760);
xnor U14226 (N_14226,N_13523,N_13843);
nor U14227 (N_14227,N_13721,N_13958);
or U14228 (N_14228,N_13683,N_13735);
and U14229 (N_14229,N_13621,N_13647);
or U14230 (N_14230,N_13753,N_13976);
nor U14231 (N_14231,N_13740,N_13856);
and U14232 (N_14232,N_13726,N_13927);
xnor U14233 (N_14233,N_13554,N_13546);
xor U14234 (N_14234,N_13599,N_13804);
nand U14235 (N_14235,N_13536,N_13636);
or U14236 (N_14236,N_13665,N_13820);
nand U14237 (N_14237,N_13516,N_13661);
nand U14238 (N_14238,N_13693,N_13587);
xnor U14239 (N_14239,N_13772,N_13829);
xnor U14240 (N_14240,N_13649,N_13520);
and U14241 (N_14241,N_13811,N_13919);
xnor U14242 (N_14242,N_13517,N_13671);
or U14243 (N_14243,N_13739,N_13872);
nand U14244 (N_14244,N_13555,N_13597);
or U14245 (N_14245,N_13757,N_13949);
or U14246 (N_14246,N_13570,N_13797);
or U14247 (N_14247,N_13755,N_13613);
or U14248 (N_14248,N_13838,N_13835);
nor U14249 (N_14249,N_13779,N_13568);
nand U14250 (N_14250,N_13645,N_13826);
nand U14251 (N_14251,N_13906,N_13988);
nand U14252 (N_14252,N_13923,N_13563);
nand U14253 (N_14253,N_13919,N_13845);
xnor U14254 (N_14254,N_13862,N_13647);
and U14255 (N_14255,N_13867,N_13897);
nor U14256 (N_14256,N_13563,N_13953);
nand U14257 (N_14257,N_13945,N_13956);
nor U14258 (N_14258,N_13987,N_13953);
and U14259 (N_14259,N_13725,N_13696);
nand U14260 (N_14260,N_13824,N_13863);
xnor U14261 (N_14261,N_13834,N_13634);
and U14262 (N_14262,N_13817,N_13677);
and U14263 (N_14263,N_13909,N_13798);
xor U14264 (N_14264,N_13946,N_13889);
nor U14265 (N_14265,N_13878,N_13783);
and U14266 (N_14266,N_13836,N_13972);
xor U14267 (N_14267,N_13848,N_13522);
and U14268 (N_14268,N_13692,N_13958);
nor U14269 (N_14269,N_13602,N_13708);
and U14270 (N_14270,N_13667,N_13773);
or U14271 (N_14271,N_13892,N_13706);
xor U14272 (N_14272,N_13831,N_13640);
nand U14273 (N_14273,N_13854,N_13543);
xor U14274 (N_14274,N_13842,N_13787);
or U14275 (N_14275,N_13891,N_13770);
and U14276 (N_14276,N_13831,N_13634);
xnor U14277 (N_14277,N_13634,N_13931);
or U14278 (N_14278,N_13815,N_13945);
nor U14279 (N_14279,N_13692,N_13630);
nor U14280 (N_14280,N_13535,N_13869);
xor U14281 (N_14281,N_13837,N_13504);
xor U14282 (N_14282,N_13973,N_13622);
and U14283 (N_14283,N_13842,N_13758);
xnor U14284 (N_14284,N_13566,N_13667);
nor U14285 (N_14285,N_13886,N_13795);
xnor U14286 (N_14286,N_13910,N_13678);
and U14287 (N_14287,N_13949,N_13538);
xnor U14288 (N_14288,N_13679,N_13761);
xnor U14289 (N_14289,N_13929,N_13529);
xnor U14290 (N_14290,N_13559,N_13948);
or U14291 (N_14291,N_13951,N_13548);
xnor U14292 (N_14292,N_13747,N_13969);
and U14293 (N_14293,N_13973,N_13647);
xnor U14294 (N_14294,N_13627,N_13816);
xor U14295 (N_14295,N_13930,N_13603);
nand U14296 (N_14296,N_13588,N_13626);
nand U14297 (N_14297,N_13654,N_13973);
nand U14298 (N_14298,N_13941,N_13609);
nor U14299 (N_14299,N_13785,N_13529);
or U14300 (N_14300,N_13755,N_13629);
nor U14301 (N_14301,N_13680,N_13884);
and U14302 (N_14302,N_13831,N_13825);
or U14303 (N_14303,N_13735,N_13632);
xnor U14304 (N_14304,N_13621,N_13501);
or U14305 (N_14305,N_13811,N_13761);
nor U14306 (N_14306,N_13909,N_13544);
xor U14307 (N_14307,N_13630,N_13966);
or U14308 (N_14308,N_13713,N_13829);
xnor U14309 (N_14309,N_13529,N_13927);
nand U14310 (N_14310,N_13577,N_13607);
nor U14311 (N_14311,N_13533,N_13871);
or U14312 (N_14312,N_13655,N_13507);
and U14313 (N_14313,N_13961,N_13756);
or U14314 (N_14314,N_13620,N_13982);
or U14315 (N_14315,N_13992,N_13780);
xnor U14316 (N_14316,N_13942,N_13533);
and U14317 (N_14317,N_13684,N_13830);
or U14318 (N_14318,N_13892,N_13523);
xnor U14319 (N_14319,N_13700,N_13822);
or U14320 (N_14320,N_13768,N_13639);
xor U14321 (N_14321,N_13954,N_13673);
xor U14322 (N_14322,N_13973,N_13725);
xnor U14323 (N_14323,N_13655,N_13964);
xnor U14324 (N_14324,N_13826,N_13531);
nand U14325 (N_14325,N_13929,N_13918);
or U14326 (N_14326,N_13964,N_13843);
nor U14327 (N_14327,N_13634,N_13891);
and U14328 (N_14328,N_13622,N_13603);
or U14329 (N_14329,N_13673,N_13984);
xnor U14330 (N_14330,N_13571,N_13761);
or U14331 (N_14331,N_13500,N_13711);
xor U14332 (N_14332,N_13725,N_13947);
nor U14333 (N_14333,N_13500,N_13808);
nand U14334 (N_14334,N_13583,N_13598);
nor U14335 (N_14335,N_13833,N_13612);
nor U14336 (N_14336,N_13606,N_13593);
xnor U14337 (N_14337,N_13758,N_13812);
nor U14338 (N_14338,N_13537,N_13651);
nor U14339 (N_14339,N_13890,N_13729);
or U14340 (N_14340,N_13922,N_13984);
nor U14341 (N_14341,N_13970,N_13996);
and U14342 (N_14342,N_13945,N_13599);
or U14343 (N_14343,N_13636,N_13692);
xnor U14344 (N_14344,N_13951,N_13667);
nand U14345 (N_14345,N_13728,N_13940);
xor U14346 (N_14346,N_13798,N_13910);
and U14347 (N_14347,N_13500,N_13964);
xnor U14348 (N_14348,N_13953,N_13753);
nand U14349 (N_14349,N_13502,N_13794);
nor U14350 (N_14350,N_13597,N_13846);
nand U14351 (N_14351,N_13778,N_13963);
and U14352 (N_14352,N_13620,N_13892);
and U14353 (N_14353,N_13605,N_13559);
or U14354 (N_14354,N_13533,N_13863);
nor U14355 (N_14355,N_13779,N_13860);
xnor U14356 (N_14356,N_13749,N_13950);
xor U14357 (N_14357,N_13869,N_13913);
or U14358 (N_14358,N_13884,N_13525);
nand U14359 (N_14359,N_13740,N_13712);
xor U14360 (N_14360,N_13539,N_13580);
and U14361 (N_14361,N_13726,N_13784);
nand U14362 (N_14362,N_13525,N_13654);
and U14363 (N_14363,N_13783,N_13581);
and U14364 (N_14364,N_13616,N_13905);
or U14365 (N_14365,N_13716,N_13894);
and U14366 (N_14366,N_13659,N_13985);
and U14367 (N_14367,N_13729,N_13936);
and U14368 (N_14368,N_13519,N_13904);
or U14369 (N_14369,N_13511,N_13924);
nand U14370 (N_14370,N_13882,N_13960);
nor U14371 (N_14371,N_13884,N_13873);
nor U14372 (N_14372,N_13998,N_13729);
or U14373 (N_14373,N_13725,N_13785);
nand U14374 (N_14374,N_13582,N_13870);
xor U14375 (N_14375,N_13677,N_13946);
nand U14376 (N_14376,N_13721,N_13797);
and U14377 (N_14377,N_13781,N_13881);
xor U14378 (N_14378,N_13805,N_13646);
or U14379 (N_14379,N_13596,N_13920);
or U14380 (N_14380,N_13741,N_13638);
nand U14381 (N_14381,N_13758,N_13685);
xor U14382 (N_14382,N_13800,N_13521);
and U14383 (N_14383,N_13641,N_13767);
or U14384 (N_14384,N_13930,N_13861);
and U14385 (N_14385,N_13763,N_13583);
and U14386 (N_14386,N_13990,N_13559);
nand U14387 (N_14387,N_13688,N_13786);
xnor U14388 (N_14388,N_13694,N_13865);
xor U14389 (N_14389,N_13684,N_13827);
nand U14390 (N_14390,N_13718,N_13587);
xor U14391 (N_14391,N_13575,N_13809);
nor U14392 (N_14392,N_13911,N_13691);
nand U14393 (N_14393,N_13999,N_13649);
nand U14394 (N_14394,N_13831,N_13851);
xor U14395 (N_14395,N_13562,N_13987);
xnor U14396 (N_14396,N_13815,N_13882);
and U14397 (N_14397,N_13788,N_13931);
nand U14398 (N_14398,N_13877,N_13947);
nand U14399 (N_14399,N_13834,N_13504);
xnor U14400 (N_14400,N_13843,N_13660);
nand U14401 (N_14401,N_13810,N_13723);
or U14402 (N_14402,N_13932,N_13679);
nor U14403 (N_14403,N_13914,N_13655);
or U14404 (N_14404,N_13717,N_13882);
nor U14405 (N_14405,N_13750,N_13877);
xor U14406 (N_14406,N_13929,N_13783);
nor U14407 (N_14407,N_13973,N_13926);
xor U14408 (N_14408,N_13501,N_13616);
nor U14409 (N_14409,N_13988,N_13885);
xnor U14410 (N_14410,N_13595,N_13811);
nor U14411 (N_14411,N_13611,N_13699);
xnor U14412 (N_14412,N_13973,N_13861);
and U14413 (N_14413,N_13630,N_13737);
nand U14414 (N_14414,N_13642,N_13937);
xnor U14415 (N_14415,N_13822,N_13705);
nand U14416 (N_14416,N_13929,N_13894);
nor U14417 (N_14417,N_13712,N_13835);
or U14418 (N_14418,N_13887,N_13737);
or U14419 (N_14419,N_13773,N_13586);
xnor U14420 (N_14420,N_13806,N_13534);
nand U14421 (N_14421,N_13725,N_13660);
xnor U14422 (N_14422,N_13523,N_13681);
xnor U14423 (N_14423,N_13829,N_13584);
or U14424 (N_14424,N_13866,N_13709);
nand U14425 (N_14425,N_13836,N_13885);
and U14426 (N_14426,N_13635,N_13538);
xnor U14427 (N_14427,N_13573,N_13533);
nor U14428 (N_14428,N_13883,N_13764);
or U14429 (N_14429,N_13717,N_13808);
nand U14430 (N_14430,N_13907,N_13793);
xor U14431 (N_14431,N_13646,N_13806);
nand U14432 (N_14432,N_13719,N_13916);
or U14433 (N_14433,N_13699,N_13609);
xor U14434 (N_14434,N_13514,N_13895);
nor U14435 (N_14435,N_13950,N_13650);
or U14436 (N_14436,N_13828,N_13835);
or U14437 (N_14437,N_13701,N_13649);
and U14438 (N_14438,N_13539,N_13642);
nand U14439 (N_14439,N_13668,N_13547);
xor U14440 (N_14440,N_13919,N_13694);
nand U14441 (N_14441,N_13500,N_13876);
nor U14442 (N_14442,N_13768,N_13727);
and U14443 (N_14443,N_13683,N_13990);
or U14444 (N_14444,N_13717,N_13832);
xnor U14445 (N_14445,N_13654,N_13531);
xor U14446 (N_14446,N_13663,N_13768);
xor U14447 (N_14447,N_13613,N_13937);
xnor U14448 (N_14448,N_13619,N_13554);
nor U14449 (N_14449,N_13578,N_13819);
and U14450 (N_14450,N_13975,N_13726);
nand U14451 (N_14451,N_13889,N_13873);
nor U14452 (N_14452,N_13664,N_13860);
nand U14453 (N_14453,N_13662,N_13905);
nand U14454 (N_14454,N_13932,N_13738);
or U14455 (N_14455,N_13596,N_13603);
and U14456 (N_14456,N_13579,N_13652);
or U14457 (N_14457,N_13568,N_13862);
or U14458 (N_14458,N_13555,N_13544);
xor U14459 (N_14459,N_13727,N_13918);
xor U14460 (N_14460,N_13665,N_13831);
xnor U14461 (N_14461,N_13738,N_13854);
xor U14462 (N_14462,N_13640,N_13704);
or U14463 (N_14463,N_13571,N_13607);
nor U14464 (N_14464,N_13877,N_13662);
nand U14465 (N_14465,N_13977,N_13843);
xor U14466 (N_14466,N_13873,N_13511);
and U14467 (N_14467,N_13745,N_13695);
and U14468 (N_14468,N_13863,N_13967);
or U14469 (N_14469,N_13663,N_13559);
nor U14470 (N_14470,N_13886,N_13542);
or U14471 (N_14471,N_13608,N_13984);
nand U14472 (N_14472,N_13815,N_13537);
nand U14473 (N_14473,N_13700,N_13792);
and U14474 (N_14474,N_13872,N_13614);
and U14475 (N_14475,N_13697,N_13858);
nand U14476 (N_14476,N_13812,N_13596);
or U14477 (N_14477,N_13887,N_13550);
and U14478 (N_14478,N_13684,N_13897);
or U14479 (N_14479,N_13834,N_13873);
or U14480 (N_14480,N_13712,N_13542);
or U14481 (N_14481,N_13939,N_13514);
and U14482 (N_14482,N_13523,N_13822);
and U14483 (N_14483,N_13752,N_13595);
nand U14484 (N_14484,N_13965,N_13574);
or U14485 (N_14485,N_13894,N_13949);
nor U14486 (N_14486,N_13585,N_13759);
nand U14487 (N_14487,N_13579,N_13687);
nor U14488 (N_14488,N_13835,N_13646);
nand U14489 (N_14489,N_13674,N_13690);
nor U14490 (N_14490,N_13888,N_13660);
xnor U14491 (N_14491,N_13753,N_13754);
nor U14492 (N_14492,N_13502,N_13656);
and U14493 (N_14493,N_13645,N_13812);
nor U14494 (N_14494,N_13531,N_13894);
xnor U14495 (N_14495,N_13796,N_13695);
and U14496 (N_14496,N_13541,N_13749);
nor U14497 (N_14497,N_13905,N_13899);
or U14498 (N_14498,N_13990,N_13557);
or U14499 (N_14499,N_13691,N_13953);
nand U14500 (N_14500,N_14136,N_14013);
xor U14501 (N_14501,N_14321,N_14303);
and U14502 (N_14502,N_14102,N_14278);
and U14503 (N_14503,N_14298,N_14283);
or U14504 (N_14504,N_14490,N_14290);
and U14505 (N_14505,N_14109,N_14078);
or U14506 (N_14506,N_14235,N_14373);
nand U14507 (N_14507,N_14268,N_14436);
nor U14508 (N_14508,N_14020,N_14085);
xor U14509 (N_14509,N_14249,N_14306);
and U14510 (N_14510,N_14056,N_14291);
nand U14511 (N_14511,N_14000,N_14003);
nor U14512 (N_14512,N_14361,N_14089);
nor U14513 (N_14513,N_14417,N_14066);
nor U14514 (N_14514,N_14253,N_14051);
nand U14515 (N_14515,N_14449,N_14451);
nor U14516 (N_14516,N_14270,N_14391);
nand U14517 (N_14517,N_14299,N_14478);
xnor U14518 (N_14518,N_14316,N_14172);
nand U14519 (N_14519,N_14471,N_14009);
nand U14520 (N_14520,N_14080,N_14352);
or U14521 (N_14521,N_14222,N_14227);
or U14522 (N_14522,N_14395,N_14351);
and U14523 (N_14523,N_14138,N_14221);
or U14524 (N_14524,N_14468,N_14072);
nand U14525 (N_14525,N_14076,N_14384);
xnor U14526 (N_14526,N_14209,N_14036);
nor U14527 (N_14527,N_14021,N_14480);
and U14528 (N_14528,N_14068,N_14446);
or U14529 (N_14529,N_14210,N_14272);
or U14530 (N_14530,N_14444,N_14014);
nand U14531 (N_14531,N_14035,N_14063);
and U14532 (N_14532,N_14282,N_14314);
or U14533 (N_14533,N_14359,N_14263);
or U14534 (N_14534,N_14156,N_14028);
nor U14535 (N_14535,N_14019,N_14259);
or U14536 (N_14536,N_14079,N_14269);
nor U14537 (N_14537,N_14344,N_14192);
nand U14538 (N_14538,N_14034,N_14477);
nor U14539 (N_14539,N_14055,N_14470);
nand U14540 (N_14540,N_14482,N_14117);
and U14541 (N_14541,N_14201,N_14120);
xor U14542 (N_14542,N_14100,N_14419);
nand U14543 (N_14543,N_14140,N_14365);
and U14544 (N_14544,N_14440,N_14231);
nor U14545 (N_14545,N_14075,N_14010);
nand U14546 (N_14546,N_14129,N_14312);
or U14547 (N_14547,N_14145,N_14099);
and U14548 (N_14548,N_14062,N_14325);
or U14549 (N_14549,N_14105,N_14040);
xor U14550 (N_14550,N_14454,N_14179);
nor U14551 (N_14551,N_14159,N_14065);
nor U14552 (N_14552,N_14043,N_14354);
nand U14553 (N_14553,N_14012,N_14305);
and U14554 (N_14554,N_14264,N_14077);
and U14555 (N_14555,N_14252,N_14381);
nand U14556 (N_14556,N_14459,N_14465);
or U14557 (N_14557,N_14050,N_14185);
nor U14558 (N_14558,N_14377,N_14411);
nand U14559 (N_14559,N_14168,N_14489);
or U14560 (N_14560,N_14232,N_14111);
xnor U14561 (N_14561,N_14261,N_14341);
nor U14562 (N_14562,N_14154,N_14293);
xnor U14563 (N_14563,N_14097,N_14251);
and U14564 (N_14564,N_14127,N_14011);
nand U14565 (N_14565,N_14375,N_14432);
and U14566 (N_14566,N_14453,N_14132);
and U14567 (N_14567,N_14326,N_14474);
or U14568 (N_14568,N_14024,N_14498);
nor U14569 (N_14569,N_14216,N_14171);
or U14570 (N_14570,N_14318,N_14425);
xnor U14571 (N_14571,N_14170,N_14368);
xnor U14572 (N_14572,N_14492,N_14026);
xnor U14573 (N_14573,N_14193,N_14307);
xnor U14574 (N_14574,N_14379,N_14180);
nand U14575 (N_14575,N_14445,N_14484);
nand U14576 (N_14576,N_14485,N_14265);
nand U14577 (N_14577,N_14176,N_14023);
or U14578 (N_14578,N_14398,N_14096);
and U14579 (N_14579,N_14315,N_14336);
and U14580 (N_14580,N_14236,N_14048);
nor U14581 (N_14581,N_14133,N_14110);
xnor U14582 (N_14582,N_14281,N_14197);
nand U14583 (N_14583,N_14450,N_14430);
and U14584 (N_14584,N_14435,N_14181);
and U14585 (N_14585,N_14401,N_14456);
and U14586 (N_14586,N_14403,N_14289);
xor U14587 (N_14587,N_14311,N_14335);
or U14588 (N_14588,N_14428,N_14057);
xor U14589 (N_14589,N_14266,N_14362);
or U14590 (N_14590,N_14390,N_14328);
xor U14591 (N_14591,N_14383,N_14422);
nor U14592 (N_14592,N_14286,N_14412);
and U14593 (N_14593,N_14487,N_14092);
nand U14594 (N_14594,N_14112,N_14413);
nand U14595 (N_14595,N_14360,N_14386);
or U14596 (N_14596,N_14346,N_14084);
or U14597 (N_14597,N_14073,N_14276);
xnor U14598 (N_14598,N_14190,N_14044);
and U14599 (N_14599,N_14329,N_14349);
or U14600 (N_14600,N_14423,N_14150);
xor U14601 (N_14601,N_14439,N_14144);
or U14602 (N_14602,N_14108,N_14217);
or U14603 (N_14603,N_14095,N_14322);
and U14604 (N_14604,N_14483,N_14228);
xnor U14605 (N_14605,N_14119,N_14205);
xnor U14606 (N_14606,N_14256,N_14388);
and U14607 (N_14607,N_14015,N_14158);
xnor U14608 (N_14608,N_14402,N_14017);
nor U14609 (N_14609,N_14189,N_14218);
nand U14610 (N_14610,N_14183,N_14476);
xnor U14611 (N_14611,N_14199,N_14142);
or U14612 (N_14612,N_14300,N_14196);
and U14613 (N_14613,N_14016,N_14162);
nor U14614 (N_14614,N_14247,N_14397);
nor U14615 (N_14615,N_14018,N_14271);
nand U14616 (N_14616,N_14086,N_14358);
nand U14617 (N_14617,N_14087,N_14031);
nand U14618 (N_14618,N_14047,N_14284);
xor U14619 (N_14619,N_14022,N_14125);
or U14620 (N_14620,N_14455,N_14025);
nand U14621 (N_14621,N_14369,N_14037);
or U14622 (N_14622,N_14155,N_14338);
or U14623 (N_14623,N_14363,N_14103);
or U14624 (N_14624,N_14319,N_14098);
nor U14625 (N_14625,N_14239,N_14128);
and U14626 (N_14626,N_14320,N_14039);
nor U14627 (N_14627,N_14131,N_14491);
or U14628 (N_14628,N_14118,N_14163);
xor U14629 (N_14629,N_14473,N_14400);
and U14630 (N_14630,N_14121,N_14134);
nand U14631 (N_14631,N_14246,N_14030);
nor U14632 (N_14632,N_14313,N_14149);
and U14633 (N_14633,N_14059,N_14195);
and U14634 (N_14634,N_14241,N_14052);
or U14635 (N_14635,N_14409,N_14093);
nor U14636 (N_14636,N_14090,N_14370);
nor U14637 (N_14637,N_14333,N_14153);
xor U14638 (N_14638,N_14211,N_14257);
nor U14639 (N_14639,N_14135,N_14467);
or U14640 (N_14640,N_14174,N_14466);
nor U14641 (N_14641,N_14464,N_14296);
nor U14642 (N_14642,N_14255,N_14394);
nor U14643 (N_14643,N_14137,N_14045);
or U14644 (N_14644,N_14304,N_14160);
and U14645 (N_14645,N_14273,N_14214);
xnor U14646 (N_14646,N_14353,N_14187);
or U14647 (N_14647,N_14324,N_14122);
nor U14648 (N_14648,N_14165,N_14007);
nand U14649 (N_14649,N_14206,N_14238);
xor U14650 (N_14650,N_14294,N_14405);
and U14651 (N_14651,N_14433,N_14173);
or U14652 (N_14652,N_14237,N_14130);
or U14653 (N_14653,N_14475,N_14058);
xor U14654 (N_14654,N_14069,N_14385);
nor U14655 (N_14655,N_14393,N_14429);
or U14656 (N_14656,N_14458,N_14207);
xnor U14657 (N_14657,N_14447,N_14027);
xor U14658 (N_14658,N_14461,N_14177);
nor U14659 (N_14659,N_14469,N_14443);
or U14660 (N_14660,N_14060,N_14399);
or U14661 (N_14661,N_14107,N_14343);
or U14662 (N_14662,N_14410,N_14226);
xnor U14663 (N_14663,N_14033,N_14038);
and U14664 (N_14664,N_14230,N_14175);
and U14665 (N_14665,N_14215,N_14242);
nand U14666 (N_14666,N_14442,N_14094);
nor U14667 (N_14667,N_14054,N_14345);
xnor U14668 (N_14668,N_14167,N_14248);
nor U14669 (N_14669,N_14371,N_14146);
or U14670 (N_14670,N_14441,N_14437);
and U14671 (N_14671,N_14367,N_14389);
or U14672 (N_14672,N_14148,N_14332);
nand U14673 (N_14673,N_14355,N_14295);
nor U14674 (N_14674,N_14041,N_14151);
nor U14675 (N_14675,N_14074,N_14113);
or U14676 (N_14676,N_14223,N_14481);
or U14677 (N_14677,N_14347,N_14274);
and U14678 (N_14678,N_14225,N_14002);
nand U14679 (N_14679,N_14188,N_14277);
xor U14680 (N_14680,N_14292,N_14364);
xnor U14681 (N_14681,N_14004,N_14166);
nor U14682 (N_14682,N_14310,N_14082);
and U14683 (N_14683,N_14184,N_14123);
nand U14684 (N_14684,N_14067,N_14104);
nand U14685 (N_14685,N_14053,N_14488);
nor U14686 (N_14686,N_14460,N_14424);
nand U14687 (N_14687,N_14406,N_14331);
xnor U14688 (N_14688,N_14101,N_14418);
or U14689 (N_14689,N_14323,N_14380);
nand U14690 (N_14690,N_14233,N_14357);
nor U14691 (N_14691,N_14064,N_14486);
nor U14692 (N_14692,N_14126,N_14496);
and U14693 (N_14693,N_14438,N_14240);
or U14694 (N_14694,N_14414,N_14115);
xnor U14695 (N_14695,N_14139,N_14042);
nor U14696 (N_14696,N_14494,N_14356);
nand U14697 (N_14697,N_14285,N_14220);
nand U14698 (N_14698,N_14203,N_14194);
nand U14699 (N_14699,N_14279,N_14152);
nand U14700 (N_14700,N_14229,N_14254);
nor U14701 (N_14701,N_14260,N_14267);
nor U14702 (N_14702,N_14407,N_14415);
xor U14703 (N_14703,N_14071,N_14046);
and U14704 (N_14704,N_14262,N_14178);
nand U14705 (N_14705,N_14378,N_14392);
nand U14706 (N_14706,N_14308,N_14088);
nand U14707 (N_14707,N_14114,N_14182);
and U14708 (N_14708,N_14204,N_14499);
or U14709 (N_14709,N_14191,N_14427);
xnor U14710 (N_14710,N_14202,N_14061);
nand U14711 (N_14711,N_14337,N_14164);
or U14712 (N_14712,N_14029,N_14200);
xor U14713 (N_14713,N_14258,N_14081);
xor U14714 (N_14714,N_14387,N_14169);
or U14715 (N_14715,N_14334,N_14348);
nand U14716 (N_14716,N_14245,N_14124);
and U14717 (N_14717,N_14083,N_14366);
xor U14718 (N_14718,N_14161,N_14244);
and U14719 (N_14719,N_14141,N_14186);
xor U14720 (N_14720,N_14143,N_14049);
xor U14721 (N_14721,N_14434,N_14404);
nor U14722 (N_14722,N_14420,N_14495);
and U14723 (N_14723,N_14376,N_14287);
xnor U14724 (N_14724,N_14275,N_14250);
nor U14725 (N_14725,N_14339,N_14457);
or U14726 (N_14726,N_14479,N_14431);
or U14727 (N_14727,N_14208,N_14070);
nand U14728 (N_14728,N_14157,N_14374);
or U14729 (N_14729,N_14426,N_14005);
nor U14730 (N_14730,N_14032,N_14198);
nor U14731 (N_14731,N_14416,N_14212);
xor U14732 (N_14732,N_14116,N_14493);
nand U14733 (N_14733,N_14396,N_14309);
xnor U14734 (N_14734,N_14147,N_14301);
nor U14735 (N_14735,N_14421,N_14340);
or U14736 (N_14736,N_14234,N_14350);
and U14737 (N_14737,N_14327,N_14317);
or U14738 (N_14738,N_14302,N_14243);
nand U14739 (N_14739,N_14448,N_14280);
or U14740 (N_14740,N_14001,N_14342);
nor U14741 (N_14741,N_14408,N_14219);
nor U14742 (N_14742,N_14452,N_14091);
xnor U14743 (N_14743,N_14463,N_14497);
xnor U14744 (N_14744,N_14462,N_14224);
nor U14745 (N_14745,N_14006,N_14382);
nor U14746 (N_14746,N_14472,N_14297);
or U14747 (N_14747,N_14008,N_14372);
xnor U14748 (N_14748,N_14288,N_14330);
and U14749 (N_14749,N_14213,N_14106);
nor U14750 (N_14750,N_14329,N_14484);
nor U14751 (N_14751,N_14114,N_14033);
or U14752 (N_14752,N_14013,N_14163);
nor U14753 (N_14753,N_14274,N_14229);
xnor U14754 (N_14754,N_14459,N_14015);
xor U14755 (N_14755,N_14115,N_14260);
xnor U14756 (N_14756,N_14026,N_14217);
nand U14757 (N_14757,N_14274,N_14188);
nor U14758 (N_14758,N_14144,N_14003);
nand U14759 (N_14759,N_14174,N_14167);
or U14760 (N_14760,N_14476,N_14088);
and U14761 (N_14761,N_14373,N_14439);
nand U14762 (N_14762,N_14081,N_14250);
xor U14763 (N_14763,N_14273,N_14446);
nor U14764 (N_14764,N_14186,N_14095);
nor U14765 (N_14765,N_14454,N_14415);
and U14766 (N_14766,N_14014,N_14263);
nor U14767 (N_14767,N_14468,N_14015);
nand U14768 (N_14768,N_14352,N_14196);
or U14769 (N_14769,N_14421,N_14241);
nor U14770 (N_14770,N_14183,N_14361);
nor U14771 (N_14771,N_14340,N_14317);
and U14772 (N_14772,N_14162,N_14414);
nand U14773 (N_14773,N_14131,N_14028);
xor U14774 (N_14774,N_14391,N_14180);
nor U14775 (N_14775,N_14095,N_14213);
or U14776 (N_14776,N_14459,N_14080);
xor U14777 (N_14777,N_14008,N_14013);
and U14778 (N_14778,N_14249,N_14014);
nand U14779 (N_14779,N_14024,N_14017);
nand U14780 (N_14780,N_14146,N_14433);
or U14781 (N_14781,N_14268,N_14090);
nor U14782 (N_14782,N_14312,N_14019);
nand U14783 (N_14783,N_14204,N_14484);
xor U14784 (N_14784,N_14201,N_14477);
or U14785 (N_14785,N_14338,N_14219);
nand U14786 (N_14786,N_14063,N_14435);
or U14787 (N_14787,N_14002,N_14014);
and U14788 (N_14788,N_14356,N_14018);
nand U14789 (N_14789,N_14411,N_14382);
nor U14790 (N_14790,N_14438,N_14047);
xor U14791 (N_14791,N_14278,N_14153);
nor U14792 (N_14792,N_14009,N_14215);
nor U14793 (N_14793,N_14153,N_14331);
nand U14794 (N_14794,N_14316,N_14315);
or U14795 (N_14795,N_14430,N_14336);
and U14796 (N_14796,N_14420,N_14312);
nor U14797 (N_14797,N_14101,N_14031);
xor U14798 (N_14798,N_14059,N_14457);
and U14799 (N_14799,N_14412,N_14069);
xor U14800 (N_14800,N_14023,N_14240);
nor U14801 (N_14801,N_14430,N_14221);
and U14802 (N_14802,N_14105,N_14138);
and U14803 (N_14803,N_14119,N_14259);
nand U14804 (N_14804,N_14346,N_14265);
nand U14805 (N_14805,N_14071,N_14346);
or U14806 (N_14806,N_14425,N_14457);
or U14807 (N_14807,N_14286,N_14459);
and U14808 (N_14808,N_14318,N_14219);
nand U14809 (N_14809,N_14297,N_14390);
nand U14810 (N_14810,N_14196,N_14124);
or U14811 (N_14811,N_14138,N_14329);
nand U14812 (N_14812,N_14094,N_14434);
xnor U14813 (N_14813,N_14097,N_14042);
nor U14814 (N_14814,N_14367,N_14160);
nor U14815 (N_14815,N_14010,N_14286);
nand U14816 (N_14816,N_14196,N_14191);
or U14817 (N_14817,N_14461,N_14259);
and U14818 (N_14818,N_14220,N_14188);
and U14819 (N_14819,N_14429,N_14361);
nor U14820 (N_14820,N_14217,N_14494);
or U14821 (N_14821,N_14266,N_14265);
nand U14822 (N_14822,N_14327,N_14276);
nand U14823 (N_14823,N_14440,N_14170);
or U14824 (N_14824,N_14009,N_14455);
nand U14825 (N_14825,N_14362,N_14246);
nand U14826 (N_14826,N_14096,N_14374);
xor U14827 (N_14827,N_14326,N_14387);
and U14828 (N_14828,N_14198,N_14370);
nand U14829 (N_14829,N_14199,N_14265);
and U14830 (N_14830,N_14044,N_14457);
or U14831 (N_14831,N_14214,N_14372);
or U14832 (N_14832,N_14064,N_14347);
nand U14833 (N_14833,N_14277,N_14463);
nand U14834 (N_14834,N_14370,N_14088);
and U14835 (N_14835,N_14085,N_14206);
and U14836 (N_14836,N_14022,N_14141);
and U14837 (N_14837,N_14205,N_14392);
nor U14838 (N_14838,N_14405,N_14179);
and U14839 (N_14839,N_14365,N_14026);
xor U14840 (N_14840,N_14237,N_14391);
nand U14841 (N_14841,N_14028,N_14069);
or U14842 (N_14842,N_14056,N_14182);
and U14843 (N_14843,N_14174,N_14114);
nor U14844 (N_14844,N_14322,N_14028);
nand U14845 (N_14845,N_14368,N_14477);
and U14846 (N_14846,N_14132,N_14393);
xnor U14847 (N_14847,N_14247,N_14302);
nand U14848 (N_14848,N_14409,N_14325);
xnor U14849 (N_14849,N_14488,N_14262);
nor U14850 (N_14850,N_14341,N_14288);
xor U14851 (N_14851,N_14380,N_14168);
or U14852 (N_14852,N_14201,N_14494);
xor U14853 (N_14853,N_14027,N_14084);
and U14854 (N_14854,N_14249,N_14162);
nand U14855 (N_14855,N_14111,N_14400);
or U14856 (N_14856,N_14203,N_14381);
or U14857 (N_14857,N_14057,N_14288);
xnor U14858 (N_14858,N_14353,N_14097);
or U14859 (N_14859,N_14179,N_14343);
xnor U14860 (N_14860,N_14302,N_14403);
and U14861 (N_14861,N_14489,N_14216);
nor U14862 (N_14862,N_14113,N_14267);
or U14863 (N_14863,N_14475,N_14381);
nand U14864 (N_14864,N_14145,N_14413);
nand U14865 (N_14865,N_14094,N_14061);
and U14866 (N_14866,N_14174,N_14395);
nor U14867 (N_14867,N_14234,N_14491);
xnor U14868 (N_14868,N_14115,N_14112);
nor U14869 (N_14869,N_14254,N_14029);
nand U14870 (N_14870,N_14411,N_14468);
xnor U14871 (N_14871,N_14202,N_14457);
nor U14872 (N_14872,N_14423,N_14312);
or U14873 (N_14873,N_14014,N_14115);
nand U14874 (N_14874,N_14195,N_14443);
nor U14875 (N_14875,N_14386,N_14281);
xor U14876 (N_14876,N_14080,N_14125);
and U14877 (N_14877,N_14322,N_14112);
nor U14878 (N_14878,N_14162,N_14372);
or U14879 (N_14879,N_14136,N_14189);
or U14880 (N_14880,N_14274,N_14363);
nor U14881 (N_14881,N_14261,N_14007);
nor U14882 (N_14882,N_14376,N_14371);
or U14883 (N_14883,N_14324,N_14074);
nor U14884 (N_14884,N_14195,N_14364);
nor U14885 (N_14885,N_14186,N_14213);
or U14886 (N_14886,N_14268,N_14431);
or U14887 (N_14887,N_14124,N_14136);
or U14888 (N_14888,N_14417,N_14383);
nand U14889 (N_14889,N_14402,N_14032);
and U14890 (N_14890,N_14474,N_14480);
nand U14891 (N_14891,N_14243,N_14114);
xnor U14892 (N_14892,N_14104,N_14150);
and U14893 (N_14893,N_14030,N_14163);
nor U14894 (N_14894,N_14036,N_14260);
nor U14895 (N_14895,N_14401,N_14366);
nor U14896 (N_14896,N_14113,N_14380);
and U14897 (N_14897,N_14238,N_14165);
nand U14898 (N_14898,N_14193,N_14202);
or U14899 (N_14899,N_14099,N_14083);
or U14900 (N_14900,N_14077,N_14042);
nand U14901 (N_14901,N_14335,N_14090);
xor U14902 (N_14902,N_14343,N_14401);
and U14903 (N_14903,N_14037,N_14491);
xor U14904 (N_14904,N_14256,N_14027);
and U14905 (N_14905,N_14126,N_14008);
and U14906 (N_14906,N_14411,N_14455);
xor U14907 (N_14907,N_14183,N_14303);
and U14908 (N_14908,N_14189,N_14183);
and U14909 (N_14909,N_14169,N_14449);
or U14910 (N_14910,N_14205,N_14348);
nand U14911 (N_14911,N_14179,N_14021);
and U14912 (N_14912,N_14397,N_14019);
nand U14913 (N_14913,N_14154,N_14408);
nand U14914 (N_14914,N_14101,N_14356);
and U14915 (N_14915,N_14492,N_14196);
nand U14916 (N_14916,N_14286,N_14259);
nor U14917 (N_14917,N_14309,N_14071);
or U14918 (N_14918,N_14472,N_14311);
nor U14919 (N_14919,N_14018,N_14041);
and U14920 (N_14920,N_14153,N_14299);
or U14921 (N_14921,N_14240,N_14150);
nand U14922 (N_14922,N_14225,N_14437);
and U14923 (N_14923,N_14066,N_14051);
nand U14924 (N_14924,N_14091,N_14476);
or U14925 (N_14925,N_14057,N_14253);
xor U14926 (N_14926,N_14396,N_14152);
nand U14927 (N_14927,N_14089,N_14184);
nor U14928 (N_14928,N_14063,N_14203);
and U14929 (N_14929,N_14422,N_14328);
xor U14930 (N_14930,N_14211,N_14414);
xnor U14931 (N_14931,N_14223,N_14076);
or U14932 (N_14932,N_14388,N_14414);
xor U14933 (N_14933,N_14163,N_14237);
and U14934 (N_14934,N_14320,N_14198);
nand U14935 (N_14935,N_14123,N_14127);
xor U14936 (N_14936,N_14304,N_14012);
or U14937 (N_14937,N_14489,N_14040);
nand U14938 (N_14938,N_14144,N_14494);
or U14939 (N_14939,N_14396,N_14446);
nor U14940 (N_14940,N_14119,N_14206);
nor U14941 (N_14941,N_14231,N_14248);
or U14942 (N_14942,N_14058,N_14119);
xnor U14943 (N_14943,N_14319,N_14096);
and U14944 (N_14944,N_14157,N_14201);
xor U14945 (N_14945,N_14144,N_14178);
or U14946 (N_14946,N_14150,N_14303);
nor U14947 (N_14947,N_14227,N_14114);
nand U14948 (N_14948,N_14337,N_14477);
nor U14949 (N_14949,N_14147,N_14098);
nand U14950 (N_14950,N_14192,N_14423);
nor U14951 (N_14951,N_14245,N_14023);
nand U14952 (N_14952,N_14403,N_14153);
and U14953 (N_14953,N_14064,N_14354);
and U14954 (N_14954,N_14187,N_14086);
or U14955 (N_14955,N_14320,N_14027);
and U14956 (N_14956,N_14346,N_14052);
nand U14957 (N_14957,N_14232,N_14421);
and U14958 (N_14958,N_14067,N_14335);
nor U14959 (N_14959,N_14304,N_14477);
nor U14960 (N_14960,N_14355,N_14257);
or U14961 (N_14961,N_14012,N_14055);
nand U14962 (N_14962,N_14162,N_14438);
nand U14963 (N_14963,N_14048,N_14390);
or U14964 (N_14964,N_14229,N_14115);
or U14965 (N_14965,N_14421,N_14235);
nand U14966 (N_14966,N_14141,N_14472);
and U14967 (N_14967,N_14448,N_14368);
or U14968 (N_14968,N_14205,N_14437);
nor U14969 (N_14969,N_14230,N_14007);
or U14970 (N_14970,N_14208,N_14173);
or U14971 (N_14971,N_14098,N_14078);
nand U14972 (N_14972,N_14073,N_14062);
or U14973 (N_14973,N_14069,N_14217);
and U14974 (N_14974,N_14214,N_14377);
nor U14975 (N_14975,N_14382,N_14226);
xor U14976 (N_14976,N_14185,N_14320);
and U14977 (N_14977,N_14038,N_14063);
nor U14978 (N_14978,N_14271,N_14376);
or U14979 (N_14979,N_14208,N_14308);
nor U14980 (N_14980,N_14217,N_14137);
nand U14981 (N_14981,N_14407,N_14175);
nor U14982 (N_14982,N_14156,N_14276);
nor U14983 (N_14983,N_14156,N_14151);
xnor U14984 (N_14984,N_14244,N_14469);
or U14985 (N_14985,N_14320,N_14187);
xnor U14986 (N_14986,N_14489,N_14337);
and U14987 (N_14987,N_14188,N_14345);
nand U14988 (N_14988,N_14271,N_14043);
and U14989 (N_14989,N_14139,N_14217);
or U14990 (N_14990,N_14482,N_14299);
or U14991 (N_14991,N_14075,N_14240);
nand U14992 (N_14992,N_14205,N_14042);
xor U14993 (N_14993,N_14138,N_14332);
or U14994 (N_14994,N_14277,N_14081);
nand U14995 (N_14995,N_14218,N_14347);
nor U14996 (N_14996,N_14001,N_14456);
nand U14997 (N_14997,N_14025,N_14001);
nand U14998 (N_14998,N_14008,N_14341);
nor U14999 (N_14999,N_14086,N_14318);
or U15000 (N_15000,N_14721,N_14960);
xnor U15001 (N_15001,N_14550,N_14570);
nand U15002 (N_15002,N_14852,N_14706);
xnor U15003 (N_15003,N_14518,N_14560);
nand U15004 (N_15004,N_14583,N_14548);
nor U15005 (N_15005,N_14957,N_14800);
nand U15006 (N_15006,N_14596,N_14579);
and U15007 (N_15007,N_14505,N_14746);
and U15008 (N_15008,N_14634,N_14551);
or U15009 (N_15009,N_14868,N_14576);
or U15010 (N_15010,N_14833,N_14653);
nor U15011 (N_15011,N_14669,N_14780);
xor U15012 (N_15012,N_14502,N_14811);
nand U15013 (N_15013,N_14668,N_14781);
xnor U15014 (N_15014,N_14948,N_14585);
or U15015 (N_15015,N_14783,N_14972);
nand U15016 (N_15016,N_14798,N_14999);
nor U15017 (N_15017,N_14763,N_14924);
and U15018 (N_15018,N_14542,N_14575);
or U15019 (N_15019,N_14638,N_14609);
nand U15020 (N_15020,N_14792,N_14526);
xnor U15021 (N_15021,N_14709,N_14739);
or U15022 (N_15022,N_14680,N_14693);
nand U15023 (N_15023,N_14544,N_14582);
nand U15024 (N_15024,N_14731,N_14617);
nor U15025 (N_15025,N_14807,N_14651);
xnor U15026 (N_15026,N_14779,N_14742);
xnor U15027 (N_15027,N_14590,N_14765);
nand U15028 (N_15028,N_14600,N_14987);
nand U15029 (N_15029,N_14821,N_14831);
and U15030 (N_15030,N_14993,N_14573);
or U15031 (N_15031,N_14819,N_14572);
nand U15032 (N_15032,N_14973,N_14664);
nor U15033 (N_15033,N_14768,N_14869);
nor U15034 (N_15034,N_14732,N_14877);
and U15035 (N_15035,N_14894,N_14873);
or U15036 (N_15036,N_14778,N_14881);
and U15037 (N_15037,N_14674,N_14647);
nor U15038 (N_15038,N_14809,N_14918);
and U15039 (N_15039,N_14908,N_14753);
or U15040 (N_15040,N_14541,N_14661);
or U15041 (N_15041,N_14789,N_14546);
xnor U15042 (N_15042,N_14509,N_14929);
nor U15043 (N_15043,N_14621,N_14545);
nor U15044 (N_15044,N_14979,N_14872);
xnor U15045 (N_15045,N_14747,N_14851);
or U15046 (N_15046,N_14650,N_14959);
and U15047 (N_15047,N_14662,N_14602);
or U15048 (N_15048,N_14786,N_14828);
nand U15049 (N_15049,N_14648,N_14614);
nor U15050 (N_15050,N_14755,N_14915);
nor U15051 (N_15051,N_14538,N_14752);
or U15052 (N_15052,N_14720,N_14848);
nor U15053 (N_15053,N_14727,N_14899);
xnor U15054 (N_15054,N_14967,N_14659);
nor U15055 (N_15055,N_14622,N_14595);
nand U15056 (N_15056,N_14953,N_14598);
and U15057 (N_15057,N_14611,N_14860);
nand U15058 (N_15058,N_14776,N_14904);
or U15059 (N_15059,N_14888,N_14871);
and U15060 (N_15060,N_14687,N_14939);
nand U15061 (N_15061,N_14802,N_14795);
nand U15062 (N_15062,N_14907,N_14846);
and U15063 (N_15063,N_14823,N_14503);
and U15064 (N_15064,N_14782,N_14784);
nor U15065 (N_15065,N_14707,N_14898);
nor U15066 (N_15066,N_14847,N_14603);
or U15067 (N_15067,N_14667,N_14718);
xnor U15068 (N_15068,N_14855,N_14761);
nand U15069 (N_15069,N_14961,N_14970);
nand U15070 (N_15070,N_14808,N_14760);
nor U15071 (N_15071,N_14903,N_14977);
xor U15072 (N_15072,N_14555,N_14750);
nor U15073 (N_15073,N_14552,N_14744);
nand U15074 (N_15074,N_14919,N_14946);
or U15075 (N_15075,N_14685,N_14825);
nor U15076 (N_15076,N_14604,N_14988);
nor U15077 (N_15077,N_14827,N_14559);
xor U15078 (N_15078,N_14805,N_14818);
xor U15079 (N_15079,N_14949,N_14803);
nand U15080 (N_15080,N_14564,N_14978);
nand U15081 (N_15081,N_14882,N_14917);
xnor U15082 (N_15082,N_14681,N_14719);
nor U15083 (N_15083,N_14994,N_14867);
or U15084 (N_15084,N_14769,N_14516);
nor U15085 (N_15085,N_14968,N_14722);
nor U15086 (N_15086,N_14735,N_14991);
or U15087 (N_15087,N_14649,N_14701);
and U15088 (N_15088,N_14530,N_14906);
or U15089 (N_15089,N_14601,N_14658);
and U15090 (N_15090,N_14854,N_14514);
and U15091 (N_15091,N_14500,N_14626);
or U15092 (N_15092,N_14840,N_14524);
or U15093 (N_15093,N_14952,N_14986);
or U15094 (N_15094,N_14513,N_14878);
nor U15095 (N_15095,N_14901,N_14817);
xor U15096 (N_15096,N_14686,N_14512);
nand U15097 (N_15097,N_14976,N_14921);
nand U15098 (N_15098,N_14895,N_14943);
and U15099 (N_15099,N_14858,N_14588);
xnor U15100 (N_15100,N_14511,N_14824);
and U15101 (N_15101,N_14565,N_14689);
and U15102 (N_15102,N_14510,N_14702);
nand U15103 (N_15103,N_14625,N_14504);
and U15104 (N_15104,N_14951,N_14829);
or U15105 (N_15105,N_14591,N_14711);
xnor U15106 (N_15106,N_14998,N_14554);
nand U15107 (N_15107,N_14536,N_14635);
xnor U15108 (N_15108,N_14844,N_14995);
or U15109 (N_15109,N_14937,N_14799);
and U15110 (N_15110,N_14941,N_14982);
and U15111 (N_15111,N_14640,N_14637);
xnor U15112 (N_15112,N_14631,N_14713);
nand U15113 (N_15113,N_14633,N_14944);
nand U15114 (N_15114,N_14945,N_14629);
and U15115 (N_15115,N_14695,N_14856);
and U15116 (N_15116,N_14594,N_14812);
and U15117 (N_15117,N_14521,N_14885);
nand U15118 (N_15118,N_14879,N_14745);
xnor U15119 (N_15119,N_14599,N_14643);
nand U15120 (N_15120,N_14566,N_14553);
and U15121 (N_15121,N_14734,N_14756);
nor U15122 (N_15122,N_14954,N_14835);
or U15123 (N_15123,N_14642,N_14962);
xnor U15124 (N_15124,N_14677,N_14905);
nor U15125 (N_15125,N_14955,N_14738);
and U15126 (N_15126,N_14561,N_14574);
nand U15127 (N_15127,N_14699,N_14880);
or U15128 (N_15128,N_14612,N_14933);
xor U15129 (N_15129,N_14627,N_14708);
nand U15130 (N_15130,N_14684,N_14810);
nor U15131 (N_15131,N_14717,N_14532);
xnor U15132 (N_15132,N_14777,N_14927);
and U15133 (N_15133,N_14790,N_14992);
nor U15134 (N_15134,N_14534,N_14826);
xor U15135 (N_15135,N_14989,N_14696);
or U15136 (N_15136,N_14675,N_14522);
nand U15137 (N_15137,N_14710,N_14916);
nand U15138 (N_15138,N_14730,N_14733);
nand U15139 (N_15139,N_14892,N_14922);
xnor U15140 (N_15140,N_14607,N_14682);
and U15141 (N_15141,N_14911,N_14839);
or U15142 (N_15142,N_14531,N_14690);
xnor U15143 (N_15143,N_14624,N_14587);
xor U15144 (N_15144,N_14563,N_14920);
nor U15145 (N_15145,N_14679,N_14501);
or U15146 (N_15146,N_14963,N_14766);
or U15147 (N_15147,N_14751,N_14641);
and U15148 (N_15148,N_14997,N_14608);
xnor U15149 (N_15149,N_14673,N_14985);
nand U15150 (N_15150,N_14549,N_14618);
and U15151 (N_15151,N_14645,N_14620);
or U15152 (N_15152,N_14771,N_14813);
nand U15153 (N_15153,N_14740,N_14723);
and U15154 (N_15154,N_14644,N_14515);
xor U15155 (N_15155,N_14547,N_14703);
or U15156 (N_15156,N_14764,N_14866);
xor U15157 (N_15157,N_14528,N_14666);
and U15158 (N_15158,N_14925,N_14537);
xnor U15159 (N_15159,N_14688,N_14646);
nor U15160 (N_15160,N_14796,N_14947);
nor U15161 (N_15161,N_14716,N_14527);
or U15162 (N_15162,N_14935,N_14672);
and U15163 (N_15163,N_14887,N_14671);
nor U15164 (N_15164,N_14592,N_14874);
and U15165 (N_15165,N_14950,N_14584);
and U15166 (N_15166,N_14774,N_14700);
or U15167 (N_15167,N_14902,N_14996);
xnor U15168 (N_15168,N_14577,N_14736);
or U15169 (N_15169,N_14568,N_14931);
and U15170 (N_15170,N_14581,N_14990);
and U15171 (N_15171,N_14791,N_14865);
nor U15172 (N_15172,N_14942,N_14801);
and U15173 (N_15173,N_14543,N_14593);
or U15174 (N_15174,N_14533,N_14540);
nor U15175 (N_15175,N_14926,N_14788);
nor U15176 (N_15176,N_14928,N_14849);
nand U15177 (N_15177,N_14912,N_14793);
nor U15178 (N_15178,N_14726,N_14770);
and U15179 (N_15179,N_14729,N_14670);
xor U15180 (N_15180,N_14656,N_14748);
nand U15181 (N_15181,N_14893,N_14785);
or U15182 (N_15182,N_14619,N_14694);
and U15183 (N_15183,N_14632,N_14900);
xor U15184 (N_15184,N_14862,N_14558);
or U15185 (N_15185,N_14984,N_14569);
nor U15186 (N_15186,N_14520,N_14556);
or U15187 (N_15187,N_14562,N_14571);
or U15188 (N_15188,N_14966,N_14652);
nor U15189 (N_15189,N_14930,N_14938);
nand U15190 (N_15190,N_14897,N_14870);
and U15191 (N_15191,N_14857,N_14936);
nand U15192 (N_15192,N_14842,N_14876);
nand U15193 (N_15193,N_14875,N_14657);
and U15194 (N_15194,N_14630,N_14913);
nor U15195 (N_15195,N_14525,N_14815);
and U15196 (N_15196,N_14724,N_14610);
xor U15197 (N_15197,N_14891,N_14758);
nor U15198 (N_15198,N_14822,N_14836);
xnor U15199 (N_15199,N_14741,N_14691);
and U15200 (N_15200,N_14838,N_14692);
xnor U15201 (N_15201,N_14517,N_14728);
or U15202 (N_15202,N_14883,N_14884);
and U15203 (N_15203,N_14843,N_14889);
nand U15204 (N_15204,N_14557,N_14683);
nand U15205 (N_15205,N_14712,N_14830);
nor U15206 (N_15206,N_14636,N_14697);
and U15207 (N_15207,N_14806,N_14678);
nor U15208 (N_15208,N_14923,N_14820);
nand U15209 (N_15209,N_14980,N_14845);
nand U15210 (N_15210,N_14586,N_14714);
nor U15211 (N_15211,N_14605,N_14754);
xnor U15212 (N_15212,N_14804,N_14639);
xor U15213 (N_15213,N_14589,N_14956);
and U15214 (N_15214,N_14757,N_14567);
and U15215 (N_15215,N_14759,N_14519);
nand U15216 (N_15216,N_14864,N_14861);
or U15217 (N_15217,N_14837,N_14909);
nor U15218 (N_15218,N_14794,N_14863);
or U15219 (N_15219,N_14743,N_14762);
nand U15220 (N_15220,N_14506,N_14975);
xnor U15221 (N_15221,N_14775,N_14886);
nand U15222 (N_15222,N_14705,N_14663);
xor U15223 (N_15223,N_14654,N_14969);
and U15224 (N_15224,N_14853,N_14539);
nand U15225 (N_15225,N_14725,N_14676);
and U15226 (N_15226,N_14958,N_14932);
and U15227 (N_15227,N_14597,N_14981);
and U15228 (N_15228,N_14698,N_14890);
or U15229 (N_15229,N_14841,N_14628);
xor U15230 (N_15230,N_14616,N_14974);
nor U15231 (N_15231,N_14613,N_14787);
and U15232 (N_15232,N_14529,N_14715);
and U15233 (N_15233,N_14665,N_14834);
nor U15234 (N_15234,N_14816,N_14934);
nand U15235 (N_15235,N_14523,N_14896);
nand U15236 (N_15236,N_14983,N_14965);
xor U15237 (N_15237,N_14578,N_14910);
and U15238 (N_15238,N_14773,N_14749);
and U15239 (N_15239,N_14832,N_14772);
or U15240 (N_15240,N_14660,N_14606);
nand U15241 (N_15241,N_14850,N_14580);
or U15242 (N_15242,N_14971,N_14797);
nor U15243 (N_15243,N_14507,N_14814);
and U15244 (N_15244,N_14623,N_14508);
or U15245 (N_15245,N_14940,N_14615);
nor U15246 (N_15246,N_14767,N_14914);
or U15247 (N_15247,N_14704,N_14737);
or U15248 (N_15248,N_14535,N_14655);
xnor U15249 (N_15249,N_14964,N_14859);
and U15250 (N_15250,N_14864,N_14686);
xor U15251 (N_15251,N_14950,N_14502);
nand U15252 (N_15252,N_14588,N_14711);
or U15253 (N_15253,N_14616,N_14800);
nand U15254 (N_15254,N_14987,N_14957);
xor U15255 (N_15255,N_14759,N_14507);
xor U15256 (N_15256,N_14743,N_14865);
and U15257 (N_15257,N_14701,N_14694);
or U15258 (N_15258,N_14820,N_14722);
and U15259 (N_15259,N_14690,N_14839);
xnor U15260 (N_15260,N_14541,N_14516);
and U15261 (N_15261,N_14690,N_14863);
nor U15262 (N_15262,N_14815,N_14756);
nor U15263 (N_15263,N_14537,N_14913);
xnor U15264 (N_15264,N_14601,N_14645);
nand U15265 (N_15265,N_14720,N_14823);
or U15266 (N_15266,N_14983,N_14760);
xnor U15267 (N_15267,N_14702,N_14622);
xnor U15268 (N_15268,N_14829,N_14774);
xnor U15269 (N_15269,N_14749,N_14507);
xnor U15270 (N_15270,N_14862,N_14956);
and U15271 (N_15271,N_14516,N_14936);
or U15272 (N_15272,N_14842,N_14536);
nor U15273 (N_15273,N_14619,N_14671);
nor U15274 (N_15274,N_14783,N_14851);
xor U15275 (N_15275,N_14541,N_14872);
and U15276 (N_15276,N_14582,N_14811);
xor U15277 (N_15277,N_14691,N_14831);
xor U15278 (N_15278,N_14733,N_14679);
and U15279 (N_15279,N_14551,N_14900);
nand U15280 (N_15280,N_14998,N_14763);
nor U15281 (N_15281,N_14587,N_14633);
nand U15282 (N_15282,N_14765,N_14994);
and U15283 (N_15283,N_14921,N_14518);
nor U15284 (N_15284,N_14684,N_14733);
or U15285 (N_15285,N_14593,N_14873);
and U15286 (N_15286,N_14578,N_14883);
nor U15287 (N_15287,N_14915,N_14902);
nand U15288 (N_15288,N_14924,N_14956);
or U15289 (N_15289,N_14970,N_14511);
nor U15290 (N_15290,N_14506,N_14631);
nor U15291 (N_15291,N_14801,N_14603);
nand U15292 (N_15292,N_14992,N_14947);
xnor U15293 (N_15293,N_14993,N_14524);
nor U15294 (N_15294,N_14596,N_14922);
or U15295 (N_15295,N_14869,N_14813);
nor U15296 (N_15296,N_14536,N_14762);
nor U15297 (N_15297,N_14648,N_14819);
nand U15298 (N_15298,N_14936,N_14978);
nor U15299 (N_15299,N_14658,N_14976);
and U15300 (N_15300,N_14770,N_14939);
xor U15301 (N_15301,N_14743,N_14854);
and U15302 (N_15302,N_14728,N_14742);
xnor U15303 (N_15303,N_14568,N_14538);
and U15304 (N_15304,N_14720,N_14988);
nor U15305 (N_15305,N_14531,N_14844);
or U15306 (N_15306,N_14987,N_14916);
nand U15307 (N_15307,N_14807,N_14776);
nand U15308 (N_15308,N_14501,N_14896);
xnor U15309 (N_15309,N_14844,N_14611);
or U15310 (N_15310,N_14744,N_14743);
xor U15311 (N_15311,N_14803,N_14931);
nand U15312 (N_15312,N_14578,N_14676);
and U15313 (N_15313,N_14805,N_14904);
nand U15314 (N_15314,N_14986,N_14800);
nor U15315 (N_15315,N_14753,N_14981);
xnor U15316 (N_15316,N_14910,N_14693);
and U15317 (N_15317,N_14572,N_14586);
xor U15318 (N_15318,N_14953,N_14766);
xnor U15319 (N_15319,N_14544,N_14775);
nand U15320 (N_15320,N_14836,N_14886);
nor U15321 (N_15321,N_14876,N_14780);
or U15322 (N_15322,N_14692,N_14804);
xor U15323 (N_15323,N_14891,N_14664);
nand U15324 (N_15324,N_14772,N_14812);
xnor U15325 (N_15325,N_14546,N_14669);
nor U15326 (N_15326,N_14548,N_14558);
and U15327 (N_15327,N_14682,N_14780);
xnor U15328 (N_15328,N_14573,N_14677);
or U15329 (N_15329,N_14585,N_14739);
and U15330 (N_15330,N_14852,N_14558);
and U15331 (N_15331,N_14793,N_14938);
or U15332 (N_15332,N_14916,N_14919);
nor U15333 (N_15333,N_14831,N_14982);
nand U15334 (N_15334,N_14545,N_14503);
and U15335 (N_15335,N_14812,N_14829);
xnor U15336 (N_15336,N_14770,N_14677);
and U15337 (N_15337,N_14848,N_14885);
nand U15338 (N_15338,N_14648,N_14659);
xnor U15339 (N_15339,N_14594,N_14618);
and U15340 (N_15340,N_14776,N_14520);
nor U15341 (N_15341,N_14710,N_14955);
nor U15342 (N_15342,N_14948,N_14619);
nand U15343 (N_15343,N_14825,N_14928);
nand U15344 (N_15344,N_14958,N_14709);
xor U15345 (N_15345,N_14986,N_14905);
nand U15346 (N_15346,N_14978,N_14513);
nor U15347 (N_15347,N_14629,N_14939);
or U15348 (N_15348,N_14972,N_14579);
and U15349 (N_15349,N_14687,N_14638);
nand U15350 (N_15350,N_14805,N_14733);
nor U15351 (N_15351,N_14973,N_14706);
xnor U15352 (N_15352,N_14758,N_14807);
nand U15353 (N_15353,N_14716,N_14635);
and U15354 (N_15354,N_14956,N_14867);
xor U15355 (N_15355,N_14959,N_14652);
xor U15356 (N_15356,N_14785,N_14964);
or U15357 (N_15357,N_14612,N_14558);
or U15358 (N_15358,N_14598,N_14720);
and U15359 (N_15359,N_14553,N_14554);
and U15360 (N_15360,N_14979,N_14985);
or U15361 (N_15361,N_14826,N_14647);
nor U15362 (N_15362,N_14733,N_14747);
nand U15363 (N_15363,N_14959,N_14949);
nor U15364 (N_15364,N_14927,N_14901);
nand U15365 (N_15365,N_14502,N_14618);
xnor U15366 (N_15366,N_14991,N_14602);
and U15367 (N_15367,N_14990,N_14781);
nor U15368 (N_15368,N_14967,N_14565);
and U15369 (N_15369,N_14695,N_14594);
nor U15370 (N_15370,N_14911,N_14540);
and U15371 (N_15371,N_14580,N_14615);
nor U15372 (N_15372,N_14855,N_14671);
xor U15373 (N_15373,N_14899,N_14969);
and U15374 (N_15374,N_14927,N_14735);
xor U15375 (N_15375,N_14805,N_14699);
xnor U15376 (N_15376,N_14550,N_14718);
and U15377 (N_15377,N_14793,N_14629);
or U15378 (N_15378,N_14595,N_14650);
nand U15379 (N_15379,N_14922,N_14863);
or U15380 (N_15380,N_14515,N_14661);
and U15381 (N_15381,N_14550,N_14510);
xnor U15382 (N_15382,N_14767,N_14697);
nor U15383 (N_15383,N_14978,N_14824);
nor U15384 (N_15384,N_14815,N_14528);
nor U15385 (N_15385,N_14544,N_14705);
nor U15386 (N_15386,N_14538,N_14550);
nand U15387 (N_15387,N_14751,N_14960);
and U15388 (N_15388,N_14894,N_14768);
xnor U15389 (N_15389,N_14862,N_14626);
xnor U15390 (N_15390,N_14503,N_14938);
nand U15391 (N_15391,N_14620,N_14977);
or U15392 (N_15392,N_14993,N_14545);
xnor U15393 (N_15393,N_14774,N_14594);
xor U15394 (N_15394,N_14933,N_14605);
nand U15395 (N_15395,N_14644,N_14807);
nor U15396 (N_15396,N_14542,N_14756);
nor U15397 (N_15397,N_14749,N_14525);
or U15398 (N_15398,N_14730,N_14868);
nor U15399 (N_15399,N_14728,N_14702);
and U15400 (N_15400,N_14872,N_14741);
and U15401 (N_15401,N_14831,N_14580);
and U15402 (N_15402,N_14693,N_14639);
nor U15403 (N_15403,N_14958,N_14945);
nand U15404 (N_15404,N_14970,N_14505);
or U15405 (N_15405,N_14815,N_14536);
or U15406 (N_15406,N_14715,N_14860);
nor U15407 (N_15407,N_14767,N_14671);
nor U15408 (N_15408,N_14590,N_14610);
nand U15409 (N_15409,N_14517,N_14653);
nand U15410 (N_15410,N_14632,N_14941);
xnor U15411 (N_15411,N_14508,N_14855);
xnor U15412 (N_15412,N_14966,N_14687);
xnor U15413 (N_15413,N_14554,N_14875);
and U15414 (N_15414,N_14567,N_14849);
nor U15415 (N_15415,N_14585,N_14579);
or U15416 (N_15416,N_14674,N_14984);
xor U15417 (N_15417,N_14509,N_14672);
or U15418 (N_15418,N_14799,N_14569);
xnor U15419 (N_15419,N_14848,N_14762);
or U15420 (N_15420,N_14883,N_14519);
nand U15421 (N_15421,N_14564,N_14988);
or U15422 (N_15422,N_14638,N_14680);
and U15423 (N_15423,N_14781,N_14618);
or U15424 (N_15424,N_14992,N_14915);
nor U15425 (N_15425,N_14782,N_14627);
xor U15426 (N_15426,N_14816,N_14600);
nor U15427 (N_15427,N_14870,N_14709);
nor U15428 (N_15428,N_14670,N_14907);
and U15429 (N_15429,N_14968,N_14813);
nand U15430 (N_15430,N_14539,N_14861);
nor U15431 (N_15431,N_14732,N_14520);
and U15432 (N_15432,N_14701,N_14711);
nand U15433 (N_15433,N_14791,N_14930);
xor U15434 (N_15434,N_14730,N_14572);
nand U15435 (N_15435,N_14886,N_14724);
nand U15436 (N_15436,N_14896,N_14807);
nand U15437 (N_15437,N_14708,N_14900);
and U15438 (N_15438,N_14504,N_14942);
or U15439 (N_15439,N_14747,N_14986);
or U15440 (N_15440,N_14940,N_14617);
and U15441 (N_15441,N_14861,N_14820);
xor U15442 (N_15442,N_14608,N_14875);
xnor U15443 (N_15443,N_14720,N_14760);
nor U15444 (N_15444,N_14724,N_14987);
or U15445 (N_15445,N_14538,N_14784);
nor U15446 (N_15446,N_14699,N_14545);
nand U15447 (N_15447,N_14567,N_14766);
or U15448 (N_15448,N_14597,N_14890);
xnor U15449 (N_15449,N_14721,N_14644);
and U15450 (N_15450,N_14896,N_14892);
and U15451 (N_15451,N_14993,N_14628);
nand U15452 (N_15452,N_14688,N_14849);
or U15453 (N_15453,N_14870,N_14872);
nand U15454 (N_15454,N_14793,N_14671);
xor U15455 (N_15455,N_14700,N_14595);
nor U15456 (N_15456,N_14615,N_14884);
nand U15457 (N_15457,N_14654,N_14674);
xnor U15458 (N_15458,N_14928,N_14764);
and U15459 (N_15459,N_14564,N_14762);
and U15460 (N_15460,N_14955,N_14938);
xor U15461 (N_15461,N_14773,N_14778);
nand U15462 (N_15462,N_14741,N_14547);
nor U15463 (N_15463,N_14778,N_14559);
or U15464 (N_15464,N_14549,N_14751);
xor U15465 (N_15465,N_14642,N_14946);
nand U15466 (N_15466,N_14973,N_14682);
or U15467 (N_15467,N_14673,N_14886);
or U15468 (N_15468,N_14695,N_14971);
or U15469 (N_15469,N_14667,N_14835);
or U15470 (N_15470,N_14551,N_14554);
nand U15471 (N_15471,N_14905,N_14857);
xor U15472 (N_15472,N_14878,N_14996);
nand U15473 (N_15473,N_14655,N_14732);
xor U15474 (N_15474,N_14943,N_14530);
xor U15475 (N_15475,N_14886,N_14756);
and U15476 (N_15476,N_14735,N_14969);
and U15477 (N_15477,N_14722,N_14753);
or U15478 (N_15478,N_14963,N_14967);
or U15479 (N_15479,N_14538,N_14882);
or U15480 (N_15480,N_14761,N_14947);
or U15481 (N_15481,N_14966,N_14894);
nand U15482 (N_15482,N_14658,N_14802);
and U15483 (N_15483,N_14679,N_14942);
and U15484 (N_15484,N_14724,N_14698);
nor U15485 (N_15485,N_14826,N_14723);
nor U15486 (N_15486,N_14640,N_14737);
and U15487 (N_15487,N_14708,N_14871);
xor U15488 (N_15488,N_14670,N_14514);
nand U15489 (N_15489,N_14532,N_14698);
nor U15490 (N_15490,N_14965,N_14997);
nand U15491 (N_15491,N_14694,N_14888);
nand U15492 (N_15492,N_14525,N_14542);
nor U15493 (N_15493,N_14855,N_14799);
xor U15494 (N_15494,N_14932,N_14857);
nor U15495 (N_15495,N_14585,N_14781);
and U15496 (N_15496,N_14970,N_14950);
nor U15497 (N_15497,N_14852,N_14506);
nor U15498 (N_15498,N_14992,N_14537);
xnor U15499 (N_15499,N_14787,N_14647);
xor U15500 (N_15500,N_15226,N_15340);
xor U15501 (N_15501,N_15474,N_15475);
xor U15502 (N_15502,N_15489,N_15058);
nor U15503 (N_15503,N_15210,N_15373);
or U15504 (N_15504,N_15258,N_15337);
or U15505 (N_15505,N_15155,N_15317);
nand U15506 (N_15506,N_15031,N_15493);
xor U15507 (N_15507,N_15134,N_15019);
nand U15508 (N_15508,N_15293,N_15311);
or U15509 (N_15509,N_15144,N_15096);
xor U15510 (N_15510,N_15353,N_15471);
nor U15511 (N_15511,N_15344,N_15141);
nand U15512 (N_15512,N_15001,N_15336);
and U15513 (N_15513,N_15437,N_15047);
xnor U15514 (N_15514,N_15248,N_15117);
xnor U15515 (N_15515,N_15407,N_15268);
xnor U15516 (N_15516,N_15312,N_15222);
and U15517 (N_15517,N_15168,N_15093);
xor U15518 (N_15518,N_15254,N_15402);
nor U15519 (N_15519,N_15394,N_15456);
xnor U15520 (N_15520,N_15228,N_15316);
or U15521 (N_15521,N_15035,N_15390);
and U15522 (N_15522,N_15386,N_15213);
nand U15523 (N_15523,N_15364,N_15494);
nand U15524 (N_15524,N_15188,N_15321);
and U15525 (N_15525,N_15203,N_15218);
and U15526 (N_15526,N_15010,N_15120);
and U15527 (N_15527,N_15291,N_15007);
and U15528 (N_15528,N_15448,N_15063);
or U15529 (N_15529,N_15166,N_15370);
nor U15530 (N_15530,N_15159,N_15197);
nor U15531 (N_15531,N_15043,N_15114);
nand U15532 (N_15532,N_15314,N_15215);
nor U15533 (N_15533,N_15467,N_15261);
nor U15534 (N_15534,N_15173,N_15127);
or U15535 (N_15535,N_15032,N_15412);
xor U15536 (N_15536,N_15363,N_15046);
xor U15537 (N_15537,N_15492,N_15347);
nand U15538 (N_15538,N_15068,N_15212);
xor U15539 (N_15539,N_15450,N_15267);
or U15540 (N_15540,N_15375,N_15169);
nor U15541 (N_15541,N_15334,N_15078);
nor U15542 (N_15542,N_15053,N_15231);
and U15543 (N_15543,N_15171,N_15115);
or U15544 (N_15544,N_15004,N_15149);
nand U15545 (N_15545,N_15132,N_15080);
nor U15546 (N_15546,N_15275,N_15229);
nor U15547 (N_15547,N_15138,N_15069);
and U15548 (N_15548,N_15440,N_15436);
and U15549 (N_15549,N_15287,N_15331);
and U15550 (N_15550,N_15408,N_15161);
nand U15551 (N_15551,N_15464,N_15300);
xor U15552 (N_15552,N_15000,N_15220);
nor U15553 (N_15553,N_15247,N_15410);
nor U15554 (N_15554,N_15050,N_15062);
or U15555 (N_15555,N_15199,N_15483);
nor U15556 (N_15556,N_15129,N_15301);
or U15557 (N_15557,N_15462,N_15236);
nor U15558 (N_15558,N_15131,N_15012);
nor U15559 (N_15559,N_15143,N_15189);
nor U15560 (N_15560,N_15290,N_15385);
xnor U15561 (N_15561,N_15459,N_15147);
nor U15562 (N_15562,N_15082,N_15389);
nand U15563 (N_15563,N_15187,N_15259);
or U15564 (N_15564,N_15005,N_15310);
nor U15565 (N_15565,N_15029,N_15288);
nor U15566 (N_15566,N_15191,N_15454);
xnor U15567 (N_15567,N_15427,N_15413);
nand U15568 (N_15568,N_15235,N_15011);
xor U15569 (N_15569,N_15193,N_15030);
xnor U15570 (N_15570,N_15279,N_15152);
or U15571 (N_15571,N_15328,N_15185);
or U15572 (N_15572,N_15305,N_15024);
xnor U15573 (N_15573,N_15271,N_15482);
or U15574 (N_15574,N_15049,N_15183);
and U15575 (N_15575,N_15371,N_15455);
nand U15576 (N_15576,N_15322,N_15237);
nand U15577 (N_15577,N_15438,N_15230);
and U15578 (N_15578,N_15202,N_15051);
and U15579 (N_15579,N_15404,N_15447);
nand U15580 (N_15580,N_15146,N_15280);
xnor U15581 (N_15581,N_15048,N_15054);
xnor U15582 (N_15582,N_15318,N_15052);
xnor U15583 (N_15583,N_15377,N_15177);
or U15584 (N_15584,N_15255,N_15480);
nand U15585 (N_15585,N_15164,N_15002);
and U15586 (N_15586,N_15327,N_15232);
xnor U15587 (N_15587,N_15111,N_15071);
xnor U15588 (N_15588,N_15098,N_15260);
or U15589 (N_15589,N_15362,N_15233);
nor U15590 (N_15590,N_15463,N_15495);
nor U15591 (N_15591,N_15252,N_15251);
and U15592 (N_15592,N_15179,N_15013);
or U15593 (N_15593,N_15066,N_15196);
or U15594 (N_15594,N_15468,N_15444);
and U15595 (N_15595,N_15133,N_15335);
nor U15596 (N_15596,N_15104,N_15264);
nand U15597 (N_15597,N_15217,N_15360);
xor U15598 (N_15598,N_15195,N_15442);
and U15599 (N_15599,N_15206,N_15003);
or U15600 (N_15600,N_15384,N_15369);
and U15601 (N_15601,N_15378,N_15022);
nor U15602 (N_15602,N_15446,N_15021);
xor U15603 (N_15603,N_15405,N_15278);
or U15604 (N_15604,N_15490,N_15176);
xor U15605 (N_15605,N_15285,N_15097);
nor U15606 (N_15606,N_15130,N_15006);
nand U15607 (N_15607,N_15060,N_15214);
xor U15608 (N_15608,N_15008,N_15150);
or U15609 (N_15609,N_15128,N_15044);
and U15610 (N_15610,N_15042,N_15107);
nand U15611 (N_15611,N_15067,N_15272);
xnor U15612 (N_15612,N_15239,N_15014);
nand U15613 (N_15613,N_15295,N_15245);
nor U15614 (N_15614,N_15423,N_15397);
nand U15615 (N_15615,N_15142,N_15136);
nand U15616 (N_15616,N_15470,N_15421);
and U15617 (N_15617,N_15061,N_15339);
and U15618 (N_15618,N_15365,N_15250);
nor U15619 (N_15619,N_15399,N_15017);
nand U15620 (N_15620,N_15192,N_15351);
and U15621 (N_15621,N_15056,N_15366);
nand U15622 (N_15622,N_15204,N_15289);
xnor U15623 (N_15623,N_15180,N_15497);
nand U15624 (N_15624,N_15372,N_15422);
nand U15625 (N_15625,N_15498,N_15382);
nor U15626 (N_15626,N_15329,N_15038);
or U15627 (N_15627,N_15088,N_15085);
or U15628 (N_15628,N_15121,N_15383);
and U15629 (N_15629,N_15434,N_15084);
nand U15630 (N_15630,N_15297,N_15086);
xor U15631 (N_15631,N_15087,N_15379);
nand U15632 (N_15632,N_15367,N_15381);
and U15633 (N_15633,N_15211,N_15055);
and U15634 (N_15634,N_15485,N_15154);
nor U15635 (N_15635,N_15320,N_15449);
nand U15636 (N_15636,N_15477,N_15148);
nor U15637 (N_15637,N_15354,N_15424);
nand U15638 (N_15638,N_15345,N_15368);
nor U15639 (N_15639,N_15140,N_15425);
nor U15640 (N_15640,N_15387,N_15401);
nor U15641 (N_15641,N_15110,N_15292);
xor U15642 (N_15642,N_15246,N_15432);
nor U15643 (N_15643,N_15076,N_15341);
nand U15644 (N_15644,N_15296,N_15282);
and U15645 (N_15645,N_15355,N_15253);
nand U15646 (N_15646,N_15358,N_15453);
and U15647 (N_15647,N_15298,N_15243);
or U15648 (N_15648,N_15356,N_15175);
xor U15649 (N_15649,N_15263,N_15156);
or U15650 (N_15650,N_15332,N_15323);
or U15651 (N_15651,N_15077,N_15461);
xor U15652 (N_15652,N_15201,N_15108);
or U15653 (N_15653,N_15238,N_15009);
and U15654 (N_15654,N_15426,N_15380);
nand U15655 (N_15655,N_15023,N_15122);
nand U15656 (N_15656,N_15303,N_15361);
and U15657 (N_15657,N_15304,N_15075);
xor U15658 (N_15658,N_15348,N_15324);
nor U15659 (N_15659,N_15376,N_15325);
nor U15660 (N_15660,N_15416,N_15165);
xnor U15661 (N_15661,N_15198,N_15330);
nor U15662 (N_15662,N_15205,N_15276);
nor U15663 (N_15663,N_15395,N_15105);
or U15664 (N_15664,N_15270,N_15216);
nand U15665 (N_15665,N_15207,N_15181);
and U15666 (N_15666,N_15020,N_15074);
xnor U15667 (N_15667,N_15221,N_15209);
nor U15668 (N_15668,N_15452,N_15431);
and U15669 (N_15669,N_15342,N_15499);
nand U15670 (N_15670,N_15313,N_15308);
and U15671 (N_15671,N_15094,N_15445);
xnor U15672 (N_15672,N_15103,N_15458);
xnor U15673 (N_15673,N_15099,N_15040);
and U15674 (N_15674,N_15388,N_15419);
and U15675 (N_15675,N_15439,N_15451);
and U15676 (N_15676,N_15244,N_15262);
or U15677 (N_15677,N_15433,N_15083);
xnor U15678 (N_15678,N_15118,N_15123);
nor U15679 (N_15679,N_15025,N_15403);
and U15680 (N_15680,N_15306,N_15028);
xor U15681 (N_15681,N_15036,N_15145);
or U15682 (N_15682,N_15170,N_15409);
nor U15683 (N_15683,N_15319,N_15027);
nor U15684 (N_15684,N_15476,N_15277);
and U15685 (N_15685,N_15343,N_15472);
nor U15686 (N_15686,N_15172,N_15059);
and U15687 (N_15687,N_15157,N_15112);
or U15688 (N_15688,N_15153,N_15466);
nor U15689 (N_15689,N_15234,N_15286);
or U15690 (N_15690,N_15039,N_15266);
nor U15691 (N_15691,N_15240,N_15460);
xnor U15692 (N_15692,N_15469,N_15081);
and U15693 (N_15693,N_15139,N_15249);
xnor U15694 (N_15694,N_15057,N_15352);
nand U15695 (N_15695,N_15392,N_15346);
and U15696 (N_15696,N_15411,N_15224);
or U15697 (N_15697,N_15208,N_15333);
and U15698 (N_15698,N_15225,N_15417);
nand U15699 (N_15699,N_15307,N_15491);
nand U15700 (N_15700,N_15091,N_15223);
or U15701 (N_15701,N_15269,N_15374);
or U15702 (N_15702,N_15393,N_15178);
xor U15703 (N_15703,N_15092,N_15194);
nor U15704 (N_15704,N_15315,N_15284);
nor U15705 (N_15705,N_15190,N_15026);
xnor U15706 (N_15706,N_15163,N_15359);
xor U15707 (N_15707,N_15484,N_15227);
nand U15708 (N_15708,N_15037,N_15089);
and U15709 (N_15709,N_15326,N_15414);
xnor U15710 (N_15710,N_15070,N_15184);
nor U15711 (N_15711,N_15018,N_15160);
nand U15712 (N_15712,N_15457,N_15309);
and U15713 (N_15713,N_15125,N_15443);
xor U15714 (N_15714,N_15100,N_15151);
nor U15715 (N_15715,N_15265,N_15435);
nor U15716 (N_15716,N_15429,N_15242);
nand U15717 (N_15717,N_15095,N_15126);
and U15718 (N_15718,N_15357,N_15481);
nand U15719 (N_15719,N_15400,N_15302);
nor U15720 (N_15720,N_15033,N_15116);
or U15721 (N_15721,N_15065,N_15015);
nor U15722 (N_15722,N_15219,N_15441);
nor U15723 (N_15723,N_15119,N_15488);
or U15724 (N_15724,N_15281,N_15257);
xnor U15725 (N_15725,N_15350,N_15162);
and U15726 (N_15726,N_15486,N_15167);
nor U15727 (N_15727,N_15109,N_15072);
nor U15728 (N_15728,N_15016,N_15338);
nand U15729 (N_15729,N_15473,N_15420);
xnor U15730 (N_15730,N_15102,N_15465);
xnor U15731 (N_15731,N_15415,N_15478);
xnor U15732 (N_15732,N_15294,N_15406);
nor U15733 (N_15733,N_15396,N_15174);
nor U15734 (N_15734,N_15391,N_15283);
and U15735 (N_15735,N_15045,N_15182);
or U15736 (N_15736,N_15200,N_15479);
xor U15737 (N_15737,N_15256,N_15137);
nand U15738 (N_15738,N_15079,N_15158);
or U15739 (N_15739,N_15101,N_15430);
nor U15740 (N_15740,N_15041,N_15064);
or U15741 (N_15741,N_15135,N_15428);
or U15742 (N_15742,N_15073,N_15299);
xor U15743 (N_15743,N_15418,N_15241);
xor U15744 (N_15744,N_15487,N_15113);
or U15745 (N_15745,N_15496,N_15124);
xor U15746 (N_15746,N_15274,N_15273);
nor U15747 (N_15747,N_15398,N_15034);
nand U15748 (N_15748,N_15349,N_15090);
nor U15749 (N_15749,N_15186,N_15106);
nor U15750 (N_15750,N_15079,N_15348);
nand U15751 (N_15751,N_15287,N_15012);
nor U15752 (N_15752,N_15336,N_15442);
nand U15753 (N_15753,N_15305,N_15323);
and U15754 (N_15754,N_15248,N_15309);
nand U15755 (N_15755,N_15394,N_15332);
xor U15756 (N_15756,N_15326,N_15197);
or U15757 (N_15757,N_15372,N_15122);
nand U15758 (N_15758,N_15485,N_15080);
xor U15759 (N_15759,N_15426,N_15093);
nand U15760 (N_15760,N_15149,N_15486);
and U15761 (N_15761,N_15036,N_15025);
or U15762 (N_15762,N_15233,N_15057);
nor U15763 (N_15763,N_15341,N_15391);
nor U15764 (N_15764,N_15281,N_15304);
nand U15765 (N_15765,N_15088,N_15197);
or U15766 (N_15766,N_15285,N_15131);
nand U15767 (N_15767,N_15049,N_15221);
nand U15768 (N_15768,N_15343,N_15288);
xnor U15769 (N_15769,N_15005,N_15194);
nor U15770 (N_15770,N_15059,N_15418);
nand U15771 (N_15771,N_15402,N_15163);
or U15772 (N_15772,N_15339,N_15417);
xor U15773 (N_15773,N_15359,N_15427);
xnor U15774 (N_15774,N_15228,N_15435);
xnor U15775 (N_15775,N_15448,N_15375);
xor U15776 (N_15776,N_15395,N_15459);
and U15777 (N_15777,N_15365,N_15243);
and U15778 (N_15778,N_15117,N_15309);
or U15779 (N_15779,N_15220,N_15190);
xor U15780 (N_15780,N_15355,N_15489);
nor U15781 (N_15781,N_15420,N_15009);
nor U15782 (N_15782,N_15190,N_15140);
nand U15783 (N_15783,N_15167,N_15032);
nand U15784 (N_15784,N_15465,N_15044);
nor U15785 (N_15785,N_15282,N_15278);
or U15786 (N_15786,N_15257,N_15046);
nor U15787 (N_15787,N_15090,N_15469);
or U15788 (N_15788,N_15463,N_15383);
and U15789 (N_15789,N_15063,N_15208);
and U15790 (N_15790,N_15203,N_15276);
and U15791 (N_15791,N_15323,N_15329);
xor U15792 (N_15792,N_15303,N_15036);
nand U15793 (N_15793,N_15481,N_15269);
or U15794 (N_15794,N_15341,N_15040);
or U15795 (N_15795,N_15310,N_15135);
nor U15796 (N_15796,N_15163,N_15075);
and U15797 (N_15797,N_15080,N_15064);
nand U15798 (N_15798,N_15069,N_15331);
nand U15799 (N_15799,N_15311,N_15236);
nand U15800 (N_15800,N_15311,N_15369);
nor U15801 (N_15801,N_15446,N_15382);
nor U15802 (N_15802,N_15405,N_15080);
xnor U15803 (N_15803,N_15358,N_15206);
nand U15804 (N_15804,N_15000,N_15144);
nor U15805 (N_15805,N_15439,N_15380);
or U15806 (N_15806,N_15498,N_15351);
xnor U15807 (N_15807,N_15190,N_15299);
xnor U15808 (N_15808,N_15304,N_15120);
and U15809 (N_15809,N_15020,N_15277);
and U15810 (N_15810,N_15217,N_15231);
and U15811 (N_15811,N_15476,N_15003);
or U15812 (N_15812,N_15390,N_15159);
nor U15813 (N_15813,N_15108,N_15273);
or U15814 (N_15814,N_15113,N_15132);
or U15815 (N_15815,N_15035,N_15234);
and U15816 (N_15816,N_15282,N_15371);
xor U15817 (N_15817,N_15347,N_15422);
nor U15818 (N_15818,N_15299,N_15120);
and U15819 (N_15819,N_15497,N_15287);
nor U15820 (N_15820,N_15285,N_15426);
nand U15821 (N_15821,N_15038,N_15179);
nand U15822 (N_15822,N_15083,N_15443);
nor U15823 (N_15823,N_15253,N_15272);
or U15824 (N_15824,N_15449,N_15229);
or U15825 (N_15825,N_15082,N_15338);
or U15826 (N_15826,N_15083,N_15486);
or U15827 (N_15827,N_15134,N_15169);
and U15828 (N_15828,N_15171,N_15296);
or U15829 (N_15829,N_15284,N_15217);
nor U15830 (N_15830,N_15034,N_15208);
nand U15831 (N_15831,N_15076,N_15366);
xnor U15832 (N_15832,N_15417,N_15188);
nor U15833 (N_15833,N_15187,N_15401);
or U15834 (N_15834,N_15318,N_15180);
and U15835 (N_15835,N_15144,N_15128);
or U15836 (N_15836,N_15068,N_15011);
or U15837 (N_15837,N_15350,N_15482);
xor U15838 (N_15838,N_15232,N_15417);
nand U15839 (N_15839,N_15382,N_15125);
nor U15840 (N_15840,N_15173,N_15475);
nand U15841 (N_15841,N_15467,N_15317);
nor U15842 (N_15842,N_15146,N_15267);
or U15843 (N_15843,N_15007,N_15147);
or U15844 (N_15844,N_15264,N_15406);
nand U15845 (N_15845,N_15120,N_15405);
and U15846 (N_15846,N_15312,N_15489);
and U15847 (N_15847,N_15307,N_15227);
nor U15848 (N_15848,N_15364,N_15219);
or U15849 (N_15849,N_15191,N_15443);
xor U15850 (N_15850,N_15242,N_15334);
nand U15851 (N_15851,N_15468,N_15278);
or U15852 (N_15852,N_15134,N_15220);
or U15853 (N_15853,N_15255,N_15199);
nand U15854 (N_15854,N_15261,N_15257);
xnor U15855 (N_15855,N_15307,N_15184);
nor U15856 (N_15856,N_15123,N_15388);
or U15857 (N_15857,N_15019,N_15101);
nand U15858 (N_15858,N_15139,N_15302);
nand U15859 (N_15859,N_15283,N_15068);
nand U15860 (N_15860,N_15281,N_15406);
or U15861 (N_15861,N_15094,N_15007);
nor U15862 (N_15862,N_15202,N_15094);
nor U15863 (N_15863,N_15147,N_15053);
and U15864 (N_15864,N_15229,N_15245);
xor U15865 (N_15865,N_15291,N_15257);
or U15866 (N_15866,N_15356,N_15320);
xnor U15867 (N_15867,N_15452,N_15310);
or U15868 (N_15868,N_15314,N_15155);
nor U15869 (N_15869,N_15439,N_15297);
and U15870 (N_15870,N_15401,N_15439);
nor U15871 (N_15871,N_15222,N_15427);
or U15872 (N_15872,N_15482,N_15034);
or U15873 (N_15873,N_15100,N_15160);
and U15874 (N_15874,N_15496,N_15121);
and U15875 (N_15875,N_15184,N_15407);
nand U15876 (N_15876,N_15111,N_15396);
and U15877 (N_15877,N_15460,N_15439);
or U15878 (N_15878,N_15019,N_15195);
nor U15879 (N_15879,N_15278,N_15096);
nor U15880 (N_15880,N_15088,N_15427);
nand U15881 (N_15881,N_15148,N_15182);
or U15882 (N_15882,N_15029,N_15080);
nand U15883 (N_15883,N_15477,N_15348);
nand U15884 (N_15884,N_15234,N_15237);
or U15885 (N_15885,N_15138,N_15386);
nor U15886 (N_15886,N_15276,N_15159);
xnor U15887 (N_15887,N_15365,N_15317);
nand U15888 (N_15888,N_15361,N_15207);
nor U15889 (N_15889,N_15397,N_15239);
nand U15890 (N_15890,N_15054,N_15300);
nand U15891 (N_15891,N_15300,N_15365);
nor U15892 (N_15892,N_15223,N_15152);
nand U15893 (N_15893,N_15381,N_15044);
xnor U15894 (N_15894,N_15333,N_15290);
nand U15895 (N_15895,N_15216,N_15387);
or U15896 (N_15896,N_15496,N_15283);
and U15897 (N_15897,N_15043,N_15243);
or U15898 (N_15898,N_15353,N_15019);
nand U15899 (N_15899,N_15397,N_15166);
nand U15900 (N_15900,N_15285,N_15454);
nor U15901 (N_15901,N_15092,N_15199);
and U15902 (N_15902,N_15234,N_15443);
and U15903 (N_15903,N_15212,N_15253);
and U15904 (N_15904,N_15113,N_15008);
or U15905 (N_15905,N_15062,N_15327);
xnor U15906 (N_15906,N_15224,N_15346);
xor U15907 (N_15907,N_15114,N_15472);
or U15908 (N_15908,N_15027,N_15030);
xor U15909 (N_15909,N_15224,N_15210);
xor U15910 (N_15910,N_15479,N_15103);
nor U15911 (N_15911,N_15350,N_15212);
and U15912 (N_15912,N_15219,N_15333);
xor U15913 (N_15913,N_15298,N_15133);
or U15914 (N_15914,N_15066,N_15164);
xor U15915 (N_15915,N_15100,N_15148);
and U15916 (N_15916,N_15188,N_15203);
nor U15917 (N_15917,N_15040,N_15421);
and U15918 (N_15918,N_15231,N_15135);
nand U15919 (N_15919,N_15194,N_15415);
or U15920 (N_15920,N_15131,N_15448);
nand U15921 (N_15921,N_15497,N_15173);
and U15922 (N_15922,N_15000,N_15287);
nand U15923 (N_15923,N_15083,N_15383);
nor U15924 (N_15924,N_15264,N_15467);
xor U15925 (N_15925,N_15328,N_15064);
xor U15926 (N_15926,N_15308,N_15284);
xor U15927 (N_15927,N_15017,N_15463);
and U15928 (N_15928,N_15003,N_15317);
xnor U15929 (N_15929,N_15374,N_15161);
and U15930 (N_15930,N_15482,N_15241);
or U15931 (N_15931,N_15142,N_15192);
or U15932 (N_15932,N_15241,N_15006);
xnor U15933 (N_15933,N_15224,N_15109);
and U15934 (N_15934,N_15208,N_15024);
nor U15935 (N_15935,N_15007,N_15172);
or U15936 (N_15936,N_15239,N_15292);
xnor U15937 (N_15937,N_15151,N_15282);
and U15938 (N_15938,N_15445,N_15285);
nor U15939 (N_15939,N_15266,N_15343);
nor U15940 (N_15940,N_15431,N_15393);
nand U15941 (N_15941,N_15318,N_15068);
and U15942 (N_15942,N_15363,N_15438);
nor U15943 (N_15943,N_15057,N_15201);
nor U15944 (N_15944,N_15205,N_15186);
xnor U15945 (N_15945,N_15145,N_15439);
and U15946 (N_15946,N_15321,N_15306);
nor U15947 (N_15947,N_15408,N_15478);
or U15948 (N_15948,N_15155,N_15191);
and U15949 (N_15949,N_15189,N_15251);
xor U15950 (N_15950,N_15418,N_15452);
or U15951 (N_15951,N_15092,N_15128);
or U15952 (N_15952,N_15234,N_15009);
and U15953 (N_15953,N_15061,N_15176);
xor U15954 (N_15954,N_15475,N_15464);
nand U15955 (N_15955,N_15389,N_15090);
nand U15956 (N_15956,N_15460,N_15320);
and U15957 (N_15957,N_15055,N_15489);
nand U15958 (N_15958,N_15247,N_15132);
xnor U15959 (N_15959,N_15365,N_15235);
and U15960 (N_15960,N_15301,N_15117);
nand U15961 (N_15961,N_15055,N_15294);
and U15962 (N_15962,N_15058,N_15222);
xor U15963 (N_15963,N_15420,N_15237);
or U15964 (N_15964,N_15301,N_15483);
and U15965 (N_15965,N_15460,N_15304);
or U15966 (N_15966,N_15045,N_15062);
nor U15967 (N_15967,N_15265,N_15174);
nor U15968 (N_15968,N_15436,N_15347);
or U15969 (N_15969,N_15411,N_15242);
and U15970 (N_15970,N_15376,N_15121);
or U15971 (N_15971,N_15063,N_15493);
nand U15972 (N_15972,N_15329,N_15455);
nor U15973 (N_15973,N_15146,N_15327);
nor U15974 (N_15974,N_15318,N_15399);
nand U15975 (N_15975,N_15481,N_15426);
or U15976 (N_15976,N_15248,N_15443);
nand U15977 (N_15977,N_15380,N_15080);
nand U15978 (N_15978,N_15294,N_15489);
and U15979 (N_15979,N_15426,N_15027);
nor U15980 (N_15980,N_15144,N_15067);
xnor U15981 (N_15981,N_15004,N_15001);
xnor U15982 (N_15982,N_15426,N_15320);
nand U15983 (N_15983,N_15252,N_15345);
or U15984 (N_15984,N_15168,N_15295);
xnor U15985 (N_15985,N_15440,N_15003);
nor U15986 (N_15986,N_15290,N_15383);
or U15987 (N_15987,N_15238,N_15142);
nand U15988 (N_15988,N_15427,N_15282);
nand U15989 (N_15989,N_15056,N_15423);
and U15990 (N_15990,N_15363,N_15216);
nor U15991 (N_15991,N_15033,N_15491);
nand U15992 (N_15992,N_15282,N_15415);
or U15993 (N_15993,N_15185,N_15289);
and U15994 (N_15994,N_15304,N_15252);
nand U15995 (N_15995,N_15324,N_15238);
xnor U15996 (N_15996,N_15489,N_15304);
or U15997 (N_15997,N_15201,N_15251);
and U15998 (N_15998,N_15118,N_15485);
nand U15999 (N_15999,N_15056,N_15405);
nand U16000 (N_16000,N_15571,N_15668);
nor U16001 (N_16001,N_15894,N_15904);
nand U16002 (N_16002,N_15922,N_15699);
or U16003 (N_16003,N_15909,N_15930);
nand U16004 (N_16004,N_15959,N_15993);
xor U16005 (N_16005,N_15765,N_15523);
nand U16006 (N_16006,N_15992,N_15578);
nor U16007 (N_16007,N_15961,N_15733);
or U16008 (N_16008,N_15554,N_15677);
and U16009 (N_16009,N_15689,N_15574);
xor U16010 (N_16010,N_15624,N_15817);
xor U16011 (N_16011,N_15755,N_15852);
and U16012 (N_16012,N_15715,N_15708);
and U16013 (N_16013,N_15600,N_15845);
nor U16014 (N_16014,N_15623,N_15996);
nand U16015 (N_16015,N_15550,N_15823);
nand U16016 (N_16016,N_15582,N_15692);
or U16017 (N_16017,N_15786,N_15972);
nand U16018 (N_16018,N_15512,N_15934);
and U16019 (N_16019,N_15566,N_15591);
or U16020 (N_16020,N_15772,N_15644);
nand U16021 (N_16021,N_15585,N_15545);
nor U16022 (N_16022,N_15954,N_15868);
and U16023 (N_16023,N_15581,N_15667);
nor U16024 (N_16024,N_15962,N_15750);
nand U16025 (N_16025,N_15670,N_15769);
xor U16026 (N_16026,N_15734,N_15590);
and U16027 (N_16027,N_15988,N_15595);
xnor U16028 (N_16028,N_15925,N_15560);
xor U16029 (N_16029,N_15604,N_15806);
and U16030 (N_16030,N_15913,N_15849);
nor U16031 (N_16031,N_15530,N_15830);
nand U16032 (N_16032,N_15814,N_15982);
nand U16033 (N_16033,N_15980,N_15914);
or U16034 (N_16034,N_15874,N_15851);
or U16035 (N_16035,N_15520,N_15757);
nor U16036 (N_16036,N_15516,N_15698);
and U16037 (N_16037,N_15907,N_15746);
nor U16038 (N_16038,N_15740,N_15657);
and U16039 (N_16039,N_15716,N_15597);
or U16040 (N_16040,N_15609,N_15977);
or U16041 (N_16041,N_15879,N_15727);
xor U16042 (N_16042,N_15885,N_15599);
nand U16043 (N_16043,N_15989,N_15707);
or U16044 (N_16044,N_15602,N_15529);
nor U16045 (N_16045,N_15758,N_15569);
xor U16046 (N_16046,N_15944,N_15941);
xnor U16047 (N_16047,N_15684,N_15556);
or U16048 (N_16048,N_15901,N_15762);
and U16049 (N_16049,N_15735,N_15694);
xor U16050 (N_16050,N_15853,N_15918);
or U16051 (N_16051,N_15808,N_15829);
xnor U16052 (N_16052,N_15717,N_15606);
and U16053 (N_16053,N_15946,N_15553);
xnor U16054 (N_16054,N_15513,N_15741);
and U16055 (N_16055,N_15561,N_15981);
xor U16056 (N_16056,N_15620,N_15932);
nand U16057 (N_16057,N_15552,N_15598);
nor U16058 (N_16058,N_15701,N_15749);
or U16059 (N_16059,N_15860,N_15754);
xor U16060 (N_16060,N_15965,N_15908);
and U16061 (N_16061,N_15985,N_15917);
or U16062 (N_16062,N_15821,N_15618);
or U16063 (N_16063,N_15899,N_15664);
nor U16064 (N_16064,N_15945,N_15564);
and U16065 (N_16065,N_15938,N_15942);
or U16066 (N_16066,N_15820,N_15632);
or U16067 (N_16067,N_15905,N_15887);
xnor U16068 (N_16068,N_15546,N_15575);
and U16069 (N_16069,N_15898,N_15880);
nor U16070 (N_16070,N_15589,N_15953);
xor U16071 (N_16071,N_15858,N_15654);
xnor U16072 (N_16072,N_15936,N_15973);
nand U16073 (N_16073,N_15866,N_15680);
nand U16074 (N_16074,N_15994,N_15825);
xor U16075 (N_16075,N_15524,N_15948);
nand U16076 (N_16076,N_15882,N_15779);
xnor U16077 (N_16077,N_15537,N_15759);
xor U16078 (N_16078,N_15738,N_15801);
xnor U16079 (N_16079,N_15943,N_15864);
nor U16080 (N_16080,N_15967,N_15838);
and U16081 (N_16081,N_15645,N_15607);
nand U16082 (N_16082,N_15966,N_15819);
or U16083 (N_16083,N_15951,N_15834);
nand U16084 (N_16084,N_15573,N_15731);
xnor U16085 (N_16085,N_15651,N_15924);
xnor U16086 (N_16086,N_15650,N_15842);
and U16087 (N_16087,N_15789,N_15862);
nand U16088 (N_16088,N_15509,N_15710);
nand U16089 (N_16089,N_15696,N_15826);
and U16090 (N_16090,N_15824,N_15565);
or U16091 (N_16091,N_15562,N_15592);
or U16092 (N_16092,N_15760,N_15969);
xnor U16093 (N_16093,N_15676,N_15614);
nand U16094 (N_16094,N_15732,N_15683);
and U16095 (N_16095,N_15777,N_15888);
nand U16096 (N_16096,N_15510,N_15911);
and U16097 (N_16097,N_15791,N_15563);
or U16098 (N_16098,N_15856,N_15940);
nand U16099 (N_16099,N_15807,N_15847);
nor U16100 (N_16100,N_15616,N_15634);
xor U16101 (N_16101,N_15773,N_15661);
and U16102 (N_16102,N_15896,N_15517);
nor U16103 (N_16103,N_15502,N_15892);
nand U16104 (N_16104,N_15625,N_15926);
nand U16105 (N_16105,N_15764,N_15870);
xnor U16106 (N_16106,N_15884,N_15691);
or U16107 (N_16107,N_15827,N_15712);
and U16108 (N_16108,N_15997,N_15690);
nand U16109 (N_16109,N_15580,N_15627);
nand U16110 (N_16110,N_15975,N_15906);
and U16111 (N_16111,N_15526,N_15729);
nand U16112 (N_16112,N_15635,N_15637);
and U16113 (N_16113,N_15970,N_15718);
nand U16114 (N_16114,N_15538,N_15653);
or U16115 (N_16115,N_15893,N_15877);
nand U16116 (N_16116,N_15688,N_15572);
nor U16117 (N_16117,N_15568,N_15804);
xnor U16118 (N_16118,N_15636,N_15728);
or U16119 (N_16119,N_15920,N_15532);
and U16120 (N_16120,N_15881,N_15611);
xor U16121 (N_16121,N_15551,N_15781);
or U16122 (N_16122,N_15547,N_15802);
nand U16123 (N_16123,N_15780,N_15531);
nor U16124 (N_16124,N_15872,N_15792);
nor U16125 (N_16125,N_15675,N_15919);
or U16126 (N_16126,N_15837,N_15835);
xor U16127 (N_16127,N_15915,N_15711);
nor U16128 (N_16128,N_15730,N_15744);
nor U16129 (N_16129,N_15947,N_15841);
and U16130 (N_16130,N_15846,N_15643);
nand U16131 (N_16131,N_15557,N_15739);
xnor U16132 (N_16132,N_15671,N_15833);
and U16133 (N_16133,N_15534,N_15533);
or U16134 (N_16134,N_15640,N_15987);
and U16135 (N_16135,N_15844,N_15900);
xor U16136 (N_16136,N_15998,N_15986);
or U16137 (N_16137,N_15923,N_15593);
and U16138 (N_16138,N_15794,N_15639);
nor U16139 (N_16139,N_15971,N_15891);
and U16140 (N_16140,N_15912,N_15790);
nand U16141 (N_16141,N_15958,N_15742);
xor U16142 (N_16142,N_15748,N_15652);
and U16143 (N_16143,N_15687,N_15500);
nand U16144 (N_16144,N_15766,N_15787);
xnor U16145 (N_16145,N_15700,N_15873);
xnor U16146 (N_16146,N_15605,N_15559);
or U16147 (N_16147,N_15519,N_15935);
nand U16148 (N_16148,N_15803,N_15666);
nand U16149 (N_16149,N_15782,N_15703);
or U16150 (N_16150,N_15867,N_15719);
nand U16151 (N_16151,N_15647,N_15577);
nor U16152 (N_16152,N_15642,N_15695);
nor U16153 (N_16153,N_15929,N_15674);
xor U16154 (N_16154,N_15515,N_15927);
and U16155 (N_16155,N_15843,N_15999);
or U16156 (N_16156,N_15567,N_15747);
nor U16157 (N_16157,N_15793,N_15974);
xor U16158 (N_16158,N_15736,N_15505);
and U16159 (N_16159,N_15672,N_15558);
xnor U16160 (N_16160,N_15536,N_15724);
and U16161 (N_16161,N_15576,N_15641);
and U16162 (N_16162,N_15697,N_15673);
nor U16163 (N_16163,N_15839,N_15615);
nor U16164 (N_16164,N_15704,N_15596);
nor U16165 (N_16165,N_15983,N_15933);
nand U16166 (N_16166,N_15548,N_15895);
or U16167 (N_16167,N_15756,N_15539);
xnor U16168 (N_16168,N_15528,N_15706);
xnor U16169 (N_16169,N_15795,N_15737);
xor U16170 (N_16170,N_15767,N_15950);
nand U16171 (N_16171,N_15937,N_15543);
and U16172 (N_16172,N_15809,N_15612);
nand U16173 (N_16173,N_15541,N_15656);
nand U16174 (N_16174,N_15584,N_15631);
xnor U16175 (N_16175,N_15610,N_15963);
nand U16176 (N_16176,N_15726,N_15840);
xnor U16177 (N_16177,N_15797,N_15869);
nor U16178 (N_16178,N_15660,N_15836);
or U16179 (N_16179,N_15633,N_15832);
and U16180 (N_16180,N_15861,N_15669);
or U16181 (N_16181,N_15810,N_15507);
nor U16182 (N_16182,N_15679,N_15685);
nand U16183 (N_16183,N_15800,N_15630);
and U16184 (N_16184,N_15902,N_15702);
nand U16185 (N_16185,N_15865,N_15527);
nor U16186 (N_16186,N_15990,N_15848);
or U16187 (N_16187,N_15626,N_15745);
and U16188 (N_16188,N_15681,N_15956);
xor U16189 (N_16189,N_15788,N_15763);
xor U16190 (N_16190,N_15928,N_15608);
nor U16191 (N_16191,N_15751,N_15952);
and U16192 (N_16192,N_15686,N_15783);
nor U16193 (N_16193,N_15659,N_15812);
nand U16194 (N_16194,N_15770,N_15722);
and U16195 (N_16195,N_15535,N_15663);
nand U16196 (N_16196,N_15621,N_15822);
or U16197 (N_16197,N_15854,N_15949);
or U16198 (N_16198,N_15886,N_15709);
xnor U16199 (N_16199,N_15579,N_15613);
and U16200 (N_16200,N_15542,N_15622);
nor U16201 (N_16201,N_15544,N_15713);
and U16202 (N_16202,N_15776,N_15752);
or U16203 (N_16203,N_15525,N_15658);
xnor U16204 (N_16204,N_15850,N_15628);
nand U16205 (N_16205,N_15501,N_15811);
and U16206 (N_16206,N_15883,N_15518);
nor U16207 (N_16207,N_15646,N_15720);
xor U16208 (N_16208,N_15693,N_15761);
xor U16209 (N_16209,N_15863,N_15522);
and U16210 (N_16210,N_15890,N_15775);
and U16211 (N_16211,N_15678,N_15910);
nand U16212 (N_16212,N_15875,N_15831);
and U16213 (N_16213,N_15504,N_15705);
xnor U16214 (N_16214,N_15968,N_15508);
or U16215 (N_16215,N_15665,N_15594);
xor U16216 (N_16216,N_15995,N_15784);
nand U16217 (N_16217,N_15503,N_15603);
xnor U16218 (N_16218,N_15799,N_15601);
nand U16219 (N_16219,N_15897,N_15976);
nor U16220 (N_16220,N_15655,N_15916);
nand U16221 (N_16221,N_15813,N_15774);
xor U16222 (N_16222,N_15768,N_15723);
or U16223 (N_16223,N_15521,N_15818);
and U16224 (N_16224,N_15805,N_15978);
xor U16225 (N_16225,N_15984,N_15828);
xor U16226 (N_16226,N_15991,N_15960);
xor U16227 (N_16227,N_15549,N_15796);
nand U16228 (N_16228,N_15682,N_15583);
and U16229 (N_16229,N_15648,N_15955);
or U16230 (N_16230,N_15876,N_15815);
xor U16231 (N_16231,N_15514,N_15964);
nor U16232 (N_16232,N_15570,N_15859);
or U16233 (N_16233,N_15778,N_15931);
nor U16234 (N_16234,N_15511,N_15889);
nor U16235 (N_16235,N_15587,N_15638);
nand U16236 (N_16236,N_15588,N_15540);
nor U16237 (N_16237,N_15878,N_15555);
and U16238 (N_16238,N_15662,N_15721);
and U16239 (N_16239,N_15771,N_15921);
or U16240 (N_16240,N_15586,N_15939);
and U16241 (N_16241,N_15957,N_15506);
nand U16242 (N_16242,N_15743,N_15855);
and U16243 (N_16243,N_15725,N_15798);
nor U16244 (N_16244,N_15753,N_15857);
and U16245 (N_16245,N_15619,N_15649);
or U16246 (N_16246,N_15979,N_15903);
nand U16247 (N_16247,N_15714,N_15871);
xor U16248 (N_16248,N_15785,N_15629);
nor U16249 (N_16249,N_15617,N_15816);
xnor U16250 (N_16250,N_15621,N_15973);
or U16251 (N_16251,N_15610,N_15662);
xor U16252 (N_16252,N_15689,N_15806);
or U16253 (N_16253,N_15852,N_15966);
nor U16254 (N_16254,N_15782,N_15758);
nand U16255 (N_16255,N_15709,N_15695);
nand U16256 (N_16256,N_15993,N_15593);
nor U16257 (N_16257,N_15769,N_15970);
or U16258 (N_16258,N_15512,N_15508);
and U16259 (N_16259,N_15971,N_15796);
nor U16260 (N_16260,N_15848,N_15933);
or U16261 (N_16261,N_15519,N_15524);
nor U16262 (N_16262,N_15635,N_15723);
or U16263 (N_16263,N_15810,N_15865);
nand U16264 (N_16264,N_15840,N_15807);
and U16265 (N_16265,N_15650,N_15766);
or U16266 (N_16266,N_15809,N_15920);
nand U16267 (N_16267,N_15777,N_15580);
nand U16268 (N_16268,N_15633,N_15741);
nor U16269 (N_16269,N_15555,N_15567);
nor U16270 (N_16270,N_15806,N_15664);
xnor U16271 (N_16271,N_15648,N_15882);
nor U16272 (N_16272,N_15709,N_15970);
nand U16273 (N_16273,N_15604,N_15736);
or U16274 (N_16274,N_15997,N_15819);
xnor U16275 (N_16275,N_15848,N_15979);
and U16276 (N_16276,N_15873,N_15851);
xor U16277 (N_16277,N_15929,N_15721);
and U16278 (N_16278,N_15798,N_15770);
nand U16279 (N_16279,N_15506,N_15581);
nor U16280 (N_16280,N_15873,N_15704);
xnor U16281 (N_16281,N_15704,N_15612);
or U16282 (N_16282,N_15889,N_15717);
xor U16283 (N_16283,N_15810,N_15612);
nor U16284 (N_16284,N_15892,N_15609);
xnor U16285 (N_16285,N_15942,N_15901);
or U16286 (N_16286,N_15906,N_15884);
or U16287 (N_16287,N_15938,N_15935);
nor U16288 (N_16288,N_15998,N_15529);
nor U16289 (N_16289,N_15654,N_15749);
or U16290 (N_16290,N_15769,N_15510);
nand U16291 (N_16291,N_15912,N_15638);
and U16292 (N_16292,N_15751,N_15839);
xnor U16293 (N_16293,N_15614,N_15734);
nand U16294 (N_16294,N_15852,N_15830);
nor U16295 (N_16295,N_15810,N_15750);
nand U16296 (N_16296,N_15682,N_15613);
nor U16297 (N_16297,N_15950,N_15769);
or U16298 (N_16298,N_15686,N_15813);
nand U16299 (N_16299,N_15838,N_15544);
and U16300 (N_16300,N_15567,N_15545);
nor U16301 (N_16301,N_15928,N_15820);
nand U16302 (N_16302,N_15916,N_15635);
or U16303 (N_16303,N_15862,N_15618);
and U16304 (N_16304,N_15830,N_15652);
xor U16305 (N_16305,N_15668,N_15639);
nor U16306 (N_16306,N_15537,N_15943);
nor U16307 (N_16307,N_15697,N_15687);
or U16308 (N_16308,N_15747,N_15837);
and U16309 (N_16309,N_15940,N_15613);
or U16310 (N_16310,N_15506,N_15693);
or U16311 (N_16311,N_15789,N_15801);
xor U16312 (N_16312,N_15611,N_15692);
or U16313 (N_16313,N_15777,N_15774);
nand U16314 (N_16314,N_15785,N_15586);
and U16315 (N_16315,N_15652,N_15788);
nor U16316 (N_16316,N_15696,N_15766);
nor U16317 (N_16317,N_15523,N_15891);
nor U16318 (N_16318,N_15535,N_15876);
or U16319 (N_16319,N_15783,N_15725);
xnor U16320 (N_16320,N_15982,N_15889);
nand U16321 (N_16321,N_15789,N_15644);
xnor U16322 (N_16322,N_15548,N_15522);
and U16323 (N_16323,N_15593,N_15796);
nand U16324 (N_16324,N_15629,N_15924);
or U16325 (N_16325,N_15687,N_15512);
nor U16326 (N_16326,N_15821,N_15557);
and U16327 (N_16327,N_15898,N_15638);
xor U16328 (N_16328,N_15772,N_15805);
or U16329 (N_16329,N_15594,N_15619);
or U16330 (N_16330,N_15731,N_15921);
and U16331 (N_16331,N_15713,N_15586);
or U16332 (N_16332,N_15751,N_15594);
nand U16333 (N_16333,N_15584,N_15952);
or U16334 (N_16334,N_15557,N_15504);
and U16335 (N_16335,N_15748,N_15727);
nor U16336 (N_16336,N_15837,N_15609);
or U16337 (N_16337,N_15812,N_15875);
nand U16338 (N_16338,N_15622,N_15611);
nand U16339 (N_16339,N_15931,N_15923);
nand U16340 (N_16340,N_15614,N_15768);
or U16341 (N_16341,N_15790,N_15982);
nor U16342 (N_16342,N_15996,N_15609);
nor U16343 (N_16343,N_15794,N_15759);
and U16344 (N_16344,N_15780,N_15669);
or U16345 (N_16345,N_15938,N_15554);
or U16346 (N_16346,N_15628,N_15530);
or U16347 (N_16347,N_15761,N_15824);
nand U16348 (N_16348,N_15650,N_15664);
and U16349 (N_16349,N_15819,N_15516);
nand U16350 (N_16350,N_15729,N_15504);
xor U16351 (N_16351,N_15550,N_15922);
xor U16352 (N_16352,N_15915,N_15560);
xnor U16353 (N_16353,N_15923,N_15963);
nor U16354 (N_16354,N_15614,N_15702);
nor U16355 (N_16355,N_15669,N_15613);
or U16356 (N_16356,N_15809,N_15505);
and U16357 (N_16357,N_15684,N_15967);
nor U16358 (N_16358,N_15707,N_15594);
nand U16359 (N_16359,N_15729,N_15533);
or U16360 (N_16360,N_15768,N_15786);
or U16361 (N_16361,N_15787,N_15982);
or U16362 (N_16362,N_15945,N_15719);
or U16363 (N_16363,N_15799,N_15834);
and U16364 (N_16364,N_15841,N_15552);
and U16365 (N_16365,N_15932,N_15809);
nor U16366 (N_16366,N_15710,N_15562);
or U16367 (N_16367,N_15694,N_15838);
nand U16368 (N_16368,N_15705,N_15823);
or U16369 (N_16369,N_15731,N_15595);
or U16370 (N_16370,N_15547,N_15563);
nand U16371 (N_16371,N_15689,N_15905);
nand U16372 (N_16372,N_15625,N_15780);
or U16373 (N_16373,N_15761,N_15652);
nand U16374 (N_16374,N_15571,N_15957);
or U16375 (N_16375,N_15801,N_15713);
nand U16376 (N_16376,N_15886,N_15960);
xnor U16377 (N_16377,N_15549,N_15525);
or U16378 (N_16378,N_15666,N_15976);
xnor U16379 (N_16379,N_15652,N_15976);
nor U16380 (N_16380,N_15566,N_15654);
nand U16381 (N_16381,N_15689,N_15772);
and U16382 (N_16382,N_15880,N_15775);
xnor U16383 (N_16383,N_15743,N_15627);
nor U16384 (N_16384,N_15557,N_15755);
or U16385 (N_16385,N_15845,N_15821);
or U16386 (N_16386,N_15577,N_15568);
nor U16387 (N_16387,N_15613,N_15510);
nand U16388 (N_16388,N_15780,N_15837);
and U16389 (N_16389,N_15618,N_15913);
nand U16390 (N_16390,N_15890,N_15611);
nor U16391 (N_16391,N_15623,N_15926);
nand U16392 (N_16392,N_15684,N_15723);
nand U16393 (N_16393,N_15716,N_15923);
and U16394 (N_16394,N_15643,N_15991);
xnor U16395 (N_16395,N_15701,N_15631);
and U16396 (N_16396,N_15975,N_15662);
nand U16397 (N_16397,N_15689,N_15935);
nor U16398 (N_16398,N_15633,N_15663);
nor U16399 (N_16399,N_15965,N_15888);
nand U16400 (N_16400,N_15956,N_15992);
nand U16401 (N_16401,N_15942,N_15945);
or U16402 (N_16402,N_15585,N_15577);
xor U16403 (N_16403,N_15734,N_15934);
or U16404 (N_16404,N_15816,N_15969);
xor U16405 (N_16405,N_15661,N_15563);
or U16406 (N_16406,N_15987,N_15574);
and U16407 (N_16407,N_15764,N_15564);
and U16408 (N_16408,N_15869,N_15824);
or U16409 (N_16409,N_15662,N_15503);
or U16410 (N_16410,N_15914,N_15814);
or U16411 (N_16411,N_15943,N_15992);
nor U16412 (N_16412,N_15717,N_15879);
xor U16413 (N_16413,N_15818,N_15975);
nor U16414 (N_16414,N_15608,N_15692);
or U16415 (N_16415,N_15682,N_15962);
and U16416 (N_16416,N_15590,N_15640);
and U16417 (N_16417,N_15981,N_15929);
and U16418 (N_16418,N_15578,N_15923);
nand U16419 (N_16419,N_15913,N_15526);
or U16420 (N_16420,N_15568,N_15547);
nor U16421 (N_16421,N_15950,N_15740);
nor U16422 (N_16422,N_15897,N_15510);
or U16423 (N_16423,N_15910,N_15868);
nor U16424 (N_16424,N_15984,N_15885);
or U16425 (N_16425,N_15969,N_15860);
nand U16426 (N_16426,N_15999,N_15973);
and U16427 (N_16427,N_15910,N_15859);
nand U16428 (N_16428,N_15951,N_15590);
xnor U16429 (N_16429,N_15792,N_15809);
and U16430 (N_16430,N_15682,N_15732);
nand U16431 (N_16431,N_15793,N_15853);
or U16432 (N_16432,N_15899,N_15615);
nor U16433 (N_16433,N_15531,N_15837);
or U16434 (N_16434,N_15547,N_15966);
or U16435 (N_16435,N_15848,N_15905);
xnor U16436 (N_16436,N_15516,N_15858);
or U16437 (N_16437,N_15589,N_15806);
nand U16438 (N_16438,N_15992,N_15724);
nor U16439 (N_16439,N_15785,N_15559);
and U16440 (N_16440,N_15736,N_15925);
or U16441 (N_16441,N_15983,N_15757);
xnor U16442 (N_16442,N_15986,N_15628);
nand U16443 (N_16443,N_15689,N_15910);
and U16444 (N_16444,N_15844,N_15569);
and U16445 (N_16445,N_15654,N_15700);
or U16446 (N_16446,N_15972,N_15945);
or U16447 (N_16447,N_15534,N_15747);
xnor U16448 (N_16448,N_15542,N_15522);
and U16449 (N_16449,N_15951,N_15940);
xnor U16450 (N_16450,N_15768,N_15639);
or U16451 (N_16451,N_15664,N_15961);
or U16452 (N_16452,N_15894,N_15836);
and U16453 (N_16453,N_15914,N_15677);
or U16454 (N_16454,N_15969,N_15500);
xor U16455 (N_16455,N_15969,N_15670);
nand U16456 (N_16456,N_15775,N_15958);
xnor U16457 (N_16457,N_15832,N_15988);
nor U16458 (N_16458,N_15850,N_15538);
and U16459 (N_16459,N_15926,N_15810);
nor U16460 (N_16460,N_15635,N_15983);
nor U16461 (N_16461,N_15926,N_15522);
nand U16462 (N_16462,N_15739,N_15620);
nor U16463 (N_16463,N_15716,N_15963);
nand U16464 (N_16464,N_15523,N_15804);
and U16465 (N_16465,N_15843,N_15838);
xnor U16466 (N_16466,N_15631,N_15764);
and U16467 (N_16467,N_15649,N_15526);
and U16468 (N_16468,N_15937,N_15662);
or U16469 (N_16469,N_15927,N_15674);
or U16470 (N_16470,N_15804,N_15836);
or U16471 (N_16471,N_15672,N_15525);
nor U16472 (N_16472,N_15822,N_15991);
or U16473 (N_16473,N_15553,N_15719);
or U16474 (N_16474,N_15821,N_15609);
xor U16475 (N_16475,N_15529,N_15939);
or U16476 (N_16476,N_15528,N_15535);
and U16477 (N_16477,N_15657,N_15689);
nor U16478 (N_16478,N_15801,N_15702);
and U16479 (N_16479,N_15903,N_15725);
xor U16480 (N_16480,N_15921,N_15859);
nor U16481 (N_16481,N_15980,N_15800);
xnor U16482 (N_16482,N_15636,N_15781);
xnor U16483 (N_16483,N_15562,N_15703);
xor U16484 (N_16484,N_15841,N_15764);
or U16485 (N_16485,N_15743,N_15568);
and U16486 (N_16486,N_15688,N_15660);
xnor U16487 (N_16487,N_15576,N_15502);
nor U16488 (N_16488,N_15833,N_15816);
or U16489 (N_16489,N_15535,N_15609);
or U16490 (N_16490,N_15972,N_15572);
or U16491 (N_16491,N_15677,N_15585);
xor U16492 (N_16492,N_15991,N_15522);
xor U16493 (N_16493,N_15582,N_15763);
nand U16494 (N_16494,N_15942,N_15992);
nor U16495 (N_16495,N_15624,N_15941);
xnor U16496 (N_16496,N_15724,N_15808);
xnor U16497 (N_16497,N_15754,N_15799);
and U16498 (N_16498,N_15736,N_15528);
xnor U16499 (N_16499,N_15847,N_15983);
nor U16500 (N_16500,N_16096,N_16040);
or U16501 (N_16501,N_16154,N_16289);
or U16502 (N_16502,N_16002,N_16133);
nor U16503 (N_16503,N_16212,N_16259);
nor U16504 (N_16504,N_16182,N_16023);
xnor U16505 (N_16505,N_16013,N_16239);
or U16506 (N_16506,N_16304,N_16037);
and U16507 (N_16507,N_16418,N_16063);
and U16508 (N_16508,N_16277,N_16088);
xor U16509 (N_16509,N_16399,N_16221);
nor U16510 (N_16510,N_16426,N_16347);
and U16511 (N_16511,N_16059,N_16439);
nor U16512 (N_16512,N_16476,N_16288);
or U16513 (N_16513,N_16338,N_16444);
and U16514 (N_16514,N_16472,N_16329);
xor U16515 (N_16515,N_16339,N_16163);
or U16516 (N_16516,N_16169,N_16460);
or U16517 (N_16517,N_16480,N_16084);
nor U16518 (N_16518,N_16126,N_16451);
or U16519 (N_16519,N_16072,N_16113);
xor U16520 (N_16520,N_16227,N_16408);
and U16521 (N_16521,N_16380,N_16136);
nand U16522 (N_16522,N_16211,N_16092);
xor U16523 (N_16523,N_16081,N_16103);
xor U16524 (N_16524,N_16381,N_16434);
xor U16525 (N_16525,N_16209,N_16085);
and U16526 (N_16526,N_16078,N_16445);
xnor U16527 (N_16527,N_16473,N_16387);
or U16528 (N_16528,N_16033,N_16178);
and U16529 (N_16529,N_16274,N_16406);
xnor U16530 (N_16530,N_16176,N_16374);
nand U16531 (N_16531,N_16159,N_16352);
xor U16532 (N_16532,N_16315,N_16093);
nor U16533 (N_16533,N_16357,N_16291);
nor U16534 (N_16534,N_16252,N_16055);
nand U16535 (N_16535,N_16061,N_16264);
and U16536 (N_16536,N_16022,N_16272);
xor U16537 (N_16537,N_16430,N_16358);
and U16538 (N_16538,N_16342,N_16341);
xnor U16539 (N_16539,N_16064,N_16496);
xnor U16540 (N_16540,N_16197,N_16349);
xor U16541 (N_16541,N_16371,N_16125);
nand U16542 (N_16542,N_16089,N_16309);
nand U16543 (N_16543,N_16435,N_16008);
nand U16544 (N_16544,N_16213,N_16364);
xnor U16545 (N_16545,N_16330,N_16384);
xnor U16546 (N_16546,N_16215,N_16124);
and U16547 (N_16547,N_16390,N_16208);
nor U16548 (N_16548,N_16074,N_16242);
and U16549 (N_16549,N_16255,N_16484);
nor U16550 (N_16550,N_16433,N_16017);
or U16551 (N_16551,N_16253,N_16251);
and U16552 (N_16552,N_16437,N_16118);
nor U16553 (N_16553,N_16366,N_16455);
nand U16554 (N_16554,N_16094,N_16372);
xor U16555 (N_16555,N_16312,N_16230);
nor U16556 (N_16556,N_16132,N_16150);
and U16557 (N_16557,N_16448,N_16145);
xor U16558 (N_16558,N_16207,N_16417);
and U16559 (N_16559,N_16443,N_16121);
nor U16560 (N_16560,N_16482,N_16248);
and U16561 (N_16561,N_16488,N_16232);
nor U16562 (N_16562,N_16343,N_16117);
nor U16563 (N_16563,N_16224,N_16471);
nand U16564 (N_16564,N_16246,N_16412);
nor U16565 (N_16565,N_16367,N_16317);
xor U16566 (N_16566,N_16183,N_16225);
or U16567 (N_16567,N_16337,N_16062);
or U16568 (N_16568,N_16051,N_16407);
nor U16569 (N_16569,N_16286,N_16243);
or U16570 (N_16570,N_16271,N_16067);
xor U16571 (N_16571,N_16446,N_16324);
xnor U16572 (N_16572,N_16346,N_16254);
or U16573 (N_16573,N_16100,N_16079);
and U16574 (N_16574,N_16293,N_16007);
nor U16575 (N_16575,N_16466,N_16438);
or U16576 (N_16576,N_16097,N_16368);
nand U16577 (N_16577,N_16127,N_16416);
xor U16578 (N_16578,N_16414,N_16319);
nor U16579 (N_16579,N_16415,N_16091);
nand U16580 (N_16580,N_16283,N_16042);
xor U16581 (N_16581,N_16423,N_16427);
nand U16582 (N_16582,N_16160,N_16030);
or U16583 (N_16583,N_16395,N_16205);
xor U16584 (N_16584,N_16158,N_16181);
nor U16585 (N_16585,N_16202,N_16499);
and U16586 (N_16586,N_16192,N_16486);
and U16587 (N_16587,N_16413,N_16226);
xor U16588 (N_16588,N_16168,N_16191);
nor U16589 (N_16589,N_16070,N_16012);
xnor U16590 (N_16590,N_16333,N_16497);
xor U16591 (N_16591,N_16234,N_16032);
xor U16592 (N_16592,N_16186,N_16273);
xnor U16593 (N_16593,N_16392,N_16465);
xnor U16594 (N_16594,N_16140,N_16015);
nand U16595 (N_16595,N_16355,N_16184);
xnor U16596 (N_16596,N_16004,N_16470);
xnor U16597 (N_16597,N_16441,N_16231);
or U16598 (N_16598,N_16328,N_16491);
or U16599 (N_16599,N_16490,N_16398);
nor U16600 (N_16600,N_16087,N_16044);
nand U16601 (N_16601,N_16016,N_16450);
nor U16602 (N_16602,N_16057,N_16146);
nand U16603 (N_16603,N_16452,N_16047);
nand U16604 (N_16604,N_16498,N_16107);
xnor U16605 (N_16605,N_16340,N_16130);
xnor U16606 (N_16606,N_16290,N_16334);
xor U16607 (N_16607,N_16365,N_16172);
or U16608 (N_16608,N_16082,N_16397);
and U16609 (N_16609,N_16201,N_16425);
xor U16610 (N_16610,N_16166,N_16011);
nand U16611 (N_16611,N_16149,N_16428);
and U16612 (N_16612,N_16045,N_16171);
or U16613 (N_16613,N_16469,N_16141);
nor U16614 (N_16614,N_16424,N_16218);
or U16615 (N_16615,N_16019,N_16257);
and U16616 (N_16616,N_16279,N_16038);
or U16617 (N_16617,N_16144,N_16052);
xor U16618 (N_16618,N_16335,N_16373);
or U16619 (N_16619,N_16269,N_16280);
xor U16620 (N_16620,N_16281,N_16020);
nand U16621 (N_16621,N_16263,N_16180);
or U16622 (N_16622,N_16256,N_16345);
or U16623 (N_16623,N_16101,N_16362);
and U16624 (N_16624,N_16155,N_16115);
xnor U16625 (N_16625,N_16075,N_16454);
or U16626 (N_16626,N_16058,N_16300);
and U16627 (N_16627,N_16461,N_16185);
nor U16628 (N_16628,N_16116,N_16306);
xor U16629 (N_16629,N_16036,N_16065);
nor U16630 (N_16630,N_16006,N_16147);
nor U16631 (N_16631,N_16189,N_16043);
xnor U16632 (N_16632,N_16278,N_16322);
or U16633 (N_16633,N_16109,N_16295);
xnor U16634 (N_16634,N_16129,N_16039);
and U16635 (N_16635,N_16320,N_16276);
nor U16636 (N_16636,N_16105,N_16010);
nand U16637 (N_16637,N_16108,N_16275);
nand U16638 (N_16638,N_16265,N_16421);
or U16639 (N_16639,N_16268,N_16244);
nor U16640 (N_16640,N_16098,N_16131);
nor U16641 (N_16641,N_16318,N_16195);
or U16642 (N_16642,N_16386,N_16206);
or U16643 (N_16643,N_16462,N_16440);
xnor U16644 (N_16644,N_16308,N_16420);
nor U16645 (N_16645,N_16134,N_16143);
and U16646 (N_16646,N_16220,N_16025);
nand U16647 (N_16647,N_16363,N_16233);
nor U16648 (N_16648,N_16194,N_16095);
and U16649 (N_16649,N_16053,N_16014);
or U16650 (N_16650,N_16102,N_16325);
nand U16651 (N_16651,N_16436,N_16135);
xor U16652 (N_16652,N_16463,N_16468);
nor U16653 (N_16653,N_16493,N_16219);
or U16654 (N_16654,N_16196,N_16222);
or U16655 (N_16655,N_16385,N_16282);
xor U16656 (N_16656,N_16297,N_16005);
xor U16657 (N_16657,N_16054,N_16394);
nand U16658 (N_16658,N_16138,N_16001);
nand U16659 (N_16659,N_16467,N_16241);
nor U16660 (N_16660,N_16332,N_16148);
and U16661 (N_16661,N_16331,N_16049);
nand U16662 (N_16662,N_16361,N_16179);
xnor U16663 (N_16663,N_16153,N_16111);
or U16664 (N_16664,N_16356,N_16458);
or U16665 (N_16665,N_16188,N_16249);
or U16666 (N_16666,N_16199,N_16250);
nor U16667 (N_16667,N_16475,N_16354);
xnor U16668 (N_16668,N_16348,N_16000);
nand U16669 (N_16669,N_16396,N_16301);
and U16670 (N_16670,N_16449,N_16099);
nor U16671 (N_16671,N_16432,N_16200);
or U16672 (N_16672,N_16238,N_16481);
nand U16673 (N_16673,N_16137,N_16229);
or U16674 (N_16674,N_16021,N_16266);
or U16675 (N_16675,N_16267,N_16296);
nor U16676 (N_16676,N_16485,N_16453);
or U16677 (N_16677,N_16403,N_16409);
xor U16678 (N_16678,N_16350,N_16142);
nand U16679 (N_16679,N_16228,N_16203);
or U16680 (N_16680,N_16217,N_16487);
nand U16681 (N_16681,N_16003,N_16216);
and U16682 (N_16682,N_16106,N_16442);
or U16683 (N_16683,N_16157,N_16151);
or U16684 (N_16684,N_16313,N_16139);
nor U16685 (N_16685,N_16382,N_16041);
and U16686 (N_16686,N_16270,N_16167);
nor U16687 (N_16687,N_16235,N_16214);
nor U16688 (N_16688,N_16071,N_16223);
xnor U16689 (N_16689,N_16376,N_16401);
and U16690 (N_16690,N_16457,N_16029);
or U16691 (N_16691,N_16104,N_16026);
and U16692 (N_16692,N_16299,N_16161);
and U16693 (N_16693,N_16411,N_16402);
xnor U16694 (N_16694,N_16404,N_16321);
and U16695 (N_16695,N_16193,N_16393);
nor U16696 (N_16696,N_16431,N_16240);
nor U16697 (N_16697,N_16474,N_16447);
nor U16698 (N_16698,N_16360,N_16035);
or U16699 (N_16699,N_16388,N_16210);
nand U16700 (N_16700,N_16379,N_16464);
nand U16701 (N_16701,N_16086,N_16069);
nor U16702 (N_16702,N_16080,N_16310);
and U16703 (N_16703,N_16405,N_16456);
nand U16704 (N_16704,N_16495,N_16187);
and U16705 (N_16705,N_16164,N_16034);
xnor U16706 (N_16706,N_16046,N_16351);
nor U16707 (N_16707,N_16245,N_16152);
or U16708 (N_16708,N_16162,N_16112);
nand U16709 (N_16709,N_16110,N_16344);
and U16710 (N_16710,N_16177,N_16326);
nor U16711 (N_16711,N_16173,N_16494);
nand U16712 (N_16712,N_16327,N_16294);
xnor U16713 (N_16713,N_16083,N_16198);
xnor U16714 (N_16714,N_16262,N_16377);
nor U16715 (N_16715,N_16287,N_16247);
nor U16716 (N_16716,N_16114,N_16391);
nor U16717 (N_16717,N_16056,N_16314);
xor U16718 (N_16718,N_16483,N_16077);
nor U16719 (N_16719,N_16400,N_16389);
and U16720 (N_16720,N_16353,N_16165);
or U16721 (N_16721,N_16378,N_16190);
or U16722 (N_16722,N_16027,N_16370);
nor U16723 (N_16723,N_16066,N_16292);
nand U16724 (N_16724,N_16122,N_16419);
xnor U16725 (N_16725,N_16048,N_16258);
nand U16726 (N_16726,N_16478,N_16261);
nor U16727 (N_16727,N_16073,N_16237);
and U16728 (N_16728,N_16303,N_16422);
or U16729 (N_16729,N_16076,N_16383);
and U16730 (N_16730,N_16236,N_16477);
nand U16731 (N_16731,N_16128,N_16260);
xor U16732 (N_16732,N_16174,N_16410);
nand U16733 (N_16733,N_16175,N_16336);
or U16734 (N_16734,N_16284,N_16375);
nand U16735 (N_16735,N_16369,N_16123);
nor U16736 (N_16736,N_16156,N_16170);
and U16737 (N_16737,N_16307,N_16479);
or U16738 (N_16738,N_16120,N_16302);
xnor U16739 (N_16739,N_16489,N_16492);
and U16740 (N_16740,N_16031,N_16068);
xor U16741 (N_16741,N_16429,N_16459);
or U16742 (N_16742,N_16018,N_16028);
nand U16743 (N_16743,N_16204,N_16359);
nand U16744 (N_16744,N_16009,N_16298);
nor U16745 (N_16745,N_16285,N_16050);
xor U16746 (N_16746,N_16024,N_16305);
xnor U16747 (N_16747,N_16316,N_16119);
nor U16748 (N_16748,N_16311,N_16090);
xnor U16749 (N_16749,N_16060,N_16323);
and U16750 (N_16750,N_16051,N_16038);
nor U16751 (N_16751,N_16063,N_16350);
and U16752 (N_16752,N_16218,N_16250);
xor U16753 (N_16753,N_16468,N_16085);
nand U16754 (N_16754,N_16477,N_16325);
nor U16755 (N_16755,N_16143,N_16243);
nor U16756 (N_16756,N_16432,N_16007);
or U16757 (N_16757,N_16194,N_16125);
and U16758 (N_16758,N_16141,N_16297);
and U16759 (N_16759,N_16161,N_16224);
nor U16760 (N_16760,N_16391,N_16155);
nor U16761 (N_16761,N_16388,N_16435);
nor U16762 (N_16762,N_16181,N_16271);
nor U16763 (N_16763,N_16093,N_16186);
xor U16764 (N_16764,N_16174,N_16206);
nor U16765 (N_16765,N_16438,N_16084);
or U16766 (N_16766,N_16292,N_16145);
xnor U16767 (N_16767,N_16347,N_16015);
and U16768 (N_16768,N_16172,N_16346);
xnor U16769 (N_16769,N_16075,N_16279);
nand U16770 (N_16770,N_16284,N_16436);
nand U16771 (N_16771,N_16455,N_16058);
nand U16772 (N_16772,N_16391,N_16373);
nor U16773 (N_16773,N_16133,N_16039);
and U16774 (N_16774,N_16215,N_16458);
nand U16775 (N_16775,N_16041,N_16286);
nand U16776 (N_16776,N_16093,N_16031);
nand U16777 (N_16777,N_16314,N_16273);
nand U16778 (N_16778,N_16260,N_16063);
nor U16779 (N_16779,N_16054,N_16108);
xnor U16780 (N_16780,N_16144,N_16007);
and U16781 (N_16781,N_16165,N_16448);
nor U16782 (N_16782,N_16427,N_16270);
nor U16783 (N_16783,N_16059,N_16197);
nand U16784 (N_16784,N_16009,N_16112);
and U16785 (N_16785,N_16010,N_16147);
xor U16786 (N_16786,N_16022,N_16226);
nor U16787 (N_16787,N_16278,N_16155);
and U16788 (N_16788,N_16153,N_16056);
nor U16789 (N_16789,N_16206,N_16299);
xnor U16790 (N_16790,N_16261,N_16134);
or U16791 (N_16791,N_16046,N_16251);
xnor U16792 (N_16792,N_16028,N_16436);
nor U16793 (N_16793,N_16156,N_16446);
nor U16794 (N_16794,N_16073,N_16169);
nand U16795 (N_16795,N_16347,N_16306);
nor U16796 (N_16796,N_16265,N_16049);
nor U16797 (N_16797,N_16235,N_16176);
xor U16798 (N_16798,N_16428,N_16075);
nand U16799 (N_16799,N_16176,N_16036);
xor U16800 (N_16800,N_16108,N_16291);
nor U16801 (N_16801,N_16185,N_16430);
and U16802 (N_16802,N_16181,N_16203);
nand U16803 (N_16803,N_16363,N_16456);
nor U16804 (N_16804,N_16178,N_16344);
or U16805 (N_16805,N_16412,N_16258);
and U16806 (N_16806,N_16085,N_16044);
nand U16807 (N_16807,N_16069,N_16224);
or U16808 (N_16808,N_16163,N_16289);
and U16809 (N_16809,N_16285,N_16270);
and U16810 (N_16810,N_16275,N_16382);
or U16811 (N_16811,N_16171,N_16161);
xor U16812 (N_16812,N_16004,N_16399);
or U16813 (N_16813,N_16481,N_16299);
nand U16814 (N_16814,N_16290,N_16207);
xor U16815 (N_16815,N_16323,N_16025);
or U16816 (N_16816,N_16336,N_16017);
nand U16817 (N_16817,N_16063,N_16324);
nand U16818 (N_16818,N_16415,N_16333);
or U16819 (N_16819,N_16032,N_16148);
or U16820 (N_16820,N_16132,N_16308);
nand U16821 (N_16821,N_16207,N_16236);
nand U16822 (N_16822,N_16299,N_16162);
xor U16823 (N_16823,N_16077,N_16472);
xor U16824 (N_16824,N_16046,N_16050);
nand U16825 (N_16825,N_16380,N_16227);
and U16826 (N_16826,N_16010,N_16412);
xor U16827 (N_16827,N_16085,N_16003);
and U16828 (N_16828,N_16213,N_16272);
or U16829 (N_16829,N_16258,N_16010);
or U16830 (N_16830,N_16222,N_16236);
xor U16831 (N_16831,N_16278,N_16454);
nor U16832 (N_16832,N_16259,N_16408);
or U16833 (N_16833,N_16066,N_16455);
nor U16834 (N_16834,N_16220,N_16186);
xor U16835 (N_16835,N_16263,N_16330);
and U16836 (N_16836,N_16155,N_16190);
and U16837 (N_16837,N_16469,N_16135);
nand U16838 (N_16838,N_16300,N_16104);
and U16839 (N_16839,N_16478,N_16443);
nor U16840 (N_16840,N_16080,N_16042);
nor U16841 (N_16841,N_16307,N_16350);
nor U16842 (N_16842,N_16089,N_16173);
and U16843 (N_16843,N_16485,N_16152);
nor U16844 (N_16844,N_16381,N_16097);
and U16845 (N_16845,N_16468,N_16441);
or U16846 (N_16846,N_16176,N_16049);
nor U16847 (N_16847,N_16110,N_16145);
xnor U16848 (N_16848,N_16352,N_16027);
nand U16849 (N_16849,N_16349,N_16446);
nand U16850 (N_16850,N_16432,N_16418);
nor U16851 (N_16851,N_16255,N_16496);
nand U16852 (N_16852,N_16207,N_16320);
and U16853 (N_16853,N_16369,N_16094);
or U16854 (N_16854,N_16436,N_16152);
or U16855 (N_16855,N_16447,N_16402);
or U16856 (N_16856,N_16331,N_16447);
nand U16857 (N_16857,N_16400,N_16008);
or U16858 (N_16858,N_16321,N_16061);
nand U16859 (N_16859,N_16275,N_16454);
nor U16860 (N_16860,N_16274,N_16473);
and U16861 (N_16861,N_16315,N_16171);
xor U16862 (N_16862,N_16016,N_16307);
nand U16863 (N_16863,N_16384,N_16262);
and U16864 (N_16864,N_16264,N_16355);
xor U16865 (N_16865,N_16235,N_16132);
xnor U16866 (N_16866,N_16119,N_16366);
nor U16867 (N_16867,N_16111,N_16097);
and U16868 (N_16868,N_16048,N_16298);
xnor U16869 (N_16869,N_16395,N_16032);
xnor U16870 (N_16870,N_16432,N_16229);
xnor U16871 (N_16871,N_16341,N_16006);
and U16872 (N_16872,N_16058,N_16161);
and U16873 (N_16873,N_16324,N_16473);
and U16874 (N_16874,N_16355,N_16122);
nand U16875 (N_16875,N_16250,N_16213);
nand U16876 (N_16876,N_16008,N_16399);
and U16877 (N_16877,N_16112,N_16492);
or U16878 (N_16878,N_16403,N_16014);
nand U16879 (N_16879,N_16042,N_16254);
and U16880 (N_16880,N_16049,N_16249);
and U16881 (N_16881,N_16181,N_16034);
nand U16882 (N_16882,N_16119,N_16486);
nor U16883 (N_16883,N_16406,N_16042);
or U16884 (N_16884,N_16318,N_16016);
and U16885 (N_16885,N_16449,N_16126);
or U16886 (N_16886,N_16496,N_16076);
nand U16887 (N_16887,N_16005,N_16372);
nor U16888 (N_16888,N_16499,N_16391);
and U16889 (N_16889,N_16186,N_16022);
nand U16890 (N_16890,N_16140,N_16038);
xnor U16891 (N_16891,N_16061,N_16396);
and U16892 (N_16892,N_16448,N_16091);
nand U16893 (N_16893,N_16080,N_16108);
nand U16894 (N_16894,N_16431,N_16229);
nand U16895 (N_16895,N_16427,N_16216);
xor U16896 (N_16896,N_16197,N_16367);
or U16897 (N_16897,N_16058,N_16434);
or U16898 (N_16898,N_16029,N_16044);
nor U16899 (N_16899,N_16343,N_16454);
or U16900 (N_16900,N_16376,N_16049);
and U16901 (N_16901,N_16083,N_16464);
nand U16902 (N_16902,N_16360,N_16395);
and U16903 (N_16903,N_16175,N_16033);
nor U16904 (N_16904,N_16403,N_16109);
or U16905 (N_16905,N_16377,N_16269);
nand U16906 (N_16906,N_16129,N_16289);
and U16907 (N_16907,N_16039,N_16041);
nand U16908 (N_16908,N_16240,N_16356);
and U16909 (N_16909,N_16445,N_16117);
or U16910 (N_16910,N_16000,N_16370);
xnor U16911 (N_16911,N_16175,N_16319);
nand U16912 (N_16912,N_16216,N_16195);
xnor U16913 (N_16913,N_16246,N_16347);
nor U16914 (N_16914,N_16486,N_16180);
and U16915 (N_16915,N_16072,N_16176);
and U16916 (N_16916,N_16342,N_16387);
nor U16917 (N_16917,N_16368,N_16497);
or U16918 (N_16918,N_16361,N_16196);
nor U16919 (N_16919,N_16443,N_16268);
xor U16920 (N_16920,N_16029,N_16302);
nor U16921 (N_16921,N_16264,N_16349);
xnor U16922 (N_16922,N_16058,N_16314);
or U16923 (N_16923,N_16125,N_16409);
nand U16924 (N_16924,N_16305,N_16434);
and U16925 (N_16925,N_16488,N_16066);
or U16926 (N_16926,N_16032,N_16017);
or U16927 (N_16927,N_16281,N_16143);
or U16928 (N_16928,N_16459,N_16183);
or U16929 (N_16929,N_16458,N_16034);
or U16930 (N_16930,N_16061,N_16397);
nor U16931 (N_16931,N_16300,N_16234);
and U16932 (N_16932,N_16304,N_16134);
xor U16933 (N_16933,N_16067,N_16145);
or U16934 (N_16934,N_16043,N_16356);
nand U16935 (N_16935,N_16126,N_16257);
or U16936 (N_16936,N_16277,N_16322);
nand U16937 (N_16937,N_16083,N_16096);
nor U16938 (N_16938,N_16250,N_16306);
nand U16939 (N_16939,N_16344,N_16184);
and U16940 (N_16940,N_16463,N_16466);
nand U16941 (N_16941,N_16435,N_16099);
and U16942 (N_16942,N_16399,N_16323);
nor U16943 (N_16943,N_16160,N_16017);
nand U16944 (N_16944,N_16016,N_16259);
xor U16945 (N_16945,N_16337,N_16112);
nand U16946 (N_16946,N_16137,N_16046);
nand U16947 (N_16947,N_16348,N_16245);
nand U16948 (N_16948,N_16475,N_16207);
xnor U16949 (N_16949,N_16033,N_16187);
and U16950 (N_16950,N_16301,N_16385);
or U16951 (N_16951,N_16008,N_16499);
and U16952 (N_16952,N_16364,N_16199);
nor U16953 (N_16953,N_16460,N_16150);
nor U16954 (N_16954,N_16170,N_16412);
nand U16955 (N_16955,N_16489,N_16412);
and U16956 (N_16956,N_16034,N_16409);
xor U16957 (N_16957,N_16301,N_16202);
nand U16958 (N_16958,N_16122,N_16322);
nand U16959 (N_16959,N_16406,N_16016);
xnor U16960 (N_16960,N_16104,N_16194);
and U16961 (N_16961,N_16163,N_16151);
nand U16962 (N_16962,N_16199,N_16347);
xor U16963 (N_16963,N_16188,N_16417);
or U16964 (N_16964,N_16318,N_16284);
xor U16965 (N_16965,N_16045,N_16281);
xnor U16966 (N_16966,N_16136,N_16197);
or U16967 (N_16967,N_16200,N_16346);
nor U16968 (N_16968,N_16029,N_16338);
nand U16969 (N_16969,N_16001,N_16151);
nor U16970 (N_16970,N_16098,N_16373);
nor U16971 (N_16971,N_16170,N_16048);
nor U16972 (N_16972,N_16138,N_16274);
or U16973 (N_16973,N_16096,N_16232);
nand U16974 (N_16974,N_16335,N_16321);
and U16975 (N_16975,N_16178,N_16422);
xor U16976 (N_16976,N_16404,N_16248);
nor U16977 (N_16977,N_16327,N_16093);
and U16978 (N_16978,N_16141,N_16274);
and U16979 (N_16979,N_16046,N_16412);
and U16980 (N_16980,N_16302,N_16177);
nand U16981 (N_16981,N_16404,N_16018);
and U16982 (N_16982,N_16480,N_16327);
or U16983 (N_16983,N_16437,N_16155);
nor U16984 (N_16984,N_16256,N_16469);
or U16985 (N_16985,N_16399,N_16403);
nand U16986 (N_16986,N_16295,N_16482);
xnor U16987 (N_16987,N_16400,N_16334);
or U16988 (N_16988,N_16142,N_16330);
nor U16989 (N_16989,N_16207,N_16218);
and U16990 (N_16990,N_16102,N_16055);
nand U16991 (N_16991,N_16290,N_16462);
xor U16992 (N_16992,N_16335,N_16085);
nor U16993 (N_16993,N_16185,N_16161);
xnor U16994 (N_16994,N_16327,N_16103);
or U16995 (N_16995,N_16303,N_16454);
xor U16996 (N_16996,N_16192,N_16072);
and U16997 (N_16997,N_16031,N_16371);
and U16998 (N_16998,N_16028,N_16405);
xor U16999 (N_16999,N_16441,N_16436);
or U17000 (N_17000,N_16545,N_16563);
xor U17001 (N_17001,N_16999,N_16668);
and U17002 (N_17002,N_16865,N_16663);
and U17003 (N_17003,N_16530,N_16814);
nand U17004 (N_17004,N_16797,N_16576);
nand U17005 (N_17005,N_16812,N_16929);
and U17006 (N_17006,N_16989,N_16821);
xor U17007 (N_17007,N_16686,N_16775);
or U17008 (N_17008,N_16689,N_16727);
and U17009 (N_17009,N_16592,N_16777);
or U17010 (N_17010,N_16705,N_16778);
or U17011 (N_17011,N_16849,N_16992);
and U17012 (N_17012,N_16868,N_16895);
nand U17013 (N_17013,N_16936,N_16752);
or U17014 (N_17014,N_16572,N_16794);
and U17015 (N_17015,N_16561,N_16824);
or U17016 (N_17016,N_16851,N_16957);
nor U17017 (N_17017,N_16925,N_16627);
nand U17018 (N_17018,N_16903,N_16951);
xor U17019 (N_17019,N_16599,N_16772);
xor U17020 (N_17020,N_16913,N_16610);
xor U17021 (N_17021,N_16863,N_16784);
or U17022 (N_17022,N_16507,N_16609);
and U17023 (N_17023,N_16860,N_16670);
nand U17024 (N_17024,N_16833,N_16575);
or U17025 (N_17025,N_16871,N_16807);
xor U17026 (N_17026,N_16745,N_16783);
and U17027 (N_17027,N_16964,N_16955);
nand U17028 (N_17028,N_16677,N_16901);
or U17029 (N_17029,N_16854,N_16780);
or U17030 (N_17030,N_16861,N_16946);
and U17031 (N_17031,N_16688,N_16822);
nor U17032 (N_17032,N_16562,N_16881);
nor U17033 (N_17033,N_16630,N_16574);
or U17034 (N_17034,N_16698,N_16602);
or U17035 (N_17035,N_16622,N_16603);
and U17036 (N_17036,N_16595,N_16831);
nor U17037 (N_17037,N_16921,N_16549);
xnor U17038 (N_17038,N_16884,N_16914);
or U17039 (N_17039,N_16623,N_16830);
and U17040 (N_17040,N_16737,N_16912);
xor U17041 (N_17041,N_16648,N_16748);
and U17042 (N_17042,N_16606,N_16584);
xor U17043 (N_17043,N_16766,N_16840);
or U17044 (N_17044,N_16819,N_16781);
and U17045 (N_17045,N_16974,N_16856);
and U17046 (N_17046,N_16687,N_16624);
or U17047 (N_17047,N_16501,N_16759);
nand U17048 (N_17048,N_16607,N_16618);
nor U17049 (N_17049,N_16621,N_16629);
nor U17050 (N_17050,N_16892,N_16692);
nand U17051 (N_17051,N_16911,N_16719);
nand U17052 (N_17052,N_16720,N_16960);
nor U17053 (N_17053,N_16845,N_16755);
and U17054 (N_17054,N_16581,N_16976);
and U17055 (N_17055,N_16568,N_16557);
or U17056 (N_17056,N_16724,N_16899);
and U17057 (N_17057,N_16524,N_16855);
nor U17058 (N_17058,N_16632,N_16799);
or U17059 (N_17059,N_16548,N_16986);
nand U17060 (N_17060,N_16517,N_16848);
nor U17061 (N_17061,N_16559,N_16950);
or U17062 (N_17062,N_16877,N_16674);
nor U17063 (N_17063,N_16656,N_16972);
xnor U17064 (N_17064,N_16835,N_16917);
or U17065 (N_17065,N_16829,N_16940);
xnor U17066 (N_17066,N_16850,N_16998);
or U17067 (N_17067,N_16716,N_16876);
xor U17068 (N_17068,N_16558,N_16743);
xnor U17069 (N_17069,N_16928,N_16800);
and U17070 (N_17070,N_16585,N_16506);
nand U17071 (N_17071,N_16813,N_16547);
nand U17072 (N_17072,N_16653,N_16802);
xor U17073 (N_17073,N_16565,N_16742);
or U17074 (N_17074,N_16587,N_16675);
nand U17075 (N_17075,N_16991,N_16634);
and U17076 (N_17076,N_16915,N_16662);
nor U17077 (N_17077,N_16704,N_16982);
xnor U17078 (N_17078,N_16652,N_16730);
xnor U17079 (N_17079,N_16593,N_16505);
nand U17080 (N_17080,N_16612,N_16765);
xor U17081 (N_17081,N_16700,N_16941);
nand U17082 (N_17082,N_16669,N_16939);
and U17083 (N_17083,N_16509,N_16699);
or U17084 (N_17084,N_16681,N_16514);
xnor U17085 (N_17085,N_16885,N_16927);
or U17086 (N_17086,N_16853,N_16810);
nand U17087 (N_17087,N_16805,N_16697);
xnor U17088 (N_17088,N_16749,N_16611);
nor U17089 (N_17089,N_16943,N_16747);
xor U17090 (N_17090,N_16694,N_16589);
xnor U17091 (N_17091,N_16735,N_16938);
or U17092 (N_17092,N_16537,N_16968);
nor U17093 (N_17093,N_16942,N_16932);
nand U17094 (N_17094,N_16862,N_16768);
and U17095 (N_17095,N_16842,N_16650);
or U17096 (N_17096,N_16949,N_16740);
and U17097 (N_17097,N_16937,N_16930);
or U17098 (N_17098,N_16706,N_16870);
nor U17099 (N_17099,N_16882,N_16788);
and U17100 (N_17100,N_16875,N_16619);
nor U17101 (N_17101,N_16963,N_16613);
nand U17102 (N_17102,N_16750,N_16625);
or U17103 (N_17103,N_16654,N_16732);
xnor U17104 (N_17104,N_16776,N_16808);
xnor U17105 (N_17105,N_16931,N_16744);
or U17106 (N_17106,N_16616,N_16715);
nand U17107 (N_17107,N_16515,N_16531);
and U17108 (N_17108,N_16746,N_16785);
xnor U17109 (N_17109,N_16679,N_16832);
and U17110 (N_17110,N_16544,N_16628);
xnor U17111 (N_17111,N_16534,N_16907);
or U17112 (N_17112,N_16731,N_16703);
nor U17113 (N_17113,N_16651,N_16555);
and U17114 (N_17114,N_16637,N_16773);
nand U17115 (N_17115,N_16990,N_16710);
xor U17116 (N_17116,N_16601,N_16714);
xnor U17117 (N_17117,N_16702,N_16567);
xnor U17118 (N_17118,N_16886,N_16543);
nor U17119 (N_17119,N_16933,N_16894);
and U17120 (N_17120,N_16512,N_16525);
and U17121 (N_17121,N_16864,N_16887);
nand U17122 (N_17122,N_16597,N_16987);
xnor U17123 (N_17123,N_16569,N_16527);
or U17124 (N_17124,N_16631,N_16945);
and U17125 (N_17125,N_16753,N_16958);
or U17126 (N_17126,N_16965,N_16836);
and U17127 (N_17127,N_16995,N_16539);
or U17128 (N_17128,N_16564,N_16893);
nand U17129 (N_17129,N_16996,N_16659);
nor U17130 (N_17130,N_16985,N_16980);
or U17131 (N_17131,N_16858,N_16983);
nor U17132 (N_17132,N_16869,N_16770);
nor U17133 (N_17133,N_16617,N_16902);
or U17134 (N_17134,N_16580,N_16641);
nand U17135 (N_17135,N_16672,N_16666);
nor U17136 (N_17136,N_16859,N_16510);
and U17137 (N_17137,N_16908,N_16728);
and U17138 (N_17138,N_16852,N_16791);
or U17139 (N_17139,N_16709,N_16536);
and U17140 (N_17140,N_16970,N_16708);
and U17141 (N_17141,N_16934,N_16997);
and U17142 (N_17142,N_16923,N_16690);
nand U17143 (N_17143,N_16684,N_16586);
nor U17144 (N_17144,N_16582,N_16532);
and U17145 (N_17145,N_16910,N_16533);
nor U17146 (N_17146,N_16846,N_16919);
or U17147 (N_17147,N_16896,N_16973);
and U17148 (N_17148,N_16635,N_16571);
and U17149 (N_17149,N_16947,N_16646);
and U17150 (N_17150,N_16661,N_16952);
xor U17151 (N_17151,N_16712,N_16795);
nand U17152 (N_17152,N_16838,N_16793);
xor U17153 (N_17153,N_16954,N_16796);
nor U17154 (N_17154,N_16693,N_16801);
nand U17155 (N_17155,N_16657,N_16874);
and U17156 (N_17156,N_16721,N_16751);
or U17157 (N_17157,N_16890,N_16502);
nor U17158 (N_17158,N_16639,N_16935);
nor U17159 (N_17159,N_16655,N_16615);
and U17160 (N_17160,N_16888,N_16682);
nor U17161 (N_17161,N_16516,N_16695);
or U17162 (N_17162,N_16552,N_16643);
nand U17163 (N_17163,N_16803,N_16590);
nand U17164 (N_17164,N_16790,N_16546);
xor U17165 (N_17165,N_16556,N_16879);
or U17166 (N_17166,N_16570,N_16872);
and U17167 (N_17167,N_16979,N_16667);
or U17168 (N_17168,N_16658,N_16847);
or U17169 (N_17169,N_16678,N_16878);
xor U17170 (N_17170,N_16522,N_16718);
nor U17171 (N_17171,N_16726,N_16873);
xor U17172 (N_17172,N_16905,N_16891);
nand U17173 (N_17173,N_16889,N_16900);
nand U17174 (N_17174,N_16528,N_16771);
xor U17175 (N_17175,N_16503,N_16540);
or U17176 (N_17176,N_16526,N_16897);
xnor U17177 (N_17177,N_16825,N_16823);
nand U17178 (N_17178,N_16676,N_16722);
and U17179 (N_17179,N_16511,N_16811);
nand U17180 (N_17180,N_16673,N_16787);
nor U17181 (N_17181,N_16588,N_16566);
nor U17182 (N_17182,N_16542,N_16577);
or U17183 (N_17183,N_16782,N_16649);
and U17184 (N_17184,N_16520,N_16600);
nor U17185 (N_17185,N_16620,N_16762);
xor U17186 (N_17186,N_16857,N_16806);
and U17187 (N_17187,N_16789,N_16591);
xnor U17188 (N_17188,N_16701,N_16798);
or U17189 (N_17189,N_16519,N_16984);
nand U17190 (N_17190,N_16761,N_16645);
nand U17191 (N_17191,N_16920,N_16521);
nand U17192 (N_17192,N_16779,N_16551);
xnor U17193 (N_17193,N_16841,N_16604);
and U17194 (N_17194,N_16553,N_16969);
nor U17195 (N_17195,N_16596,N_16725);
xnor U17196 (N_17196,N_16826,N_16614);
or U17197 (N_17197,N_16696,N_16792);
and U17198 (N_17198,N_16707,N_16786);
and U17199 (N_17199,N_16504,N_16729);
and U17200 (N_17200,N_16763,N_16717);
nand U17201 (N_17201,N_16583,N_16844);
xor U17202 (N_17202,N_16926,N_16839);
nor U17203 (N_17203,N_16754,N_16994);
xnor U17204 (N_17204,N_16904,N_16535);
and U17205 (N_17205,N_16883,N_16898);
nand U17206 (N_17206,N_16636,N_16817);
and U17207 (N_17207,N_16598,N_16962);
nor U17208 (N_17208,N_16541,N_16500);
nand U17209 (N_17209,N_16993,N_16594);
nand U17210 (N_17210,N_16804,N_16713);
xnor U17211 (N_17211,N_16736,N_16820);
or U17212 (N_17212,N_16948,N_16977);
nor U17213 (N_17213,N_16711,N_16605);
or U17214 (N_17214,N_16944,N_16733);
nand U17215 (N_17215,N_16834,N_16866);
xor U17216 (N_17216,N_16922,N_16573);
xnor U17217 (N_17217,N_16756,N_16918);
nand U17218 (N_17218,N_16809,N_16971);
xnor U17219 (N_17219,N_16880,N_16665);
nand U17220 (N_17220,N_16578,N_16579);
and U17221 (N_17221,N_16513,N_16757);
nand U17222 (N_17222,N_16739,N_16815);
nand U17223 (N_17223,N_16767,N_16671);
nand U17224 (N_17224,N_16550,N_16818);
or U17225 (N_17225,N_16978,N_16738);
or U17226 (N_17226,N_16538,N_16774);
or U17227 (N_17227,N_16981,N_16633);
nand U17228 (N_17228,N_16924,N_16685);
or U17229 (N_17229,N_16741,N_16660);
or U17230 (N_17230,N_16837,N_16764);
nand U17231 (N_17231,N_16640,N_16906);
or U17232 (N_17232,N_16966,N_16638);
nor U17233 (N_17233,N_16975,N_16647);
nand U17234 (N_17234,N_16827,N_16529);
and U17235 (N_17235,N_16691,N_16518);
xor U17236 (N_17236,N_16816,N_16664);
or U17237 (N_17237,N_16608,N_16644);
nor U17238 (N_17238,N_16828,N_16967);
and U17239 (N_17239,N_16916,N_16680);
nor U17240 (N_17240,N_16988,N_16867);
nor U17241 (N_17241,N_16734,N_16843);
and U17242 (N_17242,N_16554,N_16683);
xor U17243 (N_17243,N_16956,N_16769);
or U17244 (N_17244,N_16909,N_16523);
xor U17245 (N_17245,N_16760,N_16953);
and U17246 (N_17246,N_16959,N_16961);
or U17247 (N_17247,N_16626,N_16560);
or U17248 (N_17248,N_16508,N_16723);
or U17249 (N_17249,N_16642,N_16758);
nand U17250 (N_17250,N_16763,N_16723);
xnor U17251 (N_17251,N_16515,N_16751);
xnor U17252 (N_17252,N_16843,N_16618);
nand U17253 (N_17253,N_16642,N_16995);
xnor U17254 (N_17254,N_16984,N_16747);
and U17255 (N_17255,N_16984,N_16573);
nor U17256 (N_17256,N_16715,N_16930);
xor U17257 (N_17257,N_16607,N_16790);
nand U17258 (N_17258,N_16792,N_16957);
nor U17259 (N_17259,N_16940,N_16885);
xor U17260 (N_17260,N_16607,N_16999);
and U17261 (N_17261,N_16997,N_16941);
nand U17262 (N_17262,N_16514,N_16538);
nor U17263 (N_17263,N_16920,N_16675);
and U17264 (N_17264,N_16559,N_16853);
or U17265 (N_17265,N_16785,N_16740);
xnor U17266 (N_17266,N_16659,N_16987);
xor U17267 (N_17267,N_16569,N_16859);
nor U17268 (N_17268,N_16685,N_16617);
and U17269 (N_17269,N_16849,N_16671);
and U17270 (N_17270,N_16872,N_16655);
nand U17271 (N_17271,N_16869,N_16579);
nor U17272 (N_17272,N_16664,N_16894);
and U17273 (N_17273,N_16546,N_16563);
nand U17274 (N_17274,N_16640,N_16819);
xnor U17275 (N_17275,N_16746,N_16738);
nand U17276 (N_17276,N_16709,N_16925);
nand U17277 (N_17277,N_16680,N_16837);
nor U17278 (N_17278,N_16963,N_16731);
nor U17279 (N_17279,N_16515,N_16908);
xnor U17280 (N_17280,N_16736,N_16507);
or U17281 (N_17281,N_16625,N_16965);
or U17282 (N_17282,N_16797,N_16655);
nand U17283 (N_17283,N_16960,N_16716);
nand U17284 (N_17284,N_16903,N_16670);
nand U17285 (N_17285,N_16785,N_16862);
or U17286 (N_17286,N_16857,N_16647);
and U17287 (N_17287,N_16922,N_16536);
or U17288 (N_17288,N_16683,N_16943);
nor U17289 (N_17289,N_16982,N_16798);
or U17290 (N_17290,N_16584,N_16610);
nand U17291 (N_17291,N_16626,N_16765);
and U17292 (N_17292,N_16716,N_16651);
nand U17293 (N_17293,N_16652,N_16664);
and U17294 (N_17294,N_16646,N_16752);
nor U17295 (N_17295,N_16644,N_16784);
xor U17296 (N_17296,N_16667,N_16812);
nor U17297 (N_17297,N_16536,N_16955);
or U17298 (N_17298,N_16971,N_16826);
or U17299 (N_17299,N_16842,N_16874);
nand U17300 (N_17300,N_16700,N_16922);
nor U17301 (N_17301,N_16580,N_16699);
nand U17302 (N_17302,N_16821,N_16863);
xor U17303 (N_17303,N_16789,N_16704);
nor U17304 (N_17304,N_16742,N_16772);
nand U17305 (N_17305,N_16655,N_16782);
xor U17306 (N_17306,N_16737,N_16553);
nand U17307 (N_17307,N_16569,N_16954);
nand U17308 (N_17308,N_16723,N_16889);
and U17309 (N_17309,N_16876,N_16705);
nand U17310 (N_17310,N_16838,N_16661);
xor U17311 (N_17311,N_16684,N_16715);
or U17312 (N_17312,N_16932,N_16755);
or U17313 (N_17313,N_16903,N_16500);
nor U17314 (N_17314,N_16952,N_16973);
xor U17315 (N_17315,N_16635,N_16862);
nor U17316 (N_17316,N_16959,N_16887);
nand U17317 (N_17317,N_16934,N_16793);
xnor U17318 (N_17318,N_16507,N_16953);
nor U17319 (N_17319,N_16886,N_16892);
and U17320 (N_17320,N_16960,N_16568);
nand U17321 (N_17321,N_16768,N_16974);
and U17322 (N_17322,N_16655,N_16573);
and U17323 (N_17323,N_16937,N_16808);
xnor U17324 (N_17324,N_16711,N_16588);
and U17325 (N_17325,N_16844,N_16631);
or U17326 (N_17326,N_16529,N_16931);
or U17327 (N_17327,N_16864,N_16622);
nand U17328 (N_17328,N_16953,N_16860);
and U17329 (N_17329,N_16541,N_16845);
nand U17330 (N_17330,N_16794,N_16792);
xor U17331 (N_17331,N_16776,N_16604);
and U17332 (N_17332,N_16616,N_16588);
nand U17333 (N_17333,N_16841,N_16960);
nand U17334 (N_17334,N_16637,N_16633);
nand U17335 (N_17335,N_16775,N_16991);
nand U17336 (N_17336,N_16917,N_16830);
nor U17337 (N_17337,N_16612,N_16818);
nand U17338 (N_17338,N_16944,N_16823);
nor U17339 (N_17339,N_16824,N_16647);
and U17340 (N_17340,N_16597,N_16762);
or U17341 (N_17341,N_16914,N_16644);
or U17342 (N_17342,N_16854,N_16554);
nand U17343 (N_17343,N_16799,N_16747);
and U17344 (N_17344,N_16915,N_16810);
xnor U17345 (N_17345,N_16939,N_16824);
xor U17346 (N_17346,N_16805,N_16759);
and U17347 (N_17347,N_16718,N_16874);
and U17348 (N_17348,N_16908,N_16811);
nand U17349 (N_17349,N_16796,N_16977);
and U17350 (N_17350,N_16857,N_16638);
or U17351 (N_17351,N_16629,N_16760);
or U17352 (N_17352,N_16915,N_16788);
and U17353 (N_17353,N_16704,N_16798);
xor U17354 (N_17354,N_16816,N_16708);
nand U17355 (N_17355,N_16617,N_16903);
or U17356 (N_17356,N_16987,N_16819);
or U17357 (N_17357,N_16817,N_16901);
or U17358 (N_17358,N_16682,N_16551);
xnor U17359 (N_17359,N_16528,N_16936);
nor U17360 (N_17360,N_16565,N_16535);
nand U17361 (N_17361,N_16997,N_16528);
nand U17362 (N_17362,N_16679,N_16690);
or U17363 (N_17363,N_16678,N_16750);
nor U17364 (N_17364,N_16707,N_16771);
nand U17365 (N_17365,N_16803,N_16500);
nand U17366 (N_17366,N_16828,N_16549);
xor U17367 (N_17367,N_16937,N_16910);
or U17368 (N_17368,N_16676,N_16910);
or U17369 (N_17369,N_16931,N_16851);
xnor U17370 (N_17370,N_16695,N_16757);
or U17371 (N_17371,N_16592,N_16942);
nor U17372 (N_17372,N_16596,N_16522);
nand U17373 (N_17373,N_16824,N_16747);
or U17374 (N_17374,N_16605,N_16627);
nor U17375 (N_17375,N_16849,N_16961);
and U17376 (N_17376,N_16835,N_16882);
nand U17377 (N_17377,N_16546,N_16589);
or U17378 (N_17378,N_16721,N_16714);
or U17379 (N_17379,N_16724,N_16834);
or U17380 (N_17380,N_16707,N_16559);
xor U17381 (N_17381,N_16691,N_16709);
nor U17382 (N_17382,N_16526,N_16626);
xnor U17383 (N_17383,N_16963,N_16505);
or U17384 (N_17384,N_16827,N_16855);
xnor U17385 (N_17385,N_16646,N_16778);
xor U17386 (N_17386,N_16698,N_16832);
nor U17387 (N_17387,N_16742,N_16975);
or U17388 (N_17388,N_16745,N_16503);
nand U17389 (N_17389,N_16851,N_16514);
and U17390 (N_17390,N_16628,N_16888);
nor U17391 (N_17391,N_16509,N_16826);
and U17392 (N_17392,N_16936,N_16858);
nor U17393 (N_17393,N_16591,N_16888);
nand U17394 (N_17394,N_16935,N_16803);
or U17395 (N_17395,N_16638,N_16806);
xnor U17396 (N_17396,N_16783,N_16893);
and U17397 (N_17397,N_16682,N_16726);
xnor U17398 (N_17398,N_16570,N_16839);
nand U17399 (N_17399,N_16587,N_16725);
xor U17400 (N_17400,N_16523,N_16950);
xor U17401 (N_17401,N_16540,N_16832);
nor U17402 (N_17402,N_16819,N_16592);
xor U17403 (N_17403,N_16739,N_16672);
or U17404 (N_17404,N_16503,N_16699);
xnor U17405 (N_17405,N_16801,N_16772);
and U17406 (N_17406,N_16943,N_16722);
or U17407 (N_17407,N_16563,N_16933);
xor U17408 (N_17408,N_16604,N_16728);
or U17409 (N_17409,N_16952,N_16528);
or U17410 (N_17410,N_16597,N_16924);
nor U17411 (N_17411,N_16843,N_16669);
nor U17412 (N_17412,N_16724,N_16922);
xor U17413 (N_17413,N_16974,N_16844);
or U17414 (N_17414,N_16708,N_16544);
nand U17415 (N_17415,N_16989,N_16579);
nand U17416 (N_17416,N_16966,N_16994);
nor U17417 (N_17417,N_16704,N_16837);
or U17418 (N_17418,N_16675,N_16962);
and U17419 (N_17419,N_16621,N_16940);
nand U17420 (N_17420,N_16807,N_16556);
and U17421 (N_17421,N_16517,N_16622);
nor U17422 (N_17422,N_16646,N_16545);
nor U17423 (N_17423,N_16967,N_16868);
nand U17424 (N_17424,N_16995,N_16868);
nand U17425 (N_17425,N_16662,N_16568);
or U17426 (N_17426,N_16670,N_16611);
xor U17427 (N_17427,N_16784,N_16882);
nor U17428 (N_17428,N_16966,N_16889);
and U17429 (N_17429,N_16851,N_16988);
nand U17430 (N_17430,N_16965,N_16828);
xor U17431 (N_17431,N_16977,N_16922);
nor U17432 (N_17432,N_16776,N_16893);
nand U17433 (N_17433,N_16705,N_16956);
or U17434 (N_17434,N_16747,N_16529);
xnor U17435 (N_17435,N_16573,N_16892);
nand U17436 (N_17436,N_16598,N_16549);
nor U17437 (N_17437,N_16603,N_16880);
or U17438 (N_17438,N_16682,N_16591);
xnor U17439 (N_17439,N_16511,N_16814);
xnor U17440 (N_17440,N_16567,N_16565);
and U17441 (N_17441,N_16810,N_16862);
nand U17442 (N_17442,N_16665,N_16993);
nor U17443 (N_17443,N_16974,N_16928);
and U17444 (N_17444,N_16999,N_16923);
and U17445 (N_17445,N_16952,N_16648);
nand U17446 (N_17446,N_16793,N_16731);
nand U17447 (N_17447,N_16997,N_16881);
xor U17448 (N_17448,N_16560,N_16685);
and U17449 (N_17449,N_16603,N_16592);
nor U17450 (N_17450,N_16822,N_16856);
and U17451 (N_17451,N_16570,N_16714);
nor U17452 (N_17452,N_16902,N_16985);
and U17453 (N_17453,N_16747,N_16803);
xnor U17454 (N_17454,N_16912,N_16798);
nor U17455 (N_17455,N_16890,N_16712);
nand U17456 (N_17456,N_16624,N_16642);
and U17457 (N_17457,N_16825,N_16957);
xnor U17458 (N_17458,N_16936,N_16673);
or U17459 (N_17459,N_16563,N_16847);
and U17460 (N_17460,N_16861,N_16601);
and U17461 (N_17461,N_16855,N_16974);
nand U17462 (N_17462,N_16808,N_16796);
nor U17463 (N_17463,N_16648,N_16802);
or U17464 (N_17464,N_16574,N_16538);
or U17465 (N_17465,N_16593,N_16955);
and U17466 (N_17466,N_16907,N_16774);
xor U17467 (N_17467,N_16780,N_16924);
nand U17468 (N_17468,N_16829,N_16747);
and U17469 (N_17469,N_16651,N_16661);
nor U17470 (N_17470,N_16778,N_16663);
xnor U17471 (N_17471,N_16842,N_16792);
xnor U17472 (N_17472,N_16646,N_16724);
nand U17473 (N_17473,N_16892,N_16734);
nand U17474 (N_17474,N_16817,N_16683);
or U17475 (N_17475,N_16792,N_16992);
nand U17476 (N_17476,N_16730,N_16860);
nand U17477 (N_17477,N_16530,N_16807);
nor U17478 (N_17478,N_16720,N_16870);
nand U17479 (N_17479,N_16531,N_16850);
nor U17480 (N_17480,N_16563,N_16590);
and U17481 (N_17481,N_16562,N_16972);
and U17482 (N_17482,N_16966,N_16629);
or U17483 (N_17483,N_16669,N_16876);
or U17484 (N_17484,N_16784,N_16970);
xor U17485 (N_17485,N_16739,N_16632);
and U17486 (N_17486,N_16900,N_16616);
xnor U17487 (N_17487,N_16928,N_16892);
nand U17488 (N_17488,N_16742,N_16777);
and U17489 (N_17489,N_16901,N_16531);
or U17490 (N_17490,N_16721,N_16653);
or U17491 (N_17491,N_16843,N_16866);
nor U17492 (N_17492,N_16864,N_16556);
nor U17493 (N_17493,N_16607,N_16822);
xnor U17494 (N_17494,N_16985,N_16662);
and U17495 (N_17495,N_16587,N_16538);
or U17496 (N_17496,N_16795,N_16951);
and U17497 (N_17497,N_16737,N_16622);
nand U17498 (N_17498,N_16695,N_16779);
nor U17499 (N_17499,N_16626,N_16528);
nand U17500 (N_17500,N_17293,N_17247);
or U17501 (N_17501,N_17428,N_17416);
nor U17502 (N_17502,N_17227,N_17350);
nor U17503 (N_17503,N_17048,N_17029);
nand U17504 (N_17504,N_17394,N_17474);
and U17505 (N_17505,N_17456,N_17482);
or U17506 (N_17506,N_17298,N_17067);
or U17507 (N_17507,N_17290,N_17007);
nor U17508 (N_17508,N_17437,N_17452);
and U17509 (N_17509,N_17092,N_17095);
nor U17510 (N_17510,N_17008,N_17371);
and U17511 (N_17511,N_17167,N_17120);
xnor U17512 (N_17512,N_17027,N_17179);
nor U17513 (N_17513,N_17275,N_17049);
and U17514 (N_17514,N_17238,N_17003);
xor U17515 (N_17515,N_17412,N_17181);
xnor U17516 (N_17516,N_17091,N_17036);
or U17517 (N_17517,N_17471,N_17273);
or U17518 (N_17518,N_17282,N_17462);
and U17519 (N_17519,N_17388,N_17072);
or U17520 (N_17520,N_17039,N_17415);
and U17521 (N_17521,N_17132,N_17302);
nand U17522 (N_17522,N_17458,N_17487);
nor U17523 (N_17523,N_17359,N_17442);
nand U17524 (N_17524,N_17361,N_17090);
nor U17525 (N_17525,N_17080,N_17041);
and U17526 (N_17526,N_17206,N_17110);
or U17527 (N_17527,N_17079,N_17358);
nor U17528 (N_17528,N_17499,N_17387);
xor U17529 (N_17529,N_17297,N_17497);
or U17530 (N_17530,N_17009,N_17168);
xnor U17531 (N_17531,N_17362,N_17022);
and U17532 (N_17532,N_17266,N_17339);
and U17533 (N_17533,N_17429,N_17054);
nand U17534 (N_17534,N_17197,N_17444);
nor U17535 (N_17535,N_17112,N_17470);
or U17536 (N_17536,N_17130,N_17246);
or U17537 (N_17537,N_17294,N_17484);
or U17538 (N_17538,N_17017,N_17129);
nand U17539 (N_17539,N_17045,N_17177);
nor U17540 (N_17540,N_17402,N_17226);
and U17541 (N_17541,N_17146,N_17315);
and U17542 (N_17542,N_17433,N_17403);
and U17543 (N_17543,N_17195,N_17065);
nand U17544 (N_17544,N_17320,N_17400);
and U17545 (N_17545,N_17194,N_17097);
nor U17546 (N_17546,N_17062,N_17351);
and U17547 (N_17547,N_17133,N_17220);
nand U17548 (N_17548,N_17427,N_17231);
nand U17549 (N_17549,N_17114,N_17207);
xnor U17550 (N_17550,N_17439,N_17322);
nand U17551 (N_17551,N_17372,N_17461);
nor U17552 (N_17552,N_17391,N_17038);
nand U17553 (N_17553,N_17406,N_17089);
or U17554 (N_17554,N_17104,N_17043);
or U17555 (N_17555,N_17098,N_17085);
and U17556 (N_17556,N_17056,N_17453);
and U17557 (N_17557,N_17139,N_17047);
and U17558 (N_17558,N_17086,N_17128);
nor U17559 (N_17559,N_17399,N_17284);
and U17560 (N_17560,N_17386,N_17258);
xnor U17561 (N_17561,N_17448,N_17354);
nand U17562 (N_17562,N_17014,N_17311);
or U17563 (N_17563,N_17326,N_17171);
nand U17564 (N_17564,N_17279,N_17256);
or U17565 (N_17565,N_17221,N_17498);
or U17566 (N_17566,N_17236,N_17088);
nand U17567 (N_17567,N_17199,N_17389);
nand U17568 (N_17568,N_17051,N_17454);
nand U17569 (N_17569,N_17353,N_17420);
nand U17570 (N_17570,N_17137,N_17481);
nand U17571 (N_17571,N_17074,N_17223);
nand U17572 (N_17572,N_17000,N_17460);
and U17573 (N_17573,N_17449,N_17023);
xor U17574 (N_17574,N_17488,N_17064);
nor U17575 (N_17575,N_17123,N_17245);
xnor U17576 (N_17576,N_17384,N_17349);
nand U17577 (N_17577,N_17465,N_17379);
and U17578 (N_17578,N_17380,N_17176);
xnor U17579 (N_17579,N_17166,N_17100);
xor U17580 (N_17580,N_17116,N_17292);
nor U17581 (N_17581,N_17239,N_17124);
or U17582 (N_17582,N_17190,N_17476);
nand U17583 (N_17583,N_17081,N_17364);
xor U17584 (N_17584,N_17113,N_17082);
nand U17585 (N_17585,N_17333,N_17328);
or U17586 (N_17586,N_17457,N_17118);
and U17587 (N_17587,N_17327,N_17156);
xnor U17588 (N_17588,N_17288,N_17234);
or U17589 (N_17589,N_17162,N_17076);
xnor U17590 (N_17590,N_17196,N_17005);
nor U17591 (N_17591,N_17342,N_17422);
xnor U17592 (N_17592,N_17398,N_17084);
nor U17593 (N_17593,N_17489,N_17225);
xnor U17594 (N_17594,N_17493,N_17028);
and U17595 (N_17595,N_17053,N_17185);
and U17596 (N_17596,N_17230,N_17401);
and U17597 (N_17597,N_17058,N_17153);
xnor U17598 (N_17598,N_17071,N_17033);
nand U17599 (N_17599,N_17418,N_17219);
nor U17600 (N_17600,N_17381,N_17385);
or U17601 (N_17601,N_17338,N_17272);
xnor U17602 (N_17602,N_17158,N_17347);
and U17603 (N_17603,N_17435,N_17344);
nand U17604 (N_17604,N_17324,N_17021);
nor U17605 (N_17605,N_17268,N_17263);
nor U17606 (N_17606,N_17154,N_17063);
nand U17607 (N_17607,N_17308,N_17304);
nor U17608 (N_17608,N_17450,N_17485);
xnor U17609 (N_17609,N_17208,N_17424);
and U17610 (N_17610,N_17421,N_17188);
nor U17611 (N_17611,N_17287,N_17334);
and U17612 (N_17612,N_17479,N_17144);
or U17613 (N_17613,N_17228,N_17464);
or U17614 (N_17614,N_17390,N_17172);
and U17615 (N_17615,N_17224,N_17321);
xnor U17616 (N_17616,N_17306,N_17201);
and U17617 (N_17617,N_17184,N_17285);
nor U17618 (N_17618,N_17370,N_17495);
or U17619 (N_17619,N_17174,N_17410);
nor U17620 (N_17620,N_17165,N_17341);
nor U17621 (N_17621,N_17213,N_17031);
nand U17622 (N_17622,N_17303,N_17373);
and U17623 (N_17623,N_17018,N_17105);
nand U17624 (N_17624,N_17249,N_17210);
or U17625 (N_17625,N_17473,N_17001);
and U17626 (N_17626,N_17131,N_17316);
or U17627 (N_17627,N_17241,N_17271);
xnor U17628 (N_17628,N_17455,N_17286);
nor U17629 (N_17629,N_17026,N_17491);
nor U17630 (N_17630,N_17083,N_17278);
nor U17631 (N_17631,N_17127,N_17050);
nor U17632 (N_17632,N_17198,N_17269);
or U17633 (N_17633,N_17202,N_17411);
or U17634 (N_17634,N_17393,N_17161);
nor U17635 (N_17635,N_17061,N_17107);
xnor U17636 (N_17636,N_17331,N_17170);
nand U17637 (N_17637,N_17042,N_17307);
and U17638 (N_17638,N_17348,N_17235);
nor U17639 (N_17639,N_17357,N_17260);
xnor U17640 (N_17640,N_17252,N_17178);
xnor U17641 (N_17641,N_17096,N_17309);
nor U17642 (N_17642,N_17044,N_17145);
and U17643 (N_17643,N_17106,N_17164);
and U17644 (N_17644,N_17019,N_17183);
xnor U17645 (N_17645,N_17483,N_17125);
xor U17646 (N_17646,N_17265,N_17431);
nand U17647 (N_17647,N_17492,N_17392);
and U17648 (N_17648,N_17356,N_17367);
or U17649 (N_17649,N_17078,N_17451);
nand U17650 (N_17650,N_17068,N_17405);
and U17651 (N_17651,N_17121,N_17126);
nor U17652 (N_17652,N_17173,N_17330);
or U17653 (N_17653,N_17136,N_17480);
or U17654 (N_17654,N_17340,N_17016);
xnor U17655 (N_17655,N_17242,N_17382);
or U17656 (N_17656,N_17300,N_17073);
nand U17657 (N_17657,N_17329,N_17013);
xor U17658 (N_17658,N_17102,N_17376);
nor U17659 (N_17659,N_17149,N_17002);
xnor U17660 (N_17660,N_17257,N_17360);
nand U17661 (N_17661,N_17264,N_17408);
nand U17662 (N_17662,N_17205,N_17446);
or U17663 (N_17663,N_17237,N_17459);
or U17664 (N_17664,N_17283,N_17262);
nand U17665 (N_17665,N_17434,N_17024);
or U17666 (N_17666,N_17274,N_17150);
xor U17667 (N_17667,N_17200,N_17244);
nor U17668 (N_17668,N_17395,N_17261);
or U17669 (N_17669,N_17117,N_17305);
or U17670 (N_17670,N_17254,N_17187);
and U17671 (N_17671,N_17046,N_17423);
nand U17672 (N_17672,N_17383,N_17099);
xnor U17673 (N_17673,N_17267,N_17355);
and U17674 (N_17674,N_17217,N_17152);
nor U17675 (N_17675,N_17404,N_17475);
and U17676 (N_17676,N_17253,N_17122);
nor U17677 (N_17677,N_17004,N_17070);
and U17678 (N_17678,N_17368,N_17365);
nand U17679 (N_17679,N_17066,N_17012);
and U17680 (N_17680,N_17240,N_17335);
and U17681 (N_17681,N_17375,N_17138);
nand U17682 (N_17682,N_17374,N_17346);
and U17683 (N_17683,N_17323,N_17414);
nand U17684 (N_17684,N_17467,N_17163);
nand U17685 (N_17685,N_17251,N_17319);
and U17686 (N_17686,N_17055,N_17281);
nor U17687 (N_17687,N_17468,N_17135);
nand U17688 (N_17688,N_17191,N_17216);
and U17689 (N_17689,N_17343,N_17314);
and U17690 (N_17690,N_17270,N_17218);
and U17691 (N_17691,N_17378,N_17438);
and U17692 (N_17692,N_17255,N_17430);
xnor U17693 (N_17693,N_17494,N_17222);
or U17694 (N_17694,N_17087,N_17436);
or U17695 (N_17695,N_17413,N_17160);
or U17696 (N_17696,N_17119,N_17299);
nand U17697 (N_17697,N_17377,N_17151);
and U17698 (N_17698,N_17233,N_17232);
xnor U17699 (N_17699,N_17243,N_17301);
and U17700 (N_17700,N_17060,N_17463);
and U17701 (N_17701,N_17147,N_17486);
nor U17702 (N_17702,N_17317,N_17447);
nand U17703 (N_17703,N_17211,N_17396);
or U17704 (N_17704,N_17215,N_17186);
nand U17705 (N_17705,N_17496,N_17077);
or U17706 (N_17706,N_17032,N_17006);
or U17707 (N_17707,N_17214,N_17209);
nand U17708 (N_17708,N_17291,N_17182);
xor U17709 (N_17709,N_17142,N_17115);
nand U17710 (N_17710,N_17345,N_17030);
or U17711 (N_17711,N_17069,N_17094);
nand U17712 (N_17712,N_17477,N_17295);
nand U17713 (N_17713,N_17155,N_17093);
or U17714 (N_17714,N_17369,N_17250);
or U17715 (N_17715,N_17312,N_17490);
or U17716 (N_17716,N_17015,N_17148);
and U17717 (N_17717,N_17289,N_17169);
and U17718 (N_17718,N_17441,N_17011);
or U17719 (N_17719,N_17318,N_17445);
or U17720 (N_17720,N_17175,N_17366);
xor U17721 (N_17721,N_17409,N_17143);
and U17722 (N_17722,N_17332,N_17426);
xnor U17723 (N_17723,N_17280,N_17432);
nor U17724 (N_17724,N_17466,N_17397);
nand U17725 (N_17725,N_17025,N_17108);
or U17726 (N_17726,N_17192,N_17111);
and U17727 (N_17727,N_17109,N_17157);
xnor U17728 (N_17728,N_17037,N_17248);
or U17729 (N_17729,N_17276,N_17059);
nand U17730 (N_17730,N_17193,N_17189);
and U17731 (N_17731,N_17469,N_17140);
xnor U17732 (N_17732,N_17229,N_17296);
xor U17733 (N_17733,N_17313,N_17363);
nor U17734 (N_17734,N_17277,N_17419);
or U17735 (N_17735,N_17034,N_17103);
or U17736 (N_17736,N_17478,N_17407);
nand U17737 (N_17737,N_17020,N_17134);
xnor U17738 (N_17738,N_17180,N_17204);
or U17739 (N_17739,N_17212,N_17325);
and U17740 (N_17740,N_17159,N_17440);
xor U17741 (N_17741,N_17057,N_17010);
xnor U17742 (N_17742,N_17052,N_17337);
nor U17743 (N_17743,N_17310,N_17259);
nor U17744 (N_17744,N_17101,N_17443);
nor U17745 (N_17745,N_17352,N_17417);
and U17746 (N_17746,N_17425,N_17141);
xor U17747 (N_17747,N_17075,N_17472);
xnor U17748 (N_17748,N_17035,N_17203);
nand U17749 (N_17749,N_17040,N_17336);
nor U17750 (N_17750,N_17067,N_17005);
or U17751 (N_17751,N_17177,N_17281);
xor U17752 (N_17752,N_17224,N_17159);
or U17753 (N_17753,N_17106,N_17419);
xor U17754 (N_17754,N_17132,N_17209);
nor U17755 (N_17755,N_17392,N_17365);
xor U17756 (N_17756,N_17471,N_17346);
nor U17757 (N_17757,N_17109,N_17116);
nor U17758 (N_17758,N_17403,N_17189);
xor U17759 (N_17759,N_17376,N_17254);
nand U17760 (N_17760,N_17107,N_17417);
xor U17761 (N_17761,N_17427,N_17365);
and U17762 (N_17762,N_17031,N_17079);
xor U17763 (N_17763,N_17284,N_17090);
nand U17764 (N_17764,N_17089,N_17027);
nand U17765 (N_17765,N_17297,N_17245);
nand U17766 (N_17766,N_17189,N_17275);
nor U17767 (N_17767,N_17245,N_17062);
nor U17768 (N_17768,N_17343,N_17277);
or U17769 (N_17769,N_17063,N_17455);
nand U17770 (N_17770,N_17316,N_17208);
or U17771 (N_17771,N_17232,N_17401);
nand U17772 (N_17772,N_17202,N_17219);
xnor U17773 (N_17773,N_17107,N_17150);
or U17774 (N_17774,N_17328,N_17446);
nor U17775 (N_17775,N_17201,N_17451);
xor U17776 (N_17776,N_17271,N_17253);
and U17777 (N_17777,N_17186,N_17034);
xnor U17778 (N_17778,N_17167,N_17218);
xor U17779 (N_17779,N_17380,N_17272);
xnor U17780 (N_17780,N_17467,N_17145);
nor U17781 (N_17781,N_17437,N_17010);
or U17782 (N_17782,N_17095,N_17069);
nor U17783 (N_17783,N_17127,N_17454);
nand U17784 (N_17784,N_17463,N_17025);
xor U17785 (N_17785,N_17420,N_17103);
and U17786 (N_17786,N_17046,N_17145);
nand U17787 (N_17787,N_17321,N_17344);
and U17788 (N_17788,N_17427,N_17146);
nor U17789 (N_17789,N_17202,N_17083);
nor U17790 (N_17790,N_17014,N_17163);
nand U17791 (N_17791,N_17075,N_17387);
and U17792 (N_17792,N_17491,N_17351);
xnor U17793 (N_17793,N_17399,N_17155);
nand U17794 (N_17794,N_17480,N_17135);
nor U17795 (N_17795,N_17308,N_17481);
nand U17796 (N_17796,N_17210,N_17233);
nor U17797 (N_17797,N_17236,N_17215);
or U17798 (N_17798,N_17467,N_17478);
nand U17799 (N_17799,N_17256,N_17420);
or U17800 (N_17800,N_17112,N_17251);
xnor U17801 (N_17801,N_17430,N_17051);
and U17802 (N_17802,N_17189,N_17163);
nor U17803 (N_17803,N_17148,N_17370);
nand U17804 (N_17804,N_17326,N_17016);
and U17805 (N_17805,N_17167,N_17425);
or U17806 (N_17806,N_17022,N_17325);
and U17807 (N_17807,N_17093,N_17013);
or U17808 (N_17808,N_17201,N_17498);
xor U17809 (N_17809,N_17344,N_17160);
nor U17810 (N_17810,N_17198,N_17073);
nor U17811 (N_17811,N_17033,N_17355);
xor U17812 (N_17812,N_17015,N_17305);
nand U17813 (N_17813,N_17466,N_17000);
or U17814 (N_17814,N_17074,N_17201);
and U17815 (N_17815,N_17004,N_17387);
xor U17816 (N_17816,N_17403,N_17494);
nor U17817 (N_17817,N_17397,N_17182);
xnor U17818 (N_17818,N_17251,N_17068);
or U17819 (N_17819,N_17450,N_17082);
or U17820 (N_17820,N_17017,N_17004);
or U17821 (N_17821,N_17057,N_17061);
nand U17822 (N_17822,N_17173,N_17157);
nand U17823 (N_17823,N_17229,N_17415);
nand U17824 (N_17824,N_17064,N_17472);
xnor U17825 (N_17825,N_17159,N_17255);
nor U17826 (N_17826,N_17175,N_17377);
nand U17827 (N_17827,N_17106,N_17268);
xor U17828 (N_17828,N_17247,N_17191);
nor U17829 (N_17829,N_17082,N_17092);
and U17830 (N_17830,N_17462,N_17109);
xnor U17831 (N_17831,N_17453,N_17177);
and U17832 (N_17832,N_17475,N_17241);
or U17833 (N_17833,N_17077,N_17064);
nor U17834 (N_17834,N_17283,N_17464);
xor U17835 (N_17835,N_17023,N_17207);
nand U17836 (N_17836,N_17196,N_17161);
nor U17837 (N_17837,N_17323,N_17013);
xnor U17838 (N_17838,N_17044,N_17012);
nor U17839 (N_17839,N_17059,N_17032);
xor U17840 (N_17840,N_17229,N_17310);
and U17841 (N_17841,N_17071,N_17024);
and U17842 (N_17842,N_17056,N_17070);
nor U17843 (N_17843,N_17423,N_17473);
xnor U17844 (N_17844,N_17370,N_17190);
xnor U17845 (N_17845,N_17303,N_17296);
nand U17846 (N_17846,N_17270,N_17097);
xor U17847 (N_17847,N_17330,N_17391);
and U17848 (N_17848,N_17276,N_17435);
or U17849 (N_17849,N_17190,N_17458);
and U17850 (N_17850,N_17008,N_17338);
xnor U17851 (N_17851,N_17381,N_17175);
or U17852 (N_17852,N_17259,N_17062);
nor U17853 (N_17853,N_17097,N_17396);
nor U17854 (N_17854,N_17355,N_17286);
nor U17855 (N_17855,N_17189,N_17064);
nor U17856 (N_17856,N_17429,N_17421);
nand U17857 (N_17857,N_17307,N_17250);
or U17858 (N_17858,N_17102,N_17346);
and U17859 (N_17859,N_17287,N_17408);
nand U17860 (N_17860,N_17400,N_17140);
nor U17861 (N_17861,N_17115,N_17000);
or U17862 (N_17862,N_17498,N_17436);
nand U17863 (N_17863,N_17281,N_17285);
and U17864 (N_17864,N_17445,N_17144);
nor U17865 (N_17865,N_17250,N_17291);
nor U17866 (N_17866,N_17223,N_17374);
nor U17867 (N_17867,N_17490,N_17361);
nor U17868 (N_17868,N_17079,N_17194);
and U17869 (N_17869,N_17212,N_17302);
or U17870 (N_17870,N_17235,N_17336);
nor U17871 (N_17871,N_17441,N_17484);
or U17872 (N_17872,N_17313,N_17075);
xor U17873 (N_17873,N_17447,N_17403);
xnor U17874 (N_17874,N_17401,N_17264);
xnor U17875 (N_17875,N_17215,N_17088);
nand U17876 (N_17876,N_17422,N_17489);
and U17877 (N_17877,N_17282,N_17384);
or U17878 (N_17878,N_17143,N_17209);
nor U17879 (N_17879,N_17123,N_17125);
and U17880 (N_17880,N_17352,N_17158);
and U17881 (N_17881,N_17333,N_17167);
and U17882 (N_17882,N_17074,N_17052);
nor U17883 (N_17883,N_17210,N_17028);
or U17884 (N_17884,N_17089,N_17256);
and U17885 (N_17885,N_17055,N_17111);
nor U17886 (N_17886,N_17041,N_17251);
or U17887 (N_17887,N_17013,N_17425);
xor U17888 (N_17888,N_17376,N_17140);
or U17889 (N_17889,N_17394,N_17438);
nor U17890 (N_17890,N_17023,N_17420);
or U17891 (N_17891,N_17217,N_17428);
nor U17892 (N_17892,N_17381,N_17170);
and U17893 (N_17893,N_17031,N_17000);
xnor U17894 (N_17894,N_17363,N_17155);
and U17895 (N_17895,N_17036,N_17079);
nand U17896 (N_17896,N_17116,N_17137);
nand U17897 (N_17897,N_17065,N_17107);
or U17898 (N_17898,N_17065,N_17020);
and U17899 (N_17899,N_17023,N_17314);
nand U17900 (N_17900,N_17005,N_17420);
nor U17901 (N_17901,N_17047,N_17456);
nor U17902 (N_17902,N_17210,N_17396);
nand U17903 (N_17903,N_17412,N_17296);
nand U17904 (N_17904,N_17201,N_17191);
and U17905 (N_17905,N_17014,N_17374);
and U17906 (N_17906,N_17251,N_17172);
and U17907 (N_17907,N_17023,N_17240);
nand U17908 (N_17908,N_17093,N_17029);
xor U17909 (N_17909,N_17307,N_17463);
nand U17910 (N_17910,N_17135,N_17421);
or U17911 (N_17911,N_17220,N_17386);
or U17912 (N_17912,N_17192,N_17466);
or U17913 (N_17913,N_17244,N_17363);
nor U17914 (N_17914,N_17140,N_17497);
nand U17915 (N_17915,N_17369,N_17332);
nand U17916 (N_17916,N_17288,N_17362);
nand U17917 (N_17917,N_17143,N_17250);
and U17918 (N_17918,N_17285,N_17499);
and U17919 (N_17919,N_17051,N_17462);
nor U17920 (N_17920,N_17261,N_17026);
xnor U17921 (N_17921,N_17143,N_17425);
nand U17922 (N_17922,N_17467,N_17213);
nand U17923 (N_17923,N_17275,N_17169);
xor U17924 (N_17924,N_17037,N_17160);
nand U17925 (N_17925,N_17361,N_17271);
nand U17926 (N_17926,N_17147,N_17490);
nand U17927 (N_17927,N_17437,N_17050);
and U17928 (N_17928,N_17283,N_17079);
and U17929 (N_17929,N_17484,N_17162);
nor U17930 (N_17930,N_17076,N_17448);
xnor U17931 (N_17931,N_17379,N_17380);
xnor U17932 (N_17932,N_17331,N_17042);
nand U17933 (N_17933,N_17228,N_17147);
xnor U17934 (N_17934,N_17091,N_17263);
xnor U17935 (N_17935,N_17147,N_17212);
nand U17936 (N_17936,N_17252,N_17438);
or U17937 (N_17937,N_17390,N_17149);
nand U17938 (N_17938,N_17428,N_17007);
and U17939 (N_17939,N_17147,N_17150);
nor U17940 (N_17940,N_17030,N_17019);
nor U17941 (N_17941,N_17259,N_17006);
or U17942 (N_17942,N_17015,N_17404);
or U17943 (N_17943,N_17140,N_17059);
nand U17944 (N_17944,N_17366,N_17095);
and U17945 (N_17945,N_17032,N_17258);
nor U17946 (N_17946,N_17286,N_17116);
nor U17947 (N_17947,N_17152,N_17120);
and U17948 (N_17948,N_17420,N_17097);
xor U17949 (N_17949,N_17140,N_17095);
nand U17950 (N_17950,N_17350,N_17002);
nand U17951 (N_17951,N_17359,N_17386);
nand U17952 (N_17952,N_17156,N_17105);
xor U17953 (N_17953,N_17000,N_17442);
or U17954 (N_17954,N_17154,N_17146);
nor U17955 (N_17955,N_17212,N_17378);
and U17956 (N_17956,N_17061,N_17441);
nand U17957 (N_17957,N_17374,N_17230);
and U17958 (N_17958,N_17029,N_17269);
or U17959 (N_17959,N_17033,N_17414);
xor U17960 (N_17960,N_17002,N_17240);
nand U17961 (N_17961,N_17380,N_17246);
and U17962 (N_17962,N_17148,N_17261);
xor U17963 (N_17963,N_17333,N_17316);
nor U17964 (N_17964,N_17158,N_17259);
and U17965 (N_17965,N_17448,N_17347);
xor U17966 (N_17966,N_17499,N_17206);
nand U17967 (N_17967,N_17121,N_17467);
xor U17968 (N_17968,N_17084,N_17211);
and U17969 (N_17969,N_17387,N_17048);
xor U17970 (N_17970,N_17364,N_17049);
nand U17971 (N_17971,N_17268,N_17087);
nor U17972 (N_17972,N_17103,N_17304);
nor U17973 (N_17973,N_17325,N_17491);
and U17974 (N_17974,N_17229,N_17069);
xnor U17975 (N_17975,N_17256,N_17134);
nand U17976 (N_17976,N_17012,N_17222);
or U17977 (N_17977,N_17384,N_17007);
nand U17978 (N_17978,N_17358,N_17445);
and U17979 (N_17979,N_17072,N_17405);
or U17980 (N_17980,N_17210,N_17243);
nand U17981 (N_17981,N_17158,N_17431);
and U17982 (N_17982,N_17154,N_17086);
nor U17983 (N_17983,N_17383,N_17126);
or U17984 (N_17984,N_17447,N_17412);
nor U17985 (N_17985,N_17018,N_17463);
xor U17986 (N_17986,N_17347,N_17402);
and U17987 (N_17987,N_17191,N_17121);
nand U17988 (N_17988,N_17421,N_17132);
xor U17989 (N_17989,N_17088,N_17420);
nand U17990 (N_17990,N_17046,N_17187);
nor U17991 (N_17991,N_17448,N_17312);
nor U17992 (N_17992,N_17347,N_17092);
and U17993 (N_17993,N_17179,N_17424);
nor U17994 (N_17994,N_17258,N_17039);
nand U17995 (N_17995,N_17246,N_17203);
nor U17996 (N_17996,N_17468,N_17257);
nor U17997 (N_17997,N_17056,N_17267);
nor U17998 (N_17998,N_17421,N_17306);
nand U17999 (N_17999,N_17413,N_17396);
xnor U18000 (N_18000,N_17964,N_17737);
nand U18001 (N_18001,N_17808,N_17999);
or U18002 (N_18002,N_17614,N_17720);
or U18003 (N_18003,N_17899,N_17602);
nand U18004 (N_18004,N_17761,N_17634);
xor U18005 (N_18005,N_17684,N_17756);
nand U18006 (N_18006,N_17523,N_17544);
and U18007 (N_18007,N_17706,N_17975);
or U18008 (N_18008,N_17654,N_17510);
nor U18009 (N_18009,N_17838,N_17850);
and U18010 (N_18010,N_17922,N_17712);
or U18011 (N_18011,N_17960,N_17879);
xor U18012 (N_18012,N_17580,N_17653);
or U18013 (N_18013,N_17529,N_17941);
xor U18014 (N_18014,N_17525,N_17547);
and U18015 (N_18015,N_17983,N_17900);
nand U18016 (N_18016,N_17567,N_17957);
nor U18017 (N_18017,N_17500,N_17696);
nand U18018 (N_18018,N_17577,N_17767);
and U18019 (N_18019,N_17929,N_17658);
xnor U18020 (N_18020,N_17889,N_17804);
xor U18021 (N_18021,N_17616,N_17886);
nand U18022 (N_18022,N_17932,N_17652);
and U18023 (N_18023,N_17656,N_17594);
xor U18024 (N_18024,N_17662,N_17583);
xnor U18025 (N_18025,N_17512,N_17526);
nand U18026 (N_18026,N_17931,N_17503);
nand U18027 (N_18027,N_17752,N_17782);
xor U18028 (N_18028,N_17572,N_17631);
nand U18029 (N_18029,N_17518,N_17953);
nor U18030 (N_18030,N_17743,N_17686);
nor U18031 (N_18031,N_17667,N_17853);
nand U18032 (N_18032,N_17536,N_17781);
or U18033 (N_18033,N_17559,N_17777);
or U18034 (N_18034,N_17501,N_17534);
or U18035 (N_18035,N_17934,N_17611);
xor U18036 (N_18036,N_17912,N_17671);
nand U18037 (N_18037,N_17968,N_17998);
xor U18038 (N_18038,N_17540,N_17982);
or U18039 (N_18039,N_17717,N_17558);
xor U18040 (N_18040,N_17507,N_17590);
nor U18041 (N_18041,N_17660,N_17798);
nand U18042 (N_18042,N_17659,N_17877);
nand U18043 (N_18043,N_17775,N_17681);
nor U18044 (N_18044,N_17903,N_17857);
nor U18045 (N_18045,N_17817,N_17589);
xor U18046 (N_18046,N_17966,N_17704);
or U18047 (N_18047,N_17945,N_17736);
xnor U18048 (N_18048,N_17582,N_17869);
and U18049 (N_18049,N_17576,N_17876);
or U18050 (N_18050,N_17833,N_17849);
nand U18051 (N_18051,N_17919,N_17679);
or U18052 (N_18052,N_17763,N_17640);
or U18053 (N_18053,N_17649,N_17618);
or U18054 (N_18054,N_17548,N_17758);
xor U18055 (N_18055,N_17701,N_17890);
nor U18056 (N_18056,N_17783,N_17595);
xnor U18057 (N_18057,N_17861,N_17663);
nor U18058 (N_18058,N_17605,N_17848);
xor U18059 (N_18059,N_17599,N_17830);
and U18060 (N_18060,N_17753,N_17713);
xor U18061 (N_18061,N_17562,N_17601);
and U18062 (N_18062,N_17754,N_17949);
xor U18063 (N_18063,N_17623,N_17506);
and U18064 (N_18064,N_17994,N_17979);
xnor U18065 (N_18065,N_17827,N_17748);
xor U18066 (N_18066,N_17731,N_17913);
nor U18067 (N_18067,N_17944,N_17584);
nor U18068 (N_18068,N_17710,N_17722);
nand U18069 (N_18069,N_17571,N_17887);
nor U18070 (N_18070,N_17511,N_17757);
nor U18071 (N_18071,N_17788,N_17709);
nand U18072 (N_18072,N_17759,N_17627);
nor U18073 (N_18073,N_17832,N_17517);
and U18074 (N_18074,N_17780,N_17956);
or U18075 (N_18075,N_17539,N_17508);
nor U18076 (N_18076,N_17530,N_17978);
and U18077 (N_18077,N_17892,N_17764);
and U18078 (N_18078,N_17588,N_17606);
nor U18079 (N_18079,N_17930,N_17906);
nor U18080 (N_18080,N_17561,N_17772);
or U18081 (N_18081,N_17924,N_17809);
or U18082 (N_18082,N_17888,N_17778);
xor U18083 (N_18083,N_17733,N_17708);
and U18084 (N_18084,N_17823,N_17741);
nor U18085 (N_18085,N_17799,N_17825);
xnor U18086 (N_18086,N_17672,N_17883);
or U18087 (N_18087,N_17793,N_17801);
and U18088 (N_18088,N_17661,N_17625);
nand U18089 (N_18089,N_17537,N_17776);
nor U18090 (N_18090,N_17993,N_17522);
nand U18091 (N_18091,N_17624,N_17805);
and U18092 (N_18092,N_17990,N_17995);
xor U18093 (N_18093,N_17920,N_17987);
and U18094 (N_18094,N_17824,N_17894);
nor U18095 (N_18095,N_17598,N_17555);
nor U18096 (N_18096,N_17644,N_17642);
nor U18097 (N_18097,N_17845,N_17608);
and U18098 (N_18098,N_17641,N_17648);
xnor U18099 (N_18099,N_17746,N_17870);
xor U18100 (N_18100,N_17792,N_17750);
nand U18101 (N_18101,N_17976,N_17875);
xor U18102 (N_18102,N_17665,N_17586);
nor U18103 (N_18103,N_17635,N_17785);
nand U18104 (N_18104,N_17749,N_17923);
nand U18105 (N_18105,N_17666,N_17810);
or U18106 (N_18106,N_17504,N_17600);
xor U18107 (N_18107,N_17936,N_17997);
or U18108 (N_18108,N_17791,N_17981);
or U18109 (N_18109,N_17839,N_17829);
nand U18110 (N_18110,N_17779,N_17790);
and U18111 (N_18111,N_17612,N_17867);
xnor U18112 (N_18112,N_17643,N_17573);
nand U18113 (N_18113,N_17868,N_17578);
and U18114 (N_18114,N_17939,N_17692);
and U18115 (N_18115,N_17570,N_17747);
nor U18116 (N_18116,N_17543,N_17871);
or U18117 (N_18117,N_17980,N_17811);
nand U18118 (N_18118,N_17911,N_17745);
nand U18119 (N_18119,N_17732,N_17581);
nor U18120 (N_18120,N_17991,N_17961);
nor U18121 (N_18121,N_17687,N_17766);
nor U18122 (N_18122,N_17513,N_17509);
and U18123 (N_18123,N_17866,N_17755);
nor U18124 (N_18124,N_17865,N_17996);
nor U18125 (N_18125,N_17552,N_17955);
nand U18126 (N_18126,N_17514,N_17933);
xnor U18127 (N_18127,N_17771,N_17915);
xnor U18128 (N_18128,N_17768,N_17657);
nand U18129 (N_18129,N_17551,N_17637);
xor U18130 (N_18130,N_17615,N_17673);
nor U18131 (N_18131,N_17925,N_17596);
nand U18132 (N_18132,N_17770,N_17951);
nor U18133 (N_18133,N_17988,N_17650);
xnor U18134 (N_18134,N_17647,N_17854);
nor U18135 (N_18135,N_17840,N_17897);
and U18136 (N_18136,N_17632,N_17813);
and U18137 (N_18137,N_17744,N_17950);
nand U18138 (N_18138,N_17986,N_17689);
nor U18139 (N_18139,N_17505,N_17621);
and U18140 (N_18140,N_17694,N_17928);
or U18141 (N_18141,N_17693,N_17702);
and U18142 (N_18142,N_17921,N_17896);
xnor U18143 (N_18143,N_17834,N_17727);
nand U18144 (N_18144,N_17837,N_17683);
nor U18145 (N_18145,N_17715,N_17843);
nand U18146 (N_18146,N_17639,N_17729);
and U18147 (N_18147,N_17787,N_17970);
and U18148 (N_18148,N_17989,N_17553);
or U18149 (N_18149,N_17751,N_17734);
nand U18150 (N_18150,N_17730,N_17958);
or U18151 (N_18151,N_17864,N_17682);
and U18152 (N_18152,N_17893,N_17760);
nor U18153 (N_18153,N_17882,N_17620);
xor U18154 (N_18154,N_17855,N_17963);
nor U18155 (N_18155,N_17568,N_17520);
xor U18156 (N_18156,N_17532,N_17762);
or U18157 (N_18157,N_17806,N_17846);
nand U18158 (N_18158,N_17962,N_17677);
or U18159 (N_18159,N_17742,N_17971);
nand U18160 (N_18160,N_17918,N_17695);
or U18161 (N_18161,N_17528,N_17569);
nand U18162 (N_18162,N_17863,N_17566);
or U18163 (N_18163,N_17972,N_17628);
and U18164 (N_18164,N_17914,N_17985);
xnor U18165 (N_18165,N_17574,N_17784);
nor U18166 (N_18166,N_17691,N_17844);
and U18167 (N_18167,N_17698,N_17926);
and U18168 (N_18168,N_17802,N_17916);
or U18169 (N_18169,N_17585,N_17593);
nor U18170 (N_18170,N_17974,N_17820);
nor U18171 (N_18171,N_17575,N_17909);
and U18172 (N_18172,N_17527,N_17638);
xnor U18173 (N_18173,N_17674,N_17794);
xor U18174 (N_18174,N_17862,N_17554);
or U18175 (N_18175,N_17872,N_17609);
and U18176 (N_18176,N_17735,N_17795);
nor U18177 (N_18177,N_17533,N_17847);
nor U18178 (N_18178,N_17895,N_17622);
xnor U18179 (N_18179,N_17908,N_17942);
or U18180 (N_18180,N_17917,N_17685);
or U18181 (N_18181,N_17550,N_17629);
xnor U18182 (N_18182,N_17814,N_17714);
nand U18183 (N_18183,N_17797,N_17579);
or U18184 (N_18184,N_17564,N_17724);
nand U18185 (N_18185,N_17901,N_17556);
xor U18186 (N_18186,N_17828,N_17664);
or U18187 (N_18187,N_17563,N_17874);
and U18188 (N_18188,N_17856,N_17592);
nand U18189 (N_18189,N_17969,N_17852);
nor U18190 (N_18190,N_17519,N_17549);
xor U18191 (N_18191,N_17699,N_17905);
or U18192 (N_18192,N_17557,N_17947);
or U18193 (N_18193,N_17952,N_17940);
nand U18194 (N_18194,N_17954,N_17878);
xnor U18195 (N_18195,N_17819,N_17880);
nor U18196 (N_18196,N_17835,N_17705);
and U18197 (N_18197,N_17630,N_17774);
or U18198 (N_18198,N_17626,N_17617);
nand U18199 (N_18199,N_17688,N_17800);
xnor U18200 (N_18200,N_17977,N_17858);
xnor U18201 (N_18201,N_17927,N_17907);
nand U18202 (N_18202,N_17891,N_17884);
nor U18203 (N_18203,N_17984,N_17938);
nand U18204 (N_18204,N_17531,N_17822);
nand U18205 (N_18205,N_17965,N_17670);
xnor U18206 (N_18206,N_17740,N_17613);
xor U18207 (N_18207,N_17786,N_17992);
xor U18208 (N_18208,N_17807,N_17675);
nor U18209 (N_18209,N_17910,N_17946);
or U18210 (N_18210,N_17603,N_17703);
or U18211 (N_18211,N_17524,N_17812);
nand U18212 (N_18212,N_17816,N_17587);
xnor U18213 (N_18213,N_17591,N_17610);
and U18214 (N_18214,N_17726,N_17836);
and U18215 (N_18215,N_17560,N_17597);
nand U18216 (N_18216,N_17604,N_17898);
xor U18217 (N_18217,N_17765,N_17678);
xnor U18218 (N_18218,N_17697,N_17769);
or U18219 (N_18219,N_17716,N_17516);
and U18220 (N_18220,N_17859,N_17535);
or U18221 (N_18221,N_17607,N_17739);
and U18222 (N_18222,N_17789,N_17719);
nand U18223 (N_18223,N_17948,N_17860);
xor U18224 (N_18224,N_17815,N_17873);
nand U18225 (N_18225,N_17645,N_17851);
xnor U18226 (N_18226,N_17646,N_17669);
and U18227 (N_18227,N_17841,N_17668);
xnor U18228 (N_18228,N_17935,N_17651);
xnor U18229 (N_18229,N_17723,N_17636);
nand U18230 (N_18230,N_17818,N_17796);
nor U18231 (N_18231,N_17826,N_17773);
and U18232 (N_18232,N_17803,N_17902);
and U18233 (N_18233,N_17546,N_17619);
nor U18234 (N_18234,N_17515,N_17725);
and U18235 (N_18235,N_17711,N_17502);
xnor U18236 (N_18236,N_17633,N_17538);
nor U18237 (N_18237,N_17676,N_17565);
xnor U18238 (N_18238,N_17521,N_17655);
or U18239 (N_18239,N_17967,N_17821);
xor U18240 (N_18240,N_17541,N_17721);
and U18241 (N_18241,N_17700,N_17831);
nor U18242 (N_18242,N_17885,N_17937);
nand U18243 (N_18243,N_17959,N_17542);
nand U18244 (N_18244,N_17690,N_17707);
nor U18245 (N_18245,N_17973,N_17728);
or U18246 (N_18246,N_17738,N_17881);
xor U18247 (N_18247,N_17842,N_17943);
xor U18248 (N_18248,N_17904,N_17545);
and U18249 (N_18249,N_17718,N_17680);
nor U18250 (N_18250,N_17518,N_17537);
xor U18251 (N_18251,N_17613,N_17930);
or U18252 (N_18252,N_17515,N_17974);
and U18253 (N_18253,N_17664,N_17501);
or U18254 (N_18254,N_17876,N_17538);
xnor U18255 (N_18255,N_17732,N_17842);
or U18256 (N_18256,N_17789,N_17862);
xnor U18257 (N_18257,N_17687,N_17716);
nor U18258 (N_18258,N_17883,N_17839);
or U18259 (N_18259,N_17569,N_17754);
nor U18260 (N_18260,N_17564,N_17960);
or U18261 (N_18261,N_17822,N_17599);
nor U18262 (N_18262,N_17615,N_17722);
nor U18263 (N_18263,N_17751,N_17756);
and U18264 (N_18264,N_17652,N_17847);
and U18265 (N_18265,N_17827,N_17750);
or U18266 (N_18266,N_17785,N_17844);
nand U18267 (N_18267,N_17719,N_17966);
and U18268 (N_18268,N_17724,N_17826);
xnor U18269 (N_18269,N_17802,N_17678);
nand U18270 (N_18270,N_17748,N_17631);
nor U18271 (N_18271,N_17948,N_17534);
xnor U18272 (N_18272,N_17667,N_17811);
xor U18273 (N_18273,N_17604,N_17631);
or U18274 (N_18274,N_17957,N_17576);
nor U18275 (N_18275,N_17585,N_17973);
nor U18276 (N_18276,N_17748,N_17676);
xnor U18277 (N_18277,N_17620,N_17836);
or U18278 (N_18278,N_17726,N_17964);
xnor U18279 (N_18279,N_17911,N_17521);
xnor U18280 (N_18280,N_17920,N_17565);
and U18281 (N_18281,N_17849,N_17543);
nand U18282 (N_18282,N_17865,N_17746);
or U18283 (N_18283,N_17831,N_17625);
xnor U18284 (N_18284,N_17549,N_17556);
xnor U18285 (N_18285,N_17888,N_17648);
xnor U18286 (N_18286,N_17806,N_17991);
nand U18287 (N_18287,N_17540,N_17887);
and U18288 (N_18288,N_17746,N_17902);
nor U18289 (N_18289,N_17794,N_17666);
nor U18290 (N_18290,N_17789,N_17612);
and U18291 (N_18291,N_17761,N_17916);
xor U18292 (N_18292,N_17953,N_17657);
or U18293 (N_18293,N_17633,N_17881);
xnor U18294 (N_18294,N_17978,N_17888);
and U18295 (N_18295,N_17983,N_17966);
or U18296 (N_18296,N_17565,N_17890);
and U18297 (N_18297,N_17998,N_17620);
nand U18298 (N_18298,N_17836,N_17617);
nor U18299 (N_18299,N_17778,N_17514);
nand U18300 (N_18300,N_17524,N_17645);
or U18301 (N_18301,N_17734,N_17666);
xor U18302 (N_18302,N_17888,N_17753);
and U18303 (N_18303,N_17827,N_17838);
nor U18304 (N_18304,N_17658,N_17979);
xor U18305 (N_18305,N_17911,N_17798);
nor U18306 (N_18306,N_17635,N_17856);
xnor U18307 (N_18307,N_17660,N_17540);
nand U18308 (N_18308,N_17894,N_17561);
or U18309 (N_18309,N_17709,N_17862);
nand U18310 (N_18310,N_17889,N_17897);
nand U18311 (N_18311,N_17614,N_17935);
or U18312 (N_18312,N_17542,N_17982);
and U18313 (N_18313,N_17518,N_17568);
or U18314 (N_18314,N_17764,N_17596);
xnor U18315 (N_18315,N_17691,N_17627);
xnor U18316 (N_18316,N_17896,N_17922);
nand U18317 (N_18317,N_17691,N_17750);
nor U18318 (N_18318,N_17849,N_17916);
nor U18319 (N_18319,N_17951,N_17694);
and U18320 (N_18320,N_17623,N_17522);
and U18321 (N_18321,N_17753,N_17592);
and U18322 (N_18322,N_17794,N_17865);
xnor U18323 (N_18323,N_17965,N_17763);
and U18324 (N_18324,N_17770,N_17744);
and U18325 (N_18325,N_17953,N_17923);
nand U18326 (N_18326,N_17631,N_17822);
nor U18327 (N_18327,N_17825,N_17633);
xor U18328 (N_18328,N_17789,N_17889);
and U18329 (N_18329,N_17772,N_17529);
or U18330 (N_18330,N_17874,N_17745);
and U18331 (N_18331,N_17715,N_17574);
or U18332 (N_18332,N_17918,N_17686);
and U18333 (N_18333,N_17546,N_17783);
or U18334 (N_18334,N_17871,N_17933);
xor U18335 (N_18335,N_17653,N_17944);
xor U18336 (N_18336,N_17512,N_17962);
nor U18337 (N_18337,N_17955,N_17729);
and U18338 (N_18338,N_17680,N_17723);
xor U18339 (N_18339,N_17579,N_17922);
or U18340 (N_18340,N_17757,N_17575);
and U18341 (N_18341,N_17860,N_17693);
and U18342 (N_18342,N_17538,N_17857);
and U18343 (N_18343,N_17916,N_17625);
and U18344 (N_18344,N_17739,N_17654);
xor U18345 (N_18345,N_17530,N_17668);
and U18346 (N_18346,N_17570,N_17912);
and U18347 (N_18347,N_17964,N_17960);
or U18348 (N_18348,N_17822,N_17955);
nor U18349 (N_18349,N_17758,N_17713);
nand U18350 (N_18350,N_17852,N_17694);
nand U18351 (N_18351,N_17641,N_17609);
nand U18352 (N_18352,N_17689,N_17529);
or U18353 (N_18353,N_17828,N_17580);
xnor U18354 (N_18354,N_17955,N_17940);
and U18355 (N_18355,N_17825,N_17874);
nand U18356 (N_18356,N_17664,N_17913);
or U18357 (N_18357,N_17518,N_17572);
or U18358 (N_18358,N_17782,N_17873);
nand U18359 (N_18359,N_17905,N_17850);
nand U18360 (N_18360,N_17640,N_17575);
nor U18361 (N_18361,N_17534,N_17688);
or U18362 (N_18362,N_17678,N_17653);
and U18363 (N_18363,N_17788,N_17977);
nand U18364 (N_18364,N_17665,N_17944);
or U18365 (N_18365,N_17941,N_17653);
nand U18366 (N_18366,N_17856,N_17826);
or U18367 (N_18367,N_17954,N_17591);
nand U18368 (N_18368,N_17562,N_17884);
and U18369 (N_18369,N_17991,N_17528);
xnor U18370 (N_18370,N_17739,N_17876);
and U18371 (N_18371,N_17906,N_17671);
nand U18372 (N_18372,N_17764,N_17967);
nand U18373 (N_18373,N_17607,N_17558);
nor U18374 (N_18374,N_17622,N_17926);
xnor U18375 (N_18375,N_17602,N_17664);
or U18376 (N_18376,N_17568,N_17814);
xnor U18377 (N_18377,N_17614,N_17686);
nand U18378 (N_18378,N_17570,N_17513);
xnor U18379 (N_18379,N_17667,N_17845);
or U18380 (N_18380,N_17897,N_17976);
nor U18381 (N_18381,N_17991,N_17527);
nand U18382 (N_18382,N_17506,N_17518);
or U18383 (N_18383,N_17563,N_17560);
and U18384 (N_18384,N_17795,N_17777);
xor U18385 (N_18385,N_17924,N_17902);
xnor U18386 (N_18386,N_17796,N_17503);
or U18387 (N_18387,N_17903,N_17807);
nand U18388 (N_18388,N_17544,N_17646);
or U18389 (N_18389,N_17694,N_17556);
xor U18390 (N_18390,N_17530,N_17995);
and U18391 (N_18391,N_17890,N_17576);
nand U18392 (N_18392,N_17744,N_17817);
or U18393 (N_18393,N_17638,N_17738);
nand U18394 (N_18394,N_17594,N_17608);
nor U18395 (N_18395,N_17577,N_17628);
or U18396 (N_18396,N_17959,N_17879);
nor U18397 (N_18397,N_17887,N_17842);
and U18398 (N_18398,N_17806,N_17775);
or U18399 (N_18399,N_17707,N_17714);
or U18400 (N_18400,N_17772,N_17939);
and U18401 (N_18401,N_17514,N_17941);
nor U18402 (N_18402,N_17945,N_17723);
nand U18403 (N_18403,N_17697,N_17787);
nand U18404 (N_18404,N_17802,N_17999);
nand U18405 (N_18405,N_17776,N_17856);
and U18406 (N_18406,N_17656,N_17771);
nor U18407 (N_18407,N_17940,N_17553);
nor U18408 (N_18408,N_17500,N_17734);
or U18409 (N_18409,N_17860,N_17774);
xnor U18410 (N_18410,N_17836,N_17556);
or U18411 (N_18411,N_17829,N_17524);
and U18412 (N_18412,N_17974,N_17882);
or U18413 (N_18413,N_17515,N_17612);
nor U18414 (N_18414,N_17728,N_17580);
nor U18415 (N_18415,N_17531,N_17602);
or U18416 (N_18416,N_17824,N_17785);
nor U18417 (N_18417,N_17796,N_17725);
or U18418 (N_18418,N_17647,N_17612);
xnor U18419 (N_18419,N_17694,N_17595);
nand U18420 (N_18420,N_17686,N_17524);
nand U18421 (N_18421,N_17979,N_17986);
and U18422 (N_18422,N_17697,N_17556);
nor U18423 (N_18423,N_17823,N_17623);
xnor U18424 (N_18424,N_17709,N_17959);
xor U18425 (N_18425,N_17642,N_17597);
nor U18426 (N_18426,N_17595,N_17601);
nand U18427 (N_18427,N_17668,N_17615);
and U18428 (N_18428,N_17926,N_17735);
nor U18429 (N_18429,N_17749,N_17754);
nand U18430 (N_18430,N_17503,N_17849);
xnor U18431 (N_18431,N_17832,N_17608);
nand U18432 (N_18432,N_17856,N_17509);
xnor U18433 (N_18433,N_17584,N_17930);
or U18434 (N_18434,N_17810,N_17881);
xnor U18435 (N_18435,N_17801,N_17578);
nor U18436 (N_18436,N_17612,N_17538);
and U18437 (N_18437,N_17604,N_17969);
and U18438 (N_18438,N_17972,N_17960);
or U18439 (N_18439,N_17667,N_17506);
nor U18440 (N_18440,N_17557,N_17742);
or U18441 (N_18441,N_17715,N_17956);
nand U18442 (N_18442,N_17929,N_17830);
nor U18443 (N_18443,N_17869,N_17838);
nand U18444 (N_18444,N_17952,N_17885);
or U18445 (N_18445,N_17954,N_17696);
and U18446 (N_18446,N_17527,N_17835);
xnor U18447 (N_18447,N_17796,N_17891);
and U18448 (N_18448,N_17636,N_17798);
nand U18449 (N_18449,N_17813,N_17922);
nor U18450 (N_18450,N_17787,N_17790);
nor U18451 (N_18451,N_17867,N_17803);
or U18452 (N_18452,N_17830,N_17963);
xnor U18453 (N_18453,N_17718,N_17822);
xor U18454 (N_18454,N_17667,N_17891);
nor U18455 (N_18455,N_17933,N_17565);
nor U18456 (N_18456,N_17895,N_17598);
and U18457 (N_18457,N_17701,N_17863);
nand U18458 (N_18458,N_17615,N_17769);
or U18459 (N_18459,N_17937,N_17787);
nand U18460 (N_18460,N_17873,N_17536);
or U18461 (N_18461,N_17649,N_17663);
nand U18462 (N_18462,N_17977,N_17759);
or U18463 (N_18463,N_17916,N_17912);
and U18464 (N_18464,N_17910,N_17696);
or U18465 (N_18465,N_17895,N_17747);
or U18466 (N_18466,N_17966,N_17825);
xnor U18467 (N_18467,N_17621,N_17810);
nand U18468 (N_18468,N_17545,N_17533);
and U18469 (N_18469,N_17734,N_17787);
nor U18470 (N_18470,N_17782,N_17621);
nor U18471 (N_18471,N_17674,N_17973);
nor U18472 (N_18472,N_17520,N_17644);
or U18473 (N_18473,N_17648,N_17862);
nand U18474 (N_18474,N_17542,N_17616);
xnor U18475 (N_18475,N_17985,N_17956);
xnor U18476 (N_18476,N_17789,N_17670);
and U18477 (N_18477,N_17590,N_17554);
nor U18478 (N_18478,N_17875,N_17847);
xnor U18479 (N_18479,N_17848,N_17895);
or U18480 (N_18480,N_17881,N_17762);
xnor U18481 (N_18481,N_17856,N_17628);
nand U18482 (N_18482,N_17802,N_17721);
xor U18483 (N_18483,N_17698,N_17997);
xor U18484 (N_18484,N_17910,N_17528);
nor U18485 (N_18485,N_17994,N_17537);
nor U18486 (N_18486,N_17823,N_17637);
xor U18487 (N_18487,N_17874,N_17823);
or U18488 (N_18488,N_17914,N_17875);
nand U18489 (N_18489,N_17855,N_17680);
or U18490 (N_18490,N_17584,N_17658);
nand U18491 (N_18491,N_17630,N_17600);
and U18492 (N_18492,N_17770,N_17901);
nand U18493 (N_18493,N_17623,N_17894);
nand U18494 (N_18494,N_17961,N_17752);
xnor U18495 (N_18495,N_17633,N_17940);
or U18496 (N_18496,N_17546,N_17996);
nand U18497 (N_18497,N_17772,N_17517);
and U18498 (N_18498,N_17992,N_17637);
nor U18499 (N_18499,N_17639,N_17910);
xor U18500 (N_18500,N_18185,N_18393);
or U18501 (N_18501,N_18139,N_18230);
or U18502 (N_18502,N_18465,N_18389);
and U18503 (N_18503,N_18032,N_18437);
and U18504 (N_18504,N_18205,N_18324);
and U18505 (N_18505,N_18189,N_18159);
nor U18506 (N_18506,N_18434,N_18143);
nor U18507 (N_18507,N_18246,N_18461);
xor U18508 (N_18508,N_18022,N_18038);
xnor U18509 (N_18509,N_18308,N_18336);
xnor U18510 (N_18510,N_18227,N_18470);
or U18511 (N_18511,N_18337,N_18449);
nor U18512 (N_18512,N_18242,N_18454);
or U18513 (N_18513,N_18366,N_18320);
or U18514 (N_18514,N_18484,N_18253);
nand U18515 (N_18515,N_18122,N_18099);
or U18516 (N_18516,N_18313,N_18131);
nand U18517 (N_18517,N_18216,N_18351);
or U18518 (N_18518,N_18284,N_18229);
nor U18519 (N_18519,N_18091,N_18068);
nor U18520 (N_18520,N_18098,N_18128);
and U18521 (N_18521,N_18160,N_18007);
xnor U18522 (N_18522,N_18417,N_18114);
nand U18523 (N_18523,N_18499,N_18400);
and U18524 (N_18524,N_18084,N_18238);
and U18525 (N_18525,N_18163,N_18476);
and U18526 (N_18526,N_18401,N_18208);
or U18527 (N_18527,N_18148,N_18441);
nand U18528 (N_18528,N_18309,N_18075);
xor U18529 (N_18529,N_18210,N_18149);
nand U18530 (N_18530,N_18096,N_18183);
xor U18531 (N_18531,N_18325,N_18270);
nand U18532 (N_18532,N_18363,N_18331);
and U18533 (N_18533,N_18169,N_18398);
and U18534 (N_18534,N_18219,N_18140);
or U18535 (N_18535,N_18279,N_18338);
nor U18536 (N_18536,N_18498,N_18150);
xnor U18537 (N_18537,N_18359,N_18002);
nor U18538 (N_18538,N_18080,N_18187);
xnor U18539 (N_18539,N_18251,N_18490);
nand U18540 (N_18540,N_18347,N_18373);
xnor U18541 (N_18541,N_18082,N_18374);
xor U18542 (N_18542,N_18370,N_18137);
or U18543 (N_18543,N_18263,N_18299);
and U18544 (N_18544,N_18358,N_18362);
or U18545 (N_18545,N_18327,N_18381);
nand U18546 (N_18546,N_18425,N_18066);
or U18547 (N_18547,N_18377,N_18415);
xor U18548 (N_18548,N_18047,N_18269);
xnor U18549 (N_18549,N_18110,N_18028);
xor U18550 (N_18550,N_18113,N_18217);
or U18551 (N_18551,N_18408,N_18092);
and U18552 (N_18552,N_18375,N_18481);
or U18553 (N_18553,N_18164,N_18412);
and U18554 (N_18554,N_18289,N_18201);
xnor U18555 (N_18555,N_18145,N_18474);
nor U18556 (N_18556,N_18345,N_18174);
and U18557 (N_18557,N_18192,N_18206);
nand U18558 (N_18558,N_18196,N_18103);
xor U18559 (N_18559,N_18466,N_18428);
or U18560 (N_18560,N_18414,N_18323);
nor U18561 (N_18561,N_18200,N_18477);
nand U18562 (N_18562,N_18019,N_18422);
nand U18563 (N_18563,N_18410,N_18211);
nand U18564 (N_18564,N_18121,N_18055);
or U18565 (N_18565,N_18054,N_18266);
nor U18566 (N_18566,N_18286,N_18011);
xnor U18567 (N_18567,N_18456,N_18440);
xnor U18568 (N_18568,N_18322,N_18235);
nor U18569 (N_18569,N_18218,N_18067);
nor U18570 (N_18570,N_18036,N_18407);
or U18571 (N_18571,N_18195,N_18492);
xor U18572 (N_18572,N_18280,N_18162);
or U18573 (N_18573,N_18353,N_18334);
xor U18574 (N_18574,N_18311,N_18072);
or U18575 (N_18575,N_18451,N_18316);
nor U18576 (N_18576,N_18435,N_18118);
nor U18577 (N_18577,N_18312,N_18129);
nor U18578 (N_18578,N_18302,N_18467);
and U18579 (N_18579,N_18404,N_18419);
nor U18580 (N_18580,N_18180,N_18307);
nor U18581 (N_18581,N_18109,N_18383);
or U18582 (N_18582,N_18221,N_18041);
xnor U18583 (N_18583,N_18016,N_18061);
xor U18584 (N_18584,N_18368,N_18436);
nor U18585 (N_18585,N_18391,N_18431);
nor U18586 (N_18586,N_18087,N_18170);
nand U18587 (N_18587,N_18273,N_18101);
and U18588 (N_18588,N_18457,N_18485);
nor U18589 (N_18589,N_18167,N_18491);
and U18590 (N_18590,N_18247,N_18267);
and U18591 (N_18591,N_18111,N_18259);
nor U18592 (N_18592,N_18369,N_18376);
xnor U18593 (N_18593,N_18287,N_18447);
and U18594 (N_18594,N_18010,N_18319);
and U18595 (N_18595,N_18379,N_18275);
xor U18596 (N_18596,N_18283,N_18315);
and U18597 (N_18597,N_18027,N_18257);
xnor U18598 (N_18598,N_18388,N_18146);
xnor U18599 (N_18599,N_18046,N_18105);
xnor U18600 (N_18600,N_18397,N_18380);
nand U18601 (N_18601,N_18459,N_18120);
xnor U18602 (N_18602,N_18236,N_18013);
nor U18603 (N_18603,N_18458,N_18144);
nand U18604 (N_18604,N_18117,N_18494);
xor U18605 (N_18605,N_18178,N_18086);
and U18606 (N_18606,N_18043,N_18329);
and U18607 (N_18607,N_18179,N_18088);
xnor U18608 (N_18608,N_18177,N_18475);
nor U18609 (N_18609,N_18278,N_18471);
nand U18610 (N_18610,N_18119,N_18126);
nand U18611 (N_18611,N_18173,N_18290);
nor U18612 (N_18612,N_18017,N_18240);
and U18613 (N_18613,N_18300,N_18095);
nor U18614 (N_18614,N_18361,N_18153);
and U18615 (N_18615,N_18424,N_18001);
nor U18616 (N_18616,N_18035,N_18395);
and U18617 (N_18617,N_18271,N_18489);
xnor U18618 (N_18618,N_18463,N_18332);
nor U18619 (N_18619,N_18448,N_18254);
nand U18620 (N_18620,N_18045,N_18059);
and U18621 (N_18621,N_18497,N_18051);
nor U18622 (N_18622,N_18250,N_18452);
nand U18623 (N_18623,N_18094,N_18202);
or U18624 (N_18624,N_18343,N_18024);
nand U18625 (N_18625,N_18314,N_18037);
xor U18626 (N_18626,N_18203,N_18194);
nor U18627 (N_18627,N_18232,N_18156);
or U18628 (N_18628,N_18468,N_18226);
or U18629 (N_18629,N_18065,N_18049);
or U18630 (N_18630,N_18292,N_18154);
and U18631 (N_18631,N_18244,N_18249);
xor U18632 (N_18632,N_18171,N_18346);
xor U18633 (N_18633,N_18107,N_18078);
and U18634 (N_18634,N_18100,N_18193);
nor U18635 (N_18635,N_18469,N_18060);
nor U18636 (N_18636,N_18062,N_18004);
nor U18637 (N_18637,N_18392,N_18135);
nand U18638 (N_18638,N_18303,N_18326);
and U18639 (N_18639,N_18089,N_18328);
and U18640 (N_18640,N_18453,N_18018);
nand U18641 (N_18641,N_18133,N_18209);
xor U18642 (N_18642,N_18382,N_18132);
or U18643 (N_18643,N_18029,N_18198);
xnor U18644 (N_18644,N_18394,N_18124);
nor U18645 (N_18645,N_18444,N_18237);
or U18646 (N_18646,N_18405,N_18384);
or U18647 (N_18647,N_18191,N_18277);
nor U18648 (N_18648,N_18473,N_18333);
nor U18649 (N_18649,N_18411,N_18360);
nor U18650 (N_18650,N_18233,N_18023);
xnor U18651 (N_18651,N_18090,N_18225);
nand U18652 (N_18652,N_18190,N_18335);
nor U18653 (N_18653,N_18288,N_18301);
nor U18654 (N_18654,N_18387,N_18070);
or U18655 (N_18655,N_18165,N_18125);
and U18656 (N_18656,N_18056,N_18228);
and U18657 (N_18657,N_18495,N_18040);
and U18658 (N_18658,N_18222,N_18188);
nor U18659 (N_18659,N_18108,N_18483);
or U18660 (N_18660,N_18081,N_18215);
xnor U18661 (N_18661,N_18239,N_18402);
or U18662 (N_18662,N_18462,N_18304);
nor U18663 (N_18663,N_18008,N_18420);
and U18664 (N_18664,N_18241,N_18293);
and U18665 (N_18665,N_18310,N_18012);
xnor U18666 (N_18666,N_18423,N_18472);
nor U18667 (N_18667,N_18265,N_18166);
xnor U18668 (N_18668,N_18450,N_18282);
nor U18669 (N_18669,N_18354,N_18429);
and U18670 (N_18670,N_18071,N_18030);
nand U18671 (N_18671,N_18357,N_18487);
and U18672 (N_18672,N_18268,N_18344);
or U18673 (N_18673,N_18378,N_18021);
nand U18674 (N_18674,N_18014,N_18147);
or U18675 (N_18675,N_18355,N_18298);
nor U18676 (N_18676,N_18260,N_18155);
nor U18677 (N_18677,N_18349,N_18482);
or U18678 (N_18678,N_18295,N_18341);
xnor U18679 (N_18679,N_18413,N_18294);
nand U18680 (N_18680,N_18199,N_18214);
xor U18681 (N_18681,N_18297,N_18409);
and U18682 (N_18682,N_18396,N_18076);
and U18683 (N_18683,N_18256,N_18116);
or U18684 (N_18684,N_18291,N_18057);
and U18685 (N_18685,N_18479,N_18158);
nor U18686 (N_18686,N_18430,N_18356);
xor U18687 (N_18687,N_18026,N_18073);
nand U18688 (N_18688,N_18127,N_18005);
or U18689 (N_18689,N_18339,N_18403);
nand U18690 (N_18690,N_18136,N_18340);
xor U18691 (N_18691,N_18033,N_18261);
xnor U18692 (N_18692,N_18318,N_18000);
xnor U18693 (N_18693,N_18063,N_18443);
or U18694 (N_18694,N_18406,N_18385);
nand U18695 (N_18695,N_18488,N_18034);
or U18696 (N_18696,N_18161,N_18115);
nor U18697 (N_18697,N_18274,N_18348);
xnor U18698 (N_18698,N_18305,N_18438);
or U18699 (N_18699,N_18031,N_18486);
or U18700 (N_18700,N_18258,N_18104);
nand U18701 (N_18701,N_18181,N_18248);
xor U18702 (N_18702,N_18234,N_18317);
and U18703 (N_18703,N_18455,N_18399);
nor U18704 (N_18704,N_18352,N_18064);
xnor U18705 (N_18705,N_18371,N_18386);
or U18706 (N_18706,N_18390,N_18464);
nor U18707 (N_18707,N_18069,N_18042);
nor U18708 (N_18708,N_18204,N_18478);
or U18709 (N_18709,N_18123,N_18151);
or U18710 (N_18710,N_18416,N_18015);
nand U18711 (N_18711,N_18281,N_18044);
nor U18712 (N_18712,N_18252,N_18460);
xor U18713 (N_18713,N_18321,N_18262);
or U18714 (N_18714,N_18142,N_18442);
xor U18715 (N_18715,N_18097,N_18048);
xnor U18716 (N_18716,N_18182,N_18223);
and U18717 (N_18717,N_18025,N_18009);
nand U18718 (N_18718,N_18446,N_18093);
and U18719 (N_18719,N_18134,N_18306);
or U18720 (N_18720,N_18168,N_18224);
nor U18721 (N_18721,N_18112,N_18493);
xnor U18722 (N_18722,N_18243,N_18050);
nor U18723 (N_18723,N_18052,N_18427);
nand U18724 (N_18724,N_18432,N_18276);
xor U18725 (N_18725,N_18426,N_18220);
nor U18726 (N_18726,N_18197,N_18285);
nor U18727 (N_18727,N_18058,N_18245);
nand U18728 (N_18728,N_18372,N_18433);
or U18729 (N_18729,N_18130,N_18106);
xnor U18730 (N_18730,N_18350,N_18083);
nor U18731 (N_18731,N_18365,N_18231);
and U18732 (N_18732,N_18138,N_18102);
nand U18733 (N_18733,N_18439,N_18421);
nor U18734 (N_18734,N_18186,N_18330);
nand U18735 (N_18735,N_18085,N_18039);
xor U18736 (N_18736,N_18213,N_18207);
nor U18737 (N_18737,N_18184,N_18296);
or U18738 (N_18738,N_18480,N_18157);
nor U18739 (N_18739,N_18141,N_18367);
or U18740 (N_18740,N_18077,N_18496);
xnor U18741 (N_18741,N_18074,N_18212);
and U18742 (N_18742,N_18175,N_18255);
or U18743 (N_18743,N_18079,N_18172);
xor U18744 (N_18744,N_18020,N_18053);
and U18745 (N_18745,N_18003,N_18264);
nand U18746 (N_18746,N_18272,N_18152);
and U18747 (N_18747,N_18342,N_18364);
xnor U18748 (N_18748,N_18418,N_18176);
xnor U18749 (N_18749,N_18445,N_18006);
or U18750 (N_18750,N_18266,N_18458);
or U18751 (N_18751,N_18268,N_18263);
nand U18752 (N_18752,N_18032,N_18326);
and U18753 (N_18753,N_18101,N_18097);
xnor U18754 (N_18754,N_18302,N_18323);
and U18755 (N_18755,N_18326,N_18273);
or U18756 (N_18756,N_18241,N_18348);
nor U18757 (N_18757,N_18478,N_18056);
and U18758 (N_18758,N_18455,N_18061);
or U18759 (N_18759,N_18234,N_18318);
nor U18760 (N_18760,N_18242,N_18069);
xnor U18761 (N_18761,N_18477,N_18489);
and U18762 (N_18762,N_18036,N_18210);
nor U18763 (N_18763,N_18469,N_18178);
and U18764 (N_18764,N_18061,N_18431);
nor U18765 (N_18765,N_18192,N_18382);
or U18766 (N_18766,N_18344,N_18212);
and U18767 (N_18767,N_18469,N_18429);
or U18768 (N_18768,N_18443,N_18071);
xnor U18769 (N_18769,N_18075,N_18293);
xnor U18770 (N_18770,N_18451,N_18485);
xor U18771 (N_18771,N_18239,N_18312);
and U18772 (N_18772,N_18472,N_18199);
and U18773 (N_18773,N_18163,N_18165);
or U18774 (N_18774,N_18023,N_18052);
xor U18775 (N_18775,N_18296,N_18148);
or U18776 (N_18776,N_18052,N_18315);
and U18777 (N_18777,N_18467,N_18171);
and U18778 (N_18778,N_18454,N_18105);
and U18779 (N_18779,N_18338,N_18225);
and U18780 (N_18780,N_18176,N_18455);
and U18781 (N_18781,N_18481,N_18438);
nor U18782 (N_18782,N_18444,N_18485);
or U18783 (N_18783,N_18371,N_18205);
nand U18784 (N_18784,N_18014,N_18248);
xnor U18785 (N_18785,N_18111,N_18485);
or U18786 (N_18786,N_18399,N_18259);
or U18787 (N_18787,N_18331,N_18400);
nor U18788 (N_18788,N_18169,N_18087);
nor U18789 (N_18789,N_18214,N_18321);
xor U18790 (N_18790,N_18021,N_18456);
nor U18791 (N_18791,N_18296,N_18159);
nor U18792 (N_18792,N_18124,N_18468);
nor U18793 (N_18793,N_18091,N_18389);
or U18794 (N_18794,N_18347,N_18064);
xor U18795 (N_18795,N_18294,N_18304);
and U18796 (N_18796,N_18382,N_18020);
nor U18797 (N_18797,N_18231,N_18095);
and U18798 (N_18798,N_18090,N_18449);
or U18799 (N_18799,N_18423,N_18021);
and U18800 (N_18800,N_18044,N_18447);
nand U18801 (N_18801,N_18293,N_18425);
xor U18802 (N_18802,N_18211,N_18475);
nor U18803 (N_18803,N_18153,N_18386);
xnor U18804 (N_18804,N_18323,N_18480);
and U18805 (N_18805,N_18084,N_18240);
nor U18806 (N_18806,N_18422,N_18161);
and U18807 (N_18807,N_18366,N_18152);
xor U18808 (N_18808,N_18405,N_18200);
nor U18809 (N_18809,N_18148,N_18220);
xor U18810 (N_18810,N_18240,N_18111);
nor U18811 (N_18811,N_18298,N_18037);
xor U18812 (N_18812,N_18026,N_18332);
xnor U18813 (N_18813,N_18358,N_18270);
nor U18814 (N_18814,N_18041,N_18496);
or U18815 (N_18815,N_18206,N_18072);
and U18816 (N_18816,N_18200,N_18373);
and U18817 (N_18817,N_18073,N_18409);
nand U18818 (N_18818,N_18036,N_18400);
nor U18819 (N_18819,N_18147,N_18125);
nand U18820 (N_18820,N_18192,N_18053);
and U18821 (N_18821,N_18186,N_18271);
xnor U18822 (N_18822,N_18293,N_18355);
nand U18823 (N_18823,N_18421,N_18313);
or U18824 (N_18824,N_18017,N_18214);
nand U18825 (N_18825,N_18322,N_18424);
or U18826 (N_18826,N_18239,N_18013);
and U18827 (N_18827,N_18361,N_18337);
or U18828 (N_18828,N_18023,N_18476);
nor U18829 (N_18829,N_18356,N_18436);
xnor U18830 (N_18830,N_18498,N_18366);
nand U18831 (N_18831,N_18030,N_18037);
nor U18832 (N_18832,N_18142,N_18022);
nand U18833 (N_18833,N_18331,N_18487);
or U18834 (N_18834,N_18419,N_18469);
or U18835 (N_18835,N_18390,N_18193);
nor U18836 (N_18836,N_18151,N_18446);
and U18837 (N_18837,N_18141,N_18189);
and U18838 (N_18838,N_18351,N_18261);
nor U18839 (N_18839,N_18012,N_18461);
xnor U18840 (N_18840,N_18214,N_18449);
or U18841 (N_18841,N_18452,N_18034);
xor U18842 (N_18842,N_18326,N_18411);
and U18843 (N_18843,N_18377,N_18003);
nor U18844 (N_18844,N_18157,N_18321);
xnor U18845 (N_18845,N_18061,N_18180);
nand U18846 (N_18846,N_18023,N_18257);
and U18847 (N_18847,N_18097,N_18376);
xor U18848 (N_18848,N_18388,N_18160);
nand U18849 (N_18849,N_18410,N_18261);
nor U18850 (N_18850,N_18484,N_18288);
xor U18851 (N_18851,N_18114,N_18274);
nand U18852 (N_18852,N_18042,N_18220);
xor U18853 (N_18853,N_18272,N_18353);
nor U18854 (N_18854,N_18051,N_18371);
nor U18855 (N_18855,N_18347,N_18145);
or U18856 (N_18856,N_18254,N_18078);
xnor U18857 (N_18857,N_18461,N_18295);
nand U18858 (N_18858,N_18045,N_18426);
and U18859 (N_18859,N_18470,N_18499);
and U18860 (N_18860,N_18460,N_18432);
and U18861 (N_18861,N_18290,N_18380);
nand U18862 (N_18862,N_18304,N_18165);
or U18863 (N_18863,N_18037,N_18276);
and U18864 (N_18864,N_18268,N_18055);
nand U18865 (N_18865,N_18370,N_18131);
xnor U18866 (N_18866,N_18343,N_18112);
and U18867 (N_18867,N_18447,N_18426);
nor U18868 (N_18868,N_18470,N_18356);
xnor U18869 (N_18869,N_18025,N_18358);
and U18870 (N_18870,N_18420,N_18088);
xor U18871 (N_18871,N_18328,N_18264);
xnor U18872 (N_18872,N_18224,N_18056);
xnor U18873 (N_18873,N_18137,N_18187);
xnor U18874 (N_18874,N_18297,N_18333);
or U18875 (N_18875,N_18179,N_18174);
xor U18876 (N_18876,N_18072,N_18151);
or U18877 (N_18877,N_18082,N_18490);
and U18878 (N_18878,N_18021,N_18089);
nor U18879 (N_18879,N_18109,N_18353);
and U18880 (N_18880,N_18106,N_18082);
xor U18881 (N_18881,N_18216,N_18317);
nand U18882 (N_18882,N_18026,N_18316);
and U18883 (N_18883,N_18299,N_18453);
xor U18884 (N_18884,N_18184,N_18316);
nand U18885 (N_18885,N_18161,N_18037);
and U18886 (N_18886,N_18099,N_18232);
and U18887 (N_18887,N_18270,N_18142);
or U18888 (N_18888,N_18372,N_18252);
and U18889 (N_18889,N_18005,N_18320);
or U18890 (N_18890,N_18327,N_18203);
xor U18891 (N_18891,N_18307,N_18467);
or U18892 (N_18892,N_18279,N_18029);
or U18893 (N_18893,N_18197,N_18124);
and U18894 (N_18894,N_18310,N_18185);
nor U18895 (N_18895,N_18169,N_18224);
or U18896 (N_18896,N_18453,N_18424);
or U18897 (N_18897,N_18000,N_18338);
nor U18898 (N_18898,N_18263,N_18101);
xor U18899 (N_18899,N_18345,N_18299);
xnor U18900 (N_18900,N_18466,N_18160);
nand U18901 (N_18901,N_18081,N_18197);
and U18902 (N_18902,N_18343,N_18007);
nand U18903 (N_18903,N_18046,N_18298);
and U18904 (N_18904,N_18079,N_18303);
or U18905 (N_18905,N_18476,N_18469);
nand U18906 (N_18906,N_18385,N_18276);
xor U18907 (N_18907,N_18393,N_18414);
nor U18908 (N_18908,N_18251,N_18212);
or U18909 (N_18909,N_18119,N_18195);
nor U18910 (N_18910,N_18295,N_18288);
and U18911 (N_18911,N_18087,N_18335);
or U18912 (N_18912,N_18235,N_18340);
nor U18913 (N_18913,N_18185,N_18486);
or U18914 (N_18914,N_18278,N_18341);
or U18915 (N_18915,N_18132,N_18363);
or U18916 (N_18916,N_18103,N_18311);
nor U18917 (N_18917,N_18370,N_18326);
nand U18918 (N_18918,N_18406,N_18062);
or U18919 (N_18919,N_18484,N_18416);
nand U18920 (N_18920,N_18353,N_18186);
or U18921 (N_18921,N_18438,N_18155);
or U18922 (N_18922,N_18423,N_18149);
or U18923 (N_18923,N_18259,N_18172);
and U18924 (N_18924,N_18193,N_18048);
and U18925 (N_18925,N_18344,N_18048);
nand U18926 (N_18926,N_18113,N_18266);
xor U18927 (N_18927,N_18483,N_18462);
xor U18928 (N_18928,N_18158,N_18311);
or U18929 (N_18929,N_18311,N_18297);
nand U18930 (N_18930,N_18461,N_18191);
xnor U18931 (N_18931,N_18424,N_18179);
nor U18932 (N_18932,N_18080,N_18102);
and U18933 (N_18933,N_18356,N_18361);
xnor U18934 (N_18934,N_18012,N_18047);
nand U18935 (N_18935,N_18190,N_18312);
and U18936 (N_18936,N_18229,N_18459);
nand U18937 (N_18937,N_18397,N_18019);
xnor U18938 (N_18938,N_18092,N_18266);
xnor U18939 (N_18939,N_18113,N_18442);
and U18940 (N_18940,N_18479,N_18077);
and U18941 (N_18941,N_18481,N_18376);
nor U18942 (N_18942,N_18147,N_18130);
and U18943 (N_18943,N_18237,N_18265);
nor U18944 (N_18944,N_18111,N_18193);
nor U18945 (N_18945,N_18117,N_18111);
xor U18946 (N_18946,N_18286,N_18166);
xor U18947 (N_18947,N_18109,N_18258);
and U18948 (N_18948,N_18182,N_18128);
and U18949 (N_18949,N_18447,N_18385);
and U18950 (N_18950,N_18066,N_18064);
nand U18951 (N_18951,N_18335,N_18395);
or U18952 (N_18952,N_18266,N_18143);
nand U18953 (N_18953,N_18193,N_18222);
and U18954 (N_18954,N_18416,N_18186);
xor U18955 (N_18955,N_18273,N_18160);
xnor U18956 (N_18956,N_18354,N_18100);
and U18957 (N_18957,N_18037,N_18418);
or U18958 (N_18958,N_18432,N_18338);
or U18959 (N_18959,N_18268,N_18085);
xnor U18960 (N_18960,N_18067,N_18340);
nor U18961 (N_18961,N_18492,N_18407);
nor U18962 (N_18962,N_18212,N_18061);
nor U18963 (N_18963,N_18215,N_18166);
and U18964 (N_18964,N_18176,N_18020);
and U18965 (N_18965,N_18470,N_18204);
nor U18966 (N_18966,N_18413,N_18225);
or U18967 (N_18967,N_18046,N_18125);
or U18968 (N_18968,N_18241,N_18390);
and U18969 (N_18969,N_18307,N_18092);
and U18970 (N_18970,N_18280,N_18383);
and U18971 (N_18971,N_18326,N_18399);
nor U18972 (N_18972,N_18231,N_18367);
and U18973 (N_18973,N_18340,N_18266);
nor U18974 (N_18974,N_18430,N_18061);
nand U18975 (N_18975,N_18499,N_18322);
nor U18976 (N_18976,N_18134,N_18152);
nand U18977 (N_18977,N_18169,N_18080);
and U18978 (N_18978,N_18077,N_18106);
or U18979 (N_18979,N_18278,N_18440);
or U18980 (N_18980,N_18017,N_18409);
xor U18981 (N_18981,N_18209,N_18182);
xnor U18982 (N_18982,N_18252,N_18354);
nand U18983 (N_18983,N_18068,N_18249);
nor U18984 (N_18984,N_18295,N_18040);
nand U18985 (N_18985,N_18399,N_18070);
nand U18986 (N_18986,N_18136,N_18283);
xor U18987 (N_18987,N_18127,N_18067);
nor U18988 (N_18988,N_18435,N_18041);
nor U18989 (N_18989,N_18450,N_18123);
nor U18990 (N_18990,N_18414,N_18145);
nand U18991 (N_18991,N_18038,N_18114);
nand U18992 (N_18992,N_18347,N_18487);
xor U18993 (N_18993,N_18013,N_18041);
xor U18994 (N_18994,N_18488,N_18450);
and U18995 (N_18995,N_18443,N_18089);
or U18996 (N_18996,N_18092,N_18004);
nand U18997 (N_18997,N_18061,N_18334);
and U18998 (N_18998,N_18241,N_18369);
and U18999 (N_18999,N_18262,N_18082);
or U19000 (N_19000,N_18576,N_18710);
nor U19001 (N_19001,N_18997,N_18791);
nand U19002 (N_19002,N_18998,N_18583);
nand U19003 (N_19003,N_18915,N_18613);
xor U19004 (N_19004,N_18758,N_18502);
xnor U19005 (N_19005,N_18985,N_18850);
xnor U19006 (N_19006,N_18786,N_18578);
and U19007 (N_19007,N_18925,N_18674);
or U19008 (N_19008,N_18824,N_18881);
xor U19009 (N_19009,N_18887,N_18618);
and U19010 (N_19010,N_18923,N_18875);
xnor U19011 (N_19011,N_18784,N_18785);
nand U19012 (N_19012,N_18564,N_18837);
xor U19013 (N_19013,N_18566,N_18862);
xnor U19014 (N_19014,N_18794,N_18760);
or U19015 (N_19015,N_18528,N_18619);
or U19016 (N_19016,N_18606,N_18677);
nor U19017 (N_19017,N_18901,N_18680);
nand U19018 (N_19018,N_18732,N_18649);
xnor U19019 (N_19019,N_18695,N_18951);
or U19020 (N_19020,N_18724,N_18937);
and U19021 (N_19021,N_18535,N_18888);
or U19022 (N_19022,N_18776,N_18857);
nand U19023 (N_19023,N_18636,N_18629);
or U19024 (N_19024,N_18505,N_18729);
or U19025 (N_19025,N_18867,N_18775);
and U19026 (N_19026,N_18828,N_18879);
or U19027 (N_19027,N_18911,N_18814);
xnor U19028 (N_19028,N_18548,N_18627);
nor U19029 (N_19029,N_18598,N_18694);
and U19030 (N_19030,N_18831,N_18780);
or U19031 (N_19031,N_18861,N_18610);
nor U19032 (N_19032,N_18543,N_18733);
nand U19033 (N_19033,N_18756,N_18631);
nor U19034 (N_19034,N_18704,N_18999);
nand U19035 (N_19035,N_18500,N_18616);
or U19036 (N_19036,N_18928,N_18759);
xor U19037 (N_19037,N_18736,N_18565);
and U19038 (N_19038,N_18559,N_18774);
and U19039 (N_19039,N_18897,N_18910);
or U19040 (N_19040,N_18839,N_18864);
nor U19041 (N_19041,N_18676,N_18844);
or U19042 (N_19042,N_18660,N_18795);
xnor U19043 (N_19043,N_18555,N_18821);
and U19044 (N_19044,N_18642,N_18983);
nand U19045 (N_19045,N_18843,N_18971);
nor U19046 (N_19046,N_18949,N_18718);
nand U19047 (N_19047,N_18917,N_18707);
and U19048 (N_19048,N_18700,N_18580);
xnor U19049 (N_19049,N_18865,N_18682);
or U19050 (N_19050,N_18913,N_18653);
nor U19051 (N_19051,N_18830,N_18777);
xor U19052 (N_19052,N_18863,N_18966);
xnor U19053 (N_19053,N_18815,N_18907);
xnor U19054 (N_19054,N_18972,N_18800);
xnor U19055 (N_19055,N_18894,N_18670);
nor U19056 (N_19056,N_18932,N_18679);
xnor U19057 (N_19057,N_18571,N_18833);
or U19058 (N_19058,N_18793,N_18572);
or U19059 (N_19059,N_18961,N_18939);
or U19060 (N_19060,N_18628,N_18678);
nand U19061 (N_19061,N_18841,N_18518);
or U19062 (N_19062,N_18902,N_18904);
and U19063 (N_19063,N_18757,N_18820);
xnor U19064 (N_19064,N_18720,N_18770);
xor U19065 (N_19065,N_18715,N_18573);
or U19066 (N_19066,N_18935,N_18582);
xnor U19067 (N_19067,N_18974,N_18990);
nor U19068 (N_19068,N_18506,N_18866);
and U19069 (N_19069,N_18955,N_18803);
and U19070 (N_19070,N_18727,N_18798);
xnor U19071 (N_19071,N_18664,N_18731);
xnor U19072 (N_19072,N_18943,N_18801);
or U19073 (N_19073,N_18809,N_18845);
xor U19074 (N_19074,N_18507,N_18751);
nor U19075 (N_19075,N_18623,N_18714);
nor U19076 (N_19076,N_18813,N_18931);
or U19077 (N_19077,N_18953,N_18644);
nand U19078 (N_19078,N_18970,N_18869);
nand U19079 (N_19079,N_18764,N_18877);
xnor U19080 (N_19080,N_18878,N_18895);
nor U19081 (N_19081,N_18773,N_18744);
and U19082 (N_19082,N_18522,N_18659);
xnor U19083 (N_19083,N_18551,N_18818);
and U19084 (N_19084,N_18969,N_18842);
xnor U19085 (N_19085,N_18789,N_18602);
or U19086 (N_19086,N_18908,N_18635);
nand U19087 (N_19087,N_18790,N_18730);
and U19088 (N_19088,N_18728,N_18717);
or U19089 (N_19089,N_18766,N_18920);
nor U19090 (N_19090,N_18554,N_18747);
and U19091 (N_19091,N_18981,N_18647);
or U19092 (N_19092,N_18827,N_18600);
or U19093 (N_19093,N_18944,N_18782);
nand U19094 (N_19094,N_18698,N_18889);
nor U19095 (N_19095,N_18745,N_18640);
and U19096 (N_19096,N_18769,N_18652);
or U19097 (N_19097,N_18504,N_18846);
xor U19098 (N_19098,N_18550,N_18662);
nor U19099 (N_19099,N_18805,N_18542);
or U19100 (N_19100,N_18614,N_18853);
nand U19101 (N_19101,N_18787,N_18632);
or U19102 (N_19102,N_18592,N_18586);
nand U19103 (N_19103,N_18609,N_18595);
nor U19104 (N_19104,N_18952,N_18557);
nor U19105 (N_19105,N_18980,N_18826);
nor U19106 (N_19106,N_18617,N_18658);
nor U19107 (N_19107,N_18549,N_18856);
xor U19108 (N_19108,N_18840,N_18964);
xnor U19109 (N_19109,N_18611,N_18941);
xnor U19110 (N_19110,N_18989,N_18692);
nand U19111 (N_19111,N_18763,N_18924);
nor U19112 (N_19112,N_18973,N_18533);
nor U19113 (N_19113,N_18979,N_18643);
and U19114 (N_19114,N_18712,N_18544);
nor U19115 (N_19115,N_18645,N_18574);
xnor U19116 (N_19116,N_18577,N_18581);
nand U19117 (N_19117,N_18591,N_18906);
nor U19118 (N_19118,N_18936,N_18933);
xor U19119 (N_19119,N_18510,N_18772);
xor U19120 (N_19120,N_18858,N_18752);
nand U19121 (N_19121,N_18958,N_18768);
nand U19122 (N_19122,N_18948,N_18596);
nor U19123 (N_19123,N_18537,N_18739);
xor U19124 (N_19124,N_18625,N_18553);
and U19125 (N_19125,N_18651,N_18806);
xnor U19126 (N_19126,N_18512,N_18967);
nor U19127 (N_19127,N_18575,N_18713);
and U19128 (N_19128,N_18854,N_18956);
and U19129 (N_19129,N_18808,N_18668);
or U19130 (N_19130,N_18994,N_18959);
xor U19131 (N_19131,N_18532,N_18716);
nand U19132 (N_19132,N_18799,N_18527);
xor U19133 (N_19133,N_18918,N_18657);
or U19134 (N_19134,N_18876,N_18562);
or U19135 (N_19135,N_18886,N_18517);
nand U19136 (N_19136,N_18579,N_18940);
and U19137 (N_19137,N_18835,N_18634);
or U19138 (N_19138,N_18539,N_18742);
nand U19139 (N_19139,N_18802,N_18987);
nand U19140 (N_19140,N_18765,N_18811);
or U19141 (N_19141,N_18741,N_18546);
xnor U19142 (N_19142,N_18706,N_18882);
nand U19143 (N_19143,N_18673,N_18992);
or U19144 (N_19144,N_18639,N_18892);
nor U19145 (N_19145,N_18822,N_18991);
or U19146 (N_19146,N_18558,N_18515);
or U19147 (N_19147,N_18519,N_18514);
or U19148 (N_19148,N_18501,N_18666);
nor U19149 (N_19149,N_18738,N_18708);
or U19150 (N_19150,N_18750,N_18912);
nor U19151 (N_19151,N_18691,N_18900);
nor U19152 (N_19152,N_18965,N_18667);
xnor U19153 (N_19153,N_18737,N_18870);
or U19154 (N_19154,N_18624,N_18860);
xor U19155 (N_19155,N_18536,N_18905);
or U19156 (N_19156,N_18511,N_18753);
nor U19157 (N_19157,N_18597,N_18584);
nand U19158 (N_19158,N_18899,N_18977);
or U19159 (N_19159,N_18589,N_18561);
or U19160 (N_19160,N_18819,N_18656);
nor U19161 (N_19161,N_18817,N_18761);
nand U19162 (N_19162,N_18848,N_18754);
nand U19163 (N_19163,N_18690,N_18547);
xnor U19164 (N_19164,N_18671,N_18693);
or U19165 (N_19165,N_18622,N_18612);
nand U19166 (N_19166,N_18962,N_18723);
nand U19167 (N_19167,N_18783,N_18823);
nand U19168 (N_19168,N_18705,N_18567);
nor U19169 (N_19169,N_18563,N_18930);
or U19170 (N_19170,N_18748,N_18946);
and U19171 (N_19171,N_18540,N_18909);
nand U19172 (N_19172,N_18688,N_18755);
nand U19173 (N_19173,N_18681,N_18655);
xor U19174 (N_19174,N_18697,N_18781);
or U19175 (N_19175,N_18641,N_18880);
nor U19176 (N_19176,N_18725,N_18792);
and U19177 (N_19177,N_18740,N_18588);
or U19178 (N_19178,N_18702,N_18829);
and U19179 (N_19179,N_18638,N_18749);
nand U19180 (N_19180,N_18885,N_18849);
xor U19181 (N_19181,N_18891,N_18903);
nor U19182 (N_19182,N_18927,N_18868);
and U19183 (N_19183,N_18838,N_18804);
and U19184 (N_19184,N_18734,N_18986);
nor U19185 (N_19185,N_18855,N_18921);
nand U19186 (N_19186,N_18778,N_18834);
xnor U19187 (N_19187,N_18529,N_18685);
or U19188 (N_19188,N_18509,N_18569);
and U19189 (N_19189,N_18599,N_18711);
and U19190 (N_19190,N_18703,N_18916);
or U19191 (N_19191,N_18534,N_18545);
and U19192 (N_19192,N_18978,N_18984);
nor U19193 (N_19193,N_18661,N_18663);
and U19194 (N_19194,N_18648,N_18767);
nor U19195 (N_19195,N_18556,N_18746);
or U19196 (N_19196,N_18995,N_18701);
or U19197 (N_19197,N_18513,N_18669);
or U19198 (N_19198,N_18689,N_18893);
or U19199 (N_19199,N_18552,N_18568);
nand U19200 (N_19200,N_18807,N_18859);
or U19201 (N_19201,N_18968,N_18630);
xnor U19202 (N_19202,N_18779,N_18926);
and U19203 (N_19203,N_18947,N_18621);
xnor U19204 (N_19204,N_18996,N_18594);
nand U19205 (N_19205,N_18637,N_18722);
nand U19206 (N_19206,N_18883,N_18988);
and U19207 (N_19207,N_18873,N_18520);
or U19208 (N_19208,N_18922,N_18560);
nand U19209 (N_19209,N_18654,N_18684);
nand U19210 (N_19210,N_18735,N_18696);
nor U19211 (N_19211,N_18646,N_18872);
xnor U19212 (N_19212,N_18603,N_18508);
xnor U19213 (N_19213,N_18538,N_18871);
and U19214 (N_19214,N_18743,N_18797);
xor U19215 (N_19215,N_18650,N_18709);
nand U19216 (N_19216,N_18851,N_18929);
or U19217 (N_19217,N_18525,N_18963);
nor U19218 (N_19218,N_18687,N_18950);
and U19219 (N_19219,N_18605,N_18541);
and U19220 (N_19220,N_18608,N_18523);
xor U19221 (N_19221,N_18590,N_18812);
and U19222 (N_19222,N_18852,N_18607);
nand U19223 (N_19223,N_18976,N_18810);
or U19224 (N_19224,N_18516,N_18593);
or U19225 (N_19225,N_18699,N_18816);
nand U19226 (N_19226,N_18771,N_18530);
nand U19227 (N_19227,N_18726,N_18954);
xor U19228 (N_19228,N_18604,N_18665);
nand U19229 (N_19229,N_18982,N_18531);
or U19230 (N_19230,N_18683,N_18686);
xnor U19231 (N_19231,N_18633,N_18874);
xnor U19232 (N_19232,N_18914,N_18898);
and U19233 (N_19233,N_18719,N_18884);
or U19234 (N_19234,N_18615,N_18890);
nand U19235 (N_19235,N_18934,N_18524);
nand U19236 (N_19236,N_18896,N_18585);
xor U19237 (N_19237,N_18919,N_18762);
nor U19238 (N_19238,N_18620,N_18836);
xnor U19239 (N_19239,N_18825,N_18847);
nand U19240 (N_19240,N_18796,N_18788);
xor U19241 (N_19241,N_18521,N_18938);
nor U19242 (N_19242,N_18721,N_18832);
nor U19243 (N_19243,N_18570,N_18957);
and U19244 (N_19244,N_18993,N_18945);
nor U19245 (N_19245,N_18503,N_18601);
or U19246 (N_19246,N_18672,N_18587);
and U19247 (N_19247,N_18526,N_18975);
and U19248 (N_19248,N_18942,N_18960);
or U19249 (N_19249,N_18675,N_18626);
nor U19250 (N_19250,N_18582,N_18811);
or U19251 (N_19251,N_18684,N_18603);
or U19252 (N_19252,N_18861,N_18764);
or U19253 (N_19253,N_18771,N_18952);
and U19254 (N_19254,N_18854,N_18778);
and U19255 (N_19255,N_18767,N_18625);
or U19256 (N_19256,N_18510,N_18797);
and U19257 (N_19257,N_18652,N_18802);
or U19258 (N_19258,N_18870,N_18577);
or U19259 (N_19259,N_18702,N_18630);
nor U19260 (N_19260,N_18725,N_18846);
or U19261 (N_19261,N_18778,N_18926);
nand U19262 (N_19262,N_18843,N_18557);
and U19263 (N_19263,N_18682,N_18804);
nor U19264 (N_19264,N_18649,N_18507);
or U19265 (N_19265,N_18815,N_18582);
nor U19266 (N_19266,N_18768,N_18556);
and U19267 (N_19267,N_18696,N_18719);
nand U19268 (N_19268,N_18834,N_18805);
or U19269 (N_19269,N_18993,N_18871);
nor U19270 (N_19270,N_18964,N_18812);
nor U19271 (N_19271,N_18581,N_18944);
nand U19272 (N_19272,N_18656,N_18543);
nor U19273 (N_19273,N_18991,N_18778);
or U19274 (N_19274,N_18614,N_18524);
xor U19275 (N_19275,N_18918,N_18577);
and U19276 (N_19276,N_18778,N_18754);
nand U19277 (N_19277,N_18868,N_18658);
xor U19278 (N_19278,N_18591,N_18984);
or U19279 (N_19279,N_18960,N_18635);
nor U19280 (N_19280,N_18907,N_18533);
or U19281 (N_19281,N_18934,N_18812);
and U19282 (N_19282,N_18771,N_18646);
and U19283 (N_19283,N_18730,N_18733);
nor U19284 (N_19284,N_18647,N_18678);
nor U19285 (N_19285,N_18854,N_18732);
and U19286 (N_19286,N_18552,N_18798);
xnor U19287 (N_19287,N_18777,N_18626);
nor U19288 (N_19288,N_18700,N_18766);
or U19289 (N_19289,N_18957,N_18789);
nor U19290 (N_19290,N_18753,N_18776);
xor U19291 (N_19291,N_18763,N_18772);
xor U19292 (N_19292,N_18975,N_18694);
and U19293 (N_19293,N_18907,N_18765);
nor U19294 (N_19294,N_18611,N_18610);
nand U19295 (N_19295,N_18873,N_18917);
xnor U19296 (N_19296,N_18641,N_18992);
nor U19297 (N_19297,N_18563,N_18765);
or U19298 (N_19298,N_18988,N_18641);
or U19299 (N_19299,N_18874,N_18655);
xor U19300 (N_19300,N_18954,N_18573);
nand U19301 (N_19301,N_18630,N_18576);
and U19302 (N_19302,N_18982,N_18942);
nand U19303 (N_19303,N_18502,N_18576);
or U19304 (N_19304,N_18870,N_18588);
and U19305 (N_19305,N_18901,N_18906);
or U19306 (N_19306,N_18524,N_18829);
xnor U19307 (N_19307,N_18797,N_18683);
nor U19308 (N_19308,N_18588,N_18878);
and U19309 (N_19309,N_18968,N_18923);
nand U19310 (N_19310,N_18696,N_18894);
nand U19311 (N_19311,N_18887,N_18765);
or U19312 (N_19312,N_18917,N_18916);
nor U19313 (N_19313,N_18902,N_18765);
nand U19314 (N_19314,N_18856,N_18506);
xor U19315 (N_19315,N_18526,N_18926);
xnor U19316 (N_19316,N_18631,N_18933);
xnor U19317 (N_19317,N_18821,N_18838);
nand U19318 (N_19318,N_18732,N_18562);
and U19319 (N_19319,N_18511,N_18712);
and U19320 (N_19320,N_18744,N_18866);
nor U19321 (N_19321,N_18701,N_18507);
or U19322 (N_19322,N_18773,N_18565);
nor U19323 (N_19323,N_18539,N_18793);
nand U19324 (N_19324,N_18533,N_18557);
and U19325 (N_19325,N_18984,N_18727);
xor U19326 (N_19326,N_18715,N_18686);
nor U19327 (N_19327,N_18679,N_18705);
and U19328 (N_19328,N_18918,N_18864);
and U19329 (N_19329,N_18769,N_18559);
xnor U19330 (N_19330,N_18904,N_18532);
and U19331 (N_19331,N_18995,N_18653);
nor U19332 (N_19332,N_18965,N_18684);
or U19333 (N_19333,N_18714,N_18663);
nor U19334 (N_19334,N_18982,N_18851);
xor U19335 (N_19335,N_18756,N_18736);
or U19336 (N_19336,N_18778,N_18501);
or U19337 (N_19337,N_18952,N_18592);
and U19338 (N_19338,N_18816,N_18515);
nand U19339 (N_19339,N_18888,N_18829);
and U19340 (N_19340,N_18660,N_18692);
nand U19341 (N_19341,N_18632,N_18515);
or U19342 (N_19342,N_18673,N_18564);
nor U19343 (N_19343,N_18766,N_18889);
nor U19344 (N_19344,N_18913,N_18656);
nand U19345 (N_19345,N_18713,N_18848);
nor U19346 (N_19346,N_18736,N_18958);
or U19347 (N_19347,N_18529,N_18864);
or U19348 (N_19348,N_18949,N_18827);
xor U19349 (N_19349,N_18857,N_18915);
nor U19350 (N_19350,N_18596,N_18749);
nor U19351 (N_19351,N_18891,N_18921);
nand U19352 (N_19352,N_18899,N_18886);
nor U19353 (N_19353,N_18711,N_18829);
or U19354 (N_19354,N_18971,N_18970);
nor U19355 (N_19355,N_18645,N_18913);
nor U19356 (N_19356,N_18992,N_18630);
or U19357 (N_19357,N_18797,N_18705);
and U19358 (N_19358,N_18870,N_18914);
and U19359 (N_19359,N_18924,N_18868);
nor U19360 (N_19360,N_18661,N_18815);
nand U19361 (N_19361,N_18966,N_18684);
and U19362 (N_19362,N_18791,N_18824);
and U19363 (N_19363,N_18753,N_18612);
xnor U19364 (N_19364,N_18952,N_18733);
nand U19365 (N_19365,N_18959,N_18887);
or U19366 (N_19366,N_18900,N_18895);
nor U19367 (N_19367,N_18687,N_18603);
nor U19368 (N_19368,N_18504,N_18619);
nand U19369 (N_19369,N_18858,N_18845);
nor U19370 (N_19370,N_18927,N_18975);
and U19371 (N_19371,N_18620,N_18968);
or U19372 (N_19372,N_18831,N_18613);
xnor U19373 (N_19373,N_18744,N_18721);
nor U19374 (N_19374,N_18769,N_18843);
or U19375 (N_19375,N_18584,N_18675);
nor U19376 (N_19376,N_18582,N_18519);
or U19377 (N_19377,N_18657,N_18715);
or U19378 (N_19378,N_18730,N_18879);
nand U19379 (N_19379,N_18989,N_18951);
nand U19380 (N_19380,N_18703,N_18569);
nor U19381 (N_19381,N_18800,N_18731);
nand U19382 (N_19382,N_18993,N_18759);
nor U19383 (N_19383,N_18844,N_18857);
and U19384 (N_19384,N_18750,N_18677);
xnor U19385 (N_19385,N_18678,N_18780);
and U19386 (N_19386,N_18991,N_18558);
nand U19387 (N_19387,N_18780,N_18749);
and U19388 (N_19388,N_18582,N_18769);
nand U19389 (N_19389,N_18591,N_18794);
xnor U19390 (N_19390,N_18533,N_18673);
nor U19391 (N_19391,N_18981,N_18823);
or U19392 (N_19392,N_18667,N_18814);
nor U19393 (N_19393,N_18922,N_18550);
nand U19394 (N_19394,N_18813,N_18638);
or U19395 (N_19395,N_18780,N_18631);
nand U19396 (N_19396,N_18504,N_18550);
nand U19397 (N_19397,N_18677,N_18716);
or U19398 (N_19398,N_18787,N_18610);
and U19399 (N_19399,N_18532,N_18753);
nor U19400 (N_19400,N_18627,N_18756);
or U19401 (N_19401,N_18911,N_18710);
xnor U19402 (N_19402,N_18735,N_18648);
and U19403 (N_19403,N_18824,N_18776);
nor U19404 (N_19404,N_18722,N_18696);
nor U19405 (N_19405,N_18538,N_18988);
and U19406 (N_19406,N_18789,N_18935);
nor U19407 (N_19407,N_18517,N_18504);
nor U19408 (N_19408,N_18862,N_18702);
or U19409 (N_19409,N_18857,N_18624);
xor U19410 (N_19410,N_18861,N_18691);
or U19411 (N_19411,N_18943,N_18969);
nor U19412 (N_19412,N_18599,N_18825);
or U19413 (N_19413,N_18959,N_18681);
nor U19414 (N_19414,N_18871,N_18650);
xor U19415 (N_19415,N_18749,N_18841);
xor U19416 (N_19416,N_18741,N_18651);
and U19417 (N_19417,N_18976,N_18600);
xnor U19418 (N_19418,N_18919,N_18835);
xnor U19419 (N_19419,N_18780,N_18924);
and U19420 (N_19420,N_18715,N_18737);
or U19421 (N_19421,N_18789,N_18509);
nand U19422 (N_19422,N_18659,N_18538);
nor U19423 (N_19423,N_18758,N_18816);
xnor U19424 (N_19424,N_18928,N_18729);
nand U19425 (N_19425,N_18665,N_18853);
or U19426 (N_19426,N_18535,N_18797);
xnor U19427 (N_19427,N_18907,N_18545);
and U19428 (N_19428,N_18826,N_18549);
nand U19429 (N_19429,N_18733,N_18613);
and U19430 (N_19430,N_18988,N_18629);
xnor U19431 (N_19431,N_18686,N_18947);
nor U19432 (N_19432,N_18650,N_18830);
or U19433 (N_19433,N_18529,N_18649);
nor U19434 (N_19434,N_18653,N_18697);
nand U19435 (N_19435,N_18753,N_18601);
nor U19436 (N_19436,N_18642,N_18871);
nand U19437 (N_19437,N_18618,N_18932);
or U19438 (N_19438,N_18784,N_18583);
nor U19439 (N_19439,N_18753,N_18735);
or U19440 (N_19440,N_18708,N_18847);
or U19441 (N_19441,N_18664,N_18951);
nor U19442 (N_19442,N_18941,N_18717);
nand U19443 (N_19443,N_18953,N_18957);
nand U19444 (N_19444,N_18666,N_18943);
nand U19445 (N_19445,N_18987,N_18796);
and U19446 (N_19446,N_18643,N_18578);
xor U19447 (N_19447,N_18592,N_18895);
xnor U19448 (N_19448,N_18801,N_18873);
and U19449 (N_19449,N_18834,N_18789);
and U19450 (N_19450,N_18503,N_18556);
xor U19451 (N_19451,N_18537,N_18969);
nand U19452 (N_19452,N_18590,N_18974);
xor U19453 (N_19453,N_18555,N_18946);
xor U19454 (N_19454,N_18992,N_18681);
or U19455 (N_19455,N_18590,N_18655);
nand U19456 (N_19456,N_18649,N_18915);
xnor U19457 (N_19457,N_18792,N_18846);
nand U19458 (N_19458,N_18833,N_18864);
nor U19459 (N_19459,N_18534,N_18644);
and U19460 (N_19460,N_18717,N_18854);
or U19461 (N_19461,N_18736,N_18690);
nand U19462 (N_19462,N_18736,N_18868);
and U19463 (N_19463,N_18945,N_18766);
xor U19464 (N_19464,N_18925,N_18616);
and U19465 (N_19465,N_18933,N_18672);
xnor U19466 (N_19466,N_18542,N_18760);
nor U19467 (N_19467,N_18573,N_18541);
or U19468 (N_19468,N_18919,N_18908);
xor U19469 (N_19469,N_18608,N_18940);
and U19470 (N_19470,N_18813,N_18814);
and U19471 (N_19471,N_18719,N_18674);
nand U19472 (N_19472,N_18917,N_18797);
nand U19473 (N_19473,N_18597,N_18827);
xnor U19474 (N_19474,N_18936,N_18554);
or U19475 (N_19475,N_18706,N_18605);
xnor U19476 (N_19476,N_18773,N_18537);
xor U19477 (N_19477,N_18885,N_18754);
nor U19478 (N_19478,N_18563,N_18986);
nand U19479 (N_19479,N_18913,N_18748);
or U19480 (N_19480,N_18593,N_18770);
xnor U19481 (N_19481,N_18829,N_18642);
or U19482 (N_19482,N_18671,N_18587);
and U19483 (N_19483,N_18838,N_18672);
and U19484 (N_19484,N_18946,N_18920);
and U19485 (N_19485,N_18965,N_18757);
or U19486 (N_19486,N_18563,N_18507);
xnor U19487 (N_19487,N_18777,N_18617);
or U19488 (N_19488,N_18872,N_18811);
and U19489 (N_19489,N_18752,N_18728);
and U19490 (N_19490,N_18764,N_18681);
nor U19491 (N_19491,N_18832,N_18653);
nor U19492 (N_19492,N_18982,N_18682);
nor U19493 (N_19493,N_18681,N_18928);
and U19494 (N_19494,N_18981,N_18938);
nand U19495 (N_19495,N_18540,N_18761);
or U19496 (N_19496,N_18860,N_18997);
and U19497 (N_19497,N_18833,N_18859);
and U19498 (N_19498,N_18568,N_18546);
xnor U19499 (N_19499,N_18622,N_18635);
or U19500 (N_19500,N_19112,N_19413);
nand U19501 (N_19501,N_19405,N_19020);
and U19502 (N_19502,N_19293,N_19389);
and U19503 (N_19503,N_19437,N_19295);
and U19504 (N_19504,N_19249,N_19376);
or U19505 (N_19505,N_19266,N_19178);
nor U19506 (N_19506,N_19264,N_19019);
nand U19507 (N_19507,N_19077,N_19425);
nand U19508 (N_19508,N_19270,N_19487);
nand U19509 (N_19509,N_19001,N_19203);
nor U19510 (N_19510,N_19248,N_19464);
and U19511 (N_19511,N_19120,N_19118);
or U19512 (N_19512,N_19371,N_19158);
nand U19513 (N_19513,N_19333,N_19335);
nor U19514 (N_19514,N_19100,N_19435);
nor U19515 (N_19515,N_19367,N_19091);
xnor U19516 (N_19516,N_19407,N_19244);
nor U19517 (N_19517,N_19459,N_19466);
xor U19518 (N_19518,N_19281,N_19300);
xnor U19519 (N_19519,N_19320,N_19237);
nand U19520 (N_19520,N_19059,N_19103);
xnor U19521 (N_19521,N_19150,N_19061);
nand U19522 (N_19522,N_19067,N_19155);
nand U19523 (N_19523,N_19206,N_19431);
nand U19524 (N_19524,N_19280,N_19218);
xor U19525 (N_19525,N_19406,N_19098);
and U19526 (N_19526,N_19176,N_19054);
or U19527 (N_19527,N_19330,N_19325);
nor U19528 (N_19528,N_19065,N_19488);
nor U19529 (N_19529,N_19354,N_19148);
nor U19530 (N_19530,N_19250,N_19201);
nand U19531 (N_19531,N_19399,N_19035);
nor U19532 (N_19532,N_19381,N_19398);
and U19533 (N_19533,N_19424,N_19029);
or U19534 (N_19534,N_19334,N_19274);
nor U19535 (N_19535,N_19440,N_19132);
xor U19536 (N_19536,N_19047,N_19272);
or U19537 (N_19537,N_19338,N_19439);
nor U19538 (N_19538,N_19179,N_19004);
nor U19539 (N_19539,N_19472,N_19277);
nand U19540 (N_19540,N_19324,N_19495);
and U19541 (N_19541,N_19049,N_19257);
nand U19542 (N_19542,N_19013,N_19071);
nor U19543 (N_19543,N_19225,N_19379);
xor U19544 (N_19544,N_19349,N_19093);
xnor U19545 (N_19545,N_19370,N_19129);
and U19546 (N_19546,N_19243,N_19471);
and U19547 (N_19547,N_19139,N_19119);
nor U19548 (N_19548,N_19468,N_19457);
and U19549 (N_19549,N_19219,N_19197);
and U19550 (N_19550,N_19473,N_19090);
nor U19551 (N_19551,N_19023,N_19142);
xnor U19552 (N_19552,N_19469,N_19362);
nor U19553 (N_19553,N_19111,N_19068);
nand U19554 (N_19554,N_19253,N_19000);
nand U19555 (N_19555,N_19105,N_19316);
and U19556 (N_19556,N_19092,N_19127);
and U19557 (N_19557,N_19454,N_19131);
xnor U19558 (N_19558,N_19496,N_19391);
and U19559 (N_19559,N_19213,N_19251);
or U19560 (N_19560,N_19221,N_19200);
xnor U19561 (N_19561,N_19319,N_19121);
xor U19562 (N_19562,N_19322,N_19348);
nor U19563 (N_19563,N_19263,N_19076);
nor U19564 (N_19564,N_19169,N_19028);
and U19565 (N_19565,N_19477,N_19339);
nand U19566 (N_19566,N_19368,N_19246);
or U19567 (N_19567,N_19006,N_19073);
and U19568 (N_19568,N_19202,N_19027);
xor U19569 (N_19569,N_19140,N_19446);
nand U19570 (N_19570,N_19040,N_19401);
and U19571 (N_19571,N_19494,N_19184);
xnor U19572 (N_19572,N_19198,N_19475);
or U19573 (N_19573,N_19123,N_19145);
nor U19574 (N_19574,N_19384,N_19448);
and U19575 (N_19575,N_19375,N_19144);
or U19576 (N_19576,N_19080,N_19043);
nor U19577 (N_19577,N_19408,N_19192);
and U19578 (N_19578,N_19404,N_19358);
xor U19579 (N_19579,N_19302,N_19493);
and U19580 (N_19580,N_19180,N_19018);
or U19581 (N_19581,N_19008,N_19151);
nand U19582 (N_19582,N_19104,N_19419);
nor U19583 (N_19583,N_19489,N_19102);
nand U19584 (N_19584,N_19294,N_19069);
nand U19585 (N_19585,N_19474,N_19188);
or U19586 (N_19586,N_19329,N_19356);
and U19587 (N_19587,N_19327,N_19409);
nand U19588 (N_19588,N_19438,N_19156);
nand U19589 (N_19589,N_19113,N_19177);
nand U19590 (N_19590,N_19441,N_19212);
xnor U19591 (N_19591,N_19481,N_19296);
or U19592 (N_19592,N_19117,N_19497);
and U19593 (N_19593,N_19275,N_19285);
nor U19594 (N_19594,N_19074,N_19014);
and U19595 (N_19595,N_19462,N_19088);
xnor U19596 (N_19596,N_19394,N_19268);
nor U19597 (N_19597,N_19411,N_19422);
and U19598 (N_19598,N_19057,N_19314);
and U19599 (N_19599,N_19216,N_19174);
xor U19600 (N_19600,N_19421,N_19323);
nor U19601 (N_19601,N_19133,N_19382);
nor U19602 (N_19602,N_19208,N_19012);
xor U19603 (N_19603,N_19051,N_19031);
and U19604 (N_19604,N_19101,N_19491);
nand U19605 (N_19605,N_19415,N_19352);
nand U19606 (N_19606,N_19366,N_19038);
and U19607 (N_19607,N_19254,N_19340);
xnor U19608 (N_19608,N_19490,N_19153);
nand U19609 (N_19609,N_19172,N_19055);
xor U19610 (N_19610,N_19189,N_19351);
nand U19611 (N_19611,N_19380,N_19220);
and U19612 (N_19612,N_19239,N_19159);
nor U19613 (N_19613,N_19154,N_19373);
or U19614 (N_19614,N_19483,N_19363);
and U19615 (N_19615,N_19041,N_19060);
xor U19616 (N_19616,N_19233,N_19171);
nor U19617 (N_19617,N_19279,N_19194);
nor U19618 (N_19618,N_19222,N_19265);
nor U19619 (N_19619,N_19304,N_19024);
nand U19620 (N_19620,N_19343,N_19393);
nand U19621 (N_19621,N_19010,N_19412);
nor U19622 (N_19622,N_19321,N_19478);
and U19623 (N_19623,N_19070,N_19433);
xor U19624 (N_19624,N_19007,N_19183);
xor U19625 (N_19625,N_19033,N_19094);
and U19626 (N_19626,N_19303,N_19453);
nor U19627 (N_19627,N_19455,N_19463);
nor U19628 (N_19628,N_19242,N_19350);
nor U19629 (N_19629,N_19204,N_19479);
xor U19630 (N_19630,N_19449,N_19291);
or U19631 (N_19631,N_19283,N_19387);
and U19632 (N_19632,N_19317,N_19149);
and U19633 (N_19633,N_19465,N_19097);
nand U19634 (N_19634,N_19143,N_19232);
or U19635 (N_19635,N_19357,N_19223);
xor U19636 (N_19636,N_19480,N_19025);
nor U19637 (N_19637,N_19026,N_19130);
xnor U19638 (N_19638,N_19122,N_19498);
nor U19639 (N_19639,N_19191,N_19185);
xnor U19640 (N_19640,N_19482,N_19138);
xor U19641 (N_19641,N_19075,N_19116);
or U19642 (N_19642,N_19445,N_19361);
nor U19643 (N_19643,N_19467,N_19128);
nor U19644 (N_19644,N_19241,N_19209);
nand U19645 (N_19645,N_19452,N_19199);
nand U19646 (N_19646,N_19499,N_19292);
and U19647 (N_19647,N_19282,N_19084);
nand U19648 (N_19648,N_19400,N_19476);
xor U19649 (N_19649,N_19460,N_19211);
nand U19650 (N_19650,N_19353,N_19360);
nand U19651 (N_19651,N_19332,N_19364);
and U19652 (N_19652,N_19346,N_19426);
xnor U19653 (N_19653,N_19196,N_19125);
and U19654 (N_19654,N_19255,N_19078);
nor U19655 (N_19655,N_19427,N_19458);
or U19656 (N_19656,N_19227,N_19372);
nor U19657 (N_19657,N_19044,N_19450);
or U19658 (N_19658,N_19082,N_19141);
xnor U19659 (N_19659,N_19170,N_19388);
nand U19660 (N_19660,N_19456,N_19416);
or U19661 (N_19661,N_19053,N_19048);
and U19662 (N_19662,N_19215,N_19072);
or U19663 (N_19663,N_19085,N_19087);
and U19664 (N_19664,N_19245,N_19374);
xor U19665 (N_19665,N_19305,N_19229);
nor U19666 (N_19666,N_19036,N_19318);
nor U19667 (N_19667,N_19443,N_19066);
nand U19668 (N_19668,N_19236,N_19336);
and U19669 (N_19669,N_19058,N_19287);
nand U19670 (N_19670,N_19286,N_19418);
nor U19671 (N_19671,N_19308,N_19157);
and U19672 (N_19672,N_19434,N_19230);
nor U19673 (N_19673,N_19261,N_19423);
nand U19674 (N_19674,N_19345,N_19039);
and U19675 (N_19675,N_19052,N_19392);
or U19676 (N_19676,N_19262,N_19310);
nor U19677 (N_19677,N_19313,N_19195);
or U19678 (N_19678,N_19108,N_19432);
nor U19679 (N_19679,N_19484,N_19276);
or U19680 (N_19680,N_19390,N_19311);
xnor U19681 (N_19681,N_19003,N_19420);
nor U19682 (N_19682,N_19086,N_19163);
and U19683 (N_19683,N_19217,N_19385);
and U19684 (N_19684,N_19021,N_19240);
xnor U19685 (N_19685,N_19032,N_19114);
nand U19686 (N_19686,N_19009,N_19386);
or U19687 (N_19687,N_19395,N_19298);
or U19688 (N_19688,N_19016,N_19147);
or U19689 (N_19689,N_19429,N_19259);
nor U19690 (N_19690,N_19377,N_19289);
and U19691 (N_19691,N_19344,N_19436);
nand U19692 (N_19692,N_19110,N_19260);
xnor U19693 (N_19693,N_19030,N_19290);
xor U19694 (N_19694,N_19252,N_19359);
nor U19695 (N_19695,N_19089,N_19042);
nand U19696 (N_19696,N_19306,N_19461);
or U19697 (N_19697,N_19485,N_19050);
nor U19698 (N_19698,N_19447,N_19005);
nand U19699 (N_19699,N_19397,N_19383);
or U19700 (N_19700,N_19083,N_19312);
nor U19701 (N_19701,N_19107,N_19079);
nand U19702 (N_19702,N_19095,N_19267);
and U19703 (N_19703,N_19224,N_19161);
nor U19704 (N_19704,N_19164,N_19045);
nor U19705 (N_19705,N_19297,N_19328);
nand U19706 (N_19706,N_19109,N_19247);
and U19707 (N_19707,N_19002,N_19062);
nor U19708 (N_19708,N_19037,N_19126);
nor U19709 (N_19709,N_19234,N_19081);
and U19710 (N_19710,N_19315,N_19167);
or U19711 (N_19711,N_19063,N_19428);
or U19712 (N_19712,N_19168,N_19430);
nor U19713 (N_19713,N_19355,N_19369);
nand U19714 (N_19714,N_19137,N_19205);
nand U19715 (N_19715,N_19064,N_19011);
nor U19716 (N_19716,N_19403,N_19106);
or U19717 (N_19717,N_19175,N_19410);
or U19718 (N_19718,N_19046,N_19166);
nor U19719 (N_19719,N_19417,N_19347);
nor U19720 (N_19720,N_19326,N_19442);
nor U19721 (N_19721,N_19470,N_19288);
and U19722 (N_19722,N_19301,N_19022);
or U19723 (N_19723,N_19182,N_19056);
or U19724 (N_19724,N_19226,N_19258);
and U19725 (N_19725,N_19181,N_19269);
and U19726 (N_19726,N_19271,N_19238);
and U19727 (N_19727,N_19378,N_19309);
xor U19728 (N_19728,N_19214,N_19273);
nand U19729 (N_19729,N_19451,N_19187);
nand U19730 (N_19730,N_19190,N_19402);
xnor U19731 (N_19731,N_19331,N_19486);
or U19732 (N_19732,N_19207,N_19256);
or U19733 (N_19733,N_19228,N_19165);
or U19734 (N_19734,N_19342,N_19135);
xor U19735 (N_19735,N_19160,N_19015);
nor U19736 (N_19736,N_19115,N_19186);
or U19737 (N_19737,N_19096,N_19134);
nor U19738 (N_19738,N_19492,N_19365);
and U19739 (N_19739,N_19210,N_19396);
and U19740 (N_19740,N_19337,N_19136);
and U19741 (N_19741,N_19444,N_19173);
or U19742 (N_19742,N_19299,N_19278);
nor U19743 (N_19743,N_19162,N_19284);
nand U19744 (N_19744,N_19099,N_19152);
and U19745 (N_19745,N_19307,N_19414);
nor U19746 (N_19746,N_19146,N_19231);
nand U19747 (N_19747,N_19193,N_19017);
nor U19748 (N_19748,N_19235,N_19341);
xnor U19749 (N_19749,N_19034,N_19124);
nand U19750 (N_19750,N_19001,N_19312);
nor U19751 (N_19751,N_19174,N_19078);
nand U19752 (N_19752,N_19047,N_19196);
and U19753 (N_19753,N_19400,N_19242);
xor U19754 (N_19754,N_19211,N_19188);
nand U19755 (N_19755,N_19399,N_19236);
and U19756 (N_19756,N_19062,N_19200);
or U19757 (N_19757,N_19427,N_19275);
nor U19758 (N_19758,N_19035,N_19096);
and U19759 (N_19759,N_19230,N_19496);
xnor U19760 (N_19760,N_19127,N_19417);
nor U19761 (N_19761,N_19200,N_19276);
xnor U19762 (N_19762,N_19348,N_19155);
xnor U19763 (N_19763,N_19132,N_19179);
xor U19764 (N_19764,N_19088,N_19316);
and U19765 (N_19765,N_19376,N_19018);
nand U19766 (N_19766,N_19035,N_19197);
nor U19767 (N_19767,N_19023,N_19166);
or U19768 (N_19768,N_19410,N_19038);
xor U19769 (N_19769,N_19009,N_19214);
and U19770 (N_19770,N_19234,N_19143);
xnor U19771 (N_19771,N_19119,N_19375);
xor U19772 (N_19772,N_19326,N_19367);
nand U19773 (N_19773,N_19470,N_19037);
nor U19774 (N_19774,N_19172,N_19236);
and U19775 (N_19775,N_19185,N_19192);
or U19776 (N_19776,N_19306,N_19498);
nand U19777 (N_19777,N_19281,N_19397);
nor U19778 (N_19778,N_19020,N_19366);
nor U19779 (N_19779,N_19052,N_19326);
or U19780 (N_19780,N_19247,N_19260);
nand U19781 (N_19781,N_19060,N_19275);
or U19782 (N_19782,N_19115,N_19444);
or U19783 (N_19783,N_19057,N_19187);
and U19784 (N_19784,N_19010,N_19009);
or U19785 (N_19785,N_19199,N_19352);
or U19786 (N_19786,N_19371,N_19426);
nand U19787 (N_19787,N_19095,N_19446);
xnor U19788 (N_19788,N_19289,N_19332);
nand U19789 (N_19789,N_19166,N_19027);
or U19790 (N_19790,N_19073,N_19121);
xor U19791 (N_19791,N_19216,N_19138);
nor U19792 (N_19792,N_19454,N_19019);
and U19793 (N_19793,N_19176,N_19301);
nor U19794 (N_19794,N_19337,N_19353);
or U19795 (N_19795,N_19221,N_19458);
nand U19796 (N_19796,N_19255,N_19140);
or U19797 (N_19797,N_19442,N_19031);
and U19798 (N_19798,N_19010,N_19047);
nand U19799 (N_19799,N_19144,N_19497);
or U19800 (N_19800,N_19252,N_19117);
xnor U19801 (N_19801,N_19229,N_19440);
and U19802 (N_19802,N_19459,N_19360);
nand U19803 (N_19803,N_19061,N_19456);
xor U19804 (N_19804,N_19497,N_19344);
nand U19805 (N_19805,N_19363,N_19486);
xor U19806 (N_19806,N_19288,N_19422);
or U19807 (N_19807,N_19195,N_19241);
nand U19808 (N_19808,N_19227,N_19088);
and U19809 (N_19809,N_19173,N_19430);
nand U19810 (N_19810,N_19434,N_19228);
nand U19811 (N_19811,N_19272,N_19114);
nor U19812 (N_19812,N_19463,N_19025);
nand U19813 (N_19813,N_19160,N_19366);
xnor U19814 (N_19814,N_19069,N_19129);
nor U19815 (N_19815,N_19254,N_19399);
nand U19816 (N_19816,N_19089,N_19021);
xnor U19817 (N_19817,N_19104,N_19329);
and U19818 (N_19818,N_19474,N_19403);
and U19819 (N_19819,N_19439,N_19480);
or U19820 (N_19820,N_19322,N_19021);
nand U19821 (N_19821,N_19346,N_19117);
nor U19822 (N_19822,N_19128,N_19471);
nand U19823 (N_19823,N_19405,N_19135);
or U19824 (N_19824,N_19209,N_19230);
nand U19825 (N_19825,N_19224,N_19419);
nor U19826 (N_19826,N_19141,N_19467);
and U19827 (N_19827,N_19414,N_19449);
and U19828 (N_19828,N_19252,N_19387);
xor U19829 (N_19829,N_19249,N_19487);
nor U19830 (N_19830,N_19112,N_19369);
and U19831 (N_19831,N_19317,N_19269);
xor U19832 (N_19832,N_19295,N_19061);
nand U19833 (N_19833,N_19121,N_19341);
and U19834 (N_19834,N_19179,N_19083);
and U19835 (N_19835,N_19417,N_19449);
and U19836 (N_19836,N_19251,N_19294);
xnor U19837 (N_19837,N_19427,N_19351);
nor U19838 (N_19838,N_19334,N_19056);
or U19839 (N_19839,N_19318,N_19165);
xnor U19840 (N_19840,N_19000,N_19384);
nor U19841 (N_19841,N_19087,N_19465);
nand U19842 (N_19842,N_19357,N_19192);
xor U19843 (N_19843,N_19119,N_19104);
or U19844 (N_19844,N_19497,N_19197);
and U19845 (N_19845,N_19331,N_19005);
and U19846 (N_19846,N_19084,N_19476);
xnor U19847 (N_19847,N_19010,N_19033);
and U19848 (N_19848,N_19199,N_19283);
nand U19849 (N_19849,N_19189,N_19043);
and U19850 (N_19850,N_19138,N_19215);
nand U19851 (N_19851,N_19313,N_19479);
or U19852 (N_19852,N_19128,N_19191);
or U19853 (N_19853,N_19147,N_19264);
or U19854 (N_19854,N_19202,N_19099);
nor U19855 (N_19855,N_19197,N_19098);
or U19856 (N_19856,N_19320,N_19187);
nand U19857 (N_19857,N_19068,N_19325);
xnor U19858 (N_19858,N_19479,N_19169);
and U19859 (N_19859,N_19025,N_19383);
or U19860 (N_19860,N_19316,N_19278);
nand U19861 (N_19861,N_19344,N_19025);
nor U19862 (N_19862,N_19158,N_19012);
and U19863 (N_19863,N_19120,N_19185);
and U19864 (N_19864,N_19451,N_19055);
and U19865 (N_19865,N_19439,N_19399);
nand U19866 (N_19866,N_19455,N_19413);
nor U19867 (N_19867,N_19077,N_19131);
or U19868 (N_19868,N_19118,N_19386);
nand U19869 (N_19869,N_19309,N_19085);
nand U19870 (N_19870,N_19485,N_19498);
and U19871 (N_19871,N_19069,N_19483);
or U19872 (N_19872,N_19123,N_19373);
nor U19873 (N_19873,N_19093,N_19460);
xor U19874 (N_19874,N_19034,N_19328);
nand U19875 (N_19875,N_19470,N_19088);
and U19876 (N_19876,N_19242,N_19453);
nand U19877 (N_19877,N_19097,N_19217);
nor U19878 (N_19878,N_19189,N_19242);
xor U19879 (N_19879,N_19390,N_19204);
nor U19880 (N_19880,N_19123,N_19014);
nand U19881 (N_19881,N_19021,N_19109);
nand U19882 (N_19882,N_19313,N_19259);
or U19883 (N_19883,N_19156,N_19221);
or U19884 (N_19884,N_19034,N_19247);
and U19885 (N_19885,N_19219,N_19246);
xor U19886 (N_19886,N_19400,N_19025);
xor U19887 (N_19887,N_19364,N_19290);
and U19888 (N_19888,N_19418,N_19497);
nand U19889 (N_19889,N_19140,N_19035);
and U19890 (N_19890,N_19398,N_19318);
xnor U19891 (N_19891,N_19247,N_19076);
and U19892 (N_19892,N_19225,N_19369);
nor U19893 (N_19893,N_19178,N_19049);
or U19894 (N_19894,N_19469,N_19064);
and U19895 (N_19895,N_19097,N_19489);
xnor U19896 (N_19896,N_19226,N_19026);
nor U19897 (N_19897,N_19353,N_19454);
xnor U19898 (N_19898,N_19103,N_19390);
nor U19899 (N_19899,N_19322,N_19402);
nor U19900 (N_19900,N_19411,N_19470);
xor U19901 (N_19901,N_19301,N_19401);
nor U19902 (N_19902,N_19133,N_19344);
nor U19903 (N_19903,N_19117,N_19290);
or U19904 (N_19904,N_19325,N_19432);
nand U19905 (N_19905,N_19411,N_19427);
xor U19906 (N_19906,N_19202,N_19106);
xnor U19907 (N_19907,N_19452,N_19471);
or U19908 (N_19908,N_19021,N_19332);
nand U19909 (N_19909,N_19178,N_19126);
or U19910 (N_19910,N_19108,N_19271);
nand U19911 (N_19911,N_19006,N_19318);
nand U19912 (N_19912,N_19369,N_19438);
and U19913 (N_19913,N_19400,N_19321);
nand U19914 (N_19914,N_19022,N_19317);
nand U19915 (N_19915,N_19417,N_19400);
nor U19916 (N_19916,N_19150,N_19346);
xnor U19917 (N_19917,N_19058,N_19304);
nand U19918 (N_19918,N_19343,N_19021);
nor U19919 (N_19919,N_19278,N_19137);
nand U19920 (N_19920,N_19167,N_19052);
or U19921 (N_19921,N_19185,N_19004);
nand U19922 (N_19922,N_19332,N_19280);
nand U19923 (N_19923,N_19449,N_19424);
xnor U19924 (N_19924,N_19290,N_19051);
xnor U19925 (N_19925,N_19427,N_19449);
or U19926 (N_19926,N_19426,N_19340);
nor U19927 (N_19927,N_19034,N_19153);
nor U19928 (N_19928,N_19313,N_19425);
and U19929 (N_19929,N_19402,N_19248);
or U19930 (N_19930,N_19433,N_19026);
or U19931 (N_19931,N_19284,N_19059);
nor U19932 (N_19932,N_19066,N_19189);
and U19933 (N_19933,N_19267,N_19262);
nor U19934 (N_19934,N_19136,N_19113);
nand U19935 (N_19935,N_19141,N_19415);
nand U19936 (N_19936,N_19342,N_19333);
nor U19937 (N_19937,N_19038,N_19093);
or U19938 (N_19938,N_19473,N_19487);
nor U19939 (N_19939,N_19326,N_19058);
xor U19940 (N_19940,N_19452,N_19031);
or U19941 (N_19941,N_19484,N_19032);
xor U19942 (N_19942,N_19267,N_19284);
or U19943 (N_19943,N_19393,N_19142);
xor U19944 (N_19944,N_19221,N_19185);
or U19945 (N_19945,N_19218,N_19191);
nand U19946 (N_19946,N_19067,N_19097);
nand U19947 (N_19947,N_19198,N_19038);
nand U19948 (N_19948,N_19349,N_19064);
nor U19949 (N_19949,N_19360,N_19201);
xor U19950 (N_19950,N_19382,N_19347);
or U19951 (N_19951,N_19439,N_19103);
and U19952 (N_19952,N_19189,N_19170);
and U19953 (N_19953,N_19026,N_19262);
nor U19954 (N_19954,N_19120,N_19153);
nor U19955 (N_19955,N_19304,N_19447);
and U19956 (N_19956,N_19037,N_19286);
or U19957 (N_19957,N_19110,N_19395);
nand U19958 (N_19958,N_19255,N_19404);
and U19959 (N_19959,N_19060,N_19161);
xor U19960 (N_19960,N_19364,N_19411);
or U19961 (N_19961,N_19360,N_19396);
and U19962 (N_19962,N_19375,N_19280);
and U19963 (N_19963,N_19169,N_19319);
nor U19964 (N_19964,N_19447,N_19329);
nand U19965 (N_19965,N_19063,N_19211);
and U19966 (N_19966,N_19103,N_19489);
and U19967 (N_19967,N_19056,N_19442);
or U19968 (N_19968,N_19491,N_19470);
or U19969 (N_19969,N_19045,N_19331);
nor U19970 (N_19970,N_19370,N_19222);
xnor U19971 (N_19971,N_19487,N_19406);
nor U19972 (N_19972,N_19265,N_19163);
and U19973 (N_19973,N_19386,N_19154);
nor U19974 (N_19974,N_19077,N_19430);
xor U19975 (N_19975,N_19229,N_19065);
nand U19976 (N_19976,N_19215,N_19286);
nor U19977 (N_19977,N_19409,N_19287);
or U19978 (N_19978,N_19020,N_19290);
xnor U19979 (N_19979,N_19420,N_19247);
or U19980 (N_19980,N_19274,N_19062);
and U19981 (N_19981,N_19312,N_19092);
and U19982 (N_19982,N_19208,N_19387);
or U19983 (N_19983,N_19410,N_19037);
nor U19984 (N_19984,N_19023,N_19360);
or U19985 (N_19985,N_19372,N_19337);
xor U19986 (N_19986,N_19485,N_19360);
nor U19987 (N_19987,N_19020,N_19252);
nand U19988 (N_19988,N_19479,N_19298);
nand U19989 (N_19989,N_19444,N_19237);
or U19990 (N_19990,N_19197,N_19459);
nand U19991 (N_19991,N_19248,N_19341);
or U19992 (N_19992,N_19469,N_19340);
xor U19993 (N_19993,N_19070,N_19394);
xnor U19994 (N_19994,N_19196,N_19383);
nor U19995 (N_19995,N_19164,N_19093);
and U19996 (N_19996,N_19100,N_19036);
nand U19997 (N_19997,N_19499,N_19058);
xor U19998 (N_19998,N_19417,N_19268);
nor U19999 (N_19999,N_19306,N_19464);
nand UO_0 (O_0,N_19699,N_19665);
xnor UO_1 (O_1,N_19920,N_19502);
nand UO_2 (O_2,N_19565,N_19796);
and UO_3 (O_3,N_19926,N_19939);
nand UO_4 (O_4,N_19652,N_19521);
nor UO_5 (O_5,N_19578,N_19823);
nand UO_6 (O_6,N_19810,N_19558);
nor UO_7 (O_7,N_19932,N_19539);
nand UO_8 (O_8,N_19529,N_19595);
nor UO_9 (O_9,N_19639,N_19621);
nand UO_10 (O_10,N_19566,N_19725);
xnor UO_11 (O_11,N_19936,N_19772);
nor UO_12 (O_12,N_19960,N_19569);
and UO_13 (O_13,N_19694,N_19604);
nor UO_14 (O_14,N_19682,N_19750);
nor UO_15 (O_15,N_19907,N_19802);
xnor UO_16 (O_16,N_19943,N_19633);
nor UO_17 (O_17,N_19818,N_19861);
and UO_18 (O_18,N_19528,N_19648);
or UO_19 (O_19,N_19698,N_19641);
and UO_20 (O_20,N_19608,N_19613);
or UO_21 (O_21,N_19540,N_19852);
and UO_22 (O_22,N_19935,N_19617);
and UO_23 (O_23,N_19544,N_19782);
or UO_24 (O_24,N_19841,N_19792);
xnor UO_25 (O_25,N_19771,N_19689);
and UO_26 (O_26,N_19761,N_19680);
xnor UO_27 (O_27,N_19560,N_19535);
nor UO_28 (O_28,N_19649,N_19924);
xnor UO_29 (O_29,N_19630,N_19514);
and UO_30 (O_30,N_19914,N_19501);
and UO_31 (O_31,N_19770,N_19610);
nor UO_32 (O_32,N_19599,N_19942);
xnor UO_33 (O_33,N_19571,N_19657);
nand UO_34 (O_34,N_19500,N_19773);
xnor UO_35 (O_35,N_19508,N_19755);
and UO_36 (O_36,N_19865,N_19996);
nor UO_37 (O_37,N_19855,N_19780);
or UO_38 (O_38,N_19874,N_19575);
nand UO_39 (O_39,N_19949,N_19702);
or UO_40 (O_40,N_19668,N_19846);
and UO_41 (O_41,N_19828,N_19813);
nor UO_42 (O_42,N_19509,N_19741);
nand UO_43 (O_43,N_19888,N_19614);
and UO_44 (O_44,N_19644,N_19534);
nand UO_45 (O_45,N_19588,N_19891);
xor UO_46 (O_46,N_19646,N_19748);
nor UO_47 (O_47,N_19800,N_19906);
xnor UO_48 (O_48,N_19990,N_19765);
xor UO_49 (O_49,N_19854,N_19980);
and UO_50 (O_50,N_19851,N_19834);
xor UO_51 (O_51,N_19701,N_19915);
nor UO_52 (O_52,N_19515,N_19928);
nor UO_53 (O_53,N_19808,N_19954);
nor UO_54 (O_54,N_19863,N_19760);
and UO_55 (O_55,N_19551,N_19688);
nor UO_56 (O_56,N_19783,N_19628);
xor UO_57 (O_57,N_19871,N_19972);
xnor UO_58 (O_58,N_19903,N_19594);
nand UO_59 (O_59,N_19849,N_19913);
nor UO_60 (O_60,N_19733,N_19971);
and UO_61 (O_61,N_19807,N_19909);
or UO_62 (O_62,N_19975,N_19732);
and UO_63 (O_63,N_19611,N_19864);
nand UO_64 (O_64,N_19884,N_19685);
nor UO_65 (O_65,N_19712,N_19693);
and UO_66 (O_66,N_19775,N_19713);
and UO_67 (O_67,N_19727,N_19723);
and UO_68 (O_68,N_19679,N_19798);
nor UO_69 (O_69,N_19793,N_19862);
nand UO_70 (O_70,N_19634,N_19526);
and UO_71 (O_71,N_19989,N_19919);
and UO_72 (O_72,N_19692,N_19969);
or UO_73 (O_73,N_19553,N_19885);
nor UO_74 (O_74,N_19892,N_19684);
or UO_75 (O_75,N_19708,N_19764);
nor UO_76 (O_76,N_19756,N_19647);
or UO_77 (O_77,N_19979,N_19606);
xor UO_78 (O_78,N_19872,N_19923);
nand UO_79 (O_79,N_19774,N_19769);
and UO_80 (O_80,N_19779,N_19789);
or UO_81 (O_81,N_19816,N_19519);
nand UO_82 (O_82,N_19520,N_19934);
xnor UO_83 (O_83,N_19958,N_19522);
and UO_84 (O_84,N_19794,N_19597);
xnor UO_85 (O_85,N_19678,N_19850);
and UO_86 (O_86,N_19687,N_19746);
xnor UO_87 (O_87,N_19838,N_19981);
xnor UO_88 (O_88,N_19695,N_19632);
xnor UO_89 (O_89,N_19592,N_19690);
nor UO_90 (O_90,N_19982,N_19504);
or UO_91 (O_91,N_19985,N_19955);
and UO_92 (O_92,N_19973,N_19567);
and UO_93 (O_93,N_19587,N_19922);
or UO_94 (O_94,N_19977,N_19559);
and UO_95 (O_95,N_19556,N_19615);
and UO_96 (O_96,N_19803,N_19601);
and UO_97 (O_97,N_19825,N_19811);
and UO_98 (O_98,N_19564,N_19758);
nand UO_99 (O_99,N_19676,N_19661);
or UO_100 (O_100,N_19867,N_19966);
nand UO_101 (O_101,N_19552,N_19759);
nor UO_102 (O_102,N_19877,N_19666);
nor UO_103 (O_103,N_19511,N_19591);
nor UO_104 (O_104,N_19660,N_19705);
nand UO_105 (O_105,N_19635,N_19786);
nand UO_106 (O_106,N_19921,N_19523);
nor UO_107 (O_107,N_19768,N_19625);
xnor UO_108 (O_108,N_19876,N_19734);
nor UO_109 (O_109,N_19506,N_19925);
or UO_110 (O_110,N_19663,N_19656);
xor UO_111 (O_111,N_19724,N_19557);
and UO_112 (O_112,N_19518,N_19787);
or UO_113 (O_113,N_19911,N_19716);
and UO_114 (O_114,N_19722,N_19711);
or UO_115 (O_115,N_19815,N_19795);
and UO_116 (O_116,N_19858,N_19549);
nand UO_117 (O_117,N_19869,N_19817);
and UO_118 (O_118,N_19561,N_19857);
and UO_119 (O_119,N_19707,N_19910);
nor UO_120 (O_120,N_19930,N_19550);
nand UO_121 (O_121,N_19507,N_19653);
nand UO_122 (O_122,N_19714,N_19642);
nand UO_123 (O_123,N_19554,N_19754);
xor UO_124 (O_124,N_19898,N_19670);
and UO_125 (O_125,N_19726,N_19976);
or UO_126 (O_126,N_19753,N_19840);
or UO_127 (O_127,N_19586,N_19944);
xor UO_128 (O_128,N_19805,N_19933);
nand UO_129 (O_129,N_19721,N_19555);
nor UO_130 (O_130,N_19681,N_19839);
nor UO_131 (O_131,N_19883,N_19636);
or UO_132 (O_132,N_19709,N_19875);
and UO_133 (O_133,N_19640,N_19917);
nor UO_134 (O_134,N_19728,N_19988);
xnor UO_135 (O_135,N_19720,N_19737);
or UO_136 (O_136,N_19941,N_19532);
and UO_137 (O_137,N_19645,N_19579);
nand UO_138 (O_138,N_19997,N_19938);
nand UO_139 (O_139,N_19835,N_19847);
or UO_140 (O_140,N_19882,N_19710);
or UO_141 (O_141,N_19804,N_19964);
or UO_142 (O_142,N_19991,N_19947);
nor UO_143 (O_143,N_19583,N_19577);
xor UO_144 (O_144,N_19967,N_19951);
nand UO_145 (O_145,N_19890,N_19931);
nand UO_146 (O_146,N_19729,N_19992);
or UO_147 (O_147,N_19512,N_19830);
xor UO_148 (O_148,N_19836,N_19821);
nand UO_149 (O_149,N_19912,N_19516);
or UO_150 (O_150,N_19777,N_19744);
and UO_151 (O_151,N_19616,N_19873);
nor UO_152 (O_152,N_19669,N_19686);
or UO_153 (O_153,N_19600,N_19730);
nor UO_154 (O_154,N_19881,N_19700);
or UO_155 (O_155,N_19570,N_19905);
xor UO_156 (O_156,N_19580,N_19747);
and UO_157 (O_157,N_19643,N_19650);
nand UO_158 (O_158,N_19843,N_19607);
or UO_159 (O_159,N_19901,N_19609);
and UO_160 (O_160,N_19887,N_19831);
and UO_161 (O_161,N_19987,N_19762);
and UO_162 (O_162,N_19833,N_19696);
nor UO_163 (O_163,N_19745,N_19856);
nor UO_164 (O_164,N_19844,N_19829);
xnor UO_165 (O_165,N_19538,N_19781);
and UO_166 (O_166,N_19627,N_19624);
nand UO_167 (O_167,N_19530,N_19826);
and UO_168 (O_168,N_19859,N_19743);
and UO_169 (O_169,N_19623,N_19809);
and UO_170 (O_170,N_19791,N_19602);
and UO_171 (O_171,N_19605,N_19918);
nor UO_172 (O_172,N_19510,N_19766);
xor UO_173 (O_173,N_19984,N_19902);
nand UO_174 (O_174,N_19596,N_19590);
xnor UO_175 (O_175,N_19889,N_19658);
nor UO_176 (O_176,N_19806,N_19986);
and UO_177 (O_177,N_19799,N_19675);
nand UO_178 (O_178,N_19894,N_19998);
nor UO_179 (O_179,N_19896,N_19574);
nand UO_180 (O_180,N_19582,N_19790);
and UO_181 (O_181,N_19563,N_19593);
or UO_182 (O_182,N_19797,N_19963);
and UO_183 (O_183,N_19525,N_19814);
and UO_184 (O_184,N_19788,N_19572);
and UO_185 (O_185,N_19820,N_19697);
nor UO_186 (O_186,N_19671,N_19629);
xor UO_187 (O_187,N_19654,N_19703);
nand UO_188 (O_188,N_19893,N_19897);
xor UO_189 (O_189,N_19900,N_19505);
and UO_190 (O_190,N_19959,N_19824);
nor UO_191 (O_191,N_19965,N_19704);
nor UO_192 (O_192,N_19585,N_19503);
or UO_193 (O_193,N_19749,N_19545);
nand UO_194 (O_194,N_19738,N_19739);
nand UO_195 (O_195,N_19848,N_19940);
nor UO_196 (O_196,N_19784,N_19620);
or UO_197 (O_197,N_19879,N_19717);
xnor UO_198 (O_198,N_19853,N_19576);
and UO_199 (O_199,N_19763,N_19546);
nand UO_200 (O_200,N_19736,N_19677);
or UO_201 (O_201,N_19706,N_19880);
xnor UO_202 (O_202,N_19537,N_19752);
and UO_203 (O_203,N_19999,N_19719);
nor UO_204 (O_204,N_19995,N_19673);
nor UO_205 (O_205,N_19908,N_19742);
nand UO_206 (O_206,N_19812,N_19916);
nor UO_207 (O_207,N_19832,N_19672);
nand UO_208 (O_208,N_19598,N_19568);
nand UO_209 (O_209,N_19626,N_19562);
or UO_210 (O_210,N_19952,N_19637);
nor UO_211 (O_211,N_19983,N_19950);
and UO_212 (O_212,N_19664,N_19524);
xnor UO_213 (O_213,N_19767,N_19870);
nand UO_214 (O_214,N_19536,N_19584);
or UO_215 (O_215,N_19819,N_19622);
xnor UO_216 (O_216,N_19993,N_19822);
nor UO_217 (O_217,N_19937,N_19899);
nor UO_218 (O_218,N_19740,N_19929);
and UO_219 (O_219,N_19651,N_19776);
nor UO_220 (O_220,N_19927,N_19785);
nand UO_221 (O_221,N_19718,N_19837);
xor UO_222 (O_222,N_19527,N_19970);
or UO_223 (O_223,N_19751,N_19827);
or UO_224 (O_224,N_19619,N_19543);
nor UO_225 (O_225,N_19994,N_19962);
or UO_226 (O_226,N_19757,N_19589);
nor UO_227 (O_227,N_19956,N_19662);
and UO_228 (O_228,N_19581,N_19612);
or UO_229 (O_229,N_19961,N_19631);
nand UO_230 (O_230,N_19517,N_19674);
nand UO_231 (O_231,N_19603,N_19638);
or UO_232 (O_232,N_19978,N_19957);
nor UO_233 (O_233,N_19683,N_19968);
or UO_234 (O_234,N_19618,N_19659);
and UO_235 (O_235,N_19573,N_19895);
nand UO_236 (O_236,N_19731,N_19845);
nand UO_237 (O_237,N_19667,N_19904);
and UO_238 (O_238,N_19542,N_19878);
nand UO_239 (O_239,N_19541,N_19868);
or UO_240 (O_240,N_19691,N_19778);
nor UO_241 (O_241,N_19547,N_19715);
xnor UO_242 (O_242,N_19842,N_19513);
xor UO_243 (O_243,N_19953,N_19948);
nand UO_244 (O_244,N_19945,N_19886);
nor UO_245 (O_245,N_19655,N_19860);
and UO_246 (O_246,N_19533,N_19866);
and UO_247 (O_247,N_19801,N_19531);
or UO_248 (O_248,N_19735,N_19548);
nor UO_249 (O_249,N_19946,N_19974);
and UO_250 (O_250,N_19904,N_19761);
nand UO_251 (O_251,N_19587,N_19865);
and UO_252 (O_252,N_19708,N_19525);
xnor UO_253 (O_253,N_19945,N_19796);
xnor UO_254 (O_254,N_19803,N_19804);
nor UO_255 (O_255,N_19794,N_19911);
and UO_256 (O_256,N_19873,N_19733);
and UO_257 (O_257,N_19595,N_19505);
nor UO_258 (O_258,N_19815,N_19722);
nor UO_259 (O_259,N_19860,N_19526);
nor UO_260 (O_260,N_19631,N_19899);
nand UO_261 (O_261,N_19765,N_19616);
nand UO_262 (O_262,N_19955,N_19819);
xor UO_263 (O_263,N_19871,N_19656);
or UO_264 (O_264,N_19522,N_19592);
xnor UO_265 (O_265,N_19996,N_19725);
or UO_266 (O_266,N_19672,N_19946);
nand UO_267 (O_267,N_19942,N_19555);
nor UO_268 (O_268,N_19700,N_19950);
xor UO_269 (O_269,N_19969,N_19977);
nor UO_270 (O_270,N_19771,N_19709);
xnor UO_271 (O_271,N_19798,N_19778);
xor UO_272 (O_272,N_19884,N_19780);
nand UO_273 (O_273,N_19940,N_19698);
or UO_274 (O_274,N_19949,N_19892);
nand UO_275 (O_275,N_19562,N_19591);
nand UO_276 (O_276,N_19710,N_19659);
and UO_277 (O_277,N_19563,N_19542);
or UO_278 (O_278,N_19707,N_19712);
nor UO_279 (O_279,N_19978,N_19559);
or UO_280 (O_280,N_19667,N_19571);
or UO_281 (O_281,N_19790,N_19688);
or UO_282 (O_282,N_19791,N_19581);
nor UO_283 (O_283,N_19695,N_19861);
and UO_284 (O_284,N_19963,N_19777);
or UO_285 (O_285,N_19672,N_19551);
and UO_286 (O_286,N_19548,N_19627);
xnor UO_287 (O_287,N_19635,N_19682);
and UO_288 (O_288,N_19910,N_19781);
nor UO_289 (O_289,N_19836,N_19505);
nor UO_290 (O_290,N_19889,N_19558);
nand UO_291 (O_291,N_19689,N_19682);
nor UO_292 (O_292,N_19870,N_19895);
xnor UO_293 (O_293,N_19571,N_19890);
nor UO_294 (O_294,N_19876,N_19792);
xnor UO_295 (O_295,N_19947,N_19751);
and UO_296 (O_296,N_19574,N_19954);
or UO_297 (O_297,N_19940,N_19717);
xnor UO_298 (O_298,N_19548,N_19609);
and UO_299 (O_299,N_19845,N_19987);
xnor UO_300 (O_300,N_19801,N_19525);
nand UO_301 (O_301,N_19785,N_19697);
nor UO_302 (O_302,N_19923,N_19848);
nand UO_303 (O_303,N_19977,N_19692);
and UO_304 (O_304,N_19991,N_19690);
or UO_305 (O_305,N_19761,N_19567);
nor UO_306 (O_306,N_19563,N_19734);
xnor UO_307 (O_307,N_19647,N_19927);
xnor UO_308 (O_308,N_19749,N_19655);
or UO_309 (O_309,N_19606,N_19953);
and UO_310 (O_310,N_19566,N_19809);
xor UO_311 (O_311,N_19610,N_19644);
nor UO_312 (O_312,N_19862,N_19601);
nor UO_313 (O_313,N_19625,N_19832);
nand UO_314 (O_314,N_19717,N_19935);
nand UO_315 (O_315,N_19981,N_19630);
or UO_316 (O_316,N_19796,N_19709);
and UO_317 (O_317,N_19902,N_19531);
xor UO_318 (O_318,N_19657,N_19534);
or UO_319 (O_319,N_19993,N_19963);
and UO_320 (O_320,N_19913,N_19539);
xnor UO_321 (O_321,N_19794,N_19548);
xnor UO_322 (O_322,N_19532,N_19528);
nand UO_323 (O_323,N_19500,N_19762);
nor UO_324 (O_324,N_19926,N_19960);
and UO_325 (O_325,N_19930,N_19768);
nand UO_326 (O_326,N_19581,N_19950);
and UO_327 (O_327,N_19796,N_19830);
nor UO_328 (O_328,N_19633,N_19741);
and UO_329 (O_329,N_19738,N_19661);
xnor UO_330 (O_330,N_19897,N_19842);
nor UO_331 (O_331,N_19789,N_19749);
or UO_332 (O_332,N_19540,N_19908);
nor UO_333 (O_333,N_19927,N_19556);
and UO_334 (O_334,N_19969,N_19564);
or UO_335 (O_335,N_19694,N_19723);
or UO_336 (O_336,N_19973,N_19698);
nor UO_337 (O_337,N_19960,N_19858);
or UO_338 (O_338,N_19719,N_19672);
xnor UO_339 (O_339,N_19997,N_19903);
nor UO_340 (O_340,N_19558,N_19976);
nand UO_341 (O_341,N_19551,N_19775);
or UO_342 (O_342,N_19726,N_19655);
nand UO_343 (O_343,N_19932,N_19848);
nor UO_344 (O_344,N_19724,N_19739);
xor UO_345 (O_345,N_19527,N_19803);
xnor UO_346 (O_346,N_19968,N_19780);
nand UO_347 (O_347,N_19636,N_19888);
xnor UO_348 (O_348,N_19588,N_19999);
nand UO_349 (O_349,N_19882,N_19779);
and UO_350 (O_350,N_19856,N_19814);
and UO_351 (O_351,N_19605,N_19984);
xor UO_352 (O_352,N_19986,N_19657);
nor UO_353 (O_353,N_19814,N_19773);
and UO_354 (O_354,N_19681,N_19507);
nand UO_355 (O_355,N_19901,N_19656);
and UO_356 (O_356,N_19806,N_19560);
nand UO_357 (O_357,N_19543,N_19913);
and UO_358 (O_358,N_19556,N_19713);
xor UO_359 (O_359,N_19830,N_19921);
nand UO_360 (O_360,N_19511,N_19866);
nor UO_361 (O_361,N_19717,N_19557);
or UO_362 (O_362,N_19926,N_19794);
xor UO_363 (O_363,N_19558,N_19844);
or UO_364 (O_364,N_19810,N_19895);
xnor UO_365 (O_365,N_19540,N_19529);
xnor UO_366 (O_366,N_19602,N_19521);
xnor UO_367 (O_367,N_19857,N_19744);
and UO_368 (O_368,N_19787,N_19894);
or UO_369 (O_369,N_19533,N_19778);
and UO_370 (O_370,N_19653,N_19940);
xor UO_371 (O_371,N_19837,N_19509);
or UO_372 (O_372,N_19607,N_19656);
nand UO_373 (O_373,N_19576,N_19923);
and UO_374 (O_374,N_19749,N_19847);
or UO_375 (O_375,N_19882,N_19649);
or UO_376 (O_376,N_19658,N_19811);
nor UO_377 (O_377,N_19657,N_19582);
nor UO_378 (O_378,N_19737,N_19641);
or UO_379 (O_379,N_19817,N_19717);
nand UO_380 (O_380,N_19517,N_19980);
or UO_381 (O_381,N_19545,N_19842);
xor UO_382 (O_382,N_19799,N_19638);
xor UO_383 (O_383,N_19739,N_19968);
nor UO_384 (O_384,N_19685,N_19803);
xor UO_385 (O_385,N_19726,N_19706);
and UO_386 (O_386,N_19519,N_19729);
or UO_387 (O_387,N_19796,N_19822);
and UO_388 (O_388,N_19711,N_19737);
nor UO_389 (O_389,N_19922,N_19881);
nand UO_390 (O_390,N_19949,N_19917);
or UO_391 (O_391,N_19536,N_19804);
nand UO_392 (O_392,N_19891,N_19647);
xnor UO_393 (O_393,N_19936,N_19820);
xnor UO_394 (O_394,N_19663,N_19925);
nand UO_395 (O_395,N_19669,N_19624);
nand UO_396 (O_396,N_19738,N_19830);
nand UO_397 (O_397,N_19898,N_19617);
or UO_398 (O_398,N_19997,N_19720);
or UO_399 (O_399,N_19968,N_19606);
nand UO_400 (O_400,N_19854,N_19904);
xor UO_401 (O_401,N_19964,N_19676);
nand UO_402 (O_402,N_19847,N_19805);
and UO_403 (O_403,N_19700,N_19535);
and UO_404 (O_404,N_19922,N_19959);
or UO_405 (O_405,N_19924,N_19659);
or UO_406 (O_406,N_19916,N_19993);
and UO_407 (O_407,N_19934,N_19845);
nand UO_408 (O_408,N_19559,N_19560);
and UO_409 (O_409,N_19989,N_19644);
nand UO_410 (O_410,N_19687,N_19823);
xnor UO_411 (O_411,N_19815,N_19685);
and UO_412 (O_412,N_19608,N_19848);
and UO_413 (O_413,N_19982,N_19839);
or UO_414 (O_414,N_19903,N_19716);
xnor UO_415 (O_415,N_19877,N_19584);
nor UO_416 (O_416,N_19789,N_19917);
and UO_417 (O_417,N_19994,N_19512);
xnor UO_418 (O_418,N_19991,N_19788);
and UO_419 (O_419,N_19752,N_19548);
nand UO_420 (O_420,N_19720,N_19543);
nand UO_421 (O_421,N_19529,N_19605);
nand UO_422 (O_422,N_19961,N_19727);
or UO_423 (O_423,N_19732,N_19958);
nor UO_424 (O_424,N_19978,N_19693);
or UO_425 (O_425,N_19983,N_19695);
nor UO_426 (O_426,N_19807,N_19836);
or UO_427 (O_427,N_19675,N_19973);
nor UO_428 (O_428,N_19703,N_19924);
nor UO_429 (O_429,N_19750,N_19881);
nand UO_430 (O_430,N_19585,N_19569);
nor UO_431 (O_431,N_19682,N_19820);
xor UO_432 (O_432,N_19946,N_19905);
nor UO_433 (O_433,N_19863,N_19852);
or UO_434 (O_434,N_19633,N_19731);
or UO_435 (O_435,N_19734,N_19713);
or UO_436 (O_436,N_19806,N_19971);
and UO_437 (O_437,N_19692,N_19837);
xor UO_438 (O_438,N_19925,N_19764);
xnor UO_439 (O_439,N_19687,N_19579);
and UO_440 (O_440,N_19605,N_19666);
xor UO_441 (O_441,N_19876,N_19744);
nor UO_442 (O_442,N_19524,N_19970);
nand UO_443 (O_443,N_19975,N_19656);
nor UO_444 (O_444,N_19653,N_19707);
xnor UO_445 (O_445,N_19796,N_19542);
nand UO_446 (O_446,N_19701,N_19710);
nor UO_447 (O_447,N_19511,N_19805);
or UO_448 (O_448,N_19776,N_19744);
or UO_449 (O_449,N_19858,N_19969);
nand UO_450 (O_450,N_19843,N_19675);
and UO_451 (O_451,N_19796,N_19711);
nand UO_452 (O_452,N_19698,N_19754);
or UO_453 (O_453,N_19919,N_19688);
nor UO_454 (O_454,N_19524,N_19784);
or UO_455 (O_455,N_19621,N_19863);
and UO_456 (O_456,N_19641,N_19865);
xor UO_457 (O_457,N_19644,N_19504);
xor UO_458 (O_458,N_19862,N_19812);
and UO_459 (O_459,N_19733,N_19635);
or UO_460 (O_460,N_19834,N_19725);
nor UO_461 (O_461,N_19500,N_19820);
or UO_462 (O_462,N_19705,N_19846);
nand UO_463 (O_463,N_19597,N_19779);
or UO_464 (O_464,N_19959,N_19602);
nand UO_465 (O_465,N_19573,N_19768);
nand UO_466 (O_466,N_19809,N_19515);
and UO_467 (O_467,N_19839,N_19640);
and UO_468 (O_468,N_19813,N_19554);
nand UO_469 (O_469,N_19640,N_19761);
xor UO_470 (O_470,N_19972,N_19764);
and UO_471 (O_471,N_19891,N_19601);
or UO_472 (O_472,N_19696,N_19890);
and UO_473 (O_473,N_19821,N_19609);
and UO_474 (O_474,N_19880,N_19565);
xor UO_475 (O_475,N_19557,N_19543);
and UO_476 (O_476,N_19724,N_19627);
xnor UO_477 (O_477,N_19635,N_19852);
or UO_478 (O_478,N_19847,N_19720);
or UO_479 (O_479,N_19665,N_19995);
or UO_480 (O_480,N_19833,N_19815);
and UO_481 (O_481,N_19826,N_19891);
xnor UO_482 (O_482,N_19810,N_19736);
xnor UO_483 (O_483,N_19801,N_19888);
nor UO_484 (O_484,N_19761,N_19889);
or UO_485 (O_485,N_19968,N_19850);
nor UO_486 (O_486,N_19618,N_19991);
and UO_487 (O_487,N_19559,N_19724);
nand UO_488 (O_488,N_19654,N_19781);
and UO_489 (O_489,N_19872,N_19875);
nand UO_490 (O_490,N_19526,N_19849);
and UO_491 (O_491,N_19806,N_19954);
and UO_492 (O_492,N_19611,N_19876);
and UO_493 (O_493,N_19505,N_19666);
nand UO_494 (O_494,N_19766,N_19661);
xor UO_495 (O_495,N_19556,N_19624);
or UO_496 (O_496,N_19594,N_19715);
or UO_497 (O_497,N_19856,N_19608);
xor UO_498 (O_498,N_19661,N_19985);
xnor UO_499 (O_499,N_19871,N_19635);
nand UO_500 (O_500,N_19555,N_19639);
and UO_501 (O_501,N_19944,N_19647);
xnor UO_502 (O_502,N_19618,N_19901);
nand UO_503 (O_503,N_19952,N_19517);
and UO_504 (O_504,N_19596,N_19535);
nand UO_505 (O_505,N_19884,N_19960);
and UO_506 (O_506,N_19603,N_19796);
nand UO_507 (O_507,N_19882,N_19615);
nor UO_508 (O_508,N_19976,N_19902);
nor UO_509 (O_509,N_19933,N_19915);
nor UO_510 (O_510,N_19587,N_19618);
xnor UO_511 (O_511,N_19824,N_19540);
nand UO_512 (O_512,N_19706,N_19539);
nand UO_513 (O_513,N_19887,N_19914);
xnor UO_514 (O_514,N_19512,N_19588);
nor UO_515 (O_515,N_19709,N_19846);
nor UO_516 (O_516,N_19526,N_19754);
nand UO_517 (O_517,N_19741,N_19887);
or UO_518 (O_518,N_19827,N_19525);
or UO_519 (O_519,N_19612,N_19618);
xor UO_520 (O_520,N_19643,N_19946);
nor UO_521 (O_521,N_19832,N_19609);
xnor UO_522 (O_522,N_19687,N_19837);
xnor UO_523 (O_523,N_19542,N_19877);
and UO_524 (O_524,N_19776,N_19731);
xor UO_525 (O_525,N_19656,N_19784);
xnor UO_526 (O_526,N_19564,N_19954);
nand UO_527 (O_527,N_19963,N_19749);
or UO_528 (O_528,N_19733,N_19549);
xor UO_529 (O_529,N_19997,N_19711);
xor UO_530 (O_530,N_19644,N_19683);
xnor UO_531 (O_531,N_19833,N_19676);
nand UO_532 (O_532,N_19990,N_19521);
and UO_533 (O_533,N_19899,N_19559);
xor UO_534 (O_534,N_19694,N_19747);
xnor UO_535 (O_535,N_19931,N_19831);
nand UO_536 (O_536,N_19554,N_19517);
nand UO_537 (O_537,N_19715,N_19626);
and UO_538 (O_538,N_19792,N_19548);
or UO_539 (O_539,N_19743,N_19793);
xnor UO_540 (O_540,N_19766,N_19956);
or UO_541 (O_541,N_19637,N_19971);
nand UO_542 (O_542,N_19718,N_19759);
nand UO_543 (O_543,N_19949,N_19999);
and UO_544 (O_544,N_19587,N_19523);
nand UO_545 (O_545,N_19774,N_19694);
xnor UO_546 (O_546,N_19743,N_19992);
nor UO_547 (O_547,N_19642,N_19618);
nand UO_548 (O_548,N_19581,N_19645);
nand UO_549 (O_549,N_19880,N_19792);
xor UO_550 (O_550,N_19601,N_19569);
nand UO_551 (O_551,N_19870,N_19804);
nor UO_552 (O_552,N_19801,N_19940);
xor UO_553 (O_553,N_19507,N_19873);
xnor UO_554 (O_554,N_19805,N_19549);
or UO_555 (O_555,N_19903,N_19680);
nor UO_556 (O_556,N_19821,N_19720);
and UO_557 (O_557,N_19824,N_19820);
nand UO_558 (O_558,N_19521,N_19786);
xor UO_559 (O_559,N_19859,N_19565);
nor UO_560 (O_560,N_19772,N_19900);
nor UO_561 (O_561,N_19653,N_19770);
and UO_562 (O_562,N_19770,N_19908);
nor UO_563 (O_563,N_19513,N_19640);
xor UO_564 (O_564,N_19936,N_19998);
nand UO_565 (O_565,N_19772,N_19940);
nand UO_566 (O_566,N_19974,N_19714);
nand UO_567 (O_567,N_19805,N_19569);
nor UO_568 (O_568,N_19885,N_19834);
and UO_569 (O_569,N_19921,N_19963);
nand UO_570 (O_570,N_19888,N_19995);
xnor UO_571 (O_571,N_19577,N_19744);
or UO_572 (O_572,N_19625,N_19836);
or UO_573 (O_573,N_19685,N_19730);
nor UO_574 (O_574,N_19993,N_19891);
and UO_575 (O_575,N_19511,N_19752);
xor UO_576 (O_576,N_19637,N_19853);
and UO_577 (O_577,N_19986,N_19540);
or UO_578 (O_578,N_19806,N_19813);
nand UO_579 (O_579,N_19625,N_19960);
or UO_580 (O_580,N_19639,N_19500);
nand UO_581 (O_581,N_19785,N_19988);
and UO_582 (O_582,N_19629,N_19976);
nor UO_583 (O_583,N_19959,N_19698);
and UO_584 (O_584,N_19725,N_19656);
nand UO_585 (O_585,N_19587,N_19892);
xor UO_586 (O_586,N_19885,N_19563);
and UO_587 (O_587,N_19848,N_19629);
nand UO_588 (O_588,N_19753,N_19569);
nand UO_589 (O_589,N_19839,N_19897);
and UO_590 (O_590,N_19802,N_19760);
and UO_591 (O_591,N_19548,N_19882);
and UO_592 (O_592,N_19711,N_19512);
and UO_593 (O_593,N_19679,N_19726);
or UO_594 (O_594,N_19697,N_19681);
and UO_595 (O_595,N_19518,N_19585);
nor UO_596 (O_596,N_19793,N_19822);
and UO_597 (O_597,N_19905,N_19723);
xnor UO_598 (O_598,N_19960,N_19986);
xor UO_599 (O_599,N_19720,N_19500);
nand UO_600 (O_600,N_19709,N_19952);
xor UO_601 (O_601,N_19598,N_19889);
xor UO_602 (O_602,N_19838,N_19721);
and UO_603 (O_603,N_19876,N_19680);
or UO_604 (O_604,N_19859,N_19867);
nand UO_605 (O_605,N_19585,N_19959);
nor UO_606 (O_606,N_19612,N_19820);
or UO_607 (O_607,N_19882,N_19522);
nor UO_608 (O_608,N_19950,N_19881);
and UO_609 (O_609,N_19692,N_19912);
nand UO_610 (O_610,N_19962,N_19662);
or UO_611 (O_611,N_19988,N_19665);
and UO_612 (O_612,N_19554,N_19512);
nand UO_613 (O_613,N_19524,N_19723);
xor UO_614 (O_614,N_19829,N_19637);
nor UO_615 (O_615,N_19992,N_19961);
and UO_616 (O_616,N_19701,N_19524);
or UO_617 (O_617,N_19946,N_19806);
xnor UO_618 (O_618,N_19963,N_19781);
nand UO_619 (O_619,N_19623,N_19664);
xor UO_620 (O_620,N_19729,N_19775);
and UO_621 (O_621,N_19899,N_19756);
nand UO_622 (O_622,N_19536,N_19612);
xor UO_623 (O_623,N_19748,N_19996);
xnor UO_624 (O_624,N_19670,N_19889);
xnor UO_625 (O_625,N_19731,N_19678);
xnor UO_626 (O_626,N_19867,N_19669);
xor UO_627 (O_627,N_19522,N_19702);
or UO_628 (O_628,N_19803,N_19594);
and UO_629 (O_629,N_19784,N_19578);
or UO_630 (O_630,N_19735,N_19982);
nor UO_631 (O_631,N_19532,N_19542);
and UO_632 (O_632,N_19959,N_19623);
nand UO_633 (O_633,N_19640,N_19679);
nor UO_634 (O_634,N_19804,N_19664);
nor UO_635 (O_635,N_19765,N_19760);
or UO_636 (O_636,N_19927,N_19922);
and UO_637 (O_637,N_19895,N_19726);
or UO_638 (O_638,N_19589,N_19769);
nand UO_639 (O_639,N_19730,N_19809);
nand UO_640 (O_640,N_19552,N_19576);
or UO_641 (O_641,N_19779,N_19590);
nor UO_642 (O_642,N_19741,N_19598);
nand UO_643 (O_643,N_19519,N_19750);
xor UO_644 (O_644,N_19971,N_19711);
nand UO_645 (O_645,N_19603,N_19731);
nand UO_646 (O_646,N_19956,N_19951);
nand UO_647 (O_647,N_19604,N_19933);
nor UO_648 (O_648,N_19535,N_19563);
nand UO_649 (O_649,N_19944,N_19879);
nor UO_650 (O_650,N_19659,N_19810);
and UO_651 (O_651,N_19648,N_19780);
or UO_652 (O_652,N_19558,N_19578);
or UO_653 (O_653,N_19915,N_19614);
xor UO_654 (O_654,N_19708,N_19816);
and UO_655 (O_655,N_19646,N_19506);
xnor UO_656 (O_656,N_19825,N_19961);
and UO_657 (O_657,N_19844,N_19516);
xnor UO_658 (O_658,N_19904,N_19724);
nor UO_659 (O_659,N_19601,N_19689);
and UO_660 (O_660,N_19945,N_19807);
nand UO_661 (O_661,N_19910,N_19776);
or UO_662 (O_662,N_19817,N_19586);
or UO_663 (O_663,N_19674,N_19556);
nand UO_664 (O_664,N_19572,N_19950);
nand UO_665 (O_665,N_19974,N_19720);
or UO_666 (O_666,N_19574,N_19815);
or UO_667 (O_667,N_19669,N_19719);
and UO_668 (O_668,N_19762,N_19755);
and UO_669 (O_669,N_19794,N_19593);
nand UO_670 (O_670,N_19786,N_19933);
xor UO_671 (O_671,N_19670,N_19809);
and UO_672 (O_672,N_19740,N_19871);
nor UO_673 (O_673,N_19606,N_19690);
nor UO_674 (O_674,N_19649,N_19815);
nand UO_675 (O_675,N_19541,N_19733);
nand UO_676 (O_676,N_19573,N_19823);
nand UO_677 (O_677,N_19577,N_19630);
or UO_678 (O_678,N_19617,N_19972);
xnor UO_679 (O_679,N_19528,N_19643);
or UO_680 (O_680,N_19785,N_19947);
and UO_681 (O_681,N_19772,N_19934);
nand UO_682 (O_682,N_19591,N_19604);
nand UO_683 (O_683,N_19767,N_19979);
and UO_684 (O_684,N_19716,N_19888);
nand UO_685 (O_685,N_19883,N_19855);
and UO_686 (O_686,N_19657,N_19823);
or UO_687 (O_687,N_19632,N_19796);
nor UO_688 (O_688,N_19878,N_19596);
xnor UO_689 (O_689,N_19753,N_19960);
or UO_690 (O_690,N_19789,N_19777);
xnor UO_691 (O_691,N_19838,N_19705);
xor UO_692 (O_692,N_19873,N_19885);
xnor UO_693 (O_693,N_19947,N_19635);
or UO_694 (O_694,N_19750,N_19715);
or UO_695 (O_695,N_19750,N_19962);
nor UO_696 (O_696,N_19973,N_19729);
nor UO_697 (O_697,N_19591,N_19846);
and UO_698 (O_698,N_19558,N_19859);
and UO_699 (O_699,N_19805,N_19922);
and UO_700 (O_700,N_19579,N_19919);
and UO_701 (O_701,N_19998,N_19625);
nand UO_702 (O_702,N_19836,N_19707);
xnor UO_703 (O_703,N_19945,N_19639);
nor UO_704 (O_704,N_19971,N_19796);
nor UO_705 (O_705,N_19621,N_19583);
xnor UO_706 (O_706,N_19677,N_19758);
and UO_707 (O_707,N_19883,N_19721);
nor UO_708 (O_708,N_19878,N_19714);
nand UO_709 (O_709,N_19683,N_19873);
nor UO_710 (O_710,N_19616,N_19663);
or UO_711 (O_711,N_19661,N_19857);
xor UO_712 (O_712,N_19769,N_19923);
and UO_713 (O_713,N_19783,N_19734);
or UO_714 (O_714,N_19657,N_19574);
nand UO_715 (O_715,N_19945,N_19795);
nor UO_716 (O_716,N_19889,N_19847);
nor UO_717 (O_717,N_19960,N_19897);
xnor UO_718 (O_718,N_19803,N_19816);
xor UO_719 (O_719,N_19600,N_19614);
nand UO_720 (O_720,N_19749,N_19950);
and UO_721 (O_721,N_19856,N_19936);
nor UO_722 (O_722,N_19996,N_19736);
xor UO_723 (O_723,N_19731,N_19526);
nor UO_724 (O_724,N_19568,N_19974);
xnor UO_725 (O_725,N_19790,N_19976);
nand UO_726 (O_726,N_19619,N_19919);
and UO_727 (O_727,N_19734,N_19653);
xor UO_728 (O_728,N_19830,N_19757);
and UO_729 (O_729,N_19729,N_19728);
nand UO_730 (O_730,N_19559,N_19598);
nor UO_731 (O_731,N_19561,N_19695);
nor UO_732 (O_732,N_19859,N_19681);
nor UO_733 (O_733,N_19766,N_19868);
or UO_734 (O_734,N_19648,N_19984);
xnor UO_735 (O_735,N_19927,N_19523);
xnor UO_736 (O_736,N_19940,N_19943);
xor UO_737 (O_737,N_19512,N_19678);
and UO_738 (O_738,N_19670,N_19620);
or UO_739 (O_739,N_19609,N_19870);
or UO_740 (O_740,N_19711,N_19695);
and UO_741 (O_741,N_19703,N_19895);
nor UO_742 (O_742,N_19771,N_19762);
or UO_743 (O_743,N_19589,N_19576);
xnor UO_744 (O_744,N_19798,N_19828);
nor UO_745 (O_745,N_19892,N_19784);
xnor UO_746 (O_746,N_19563,N_19894);
nor UO_747 (O_747,N_19680,N_19987);
and UO_748 (O_748,N_19607,N_19889);
nor UO_749 (O_749,N_19740,N_19631);
nand UO_750 (O_750,N_19789,N_19990);
nand UO_751 (O_751,N_19935,N_19604);
xnor UO_752 (O_752,N_19879,N_19989);
nand UO_753 (O_753,N_19785,N_19878);
or UO_754 (O_754,N_19618,N_19860);
xor UO_755 (O_755,N_19640,N_19857);
xor UO_756 (O_756,N_19992,N_19900);
xnor UO_757 (O_757,N_19908,N_19565);
nand UO_758 (O_758,N_19652,N_19819);
nand UO_759 (O_759,N_19631,N_19809);
nor UO_760 (O_760,N_19998,N_19596);
nand UO_761 (O_761,N_19754,N_19671);
nor UO_762 (O_762,N_19575,N_19900);
and UO_763 (O_763,N_19610,N_19688);
nor UO_764 (O_764,N_19934,N_19930);
or UO_765 (O_765,N_19805,N_19911);
nand UO_766 (O_766,N_19972,N_19584);
or UO_767 (O_767,N_19647,N_19959);
xor UO_768 (O_768,N_19597,N_19629);
xor UO_769 (O_769,N_19874,N_19989);
or UO_770 (O_770,N_19596,N_19996);
and UO_771 (O_771,N_19986,N_19611);
and UO_772 (O_772,N_19858,N_19556);
or UO_773 (O_773,N_19863,N_19776);
or UO_774 (O_774,N_19803,N_19609);
nand UO_775 (O_775,N_19734,N_19637);
and UO_776 (O_776,N_19745,N_19503);
nor UO_777 (O_777,N_19830,N_19922);
and UO_778 (O_778,N_19953,N_19612);
or UO_779 (O_779,N_19819,N_19731);
xnor UO_780 (O_780,N_19558,N_19861);
nand UO_781 (O_781,N_19922,N_19758);
nor UO_782 (O_782,N_19879,N_19549);
or UO_783 (O_783,N_19903,N_19629);
or UO_784 (O_784,N_19976,N_19715);
nor UO_785 (O_785,N_19838,N_19809);
xnor UO_786 (O_786,N_19891,N_19665);
or UO_787 (O_787,N_19572,N_19868);
nor UO_788 (O_788,N_19543,N_19794);
or UO_789 (O_789,N_19622,N_19936);
or UO_790 (O_790,N_19522,N_19611);
and UO_791 (O_791,N_19632,N_19660);
nor UO_792 (O_792,N_19579,N_19690);
nor UO_793 (O_793,N_19806,N_19541);
or UO_794 (O_794,N_19817,N_19564);
xor UO_795 (O_795,N_19818,N_19565);
or UO_796 (O_796,N_19767,N_19778);
nand UO_797 (O_797,N_19897,N_19639);
or UO_798 (O_798,N_19936,N_19565);
xor UO_799 (O_799,N_19879,N_19638);
nor UO_800 (O_800,N_19642,N_19937);
xor UO_801 (O_801,N_19766,N_19916);
nor UO_802 (O_802,N_19840,N_19550);
nor UO_803 (O_803,N_19674,N_19536);
or UO_804 (O_804,N_19948,N_19752);
nor UO_805 (O_805,N_19562,N_19940);
and UO_806 (O_806,N_19752,N_19703);
and UO_807 (O_807,N_19755,N_19685);
nand UO_808 (O_808,N_19548,N_19654);
and UO_809 (O_809,N_19643,N_19905);
xnor UO_810 (O_810,N_19589,N_19727);
and UO_811 (O_811,N_19722,N_19986);
xnor UO_812 (O_812,N_19841,N_19534);
or UO_813 (O_813,N_19626,N_19687);
or UO_814 (O_814,N_19979,N_19517);
nand UO_815 (O_815,N_19616,N_19966);
nand UO_816 (O_816,N_19808,N_19829);
xor UO_817 (O_817,N_19541,N_19842);
xnor UO_818 (O_818,N_19843,N_19907);
and UO_819 (O_819,N_19605,N_19769);
and UO_820 (O_820,N_19694,N_19956);
xnor UO_821 (O_821,N_19639,N_19611);
nor UO_822 (O_822,N_19938,N_19622);
or UO_823 (O_823,N_19715,N_19969);
nor UO_824 (O_824,N_19521,N_19636);
nor UO_825 (O_825,N_19786,N_19913);
nor UO_826 (O_826,N_19671,N_19922);
and UO_827 (O_827,N_19673,N_19776);
xnor UO_828 (O_828,N_19947,N_19985);
nor UO_829 (O_829,N_19996,N_19912);
and UO_830 (O_830,N_19545,N_19990);
xor UO_831 (O_831,N_19726,N_19938);
nor UO_832 (O_832,N_19640,N_19646);
xnor UO_833 (O_833,N_19839,N_19961);
or UO_834 (O_834,N_19850,N_19694);
and UO_835 (O_835,N_19760,N_19778);
nor UO_836 (O_836,N_19571,N_19733);
nand UO_837 (O_837,N_19762,N_19569);
nand UO_838 (O_838,N_19552,N_19924);
xor UO_839 (O_839,N_19586,N_19715);
or UO_840 (O_840,N_19818,N_19657);
nand UO_841 (O_841,N_19991,N_19547);
and UO_842 (O_842,N_19654,N_19712);
nand UO_843 (O_843,N_19934,N_19839);
nor UO_844 (O_844,N_19771,N_19732);
xnor UO_845 (O_845,N_19560,N_19705);
or UO_846 (O_846,N_19740,N_19613);
or UO_847 (O_847,N_19656,N_19515);
nor UO_848 (O_848,N_19685,N_19701);
xor UO_849 (O_849,N_19878,N_19851);
xor UO_850 (O_850,N_19699,N_19536);
and UO_851 (O_851,N_19941,N_19585);
nand UO_852 (O_852,N_19635,N_19942);
nor UO_853 (O_853,N_19520,N_19773);
nand UO_854 (O_854,N_19632,N_19738);
xor UO_855 (O_855,N_19937,N_19756);
and UO_856 (O_856,N_19817,N_19835);
nand UO_857 (O_857,N_19648,N_19691);
nand UO_858 (O_858,N_19732,N_19879);
and UO_859 (O_859,N_19694,N_19895);
nor UO_860 (O_860,N_19873,N_19898);
nor UO_861 (O_861,N_19815,N_19660);
or UO_862 (O_862,N_19751,N_19860);
nand UO_863 (O_863,N_19708,N_19796);
or UO_864 (O_864,N_19840,N_19970);
xnor UO_865 (O_865,N_19935,N_19796);
nand UO_866 (O_866,N_19612,N_19573);
xor UO_867 (O_867,N_19947,N_19979);
xnor UO_868 (O_868,N_19559,N_19699);
xor UO_869 (O_869,N_19912,N_19918);
or UO_870 (O_870,N_19999,N_19740);
and UO_871 (O_871,N_19898,N_19847);
nand UO_872 (O_872,N_19602,N_19756);
nor UO_873 (O_873,N_19779,N_19960);
and UO_874 (O_874,N_19847,N_19553);
nand UO_875 (O_875,N_19660,N_19652);
xnor UO_876 (O_876,N_19567,N_19641);
nor UO_877 (O_877,N_19806,N_19783);
and UO_878 (O_878,N_19904,N_19862);
xnor UO_879 (O_879,N_19777,N_19526);
xnor UO_880 (O_880,N_19625,N_19701);
nor UO_881 (O_881,N_19518,N_19983);
or UO_882 (O_882,N_19516,N_19862);
xnor UO_883 (O_883,N_19930,N_19517);
or UO_884 (O_884,N_19882,N_19815);
nor UO_885 (O_885,N_19680,N_19952);
xnor UO_886 (O_886,N_19892,N_19739);
nor UO_887 (O_887,N_19844,N_19993);
and UO_888 (O_888,N_19582,N_19714);
nor UO_889 (O_889,N_19959,N_19637);
and UO_890 (O_890,N_19809,N_19813);
nand UO_891 (O_891,N_19543,N_19595);
and UO_892 (O_892,N_19946,N_19845);
xnor UO_893 (O_893,N_19783,N_19744);
xnor UO_894 (O_894,N_19984,N_19624);
or UO_895 (O_895,N_19911,N_19562);
or UO_896 (O_896,N_19556,N_19831);
and UO_897 (O_897,N_19970,N_19879);
xnor UO_898 (O_898,N_19569,N_19642);
or UO_899 (O_899,N_19501,N_19656);
nor UO_900 (O_900,N_19932,N_19819);
nor UO_901 (O_901,N_19811,N_19631);
and UO_902 (O_902,N_19966,N_19503);
or UO_903 (O_903,N_19944,N_19938);
or UO_904 (O_904,N_19694,N_19599);
nand UO_905 (O_905,N_19934,N_19692);
nor UO_906 (O_906,N_19666,N_19972);
nor UO_907 (O_907,N_19681,N_19949);
nor UO_908 (O_908,N_19773,N_19516);
xnor UO_909 (O_909,N_19983,N_19894);
nor UO_910 (O_910,N_19813,N_19705);
or UO_911 (O_911,N_19504,N_19627);
or UO_912 (O_912,N_19916,N_19987);
or UO_913 (O_913,N_19776,N_19767);
and UO_914 (O_914,N_19760,N_19616);
xnor UO_915 (O_915,N_19705,N_19520);
nand UO_916 (O_916,N_19664,N_19609);
nor UO_917 (O_917,N_19590,N_19524);
xnor UO_918 (O_918,N_19601,N_19705);
xor UO_919 (O_919,N_19554,N_19843);
and UO_920 (O_920,N_19791,N_19939);
xor UO_921 (O_921,N_19698,N_19517);
and UO_922 (O_922,N_19643,N_19684);
nand UO_923 (O_923,N_19678,N_19734);
and UO_924 (O_924,N_19910,N_19889);
or UO_925 (O_925,N_19615,N_19871);
nand UO_926 (O_926,N_19615,N_19617);
xnor UO_927 (O_927,N_19968,N_19756);
nor UO_928 (O_928,N_19556,N_19500);
nand UO_929 (O_929,N_19777,N_19872);
xor UO_930 (O_930,N_19567,N_19786);
xor UO_931 (O_931,N_19647,N_19519);
nor UO_932 (O_932,N_19941,N_19667);
nand UO_933 (O_933,N_19932,N_19851);
or UO_934 (O_934,N_19862,N_19590);
nor UO_935 (O_935,N_19559,N_19833);
nand UO_936 (O_936,N_19771,N_19863);
nand UO_937 (O_937,N_19544,N_19791);
nor UO_938 (O_938,N_19589,N_19902);
and UO_939 (O_939,N_19658,N_19848);
nor UO_940 (O_940,N_19889,N_19985);
and UO_941 (O_941,N_19737,N_19963);
xnor UO_942 (O_942,N_19973,N_19816);
nand UO_943 (O_943,N_19594,N_19879);
or UO_944 (O_944,N_19786,N_19810);
nor UO_945 (O_945,N_19664,N_19691);
and UO_946 (O_946,N_19951,N_19878);
or UO_947 (O_947,N_19721,N_19667);
xor UO_948 (O_948,N_19588,N_19823);
or UO_949 (O_949,N_19818,N_19762);
or UO_950 (O_950,N_19523,N_19804);
nor UO_951 (O_951,N_19574,N_19874);
xnor UO_952 (O_952,N_19678,N_19527);
and UO_953 (O_953,N_19862,N_19744);
or UO_954 (O_954,N_19706,N_19563);
and UO_955 (O_955,N_19874,N_19525);
nor UO_956 (O_956,N_19832,N_19866);
xnor UO_957 (O_957,N_19567,N_19940);
nand UO_958 (O_958,N_19601,N_19908);
nor UO_959 (O_959,N_19740,N_19721);
or UO_960 (O_960,N_19553,N_19617);
nand UO_961 (O_961,N_19758,N_19689);
or UO_962 (O_962,N_19851,N_19550);
or UO_963 (O_963,N_19576,N_19973);
or UO_964 (O_964,N_19754,N_19635);
or UO_965 (O_965,N_19971,N_19705);
nor UO_966 (O_966,N_19965,N_19848);
or UO_967 (O_967,N_19747,N_19753);
or UO_968 (O_968,N_19612,N_19806);
nor UO_969 (O_969,N_19756,N_19522);
nor UO_970 (O_970,N_19978,N_19570);
or UO_971 (O_971,N_19958,N_19844);
or UO_972 (O_972,N_19680,N_19602);
or UO_973 (O_973,N_19734,N_19959);
or UO_974 (O_974,N_19857,N_19789);
or UO_975 (O_975,N_19601,N_19653);
nand UO_976 (O_976,N_19608,N_19907);
xnor UO_977 (O_977,N_19668,N_19566);
xor UO_978 (O_978,N_19513,N_19786);
or UO_979 (O_979,N_19944,N_19950);
xnor UO_980 (O_980,N_19751,N_19953);
xnor UO_981 (O_981,N_19781,N_19630);
or UO_982 (O_982,N_19786,N_19551);
xnor UO_983 (O_983,N_19986,N_19633);
and UO_984 (O_984,N_19873,N_19934);
nor UO_985 (O_985,N_19893,N_19575);
nor UO_986 (O_986,N_19711,N_19506);
xnor UO_987 (O_987,N_19847,N_19879);
nand UO_988 (O_988,N_19563,N_19905);
nor UO_989 (O_989,N_19991,N_19726);
and UO_990 (O_990,N_19704,N_19683);
xor UO_991 (O_991,N_19573,N_19571);
and UO_992 (O_992,N_19960,N_19870);
nand UO_993 (O_993,N_19760,N_19663);
and UO_994 (O_994,N_19602,N_19501);
nand UO_995 (O_995,N_19591,N_19649);
and UO_996 (O_996,N_19789,N_19891);
nor UO_997 (O_997,N_19751,N_19740);
nor UO_998 (O_998,N_19903,N_19502);
nor UO_999 (O_999,N_19946,N_19656);
nor UO_1000 (O_1000,N_19856,N_19545);
or UO_1001 (O_1001,N_19690,N_19707);
nand UO_1002 (O_1002,N_19784,N_19875);
or UO_1003 (O_1003,N_19883,N_19538);
nand UO_1004 (O_1004,N_19609,N_19735);
xnor UO_1005 (O_1005,N_19663,N_19929);
nor UO_1006 (O_1006,N_19649,N_19803);
nand UO_1007 (O_1007,N_19715,N_19712);
xor UO_1008 (O_1008,N_19775,N_19516);
nor UO_1009 (O_1009,N_19574,N_19539);
nand UO_1010 (O_1010,N_19764,N_19516);
nand UO_1011 (O_1011,N_19831,N_19957);
nand UO_1012 (O_1012,N_19787,N_19634);
nand UO_1013 (O_1013,N_19815,N_19851);
nor UO_1014 (O_1014,N_19931,N_19752);
or UO_1015 (O_1015,N_19929,N_19664);
xnor UO_1016 (O_1016,N_19946,N_19943);
or UO_1017 (O_1017,N_19926,N_19634);
or UO_1018 (O_1018,N_19760,N_19661);
and UO_1019 (O_1019,N_19658,N_19524);
nand UO_1020 (O_1020,N_19936,N_19866);
and UO_1021 (O_1021,N_19543,N_19918);
or UO_1022 (O_1022,N_19556,N_19509);
or UO_1023 (O_1023,N_19677,N_19916);
nor UO_1024 (O_1024,N_19829,N_19507);
and UO_1025 (O_1025,N_19572,N_19508);
and UO_1026 (O_1026,N_19749,N_19983);
xor UO_1027 (O_1027,N_19705,N_19800);
nand UO_1028 (O_1028,N_19791,N_19585);
or UO_1029 (O_1029,N_19504,N_19802);
nand UO_1030 (O_1030,N_19864,N_19878);
or UO_1031 (O_1031,N_19773,N_19780);
or UO_1032 (O_1032,N_19797,N_19645);
and UO_1033 (O_1033,N_19611,N_19523);
nand UO_1034 (O_1034,N_19829,N_19589);
xor UO_1035 (O_1035,N_19965,N_19662);
nand UO_1036 (O_1036,N_19966,N_19868);
xnor UO_1037 (O_1037,N_19580,N_19901);
or UO_1038 (O_1038,N_19985,N_19795);
xnor UO_1039 (O_1039,N_19897,N_19725);
nand UO_1040 (O_1040,N_19842,N_19663);
or UO_1041 (O_1041,N_19565,N_19508);
and UO_1042 (O_1042,N_19833,N_19617);
xnor UO_1043 (O_1043,N_19953,N_19949);
nand UO_1044 (O_1044,N_19883,N_19769);
nor UO_1045 (O_1045,N_19898,N_19612);
xnor UO_1046 (O_1046,N_19837,N_19587);
or UO_1047 (O_1047,N_19823,N_19908);
nor UO_1048 (O_1048,N_19639,N_19904);
xnor UO_1049 (O_1049,N_19834,N_19546);
and UO_1050 (O_1050,N_19803,N_19794);
or UO_1051 (O_1051,N_19660,N_19742);
and UO_1052 (O_1052,N_19894,N_19577);
or UO_1053 (O_1053,N_19787,N_19738);
nor UO_1054 (O_1054,N_19501,N_19815);
and UO_1055 (O_1055,N_19547,N_19935);
and UO_1056 (O_1056,N_19693,N_19917);
nand UO_1057 (O_1057,N_19888,N_19565);
nand UO_1058 (O_1058,N_19563,N_19765);
and UO_1059 (O_1059,N_19853,N_19659);
or UO_1060 (O_1060,N_19716,N_19922);
or UO_1061 (O_1061,N_19744,N_19827);
and UO_1062 (O_1062,N_19989,N_19576);
or UO_1063 (O_1063,N_19577,N_19644);
nor UO_1064 (O_1064,N_19927,N_19810);
or UO_1065 (O_1065,N_19691,N_19516);
xor UO_1066 (O_1066,N_19618,N_19502);
and UO_1067 (O_1067,N_19877,N_19911);
or UO_1068 (O_1068,N_19653,N_19998);
xnor UO_1069 (O_1069,N_19899,N_19951);
xor UO_1070 (O_1070,N_19595,N_19985);
or UO_1071 (O_1071,N_19936,N_19568);
nor UO_1072 (O_1072,N_19732,N_19760);
nor UO_1073 (O_1073,N_19994,N_19526);
xnor UO_1074 (O_1074,N_19958,N_19833);
nor UO_1075 (O_1075,N_19668,N_19821);
or UO_1076 (O_1076,N_19736,N_19885);
and UO_1077 (O_1077,N_19739,N_19632);
xor UO_1078 (O_1078,N_19807,N_19888);
nor UO_1079 (O_1079,N_19566,N_19694);
and UO_1080 (O_1080,N_19920,N_19722);
nor UO_1081 (O_1081,N_19821,N_19845);
nand UO_1082 (O_1082,N_19902,N_19918);
nand UO_1083 (O_1083,N_19945,N_19925);
nor UO_1084 (O_1084,N_19896,N_19825);
xnor UO_1085 (O_1085,N_19735,N_19632);
and UO_1086 (O_1086,N_19675,N_19690);
nand UO_1087 (O_1087,N_19752,N_19926);
and UO_1088 (O_1088,N_19804,N_19806);
xnor UO_1089 (O_1089,N_19684,N_19504);
or UO_1090 (O_1090,N_19961,N_19942);
xnor UO_1091 (O_1091,N_19871,N_19641);
nand UO_1092 (O_1092,N_19975,N_19729);
or UO_1093 (O_1093,N_19744,N_19947);
nand UO_1094 (O_1094,N_19903,N_19515);
nor UO_1095 (O_1095,N_19658,N_19710);
nand UO_1096 (O_1096,N_19645,N_19885);
and UO_1097 (O_1097,N_19512,N_19672);
and UO_1098 (O_1098,N_19593,N_19857);
xor UO_1099 (O_1099,N_19539,N_19751);
xnor UO_1100 (O_1100,N_19698,N_19904);
nand UO_1101 (O_1101,N_19532,N_19855);
xor UO_1102 (O_1102,N_19983,N_19638);
nor UO_1103 (O_1103,N_19526,N_19652);
xor UO_1104 (O_1104,N_19827,N_19515);
and UO_1105 (O_1105,N_19976,N_19724);
and UO_1106 (O_1106,N_19859,N_19914);
and UO_1107 (O_1107,N_19763,N_19654);
and UO_1108 (O_1108,N_19946,N_19793);
nand UO_1109 (O_1109,N_19758,N_19597);
nor UO_1110 (O_1110,N_19522,N_19868);
nand UO_1111 (O_1111,N_19616,N_19747);
nor UO_1112 (O_1112,N_19632,N_19843);
and UO_1113 (O_1113,N_19705,N_19607);
or UO_1114 (O_1114,N_19608,N_19893);
nand UO_1115 (O_1115,N_19970,N_19774);
nor UO_1116 (O_1116,N_19698,N_19623);
and UO_1117 (O_1117,N_19880,N_19866);
or UO_1118 (O_1118,N_19611,N_19987);
or UO_1119 (O_1119,N_19883,N_19577);
nor UO_1120 (O_1120,N_19757,N_19630);
xor UO_1121 (O_1121,N_19869,N_19629);
nand UO_1122 (O_1122,N_19946,N_19964);
and UO_1123 (O_1123,N_19944,N_19660);
xor UO_1124 (O_1124,N_19578,N_19512);
nand UO_1125 (O_1125,N_19746,N_19709);
or UO_1126 (O_1126,N_19753,N_19693);
nand UO_1127 (O_1127,N_19690,N_19559);
and UO_1128 (O_1128,N_19920,N_19867);
nand UO_1129 (O_1129,N_19714,N_19981);
nor UO_1130 (O_1130,N_19753,N_19650);
or UO_1131 (O_1131,N_19733,N_19745);
or UO_1132 (O_1132,N_19537,N_19916);
nand UO_1133 (O_1133,N_19676,N_19620);
nor UO_1134 (O_1134,N_19917,N_19871);
xor UO_1135 (O_1135,N_19779,N_19629);
and UO_1136 (O_1136,N_19519,N_19515);
or UO_1137 (O_1137,N_19628,N_19854);
xnor UO_1138 (O_1138,N_19665,N_19700);
or UO_1139 (O_1139,N_19992,N_19956);
nand UO_1140 (O_1140,N_19933,N_19822);
or UO_1141 (O_1141,N_19864,N_19737);
and UO_1142 (O_1142,N_19562,N_19506);
or UO_1143 (O_1143,N_19704,N_19741);
or UO_1144 (O_1144,N_19823,N_19878);
and UO_1145 (O_1145,N_19827,N_19690);
or UO_1146 (O_1146,N_19515,N_19994);
or UO_1147 (O_1147,N_19747,N_19521);
and UO_1148 (O_1148,N_19831,N_19820);
xnor UO_1149 (O_1149,N_19943,N_19939);
xnor UO_1150 (O_1150,N_19904,N_19723);
xnor UO_1151 (O_1151,N_19932,N_19840);
nor UO_1152 (O_1152,N_19544,N_19555);
or UO_1153 (O_1153,N_19729,N_19677);
nor UO_1154 (O_1154,N_19720,N_19706);
nand UO_1155 (O_1155,N_19837,N_19936);
xor UO_1156 (O_1156,N_19678,N_19967);
xor UO_1157 (O_1157,N_19890,N_19620);
nand UO_1158 (O_1158,N_19985,N_19972);
nand UO_1159 (O_1159,N_19628,N_19932);
nand UO_1160 (O_1160,N_19618,N_19633);
nand UO_1161 (O_1161,N_19731,N_19843);
or UO_1162 (O_1162,N_19844,N_19850);
nor UO_1163 (O_1163,N_19672,N_19507);
and UO_1164 (O_1164,N_19951,N_19975);
nor UO_1165 (O_1165,N_19840,N_19592);
and UO_1166 (O_1166,N_19591,N_19865);
or UO_1167 (O_1167,N_19566,N_19789);
nor UO_1168 (O_1168,N_19706,N_19615);
nor UO_1169 (O_1169,N_19960,N_19626);
nand UO_1170 (O_1170,N_19883,N_19917);
xnor UO_1171 (O_1171,N_19573,N_19787);
nand UO_1172 (O_1172,N_19911,N_19638);
or UO_1173 (O_1173,N_19991,N_19560);
nand UO_1174 (O_1174,N_19896,N_19971);
xnor UO_1175 (O_1175,N_19804,N_19899);
nor UO_1176 (O_1176,N_19810,N_19835);
and UO_1177 (O_1177,N_19687,N_19754);
or UO_1178 (O_1178,N_19841,N_19678);
xor UO_1179 (O_1179,N_19964,N_19590);
xnor UO_1180 (O_1180,N_19724,N_19877);
nand UO_1181 (O_1181,N_19760,N_19630);
nor UO_1182 (O_1182,N_19885,N_19651);
nand UO_1183 (O_1183,N_19982,N_19946);
xor UO_1184 (O_1184,N_19854,N_19703);
and UO_1185 (O_1185,N_19890,N_19706);
or UO_1186 (O_1186,N_19602,N_19529);
and UO_1187 (O_1187,N_19830,N_19788);
or UO_1188 (O_1188,N_19503,N_19654);
or UO_1189 (O_1189,N_19807,N_19958);
or UO_1190 (O_1190,N_19989,N_19707);
and UO_1191 (O_1191,N_19962,N_19916);
nor UO_1192 (O_1192,N_19649,N_19858);
nand UO_1193 (O_1193,N_19653,N_19620);
nor UO_1194 (O_1194,N_19730,N_19966);
xor UO_1195 (O_1195,N_19720,N_19570);
or UO_1196 (O_1196,N_19807,N_19897);
and UO_1197 (O_1197,N_19716,N_19687);
nand UO_1198 (O_1198,N_19775,N_19914);
and UO_1199 (O_1199,N_19610,N_19802);
nor UO_1200 (O_1200,N_19801,N_19856);
or UO_1201 (O_1201,N_19726,N_19829);
and UO_1202 (O_1202,N_19765,N_19827);
and UO_1203 (O_1203,N_19850,N_19741);
or UO_1204 (O_1204,N_19718,N_19598);
xnor UO_1205 (O_1205,N_19677,N_19809);
xor UO_1206 (O_1206,N_19718,N_19707);
nand UO_1207 (O_1207,N_19851,N_19539);
and UO_1208 (O_1208,N_19892,N_19811);
nand UO_1209 (O_1209,N_19798,N_19674);
nor UO_1210 (O_1210,N_19903,N_19524);
and UO_1211 (O_1211,N_19883,N_19592);
nand UO_1212 (O_1212,N_19685,N_19945);
and UO_1213 (O_1213,N_19531,N_19621);
xor UO_1214 (O_1214,N_19522,N_19776);
and UO_1215 (O_1215,N_19963,N_19640);
xnor UO_1216 (O_1216,N_19805,N_19876);
nor UO_1217 (O_1217,N_19651,N_19980);
xnor UO_1218 (O_1218,N_19524,N_19829);
or UO_1219 (O_1219,N_19978,N_19877);
and UO_1220 (O_1220,N_19922,N_19935);
nor UO_1221 (O_1221,N_19569,N_19950);
xor UO_1222 (O_1222,N_19964,N_19907);
or UO_1223 (O_1223,N_19733,N_19743);
or UO_1224 (O_1224,N_19519,N_19858);
xor UO_1225 (O_1225,N_19883,N_19976);
nor UO_1226 (O_1226,N_19885,N_19815);
nor UO_1227 (O_1227,N_19647,N_19631);
and UO_1228 (O_1228,N_19515,N_19657);
or UO_1229 (O_1229,N_19802,N_19858);
nand UO_1230 (O_1230,N_19792,N_19737);
xor UO_1231 (O_1231,N_19804,N_19582);
nor UO_1232 (O_1232,N_19537,N_19755);
xnor UO_1233 (O_1233,N_19967,N_19666);
xnor UO_1234 (O_1234,N_19807,N_19995);
or UO_1235 (O_1235,N_19650,N_19817);
and UO_1236 (O_1236,N_19773,N_19969);
nor UO_1237 (O_1237,N_19681,N_19710);
or UO_1238 (O_1238,N_19519,N_19939);
xnor UO_1239 (O_1239,N_19639,N_19661);
nor UO_1240 (O_1240,N_19884,N_19714);
or UO_1241 (O_1241,N_19543,N_19697);
or UO_1242 (O_1242,N_19714,N_19525);
xor UO_1243 (O_1243,N_19923,N_19739);
xnor UO_1244 (O_1244,N_19512,N_19603);
xnor UO_1245 (O_1245,N_19639,N_19529);
and UO_1246 (O_1246,N_19506,N_19543);
xor UO_1247 (O_1247,N_19662,N_19931);
and UO_1248 (O_1248,N_19696,N_19961);
or UO_1249 (O_1249,N_19607,N_19847);
nor UO_1250 (O_1250,N_19906,N_19647);
or UO_1251 (O_1251,N_19981,N_19703);
nor UO_1252 (O_1252,N_19941,N_19819);
nand UO_1253 (O_1253,N_19530,N_19577);
xnor UO_1254 (O_1254,N_19985,N_19783);
nor UO_1255 (O_1255,N_19788,N_19558);
and UO_1256 (O_1256,N_19756,N_19539);
xor UO_1257 (O_1257,N_19969,N_19917);
nand UO_1258 (O_1258,N_19595,N_19969);
nand UO_1259 (O_1259,N_19895,N_19741);
or UO_1260 (O_1260,N_19648,N_19874);
and UO_1261 (O_1261,N_19633,N_19865);
nand UO_1262 (O_1262,N_19513,N_19583);
and UO_1263 (O_1263,N_19925,N_19649);
nor UO_1264 (O_1264,N_19668,N_19974);
nor UO_1265 (O_1265,N_19784,N_19550);
nand UO_1266 (O_1266,N_19674,N_19944);
nor UO_1267 (O_1267,N_19669,N_19991);
xor UO_1268 (O_1268,N_19786,N_19569);
nor UO_1269 (O_1269,N_19696,N_19990);
xor UO_1270 (O_1270,N_19626,N_19676);
nor UO_1271 (O_1271,N_19539,N_19581);
and UO_1272 (O_1272,N_19657,N_19547);
nor UO_1273 (O_1273,N_19902,N_19711);
xor UO_1274 (O_1274,N_19972,N_19561);
or UO_1275 (O_1275,N_19991,N_19555);
nor UO_1276 (O_1276,N_19750,N_19926);
or UO_1277 (O_1277,N_19903,N_19620);
and UO_1278 (O_1278,N_19707,N_19943);
nor UO_1279 (O_1279,N_19902,N_19735);
xor UO_1280 (O_1280,N_19844,N_19786);
and UO_1281 (O_1281,N_19561,N_19685);
and UO_1282 (O_1282,N_19850,N_19995);
and UO_1283 (O_1283,N_19845,N_19704);
and UO_1284 (O_1284,N_19592,N_19784);
nand UO_1285 (O_1285,N_19787,N_19773);
nand UO_1286 (O_1286,N_19550,N_19733);
nand UO_1287 (O_1287,N_19967,N_19517);
nand UO_1288 (O_1288,N_19691,N_19525);
and UO_1289 (O_1289,N_19617,N_19706);
or UO_1290 (O_1290,N_19623,N_19543);
xnor UO_1291 (O_1291,N_19760,N_19819);
or UO_1292 (O_1292,N_19915,N_19846);
or UO_1293 (O_1293,N_19747,N_19523);
and UO_1294 (O_1294,N_19942,N_19755);
and UO_1295 (O_1295,N_19956,N_19939);
or UO_1296 (O_1296,N_19811,N_19537);
xnor UO_1297 (O_1297,N_19581,N_19620);
and UO_1298 (O_1298,N_19512,N_19546);
nor UO_1299 (O_1299,N_19663,N_19970);
nor UO_1300 (O_1300,N_19912,N_19640);
nor UO_1301 (O_1301,N_19653,N_19739);
xnor UO_1302 (O_1302,N_19575,N_19616);
nand UO_1303 (O_1303,N_19991,N_19511);
xor UO_1304 (O_1304,N_19927,N_19970);
or UO_1305 (O_1305,N_19631,N_19797);
nor UO_1306 (O_1306,N_19640,N_19527);
nor UO_1307 (O_1307,N_19883,N_19781);
nor UO_1308 (O_1308,N_19900,N_19853);
xor UO_1309 (O_1309,N_19710,N_19952);
and UO_1310 (O_1310,N_19859,N_19707);
nor UO_1311 (O_1311,N_19532,N_19518);
nor UO_1312 (O_1312,N_19521,N_19536);
nand UO_1313 (O_1313,N_19657,N_19852);
xnor UO_1314 (O_1314,N_19902,N_19680);
and UO_1315 (O_1315,N_19849,N_19937);
nor UO_1316 (O_1316,N_19546,N_19531);
xnor UO_1317 (O_1317,N_19937,N_19873);
nor UO_1318 (O_1318,N_19734,N_19888);
or UO_1319 (O_1319,N_19525,N_19545);
or UO_1320 (O_1320,N_19939,N_19785);
nor UO_1321 (O_1321,N_19812,N_19643);
nand UO_1322 (O_1322,N_19573,N_19798);
nand UO_1323 (O_1323,N_19525,N_19790);
xor UO_1324 (O_1324,N_19681,N_19805);
nor UO_1325 (O_1325,N_19636,N_19656);
and UO_1326 (O_1326,N_19875,N_19827);
xor UO_1327 (O_1327,N_19756,N_19625);
nand UO_1328 (O_1328,N_19586,N_19584);
xnor UO_1329 (O_1329,N_19614,N_19714);
or UO_1330 (O_1330,N_19696,N_19972);
or UO_1331 (O_1331,N_19574,N_19684);
xnor UO_1332 (O_1332,N_19749,N_19517);
and UO_1333 (O_1333,N_19655,N_19748);
nor UO_1334 (O_1334,N_19684,N_19641);
xor UO_1335 (O_1335,N_19704,N_19517);
nand UO_1336 (O_1336,N_19963,N_19916);
xnor UO_1337 (O_1337,N_19502,N_19832);
or UO_1338 (O_1338,N_19533,N_19907);
nor UO_1339 (O_1339,N_19760,N_19761);
nor UO_1340 (O_1340,N_19805,N_19757);
and UO_1341 (O_1341,N_19864,N_19794);
or UO_1342 (O_1342,N_19926,N_19820);
xnor UO_1343 (O_1343,N_19772,N_19870);
nor UO_1344 (O_1344,N_19585,N_19762);
xor UO_1345 (O_1345,N_19595,N_19552);
xor UO_1346 (O_1346,N_19741,N_19988);
and UO_1347 (O_1347,N_19700,N_19967);
and UO_1348 (O_1348,N_19837,N_19689);
nor UO_1349 (O_1349,N_19506,N_19664);
and UO_1350 (O_1350,N_19994,N_19646);
nand UO_1351 (O_1351,N_19898,N_19751);
nand UO_1352 (O_1352,N_19551,N_19556);
and UO_1353 (O_1353,N_19646,N_19885);
or UO_1354 (O_1354,N_19742,N_19990);
xor UO_1355 (O_1355,N_19609,N_19601);
nor UO_1356 (O_1356,N_19897,N_19724);
nor UO_1357 (O_1357,N_19925,N_19786);
nor UO_1358 (O_1358,N_19596,N_19955);
nand UO_1359 (O_1359,N_19841,N_19565);
nand UO_1360 (O_1360,N_19687,N_19598);
xnor UO_1361 (O_1361,N_19983,N_19871);
or UO_1362 (O_1362,N_19503,N_19851);
or UO_1363 (O_1363,N_19718,N_19740);
and UO_1364 (O_1364,N_19749,N_19529);
and UO_1365 (O_1365,N_19827,N_19644);
nand UO_1366 (O_1366,N_19984,N_19674);
nor UO_1367 (O_1367,N_19833,N_19506);
nor UO_1368 (O_1368,N_19530,N_19688);
xor UO_1369 (O_1369,N_19703,N_19641);
and UO_1370 (O_1370,N_19792,N_19821);
nand UO_1371 (O_1371,N_19879,N_19927);
nand UO_1372 (O_1372,N_19969,N_19714);
nand UO_1373 (O_1373,N_19808,N_19940);
xnor UO_1374 (O_1374,N_19553,N_19918);
nor UO_1375 (O_1375,N_19584,N_19534);
and UO_1376 (O_1376,N_19538,N_19616);
xnor UO_1377 (O_1377,N_19784,N_19650);
nor UO_1378 (O_1378,N_19943,N_19836);
nand UO_1379 (O_1379,N_19644,N_19713);
xor UO_1380 (O_1380,N_19630,N_19817);
and UO_1381 (O_1381,N_19586,N_19957);
nor UO_1382 (O_1382,N_19825,N_19975);
xnor UO_1383 (O_1383,N_19984,N_19724);
nand UO_1384 (O_1384,N_19850,N_19626);
and UO_1385 (O_1385,N_19636,N_19548);
nor UO_1386 (O_1386,N_19986,N_19878);
and UO_1387 (O_1387,N_19523,N_19710);
nor UO_1388 (O_1388,N_19827,N_19992);
xor UO_1389 (O_1389,N_19839,N_19651);
xor UO_1390 (O_1390,N_19635,N_19652);
nor UO_1391 (O_1391,N_19756,N_19502);
or UO_1392 (O_1392,N_19893,N_19989);
and UO_1393 (O_1393,N_19777,N_19838);
nand UO_1394 (O_1394,N_19603,N_19506);
xor UO_1395 (O_1395,N_19557,N_19564);
nor UO_1396 (O_1396,N_19639,N_19618);
xor UO_1397 (O_1397,N_19840,N_19908);
or UO_1398 (O_1398,N_19783,N_19550);
and UO_1399 (O_1399,N_19890,N_19887);
or UO_1400 (O_1400,N_19828,N_19674);
nand UO_1401 (O_1401,N_19897,N_19926);
and UO_1402 (O_1402,N_19828,N_19667);
nand UO_1403 (O_1403,N_19810,N_19572);
xnor UO_1404 (O_1404,N_19610,N_19576);
xnor UO_1405 (O_1405,N_19501,N_19523);
xor UO_1406 (O_1406,N_19962,N_19912);
and UO_1407 (O_1407,N_19848,N_19829);
nor UO_1408 (O_1408,N_19588,N_19895);
nor UO_1409 (O_1409,N_19826,N_19507);
and UO_1410 (O_1410,N_19571,N_19603);
xnor UO_1411 (O_1411,N_19568,N_19832);
nand UO_1412 (O_1412,N_19863,N_19595);
xor UO_1413 (O_1413,N_19788,N_19786);
xor UO_1414 (O_1414,N_19748,N_19716);
and UO_1415 (O_1415,N_19726,N_19838);
nand UO_1416 (O_1416,N_19783,N_19729);
and UO_1417 (O_1417,N_19989,N_19749);
xnor UO_1418 (O_1418,N_19998,N_19690);
xnor UO_1419 (O_1419,N_19653,N_19977);
nand UO_1420 (O_1420,N_19921,N_19650);
and UO_1421 (O_1421,N_19604,N_19597);
and UO_1422 (O_1422,N_19931,N_19684);
nand UO_1423 (O_1423,N_19542,N_19566);
nor UO_1424 (O_1424,N_19894,N_19826);
xnor UO_1425 (O_1425,N_19553,N_19696);
nand UO_1426 (O_1426,N_19554,N_19513);
or UO_1427 (O_1427,N_19542,N_19528);
and UO_1428 (O_1428,N_19999,N_19861);
nor UO_1429 (O_1429,N_19922,N_19564);
nor UO_1430 (O_1430,N_19789,N_19702);
or UO_1431 (O_1431,N_19535,N_19865);
nor UO_1432 (O_1432,N_19858,N_19684);
nor UO_1433 (O_1433,N_19729,N_19618);
or UO_1434 (O_1434,N_19894,N_19661);
xor UO_1435 (O_1435,N_19742,N_19568);
nand UO_1436 (O_1436,N_19825,N_19818);
or UO_1437 (O_1437,N_19647,N_19502);
nand UO_1438 (O_1438,N_19603,N_19991);
or UO_1439 (O_1439,N_19699,N_19554);
nor UO_1440 (O_1440,N_19815,N_19888);
or UO_1441 (O_1441,N_19697,N_19649);
nor UO_1442 (O_1442,N_19602,N_19590);
nand UO_1443 (O_1443,N_19933,N_19983);
xnor UO_1444 (O_1444,N_19612,N_19954);
and UO_1445 (O_1445,N_19646,N_19678);
nor UO_1446 (O_1446,N_19887,N_19513);
nand UO_1447 (O_1447,N_19686,N_19728);
nand UO_1448 (O_1448,N_19938,N_19784);
xor UO_1449 (O_1449,N_19676,N_19813);
nand UO_1450 (O_1450,N_19726,N_19769);
and UO_1451 (O_1451,N_19822,N_19874);
or UO_1452 (O_1452,N_19693,N_19867);
nor UO_1453 (O_1453,N_19869,N_19819);
nand UO_1454 (O_1454,N_19812,N_19993);
xnor UO_1455 (O_1455,N_19612,N_19624);
or UO_1456 (O_1456,N_19857,N_19736);
and UO_1457 (O_1457,N_19834,N_19586);
xor UO_1458 (O_1458,N_19941,N_19569);
or UO_1459 (O_1459,N_19866,N_19679);
nor UO_1460 (O_1460,N_19620,N_19591);
or UO_1461 (O_1461,N_19619,N_19676);
or UO_1462 (O_1462,N_19648,N_19599);
nor UO_1463 (O_1463,N_19587,N_19874);
or UO_1464 (O_1464,N_19524,N_19599);
nor UO_1465 (O_1465,N_19508,N_19618);
nor UO_1466 (O_1466,N_19864,N_19607);
xnor UO_1467 (O_1467,N_19621,N_19607);
and UO_1468 (O_1468,N_19858,N_19507);
or UO_1469 (O_1469,N_19639,N_19562);
nor UO_1470 (O_1470,N_19693,N_19959);
nand UO_1471 (O_1471,N_19713,N_19629);
and UO_1472 (O_1472,N_19536,N_19644);
nor UO_1473 (O_1473,N_19961,N_19970);
nor UO_1474 (O_1474,N_19636,N_19760);
or UO_1475 (O_1475,N_19574,N_19681);
or UO_1476 (O_1476,N_19593,N_19723);
nor UO_1477 (O_1477,N_19949,N_19928);
or UO_1478 (O_1478,N_19579,N_19513);
xor UO_1479 (O_1479,N_19917,N_19973);
xnor UO_1480 (O_1480,N_19720,N_19959);
or UO_1481 (O_1481,N_19759,N_19810);
nand UO_1482 (O_1482,N_19634,N_19847);
or UO_1483 (O_1483,N_19571,N_19864);
or UO_1484 (O_1484,N_19511,N_19667);
or UO_1485 (O_1485,N_19752,N_19908);
nand UO_1486 (O_1486,N_19685,N_19712);
xor UO_1487 (O_1487,N_19611,N_19672);
nor UO_1488 (O_1488,N_19703,N_19980);
or UO_1489 (O_1489,N_19720,N_19609);
nand UO_1490 (O_1490,N_19530,N_19949);
nor UO_1491 (O_1491,N_19835,N_19523);
and UO_1492 (O_1492,N_19518,N_19592);
or UO_1493 (O_1493,N_19525,N_19689);
or UO_1494 (O_1494,N_19783,N_19538);
xnor UO_1495 (O_1495,N_19733,N_19525);
nand UO_1496 (O_1496,N_19834,N_19555);
xor UO_1497 (O_1497,N_19831,N_19554);
xnor UO_1498 (O_1498,N_19822,N_19962);
nor UO_1499 (O_1499,N_19673,N_19537);
or UO_1500 (O_1500,N_19552,N_19581);
or UO_1501 (O_1501,N_19966,N_19517);
xor UO_1502 (O_1502,N_19976,N_19692);
nand UO_1503 (O_1503,N_19815,N_19967);
xnor UO_1504 (O_1504,N_19628,N_19626);
xor UO_1505 (O_1505,N_19986,N_19664);
and UO_1506 (O_1506,N_19747,N_19817);
nand UO_1507 (O_1507,N_19965,N_19782);
xnor UO_1508 (O_1508,N_19921,N_19965);
or UO_1509 (O_1509,N_19842,N_19993);
xor UO_1510 (O_1510,N_19606,N_19712);
or UO_1511 (O_1511,N_19723,N_19913);
nand UO_1512 (O_1512,N_19554,N_19857);
nor UO_1513 (O_1513,N_19650,N_19935);
nor UO_1514 (O_1514,N_19568,N_19695);
nor UO_1515 (O_1515,N_19821,N_19951);
xor UO_1516 (O_1516,N_19569,N_19808);
nor UO_1517 (O_1517,N_19925,N_19878);
and UO_1518 (O_1518,N_19569,N_19947);
and UO_1519 (O_1519,N_19698,N_19571);
or UO_1520 (O_1520,N_19550,N_19785);
or UO_1521 (O_1521,N_19543,N_19585);
or UO_1522 (O_1522,N_19681,N_19808);
nand UO_1523 (O_1523,N_19814,N_19648);
or UO_1524 (O_1524,N_19570,N_19866);
nor UO_1525 (O_1525,N_19728,N_19672);
nand UO_1526 (O_1526,N_19846,N_19519);
nand UO_1527 (O_1527,N_19569,N_19674);
xnor UO_1528 (O_1528,N_19954,N_19896);
or UO_1529 (O_1529,N_19731,N_19877);
or UO_1530 (O_1530,N_19692,N_19972);
nand UO_1531 (O_1531,N_19848,N_19604);
and UO_1532 (O_1532,N_19537,N_19938);
or UO_1533 (O_1533,N_19904,N_19858);
xnor UO_1534 (O_1534,N_19684,N_19950);
and UO_1535 (O_1535,N_19709,N_19503);
nand UO_1536 (O_1536,N_19605,N_19756);
xor UO_1537 (O_1537,N_19518,N_19508);
xnor UO_1538 (O_1538,N_19529,N_19956);
and UO_1539 (O_1539,N_19943,N_19897);
nand UO_1540 (O_1540,N_19975,N_19562);
xnor UO_1541 (O_1541,N_19558,N_19502);
xnor UO_1542 (O_1542,N_19930,N_19545);
and UO_1543 (O_1543,N_19777,N_19602);
and UO_1544 (O_1544,N_19730,N_19614);
xor UO_1545 (O_1545,N_19532,N_19874);
and UO_1546 (O_1546,N_19564,N_19632);
xor UO_1547 (O_1547,N_19840,N_19683);
xor UO_1548 (O_1548,N_19872,N_19592);
nor UO_1549 (O_1549,N_19987,N_19969);
nor UO_1550 (O_1550,N_19890,N_19595);
and UO_1551 (O_1551,N_19564,N_19753);
or UO_1552 (O_1552,N_19718,N_19873);
nand UO_1553 (O_1553,N_19726,N_19559);
or UO_1554 (O_1554,N_19786,N_19746);
or UO_1555 (O_1555,N_19547,N_19568);
and UO_1556 (O_1556,N_19559,N_19795);
nor UO_1557 (O_1557,N_19719,N_19843);
and UO_1558 (O_1558,N_19794,N_19951);
nand UO_1559 (O_1559,N_19638,N_19660);
xor UO_1560 (O_1560,N_19975,N_19813);
nor UO_1561 (O_1561,N_19701,N_19843);
nor UO_1562 (O_1562,N_19615,N_19531);
and UO_1563 (O_1563,N_19691,N_19658);
or UO_1564 (O_1564,N_19548,N_19715);
xnor UO_1565 (O_1565,N_19933,N_19807);
nor UO_1566 (O_1566,N_19946,N_19791);
or UO_1567 (O_1567,N_19698,N_19504);
nand UO_1568 (O_1568,N_19502,N_19872);
xor UO_1569 (O_1569,N_19963,N_19931);
nor UO_1570 (O_1570,N_19954,N_19692);
xor UO_1571 (O_1571,N_19626,N_19747);
xor UO_1572 (O_1572,N_19538,N_19759);
and UO_1573 (O_1573,N_19541,N_19954);
and UO_1574 (O_1574,N_19520,N_19971);
or UO_1575 (O_1575,N_19810,N_19610);
xnor UO_1576 (O_1576,N_19919,N_19502);
or UO_1577 (O_1577,N_19923,N_19773);
and UO_1578 (O_1578,N_19729,N_19670);
xor UO_1579 (O_1579,N_19847,N_19828);
nor UO_1580 (O_1580,N_19989,N_19548);
xor UO_1581 (O_1581,N_19714,N_19856);
xnor UO_1582 (O_1582,N_19598,N_19880);
and UO_1583 (O_1583,N_19617,N_19547);
and UO_1584 (O_1584,N_19754,N_19972);
or UO_1585 (O_1585,N_19655,N_19944);
xor UO_1586 (O_1586,N_19998,N_19963);
nand UO_1587 (O_1587,N_19902,N_19529);
and UO_1588 (O_1588,N_19731,N_19711);
nor UO_1589 (O_1589,N_19727,N_19812);
nor UO_1590 (O_1590,N_19855,N_19813);
xnor UO_1591 (O_1591,N_19785,N_19668);
xnor UO_1592 (O_1592,N_19909,N_19898);
and UO_1593 (O_1593,N_19534,N_19993);
and UO_1594 (O_1594,N_19936,N_19992);
nor UO_1595 (O_1595,N_19691,N_19675);
xnor UO_1596 (O_1596,N_19882,N_19762);
xnor UO_1597 (O_1597,N_19859,N_19596);
or UO_1598 (O_1598,N_19804,N_19801);
and UO_1599 (O_1599,N_19764,N_19598);
nand UO_1600 (O_1600,N_19792,N_19772);
xor UO_1601 (O_1601,N_19830,N_19562);
nor UO_1602 (O_1602,N_19584,N_19802);
xnor UO_1603 (O_1603,N_19645,N_19941);
or UO_1604 (O_1604,N_19519,N_19641);
and UO_1605 (O_1605,N_19927,N_19989);
and UO_1606 (O_1606,N_19905,N_19709);
and UO_1607 (O_1607,N_19690,N_19667);
and UO_1608 (O_1608,N_19976,N_19708);
or UO_1609 (O_1609,N_19820,N_19507);
xnor UO_1610 (O_1610,N_19818,N_19732);
nor UO_1611 (O_1611,N_19673,N_19751);
nor UO_1612 (O_1612,N_19849,N_19768);
nor UO_1613 (O_1613,N_19919,N_19653);
or UO_1614 (O_1614,N_19623,N_19662);
or UO_1615 (O_1615,N_19975,N_19791);
nor UO_1616 (O_1616,N_19864,N_19770);
xor UO_1617 (O_1617,N_19667,N_19893);
and UO_1618 (O_1618,N_19702,N_19650);
nor UO_1619 (O_1619,N_19690,N_19907);
nand UO_1620 (O_1620,N_19676,N_19848);
nand UO_1621 (O_1621,N_19697,N_19865);
nor UO_1622 (O_1622,N_19784,N_19818);
xnor UO_1623 (O_1623,N_19689,N_19926);
xnor UO_1624 (O_1624,N_19945,N_19819);
nor UO_1625 (O_1625,N_19976,N_19807);
nor UO_1626 (O_1626,N_19784,N_19625);
nand UO_1627 (O_1627,N_19697,N_19657);
nand UO_1628 (O_1628,N_19646,N_19568);
and UO_1629 (O_1629,N_19973,N_19743);
xnor UO_1630 (O_1630,N_19580,N_19708);
nor UO_1631 (O_1631,N_19982,N_19625);
nor UO_1632 (O_1632,N_19552,N_19863);
nor UO_1633 (O_1633,N_19589,N_19547);
xnor UO_1634 (O_1634,N_19517,N_19874);
nor UO_1635 (O_1635,N_19895,N_19832);
nor UO_1636 (O_1636,N_19744,N_19864);
and UO_1637 (O_1637,N_19510,N_19873);
nor UO_1638 (O_1638,N_19880,N_19527);
and UO_1639 (O_1639,N_19952,N_19822);
nand UO_1640 (O_1640,N_19773,N_19856);
or UO_1641 (O_1641,N_19628,N_19665);
or UO_1642 (O_1642,N_19552,N_19870);
xor UO_1643 (O_1643,N_19811,N_19916);
nand UO_1644 (O_1644,N_19686,N_19613);
nand UO_1645 (O_1645,N_19980,N_19891);
nor UO_1646 (O_1646,N_19738,N_19673);
or UO_1647 (O_1647,N_19801,N_19598);
nand UO_1648 (O_1648,N_19896,N_19965);
and UO_1649 (O_1649,N_19575,N_19896);
xnor UO_1650 (O_1650,N_19833,N_19545);
xnor UO_1651 (O_1651,N_19711,N_19981);
and UO_1652 (O_1652,N_19994,N_19909);
and UO_1653 (O_1653,N_19825,N_19572);
and UO_1654 (O_1654,N_19844,N_19527);
nor UO_1655 (O_1655,N_19693,N_19708);
or UO_1656 (O_1656,N_19876,N_19509);
and UO_1657 (O_1657,N_19776,N_19867);
or UO_1658 (O_1658,N_19797,N_19829);
nor UO_1659 (O_1659,N_19803,N_19660);
and UO_1660 (O_1660,N_19834,N_19943);
or UO_1661 (O_1661,N_19771,N_19870);
nand UO_1662 (O_1662,N_19602,N_19632);
and UO_1663 (O_1663,N_19995,N_19749);
nand UO_1664 (O_1664,N_19796,N_19648);
nor UO_1665 (O_1665,N_19663,N_19520);
or UO_1666 (O_1666,N_19502,N_19658);
nor UO_1667 (O_1667,N_19843,N_19570);
xor UO_1668 (O_1668,N_19928,N_19811);
or UO_1669 (O_1669,N_19538,N_19897);
nand UO_1670 (O_1670,N_19942,N_19931);
nor UO_1671 (O_1671,N_19949,N_19515);
nand UO_1672 (O_1672,N_19838,N_19584);
or UO_1673 (O_1673,N_19527,N_19882);
xor UO_1674 (O_1674,N_19501,N_19906);
nand UO_1675 (O_1675,N_19611,N_19950);
xnor UO_1676 (O_1676,N_19910,N_19867);
or UO_1677 (O_1677,N_19798,N_19860);
xor UO_1678 (O_1678,N_19626,N_19989);
xnor UO_1679 (O_1679,N_19752,N_19759);
nand UO_1680 (O_1680,N_19832,N_19642);
nor UO_1681 (O_1681,N_19654,N_19631);
or UO_1682 (O_1682,N_19722,N_19852);
xor UO_1683 (O_1683,N_19576,N_19659);
and UO_1684 (O_1684,N_19907,N_19718);
nand UO_1685 (O_1685,N_19772,N_19586);
and UO_1686 (O_1686,N_19802,N_19873);
nor UO_1687 (O_1687,N_19535,N_19722);
nor UO_1688 (O_1688,N_19899,N_19660);
nand UO_1689 (O_1689,N_19502,N_19521);
xnor UO_1690 (O_1690,N_19988,N_19943);
xnor UO_1691 (O_1691,N_19607,N_19745);
or UO_1692 (O_1692,N_19959,N_19835);
nor UO_1693 (O_1693,N_19722,N_19620);
xor UO_1694 (O_1694,N_19659,N_19566);
nand UO_1695 (O_1695,N_19708,N_19804);
xor UO_1696 (O_1696,N_19531,N_19650);
nand UO_1697 (O_1697,N_19824,N_19846);
and UO_1698 (O_1698,N_19904,N_19707);
and UO_1699 (O_1699,N_19511,N_19664);
nor UO_1700 (O_1700,N_19692,N_19947);
nor UO_1701 (O_1701,N_19938,N_19544);
or UO_1702 (O_1702,N_19543,N_19673);
and UO_1703 (O_1703,N_19891,N_19715);
xor UO_1704 (O_1704,N_19548,N_19769);
xor UO_1705 (O_1705,N_19668,N_19926);
nor UO_1706 (O_1706,N_19604,N_19657);
and UO_1707 (O_1707,N_19974,N_19826);
or UO_1708 (O_1708,N_19635,N_19535);
and UO_1709 (O_1709,N_19842,N_19574);
xnor UO_1710 (O_1710,N_19870,N_19550);
nand UO_1711 (O_1711,N_19963,N_19619);
xnor UO_1712 (O_1712,N_19852,N_19959);
or UO_1713 (O_1713,N_19969,N_19644);
or UO_1714 (O_1714,N_19564,N_19750);
xor UO_1715 (O_1715,N_19896,N_19803);
and UO_1716 (O_1716,N_19873,N_19716);
and UO_1717 (O_1717,N_19725,N_19670);
nor UO_1718 (O_1718,N_19976,N_19809);
and UO_1719 (O_1719,N_19771,N_19792);
and UO_1720 (O_1720,N_19848,N_19825);
nor UO_1721 (O_1721,N_19980,N_19996);
and UO_1722 (O_1722,N_19877,N_19569);
and UO_1723 (O_1723,N_19767,N_19900);
or UO_1724 (O_1724,N_19746,N_19532);
nand UO_1725 (O_1725,N_19910,N_19536);
xnor UO_1726 (O_1726,N_19547,N_19810);
xor UO_1727 (O_1727,N_19557,N_19542);
nor UO_1728 (O_1728,N_19536,N_19532);
nand UO_1729 (O_1729,N_19598,N_19900);
nand UO_1730 (O_1730,N_19997,N_19767);
or UO_1731 (O_1731,N_19845,N_19945);
xnor UO_1732 (O_1732,N_19545,N_19818);
xor UO_1733 (O_1733,N_19721,N_19758);
and UO_1734 (O_1734,N_19553,N_19515);
or UO_1735 (O_1735,N_19537,N_19608);
and UO_1736 (O_1736,N_19630,N_19767);
and UO_1737 (O_1737,N_19671,N_19851);
and UO_1738 (O_1738,N_19818,N_19505);
xnor UO_1739 (O_1739,N_19936,N_19984);
xnor UO_1740 (O_1740,N_19564,N_19580);
nand UO_1741 (O_1741,N_19533,N_19835);
nor UO_1742 (O_1742,N_19858,N_19992);
xnor UO_1743 (O_1743,N_19685,N_19615);
or UO_1744 (O_1744,N_19634,N_19602);
nor UO_1745 (O_1745,N_19968,N_19678);
nand UO_1746 (O_1746,N_19661,N_19853);
nor UO_1747 (O_1747,N_19954,N_19670);
xor UO_1748 (O_1748,N_19599,N_19690);
nand UO_1749 (O_1749,N_19585,N_19743);
nand UO_1750 (O_1750,N_19981,N_19583);
nor UO_1751 (O_1751,N_19774,N_19936);
nor UO_1752 (O_1752,N_19521,N_19560);
nand UO_1753 (O_1753,N_19529,N_19829);
xor UO_1754 (O_1754,N_19676,N_19565);
xor UO_1755 (O_1755,N_19572,N_19559);
and UO_1756 (O_1756,N_19593,N_19810);
nor UO_1757 (O_1757,N_19708,N_19632);
nand UO_1758 (O_1758,N_19539,N_19502);
and UO_1759 (O_1759,N_19802,N_19918);
and UO_1760 (O_1760,N_19685,N_19585);
or UO_1761 (O_1761,N_19935,N_19568);
and UO_1762 (O_1762,N_19548,N_19925);
nand UO_1763 (O_1763,N_19608,N_19601);
nand UO_1764 (O_1764,N_19916,N_19526);
and UO_1765 (O_1765,N_19689,N_19868);
nor UO_1766 (O_1766,N_19993,N_19821);
nor UO_1767 (O_1767,N_19584,N_19525);
nand UO_1768 (O_1768,N_19735,N_19634);
nor UO_1769 (O_1769,N_19962,N_19800);
nand UO_1770 (O_1770,N_19517,N_19759);
nand UO_1771 (O_1771,N_19832,N_19859);
and UO_1772 (O_1772,N_19773,N_19504);
xnor UO_1773 (O_1773,N_19681,N_19522);
or UO_1774 (O_1774,N_19826,N_19589);
nor UO_1775 (O_1775,N_19962,N_19859);
or UO_1776 (O_1776,N_19638,N_19694);
nor UO_1777 (O_1777,N_19617,N_19841);
xnor UO_1778 (O_1778,N_19938,N_19670);
nor UO_1779 (O_1779,N_19965,N_19636);
nand UO_1780 (O_1780,N_19690,N_19700);
and UO_1781 (O_1781,N_19639,N_19984);
nor UO_1782 (O_1782,N_19854,N_19882);
xor UO_1783 (O_1783,N_19909,N_19794);
nand UO_1784 (O_1784,N_19940,N_19826);
or UO_1785 (O_1785,N_19737,N_19663);
nor UO_1786 (O_1786,N_19586,N_19735);
nand UO_1787 (O_1787,N_19612,N_19809);
nand UO_1788 (O_1788,N_19918,N_19794);
nand UO_1789 (O_1789,N_19812,N_19871);
nand UO_1790 (O_1790,N_19625,N_19711);
xor UO_1791 (O_1791,N_19541,N_19752);
nand UO_1792 (O_1792,N_19809,N_19704);
nor UO_1793 (O_1793,N_19870,N_19893);
xor UO_1794 (O_1794,N_19774,N_19687);
and UO_1795 (O_1795,N_19796,N_19657);
nor UO_1796 (O_1796,N_19906,N_19525);
xnor UO_1797 (O_1797,N_19880,N_19699);
nor UO_1798 (O_1798,N_19673,N_19803);
nand UO_1799 (O_1799,N_19995,N_19785);
nor UO_1800 (O_1800,N_19634,N_19961);
nand UO_1801 (O_1801,N_19768,N_19703);
nand UO_1802 (O_1802,N_19614,N_19902);
or UO_1803 (O_1803,N_19722,N_19885);
nor UO_1804 (O_1804,N_19986,N_19615);
xor UO_1805 (O_1805,N_19842,N_19973);
or UO_1806 (O_1806,N_19567,N_19566);
xnor UO_1807 (O_1807,N_19656,N_19860);
nand UO_1808 (O_1808,N_19731,N_19930);
nor UO_1809 (O_1809,N_19951,N_19921);
xnor UO_1810 (O_1810,N_19568,N_19620);
nand UO_1811 (O_1811,N_19964,N_19825);
xnor UO_1812 (O_1812,N_19767,N_19948);
and UO_1813 (O_1813,N_19662,N_19972);
nand UO_1814 (O_1814,N_19803,N_19842);
nor UO_1815 (O_1815,N_19617,N_19640);
or UO_1816 (O_1816,N_19803,N_19906);
nand UO_1817 (O_1817,N_19839,N_19594);
or UO_1818 (O_1818,N_19805,N_19694);
nor UO_1819 (O_1819,N_19625,N_19609);
xnor UO_1820 (O_1820,N_19662,N_19656);
or UO_1821 (O_1821,N_19942,N_19512);
nor UO_1822 (O_1822,N_19719,N_19606);
or UO_1823 (O_1823,N_19972,N_19947);
nand UO_1824 (O_1824,N_19677,N_19697);
or UO_1825 (O_1825,N_19762,N_19777);
nor UO_1826 (O_1826,N_19739,N_19979);
or UO_1827 (O_1827,N_19973,N_19600);
xor UO_1828 (O_1828,N_19722,N_19957);
xnor UO_1829 (O_1829,N_19872,N_19501);
xnor UO_1830 (O_1830,N_19552,N_19535);
nand UO_1831 (O_1831,N_19857,N_19951);
xnor UO_1832 (O_1832,N_19787,N_19873);
and UO_1833 (O_1833,N_19962,N_19864);
xnor UO_1834 (O_1834,N_19716,N_19957);
xor UO_1835 (O_1835,N_19739,N_19643);
nor UO_1836 (O_1836,N_19688,N_19581);
or UO_1837 (O_1837,N_19896,N_19789);
or UO_1838 (O_1838,N_19967,N_19611);
and UO_1839 (O_1839,N_19720,N_19993);
xnor UO_1840 (O_1840,N_19715,N_19541);
and UO_1841 (O_1841,N_19896,N_19557);
xor UO_1842 (O_1842,N_19570,N_19641);
xor UO_1843 (O_1843,N_19785,N_19982);
or UO_1844 (O_1844,N_19902,N_19583);
and UO_1845 (O_1845,N_19968,N_19943);
nor UO_1846 (O_1846,N_19655,N_19819);
nor UO_1847 (O_1847,N_19801,N_19724);
and UO_1848 (O_1848,N_19869,N_19584);
xor UO_1849 (O_1849,N_19860,N_19891);
nand UO_1850 (O_1850,N_19609,N_19852);
nor UO_1851 (O_1851,N_19915,N_19817);
and UO_1852 (O_1852,N_19881,N_19730);
or UO_1853 (O_1853,N_19679,N_19913);
nand UO_1854 (O_1854,N_19780,N_19686);
or UO_1855 (O_1855,N_19535,N_19772);
nand UO_1856 (O_1856,N_19999,N_19738);
xor UO_1857 (O_1857,N_19805,N_19700);
and UO_1858 (O_1858,N_19708,N_19837);
nor UO_1859 (O_1859,N_19600,N_19961);
xnor UO_1860 (O_1860,N_19530,N_19564);
and UO_1861 (O_1861,N_19642,N_19726);
or UO_1862 (O_1862,N_19842,N_19888);
nand UO_1863 (O_1863,N_19689,N_19680);
nand UO_1864 (O_1864,N_19723,N_19584);
and UO_1865 (O_1865,N_19974,N_19980);
and UO_1866 (O_1866,N_19878,N_19824);
xnor UO_1867 (O_1867,N_19890,N_19803);
nor UO_1868 (O_1868,N_19657,N_19920);
nand UO_1869 (O_1869,N_19855,N_19637);
nor UO_1870 (O_1870,N_19960,N_19789);
and UO_1871 (O_1871,N_19901,N_19724);
or UO_1872 (O_1872,N_19921,N_19930);
and UO_1873 (O_1873,N_19798,N_19641);
xnor UO_1874 (O_1874,N_19924,N_19719);
xor UO_1875 (O_1875,N_19850,N_19598);
nand UO_1876 (O_1876,N_19772,N_19500);
xor UO_1877 (O_1877,N_19645,N_19506);
and UO_1878 (O_1878,N_19921,N_19892);
or UO_1879 (O_1879,N_19998,N_19662);
xnor UO_1880 (O_1880,N_19608,N_19557);
xnor UO_1881 (O_1881,N_19884,N_19959);
nand UO_1882 (O_1882,N_19938,N_19941);
and UO_1883 (O_1883,N_19871,N_19649);
xor UO_1884 (O_1884,N_19845,N_19699);
or UO_1885 (O_1885,N_19819,N_19982);
xor UO_1886 (O_1886,N_19703,N_19957);
and UO_1887 (O_1887,N_19942,N_19937);
xnor UO_1888 (O_1888,N_19936,N_19765);
nor UO_1889 (O_1889,N_19532,N_19749);
nor UO_1890 (O_1890,N_19737,N_19988);
or UO_1891 (O_1891,N_19665,N_19602);
and UO_1892 (O_1892,N_19601,N_19555);
nor UO_1893 (O_1893,N_19755,N_19854);
xor UO_1894 (O_1894,N_19941,N_19720);
xor UO_1895 (O_1895,N_19528,N_19905);
xor UO_1896 (O_1896,N_19596,N_19939);
xnor UO_1897 (O_1897,N_19605,N_19886);
xor UO_1898 (O_1898,N_19548,N_19875);
and UO_1899 (O_1899,N_19600,N_19646);
nor UO_1900 (O_1900,N_19716,N_19502);
nand UO_1901 (O_1901,N_19994,N_19965);
and UO_1902 (O_1902,N_19850,N_19523);
nor UO_1903 (O_1903,N_19592,N_19873);
and UO_1904 (O_1904,N_19782,N_19581);
nand UO_1905 (O_1905,N_19873,N_19602);
and UO_1906 (O_1906,N_19962,N_19708);
and UO_1907 (O_1907,N_19914,N_19723);
nor UO_1908 (O_1908,N_19910,N_19563);
or UO_1909 (O_1909,N_19726,N_19634);
and UO_1910 (O_1910,N_19870,N_19587);
nor UO_1911 (O_1911,N_19794,N_19849);
nand UO_1912 (O_1912,N_19695,N_19746);
and UO_1913 (O_1913,N_19775,N_19875);
or UO_1914 (O_1914,N_19984,N_19908);
or UO_1915 (O_1915,N_19895,N_19502);
nor UO_1916 (O_1916,N_19913,N_19633);
or UO_1917 (O_1917,N_19574,N_19571);
and UO_1918 (O_1918,N_19866,N_19829);
xnor UO_1919 (O_1919,N_19790,N_19886);
nor UO_1920 (O_1920,N_19560,N_19541);
nor UO_1921 (O_1921,N_19771,N_19500);
nor UO_1922 (O_1922,N_19836,N_19739);
xor UO_1923 (O_1923,N_19677,N_19818);
nor UO_1924 (O_1924,N_19872,N_19572);
nand UO_1925 (O_1925,N_19625,N_19773);
nand UO_1926 (O_1926,N_19985,N_19557);
nor UO_1927 (O_1927,N_19860,N_19936);
and UO_1928 (O_1928,N_19522,N_19836);
and UO_1929 (O_1929,N_19562,N_19999);
nor UO_1930 (O_1930,N_19820,N_19997);
nand UO_1931 (O_1931,N_19999,N_19715);
nor UO_1932 (O_1932,N_19803,N_19538);
xor UO_1933 (O_1933,N_19691,N_19696);
and UO_1934 (O_1934,N_19775,N_19517);
and UO_1935 (O_1935,N_19758,N_19608);
nand UO_1936 (O_1936,N_19784,N_19785);
nor UO_1937 (O_1937,N_19633,N_19623);
nor UO_1938 (O_1938,N_19849,N_19619);
nor UO_1939 (O_1939,N_19600,N_19688);
nand UO_1940 (O_1940,N_19872,N_19892);
nor UO_1941 (O_1941,N_19543,N_19547);
xnor UO_1942 (O_1942,N_19587,N_19647);
nor UO_1943 (O_1943,N_19734,N_19957);
nor UO_1944 (O_1944,N_19822,N_19708);
or UO_1945 (O_1945,N_19615,N_19717);
nand UO_1946 (O_1946,N_19762,N_19796);
nor UO_1947 (O_1947,N_19828,N_19717);
or UO_1948 (O_1948,N_19773,N_19589);
and UO_1949 (O_1949,N_19982,N_19926);
nor UO_1950 (O_1950,N_19717,N_19523);
or UO_1951 (O_1951,N_19558,N_19728);
xnor UO_1952 (O_1952,N_19851,N_19619);
and UO_1953 (O_1953,N_19945,N_19794);
or UO_1954 (O_1954,N_19715,N_19805);
nand UO_1955 (O_1955,N_19855,N_19889);
xnor UO_1956 (O_1956,N_19694,N_19527);
xor UO_1957 (O_1957,N_19979,N_19564);
or UO_1958 (O_1958,N_19882,N_19802);
nand UO_1959 (O_1959,N_19714,N_19890);
or UO_1960 (O_1960,N_19744,N_19849);
nor UO_1961 (O_1961,N_19686,N_19515);
nor UO_1962 (O_1962,N_19740,N_19602);
nor UO_1963 (O_1963,N_19787,N_19760);
nand UO_1964 (O_1964,N_19753,N_19508);
xnor UO_1965 (O_1965,N_19854,N_19963);
xor UO_1966 (O_1966,N_19949,N_19529);
or UO_1967 (O_1967,N_19952,N_19755);
and UO_1968 (O_1968,N_19850,N_19639);
nand UO_1969 (O_1969,N_19907,N_19524);
xor UO_1970 (O_1970,N_19626,N_19756);
and UO_1971 (O_1971,N_19592,N_19554);
and UO_1972 (O_1972,N_19824,N_19583);
nor UO_1973 (O_1973,N_19831,N_19965);
and UO_1974 (O_1974,N_19988,N_19568);
xor UO_1975 (O_1975,N_19995,N_19823);
nor UO_1976 (O_1976,N_19810,N_19656);
and UO_1977 (O_1977,N_19562,N_19785);
and UO_1978 (O_1978,N_19733,N_19984);
xor UO_1979 (O_1979,N_19980,N_19825);
nand UO_1980 (O_1980,N_19808,N_19989);
xor UO_1981 (O_1981,N_19683,N_19846);
xor UO_1982 (O_1982,N_19609,N_19687);
or UO_1983 (O_1983,N_19795,N_19554);
nand UO_1984 (O_1984,N_19655,N_19918);
and UO_1985 (O_1985,N_19951,N_19939);
and UO_1986 (O_1986,N_19502,N_19525);
nand UO_1987 (O_1987,N_19865,N_19705);
nand UO_1988 (O_1988,N_19868,N_19667);
nand UO_1989 (O_1989,N_19745,N_19752);
or UO_1990 (O_1990,N_19915,N_19921);
nand UO_1991 (O_1991,N_19832,N_19995);
xor UO_1992 (O_1992,N_19745,N_19633);
xor UO_1993 (O_1993,N_19738,N_19558);
xnor UO_1994 (O_1994,N_19722,N_19897);
xor UO_1995 (O_1995,N_19998,N_19788);
nand UO_1996 (O_1996,N_19832,N_19575);
nand UO_1997 (O_1997,N_19953,N_19929);
nand UO_1998 (O_1998,N_19882,N_19724);
or UO_1999 (O_1999,N_19512,N_19872);
and UO_2000 (O_2000,N_19961,N_19647);
nand UO_2001 (O_2001,N_19770,N_19764);
nand UO_2002 (O_2002,N_19973,N_19938);
nand UO_2003 (O_2003,N_19620,N_19572);
and UO_2004 (O_2004,N_19833,N_19556);
or UO_2005 (O_2005,N_19668,N_19697);
xnor UO_2006 (O_2006,N_19635,N_19530);
nand UO_2007 (O_2007,N_19554,N_19616);
xnor UO_2008 (O_2008,N_19640,N_19685);
nand UO_2009 (O_2009,N_19814,N_19864);
or UO_2010 (O_2010,N_19681,N_19848);
or UO_2011 (O_2011,N_19700,N_19756);
or UO_2012 (O_2012,N_19700,N_19936);
nand UO_2013 (O_2013,N_19853,N_19851);
nor UO_2014 (O_2014,N_19799,N_19995);
xnor UO_2015 (O_2015,N_19559,N_19610);
xor UO_2016 (O_2016,N_19929,N_19699);
nor UO_2017 (O_2017,N_19514,N_19578);
xnor UO_2018 (O_2018,N_19854,N_19903);
nor UO_2019 (O_2019,N_19700,N_19989);
nor UO_2020 (O_2020,N_19698,N_19687);
nor UO_2021 (O_2021,N_19962,N_19972);
nor UO_2022 (O_2022,N_19602,N_19600);
nor UO_2023 (O_2023,N_19846,N_19664);
and UO_2024 (O_2024,N_19941,N_19983);
nand UO_2025 (O_2025,N_19561,N_19927);
nor UO_2026 (O_2026,N_19940,N_19864);
nand UO_2027 (O_2027,N_19656,N_19563);
nand UO_2028 (O_2028,N_19973,N_19501);
nor UO_2029 (O_2029,N_19754,N_19929);
nand UO_2030 (O_2030,N_19924,N_19622);
or UO_2031 (O_2031,N_19807,N_19834);
nor UO_2032 (O_2032,N_19864,N_19990);
nand UO_2033 (O_2033,N_19630,N_19548);
nor UO_2034 (O_2034,N_19923,N_19837);
or UO_2035 (O_2035,N_19835,N_19658);
xor UO_2036 (O_2036,N_19784,N_19607);
xor UO_2037 (O_2037,N_19890,N_19808);
and UO_2038 (O_2038,N_19967,N_19960);
nor UO_2039 (O_2039,N_19657,N_19612);
and UO_2040 (O_2040,N_19761,N_19721);
or UO_2041 (O_2041,N_19723,N_19954);
or UO_2042 (O_2042,N_19769,N_19721);
nor UO_2043 (O_2043,N_19784,N_19673);
and UO_2044 (O_2044,N_19900,N_19924);
or UO_2045 (O_2045,N_19715,N_19739);
and UO_2046 (O_2046,N_19885,N_19868);
nor UO_2047 (O_2047,N_19874,N_19536);
nor UO_2048 (O_2048,N_19863,N_19820);
and UO_2049 (O_2049,N_19733,N_19773);
nor UO_2050 (O_2050,N_19634,N_19809);
xor UO_2051 (O_2051,N_19574,N_19718);
or UO_2052 (O_2052,N_19839,N_19511);
xor UO_2053 (O_2053,N_19591,N_19787);
or UO_2054 (O_2054,N_19562,N_19815);
and UO_2055 (O_2055,N_19516,N_19742);
xnor UO_2056 (O_2056,N_19744,N_19941);
or UO_2057 (O_2057,N_19811,N_19888);
and UO_2058 (O_2058,N_19964,N_19597);
and UO_2059 (O_2059,N_19685,N_19795);
and UO_2060 (O_2060,N_19625,N_19898);
nand UO_2061 (O_2061,N_19930,N_19900);
nand UO_2062 (O_2062,N_19701,N_19753);
xor UO_2063 (O_2063,N_19919,N_19640);
xnor UO_2064 (O_2064,N_19882,N_19950);
nor UO_2065 (O_2065,N_19709,N_19541);
nand UO_2066 (O_2066,N_19816,N_19628);
and UO_2067 (O_2067,N_19698,N_19789);
and UO_2068 (O_2068,N_19947,N_19721);
or UO_2069 (O_2069,N_19840,N_19656);
and UO_2070 (O_2070,N_19998,N_19608);
nor UO_2071 (O_2071,N_19763,N_19904);
xor UO_2072 (O_2072,N_19979,N_19594);
or UO_2073 (O_2073,N_19858,N_19936);
nand UO_2074 (O_2074,N_19892,N_19671);
or UO_2075 (O_2075,N_19754,N_19987);
nand UO_2076 (O_2076,N_19519,N_19849);
nor UO_2077 (O_2077,N_19992,N_19562);
and UO_2078 (O_2078,N_19516,N_19727);
nor UO_2079 (O_2079,N_19587,N_19611);
and UO_2080 (O_2080,N_19746,N_19854);
nand UO_2081 (O_2081,N_19707,N_19834);
nand UO_2082 (O_2082,N_19773,N_19930);
xnor UO_2083 (O_2083,N_19599,N_19745);
nor UO_2084 (O_2084,N_19534,N_19979);
nand UO_2085 (O_2085,N_19607,N_19573);
nand UO_2086 (O_2086,N_19539,N_19889);
or UO_2087 (O_2087,N_19552,N_19952);
or UO_2088 (O_2088,N_19760,N_19712);
nand UO_2089 (O_2089,N_19560,N_19531);
xnor UO_2090 (O_2090,N_19710,N_19693);
nor UO_2091 (O_2091,N_19884,N_19992);
xor UO_2092 (O_2092,N_19550,N_19945);
nand UO_2093 (O_2093,N_19716,N_19895);
or UO_2094 (O_2094,N_19735,N_19930);
xor UO_2095 (O_2095,N_19831,N_19732);
xnor UO_2096 (O_2096,N_19528,N_19828);
and UO_2097 (O_2097,N_19949,N_19631);
nand UO_2098 (O_2098,N_19941,N_19680);
nand UO_2099 (O_2099,N_19864,N_19837);
and UO_2100 (O_2100,N_19545,N_19979);
and UO_2101 (O_2101,N_19679,N_19718);
xor UO_2102 (O_2102,N_19655,N_19877);
nor UO_2103 (O_2103,N_19827,N_19608);
nand UO_2104 (O_2104,N_19599,N_19803);
or UO_2105 (O_2105,N_19668,N_19693);
or UO_2106 (O_2106,N_19708,N_19603);
or UO_2107 (O_2107,N_19640,N_19941);
xnor UO_2108 (O_2108,N_19937,N_19670);
nand UO_2109 (O_2109,N_19739,N_19741);
nor UO_2110 (O_2110,N_19942,N_19844);
nand UO_2111 (O_2111,N_19653,N_19911);
nand UO_2112 (O_2112,N_19535,N_19937);
xnor UO_2113 (O_2113,N_19622,N_19850);
nor UO_2114 (O_2114,N_19615,N_19640);
nor UO_2115 (O_2115,N_19912,N_19904);
and UO_2116 (O_2116,N_19799,N_19984);
nand UO_2117 (O_2117,N_19738,N_19792);
nor UO_2118 (O_2118,N_19817,N_19918);
and UO_2119 (O_2119,N_19853,N_19695);
nand UO_2120 (O_2120,N_19892,N_19643);
nor UO_2121 (O_2121,N_19503,N_19527);
and UO_2122 (O_2122,N_19745,N_19872);
and UO_2123 (O_2123,N_19612,N_19729);
nand UO_2124 (O_2124,N_19712,N_19915);
nor UO_2125 (O_2125,N_19700,N_19879);
nand UO_2126 (O_2126,N_19589,N_19794);
and UO_2127 (O_2127,N_19922,N_19999);
nand UO_2128 (O_2128,N_19552,N_19545);
or UO_2129 (O_2129,N_19940,N_19844);
nor UO_2130 (O_2130,N_19847,N_19801);
xor UO_2131 (O_2131,N_19672,N_19814);
nand UO_2132 (O_2132,N_19654,N_19780);
nor UO_2133 (O_2133,N_19897,N_19775);
nor UO_2134 (O_2134,N_19748,N_19708);
or UO_2135 (O_2135,N_19807,N_19670);
xnor UO_2136 (O_2136,N_19626,N_19987);
xnor UO_2137 (O_2137,N_19860,N_19640);
and UO_2138 (O_2138,N_19965,N_19822);
xor UO_2139 (O_2139,N_19616,N_19841);
nand UO_2140 (O_2140,N_19824,N_19703);
or UO_2141 (O_2141,N_19983,N_19847);
nand UO_2142 (O_2142,N_19619,N_19893);
and UO_2143 (O_2143,N_19702,N_19968);
and UO_2144 (O_2144,N_19575,N_19618);
xnor UO_2145 (O_2145,N_19625,N_19721);
and UO_2146 (O_2146,N_19771,N_19834);
or UO_2147 (O_2147,N_19874,N_19769);
nor UO_2148 (O_2148,N_19603,N_19928);
and UO_2149 (O_2149,N_19694,N_19965);
or UO_2150 (O_2150,N_19601,N_19515);
xor UO_2151 (O_2151,N_19610,N_19868);
or UO_2152 (O_2152,N_19782,N_19954);
or UO_2153 (O_2153,N_19742,N_19513);
or UO_2154 (O_2154,N_19806,N_19580);
or UO_2155 (O_2155,N_19787,N_19900);
or UO_2156 (O_2156,N_19865,N_19632);
xnor UO_2157 (O_2157,N_19936,N_19982);
or UO_2158 (O_2158,N_19718,N_19889);
and UO_2159 (O_2159,N_19687,N_19809);
xor UO_2160 (O_2160,N_19885,N_19624);
nand UO_2161 (O_2161,N_19510,N_19858);
nor UO_2162 (O_2162,N_19935,N_19862);
nand UO_2163 (O_2163,N_19856,N_19645);
nand UO_2164 (O_2164,N_19778,N_19747);
or UO_2165 (O_2165,N_19742,N_19745);
xor UO_2166 (O_2166,N_19760,N_19598);
xnor UO_2167 (O_2167,N_19802,N_19601);
and UO_2168 (O_2168,N_19708,N_19755);
nand UO_2169 (O_2169,N_19691,N_19872);
or UO_2170 (O_2170,N_19528,N_19815);
nand UO_2171 (O_2171,N_19558,N_19528);
nor UO_2172 (O_2172,N_19964,N_19634);
and UO_2173 (O_2173,N_19816,N_19605);
nand UO_2174 (O_2174,N_19728,N_19892);
xnor UO_2175 (O_2175,N_19652,N_19518);
or UO_2176 (O_2176,N_19845,N_19762);
xnor UO_2177 (O_2177,N_19705,N_19612);
and UO_2178 (O_2178,N_19956,N_19526);
xnor UO_2179 (O_2179,N_19856,N_19504);
xor UO_2180 (O_2180,N_19888,N_19703);
and UO_2181 (O_2181,N_19791,N_19837);
nand UO_2182 (O_2182,N_19841,N_19633);
nor UO_2183 (O_2183,N_19969,N_19537);
xnor UO_2184 (O_2184,N_19849,N_19511);
xnor UO_2185 (O_2185,N_19513,N_19624);
nor UO_2186 (O_2186,N_19637,N_19507);
xor UO_2187 (O_2187,N_19528,N_19569);
nand UO_2188 (O_2188,N_19541,N_19644);
nor UO_2189 (O_2189,N_19735,N_19830);
or UO_2190 (O_2190,N_19912,N_19781);
or UO_2191 (O_2191,N_19565,N_19825);
and UO_2192 (O_2192,N_19981,N_19748);
nor UO_2193 (O_2193,N_19774,N_19875);
nor UO_2194 (O_2194,N_19740,N_19919);
or UO_2195 (O_2195,N_19600,N_19741);
and UO_2196 (O_2196,N_19657,N_19769);
nor UO_2197 (O_2197,N_19949,N_19648);
or UO_2198 (O_2198,N_19996,N_19551);
or UO_2199 (O_2199,N_19874,N_19732);
nor UO_2200 (O_2200,N_19758,N_19776);
nand UO_2201 (O_2201,N_19756,N_19731);
or UO_2202 (O_2202,N_19808,N_19696);
and UO_2203 (O_2203,N_19768,N_19776);
nand UO_2204 (O_2204,N_19531,N_19770);
nor UO_2205 (O_2205,N_19943,N_19733);
xor UO_2206 (O_2206,N_19807,N_19744);
nand UO_2207 (O_2207,N_19917,N_19703);
nand UO_2208 (O_2208,N_19620,N_19821);
and UO_2209 (O_2209,N_19868,N_19812);
or UO_2210 (O_2210,N_19699,N_19598);
nor UO_2211 (O_2211,N_19840,N_19775);
and UO_2212 (O_2212,N_19672,N_19917);
and UO_2213 (O_2213,N_19707,N_19870);
nand UO_2214 (O_2214,N_19816,N_19931);
nor UO_2215 (O_2215,N_19674,N_19856);
nor UO_2216 (O_2216,N_19953,N_19862);
nand UO_2217 (O_2217,N_19642,N_19614);
xnor UO_2218 (O_2218,N_19552,N_19976);
xor UO_2219 (O_2219,N_19715,N_19786);
xor UO_2220 (O_2220,N_19977,N_19721);
or UO_2221 (O_2221,N_19737,N_19525);
xnor UO_2222 (O_2222,N_19955,N_19610);
xor UO_2223 (O_2223,N_19780,N_19807);
nand UO_2224 (O_2224,N_19637,N_19524);
xor UO_2225 (O_2225,N_19798,N_19592);
or UO_2226 (O_2226,N_19868,N_19727);
nor UO_2227 (O_2227,N_19927,N_19729);
nor UO_2228 (O_2228,N_19616,N_19550);
or UO_2229 (O_2229,N_19591,N_19942);
or UO_2230 (O_2230,N_19611,N_19588);
and UO_2231 (O_2231,N_19899,N_19958);
nor UO_2232 (O_2232,N_19623,N_19667);
or UO_2233 (O_2233,N_19869,N_19721);
and UO_2234 (O_2234,N_19566,N_19846);
and UO_2235 (O_2235,N_19750,N_19563);
and UO_2236 (O_2236,N_19785,N_19558);
or UO_2237 (O_2237,N_19564,N_19514);
and UO_2238 (O_2238,N_19561,N_19938);
xnor UO_2239 (O_2239,N_19710,N_19715);
and UO_2240 (O_2240,N_19952,N_19867);
and UO_2241 (O_2241,N_19711,N_19825);
or UO_2242 (O_2242,N_19670,N_19545);
or UO_2243 (O_2243,N_19972,N_19560);
or UO_2244 (O_2244,N_19727,N_19865);
xor UO_2245 (O_2245,N_19963,N_19576);
and UO_2246 (O_2246,N_19967,N_19959);
nand UO_2247 (O_2247,N_19942,N_19842);
or UO_2248 (O_2248,N_19576,N_19588);
nor UO_2249 (O_2249,N_19677,N_19966);
nand UO_2250 (O_2250,N_19818,N_19595);
and UO_2251 (O_2251,N_19664,N_19830);
nand UO_2252 (O_2252,N_19712,N_19709);
xor UO_2253 (O_2253,N_19672,N_19896);
xor UO_2254 (O_2254,N_19621,N_19942);
nor UO_2255 (O_2255,N_19567,N_19918);
nand UO_2256 (O_2256,N_19748,N_19809);
nand UO_2257 (O_2257,N_19858,N_19721);
nor UO_2258 (O_2258,N_19858,N_19833);
or UO_2259 (O_2259,N_19838,N_19577);
and UO_2260 (O_2260,N_19957,N_19571);
or UO_2261 (O_2261,N_19649,N_19902);
nor UO_2262 (O_2262,N_19766,N_19705);
nand UO_2263 (O_2263,N_19672,N_19554);
and UO_2264 (O_2264,N_19719,N_19908);
nand UO_2265 (O_2265,N_19975,N_19607);
nand UO_2266 (O_2266,N_19918,N_19512);
xnor UO_2267 (O_2267,N_19851,N_19690);
nor UO_2268 (O_2268,N_19728,N_19652);
xnor UO_2269 (O_2269,N_19975,N_19971);
nand UO_2270 (O_2270,N_19500,N_19821);
nand UO_2271 (O_2271,N_19651,N_19508);
nor UO_2272 (O_2272,N_19992,N_19708);
xnor UO_2273 (O_2273,N_19829,N_19657);
nand UO_2274 (O_2274,N_19599,N_19652);
nor UO_2275 (O_2275,N_19756,N_19904);
nor UO_2276 (O_2276,N_19978,N_19884);
nor UO_2277 (O_2277,N_19812,N_19724);
and UO_2278 (O_2278,N_19871,N_19648);
nor UO_2279 (O_2279,N_19520,N_19913);
xnor UO_2280 (O_2280,N_19893,N_19526);
nor UO_2281 (O_2281,N_19890,N_19882);
nand UO_2282 (O_2282,N_19977,N_19947);
nor UO_2283 (O_2283,N_19593,N_19523);
xor UO_2284 (O_2284,N_19591,N_19553);
xnor UO_2285 (O_2285,N_19940,N_19588);
and UO_2286 (O_2286,N_19590,N_19555);
nor UO_2287 (O_2287,N_19852,N_19690);
nor UO_2288 (O_2288,N_19945,N_19801);
nand UO_2289 (O_2289,N_19960,N_19848);
nor UO_2290 (O_2290,N_19551,N_19636);
or UO_2291 (O_2291,N_19824,N_19544);
nand UO_2292 (O_2292,N_19738,N_19554);
nand UO_2293 (O_2293,N_19788,N_19883);
or UO_2294 (O_2294,N_19784,N_19611);
and UO_2295 (O_2295,N_19528,N_19618);
or UO_2296 (O_2296,N_19720,N_19562);
nor UO_2297 (O_2297,N_19566,N_19642);
nand UO_2298 (O_2298,N_19630,N_19709);
or UO_2299 (O_2299,N_19938,N_19545);
nand UO_2300 (O_2300,N_19603,N_19684);
nor UO_2301 (O_2301,N_19662,N_19704);
and UO_2302 (O_2302,N_19816,N_19855);
nand UO_2303 (O_2303,N_19784,N_19600);
xnor UO_2304 (O_2304,N_19678,N_19736);
nor UO_2305 (O_2305,N_19675,N_19770);
nor UO_2306 (O_2306,N_19888,N_19772);
nor UO_2307 (O_2307,N_19911,N_19567);
xnor UO_2308 (O_2308,N_19888,N_19825);
and UO_2309 (O_2309,N_19687,N_19718);
nand UO_2310 (O_2310,N_19848,N_19905);
nand UO_2311 (O_2311,N_19769,N_19640);
nor UO_2312 (O_2312,N_19685,N_19919);
or UO_2313 (O_2313,N_19525,N_19554);
and UO_2314 (O_2314,N_19983,N_19665);
or UO_2315 (O_2315,N_19954,N_19575);
xor UO_2316 (O_2316,N_19744,N_19972);
xnor UO_2317 (O_2317,N_19883,N_19865);
and UO_2318 (O_2318,N_19816,N_19632);
xnor UO_2319 (O_2319,N_19764,N_19650);
nand UO_2320 (O_2320,N_19561,N_19593);
nand UO_2321 (O_2321,N_19878,N_19975);
and UO_2322 (O_2322,N_19910,N_19926);
nand UO_2323 (O_2323,N_19871,N_19773);
or UO_2324 (O_2324,N_19779,N_19559);
or UO_2325 (O_2325,N_19782,N_19690);
nand UO_2326 (O_2326,N_19552,N_19914);
and UO_2327 (O_2327,N_19620,N_19893);
nor UO_2328 (O_2328,N_19695,N_19630);
nand UO_2329 (O_2329,N_19824,N_19557);
or UO_2330 (O_2330,N_19973,N_19792);
or UO_2331 (O_2331,N_19502,N_19670);
and UO_2332 (O_2332,N_19947,N_19643);
and UO_2333 (O_2333,N_19520,N_19583);
xnor UO_2334 (O_2334,N_19992,N_19901);
or UO_2335 (O_2335,N_19858,N_19546);
nand UO_2336 (O_2336,N_19798,N_19996);
nor UO_2337 (O_2337,N_19678,N_19900);
or UO_2338 (O_2338,N_19691,N_19711);
and UO_2339 (O_2339,N_19666,N_19659);
nand UO_2340 (O_2340,N_19994,N_19868);
nand UO_2341 (O_2341,N_19911,N_19954);
nor UO_2342 (O_2342,N_19524,N_19508);
nor UO_2343 (O_2343,N_19776,N_19646);
nand UO_2344 (O_2344,N_19635,N_19951);
or UO_2345 (O_2345,N_19614,N_19689);
xnor UO_2346 (O_2346,N_19746,N_19819);
nor UO_2347 (O_2347,N_19622,N_19989);
nor UO_2348 (O_2348,N_19670,N_19789);
xor UO_2349 (O_2349,N_19843,N_19987);
nor UO_2350 (O_2350,N_19730,N_19532);
or UO_2351 (O_2351,N_19910,N_19701);
xor UO_2352 (O_2352,N_19742,N_19656);
or UO_2353 (O_2353,N_19637,N_19960);
nand UO_2354 (O_2354,N_19610,N_19947);
xnor UO_2355 (O_2355,N_19586,N_19689);
nor UO_2356 (O_2356,N_19646,N_19847);
xnor UO_2357 (O_2357,N_19710,N_19583);
or UO_2358 (O_2358,N_19863,N_19577);
and UO_2359 (O_2359,N_19636,N_19881);
and UO_2360 (O_2360,N_19854,N_19828);
or UO_2361 (O_2361,N_19803,N_19578);
and UO_2362 (O_2362,N_19940,N_19526);
and UO_2363 (O_2363,N_19836,N_19556);
xor UO_2364 (O_2364,N_19753,N_19958);
nand UO_2365 (O_2365,N_19718,N_19642);
nor UO_2366 (O_2366,N_19642,N_19551);
xnor UO_2367 (O_2367,N_19840,N_19990);
or UO_2368 (O_2368,N_19572,N_19871);
or UO_2369 (O_2369,N_19598,N_19755);
xor UO_2370 (O_2370,N_19584,N_19694);
nand UO_2371 (O_2371,N_19805,N_19898);
nor UO_2372 (O_2372,N_19998,N_19720);
nand UO_2373 (O_2373,N_19856,N_19736);
and UO_2374 (O_2374,N_19866,N_19907);
and UO_2375 (O_2375,N_19672,N_19918);
nor UO_2376 (O_2376,N_19844,N_19508);
nand UO_2377 (O_2377,N_19791,N_19961);
or UO_2378 (O_2378,N_19573,N_19750);
nor UO_2379 (O_2379,N_19588,N_19624);
xor UO_2380 (O_2380,N_19595,N_19729);
and UO_2381 (O_2381,N_19918,N_19880);
xor UO_2382 (O_2382,N_19981,N_19817);
nor UO_2383 (O_2383,N_19934,N_19795);
and UO_2384 (O_2384,N_19613,N_19776);
or UO_2385 (O_2385,N_19994,N_19619);
xor UO_2386 (O_2386,N_19584,N_19636);
nand UO_2387 (O_2387,N_19783,N_19566);
nand UO_2388 (O_2388,N_19769,N_19905);
xnor UO_2389 (O_2389,N_19697,N_19592);
xnor UO_2390 (O_2390,N_19937,N_19847);
or UO_2391 (O_2391,N_19676,N_19898);
nor UO_2392 (O_2392,N_19505,N_19541);
and UO_2393 (O_2393,N_19511,N_19663);
and UO_2394 (O_2394,N_19700,N_19734);
xnor UO_2395 (O_2395,N_19920,N_19907);
nand UO_2396 (O_2396,N_19618,N_19723);
nand UO_2397 (O_2397,N_19770,N_19650);
xnor UO_2398 (O_2398,N_19899,N_19755);
or UO_2399 (O_2399,N_19737,N_19704);
nand UO_2400 (O_2400,N_19531,N_19875);
nand UO_2401 (O_2401,N_19830,N_19621);
nand UO_2402 (O_2402,N_19653,N_19646);
nor UO_2403 (O_2403,N_19923,N_19534);
nor UO_2404 (O_2404,N_19915,N_19506);
nand UO_2405 (O_2405,N_19627,N_19899);
nor UO_2406 (O_2406,N_19727,N_19724);
nand UO_2407 (O_2407,N_19614,N_19613);
xor UO_2408 (O_2408,N_19994,N_19634);
and UO_2409 (O_2409,N_19859,N_19854);
and UO_2410 (O_2410,N_19784,N_19634);
xor UO_2411 (O_2411,N_19517,N_19985);
or UO_2412 (O_2412,N_19720,N_19634);
or UO_2413 (O_2413,N_19882,N_19900);
nand UO_2414 (O_2414,N_19634,N_19956);
xnor UO_2415 (O_2415,N_19694,N_19800);
nand UO_2416 (O_2416,N_19546,N_19594);
xor UO_2417 (O_2417,N_19914,N_19855);
nor UO_2418 (O_2418,N_19747,N_19933);
xor UO_2419 (O_2419,N_19555,N_19589);
xnor UO_2420 (O_2420,N_19838,N_19954);
nand UO_2421 (O_2421,N_19911,N_19645);
nor UO_2422 (O_2422,N_19636,N_19509);
xor UO_2423 (O_2423,N_19735,N_19941);
xnor UO_2424 (O_2424,N_19637,N_19723);
or UO_2425 (O_2425,N_19646,N_19991);
nor UO_2426 (O_2426,N_19672,N_19534);
xor UO_2427 (O_2427,N_19809,N_19820);
nand UO_2428 (O_2428,N_19973,N_19508);
xnor UO_2429 (O_2429,N_19928,N_19760);
nor UO_2430 (O_2430,N_19767,N_19743);
nor UO_2431 (O_2431,N_19761,N_19672);
and UO_2432 (O_2432,N_19779,N_19785);
nand UO_2433 (O_2433,N_19510,N_19652);
nand UO_2434 (O_2434,N_19833,N_19549);
nor UO_2435 (O_2435,N_19542,N_19734);
nor UO_2436 (O_2436,N_19749,N_19701);
nor UO_2437 (O_2437,N_19929,N_19737);
xnor UO_2438 (O_2438,N_19805,N_19615);
nor UO_2439 (O_2439,N_19713,N_19671);
nor UO_2440 (O_2440,N_19837,N_19852);
or UO_2441 (O_2441,N_19632,N_19780);
and UO_2442 (O_2442,N_19666,N_19865);
nand UO_2443 (O_2443,N_19727,N_19726);
or UO_2444 (O_2444,N_19842,N_19655);
nor UO_2445 (O_2445,N_19887,N_19852);
and UO_2446 (O_2446,N_19681,N_19985);
nor UO_2447 (O_2447,N_19945,N_19881);
or UO_2448 (O_2448,N_19561,N_19900);
and UO_2449 (O_2449,N_19710,N_19971);
or UO_2450 (O_2450,N_19918,N_19971);
and UO_2451 (O_2451,N_19675,N_19506);
nor UO_2452 (O_2452,N_19579,N_19689);
xor UO_2453 (O_2453,N_19530,N_19758);
xor UO_2454 (O_2454,N_19571,N_19854);
and UO_2455 (O_2455,N_19749,N_19772);
nor UO_2456 (O_2456,N_19910,N_19523);
xor UO_2457 (O_2457,N_19607,N_19894);
nor UO_2458 (O_2458,N_19945,N_19974);
nand UO_2459 (O_2459,N_19554,N_19888);
or UO_2460 (O_2460,N_19572,N_19580);
xnor UO_2461 (O_2461,N_19800,N_19999);
or UO_2462 (O_2462,N_19559,N_19804);
and UO_2463 (O_2463,N_19878,N_19993);
or UO_2464 (O_2464,N_19649,N_19559);
and UO_2465 (O_2465,N_19719,N_19870);
nand UO_2466 (O_2466,N_19556,N_19779);
and UO_2467 (O_2467,N_19678,N_19868);
nor UO_2468 (O_2468,N_19572,N_19695);
nand UO_2469 (O_2469,N_19823,N_19932);
nor UO_2470 (O_2470,N_19698,N_19603);
nor UO_2471 (O_2471,N_19706,N_19850);
and UO_2472 (O_2472,N_19593,N_19668);
or UO_2473 (O_2473,N_19568,N_19986);
and UO_2474 (O_2474,N_19805,N_19573);
and UO_2475 (O_2475,N_19734,N_19761);
and UO_2476 (O_2476,N_19668,N_19833);
or UO_2477 (O_2477,N_19538,N_19624);
or UO_2478 (O_2478,N_19852,N_19627);
nor UO_2479 (O_2479,N_19617,N_19789);
nand UO_2480 (O_2480,N_19952,N_19904);
or UO_2481 (O_2481,N_19620,N_19699);
nor UO_2482 (O_2482,N_19740,N_19547);
and UO_2483 (O_2483,N_19520,N_19672);
and UO_2484 (O_2484,N_19553,N_19959);
nor UO_2485 (O_2485,N_19730,N_19823);
or UO_2486 (O_2486,N_19940,N_19746);
and UO_2487 (O_2487,N_19658,N_19679);
or UO_2488 (O_2488,N_19797,N_19579);
or UO_2489 (O_2489,N_19947,N_19884);
and UO_2490 (O_2490,N_19719,N_19566);
xnor UO_2491 (O_2491,N_19909,N_19634);
nor UO_2492 (O_2492,N_19612,N_19777);
nand UO_2493 (O_2493,N_19563,N_19517);
and UO_2494 (O_2494,N_19999,N_19541);
nor UO_2495 (O_2495,N_19766,N_19796);
or UO_2496 (O_2496,N_19997,N_19537);
nand UO_2497 (O_2497,N_19711,N_19953);
xor UO_2498 (O_2498,N_19869,N_19518);
nand UO_2499 (O_2499,N_19775,N_19864);
endmodule