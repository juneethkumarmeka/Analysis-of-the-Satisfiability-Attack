module basic_2000_20000_2500_4_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
xor U0 (N_0,In_1508,In_1962);
and U1 (N_1,In_71,In_1580);
nand U2 (N_2,In_676,In_1897);
nand U3 (N_3,In_1726,In_487);
nor U4 (N_4,In_1949,In_1947);
nor U5 (N_5,In_640,In_1226);
nand U6 (N_6,In_45,In_357);
and U7 (N_7,In_1078,In_792);
nand U8 (N_8,In_1910,In_617);
and U9 (N_9,In_540,In_97);
or U10 (N_10,In_1400,In_1921);
and U11 (N_11,In_1925,In_393);
nand U12 (N_12,In_1570,In_212);
xnor U13 (N_13,In_1835,In_1082);
and U14 (N_14,In_1868,In_508);
nand U15 (N_15,In_1061,In_529);
nor U16 (N_16,In_951,In_671);
nor U17 (N_17,In_1653,In_448);
nand U18 (N_18,In_1292,In_1877);
nor U19 (N_19,In_1687,In_1118);
nor U20 (N_20,In_1094,In_1373);
nand U21 (N_21,In_1225,In_124);
nand U22 (N_22,In_1756,In_477);
or U23 (N_23,In_1267,In_492);
and U24 (N_24,In_713,In_26);
nand U25 (N_25,In_457,In_317);
nand U26 (N_26,In_145,In_956);
or U27 (N_27,In_1655,In_256);
or U28 (N_28,In_615,In_1755);
and U29 (N_29,In_331,In_1814);
and U30 (N_30,In_670,In_1338);
xor U31 (N_31,In_63,In_1608);
or U32 (N_32,In_942,In_922);
nand U33 (N_33,In_1629,In_368);
nand U34 (N_34,In_948,In_316);
or U35 (N_35,In_1932,In_1989);
nor U36 (N_36,In_680,In_734);
or U37 (N_37,In_963,In_702);
and U38 (N_38,In_1283,In_335);
or U39 (N_39,In_1873,In_1818);
nor U40 (N_40,In_892,In_1144);
or U41 (N_41,In_631,In_1208);
nand U42 (N_42,In_1209,In_1642);
and U43 (N_43,In_285,In_1434);
nor U44 (N_44,In_218,In_698);
xnor U45 (N_45,In_36,In_1132);
nor U46 (N_46,In_49,In_1811);
and U47 (N_47,In_1996,In_496);
or U48 (N_48,In_1831,In_310);
nor U49 (N_49,In_428,In_1048);
or U50 (N_50,In_987,In_1488);
nand U51 (N_51,In_1360,In_226);
nand U52 (N_52,In_1673,In_297);
xnor U53 (N_53,In_1821,In_501);
nor U54 (N_54,In_195,In_1843);
and U55 (N_55,In_1768,In_1201);
nand U56 (N_56,In_154,In_585);
nor U57 (N_57,In_1593,In_1858);
or U58 (N_58,In_211,In_382);
or U59 (N_59,In_1364,In_243);
and U60 (N_60,In_486,In_1515);
nor U61 (N_61,In_967,In_1969);
nor U62 (N_62,In_1241,In_128);
nor U63 (N_63,In_1119,In_1869);
nand U64 (N_64,In_1248,In_525);
xor U65 (N_65,In_887,In_1540);
and U66 (N_66,In_665,In_1047);
nand U67 (N_67,In_1813,In_715);
nor U68 (N_68,In_449,In_1046);
nor U69 (N_69,In_1020,In_338);
or U70 (N_70,In_1345,In_1291);
nand U71 (N_71,In_1310,In_445);
nor U72 (N_72,In_1139,In_242);
nand U73 (N_73,In_111,In_1923);
nand U74 (N_74,In_1466,In_855);
and U75 (N_75,In_1342,In_1546);
nand U76 (N_76,In_1734,In_365);
nor U77 (N_77,In_58,In_1514);
or U78 (N_78,In_882,In_1142);
and U79 (N_79,In_977,In_608);
and U80 (N_80,In_1716,In_1494);
or U81 (N_81,In_348,In_541);
or U82 (N_82,In_270,In_153);
xnor U83 (N_83,In_1808,In_1203);
nor U84 (N_84,In_1958,In_371);
nor U85 (N_85,In_1304,In_1387);
nor U86 (N_86,In_591,In_839);
nor U87 (N_87,In_1924,In_996);
and U88 (N_88,In_325,In_1929);
nor U89 (N_89,In_1912,In_1100);
nand U90 (N_90,In_1557,In_1052);
and U91 (N_91,In_1883,In_1442);
or U92 (N_92,In_602,In_1529);
nor U93 (N_93,In_1715,In_244);
or U94 (N_94,In_1143,In_1101);
xnor U95 (N_95,In_1424,In_1522);
and U96 (N_96,In_328,In_345);
and U97 (N_97,In_1952,In_1177);
nor U98 (N_98,In_970,In_51);
or U99 (N_99,In_912,In_572);
and U100 (N_100,In_1109,In_272);
and U101 (N_101,In_902,In_353);
nor U102 (N_102,In_140,In_616);
nand U103 (N_103,In_1102,In_532);
or U104 (N_104,In_710,In_421);
or U105 (N_105,In_198,In_1192);
nor U106 (N_106,In_1141,In_1327);
and U107 (N_107,In_1121,In_693);
nand U108 (N_108,In_1464,In_1917);
nor U109 (N_109,In_1946,In_1002);
and U110 (N_110,In_1484,In_1988);
and U111 (N_111,In_598,In_1185);
xor U112 (N_112,In_1658,In_1718);
and U113 (N_113,In_1809,In_994);
nor U114 (N_114,In_1797,In_594);
and U115 (N_115,In_663,In_980);
nor U116 (N_116,In_835,In_966);
xor U117 (N_117,In_1122,In_629);
or U118 (N_118,In_1487,In_379);
nor U119 (N_119,In_387,In_1272);
or U120 (N_120,In_104,In_318);
nor U121 (N_121,In_1049,In_1152);
or U122 (N_122,In_928,In_610);
xor U123 (N_123,In_1156,In_696);
nor U124 (N_124,In_68,In_664);
xor U125 (N_125,In_386,In_740);
and U126 (N_126,In_1781,In_189);
or U127 (N_127,In_1258,In_162);
or U128 (N_128,In_1224,In_1375);
xnor U129 (N_129,In_1426,In_1728);
nor U130 (N_130,In_1125,In_511);
and U131 (N_131,In_1008,In_814);
nor U132 (N_132,In_899,In_202);
nand U133 (N_133,In_1855,In_419);
and U134 (N_134,In_397,In_406);
nand U135 (N_135,In_19,In_785);
nand U136 (N_136,In_109,In_389);
xor U137 (N_137,In_1159,In_815);
nor U138 (N_138,In_1182,In_1903);
nor U139 (N_139,In_1787,In_76);
or U140 (N_140,In_60,In_574);
nor U141 (N_141,In_1034,In_582);
and U142 (N_142,In_1675,In_1535);
nor U143 (N_143,In_1922,In_846);
nor U144 (N_144,In_1127,In_105);
nand U145 (N_145,In_1348,In_116);
nor U146 (N_146,In_1908,In_777);
nand U147 (N_147,In_1422,In_1184);
xnor U148 (N_148,In_1276,In_1454);
nand U149 (N_149,In_1550,In_168);
xnor U150 (N_150,In_377,In_1215);
nor U151 (N_151,In_1363,In_3);
xor U152 (N_152,In_979,In_1386);
or U153 (N_153,In_993,In_1758);
or U154 (N_154,In_422,In_1321);
or U155 (N_155,In_1945,In_1703);
nand U156 (N_156,In_903,In_954);
nand U157 (N_157,In_1914,In_1277);
or U158 (N_158,In_1108,In_866);
and U159 (N_159,In_697,In_199);
xnor U160 (N_160,In_56,In_200);
nand U161 (N_161,In_20,In_1245);
and U162 (N_162,In_1445,In_1104);
and U163 (N_163,In_1096,In_1071);
xnor U164 (N_164,In_834,In_1722);
nor U165 (N_165,In_427,In_571);
nor U166 (N_166,In_1263,In_1157);
or U167 (N_167,In_864,In_874);
and U168 (N_168,In_867,In_502);
nand U169 (N_169,In_166,In_364);
nand U170 (N_170,In_1898,In_305);
or U171 (N_171,In_1776,In_1577);
or U172 (N_172,In_132,In_978);
nand U173 (N_173,In_1618,In_1833);
nor U174 (N_174,In_1039,In_726);
nand U175 (N_175,In_66,In_648);
xor U176 (N_176,In_612,In_471);
nor U177 (N_177,In_915,In_296);
nor U178 (N_178,In_1767,In_1693);
and U179 (N_179,In_1980,In_797);
or U180 (N_180,In_1895,In_192);
xor U181 (N_181,In_1714,In_120);
nand U182 (N_182,In_373,In_398);
nor U183 (N_183,In_1872,In_39);
nand U184 (N_184,In_183,In_1406);
or U185 (N_185,In_286,In_760);
and U186 (N_186,In_235,In_580);
or U187 (N_187,In_96,In_1347);
or U188 (N_188,In_1700,In_22);
nor U189 (N_189,In_1396,In_868);
nor U190 (N_190,In_588,In_1053);
and U191 (N_191,In_558,In_1165);
nand U192 (N_192,In_1469,In_1777);
or U193 (N_193,In_330,In_1836);
nand U194 (N_194,In_1556,In_1978);
nand U195 (N_195,In_1323,In_210);
nor U196 (N_196,In_281,In_841);
nand U197 (N_197,In_1240,In_441);
and U198 (N_198,In_454,In_1727);
nor U199 (N_199,In_1024,In_493);
and U200 (N_200,In_1249,In_374);
or U201 (N_201,In_826,In_1555);
and U202 (N_202,In_765,In_1187);
or U203 (N_203,In_55,In_40);
or U204 (N_204,In_504,In_1006);
nor U205 (N_205,In_118,In_1664);
or U206 (N_206,In_9,In_99);
and U207 (N_207,In_274,In_1234);
and U208 (N_208,In_711,In_1784);
or U209 (N_209,In_636,In_692);
nor U210 (N_210,In_384,In_681);
or U211 (N_211,In_947,In_847);
nand U212 (N_212,In_1497,In_1227);
or U213 (N_213,In_1317,In_910);
nand U214 (N_214,In_264,In_528);
or U215 (N_215,In_350,In_849);
and U216 (N_216,In_1750,In_340);
nor U217 (N_217,In_1232,In_1896);
nand U218 (N_218,In_137,In_907);
or U219 (N_219,In_1243,In_1260);
or U220 (N_220,In_921,In_1072);
or U221 (N_221,In_1188,In_1564);
or U222 (N_222,In_1154,In_1198);
or U223 (N_223,In_1155,In_415);
nand U224 (N_224,In_1711,In_682);
or U225 (N_225,In_1218,In_1805);
xnor U226 (N_226,In_47,In_906);
and U227 (N_227,In_1647,In_1000);
and U228 (N_228,In_1899,In_997);
nand U229 (N_229,In_1889,In_613);
nor U230 (N_230,In_819,In_1220);
and U231 (N_231,In_871,In_1967);
nand U232 (N_232,In_568,In_781);
or U233 (N_233,In_1247,In_1230);
nor U234 (N_234,In_1014,In_1650);
or U235 (N_235,In_779,In_1374);
xnor U236 (N_236,In_1992,In_1754);
nand U237 (N_237,In_577,In_1438);
nand U238 (N_238,In_1600,In_919);
or U239 (N_239,In_1649,In_207);
xnor U240 (N_240,In_753,In_57);
nand U241 (N_241,In_821,In_1679);
nor U242 (N_242,In_412,In_731);
nand U243 (N_243,In_1786,In_1850);
nand U244 (N_244,In_684,In_1130);
nor U245 (N_245,In_115,In_78);
nand U246 (N_246,In_181,In_1738);
nand U247 (N_247,In_1448,In_1874);
xnor U248 (N_248,In_70,In_1940);
or U249 (N_249,In_1181,In_565);
nor U250 (N_250,In_534,In_190);
and U251 (N_251,In_112,In_1775);
or U252 (N_252,In_1035,In_667);
and U253 (N_253,In_800,In_845);
nor U254 (N_254,In_859,In_1991);
or U255 (N_255,In_1079,In_1830);
xor U256 (N_256,In_273,In_1571);
nor U257 (N_257,In_512,In_893);
nor U258 (N_258,In_157,In_336);
nor U259 (N_259,In_1765,In_435);
and U260 (N_260,In_806,In_1512);
nand U261 (N_261,In_231,In_15);
or U262 (N_262,In_929,In_769);
nand U263 (N_263,In_911,In_802);
or U264 (N_264,In_1216,In_1431);
nor U265 (N_265,In_790,In_436);
and U266 (N_266,In_254,In_156);
nand U267 (N_267,In_596,In_1605);
and U268 (N_268,In_288,In_1876);
nand U269 (N_269,In_958,In_1068);
xor U270 (N_270,In_444,In_1541);
or U271 (N_271,In_556,In_625);
and U272 (N_272,In_925,In_1340);
nand U273 (N_273,In_1799,In_635);
or U274 (N_274,In_1030,In_1166);
and U275 (N_275,In_1628,In_1525);
nor U276 (N_276,In_619,In_110);
and U277 (N_277,In_633,In_1657);
and U278 (N_278,In_879,In_1388);
and U279 (N_279,In_1968,In_4);
nor U280 (N_280,In_1288,In_136);
nor U281 (N_281,In_1579,In_1942);
and U282 (N_282,In_601,In_595);
or U283 (N_283,In_934,In_361);
nor U284 (N_284,In_688,In_1252);
or U285 (N_285,In_1357,In_1519);
or U286 (N_286,In_1662,In_312);
nand U287 (N_287,In_1999,In_1973);
and U288 (N_288,In_941,In_1379);
and U289 (N_289,In_1837,In_1468);
xor U290 (N_290,In_1278,In_1933);
nand U291 (N_291,In_1759,In_704);
nor U292 (N_292,In_299,In_1113);
nor U293 (N_293,In_1528,In_1206);
or U294 (N_294,In_117,In_733);
xor U295 (N_295,In_359,In_1018);
nor U296 (N_296,In_1670,In_1381);
or U297 (N_297,In_1097,In_1861);
nand U298 (N_298,In_59,In_1599);
nand U299 (N_299,In_1548,In_727);
and U300 (N_300,In_1796,In_342);
nor U301 (N_301,In_1058,In_407);
and U302 (N_302,In_423,In_257);
nor U303 (N_303,In_164,In_644);
xor U304 (N_304,In_762,In_1212);
nor U305 (N_305,In_1133,In_858);
xor U306 (N_306,In_319,In_1280);
nor U307 (N_307,In_531,In_623);
or U308 (N_308,In_133,In_1871);
nand U309 (N_309,In_13,In_1164);
nor U310 (N_310,In_1696,In_1839);
or U311 (N_311,In_1418,In_1884);
or U312 (N_312,In_1394,In_940);
nand U313 (N_313,In_440,In_643);
or U314 (N_314,In_1421,In_510);
nand U315 (N_315,In_1708,In_1346);
nor U316 (N_316,In_1669,In_624);
nor U317 (N_317,In_1539,In_1054);
nor U318 (N_318,In_1630,In_403);
xnor U319 (N_319,In_971,In_721);
or U320 (N_320,In_380,In_981);
nand U321 (N_321,In_1335,In_587);
or U322 (N_322,In_1651,In_1480);
nand U323 (N_323,In_1812,In_527);
xor U324 (N_324,In_772,In_1848);
nand U325 (N_325,In_1825,In_466);
nand U326 (N_326,In_282,In_37);
nand U327 (N_327,In_570,In_84);
and U328 (N_328,In_1233,In_805);
or U329 (N_329,In_1376,In_1120);
or U330 (N_330,In_1724,In_1641);
nor U331 (N_331,In_327,In_1025);
nor U332 (N_332,In_33,In_34);
nand U333 (N_333,In_1455,In_102);
or U334 (N_334,In_969,In_1692);
or U335 (N_335,In_182,In_536);
nand U336 (N_336,In_322,In_1881);
and U337 (N_337,In_1916,In_355);
xnor U338 (N_338,In_283,In_952);
nand U339 (N_339,In_1616,In_1560);
and U340 (N_340,In_523,In_652);
nor U341 (N_341,In_545,In_31);
nand U342 (N_342,In_10,In_1299);
and U343 (N_343,In_62,In_234);
or U344 (N_344,In_1211,In_1023);
and U345 (N_345,In_1472,In_103);
or U346 (N_346,In_1126,In_1251);
and U347 (N_347,In_468,In_1372);
nand U348 (N_348,In_551,In_366);
xor U349 (N_349,In_72,In_1547);
and U350 (N_350,In_1524,In_0);
or U351 (N_351,In_784,In_1719);
nand U352 (N_352,In_1084,In_553);
nor U353 (N_353,In_179,In_1959);
or U354 (N_354,In_144,In_352);
and U355 (N_355,In_773,In_854);
nor U356 (N_356,In_1510,In_1928);
xnor U357 (N_357,In_1576,In_1773);
and U358 (N_358,In_1285,In_524);
nor U359 (N_359,In_1385,In_370);
or U360 (N_360,In_152,In_505);
nand U361 (N_361,In_1341,In_808);
and U362 (N_362,In_1984,In_134);
and U363 (N_363,In_1197,In_1764);
or U364 (N_364,In_1467,In_32);
xor U365 (N_365,In_844,In_1795);
nor U366 (N_366,In_1516,In_1195);
or U367 (N_367,In_1935,In_432);
and U368 (N_368,In_453,In_509);
and U369 (N_369,In_95,In_1931);
or U370 (N_370,In_1575,In_1383);
or U371 (N_371,In_1485,In_1066);
xor U372 (N_372,In_810,In_961);
nand U373 (N_373,In_775,In_869);
nor U374 (N_374,In_425,In_1834);
and U375 (N_375,In_798,In_1013);
nor U376 (N_376,In_1532,In_1789);
and U377 (N_377,In_131,In_1584);
and U378 (N_378,In_1880,In_1213);
or U379 (N_379,In_1117,In_1879);
and U380 (N_380,In_1410,In_573);
or U381 (N_381,In_1167,In_443);
and U382 (N_382,In_817,In_1029);
nand U383 (N_383,In_430,In_660);
nand U384 (N_384,In_1915,In_1875);
nand U385 (N_385,In_402,In_439);
nor U386 (N_386,In_271,In_1934);
nand U387 (N_387,In_1436,In_668);
or U388 (N_388,In_1685,In_888);
xnor U389 (N_389,In_935,In_1255);
nor U390 (N_390,In_861,In_985);
or U391 (N_391,In_840,In_1287);
xnor U392 (N_392,In_1302,In_146);
nand U393 (N_393,In_173,In_1806);
nor U394 (N_394,In_1736,In_1087);
nor U395 (N_395,In_860,In_1561);
nand U396 (N_396,In_246,In_1003);
and U397 (N_397,In_404,In_1511);
and U398 (N_398,In_475,In_227);
nor U399 (N_399,In_1802,In_1456);
nand U400 (N_400,In_507,In_1533);
nand U401 (N_401,In_576,In_1778);
xnor U402 (N_402,In_836,In_1085);
or U403 (N_403,In_1960,In_148);
or U404 (N_404,In_184,In_1526);
and U405 (N_405,In_1744,In_1256);
nand U406 (N_406,In_219,In_1452);
and U407 (N_407,In_1965,In_724);
nor U408 (N_408,In_1862,In_339);
xnor U409 (N_409,In_160,In_1955);
nor U410 (N_410,In_1891,In_91);
and U411 (N_411,In_1706,In_630);
nor U412 (N_412,In_991,In_75);
xnor U413 (N_413,In_1970,In_1572);
nand U414 (N_414,In_627,In_142);
nor U415 (N_415,In_490,In_424);
nor U416 (N_416,In_44,In_1659);
nor U417 (N_417,In_522,In_794);
and U418 (N_418,In_1042,In_266);
or U419 (N_419,In_1076,In_369);
and U420 (N_420,In_1289,In_1595);
nand U421 (N_421,In_1851,In_544);
nand U422 (N_422,In_1660,In_1766);
nand U423 (N_423,In_1366,In_637);
and U424 (N_424,In_685,In_1179);
nor U425 (N_425,In_1151,In_125);
and U426 (N_426,In_16,In_161);
and U427 (N_427,In_677,In_1950);
or U428 (N_428,In_807,In_459);
nor U429 (N_429,In_1749,In_1325);
nor U430 (N_430,In_926,In_1471);
xnor U431 (N_431,In_1146,In_1017);
nor U432 (N_432,In_138,In_1483);
nand U433 (N_433,In_18,In_1699);
and U434 (N_434,In_88,In_1390);
and U435 (N_435,In_1619,In_795);
and U436 (N_436,In_298,In_1476);
nor U437 (N_437,In_1936,In_1045);
nor U438 (N_438,In_1663,In_1189);
or U439 (N_439,In_1404,In_774);
and U440 (N_440,In_1238,In_691);
xor U441 (N_441,In_1769,In_825);
nor U442 (N_442,In_965,In_533);
xor U443 (N_443,In_1845,In_1490);
or U444 (N_444,In_962,In_885);
nor U445 (N_445,In_896,In_65);
nand U446 (N_446,In_1731,In_1183);
nand U447 (N_447,In_1905,In_188);
nand U448 (N_448,In_277,In_889);
and U449 (N_449,In_354,In_1073);
nor U450 (N_450,In_1543,In_294);
xor U451 (N_451,In_1757,In_1505);
and U452 (N_452,In_535,In_1517);
xnor U453 (N_453,In_141,In_346);
and U454 (N_454,In_1038,In_1681);
nand U455 (N_455,In_707,In_1328);
nand U456 (N_456,In_1717,In_221);
or U457 (N_457,In_1083,In_669);
or U458 (N_458,In_1611,In_728);
nor U459 (N_459,In_260,In_1506);
and U460 (N_460,In_933,In_518);
or U461 (N_461,In_597,In_708);
xor U462 (N_462,In_1606,In_1175);
xnor U463 (N_463,In_549,In_1173);
xnor U464 (N_464,In_267,In_1665);
or U465 (N_465,In_1723,In_1844);
or U466 (N_466,In_1244,In_1041);
or U467 (N_467,In_870,In_291);
nand U468 (N_468,In_1334,In_1919);
nand U469 (N_469,In_848,In_600);
and U470 (N_470,In_1191,In_590);
xor U471 (N_471,In_1378,In_1680);
nand U472 (N_472,In_12,In_1743);
or U473 (N_473,In_1282,In_695);
nand U474 (N_474,In_1171,In_519);
and U475 (N_475,In_1405,In_583);
nand U476 (N_476,In_1637,In_1852);
xnor U477 (N_477,In_832,In_1523);
nand U478 (N_478,In_1951,In_537);
nor U479 (N_479,In_1210,In_209);
and U480 (N_480,In_1586,In_530);
nor U481 (N_481,In_1826,In_1823);
nor U482 (N_482,In_675,In_898);
and U483 (N_483,In_42,In_1648);
or U484 (N_484,In_1051,In_1086);
and U485 (N_485,In_1237,In_1242);
nand U486 (N_486,In_1856,In_811);
nor U487 (N_487,In_1816,In_1358);
nor U488 (N_488,In_1943,In_1273);
or U489 (N_489,In_706,In_838);
or U490 (N_490,In_959,In_569);
or U491 (N_491,In_483,In_1269);
nor U492 (N_492,In_526,In_240);
and U493 (N_493,In_478,In_1791);
and U494 (N_494,In_1704,In_313);
and U495 (N_495,In_1666,In_1573);
xor U496 (N_496,In_479,In_1033);
nand U497 (N_497,In_986,In_932);
nand U498 (N_498,In_1080,In_147);
xnor U499 (N_499,In_1676,In_1332);
nor U500 (N_500,In_1939,In_383);
nand U501 (N_501,In_546,In_334);
nor U502 (N_502,In_1067,In_349);
and U503 (N_503,In_484,In_1309);
and U504 (N_504,In_662,In_873);
nor U505 (N_505,In_1646,In_201);
nor U506 (N_506,In_1721,In_333);
or U507 (N_507,In_94,In_1205);
or U508 (N_508,In_614,In_564);
nand U509 (N_509,In_749,In_372);
nor U510 (N_510,In_801,In_1592);
nand U511 (N_511,In_1057,In_1239);
xnor U512 (N_512,In_1730,In_381);
xor U513 (N_513,In_280,In_1597);
nor U514 (N_514,In_1793,In_1368);
or U515 (N_515,In_385,In_1574);
xnor U516 (N_516,In_176,In_976);
nor U517 (N_517,In_1678,In_2);
nor U518 (N_518,In_1301,In_464);
nand U519 (N_519,In_757,In_362);
and U520 (N_520,In_121,In_1859);
and U521 (N_521,In_1990,In_1697);
or U522 (N_522,In_399,In_1303);
and U523 (N_523,In_1420,In_48);
xnor U524 (N_524,In_321,In_901);
or U525 (N_525,In_914,In_1075);
or U526 (N_526,In_1223,In_1864);
xnor U527 (N_527,In_875,In_1507);
or U528 (N_528,In_1863,In_1111);
xor U529 (N_529,In_497,In_1036);
nand U530 (N_530,In_420,In_542);
or U531 (N_531,In_1496,In_417);
nand U532 (N_532,In_1832,In_968);
or U533 (N_533,In_151,In_1565);
nor U534 (N_534,In_1846,In_79);
nor U535 (N_535,In_50,In_812);
nor U536 (N_536,In_649,In_401);
or U537 (N_537,In_1429,In_1631);
or U538 (N_538,In_718,In_1004);
or U539 (N_539,In_1316,In_1740);
nand U540 (N_540,In_1686,In_562);
nand U541 (N_541,In_1169,In_1362);
and U542 (N_542,In_1563,In_438);
and U543 (N_543,In_1581,In_1892);
nand U544 (N_544,In_378,In_559);
or U545 (N_545,In_38,In_139);
xor U546 (N_546,In_581,In_1098);
nor U547 (N_547,In_324,In_1114);
nand U548 (N_548,In_1792,In_1158);
or U549 (N_549,In_1865,In_1392);
nand U550 (N_550,In_252,In_732);
and U551 (N_551,In_689,In_1369);
and U552 (N_552,In_1402,In_1694);
and U553 (N_553,In_964,In_1643);
nand U554 (N_554,In_1906,In_238);
nand U555 (N_555,In_229,In_823);
or U556 (N_556,In_255,In_856);
nand U557 (N_557,In_842,In_1894);
nor U558 (N_558,In_1957,In_1370);
and U559 (N_559,In_661,In_170);
or U560 (N_560,In_1026,In_1265);
and U561 (N_561,In_216,In_1077);
nand U562 (N_562,In_1401,In_289);
nor U563 (N_563,In_416,In_1295);
or U564 (N_564,In_1415,In_857);
nor U565 (N_565,In_754,In_119);
nor U566 (N_566,In_984,In_326);
nor U567 (N_567,In_758,In_1986);
xnor U568 (N_568,In_1902,In_409);
nor U569 (N_569,In_1162,In_1491);
or U570 (N_570,In_1620,In_626);
nor U571 (N_571,In_1994,In_172);
xnor U572 (N_572,In_46,In_1389);
nor U573 (N_573,In_1305,In_804);
nor U574 (N_574,In_113,In_744);
nor U575 (N_575,In_990,In_1103);
nand U576 (N_576,In_1788,In_208);
and U577 (N_577,In_1683,In_1088);
xor U578 (N_578,In_586,In_1798);
nor U579 (N_579,In_1353,In_567);
nand U580 (N_580,In_1780,In_1981);
xnor U581 (N_581,In_1219,In_311);
or U582 (N_582,In_265,In_995);
or U583 (N_583,In_1435,In_69);
nor U584 (N_584,In_1603,In_788);
nand U585 (N_585,In_391,In_500);
nor U586 (N_586,In_960,In_917);
nand U587 (N_587,In_1089,In_1748);
nand U588 (N_588,In_363,In_1160);
and U589 (N_589,In_1785,In_1674);
xor U590 (N_590,In_130,In_552);
xnor U591 (N_591,In_344,In_1333);
or U592 (N_592,In_1492,In_1772);
and U593 (N_593,In_1737,In_1266);
nor U594 (N_594,In_98,In_1930);
and U595 (N_595,In_1974,In_1995);
nor U596 (N_596,In_621,In_1531);
xnor U597 (N_597,In_1326,In_1055);
or U598 (N_598,In_853,In_1259);
and U599 (N_599,In_1411,In_1887);
nand U600 (N_600,In_750,In_1847);
nor U601 (N_601,In_827,In_1450);
and U602 (N_602,In_250,In_555);
and U603 (N_603,In_1178,In_1070);
nor U604 (N_604,In_237,In_114);
nor U605 (N_605,In_1322,In_1090);
or U606 (N_606,In_1607,In_989);
nor U607 (N_607,In_107,In_452);
nand U608 (N_608,In_1199,In_1566);
nand U609 (N_609,In_1352,In_447);
nand U610 (N_610,In_1752,In_822);
and U611 (N_611,In_1617,In_1559);
nor U612 (N_612,In_1417,In_220);
nor U613 (N_613,In_177,In_450);
or U614 (N_614,In_737,In_657);
nand U615 (N_615,In_939,In_405);
nor U616 (N_616,In_284,In_787);
nand U617 (N_617,In_1691,In_1638);
and U618 (N_618,In_186,In_924);
and U619 (N_619,In_1110,In_5);
nor U620 (N_620,In_269,In_833);
nand U621 (N_621,In_1633,In_1343);
and U622 (N_622,In_1459,In_606);
or U623 (N_623,In_143,In_908);
nor U624 (N_624,In_300,In_1202);
and U625 (N_625,In_123,In_1268);
xnor U626 (N_626,In_1938,In_1954);
xor U627 (N_627,In_1558,In_1479);
or U628 (N_628,In_778,In_1590);
or U629 (N_629,In_275,In_1028);
and U630 (N_630,In_1475,In_658);
nor U631 (N_631,In_1794,In_589);
and U632 (N_632,In_1451,In_793);
nand U633 (N_633,In_1589,In_1622);
and U634 (N_634,In_469,In_470);
and U635 (N_635,In_1311,In_927);
nand U636 (N_636,In_499,In_1713);
nand U637 (N_637,In_197,In_1462);
nor U638 (N_638,In_276,In_1056);
or U639 (N_639,In_332,In_756);
or U640 (N_640,In_1596,In_320);
nand U641 (N_641,In_1609,In_301);
or U642 (N_642,In_557,In_1419);
and U643 (N_643,In_548,In_566);
nor U644 (N_644,In_803,In_1319);
and U645 (N_645,In_863,In_67);
nor U646 (N_646,In_739,In_974);
nand U647 (N_647,In_786,In_1147);
nand U648 (N_648,In_1710,In_584);
and U649 (N_649,In_1384,In_1520);
nor U650 (N_650,In_1904,In_1395);
nor U651 (N_651,In_1937,In_93);
nand U652 (N_652,In_158,In_1828);
or U653 (N_653,In_87,In_1652);
and U654 (N_654,In_1200,In_865);
nand U655 (N_655,In_1439,In_329);
xnor U656 (N_656,In_1725,In_86);
and U657 (N_657,In_1885,In_755);
nand U658 (N_658,In_193,In_890);
nor U659 (N_659,In_1639,In_410);
nand U660 (N_660,In_1842,In_547);
and U661 (N_661,In_1300,In_307);
or U662 (N_662,In_1355,In_1977);
and U663 (N_663,In_1408,In_1069);
and U664 (N_664,In_1913,In_1677);
and U665 (N_665,In_1636,In_818);
nand U666 (N_666,In_1235,In_593);
nand U667 (N_667,In_1878,In_323);
xnor U668 (N_668,In_909,In_1782);
and U669 (N_669,In_780,In_1275);
nand U670 (N_670,In_1449,In_1854);
nand U671 (N_671,In_194,In_388);
nor U672 (N_672,In_884,In_224);
and U673 (N_673,In_752,In_1284);
or U674 (N_674,In_1246,In_251);
or U675 (N_675,In_716,In_1180);
or U676 (N_676,In_52,In_1554);
or U677 (N_677,In_1804,In_1063);
or U678 (N_678,In_955,In_1583);
and U679 (N_679,In_456,In_1397);
nor U680 (N_680,In_1481,In_442);
nand U681 (N_681,In_1331,In_515);
and U682 (N_682,In_263,In_957);
and U683 (N_683,In_1746,In_1870);
or U684 (N_684,In_766,In_1207);
nand U685 (N_685,In_830,In_712);
xor U686 (N_686,In_1037,In_771);
or U687 (N_687,In_1441,In_30);
xnor U688 (N_688,In_434,In_1294);
nand U689 (N_689,In_1941,In_204);
or U690 (N_690,In_1890,In_1613);
and U691 (N_691,In_824,In_1460);
nor U692 (N_692,In_287,In_249);
and U693 (N_693,In_1975,In_1329);
nor U694 (N_694,In_767,In_1261);
nand U695 (N_695,In_43,In_1963);
or U696 (N_696,In_232,In_720);
xnor U697 (N_697,In_206,In_1568);
xor U698 (N_698,In_820,In_1339);
nor U699 (N_699,In_1477,In_1136);
xor U700 (N_700,In_1542,In_28);
and U701 (N_701,In_106,In_1698);
nand U702 (N_702,In_1552,In_262);
or U703 (N_703,In_905,In_1544);
nand U704 (N_704,In_659,In_1153);
or U705 (N_705,In_1027,In_1105);
and U706 (N_706,In_746,In_1250);
and U707 (N_707,In_1762,In_461);
or U708 (N_708,In_1763,In_717);
and U709 (N_709,In_543,In_1430);
and U710 (N_710,In_1391,In_759);
and U711 (N_711,In_1760,In_1290);
or U712 (N_712,In_414,In_1790);
nand U713 (N_713,In_1753,In_446);
and U714 (N_714,In_159,In_651);
xnor U715 (N_715,In_678,In_1900);
nor U716 (N_716,In_1458,In_673);
nand U717 (N_717,In_694,In_1015);
xor U718 (N_718,In_1186,In_1569);
or U719 (N_719,In_433,In_1465);
xor U720 (N_720,In_1367,In_23);
xnor U721 (N_721,In_1604,In_54);
nand U722 (N_722,In_308,In_1204);
and U723 (N_723,In_886,In_233);
nor U724 (N_724,In_1308,In_1382);
and U725 (N_725,In_1644,In_100);
nor U726 (N_726,In_503,In_1705);
or U727 (N_727,In_920,In_743);
nand U728 (N_728,In_1016,In_1761);
nand U729 (N_729,In_1380,In_550);
and U730 (N_730,In_605,In_169);
nand U731 (N_731,In_1901,In_1688);
or U732 (N_732,In_90,In_973);
xor U733 (N_733,In_1190,In_709);
nand U734 (N_734,In_303,In_1841);
and U735 (N_735,In_513,In_14);
or U736 (N_736,In_622,In_831);
and U737 (N_737,In_742,In_1518);
nand U738 (N_738,In_829,In_1907);
nor U739 (N_739,In_683,In_480);
or U740 (N_740,In_1474,In_563);
xnor U741 (N_741,In_1598,In_1562);
xor U742 (N_742,In_1815,In_351);
or U743 (N_743,In_1747,In_396);
or U744 (N_744,In_1803,In_413);
xor U745 (N_745,In_639,In_473);
xor U746 (N_746,In_975,In_705);
nand U747 (N_747,In_632,In_462);
nand U748 (N_748,In_1624,In_1356);
and U749 (N_749,In_1987,In_1318);
or U750 (N_750,In_603,In_1172);
nor U751 (N_751,In_1279,In_302);
nand U752 (N_752,In_1882,In_953);
or U753 (N_753,In_7,In_1625);
xor U754 (N_754,In_390,In_1031);
xor U755 (N_755,In_776,In_686);
or U756 (N_756,In_1336,In_1264);
nand U757 (N_757,In_1701,In_1513);
or U758 (N_758,In_1461,In_431);
nand U759 (N_759,In_1849,In_1602);
nand U760 (N_760,In_245,In_850);
nor U761 (N_761,In_561,In_653);
nor U762 (N_762,In_1690,In_943);
nor U763 (N_763,In_1502,In_578);
nand U764 (N_764,In_881,In_897);
nor U765 (N_765,In_1433,In_1296);
nand U766 (N_766,In_517,In_813);
nor U767 (N_767,In_53,In_1196);
nand U768 (N_768,In_1428,In_1982);
nor U769 (N_769,In_1074,In_77);
or U770 (N_770,In_1129,In_73);
and U771 (N_771,In_521,In_1948);
and U772 (N_772,In_655,In_1985);
nor U773 (N_773,In_196,In_747);
nand U774 (N_774,In_1661,In_1971);
and U775 (N_775,In_1684,In_700);
xor U776 (N_776,In_782,In_315);
or U777 (N_777,In_1820,In_894);
and U778 (N_778,In_1735,In_1222);
nand U779 (N_779,In_828,In_29);
nor U780 (N_780,In_554,In_918);
nand U781 (N_781,In_418,In_150);
and U782 (N_782,In_1093,In_1886);
and U783 (N_783,In_931,In_998);
nand U784 (N_784,In_789,In_1774);
and U785 (N_785,In_1612,In_1549);
and U786 (N_786,In_367,In_1107);
nand U787 (N_787,In_1286,In_1314);
nor U788 (N_788,In_1783,In_1221);
xor U789 (N_789,In_1829,In_1966);
and U790 (N_790,In_988,In_1081);
and U791 (N_791,In_1656,In_982);
and U792 (N_792,In_1645,In_1976);
nor U793 (N_793,In_451,In_1214);
and U794 (N_794,In_1091,In_1059);
or U795 (N_795,In_1953,In_949);
nand U796 (N_796,In_1138,In_1920);
nor U797 (N_797,In_187,In_458);
and U798 (N_798,In_191,In_1591);
nor U799 (N_799,In_1217,In_360);
xnor U800 (N_800,In_259,In_891);
or U801 (N_801,In_736,In_295);
nor U802 (N_802,In_1306,In_1911);
or U803 (N_803,In_745,In_488);
and U804 (N_804,In_1632,In_437);
and U805 (N_805,In_1635,In_127);
nand U806 (N_806,In_1337,In_1495);
nand U807 (N_807,In_592,In_1720);
nor U808 (N_808,In_1444,In_17);
and U809 (N_809,In_1551,In_1193);
nand U810 (N_810,In_1365,In_741);
or U811 (N_811,In_1623,In_155);
nor U812 (N_812,In_375,In_1956);
or U813 (N_813,In_1503,In_641);
and U814 (N_814,In_498,In_395);
and U815 (N_815,In_1409,In_1330);
nand U816 (N_816,In_1671,In_1588);
xor U817 (N_817,In_1534,In_1545);
nand U818 (N_818,In_92,In_1944);
and U819 (N_819,In_1019,In_1092);
nand U820 (N_820,In_809,In_650);
nand U821 (N_821,In_1040,In_763);
nand U822 (N_822,In_876,In_1398);
or U823 (N_823,In_278,In_520);
and U824 (N_824,In_1926,In_24);
or U825 (N_825,In_1043,In_460);
or U826 (N_826,In_647,In_1123);
or U827 (N_827,In_851,In_489);
xnor U828 (N_828,In_1972,In_21);
nand U829 (N_829,In_1707,In_268);
nand U830 (N_830,In_1827,In_638);
or U831 (N_831,In_983,In_122);
and U832 (N_832,In_1627,In_1140);
nand U833 (N_833,In_205,In_1489);
or U834 (N_834,In_923,In_225);
nand U835 (N_835,In_1998,In_672);
and U836 (N_836,In_1281,In_703);
nand U837 (N_837,In_1498,In_1964);
nand U838 (N_838,In_1324,In_516);
nor U839 (N_839,In_1423,In_253);
or U840 (N_840,In_1350,In_1499);
and U841 (N_841,In_799,In_1567);
nand U842 (N_842,In_1403,In_337);
or U843 (N_843,In_1320,In_1538);
or U844 (N_844,In_1297,In_1425);
nor U845 (N_845,In_1702,In_27);
or U846 (N_846,In_837,In_1582);
or U847 (N_847,In_1634,In_1231);
xor U848 (N_848,In_1050,In_1148);
or U849 (N_849,In_1274,In_950);
and U850 (N_850,In_1427,In_714);
nand U851 (N_851,In_203,In_64);
or U852 (N_852,In_429,In_1253);
or U853 (N_853,In_165,In_230);
or U854 (N_854,In_1095,In_1432);
nor U855 (N_855,In_1733,In_1530);
nor U856 (N_856,In_1536,In_178);
nand U857 (N_857,In_1359,In_1313);
nand U858 (N_858,In_1168,In_180);
nor U859 (N_859,In_1150,In_290);
or U860 (N_860,In_1361,In_599);
nor U861 (N_861,In_171,In_1407);
and U862 (N_862,In_1482,In_1667);
nand U863 (N_863,In_306,In_946);
nand U864 (N_864,In_1149,In_1128);
nor U865 (N_865,In_85,In_514);
and U866 (N_866,In_1262,In_491);
nor U867 (N_867,In_228,In_751);
xor U868 (N_868,In_768,In_972);
nor U869 (N_869,In_938,In_1745);
nand U870 (N_870,In_61,In_1729);
nor U871 (N_871,In_485,In_400);
xor U872 (N_872,In_1909,In_937);
nand U873 (N_873,In_1537,In_343);
xor U874 (N_874,In_729,In_1315);
nand U875 (N_875,In_1032,In_506);
nor U876 (N_876,In_358,In_1732);
nor U877 (N_877,In_1601,In_1446);
nand U878 (N_878,In_1712,In_674);
nor U879 (N_879,In_1621,In_261);
or U880 (N_880,In_356,In_1377);
nor U881 (N_881,In_83,In_796);
nand U882 (N_882,In_1413,In_699);
and U883 (N_883,In_135,In_1578);
nand U884 (N_884,In_999,In_895);
or U885 (N_885,In_1443,In_1116);
and U886 (N_886,In_1414,In_880);
and U887 (N_887,In_1062,In_1170);
or U888 (N_888,In_1779,In_1501);
nor U889 (N_889,In_1236,In_1695);
and U890 (N_890,In_1174,In_1312);
xnor U891 (N_891,In_1009,In_1860);
and U892 (N_892,In_1399,In_1412);
nand U893 (N_893,In_1585,In_394);
xnor U894 (N_894,In_1840,In_761);
and U895 (N_895,In_1115,In_236);
or U896 (N_896,In_1918,In_1927);
or U897 (N_897,In_1682,In_611);
and U898 (N_898,In_1807,In_538);
nand U899 (N_899,In_1867,In_392);
xnor U900 (N_900,In_575,In_916);
or U901 (N_901,In_341,In_654);
xor U902 (N_902,In_1440,In_1228);
or U903 (N_903,In_1161,In_126);
and U904 (N_904,In_539,In_25);
or U905 (N_905,In_185,In_239);
nand U906 (N_906,In_770,In_279);
and U907 (N_907,In_843,In_1770);
and U908 (N_908,In_1838,In_1437);
nand U909 (N_909,In_215,In_1739);
nor U910 (N_910,In_607,In_1060);
and U911 (N_911,In_6,In_149);
or U912 (N_912,In_482,In_247);
and U913 (N_913,In_723,In_1478);
xor U914 (N_914,In_791,In_877);
nor U915 (N_915,In_376,In_1106);
and U916 (N_916,In_816,In_1064);
nor U917 (N_917,In_913,In_1457);
nor U918 (N_918,In_101,In_944);
nand U919 (N_919,In_11,In_1131);
or U920 (N_920,In_1416,In_1626);
nand U921 (N_921,In_258,In_1640);
and U922 (N_922,In_1509,In_411);
or U923 (N_923,In_1672,In_620);
nand U924 (N_924,In_293,In_455);
or U925 (N_925,In_1254,In_1610);
xnor U926 (N_926,In_1065,In_1307);
xnor U927 (N_927,In_1486,In_1001);
or U928 (N_928,In_1709,In_1453);
or U929 (N_929,In_108,In_878);
or U930 (N_930,In_1853,In_1824);
or U931 (N_931,In_213,In_1344);
and U932 (N_932,In_494,In_1741);
nand U933 (N_933,In_1298,In_701);
xnor U934 (N_934,In_1124,In_292);
nor U935 (N_935,In_217,In_1527);
nor U936 (N_936,In_1007,In_163);
nor U937 (N_937,In_1822,In_1354);
xnor U938 (N_938,In_481,In_862);
nand U939 (N_939,In_1521,In_1271);
and U940 (N_940,In_1493,In_1553);
or U941 (N_941,In_347,In_1771);
nor U942 (N_942,In_1022,In_656);
nor U943 (N_943,In_783,In_174);
nand U944 (N_944,In_1012,In_883);
and U945 (N_945,In_642,In_690);
or U946 (N_946,In_1819,In_722);
nand U947 (N_947,In_1993,In_1742);
xnor U948 (N_948,In_1194,In_1);
or U949 (N_949,In_764,In_1447);
xnor U950 (N_950,In_1614,In_1751);
or U951 (N_951,In_666,In_1668);
and U952 (N_952,In_1594,In_81);
nand U953 (N_953,In_89,In_1473);
nand U954 (N_954,In_474,In_1810);
or U955 (N_955,In_35,In_1134);
and U956 (N_956,In_748,In_992);
or U957 (N_957,In_463,In_465);
nand U958 (N_958,In_1349,In_241);
nand U959 (N_959,In_74,In_476);
and U960 (N_960,In_1371,In_1979);
nand U961 (N_961,In_738,In_1801);
nand U962 (N_962,In_1504,In_467);
xnor U963 (N_963,In_1137,In_609);
nand U964 (N_964,In_634,In_1857);
nor U965 (N_965,In_8,In_426);
nor U966 (N_966,In_1393,In_1021);
nor U967 (N_967,In_930,In_852);
and U968 (N_968,In_904,In_1135);
xnor U969 (N_969,In_129,In_1005);
or U970 (N_970,In_1044,In_1112);
nand U971 (N_971,In_1010,In_560);
nand U972 (N_972,In_41,In_82);
or U973 (N_973,In_1961,In_1983);
or U974 (N_974,In_1893,In_1800);
nand U975 (N_975,In_1463,In_1099);
nand U976 (N_976,In_945,In_900);
and U977 (N_977,In_1351,In_1654);
or U978 (N_978,In_223,In_618);
and U979 (N_979,In_1470,In_735);
and U980 (N_980,In_80,In_1011);
nor U981 (N_981,In_214,In_1176);
or U982 (N_982,In_1587,In_408);
and U983 (N_983,In_1689,In_175);
and U984 (N_984,In_645,In_1145);
nand U985 (N_985,In_1888,In_1997);
or U986 (N_986,In_1229,In_304);
nand U987 (N_987,In_604,In_495);
and U988 (N_988,In_687,In_1270);
nor U989 (N_989,In_730,In_1293);
or U990 (N_990,In_167,In_719);
nor U991 (N_991,In_679,In_1615);
or U992 (N_992,In_628,In_936);
or U993 (N_993,In_1163,In_725);
and U994 (N_994,In_579,In_309);
and U995 (N_995,In_1817,In_248);
or U996 (N_996,In_314,In_1866);
nor U997 (N_997,In_872,In_646);
nand U998 (N_998,In_472,In_222);
nand U999 (N_999,In_1257,In_1500);
nor U1000 (N_1000,In_1698,In_1714);
nand U1001 (N_1001,In_1592,In_1644);
or U1002 (N_1002,In_1238,In_1893);
nand U1003 (N_1003,In_1317,In_1729);
or U1004 (N_1004,In_1748,In_1090);
xnor U1005 (N_1005,In_717,In_1543);
or U1006 (N_1006,In_1097,In_1019);
nor U1007 (N_1007,In_21,In_283);
or U1008 (N_1008,In_1545,In_1748);
xor U1009 (N_1009,In_704,In_1583);
or U1010 (N_1010,In_1853,In_621);
and U1011 (N_1011,In_1065,In_1496);
nand U1012 (N_1012,In_638,In_1898);
nand U1013 (N_1013,In_1682,In_144);
nor U1014 (N_1014,In_284,In_110);
nand U1015 (N_1015,In_574,In_1303);
nor U1016 (N_1016,In_1335,In_78);
nand U1017 (N_1017,In_585,In_1256);
and U1018 (N_1018,In_505,In_300);
or U1019 (N_1019,In_1335,In_777);
or U1020 (N_1020,In_1950,In_1592);
nand U1021 (N_1021,In_157,In_456);
or U1022 (N_1022,In_1183,In_600);
nor U1023 (N_1023,In_42,In_721);
nand U1024 (N_1024,In_1595,In_413);
nor U1025 (N_1025,In_239,In_1012);
nand U1026 (N_1026,In_508,In_201);
xnor U1027 (N_1027,In_234,In_1602);
and U1028 (N_1028,In_377,In_1338);
nand U1029 (N_1029,In_404,In_690);
and U1030 (N_1030,In_1443,In_504);
or U1031 (N_1031,In_163,In_1840);
nand U1032 (N_1032,In_131,In_136);
and U1033 (N_1033,In_934,In_1369);
and U1034 (N_1034,In_468,In_235);
nand U1035 (N_1035,In_58,In_1635);
nand U1036 (N_1036,In_1977,In_1484);
nor U1037 (N_1037,In_817,In_233);
nand U1038 (N_1038,In_1386,In_1257);
nor U1039 (N_1039,In_1703,In_807);
and U1040 (N_1040,In_1472,In_914);
and U1041 (N_1041,In_1828,In_1956);
or U1042 (N_1042,In_840,In_1139);
or U1043 (N_1043,In_627,In_776);
nor U1044 (N_1044,In_878,In_1796);
and U1045 (N_1045,In_290,In_1128);
or U1046 (N_1046,In_793,In_1834);
nand U1047 (N_1047,In_1801,In_1119);
xor U1048 (N_1048,In_471,In_1686);
nor U1049 (N_1049,In_1088,In_1615);
nand U1050 (N_1050,In_1550,In_1620);
and U1051 (N_1051,In_1078,In_1595);
and U1052 (N_1052,In_346,In_32);
nand U1053 (N_1053,In_1805,In_1127);
or U1054 (N_1054,In_1140,In_1683);
nand U1055 (N_1055,In_1226,In_174);
nand U1056 (N_1056,In_1833,In_780);
or U1057 (N_1057,In_463,In_1260);
or U1058 (N_1058,In_348,In_1269);
and U1059 (N_1059,In_340,In_1443);
or U1060 (N_1060,In_177,In_236);
nand U1061 (N_1061,In_1042,In_1385);
and U1062 (N_1062,In_242,In_261);
or U1063 (N_1063,In_99,In_465);
and U1064 (N_1064,In_48,In_1402);
and U1065 (N_1065,In_491,In_100);
and U1066 (N_1066,In_1477,In_906);
and U1067 (N_1067,In_1109,In_1819);
or U1068 (N_1068,In_1066,In_1926);
or U1069 (N_1069,In_1102,In_1279);
and U1070 (N_1070,In_1066,In_794);
nor U1071 (N_1071,In_818,In_1611);
nor U1072 (N_1072,In_956,In_1306);
nor U1073 (N_1073,In_1155,In_788);
nand U1074 (N_1074,In_1677,In_42);
and U1075 (N_1075,In_979,In_1613);
nor U1076 (N_1076,In_1504,In_907);
or U1077 (N_1077,In_1484,In_1481);
or U1078 (N_1078,In_1045,In_275);
xnor U1079 (N_1079,In_1523,In_254);
nor U1080 (N_1080,In_1327,In_300);
or U1081 (N_1081,In_1099,In_1039);
nor U1082 (N_1082,In_944,In_90);
nand U1083 (N_1083,In_6,In_1234);
nor U1084 (N_1084,In_93,In_1941);
nand U1085 (N_1085,In_385,In_149);
and U1086 (N_1086,In_505,In_1603);
nand U1087 (N_1087,In_1271,In_483);
nor U1088 (N_1088,In_472,In_1648);
and U1089 (N_1089,In_1409,In_718);
nand U1090 (N_1090,In_1723,In_416);
nand U1091 (N_1091,In_1019,In_33);
nand U1092 (N_1092,In_1960,In_980);
nor U1093 (N_1093,In_835,In_243);
nand U1094 (N_1094,In_998,In_1441);
nand U1095 (N_1095,In_1644,In_1849);
and U1096 (N_1096,In_1811,In_568);
or U1097 (N_1097,In_1629,In_955);
nand U1098 (N_1098,In_636,In_310);
xor U1099 (N_1099,In_764,In_1002);
or U1100 (N_1100,In_15,In_477);
and U1101 (N_1101,In_1584,In_1272);
nor U1102 (N_1102,In_1633,In_984);
or U1103 (N_1103,In_1454,In_129);
or U1104 (N_1104,In_444,In_1672);
nor U1105 (N_1105,In_1786,In_1246);
or U1106 (N_1106,In_388,In_321);
and U1107 (N_1107,In_1758,In_88);
nand U1108 (N_1108,In_652,In_1208);
or U1109 (N_1109,In_259,In_1756);
nand U1110 (N_1110,In_1919,In_1227);
or U1111 (N_1111,In_244,In_73);
nand U1112 (N_1112,In_77,In_929);
nand U1113 (N_1113,In_300,In_1744);
or U1114 (N_1114,In_449,In_1241);
and U1115 (N_1115,In_978,In_815);
or U1116 (N_1116,In_1996,In_962);
nor U1117 (N_1117,In_385,In_732);
or U1118 (N_1118,In_1089,In_493);
or U1119 (N_1119,In_768,In_1904);
nand U1120 (N_1120,In_1071,In_1420);
nor U1121 (N_1121,In_972,In_1424);
nand U1122 (N_1122,In_475,In_656);
xor U1123 (N_1123,In_310,In_699);
nand U1124 (N_1124,In_1832,In_1173);
nor U1125 (N_1125,In_151,In_332);
nand U1126 (N_1126,In_1022,In_1613);
and U1127 (N_1127,In_149,In_423);
and U1128 (N_1128,In_636,In_585);
and U1129 (N_1129,In_1876,In_286);
nor U1130 (N_1130,In_1679,In_1063);
nand U1131 (N_1131,In_1215,In_1417);
nor U1132 (N_1132,In_10,In_1502);
or U1133 (N_1133,In_645,In_364);
nor U1134 (N_1134,In_454,In_8);
nand U1135 (N_1135,In_1023,In_168);
nand U1136 (N_1136,In_1040,In_1761);
nor U1137 (N_1137,In_341,In_1226);
and U1138 (N_1138,In_25,In_1162);
or U1139 (N_1139,In_115,In_99);
nand U1140 (N_1140,In_567,In_1909);
nand U1141 (N_1141,In_360,In_26);
nand U1142 (N_1142,In_1720,In_1641);
or U1143 (N_1143,In_623,In_266);
nor U1144 (N_1144,In_657,In_1146);
xor U1145 (N_1145,In_179,In_252);
nand U1146 (N_1146,In_714,In_1032);
and U1147 (N_1147,In_1117,In_1428);
xnor U1148 (N_1148,In_1335,In_123);
xnor U1149 (N_1149,In_1833,In_1309);
and U1150 (N_1150,In_297,In_436);
or U1151 (N_1151,In_1663,In_198);
and U1152 (N_1152,In_1021,In_1435);
nor U1153 (N_1153,In_678,In_1951);
nor U1154 (N_1154,In_926,In_340);
nand U1155 (N_1155,In_59,In_610);
and U1156 (N_1156,In_603,In_1063);
nor U1157 (N_1157,In_38,In_871);
and U1158 (N_1158,In_1935,In_119);
nand U1159 (N_1159,In_818,In_102);
nor U1160 (N_1160,In_1823,In_269);
or U1161 (N_1161,In_989,In_362);
and U1162 (N_1162,In_827,In_1399);
and U1163 (N_1163,In_1259,In_562);
or U1164 (N_1164,In_392,In_634);
or U1165 (N_1165,In_36,In_32);
or U1166 (N_1166,In_1398,In_1986);
nor U1167 (N_1167,In_595,In_828);
or U1168 (N_1168,In_918,In_1388);
or U1169 (N_1169,In_1473,In_255);
and U1170 (N_1170,In_321,In_1238);
xnor U1171 (N_1171,In_1084,In_1958);
nand U1172 (N_1172,In_429,In_724);
and U1173 (N_1173,In_1454,In_1795);
nor U1174 (N_1174,In_538,In_1576);
nor U1175 (N_1175,In_1186,In_1022);
nand U1176 (N_1176,In_794,In_1896);
nor U1177 (N_1177,In_1645,In_1381);
nand U1178 (N_1178,In_1573,In_1693);
or U1179 (N_1179,In_1101,In_329);
and U1180 (N_1180,In_420,In_277);
and U1181 (N_1181,In_389,In_1067);
or U1182 (N_1182,In_1822,In_1724);
nor U1183 (N_1183,In_1198,In_1161);
or U1184 (N_1184,In_1010,In_1892);
and U1185 (N_1185,In_153,In_120);
nand U1186 (N_1186,In_1455,In_799);
and U1187 (N_1187,In_1011,In_359);
nand U1188 (N_1188,In_112,In_1563);
nand U1189 (N_1189,In_1050,In_1773);
xnor U1190 (N_1190,In_297,In_939);
xnor U1191 (N_1191,In_437,In_1148);
nor U1192 (N_1192,In_323,In_1755);
and U1193 (N_1193,In_524,In_1416);
or U1194 (N_1194,In_532,In_948);
or U1195 (N_1195,In_504,In_647);
nand U1196 (N_1196,In_611,In_816);
or U1197 (N_1197,In_215,In_1363);
and U1198 (N_1198,In_1869,In_524);
and U1199 (N_1199,In_1957,In_72);
nor U1200 (N_1200,In_1823,In_1820);
and U1201 (N_1201,In_64,In_21);
nand U1202 (N_1202,In_40,In_1390);
and U1203 (N_1203,In_1775,In_1871);
nand U1204 (N_1204,In_1043,In_1585);
and U1205 (N_1205,In_619,In_1852);
xor U1206 (N_1206,In_1105,In_1373);
and U1207 (N_1207,In_240,In_1878);
and U1208 (N_1208,In_326,In_713);
nand U1209 (N_1209,In_189,In_1581);
nor U1210 (N_1210,In_409,In_1394);
or U1211 (N_1211,In_437,In_1696);
or U1212 (N_1212,In_222,In_884);
xnor U1213 (N_1213,In_1304,In_822);
or U1214 (N_1214,In_114,In_1812);
nor U1215 (N_1215,In_513,In_280);
or U1216 (N_1216,In_250,In_754);
and U1217 (N_1217,In_750,In_1582);
or U1218 (N_1218,In_1391,In_1617);
or U1219 (N_1219,In_443,In_259);
xor U1220 (N_1220,In_866,In_1430);
and U1221 (N_1221,In_1305,In_597);
nor U1222 (N_1222,In_786,In_1686);
nor U1223 (N_1223,In_871,In_1398);
nor U1224 (N_1224,In_306,In_17);
or U1225 (N_1225,In_1421,In_1953);
nand U1226 (N_1226,In_1297,In_1587);
nor U1227 (N_1227,In_361,In_1831);
and U1228 (N_1228,In_1810,In_1480);
or U1229 (N_1229,In_884,In_246);
xor U1230 (N_1230,In_1197,In_1315);
and U1231 (N_1231,In_818,In_1954);
nand U1232 (N_1232,In_1386,In_1090);
and U1233 (N_1233,In_381,In_1230);
and U1234 (N_1234,In_1090,In_1948);
nor U1235 (N_1235,In_32,In_697);
nand U1236 (N_1236,In_1519,In_1184);
nor U1237 (N_1237,In_1400,In_1203);
nor U1238 (N_1238,In_1348,In_408);
nand U1239 (N_1239,In_1216,In_1988);
and U1240 (N_1240,In_1002,In_304);
and U1241 (N_1241,In_1186,In_643);
nand U1242 (N_1242,In_705,In_23);
and U1243 (N_1243,In_81,In_659);
or U1244 (N_1244,In_1285,In_699);
nor U1245 (N_1245,In_706,In_104);
or U1246 (N_1246,In_431,In_602);
nor U1247 (N_1247,In_479,In_1036);
nor U1248 (N_1248,In_576,In_376);
or U1249 (N_1249,In_1392,In_285);
nand U1250 (N_1250,In_386,In_1104);
nand U1251 (N_1251,In_888,In_958);
and U1252 (N_1252,In_984,In_1641);
or U1253 (N_1253,In_1177,In_389);
xor U1254 (N_1254,In_542,In_30);
nor U1255 (N_1255,In_143,In_1102);
xnor U1256 (N_1256,In_1112,In_987);
and U1257 (N_1257,In_527,In_1244);
and U1258 (N_1258,In_203,In_1912);
nand U1259 (N_1259,In_503,In_1288);
or U1260 (N_1260,In_1562,In_1096);
and U1261 (N_1261,In_1584,In_1929);
and U1262 (N_1262,In_730,In_10);
nor U1263 (N_1263,In_811,In_1756);
and U1264 (N_1264,In_231,In_1044);
nand U1265 (N_1265,In_766,In_1081);
nor U1266 (N_1266,In_450,In_1254);
or U1267 (N_1267,In_1505,In_1040);
nor U1268 (N_1268,In_1002,In_1516);
nor U1269 (N_1269,In_119,In_1992);
or U1270 (N_1270,In_5,In_1086);
nand U1271 (N_1271,In_3,In_647);
and U1272 (N_1272,In_1331,In_1638);
nor U1273 (N_1273,In_1977,In_867);
xnor U1274 (N_1274,In_398,In_704);
nor U1275 (N_1275,In_1306,In_163);
nand U1276 (N_1276,In_1208,In_1850);
or U1277 (N_1277,In_311,In_1225);
nand U1278 (N_1278,In_161,In_1578);
or U1279 (N_1279,In_1447,In_1665);
nor U1280 (N_1280,In_203,In_1219);
and U1281 (N_1281,In_12,In_1253);
nand U1282 (N_1282,In_1853,In_894);
nor U1283 (N_1283,In_1027,In_1498);
and U1284 (N_1284,In_1426,In_883);
nor U1285 (N_1285,In_7,In_366);
xor U1286 (N_1286,In_1400,In_1939);
nand U1287 (N_1287,In_1021,In_1174);
xor U1288 (N_1288,In_159,In_1801);
xnor U1289 (N_1289,In_1959,In_1704);
nand U1290 (N_1290,In_277,In_957);
and U1291 (N_1291,In_1194,In_941);
nand U1292 (N_1292,In_1336,In_93);
or U1293 (N_1293,In_724,In_56);
xnor U1294 (N_1294,In_1739,In_1409);
nand U1295 (N_1295,In_716,In_1579);
xor U1296 (N_1296,In_988,In_584);
or U1297 (N_1297,In_947,In_1616);
nor U1298 (N_1298,In_46,In_1884);
and U1299 (N_1299,In_1535,In_421);
nand U1300 (N_1300,In_1442,In_1281);
or U1301 (N_1301,In_1085,In_1444);
xnor U1302 (N_1302,In_1405,In_1982);
nor U1303 (N_1303,In_595,In_1837);
or U1304 (N_1304,In_1098,In_556);
nor U1305 (N_1305,In_1936,In_1949);
and U1306 (N_1306,In_989,In_1862);
or U1307 (N_1307,In_570,In_907);
nand U1308 (N_1308,In_622,In_965);
nand U1309 (N_1309,In_239,In_196);
nand U1310 (N_1310,In_249,In_806);
nor U1311 (N_1311,In_1373,In_1564);
nor U1312 (N_1312,In_168,In_489);
and U1313 (N_1313,In_1254,In_969);
nor U1314 (N_1314,In_1689,In_1654);
nand U1315 (N_1315,In_1558,In_1148);
and U1316 (N_1316,In_612,In_398);
xor U1317 (N_1317,In_1044,In_1684);
nor U1318 (N_1318,In_1123,In_1752);
or U1319 (N_1319,In_1190,In_855);
xor U1320 (N_1320,In_879,In_1650);
or U1321 (N_1321,In_1083,In_1598);
or U1322 (N_1322,In_1607,In_842);
nor U1323 (N_1323,In_1872,In_1856);
and U1324 (N_1324,In_1191,In_309);
and U1325 (N_1325,In_913,In_1504);
nor U1326 (N_1326,In_941,In_17);
nor U1327 (N_1327,In_317,In_908);
and U1328 (N_1328,In_255,In_1017);
nor U1329 (N_1329,In_992,In_1971);
nor U1330 (N_1330,In_1013,In_92);
or U1331 (N_1331,In_23,In_591);
or U1332 (N_1332,In_305,In_768);
xor U1333 (N_1333,In_1842,In_739);
nor U1334 (N_1334,In_71,In_380);
and U1335 (N_1335,In_68,In_1557);
and U1336 (N_1336,In_158,In_1123);
xor U1337 (N_1337,In_1194,In_683);
nand U1338 (N_1338,In_1910,In_1732);
nand U1339 (N_1339,In_1735,In_820);
xor U1340 (N_1340,In_674,In_1226);
nand U1341 (N_1341,In_500,In_1756);
xnor U1342 (N_1342,In_157,In_264);
nor U1343 (N_1343,In_834,In_1833);
nor U1344 (N_1344,In_200,In_1192);
nor U1345 (N_1345,In_1163,In_1739);
and U1346 (N_1346,In_297,In_465);
xnor U1347 (N_1347,In_43,In_422);
or U1348 (N_1348,In_1949,In_1431);
or U1349 (N_1349,In_1838,In_718);
and U1350 (N_1350,In_1942,In_1128);
nand U1351 (N_1351,In_495,In_242);
or U1352 (N_1352,In_1658,In_944);
or U1353 (N_1353,In_1859,In_1636);
xnor U1354 (N_1354,In_802,In_1289);
and U1355 (N_1355,In_1317,In_1089);
xor U1356 (N_1356,In_301,In_1408);
nand U1357 (N_1357,In_1791,In_321);
nor U1358 (N_1358,In_1003,In_1992);
or U1359 (N_1359,In_1818,In_1367);
xor U1360 (N_1360,In_1641,In_1977);
or U1361 (N_1361,In_1317,In_528);
nor U1362 (N_1362,In_1979,In_1582);
nand U1363 (N_1363,In_1147,In_1586);
or U1364 (N_1364,In_1694,In_1507);
or U1365 (N_1365,In_1597,In_1805);
and U1366 (N_1366,In_1344,In_22);
or U1367 (N_1367,In_1598,In_1145);
or U1368 (N_1368,In_1287,In_457);
nor U1369 (N_1369,In_1548,In_107);
nor U1370 (N_1370,In_1837,In_565);
and U1371 (N_1371,In_1386,In_886);
and U1372 (N_1372,In_451,In_1040);
xnor U1373 (N_1373,In_703,In_1635);
or U1374 (N_1374,In_1170,In_1189);
xor U1375 (N_1375,In_139,In_1095);
xnor U1376 (N_1376,In_288,In_486);
or U1377 (N_1377,In_3,In_1722);
or U1378 (N_1378,In_948,In_1776);
nor U1379 (N_1379,In_1057,In_1139);
or U1380 (N_1380,In_68,In_988);
xor U1381 (N_1381,In_1535,In_293);
nand U1382 (N_1382,In_241,In_1581);
and U1383 (N_1383,In_937,In_545);
or U1384 (N_1384,In_1595,In_1796);
nand U1385 (N_1385,In_1480,In_32);
or U1386 (N_1386,In_316,In_1242);
or U1387 (N_1387,In_118,In_1503);
and U1388 (N_1388,In_1800,In_1268);
nor U1389 (N_1389,In_91,In_1624);
or U1390 (N_1390,In_491,In_991);
nand U1391 (N_1391,In_266,In_1407);
or U1392 (N_1392,In_1741,In_302);
nor U1393 (N_1393,In_1021,In_1917);
xor U1394 (N_1394,In_1907,In_401);
xnor U1395 (N_1395,In_5,In_1112);
nor U1396 (N_1396,In_38,In_11);
or U1397 (N_1397,In_455,In_277);
nand U1398 (N_1398,In_1438,In_696);
and U1399 (N_1399,In_1267,In_570);
nor U1400 (N_1400,In_194,In_1883);
and U1401 (N_1401,In_386,In_926);
nor U1402 (N_1402,In_313,In_254);
or U1403 (N_1403,In_1309,In_1739);
nand U1404 (N_1404,In_1890,In_1699);
nand U1405 (N_1405,In_104,In_1553);
or U1406 (N_1406,In_269,In_257);
nor U1407 (N_1407,In_1787,In_1999);
nand U1408 (N_1408,In_722,In_1914);
xnor U1409 (N_1409,In_576,In_1607);
xor U1410 (N_1410,In_516,In_556);
nor U1411 (N_1411,In_1755,In_822);
nand U1412 (N_1412,In_1626,In_127);
or U1413 (N_1413,In_585,In_1261);
or U1414 (N_1414,In_1050,In_1079);
xnor U1415 (N_1415,In_1202,In_281);
nor U1416 (N_1416,In_951,In_713);
nor U1417 (N_1417,In_653,In_0);
and U1418 (N_1418,In_874,In_1101);
nor U1419 (N_1419,In_35,In_516);
xnor U1420 (N_1420,In_1270,In_902);
nor U1421 (N_1421,In_1948,In_657);
nand U1422 (N_1422,In_581,In_14);
nor U1423 (N_1423,In_1226,In_1982);
and U1424 (N_1424,In_77,In_535);
or U1425 (N_1425,In_548,In_734);
or U1426 (N_1426,In_1410,In_1188);
nand U1427 (N_1427,In_1843,In_1886);
nor U1428 (N_1428,In_1559,In_330);
or U1429 (N_1429,In_1557,In_595);
nand U1430 (N_1430,In_1689,In_745);
or U1431 (N_1431,In_903,In_1077);
or U1432 (N_1432,In_1277,In_1450);
or U1433 (N_1433,In_374,In_726);
or U1434 (N_1434,In_1016,In_429);
or U1435 (N_1435,In_1044,In_1203);
xor U1436 (N_1436,In_870,In_139);
nor U1437 (N_1437,In_704,In_493);
nor U1438 (N_1438,In_1767,In_546);
nand U1439 (N_1439,In_658,In_699);
nor U1440 (N_1440,In_602,In_15);
nand U1441 (N_1441,In_922,In_1227);
or U1442 (N_1442,In_1778,In_1208);
or U1443 (N_1443,In_997,In_1706);
and U1444 (N_1444,In_1222,In_1272);
and U1445 (N_1445,In_483,In_640);
nor U1446 (N_1446,In_576,In_1622);
xor U1447 (N_1447,In_1334,In_1674);
nor U1448 (N_1448,In_87,In_1988);
xnor U1449 (N_1449,In_1587,In_694);
or U1450 (N_1450,In_467,In_833);
or U1451 (N_1451,In_529,In_1204);
nand U1452 (N_1452,In_1860,In_1878);
xnor U1453 (N_1453,In_1750,In_428);
nor U1454 (N_1454,In_430,In_1108);
nand U1455 (N_1455,In_76,In_1595);
nand U1456 (N_1456,In_1903,In_1498);
xor U1457 (N_1457,In_1613,In_287);
and U1458 (N_1458,In_662,In_344);
or U1459 (N_1459,In_1172,In_891);
nand U1460 (N_1460,In_452,In_650);
and U1461 (N_1461,In_373,In_1193);
nand U1462 (N_1462,In_1007,In_1091);
nor U1463 (N_1463,In_1489,In_1039);
and U1464 (N_1464,In_774,In_515);
nor U1465 (N_1465,In_1239,In_1876);
and U1466 (N_1466,In_237,In_1751);
or U1467 (N_1467,In_894,In_465);
or U1468 (N_1468,In_662,In_1638);
or U1469 (N_1469,In_1972,In_382);
nand U1470 (N_1470,In_1510,In_1967);
and U1471 (N_1471,In_54,In_1799);
and U1472 (N_1472,In_1579,In_662);
or U1473 (N_1473,In_1351,In_1487);
nand U1474 (N_1474,In_61,In_1516);
or U1475 (N_1475,In_1619,In_893);
and U1476 (N_1476,In_1335,In_1206);
and U1477 (N_1477,In_1670,In_1283);
nand U1478 (N_1478,In_1634,In_119);
and U1479 (N_1479,In_1223,In_1785);
xnor U1480 (N_1480,In_97,In_1116);
xnor U1481 (N_1481,In_1267,In_1423);
xor U1482 (N_1482,In_1638,In_1882);
nor U1483 (N_1483,In_11,In_697);
and U1484 (N_1484,In_580,In_629);
or U1485 (N_1485,In_864,In_1656);
nor U1486 (N_1486,In_1469,In_7);
and U1487 (N_1487,In_1031,In_896);
nor U1488 (N_1488,In_1278,In_1454);
or U1489 (N_1489,In_561,In_1204);
nor U1490 (N_1490,In_862,In_186);
nand U1491 (N_1491,In_1270,In_151);
nor U1492 (N_1492,In_101,In_1108);
and U1493 (N_1493,In_1271,In_1088);
or U1494 (N_1494,In_66,In_1952);
nor U1495 (N_1495,In_1572,In_1496);
nand U1496 (N_1496,In_1243,In_1724);
nand U1497 (N_1497,In_153,In_716);
nor U1498 (N_1498,In_1378,In_1190);
or U1499 (N_1499,In_191,In_653);
nor U1500 (N_1500,In_1630,In_378);
and U1501 (N_1501,In_1820,In_600);
and U1502 (N_1502,In_1468,In_343);
or U1503 (N_1503,In_25,In_1720);
nor U1504 (N_1504,In_942,In_198);
or U1505 (N_1505,In_1277,In_155);
or U1506 (N_1506,In_1868,In_1217);
or U1507 (N_1507,In_803,In_479);
nor U1508 (N_1508,In_438,In_1710);
nand U1509 (N_1509,In_1377,In_1906);
or U1510 (N_1510,In_722,In_366);
or U1511 (N_1511,In_1019,In_1266);
and U1512 (N_1512,In_857,In_1912);
and U1513 (N_1513,In_670,In_273);
nand U1514 (N_1514,In_1778,In_1987);
nor U1515 (N_1515,In_1361,In_759);
nor U1516 (N_1516,In_751,In_1669);
nor U1517 (N_1517,In_1898,In_242);
nor U1518 (N_1518,In_1052,In_1128);
nand U1519 (N_1519,In_227,In_1034);
and U1520 (N_1520,In_690,In_354);
nor U1521 (N_1521,In_380,In_1178);
nor U1522 (N_1522,In_696,In_1607);
nor U1523 (N_1523,In_1871,In_1772);
nand U1524 (N_1524,In_282,In_1398);
nand U1525 (N_1525,In_1553,In_1892);
nor U1526 (N_1526,In_1829,In_1293);
nand U1527 (N_1527,In_68,In_821);
or U1528 (N_1528,In_53,In_369);
and U1529 (N_1529,In_567,In_1622);
nor U1530 (N_1530,In_1412,In_462);
or U1531 (N_1531,In_1667,In_770);
and U1532 (N_1532,In_1076,In_1710);
nand U1533 (N_1533,In_362,In_837);
and U1534 (N_1534,In_1399,In_862);
nand U1535 (N_1535,In_486,In_884);
or U1536 (N_1536,In_188,In_1015);
and U1537 (N_1537,In_218,In_1030);
nand U1538 (N_1538,In_235,In_1275);
or U1539 (N_1539,In_1440,In_170);
and U1540 (N_1540,In_512,In_871);
or U1541 (N_1541,In_1815,In_658);
and U1542 (N_1542,In_681,In_984);
or U1543 (N_1543,In_1710,In_1015);
nand U1544 (N_1544,In_1662,In_1266);
or U1545 (N_1545,In_682,In_241);
xnor U1546 (N_1546,In_1753,In_1259);
nand U1547 (N_1547,In_335,In_557);
xnor U1548 (N_1548,In_131,In_968);
and U1549 (N_1549,In_613,In_976);
nor U1550 (N_1550,In_1533,In_1938);
or U1551 (N_1551,In_493,In_505);
nand U1552 (N_1552,In_1758,In_1405);
nor U1553 (N_1553,In_1652,In_912);
nor U1554 (N_1554,In_1104,In_1726);
nand U1555 (N_1555,In_630,In_609);
and U1556 (N_1556,In_645,In_300);
nand U1557 (N_1557,In_429,In_642);
and U1558 (N_1558,In_1641,In_481);
nand U1559 (N_1559,In_657,In_1688);
nand U1560 (N_1560,In_1252,In_1959);
and U1561 (N_1561,In_106,In_1082);
nand U1562 (N_1562,In_1327,In_113);
and U1563 (N_1563,In_979,In_779);
xnor U1564 (N_1564,In_188,In_1920);
or U1565 (N_1565,In_54,In_4);
and U1566 (N_1566,In_297,In_677);
and U1567 (N_1567,In_957,In_899);
nand U1568 (N_1568,In_764,In_37);
xor U1569 (N_1569,In_64,In_490);
nor U1570 (N_1570,In_1383,In_1307);
and U1571 (N_1571,In_45,In_1691);
nand U1572 (N_1572,In_446,In_1113);
xnor U1573 (N_1573,In_1241,In_953);
and U1574 (N_1574,In_166,In_1669);
and U1575 (N_1575,In_156,In_408);
nand U1576 (N_1576,In_403,In_1622);
or U1577 (N_1577,In_341,In_158);
nor U1578 (N_1578,In_202,In_979);
and U1579 (N_1579,In_1670,In_1456);
nor U1580 (N_1580,In_655,In_599);
or U1581 (N_1581,In_419,In_919);
xnor U1582 (N_1582,In_1174,In_1232);
or U1583 (N_1583,In_1563,In_1352);
or U1584 (N_1584,In_965,In_527);
nor U1585 (N_1585,In_518,In_1108);
and U1586 (N_1586,In_47,In_1737);
xnor U1587 (N_1587,In_1529,In_1575);
nand U1588 (N_1588,In_285,In_229);
or U1589 (N_1589,In_1072,In_70);
and U1590 (N_1590,In_752,In_36);
and U1591 (N_1591,In_1345,In_1505);
and U1592 (N_1592,In_308,In_890);
nand U1593 (N_1593,In_72,In_934);
nand U1594 (N_1594,In_507,In_187);
or U1595 (N_1595,In_989,In_1485);
nand U1596 (N_1596,In_653,In_1521);
xnor U1597 (N_1597,In_902,In_935);
or U1598 (N_1598,In_901,In_1830);
nor U1599 (N_1599,In_1179,In_1570);
nand U1600 (N_1600,In_186,In_4);
or U1601 (N_1601,In_294,In_734);
nor U1602 (N_1602,In_1310,In_175);
or U1603 (N_1603,In_650,In_1042);
or U1604 (N_1604,In_590,In_535);
or U1605 (N_1605,In_910,In_1105);
and U1606 (N_1606,In_1122,In_1067);
nand U1607 (N_1607,In_872,In_84);
nand U1608 (N_1608,In_346,In_1579);
and U1609 (N_1609,In_776,In_907);
nand U1610 (N_1610,In_51,In_1682);
nand U1611 (N_1611,In_503,In_32);
xor U1612 (N_1612,In_1466,In_50);
or U1613 (N_1613,In_1958,In_1014);
or U1614 (N_1614,In_1742,In_1380);
nor U1615 (N_1615,In_371,In_1011);
nor U1616 (N_1616,In_341,In_633);
or U1617 (N_1617,In_1795,In_1662);
nand U1618 (N_1618,In_311,In_703);
nor U1619 (N_1619,In_1687,In_485);
nor U1620 (N_1620,In_1383,In_1528);
nand U1621 (N_1621,In_1861,In_109);
and U1622 (N_1622,In_1413,In_1274);
xnor U1623 (N_1623,In_721,In_459);
and U1624 (N_1624,In_1788,In_245);
or U1625 (N_1625,In_466,In_681);
or U1626 (N_1626,In_93,In_1105);
or U1627 (N_1627,In_1566,In_401);
xor U1628 (N_1628,In_695,In_1131);
nand U1629 (N_1629,In_107,In_158);
nand U1630 (N_1630,In_1905,In_294);
or U1631 (N_1631,In_1597,In_409);
and U1632 (N_1632,In_983,In_754);
nand U1633 (N_1633,In_1832,In_1329);
nand U1634 (N_1634,In_1364,In_1013);
and U1635 (N_1635,In_1500,In_1981);
or U1636 (N_1636,In_416,In_1462);
nor U1637 (N_1637,In_929,In_1007);
xnor U1638 (N_1638,In_1505,In_532);
nor U1639 (N_1639,In_590,In_935);
or U1640 (N_1640,In_1059,In_1877);
or U1641 (N_1641,In_1132,In_1740);
xnor U1642 (N_1642,In_43,In_295);
and U1643 (N_1643,In_1022,In_1783);
and U1644 (N_1644,In_750,In_1786);
nand U1645 (N_1645,In_1481,In_162);
nor U1646 (N_1646,In_1775,In_681);
nor U1647 (N_1647,In_186,In_1469);
nand U1648 (N_1648,In_344,In_641);
nor U1649 (N_1649,In_1335,In_1720);
nand U1650 (N_1650,In_1001,In_268);
or U1651 (N_1651,In_1970,In_1073);
nand U1652 (N_1652,In_891,In_422);
nor U1653 (N_1653,In_1235,In_1913);
or U1654 (N_1654,In_1119,In_864);
nor U1655 (N_1655,In_363,In_1126);
nor U1656 (N_1656,In_1922,In_1267);
nor U1657 (N_1657,In_1485,In_1316);
or U1658 (N_1658,In_958,In_892);
or U1659 (N_1659,In_919,In_1259);
nor U1660 (N_1660,In_1212,In_681);
and U1661 (N_1661,In_911,In_1654);
xor U1662 (N_1662,In_1456,In_286);
and U1663 (N_1663,In_1964,In_1974);
nand U1664 (N_1664,In_1209,In_1752);
nand U1665 (N_1665,In_1454,In_733);
nor U1666 (N_1666,In_1803,In_1223);
or U1667 (N_1667,In_1955,In_1122);
nor U1668 (N_1668,In_938,In_1811);
nor U1669 (N_1669,In_458,In_1617);
nand U1670 (N_1670,In_1583,In_537);
or U1671 (N_1671,In_1824,In_450);
and U1672 (N_1672,In_653,In_870);
nor U1673 (N_1673,In_173,In_1617);
nor U1674 (N_1674,In_254,In_1268);
and U1675 (N_1675,In_602,In_404);
and U1676 (N_1676,In_1858,In_81);
xnor U1677 (N_1677,In_691,In_1190);
or U1678 (N_1678,In_1529,In_744);
and U1679 (N_1679,In_49,In_459);
xor U1680 (N_1680,In_247,In_1657);
and U1681 (N_1681,In_1548,In_1427);
nand U1682 (N_1682,In_1707,In_1308);
and U1683 (N_1683,In_460,In_201);
nor U1684 (N_1684,In_416,In_1780);
or U1685 (N_1685,In_1117,In_25);
or U1686 (N_1686,In_1046,In_1592);
nand U1687 (N_1687,In_719,In_971);
nand U1688 (N_1688,In_1237,In_107);
and U1689 (N_1689,In_801,In_94);
and U1690 (N_1690,In_1575,In_765);
nand U1691 (N_1691,In_1551,In_481);
or U1692 (N_1692,In_1448,In_989);
xnor U1693 (N_1693,In_1081,In_1138);
nand U1694 (N_1694,In_1046,In_1052);
nor U1695 (N_1695,In_1671,In_448);
nor U1696 (N_1696,In_24,In_1726);
and U1697 (N_1697,In_1861,In_529);
nand U1698 (N_1698,In_496,In_1023);
xor U1699 (N_1699,In_1994,In_609);
xnor U1700 (N_1700,In_824,In_589);
and U1701 (N_1701,In_1805,In_645);
or U1702 (N_1702,In_567,In_1120);
or U1703 (N_1703,In_13,In_823);
or U1704 (N_1704,In_818,In_772);
nand U1705 (N_1705,In_1603,In_320);
nor U1706 (N_1706,In_755,In_1214);
or U1707 (N_1707,In_1530,In_744);
nand U1708 (N_1708,In_1637,In_1004);
and U1709 (N_1709,In_155,In_1438);
nor U1710 (N_1710,In_1570,In_159);
xor U1711 (N_1711,In_1201,In_107);
nand U1712 (N_1712,In_373,In_755);
and U1713 (N_1713,In_329,In_1038);
nor U1714 (N_1714,In_1690,In_1366);
and U1715 (N_1715,In_1194,In_324);
nand U1716 (N_1716,In_1007,In_820);
xor U1717 (N_1717,In_1488,In_885);
and U1718 (N_1718,In_1513,In_1375);
nand U1719 (N_1719,In_1299,In_1398);
or U1720 (N_1720,In_220,In_1656);
xor U1721 (N_1721,In_536,In_1617);
nor U1722 (N_1722,In_859,In_1252);
and U1723 (N_1723,In_1319,In_1459);
nor U1724 (N_1724,In_100,In_1402);
nor U1725 (N_1725,In_1201,In_699);
and U1726 (N_1726,In_1230,In_84);
and U1727 (N_1727,In_1102,In_1778);
nand U1728 (N_1728,In_511,In_493);
xnor U1729 (N_1729,In_1320,In_889);
and U1730 (N_1730,In_1325,In_850);
or U1731 (N_1731,In_1902,In_289);
nor U1732 (N_1732,In_971,In_799);
and U1733 (N_1733,In_1842,In_205);
nand U1734 (N_1734,In_203,In_128);
or U1735 (N_1735,In_77,In_1175);
or U1736 (N_1736,In_385,In_412);
nand U1737 (N_1737,In_1868,In_674);
nor U1738 (N_1738,In_1204,In_1356);
and U1739 (N_1739,In_1667,In_361);
nand U1740 (N_1740,In_141,In_967);
nor U1741 (N_1741,In_1991,In_844);
or U1742 (N_1742,In_1188,In_1129);
nand U1743 (N_1743,In_449,In_1254);
and U1744 (N_1744,In_1386,In_643);
nand U1745 (N_1745,In_1670,In_641);
xnor U1746 (N_1746,In_1705,In_1287);
or U1747 (N_1747,In_1149,In_1840);
xor U1748 (N_1748,In_1122,In_1126);
nand U1749 (N_1749,In_673,In_781);
or U1750 (N_1750,In_1395,In_1006);
or U1751 (N_1751,In_1044,In_1390);
nand U1752 (N_1752,In_861,In_386);
or U1753 (N_1753,In_1702,In_1243);
nor U1754 (N_1754,In_1,In_830);
or U1755 (N_1755,In_393,In_537);
nand U1756 (N_1756,In_798,In_979);
nor U1757 (N_1757,In_142,In_1635);
or U1758 (N_1758,In_65,In_1799);
or U1759 (N_1759,In_1178,In_1603);
and U1760 (N_1760,In_213,In_1563);
xnor U1761 (N_1761,In_1651,In_1450);
nor U1762 (N_1762,In_1573,In_902);
nor U1763 (N_1763,In_229,In_1219);
nand U1764 (N_1764,In_1311,In_1923);
nand U1765 (N_1765,In_888,In_1907);
and U1766 (N_1766,In_862,In_415);
or U1767 (N_1767,In_11,In_383);
or U1768 (N_1768,In_607,In_625);
nand U1769 (N_1769,In_931,In_396);
nand U1770 (N_1770,In_1323,In_333);
and U1771 (N_1771,In_1733,In_1446);
or U1772 (N_1772,In_1174,In_1627);
nand U1773 (N_1773,In_168,In_831);
xor U1774 (N_1774,In_52,In_1683);
nor U1775 (N_1775,In_1502,In_1913);
or U1776 (N_1776,In_1404,In_935);
and U1777 (N_1777,In_13,In_175);
and U1778 (N_1778,In_536,In_574);
and U1779 (N_1779,In_612,In_877);
and U1780 (N_1780,In_1847,In_1217);
and U1781 (N_1781,In_440,In_748);
and U1782 (N_1782,In_1687,In_1476);
nor U1783 (N_1783,In_1774,In_345);
nand U1784 (N_1784,In_1663,In_234);
or U1785 (N_1785,In_905,In_1036);
or U1786 (N_1786,In_1787,In_1413);
or U1787 (N_1787,In_978,In_892);
nand U1788 (N_1788,In_1187,In_413);
nor U1789 (N_1789,In_1597,In_180);
xor U1790 (N_1790,In_1474,In_302);
nand U1791 (N_1791,In_1663,In_1418);
or U1792 (N_1792,In_1756,In_1283);
nor U1793 (N_1793,In_865,In_434);
and U1794 (N_1794,In_1877,In_1300);
nand U1795 (N_1795,In_230,In_1521);
nand U1796 (N_1796,In_495,In_55);
nand U1797 (N_1797,In_1154,In_1180);
or U1798 (N_1798,In_904,In_929);
and U1799 (N_1799,In_985,In_1153);
and U1800 (N_1800,In_202,In_1844);
nor U1801 (N_1801,In_847,In_834);
nand U1802 (N_1802,In_1025,In_763);
or U1803 (N_1803,In_705,In_579);
or U1804 (N_1804,In_1377,In_914);
or U1805 (N_1805,In_1431,In_345);
and U1806 (N_1806,In_1103,In_1569);
and U1807 (N_1807,In_1813,In_1963);
nand U1808 (N_1808,In_470,In_1873);
xor U1809 (N_1809,In_337,In_1290);
or U1810 (N_1810,In_330,In_1972);
or U1811 (N_1811,In_1177,In_727);
or U1812 (N_1812,In_1897,In_38);
xnor U1813 (N_1813,In_1544,In_72);
and U1814 (N_1814,In_786,In_1136);
nand U1815 (N_1815,In_138,In_371);
nor U1816 (N_1816,In_981,In_699);
xnor U1817 (N_1817,In_1937,In_1424);
nor U1818 (N_1818,In_652,In_150);
nor U1819 (N_1819,In_23,In_1596);
nor U1820 (N_1820,In_1834,In_726);
nand U1821 (N_1821,In_1239,In_1573);
nand U1822 (N_1822,In_1108,In_1808);
xnor U1823 (N_1823,In_718,In_1286);
or U1824 (N_1824,In_1556,In_1320);
and U1825 (N_1825,In_231,In_506);
nand U1826 (N_1826,In_1944,In_1026);
nand U1827 (N_1827,In_1373,In_514);
or U1828 (N_1828,In_870,In_1000);
or U1829 (N_1829,In_1515,In_1641);
nand U1830 (N_1830,In_1304,In_73);
nor U1831 (N_1831,In_1713,In_1762);
nand U1832 (N_1832,In_51,In_1636);
and U1833 (N_1833,In_85,In_233);
nand U1834 (N_1834,In_1758,In_100);
xor U1835 (N_1835,In_1778,In_402);
nor U1836 (N_1836,In_440,In_1846);
nand U1837 (N_1837,In_1272,In_1607);
nand U1838 (N_1838,In_409,In_508);
nand U1839 (N_1839,In_1769,In_294);
nand U1840 (N_1840,In_331,In_122);
and U1841 (N_1841,In_741,In_1803);
nor U1842 (N_1842,In_72,In_305);
nand U1843 (N_1843,In_362,In_1720);
or U1844 (N_1844,In_943,In_62);
and U1845 (N_1845,In_1168,In_1427);
nor U1846 (N_1846,In_166,In_92);
and U1847 (N_1847,In_1669,In_1560);
nand U1848 (N_1848,In_764,In_1602);
nand U1849 (N_1849,In_186,In_278);
nand U1850 (N_1850,In_1194,In_223);
and U1851 (N_1851,In_761,In_1939);
nor U1852 (N_1852,In_1335,In_1353);
nand U1853 (N_1853,In_1120,In_41);
nor U1854 (N_1854,In_1876,In_701);
or U1855 (N_1855,In_1740,In_1272);
or U1856 (N_1856,In_1166,In_769);
and U1857 (N_1857,In_720,In_382);
and U1858 (N_1858,In_1800,In_837);
xnor U1859 (N_1859,In_453,In_966);
and U1860 (N_1860,In_1173,In_1197);
xnor U1861 (N_1861,In_84,In_22);
or U1862 (N_1862,In_1107,In_404);
nor U1863 (N_1863,In_1355,In_1684);
nand U1864 (N_1864,In_1559,In_1377);
nor U1865 (N_1865,In_722,In_569);
and U1866 (N_1866,In_1795,In_1627);
and U1867 (N_1867,In_584,In_214);
nand U1868 (N_1868,In_1795,In_1071);
and U1869 (N_1869,In_499,In_940);
xnor U1870 (N_1870,In_1268,In_472);
nor U1871 (N_1871,In_389,In_1742);
nand U1872 (N_1872,In_1238,In_1007);
xor U1873 (N_1873,In_1270,In_468);
nor U1874 (N_1874,In_502,In_681);
nor U1875 (N_1875,In_769,In_1461);
and U1876 (N_1876,In_1428,In_1778);
nand U1877 (N_1877,In_1866,In_619);
nand U1878 (N_1878,In_1293,In_460);
and U1879 (N_1879,In_1738,In_1766);
xor U1880 (N_1880,In_295,In_1318);
nor U1881 (N_1881,In_1005,In_655);
or U1882 (N_1882,In_429,In_1916);
and U1883 (N_1883,In_658,In_788);
or U1884 (N_1884,In_712,In_286);
or U1885 (N_1885,In_382,In_1618);
and U1886 (N_1886,In_915,In_1345);
and U1887 (N_1887,In_1371,In_1844);
nor U1888 (N_1888,In_0,In_1273);
or U1889 (N_1889,In_1701,In_1954);
or U1890 (N_1890,In_559,In_1947);
or U1891 (N_1891,In_809,In_785);
nor U1892 (N_1892,In_1849,In_1600);
xnor U1893 (N_1893,In_82,In_1343);
xnor U1894 (N_1894,In_675,In_1925);
nor U1895 (N_1895,In_440,In_874);
or U1896 (N_1896,In_1898,In_610);
nand U1897 (N_1897,In_948,In_1639);
or U1898 (N_1898,In_1370,In_1764);
and U1899 (N_1899,In_472,In_321);
or U1900 (N_1900,In_1057,In_1108);
xor U1901 (N_1901,In_1400,In_111);
nand U1902 (N_1902,In_1280,In_934);
nand U1903 (N_1903,In_1231,In_1607);
or U1904 (N_1904,In_1007,In_1612);
or U1905 (N_1905,In_421,In_97);
nor U1906 (N_1906,In_1763,In_177);
or U1907 (N_1907,In_590,In_362);
or U1908 (N_1908,In_623,In_827);
and U1909 (N_1909,In_89,In_156);
nor U1910 (N_1910,In_1089,In_1438);
or U1911 (N_1911,In_271,In_704);
nor U1912 (N_1912,In_971,In_1964);
and U1913 (N_1913,In_1947,In_1897);
or U1914 (N_1914,In_81,In_1796);
nor U1915 (N_1915,In_604,In_324);
nand U1916 (N_1916,In_1426,In_547);
nor U1917 (N_1917,In_885,In_1937);
and U1918 (N_1918,In_1126,In_1510);
or U1919 (N_1919,In_1175,In_495);
and U1920 (N_1920,In_1813,In_156);
or U1921 (N_1921,In_1972,In_1736);
nand U1922 (N_1922,In_15,In_702);
and U1923 (N_1923,In_1442,In_1418);
nand U1924 (N_1924,In_623,In_1459);
nor U1925 (N_1925,In_482,In_1328);
or U1926 (N_1926,In_491,In_1448);
nor U1927 (N_1927,In_1032,In_1867);
or U1928 (N_1928,In_207,In_561);
or U1929 (N_1929,In_1691,In_694);
and U1930 (N_1930,In_1000,In_282);
xor U1931 (N_1931,In_1134,In_1577);
nand U1932 (N_1932,In_160,In_297);
nand U1933 (N_1933,In_219,In_962);
xnor U1934 (N_1934,In_790,In_1216);
xnor U1935 (N_1935,In_1615,In_596);
or U1936 (N_1936,In_1033,In_370);
nand U1937 (N_1937,In_1942,In_992);
and U1938 (N_1938,In_1191,In_379);
xor U1939 (N_1939,In_839,In_1402);
and U1940 (N_1940,In_227,In_757);
nor U1941 (N_1941,In_1134,In_1775);
or U1942 (N_1942,In_215,In_1132);
nand U1943 (N_1943,In_1230,In_1888);
or U1944 (N_1944,In_1031,In_906);
and U1945 (N_1945,In_1662,In_422);
nor U1946 (N_1946,In_1450,In_1018);
nor U1947 (N_1947,In_1633,In_881);
or U1948 (N_1948,In_481,In_1556);
or U1949 (N_1949,In_534,In_1516);
or U1950 (N_1950,In_1565,In_90);
nand U1951 (N_1951,In_1124,In_669);
or U1952 (N_1952,In_28,In_348);
xor U1953 (N_1953,In_1749,In_976);
and U1954 (N_1954,In_85,In_803);
xor U1955 (N_1955,In_1969,In_1456);
nor U1956 (N_1956,In_1437,In_1001);
and U1957 (N_1957,In_1259,In_1412);
nand U1958 (N_1958,In_1381,In_1586);
and U1959 (N_1959,In_246,In_375);
and U1960 (N_1960,In_868,In_1777);
or U1961 (N_1961,In_1147,In_527);
and U1962 (N_1962,In_926,In_324);
and U1963 (N_1963,In_1653,In_361);
nand U1964 (N_1964,In_1818,In_1841);
and U1965 (N_1965,In_503,In_1462);
nor U1966 (N_1966,In_1782,In_14);
or U1967 (N_1967,In_1273,In_541);
nand U1968 (N_1968,In_1598,In_1204);
nor U1969 (N_1969,In_446,In_1650);
nor U1970 (N_1970,In_1184,In_412);
and U1971 (N_1971,In_1596,In_1472);
and U1972 (N_1972,In_1062,In_1576);
or U1973 (N_1973,In_786,In_435);
nand U1974 (N_1974,In_1595,In_20);
nor U1975 (N_1975,In_758,In_1049);
xnor U1976 (N_1976,In_1184,In_1651);
or U1977 (N_1977,In_1469,In_431);
nor U1978 (N_1978,In_885,In_1698);
or U1979 (N_1979,In_159,In_1673);
or U1980 (N_1980,In_1350,In_1017);
nor U1981 (N_1981,In_1915,In_1115);
or U1982 (N_1982,In_440,In_1146);
nand U1983 (N_1983,In_145,In_1411);
or U1984 (N_1984,In_1459,In_211);
and U1985 (N_1985,In_1679,In_761);
or U1986 (N_1986,In_364,In_581);
nand U1987 (N_1987,In_1435,In_1993);
nand U1988 (N_1988,In_1705,In_251);
nor U1989 (N_1989,In_1341,In_1384);
or U1990 (N_1990,In_1528,In_668);
or U1991 (N_1991,In_1807,In_1724);
xor U1992 (N_1992,In_1109,In_808);
nor U1993 (N_1993,In_1322,In_1389);
nor U1994 (N_1994,In_258,In_1876);
xnor U1995 (N_1995,In_369,In_755);
and U1996 (N_1996,In_237,In_1901);
and U1997 (N_1997,In_127,In_533);
nand U1998 (N_1998,In_671,In_432);
nor U1999 (N_1999,In_341,In_635);
nor U2000 (N_2000,In_378,In_1248);
nand U2001 (N_2001,In_1521,In_1);
nor U2002 (N_2002,In_1474,In_807);
nor U2003 (N_2003,In_494,In_1401);
xor U2004 (N_2004,In_228,In_1278);
or U2005 (N_2005,In_1176,In_1988);
nor U2006 (N_2006,In_199,In_1126);
nor U2007 (N_2007,In_422,In_54);
and U2008 (N_2008,In_441,In_1942);
or U2009 (N_2009,In_551,In_1915);
nor U2010 (N_2010,In_605,In_1000);
nand U2011 (N_2011,In_294,In_625);
nand U2012 (N_2012,In_645,In_1785);
nand U2013 (N_2013,In_465,In_1688);
nor U2014 (N_2014,In_1117,In_1570);
xor U2015 (N_2015,In_1789,In_1042);
nor U2016 (N_2016,In_529,In_775);
nor U2017 (N_2017,In_1261,In_1976);
or U2018 (N_2018,In_559,In_321);
nand U2019 (N_2019,In_907,In_1287);
or U2020 (N_2020,In_1663,In_116);
nand U2021 (N_2021,In_1891,In_772);
nor U2022 (N_2022,In_1333,In_786);
and U2023 (N_2023,In_1034,In_132);
and U2024 (N_2024,In_1554,In_596);
nor U2025 (N_2025,In_1894,In_1072);
and U2026 (N_2026,In_1618,In_448);
nand U2027 (N_2027,In_690,In_510);
nor U2028 (N_2028,In_1438,In_519);
and U2029 (N_2029,In_1430,In_633);
and U2030 (N_2030,In_532,In_960);
xor U2031 (N_2031,In_530,In_1389);
nand U2032 (N_2032,In_793,In_1898);
nand U2033 (N_2033,In_801,In_1710);
xnor U2034 (N_2034,In_1017,In_204);
nand U2035 (N_2035,In_510,In_402);
or U2036 (N_2036,In_1757,In_253);
nor U2037 (N_2037,In_739,In_1671);
nand U2038 (N_2038,In_1985,In_1561);
or U2039 (N_2039,In_941,In_1716);
nand U2040 (N_2040,In_365,In_7);
nand U2041 (N_2041,In_636,In_246);
or U2042 (N_2042,In_265,In_1248);
nor U2043 (N_2043,In_1852,In_460);
nor U2044 (N_2044,In_852,In_911);
and U2045 (N_2045,In_161,In_274);
or U2046 (N_2046,In_1258,In_1899);
nor U2047 (N_2047,In_717,In_684);
nand U2048 (N_2048,In_1449,In_1895);
xor U2049 (N_2049,In_23,In_1039);
nor U2050 (N_2050,In_1342,In_895);
nor U2051 (N_2051,In_444,In_535);
nor U2052 (N_2052,In_1468,In_339);
or U2053 (N_2053,In_841,In_708);
nand U2054 (N_2054,In_1684,In_353);
xor U2055 (N_2055,In_753,In_1402);
nor U2056 (N_2056,In_1884,In_1975);
or U2057 (N_2057,In_550,In_1052);
and U2058 (N_2058,In_770,In_1022);
and U2059 (N_2059,In_270,In_910);
nand U2060 (N_2060,In_875,In_940);
nand U2061 (N_2061,In_469,In_603);
nand U2062 (N_2062,In_1406,In_1359);
nor U2063 (N_2063,In_845,In_206);
or U2064 (N_2064,In_152,In_960);
or U2065 (N_2065,In_1943,In_1901);
and U2066 (N_2066,In_1664,In_721);
or U2067 (N_2067,In_1037,In_1);
nand U2068 (N_2068,In_262,In_1219);
and U2069 (N_2069,In_845,In_596);
or U2070 (N_2070,In_1225,In_1152);
nand U2071 (N_2071,In_777,In_558);
nor U2072 (N_2072,In_1874,In_801);
and U2073 (N_2073,In_450,In_1077);
nor U2074 (N_2074,In_1086,In_617);
and U2075 (N_2075,In_110,In_473);
nor U2076 (N_2076,In_923,In_1407);
nor U2077 (N_2077,In_88,In_1614);
nor U2078 (N_2078,In_1276,In_1774);
xor U2079 (N_2079,In_891,In_1249);
or U2080 (N_2080,In_1562,In_297);
and U2081 (N_2081,In_1504,In_1479);
nor U2082 (N_2082,In_1853,In_1344);
and U2083 (N_2083,In_154,In_1559);
or U2084 (N_2084,In_1464,In_1419);
and U2085 (N_2085,In_498,In_256);
nand U2086 (N_2086,In_1260,In_1253);
and U2087 (N_2087,In_429,In_1397);
or U2088 (N_2088,In_1836,In_230);
nand U2089 (N_2089,In_583,In_1158);
or U2090 (N_2090,In_1390,In_898);
or U2091 (N_2091,In_1050,In_1389);
nor U2092 (N_2092,In_1866,In_1685);
xnor U2093 (N_2093,In_785,In_1411);
nand U2094 (N_2094,In_1891,In_1765);
nor U2095 (N_2095,In_149,In_1985);
and U2096 (N_2096,In_407,In_1293);
nand U2097 (N_2097,In_148,In_372);
or U2098 (N_2098,In_65,In_556);
or U2099 (N_2099,In_74,In_1478);
nand U2100 (N_2100,In_1154,In_1869);
nor U2101 (N_2101,In_11,In_1357);
nor U2102 (N_2102,In_1069,In_25);
nor U2103 (N_2103,In_716,In_224);
xnor U2104 (N_2104,In_895,In_1562);
nand U2105 (N_2105,In_1278,In_1740);
or U2106 (N_2106,In_1140,In_954);
or U2107 (N_2107,In_1716,In_1581);
or U2108 (N_2108,In_1249,In_1213);
and U2109 (N_2109,In_932,In_974);
and U2110 (N_2110,In_1298,In_395);
nand U2111 (N_2111,In_481,In_305);
or U2112 (N_2112,In_1010,In_585);
and U2113 (N_2113,In_1762,In_27);
xor U2114 (N_2114,In_359,In_1701);
and U2115 (N_2115,In_1018,In_770);
or U2116 (N_2116,In_331,In_1533);
nand U2117 (N_2117,In_1652,In_814);
and U2118 (N_2118,In_326,In_1659);
nor U2119 (N_2119,In_191,In_1669);
nor U2120 (N_2120,In_1831,In_827);
nor U2121 (N_2121,In_60,In_1813);
or U2122 (N_2122,In_597,In_1003);
or U2123 (N_2123,In_1857,In_258);
or U2124 (N_2124,In_152,In_447);
nand U2125 (N_2125,In_1575,In_473);
and U2126 (N_2126,In_1889,In_998);
and U2127 (N_2127,In_1787,In_543);
nor U2128 (N_2128,In_1503,In_1199);
or U2129 (N_2129,In_603,In_312);
or U2130 (N_2130,In_949,In_1037);
and U2131 (N_2131,In_481,In_1149);
nand U2132 (N_2132,In_66,In_1596);
or U2133 (N_2133,In_1288,In_1332);
and U2134 (N_2134,In_1605,In_447);
and U2135 (N_2135,In_1605,In_1541);
nor U2136 (N_2136,In_662,In_1586);
nand U2137 (N_2137,In_977,In_1062);
and U2138 (N_2138,In_908,In_1661);
or U2139 (N_2139,In_1087,In_1666);
xnor U2140 (N_2140,In_1928,In_80);
nor U2141 (N_2141,In_740,In_1889);
nor U2142 (N_2142,In_1211,In_843);
xor U2143 (N_2143,In_1992,In_22);
and U2144 (N_2144,In_370,In_1614);
and U2145 (N_2145,In_1634,In_991);
and U2146 (N_2146,In_832,In_977);
and U2147 (N_2147,In_610,In_1016);
or U2148 (N_2148,In_1768,In_1360);
and U2149 (N_2149,In_428,In_1592);
nor U2150 (N_2150,In_656,In_12);
nor U2151 (N_2151,In_800,In_261);
or U2152 (N_2152,In_209,In_514);
xnor U2153 (N_2153,In_764,In_1349);
nand U2154 (N_2154,In_426,In_73);
nor U2155 (N_2155,In_1099,In_978);
nor U2156 (N_2156,In_928,In_1090);
or U2157 (N_2157,In_1676,In_85);
nor U2158 (N_2158,In_520,In_1650);
and U2159 (N_2159,In_90,In_1762);
nand U2160 (N_2160,In_775,In_1228);
nand U2161 (N_2161,In_483,In_56);
nor U2162 (N_2162,In_273,In_1119);
nor U2163 (N_2163,In_770,In_1234);
nand U2164 (N_2164,In_315,In_832);
nor U2165 (N_2165,In_993,In_1254);
and U2166 (N_2166,In_699,In_1621);
nand U2167 (N_2167,In_182,In_731);
nand U2168 (N_2168,In_1082,In_1879);
nor U2169 (N_2169,In_534,In_892);
and U2170 (N_2170,In_1841,In_1406);
or U2171 (N_2171,In_1620,In_1046);
xor U2172 (N_2172,In_1976,In_558);
and U2173 (N_2173,In_1467,In_1571);
or U2174 (N_2174,In_1540,In_1297);
or U2175 (N_2175,In_1998,In_852);
nor U2176 (N_2176,In_1377,In_146);
or U2177 (N_2177,In_600,In_213);
nor U2178 (N_2178,In_495,In_973);
nand U2179 (N_2179,In_610,In_1829);
xnor U2180 (N_2180,In_1341,In_892);
nand U2181 (N_2181,In_1009,In_1029);
and U2182 (N_2182,In_1185,In_763);
xnor U2183 (N_2183,In_1999,In_1143);
nand U2184 (N_2184,In_193,In_1147);
and U2185 (N_2185,In_1442,In_777);
and U2186 (N_2186,In_636,In_6);
nor U2187 (N_2187,In_1754,In_1281);
nand U2188 (N_2188,In_786,In_1286);
and U2189 (N_2189,In_1867,In_1851);
or U2190 (N_2190,In_913,In_1430);
nor U2191 (N_2191,In_1689,In_1154);
nand U2192 (N_2192,In_483,In_1126);
and U2193 (N_2193,In_1908,In_1402);
nor U2194 (N_2194,In_1627,In_1022);
xnor U2195 (N_2195,In_1809,In_613);
or U2196 (N_2196,In_662,In_1965);
nor U2197 (N_2197,In_3,In_1547);
and U2198 (N_2198,In_917,In_1427);
or U2199 (N_2199,In_1569,In_644);
nand U2200 (N_2200,In_1747,In_1568);
nor U2201 (N_2201,In_789,In_1959);
and U2202 (N_2202,In_1301,In_1417);
and U2203 (N_2203,In_1332,In_1730);
or U2204 (N_2204,In_674,In_1198);
nand U2205 (N_2205,In_82,In_1424);
nand U2206 (N_2206,In_465,In_1780);
and U2207 (N_2207,In_1084,In_1113);
nand U2208 (N_2208,In_1141,In_1729);
nand U2209 (N_2209,In_828,In_947);
nor U2210 (N_2210,In_1145,In_506);
nor U2211 (N_2211,In_201,In_1834);
nor U2212 (N_2212,In_1551,In_792);
or U2213 (N_2213,In_1564,In_662);
nor U2214 (N_2214,In_1050,In_1476);
and U2215 (N_2215,In_1800,In_1910);
or U2216 (N_2216,In_1894,In_73);
nor U2217 (N_2217,In_1523,In_437);
xnor U2218 (N_2218,In_753,In_1071);
and U2219 (N_2219,In_1456,In_626);
and U2220 (N_2220,In_1574,In_1967);
xnor U2221 (N_2221,In_611,In_511);
nor U2222 (N_2222,In_1097,In_1332);
or U2223 (N_2223,In_279,In_1604);
or U2224 (N_2224,In_1416,In_1171);
nor U2225 (N_2225,In_954,In_1020);
nor U2226 (N_2226,In_1659,In_1868);
and U2227 (N_2227,In_1607,In_1858);
nor U2228 (N_2228,In_319,In_1449);
nand U2229 (N_2229,In_485,In_1824);
or U2230 (N_2230,In_586,In_532);
nand U2231 (N_2231,In_840,In_1504);
and U2232 (N_2232,In_1562,In_1641);
nand U2233 (N_2233,In_757,In_1131);
and U2234 (N_2234,In_1568,In_1195);
and U2235 (N_2235,In_215,In_90);
nand U2236 (N_2236,In_51,In_1331);
or U2237 (N_2237,In_444,In_485);
and U2238 (N_2238,In_230,In_458);
nor U2239 (N_2239,In_399,In_1468);
and U2240 (N_2240,In_866,In_318);
nor U2241 (N_2241,In_1212,In_1670);
or U2242 (N_2242,In_1379,In_474);
or U2243 (N_2243,In_1876,In_1613);
and U2244 (N_2244,In_691,In_1985);
nand U2245 (N_2245,In_1854,In_1381);
xor U2246 (N_2246,In_74,In_1813);
xnor U2247 (N_2247,In_474,In_221);
and U2248 (N_2248,In_1460,In_676);
nand U2249 (N_2249,In_973,In_28);
nand U2250 (N_2250,In_44,In_1834);
or U2251 (N_2251,In_284,In_929);
nor U2252 (N_2252,In_1821,In_891);
and U2253 (N_2253,In_1909,In_1846);
and U2254 (N_2254,In_1550,In_134);
or U2255 (N_2255,In_1994,In_1280);
nand U2256 (N_2256,In_816,In_412);
or U2257 (N_2257,In_1277,In_62);
xnor U2258 (N_2258,In_609,In_668);
xor U2259 (N_2259,In_63,In_1915);
xor U2260 (N_2260,In_1628,In_33);
and U2261 (N_2261,In_628,In_1577);
or U2262 (N_2262,In_873,In_261);
nand U2263 (N_2263,In_1546,In_54);
and U2264 (N_2264,In_257,In_1383);
or U2265 (N_2265,In_1665,In_1024);
and U2266 (N_2266,In_1263,In_1380);
and U2267 (N_2267,In_1515,In_1065);
nand U2268 (N_2268,In_1829,In_150);
nand U2269 (N_2269,In_1192,In_343);
nor U2270 (N_2270,In_132,In_163);
and U2271 (N_2271,In_227,In_188);
nand U2272 (N_2272,In_611,In_1280);
and U2273 (N_2273,In_1975,In_33);
xor U2274 (N_2274,In_321,In_499);
xnor U2275 (N_2275,In_400,In_1363);
or U2276 (N_2276,In_501,In_1048);
nand U2277 (N_2277,In_854,In_1933);
and U2278 (N_2278,In_1810,In_12);
nand U2279 (N_2279,In_1931,In_1186);
and U2280 (N_2280,In_309,In_1994);
nor U2281 (N_2281,In_777,In_1688);
nor U2282 (N_2282,In_413,In_1109);
nand U2283 (N_2283,In_1941,In_343);
nor U2284 (N_2284,In_1224,In_1866);
nand U2285 (N_2285,In_915,In_642);
and U2286 (N_2286,In_1604,In_316);
and U2287 (N_2287,In_349,In_979);
nor U2288 (N_2288,In_1877,In_1728);
and U2289 (N_2289,In_673,In_1240);
xnor U2290 (N_2290,In_1065,In_771);
nor U2291 (N_2291,In_199,In_1975);
or U2292 (N_2292,In_393,In_251);
nand U2293 (N_2293,In_1769,In_1737);
nor U2294 (N_2294,In_1705,In_29);
and U2295 (N_2295,In_849,In_19);
nand U2296 (N_2296,In_1405,In_1138);
xnor U2297 (N_2297,In_1142,In_1212);
nor U2298 (N_2298,In_1403,In_3);
or U2299 (N_2299,In_629,In_1616);
xnor U2300 (N_2300,In_888,In_506);
or U2301 (N_2301,In_38,In_1267);
nor U2302 (N_2302,In_1399,In_86);
xor U2303 (N_2303,In_1241,In_369);
nand U2304 (N_2304,In_455,In_1133);
nor U2305 (N_2305,In_1878,In_774);
nand U2306 (N_2306,In_948,In_1344);
or U2307 (N_2307,In_1741,In_862);
nor U2308 (N_2308,In_829,In_530);
xnor U2309 (N_2309,In_839,In_1683);
and U2310 (N_2310,In_1207,In_1172);
nand U2311 (N_2311,In_655,In_1496);
or U2312 (N_2312,In_324,In_436);
and U2313 (N_2313,In_1290,In_739);
and U2314 (N_2314,In_1004,In_0);
or U2315 (N_2315,In_1618,In_20);
nor U2316 (N_2316,In_1917,In_1519);
or U2317 (N_2317,In_520,In_124);
xor U2318 (N_2318,In_776,In_529);
xor U2319 (N_2319,In_1978,In_313);
nor U2320 (N_2320,In_1236,In_856);
or U2321 (N_2321,In_506,In_1485);
or U2322 (N_2322,In_555,In_152);
and U2323 (N_2323,In_90,In_737);
nand U2324 (N_2324,In_1944,In_662);
nand U2325 (N_2325,In_1753,In_1382);
nor U2326 (N_2326,In_1416,In_1090);
and U2327 (N_2327,In_433,In_857);
nand U2328 (N_2328,In_18,In_125);
nor U2329 (N_2329,In_200,In_1228);
or U2330 (N_2330,In_1247,In_1493);
and U2331 (N_2331,In_1969,In_818);
nor U2332 (N_2332,In_1198,In_1024);
or U2333 (N_2333,In_1004,In_535);
nor U2334 (N_2334,In_647,In_1678);
xor U2335 (N_2335,In_490,In_1658);
and U2336 (N_2336,In_1895,In_970);
nand U2337 (N_2337,In_1241,In_139);
nand U2338 (N_2338,In_162,In_1641);
nand U2339 (N_2339,In_513,In_1036);
nand U2340 (N_2340,In_176,In_272);
and U2341 (N_2341,In_614,In_1892);
nand U2342 (N_2342,In_1757,In_1873);
nor U2343 (N_2343,In_1291,In_1190);
nand U2344 (N_2344,In_449,In_1101);
or U2345 (N_2345,In_676,In_43);
or U2346 (N_2346,In_343,In_102);
xor U2347 (N_2347,In_324,In_1411);
or U2348 (N_2348,In_633,In_1131);
xnor U2349 (N_2349,In_1852,In_344);
or U2350 (N_2350,In_1954,In_1936);
nand U2351 (N_2351,In_552,In_1167);
nand U2352 (N_2352,In_220,In_1661);
and U2353 (N_2353,In_1957,In_511);
nand U2354 (N_2354,In_1279,In_794);
or U2355 (N_2355,In_1665,In_134);
nor U2356 (N_2356,In_1450,In_1541);
nor U2357 (N_2357,In_408,In_866);
nor U2358 (N_2358,In_1565,In_494);
or U2359 (N_2359,In_1045,In_479);
xnor U2360 (N_2360,In_1859,In_1868);
or U2361 (N_2361,In_473,In_405);
nor U2362 (N_2362,In_590,In_646);
or U2363 (N_2363,In_1881,In_1219);
nor U2364 (N_2364,In_936,In_723);
or U2365 (N_2365,In_753,In_1231);
nor U2366 (N_2366,In_1246,In_892);
and U2367 (N_2367,In_928,In_1497);
or U2368 (N_2368,In_1503,In_348);
and U2369 (N_2369,In_1029,In_1018);
and U2370 (N_2370,In_508,In_521);
nand U2371 (N_2371,In_732,In_176);
nand U2372 (N_2372,In_884,In_950);
or U2373 (N_2373,In_604,In_209);
or U2374 (N_2374,In_508,In_687);
nand U2375 (N_2375,In_1226,In_1932);
and U2376 (N_2376,In_1621,In_1027);
or U2377 (N_2377,In_838,In_1568);
xor U2378 (N_2378,In_1238,In_1190);
nor U2379 (N_2379,In_455,In_449);
or U2380 (N_2380,In_1617,In_248);
and U2381 (N_2381,In_263,In_1842);
and U2382 (N_2382,In_1877,In_312);
or U2383 (N_2383,In_1746,In_776);
nand U2384 (N_2384,In_309,In_1259);
nor U2385 (N_2385,In_1729,In_1509);
or U2386 (N_2386,In_1792,In_1121);
and U2387 (N_2387,In_287,In_418);
nand U2388 (N_2388,In_339,In_158);
nand U2389 (N_2389,In_1940,In_622);
and U2390 (N_2390,In_967,In_372);
or U2391 (N_2391,In_1966,In_65);
nand U2392 (N_2392,In_397,In_88);
and U2393 (N_2393,In_383,In_929);
xor U2394 (N_2394,In_1899,In_1879);
nor U2395 (N_2395,In_118,In_687);
or U2396 (N_2396,In_1046,In_1213);
and U2397 (N_2397,In_1617,In_1576);
or U2398 (N_2398,In_1987,In_329);
nand U2399 (N_2399,In_746,In_264);
nor U2400 (N_2400,In_1354,In_608);
and U2401 (N_2401,In_1826,In_734);
and U2402 (N_2402,In_1163,In_1809);
xor U2403 (N_2403,In_1804,In_483);
nand U2404 (N_2404,In_1744,In_975);
nor U2405 (N_2405,In_165,In_222);
or U2406 (N_2406,In_33,In_1780);
or U2407 (N_2407,In_750,In_1098);
xor U2408 (N_2408,In_1099,In_1336);
nand U2409 (N_2409,In_363,In_1861);
and U2410 (N_2410,In_1045,In_168);
nor U2411 (N_2411,In_497,In_1615);
xor U2412 (N_2412,In_1053,In_1547);
and U2413 (N_2413,In_1752,In_1264);
nor U2414 (N_2414,In_1267,In_1666);
nand U2415 (N_2415,In_445,In_1694);
or U2416 (N_2416,In_1895,In_515);
and U2417 (N_2417,In_1460,In_1606);
and U2418 (N_2418,In_1243,In_372);
and U2419 (N_2419,In_1218,In_1909);
nand U2420 (N_2420,In_1491,In_1666);
nor U2421 (N_2421,In_602,In_979);
or U2422 (N_2422,In_1930,In_1845);
and U2423 (N_2423,In_123,In_890);
nand U2424 (N_2424,In_1409,In_654);
nor U2425 (N_2425,In_1012,In_1453);
or U2426 (N_2426,In_14,In_55);
nand U2427 (N_2427,In_965,In_1519);
xor U2428 (N_2428,In_1048,In_694);
or U2429 (N_2429,In_1423,In_707);
and U2430 (N_2430,In_1187,In_1850);
nand U2431 (N_2431,In_327,In_550);
nand U2432 (N_2432,In_65,In_866);
nor U2433 (N_2433,In_145,In_1089);
xor U2434 (N_2434,In_173,In_1786);
nand U2435 (N_2435,In_1691,In_1389);
nor U2436 (N_2436,In_401,In_296);
and U2437 (N_2437,In_546,In_726);
nand U2438 (N_2438,In_247,In_654);
or U2439 (N_2439,In_1164,In_625);
nor U2440 (N_2440,In_1465,In_1328);
and U2441 (N_2441,In_1354,In_181);
or U2442 (N_2442,In_1055,In_1898);
xor U2443 (N_2443,In_1026,In_1473);
xnor U2444 (N_2444,In_917,In_1341);
or U2445 (N_2445,In_656,In_1984);
nand U2446 (N_2446,In_861,In_120);
nor U2447 (N_2447,In_828,In_655);
nand U2448 (N_2448,In_1652,In_1259);
nor U2449 (N_2449,In_981,In_257);
or U2450 (N_2450,In_1594,In_364);
xor U2451 (N_2451,In_501,In_1262);
nand U2452 (N_2452,In_1027,In_367);
and U2453 (N_2453,In_1166,In_65);
or U2454 (N_2454,In_1608,In_736);
and U2455 (N_2455,In_53,In_1514);
and U2456 (N_2456,In_1885,In_1053);
or U2457 (N_2457,In_832,In_590);
nor U2458 (N_2458,In_91,In_143);
nand U2459 (N_2459,In_688,In_576);
xnor U2460 (N_2460,In_917,In_1759);
or U2461 (N_2461,In_267,In_1811);
or U2462 (N_2462,In_879,In_249);
xnor U2463 (N_2463,In_940,In_1735);
nor U2464 (N_2464,In_104,In_371);
or U2465 (N_2465,In_608,In_369);
nor U2466 (N_2466,In_658,In_1690);
and U2467 (N_2467,In_84,In_699);
and U2468 (N_2468,In_1911,In_434);
and U2469 (N_2469,In_1086,In_691);
xor U2470 (N_2470,In_1261,In_937);
or U2471 (N_2471,In_824,In_396);
or U2472 (N_2472,In_1888,In_1829);
and U2473 (N_2473,In_851,In_467);
xor U2474 (N_2474,In_1094,In_1300);
and U2475 (N_2475,In_1048,In_902);
and U2476 (N_2476,In_601,In_1857);
nor U2477 (N_2477,In_1414,In_1039);
or U2478 (N_2478,In_1558,In_875);
nor U2479 (N_2479,In_789,In_1537);
and U2480 (N_2480,In_607,In_1974);
xor U2481 (N_2481,In_8,In_813);
xnor U2482 (N_2482,In_1962,In_158);
nor U2483 (N_2483,In_269,In_1679);
nand U2484 (N_2484,In_1851,In_725);
nor U2485 (N_2485,In_268,In_229);
and U2486 (N_2486,In_504,In_1760);
and U2487 (N_2487,In_1495,In_676);
nand U2488 (N_2488,In_1476,In_1073);
or U2489 (N_2489,In_298,In_1551);
nand U2490 (N_2490,In_1613,In_569);
nor U2491 (N_2491,In_857,In_665);
or U2492 (N_2492,In_1515,In_1634);
nand U2493 (N_2493,In_985,In_1949);
or U2494 (N_2494,In_722,In_175);
or U2495 (N_2495,In_1586,In_37);
nor U2496 (N_2496,In_1086,In_840);
nor U2497 (N_2497,In_222,In_1067);
nand U2498 (N_2498,In_611,In_1219);
nand U2499 (N_2499,In_580,In_590);
nor U2500 (N_2500,In_57,In_574);
and U2501 (N_2501,In_1442,In_914);
or U2502 (N_2502,In_421,In_922);
nor U2503 (N_2503,In_1751,In_614);
nor U2504 (N_2504,In_631,In_1755);
nor U2505 (N_2505,In_1755,In_1576);
nor U2506 (N_2506,In_1703,In_975);
nor U2507 (N_2507,In_399,In_549);
nor U2508 (N_2508,In_214,In_1685);
nand U2509 (N_2509,In_1687,In_735);
or U2510 (N_2510,In_1883,In_1379);
nor U2511 (N_2511,In_640,In_1014);
nor U2512 (N_2512,In_199,In_534);
or U2513 (N_2513,In_1192,In_1873);
xor U2514 (N_2514,In_629,In_323);
and U2515 (N_2515,In_875,In_12);
and U2516 (N_2516,In_632,In_404);
nor U2517 (N_2517,In_1688,In_1820);
and U2518 (N_2518,In_1792,In_288);
and U2519 (N_2519,In_1019,In_430);
nor U2520 (N_2520,In_1014,In_927);
nor U2521 (N_2521,In_282,In_851);
nor U2522 (N_2522,In_395,In_1260);
xor U2523 (N_2523,In_600,In_32);
or U2524 (N_2524,In_312,In_53);
nor U2525 (N_2525,In_1959,In_826);
or U2526 (N_2526,In_1983,In_63);
nor U2527 (N_2527,In_949,In_1791);
nor U2528 (N_2528,In_662,In_136);
and U2529 (N_2529,In_1387,In_217);
nor U2530 (N_2530,In_564,In_472);
nand U2531 (N_2531,In_1290,In_980);
or U2532 (N_2532,In_387,In_397);
nor U2533 (N_2533,In_648,In_501);
nand U2534 (N_2534,In_1245,In_558);
nand U2535 (N_2535,In_455,In_681);
nor U2536 (N_2536,In_135,In_0);
nand U2537 (N_2537,In_623,In_1157);
xnor U2538 (N_2538,In_1689,In_392);
nor U2539 (N_2539,In_1678,In_287);
and U2540 (N_2540,In_1868,In_923);
nor U2541 (N_2541,In_312,In_544);
and U2542 (N_2542,In_822,In_101);
and U2543 (N_2543,In_175,In_1295);
and U2544 (N_2544,In_377,In_508);
nand U2545 (N_2545,In_1648,In_1946);
nor U2546 (N_2546,In_1330,In_1943);
and U2547 (N_2547,In_9,In_843);
or U2548 (N_2548,In_643,In_1018);
and U2549 (N_2549,In_210,In_214);
nand U2550 (N_2550,In_862,In_1651);
xor U2551 (N_2551,In_1048,In_1902);
and U2552 (N_2552,In_650,In_1775);
or U2553 (N_2553,In_598,In_1610);
or U2554 (N_2554,In_561,In_1626);
and U2555 (N_2555,In_25,In_1058);
or U2556 (N_2556,In_635,In_649);
nand U2557 (N_2557,In_519,In_349);
nand U2558 (N_2558,In_29,In_878);
nor U2559 (N_2559,In_1148,In_118);
nor U2560 (N_2560,In_464,In_1892);
nand U2561 (N_2561,In_391,In_1220);
nor U2562 (N_2562,In_178,In_1473);
or U2563 (N_2563,In_1522,In_1003);
nand U2564 (N_2564,In_293,In_422);
nor U2565 (N_2565,In_994,In_523);
xor U2566 (N_2566,In_1495,In_919);
nand U2567 (N_2567,In_515,In_159);
or U2568 (N_2568,In_1110,In_212);
or U2569 (N_2569,In_777,In_161);
or U2570 (N_2570,In_1100,In_372);
or U2571 (N_2571,In_1588,In_182);
nand U2572 (N_2572,In_1566,In_211);
or U2573 (N_2573,In_74,In_5);
or U2574 (N_2574,In_1329,In_1406);
nor U2575 (N_2575,In_1837,In_90);
and U2576 (N_2576,In_161,In_1030);
xor U2577 (N_2577,In_1974,In_641);
and U2578 (N_2578,In_1172,In_556);
or U2579 (N_2579,In_497,In_386);
and U2580 (N_2580,In_1358,In_572);
xnor U2581 (N_2581,In_43,In_857);
and U2582 (N_2582,In_1683,In_1889);
or U2583 (N_2583,In_1995,In_1635);
or U2584 (N_2584,In_607,In_499);
or U2585 (N_2585,In_1187,In_62);
nor U2586 (N_2586,In_108,In_927);
and U2587 (N_2587,In_1285,In_1228);
nor U2588 (N_2588,In_1770,In_1984);
nand U2589 (N_2589,In_1563,In_583);
nor U2590 (N_2590,In_1176,In_1719);
nand U2591 (N_2591,In_1466,In_1753);
and U2592 (N_2592,In_1173,In_677);
xor U2593 (N_2593,In_1115,In_150);
nor U2594 (N_2594,In_729,In_126);
nand U2595 (N_2595,In_221,In_1907);
or U2596 (N_2596,In_1085,In_413);
and U2597 (N_2597,In_1164,In_210);
and U2598 (N_2598,In_970,In_1605);
nand U2599 (N_2599,In_1246,In_1789);
nor U2600 (N_2600,In_318,In_790);
nand U2601 (N_2601,In_1932,In_1803);
nor U2602 (N_2602,In_1472,In_845);
nand U2603 (N_2603,In_301,In_1043);
nand U2604 (N_2604,In_295,In_72);
nand U2605 (N_2605,In_1090,In_1530);
nor U2606 (N_2606,In_835,In_457);
nor U2607 (N_2607,In_171,In_1345);
xnor U2608 (N_2608,In_1917,In_307);
nand U2609 (N_2609,In_195,In_789);
and U2610 (N_2610,In_865,In_1167);
or U2611 (N_2611,In_898,In_1564);
nand U2612 (N_2612,In_391,In_1208);
nor U2613 (N_2613,In_1343,In_1148);
or U2614 (N_2614,In_218,In_1510);
and U2615 (N_2615,In_733,In_1242);
or U2616 (N_2616,In_1145,In_631);
nor U2617 (N_2617,In_1698,In_1794);
or U2618 (N_2618,In_112,In_300);
or U2619 (N_2619,In_1278,In_594);
and U2620 (N_2620,In_1493,In_1592);
and U2621 (N_2621,In_167,In_1161);
nor U2622 (N_2622,In_1377,In_738);
nand U2623 (N_2623,In_285,In_1564);
and U2624 (N_2624,In_296,In_1158);
and U2625 (N_2625,In_459,In_950);
nor U2626 (N_2626,In_262,In_529);
and U2627 (N_2627,In_1619,In_781);
nand U2628 (N_2628,In_1735,In_1623);
nor U2629 (N_2629,In_1264,In_627);
nand U2630 (N_2630,In_1119,In_1080);
and U2631 (N_2631,In_73,In_994);
xnor U2632 (N_2632,In_20,In_599);
or U2633 (N_2633,In_1460,In_211);
nand U2634 (N_2634,In_238,In_1505);
or U2635 (N_2635,In_1965,In_1527);
and U2636 (N_2636,In_535,In_516);
nand U2637 (N_2637,In_1315,In_1543);
or U2638 (N_2638,In_1865,In_1089);
nand U2639 (N_2639,In_36,In_1025);
nand U2640 (N_2640,In_782,In_92);
and U2641 (N_2641,In_530,In_1332);
nor U2642 (N_2642,In_1882,In_1740);
xnor U2643 (N_2643,In_214,In_32);
nor U2644 (N_2644,In_635,In_117);
or U2645 (N_2645,In_200,In_217);
nor U2646 (N_2646,In_1615,In_1385);
or U2647 (N_2647,In_1747,In_1202);
nor U2648 (N_2648,In_1072,In_1508);
nand U2649 (N_2649,In_1215,In_1948);
or U2650 (N_2650,In_1761,In_1111);
nor U2651 (N_2651,In_1345,In_1249);
and U2652 (N_2652,In_317,In_1253);
or U2653 (N_2653,In_1349,In_1591);
nor U2654 (N_2654,In_1073,In_712);
xor U2655 (N_2655,In_237,In_1832);
nand U2656 (N_2656,In_1261,In_305);
nand U2657 (N_2657,In_257,In_207);
nand U2658 (N_2658,In_1711,In_67);
or U2659 (N_2659,In_393,In_1522);
and U2660 (N_2660,In_784,In_1235);
nor U2661 (N_2661,In_1353,In_1556);
nor U2662 (N_2662,In_1666,In_1044);
nand U2663 (N_2663,In_1908,In_357);
or U2664 (N_2664,In_1262,In_1056);
nand U2665 (N_2665,In_193,In_1819);
nand U2666 (N_2666,In_112,In_1271);
and U2667 (N_2667,In_972,In_560);
and U2668 (N_2668,In_33,In_1755);
and U2669 (N_2669,In_1605,In_1680);
and U2670 (N_2670,In_319,In_1685);
xor U2671 (N_2671,In_1850,In_1547);
nor U2672 (N_2672,In_583,In_417);
and U2673 (N_2673,In_62,In_1810);
nor U2674 (N_2674,In_1536,In_1652);
nand U2675 (N_2675,In_1638,In_1604);
or U2676 (N_2676,In_950,In_224);
nor U2677 (N_2677,In_699,In_1749);
or U2678 (N_2678,In_892,In_1174);
and U2679 (N_2679,In_1684,In_467);
or U2680 (N_2680,In_485,In_1852);
xor U2681 (N_2681,In_212,In_199);
and U2682 (N_2682,In_1480,In_1808);
and U2683 (N_2683,In_540,In_1840);
nand U2684 (N_2684,In_1459,In_124);
or U2685 (N_2685,In_536,In_1542);
nand U2686 (N_2686,In_922,In_1032);
and U2687 (N_2687,In_1034,In_1754);
or U2688 (N_2688,In_1555,In_730);
or U2689 (N_2689,In_1923,In_1376);
and U2690 (N_2690,In_1192,In_1526);
nor U2691 (N_2691,In_753,In_981);
and U2692 (N_2692,In_900,In_702);
or U2693 (N_2693,In_268,In_1654);
or U2694 (N_2694,In_1238,In_1821);
and U2695 (N_2695,In_230,In_1559);
nor U2696 (N_2696,In_1092,In_1884);
and U2697 (N_2697,In_764,In_744);
nor U2698 (N_2698,In_1766,In_802);
or U2699 (N_2699,In_11,In_905);
or U2700 (N_2700,In_1918,In_1531);
nor U2701 (N_2701,In_1939,In_1987);
and U2702 (N_2702,In_1106,In_646);
and U2703 (N_2703,In_1461,In_509);
nor U2704 (N_2704,In_1483,In_1795);
xnor U2705 (N_2705,In_1576,In_905);
and U2706 (N_2706,In_1103,In_47);
nand U2707 (N_2707,In_1211,In_1568);
nand U2708 (N_2708,In_1668,In_735);
and U2709 (N_2709,In_633,In_1316);
nand U2710 (N_2710,In_115,In_944);
and U2711 (N_2711,In_1118,In_1790);
nor U2712 (N_2712,In_1753,In_10);
or U2713 (N_2713,In_541,In_1963);
and U2714 (N_2714,In_597,In_1950);
nor U2715 (N_2715,In_903,In_190);
nor U2716 (N_2716,In_1752,In_724);
or U2717 (N_2717,In_1741,In_602);
nand U2718 (N_2718,In_1085,In_1472);
and U2719 (N_2719,In_1239,In_1779);
nor U2720 (N_2720,In_1204,In_599);
nand U2721 (N_2721,In_1341,In_1257);
nor U2722 (N_2722,In_1844,In_272);
or U2723 (N_2723,In_905,In_173);
nor U2724 (N_2724,In_1590,In_1764);
nor U2725 (N_2725,In_1991,In_390);
nand U2726 (N_2726,In_1776,In_1920);
nor U2727 (N_2727,In_1897,In_927);
nand U2728 (N_2728,In_1346,In_1377);
xnor U2729 (N_2729,In_238,In_1419);
xor U2730 (N_2730,In_616,In_898);
and U2731 (N_2731,In_1677,In_1421);
nor U2732 (N_2732,In_545,In_1840);
and U2733 (N_2733,In_1409,In_1162);
or U2734 (N_2734,In_807,In_552);
or U2735 (N_2735,In_858,In_1849);
or U2736 (N_2736,In_1302,In_264);
xor U2737 (N_2737,In_1103,In_156);
nor U2738 (N_2738,In_1596,In_69);
or U2739 (N_2739,In_623,In_847);
or U2740 (N_2740,In_198,In_1649);
and U2741 (N_2741,In_164,In_86);
and U2742 (N_2742,In_48,In_1780);
nand U2743 (N_2743,In_631,In_1609);
nor U2744 (N_2744,In_1384,In_1327);
nor U2745 (N_2745,In_325,In_1396);
and U2746 (N_2746,In_1886,In_217);
and U2747 (N_2747,In_1110,In_1241);
nor U2748 (N_2748,In_857,In_255);
nand U2749 (N_2749,In_1398,In_1719);
nand U2750 (N_2750,In_705,In_951);
and U2751 (N_2751,In_648,In_1080);
nor U2752 (N_2752,In_643,In_772);
and U2753 (N_2753,In_1085,In_1879);
and U2754 (N_2754,In_1260,In_965);
or U2755 (N_2755,In_395,In_1139);
or U2756 (N_2756,In_1596,In_544);
or U2757 (N_2757,In_497,In_1482);
or U2758 (N_2758,In_481,In_1061);
nand U2759 (N_2759,In_1954,In_133);
nor U2760 (N_2760,In_356,In_1604);
or U2761 (N_2761,In_1773,In_1322);
nand U2762 (N_2762,In_1074,In_707);
or U2763 (N_2763,In_1947,In_912);
or U2764 (N_2764,In_504,In_1401);
or U2765 (N_2765,In_886,In_1101);
and U2766 (N_2766,In_1557,In_242);
or U2767 (N_2767,In_1156,In_315);
or U2768 (N_2768,In_258,In_1183);
or U2769 (N_2769,In_747,In_417);
nor U2770 (N_2770,In_192,In_777);
nor U2771 (N_2771,In_576,In_1438);
and U2772 (N_2772,In_1050,In_890);
nand U2773 (N_2773,In_1178,In_1285);
or U2774 (N_2774,In_590,In_181);
or U2775 (N_2775,In_1331,In_1156);
nand U2776 (N_2776,In_1862,In_435);
xnor U2777 (N_2777,In_1070,In_1566);
nor U2778 (N_2778,In_1169,In_580);
nand U2779 (N_2779,In_1260,In_991);
or U2780 (N_2780,In_284,In_564);
nor U2781 (N_2781,In_1842,In_746);
or U2782 (N_2782,In_1109,In_1731);
nor U2783 (N_2783,In_1390,In_1514);
or U2784 (N_2784,In_1183,In_143);
nor U2785 (N_2785,In_1248,In_621);
nand U2786 (N_2786,In_203,In_985);
nor U2787 (N_2787,In_917,In_956);
and U2788 (N_2788,In_1772,In_723);
nor U2789 (N_2789,In_1377,In_538);
and U2790 (N_2790,In_1491,In_349);
or U2791 (N_2791,In_813,In_1628);
nand U2792 (N_2792,In_381,In_566);
nor U2793 (N_2793,In_1499,In_1814);
or U2794 (N_2794,In_802,In_1282);
xnor U2795 (N_2795,In_1964,In_1818);
xnor U2796 (N_2796,In_183,In_316);
and U2797 (N_2797,In_1727,In_139);
xor U2798 (N_2798,In_54,In_386);
or U2799 (N_2799,In_567,In_439);
nand U2800 (N_2800,In_1805,In_473);
or U2801 (N_2801,In_1900,In_1404);
and U2802 (N_2802,In_1487,In_1156);
or U2803 (N_2803,In_1621,In_814);
nor U2804 (N_2804,In_1661,In_1125);
nand U2805 (N_2805,In_1212,In_1209);
nand U2806 (N_2806,In_444,In_317);
xnor U2807 (N_2807,In_1327,In_1742);
and U2808 (N_2808,In_1588,In_711);
xor U2809 (N_2809,In_317,In_466);
or U2810 (N_2810,In_1199,In_1660);
or U2811 (N_2811,In_1963,In_1905);
nor U2812 (N_2812,In_1180,In_1382);
nand U2813 (N_2813,In_712,In_1025);
xnor U2814 (N_2814,In_950,In_543);
nand U2815 (N_2815,In_1,In_1362);
or U2816 (N_2816,In_108,In_1816);
nor U2817 (N_2817,In_917,In_519);
nor U2818 (N_2818,In_255,In_1523);
and U2819 (N_2819,In_120,In_1777);
xnor U2820 (N_2820,In_15,In_321);
xor U2821 (N_2821,In_859,In_884);
and U2822 (N_2822,In_1163,In_1805);
nand U2823 (N_2823,In_587,In_218);
nor U2824 (N_2824,In_1203,In_1739);
nand U2825 (N_2825,In_1156,In_929);
and U2826 (N_2826,In_1104,In_1273);
nor U2827 (N_2827,In_1023,In_1606);
nor U2828 (N_2828,In_27,In_828);
or U2829 (N_2829,In_1496,In_607);
nor U2830 (N_2830,In_650,In_1809);
nand U2831 (N_2831,In_1076,In_1684);
and U2832 (N_2832,In_1621,In_1802);
and U2833 (N_2833,In_1576,In_1204);
and U2834 (N_2834,In_137,In_51);
nor U2835 (N_2835,In_269,In_319);
and U2836 (N_2836,In_641,In_845);
nand U2837 (N_2837,In_1449,In_1628);
or U2838 (N_2838,In_844,In_1269);
and U2839 (N_2839,In_1317,In_1288);
nand U2840 (N_2840,In_1221,In_1139);
nor U2841 (N_2841,In_667,In_111);
or U2842 (N_2842,In_39,In_796);
and U2843 (N_2843,In_1062,In_173);
nand U2844 (N_2844,In_1979,In_1514);
xor U2845 (N_2845,In_265,In_775);
or U2846 (N_2846,In_954,In_1451);
nor U2847 (N_2847,In_1842,In_25);
or U2848 (N_2848,In_276,In_545);
or U2849 (N_2849,In_1156,In_624);
or U2850 (N_2850,In_1126,In_223);
nor U2851 (N_2851,In_1270,In_526);
nand U2852 (N_2852,In_1420,In_209);
and U2853 (N_2853,In_432,In_733);
xnor U2854 (N_2854,In_1590,In_651);
nand U2855 (N_2855,In_1638,In_91);
xor U2856 (N_2856,In_1532,In_1516);
nor U2857 (N_2857,In_659,In_461);
or U2858 (N_2858,In_618,In_688);
or U2859 (N_2859,In_426,In_1167);
or U2860 (N_2860,In_1276,In_1153);
nand U2861 (N_2861,In_490,In_174);
nor U2862 (N_2862,In_879,In_1289);
nand U2863 (N_2863,In_343,In_1107);
or U2864 (N_2864,In_1038,In_1953);
xor U2865 (N_2865,In_1767,In_1710);
and U2866 (N_2866,In_1825,In_222);
or U2867 (N_2867,In_903,In_1728);
nand U2868 (N_2868,In_1704,In_1007);
or U2869 (N_2869,In_407,In_1991);
nand U2870 (N_2870,In_1813,In_403);
or U2871 (N_2871,In_1335,In_1043);
nor U2872 (N_2872,In_97,In_795);
xor U2873 (N_2873,In_999,In_581);
nand U2874 (N_2874,In_92,In_812);
nor U2875 (N_2875,In_977,In_1028);
or U2876 (N_2876,In_1864,In_1543);
nor U2877 (N_2877,In_1553,In_1007);
and U2878 (N_2878,In_264,In_1428);
and U2879 (N_2879,In_1461,In_324);
nand U2880 (N_2880,In_633,In_1127);
nor U2881 (N_2881,In_1007,In_1899);
nand U2882 (N_2882,In_1097,In_707);
nand U2883 (N_2883,In_1428,In_937);
and U2884 (N_2884,In_1520,In_1305);
or U2885 (N_2885,In_673,In_1228);
nand U2886 (N_2886,In_728,In_1401);
nor U2887 (N_2887,In_254,In_1026);
and U2888 (N_2888,In_1904,In_843);
and U2889 (N_2889,In_502,In_798);
or U2890 (N_2890,In_564,In_1069);
and U2891 (N_2891,In_840,In_465);
nand U2892 (N_2892,In_1331,In_613);
nand U2893 (N_2893,In_812,In_645);
or U2894 (N_2894,In_1598,In_228);
or U2895 (N_2895,In_63,In_425);
or U2896 (N_2896,In_1701,In_985);
xnor U2897 (N_2897,In_304,In_1189);
nor U2898 (N_2898,In_647,In_629);
xor U2899 (N_2899,In_1386,In_494);
nor U2900 (N_2900,In_1762,In_1492);
xnor U2901 (N_2901,In_57,In_1019);
and U2902 (N_2902,In_1188,In_1);
nor U2903 (N_2903,In_1143,In_483);
nand U2904 (N_2904,In_918,In_3);
nand U2905 (N_2905,In_1908,In_297);
xor U2906 (N_2906,In_1818,In_705);
nand U2907 (N_2907,In_1593,In_1693);
nand U2908 (N_2908,In_1925,In_888);
and U2909 (N_2909,In_1737,In_1068);
nand U2910 (N_2910,In_1652,In_1840);
and U2911 (N_2911,In_33,In_1972);
and U2912 (N_2912,In_109,In_337);
nand U2913 (N_2913,In_1395,In_196);
nor U2914 (N_2914,In_1047,In_1998);
and U2915 (N_2915,In_800,In_205);
and U2916 (N_2916,In_1832,In_1897);
xor U2917 (N_2917,In_812,In_562);
nor U2918 (N_2918,In_1958,In_772);
and U2919 (N_2919,In_457,In_1269);
nor U2920 (N_2920,In_1907,In_146);
nand U2921 (N_2921,In_1925,In_938);
nand U2922 (N_2922,In_1348,In_1720);
or U2923 (N_2923,In_493,In_1193);
nand U2924 (N_2924,In_1589,In_1272);
xnor U2925 (N_2925,In_1095,In_910);
nor U2926 (N_2926,In_652,In_1742);
nand U2927 (N_2927,In_713,In_1703);
or U2928 (N_2928,In_310,In_451);
and U2929 (N_2929,In_1734,In_636);
and U2930 (N_2930,In_282,In_20);
nand U2931 (N_2931,In_205,In_1589);
nand U2932 (N_2932,In_1500,In_936);
nand U2933 (N_2933,In_990,In_389);
nand U2934 (N_2934,In_1226,In_326);
xnor U2935 (N_2935,In_1594,In_462);
or U2936 (N_2936,In_1063,In_17);
and U2937 (N_2937,In_375,In_615);
or U2938 (N_2938,In_141,In_518);
nor U2939 (N_2939,In_1715,In_1867);
or U2940 (N_2940,In_788,In_81);
nand U2941 (N_2941,In_1057,In_874);
nand U2942 (N_2942,In_1544,In_328);
or U2943 (N_2943,In_299,In_1229);
nor U2944 (N_2944,In_61,In_426);
or U2945 (N_2945,In_957,In_1251);
nand U2946 (N_2946,In_820,In_835);
nand U2947 (N_2947,In_1293,In_1783);
and U2948 (N_2948,In_143,In_680);
nor U2949 (N_2949,In_1527,In_507);
nand U2950 (N_2950,In_1109,In_477);
nor U2951 (N_2951,In_1371,In_1142);
nor U2952 (N_2952,In_1573,In_968);
nor U2953 (N_2953,In_312,In_723);
or U2954 (N_2954,In_1461,In_492);
or U2955 (N_2955,In_1356,In_1811);
xnor U2956 (N_2956,In_1152,In_1);
or U2957 (N_2957,In_868,In_210);
and U2958 (N_2958,In_188,In_862);
nor U2959 (N_2959,In_86,In_622);
nand U2960 (N_2960,In_355,In_1356);
and U2961 (N_2961,In_200,In_1222);
and U2962 (N_2962,In_1308,In_230);
xnor U2963 (N_2963,In_1031,In_402);
or U2964 (N_2964,In_154,In_1068);
and U2965 (N_2965,In_291,In_932);
and U2966 (N_2966,In_1652,In_1428);
and U2967 (N_2967,In_1067,In_874);
nand U2968 (N_2968,In_160,In_920);
or U2969 (N_2969,In_535,In_1040);
or U2970 (N_2970,In_885,In_1036);
or U2971 (N_2971,In_32,In_102);
nor U2972 (N_2972,In_1473,In_1114);
xnor U2973 (N_2973,In_896,In_1519);
nor U2974 (N_2974,In_1047,In_1800);
nand U2975 (N_2975,In_865,In_1340);
or U2976 (N_2976,In_1157,In_70);
xor U2977 (N_2977,In_1159,In_607);
and U2978 (N_2978,In_526,In_911);
nor U2979 (N_2979,In_1714,In_1607);
nand U2980 (N_2980,In_982,In_1473);
and U2981 (N_2981,In_1057,In_667);
nor U2982 (N_2982,In_934,In_1270);
and U2983 (N_2983,In_1212,In_144);
nand U2984 (N_2984,In_47,In_1136);
and U2985 (N_2985,In_1678,In_1639);
nor U2986 (N_2986,In_1384,In_1353);
nor U2987 (N_2987,In_428,In_1742);
nand U2988 (N_2988,In_1295,In_1849);
or U2989 (N_2989,In_966,In_466);
nand U2990 (N_2990,In_1979,In_1635);
nand U2991 (N_2991,In_1971,In_346);
or U2992 (N_2992,In_1873,In_596);
and U2993 (N_2993,In_583,In_745);
and U2994 (N_2994,In_989,In_1840);
nor U2995 (N_2995,In_1365,In_478);
xor U2996 (N_2996,In_1557,In_1189);
and U2997 (N_2997,In_1510,In_894);
nand U2998 (N_2998,In_136,In_502);
nand U2999 (N_2999,In_246,In_823);
or U3000 (N_3000,In_110,In_1742);
nor U3001 (N_3001,In_1075,In_363);
nor U3002 (N_3002,In_1841,In_973);
nor U3003 (N_3003,In_1583,In_1246);
or U3004 (N_3004,In_336,In_1428);
nand U3005 (N_3005,In_1697,In_202);
nand U3006 (N_3006,In_1769,In_564);
xor U3007 (N_3007,In_843,In_822);
and U3008 (N_3008,In_1843,In_991);
and U3009 (N_3009,In_1814,In_1610);
and U3010 (N_3010,In_22,In_1282);
nor U3011 (N_3011,In_123,In_456);
nand U3012 (N_3012,In_1027,In_495);
xnor U3013 (N_3013,In_1627,In_1430);
xnor U3014 (N_3014,In_1668,In_1839);
or U3015 (N_3015,In_1611,In_1058);
nand U3016 (N_3016,In_13,In_143);
nor U3017 (N_3017,In_993,In_1900);
nor U3018 (N_3018,In_1936,In_1543);
and U3019 (N_3019,In_1675,In_1166);
nand U3020 (N_3020,In_984,In_637);
and U3021 (N_3021,In_155,In_380);
nor U3022 (N_3022,In_1561,In_889);
nor U3023 (N_3023,In_400,In_814);
nand U3024 (N_3024,In_100,In_1582);
nand U3025 (N_3025,In_905,In_1212);
or U3026 (N_3026,In_1459,In_958);
xor U3027 (N_3027,In_1011,In_1799);
nand U3028 (N_3028,In_984,In_1132);
nand U3029 (N_3029,In_928,In_1629);
nor U3030 (N_3030,In_670,In_1561);
nor U3031 (N_3031,In_3,In_1978);
nor U3032 (N_3032,In_1781,In_1825);
or U3033 (N_3033,In_802,In_318);
or U3034 (N_3034,In_1818,In_58);
nor U3035 (N_3035,In_176,In_1263);
and U3036 (N_3036,In_313,In_276);
or U3037 (N_3037,In_1707,In_751);
nand U3038 (N_3038,In_1637,In_162);
or U3039 (N_3039,In_869,In_1805);
nor U3040 (N_3040,In_254,In_1861);
or U3041 (N_3041,In_1969,In_1572);
nand U3042 (N_3042,In_1491,In_1262);
nand U3043 (N_3043,In_688,In_97);
or U3044 (N_3044,In_396,In_967);
or U3045 (N_3045,In_796,In_1848);
and U3046 (N_3046,In_345,In_1854);
nand U3047 (N_3047,In_721,In_924);
and U3048 (N_3048,In_1153,In_479);
or U3049 (N_3049,In_382,In_369);
nor U3050 (N_3050,In_1886,In_1939);
nor U3051 (N_3051,In_290,In_847);
nor U3052 (N_3052,In_1479,In_1360);
or U3053 (N_3053,In_1748,In_699);
or U3054 (N_3054,In_277,In_1505);
nand U3055 (N_3055,In_206,In_970);
nand U3056 (N_3056,In_428,In_1375);
nand U3057 (N_3057,In_1992,In_140);
and U3058 (N_3058,In_1638,In_521);
nand U3059 (N_3059,In_632,In_414);
and U3060 (N_3060,In_1130,In_899);
or U3061 (N_3061,In_1346,In_1607);
and U3062 (N_3062,In_392,In_322);
nand U3063 (N_3063,In_1729,In_112);
nand U3064 (N_3064,In_1259,In_993);
xor U3065 (N_3065,In_1118,In_1953);
and U3066 (N_3066,In_349,In_1993);
and U3067 (N_3067,In_1201,In_162);
or U3068 (N_3068,In_756,In_1842);
and U3069 (N_3069,In_347,In_556);
or U3070 (N_3070,In_1557,In_1289);
nand U3071 (N_3071,In_752,In_1971);
nand U3072 (N_3072,In_1111,In_1966);
nand U3073 (N_3073,In_427,In_675);
and U3074 (N_3074,In_366,In_1908);
and U3075 (N_3075,In_810,In_1782);
and U3076 (N_3076,In_1165,In_1495);
and U3077 (N_3077,In_1214,In_1309);
nand U3078 (N_3078,In_1484,In_1884);
and U3079 (N_3079,In_768,In_1806);
and U3080 (N_3080,In_622,In_1303);
nor U3081 (N_3081,In_1030,In_1972);
nor U3082 (N_3082,In_1269,In_1172);
nand U3083 (N_3083,In_199,In_1513);
nor U3084 (N_3084,In_994,In_1698);
nor U3085 (N_3085,In_1442,In_951);
or U3086 (N_3086,In_937,In_1608);
or U3087 (N_3087,In_1862,In_1982);
and U3088 (N_3088,In_861,In_841);
and U3089 (N_3089,In_559,In_200);
nand U3090 (N_3090,In_1433,In_244);
or U3091 (N_3091,In_1654,In_1950);
and U3092 (N_3092,In_1893,In_773);
nor U3093 (N_3093,In_854,In_1279);
nor U3094 (N_3094,In_1481,In_1366);
xor U3095 (N_3095,In_196,In_1089);
xnor U3096 (N_3096,In_242,In_40);
and U3097 (N_3097,In_513,In_835);
and U3098 (N_3098,In_172,In_1479);
nand U3099 (N_3099,In_1667,In_1566);
and U3100 (N_3100,In_1888,In_1371);
and U3101 (N_3101,In_8,In_675);
and U3102 (N_3102,In_780,In_269);
nand U3103 (N_3103,In_1316,In_1475);
and U3104 (N_3104,In_202,In_622);
and U3105 (N_3105,In_707,In_1479);
and U3106 (N_3106,In_1148,In_707);
nor U3107 (N_3107,In_1774,In_842);
nand U3108 (N_3108,In_469,In_265);
nor U3109 (N_3109,In_1302,In_1193);
nand U3110 (N_3110,In_1687,In_479);
nor U3111 (N_3111,In_1800,In_824);
nand U3112 (N_3112,In_55,In_366);
or U3113 (N_3113,In_1740,In_136);
or U3114 (N_3114,In_948,In_630);
nand U3115 (N_3115,In_816,In_1987);
or U3116 (N_3116,In_1826,In_1227);
nor U3117 (N_3117,In_1239,In_919);
xor U3118 (N_3118,In_528,In_1066);
and U3119 (N_3119,In_1942,In_1066);
and U3120 (N_3120,In_1676,In_1027);
xnor U3121 (N_3121,In_72,In_801);
or U3122 (N_3122,In_1678,In_1781);
nor U3123 (N_3123,In_1180,In_1935);
or U3124 (N_3124,In_806,In_114);
xnor U3125 (N_3125,In_1,In_107);
and U3126 (N_3126,In_1944,In_676);
nor U3127 (N_3127,In_1432,In_450);
and U3128 (N_3128,In_1694,In_712);
xor U3129 (N_3129,In_970,In_579);
or U3130 (N_3130,In_440,In_1907);
nor U3131 (N_3131,In_792,In_959);
nor U3132 (N_3132,In_732,In_1835);
xor U3133 (N_3133,In_462,In_1554);
and U3134 (N_3134,In_1236,In_829);
and U3135 (N_3135,In_59,In_1618);
or U3136 (N_3136,In_400,In_148);
or U3137 (N_3137,In_1813,In_969);
and U3138 (N_3138,In_549,In_51);
nor U3139 (N_3139,In_1411,In_1464);
nor U3140 (N_3140,In_936,In_1344);
nand U3141 (N_3141,In_1864,In_971);
nand U3142 (N_3142,In_1589,In_1865);
or U3143 (N_3143,In_1313,In_1355);
nor U3144 (N_3144,In_1366,In_1373);
and U3145 (N_3145,In_769,In_1366);
nand U3146 (N_3146,In_1114,In_1859);
or U3147 (N_3147,In_1942,In_1679);
nand U3148 (N_3148,In_1619,In_1487);
and U3149 (N_3149,In_1632,In_1243);
or U3150 (N_3150,In_305,In_1018);
nand U3151 (N_3151,In_1553,In_491);
nor U3152 (N_3152,In_716,In_1574);
and U3153 (N_3153,In_666,In_756);
nand U3154 (N_3154,In_1152,In_1290);
and U3155 (N_3155,In_1103,In_1124);
nor U3156 (N_3156,In_695,In_1732);
and U3157 (N_3157,In_1167,In_1669);
nand U3158 (N_3158,In_687,In_314);
xnor U3159 (N_3159,In_1982,In_1685);
xor U3160 (N_3160,In_1086,In_1418);
and U3161 (N_3161,In_1494,In_211);
nor U3162 (N_3162,In_1812,In_1251);
or U3163 (N_3163,In_1290,In_315);
nor U3164 (N_3164,In_485,In_1710);
nor U3165 (N_3165,In_106,In_1688);
and U3166 (N_3166,In_108,In_420);
nor U3167 (N_3167,In_1359,In_1896);
nor U3168 (N_3168,In_603,In_1350);
nor U3169 (N_3169,In_520,In_1130);
or U3170 (N_3170,In_71,In_899);
nor U3171 (N_3171,In_1050,In_1408);
nor U3172 (N_3172,In_1740,In_1612);
and U3173 (N_3173,In_850,In_1439);
or U3174 (N_3174,In_1904,In_841);
nand U3175 (N_3175,In_954,In_320);
nor U3176 (N_3176,In_1545,In_1509);
nand U3177 (N_3177,In_1985,In_1481);
and U3178 (N_3178,In_133,In_982);
nor U3179 (N_3179,In_1688,In_53);
or U3180 (N_3180,In_699,In_364);
nor U3181 (N_3181,In_1096,In_1484);
and U3182 (N_3182,In_277,In_254);
and U3183 (N_3183,In_1668,In_1942);
and U3184 (N_3184,In_1744,In_1176);
nor U3185 (N_3185,In_1543,In_150);
or U3186 (N_3186,In_1638,In_1599);
and U3187 (N_3187,In_177,In_715);
xnor U3188 (N_3188,In_401,In_318);
or U3189 (N_3189,In_1265,In_1849);
xnor U3190 (N_3190,In_426,In_493);
nand U3191 (N_3191,In_420,In_898);
nor U3192 (N_3192,In_998,In_1303);
nor U3193 (N_3193,In_1370,In_588);
nand U3194 (N_3194,In_1708,In_783);
or U3195 (N_3195,In_919,In_1560);
or U3196 (N_3196,In_1438,In_864);
nand U3197 (N_3197,In_429,In_681);
xor U3198 (N_3198,In_330,In_1825);
or U3199 (N_3199,In_875,In_1289);
nand U3200 (N_3200,In_1257,In_801);
or U3201 (N_3201,In_1972,In_782);
and U3202 (N_3202,In_60,In_245);
nand U3203 (N_3203,In_208,In_556);
or U3204 (N_3204,In_1820,In_1812);
xnor U3205 (N_3205,In_1970,In_568);
or U3206 (N_3206,In_1027,In_1114);
xor U3207 (N_3207,In_1318,In_1742);
xor U3208 (N_3208,In_1266,In_1925);
nand U3209 (N_3209,In_557,In_548);
nand U3210 (N_3210,In_1098,In_164);
xnor U3211 (N_3211,In_1866,In_450);
or U3212 (N_3212,In_764,In_1819);
xnor U3213 (N_3213,In_1749,In_1984);
nor U3214 (N_3214,In_707,In_1454);
or U3215 (N_3215,In_722,In_648);
or U3216 (N_3216,In_1254,In_429);
nand U3217 (N_3217,In_303,In_1738);
and U3218 (N_3218,In_1428,In_391);
nand U3219 (N_3219,In_1086,In_736);
or U3220 (N_3220,In_1255,In_1910);
nand U3221 (N_3221,In_43,In_1311);
xor U3222 (N_3222,In_1663,In_1894);
or U3223 (N_3223,In_976,In_944);
or U3224 (N_3224,In_1497,In_279);
and U3225 (N_3225,In_146,In_754);
nand U3226 (N_3226,In_1759,In_533);
xnor U3227 (N_3227,In_257,In_1942);
nand U3228 (N_3228,In_119,In_99);
xor U3229 (N_3229,In_936,In_1098);
or U3230 (N_3230,In_651,In_1496);
and U3231 (N_3231,In_1661,In_196);
or U3232 (N_3232,In_1866,In_1951);
xor U3233 (N_3233,In_700,In_1444);
or U3234 (N_3234,In_1503,In_1208);
nor U3235 (N_3235,In_964,In_1235);
or U3236 (N_3236,In_919,In_1297);
xor U3237 (N_3237,In_1792,In_1075);
or U3238 (N_3238,In_1922,In_713);
xnor U3239 (N_3239,In_899,In_1538);
xnor U3240 (N_3240,In_1946,In_1609);
nor U3241 (N_3241,In_1066,In_1084);
xor U3242 (N_3242,In_854,In_512);
and U3243 (N_3243,In_249,In_1923);
nor U3244 (N_3244,In_309,In_391);
nor U3245 (N_3245,In_1627,In_776);
nand U3246 (N_3246,In_880,In_1100);
and U3247 (N_3247,In_1181,In_731);
and U3248 (N_3248,In_1346,In_1140);
nor U3249 (N_3249,In_1041,In_1945);
nand U3250 (N_3250,In_697,In_342);
or U3251 (N_3251,In_115,In_353);
nor U3252 (N_3252,In_1058,In_1094);
or U3253 (N_3253,In_1330,In_1017);
and U3254 (N_3254,In_279,In_1750);
nand U3255 (N_3255,In_223,In_712);
nand U3256 (N_3256,In_1024,In_46);
and U3257 (N_3257,In_250,In_1784);
and U3258 (N_3258,In_872,In_46);
nand U3259 (N_3259,In_235,In_1113);
or U3260 (N_3260,In_1784,In_1877);
and U3261 (N_3261,In_1406,In_377);
nand U3262 (N_3262,In_1491,In_34);
or U3263 (N_3263,In_820,In_576);
and U3264 (N_3264,In_733,In_1485);
nor U3265 (N_3265,In_1357,In_1496);
nor U3266 (N_3266,In_319,In_159);
and U3267 (N_3267,In_1310,In_283);
nand U3268 (N_3268,In_924,In_1727);
or U3269 (N_3269,In_798,In_1406);
nor U3270 (N_3270,In_1325,In_465);
nand U3271 (N_3271,In_474,In_74);
or U3272 (N_3272,In_409,In_925);
nand U3273 (N_3273,In_776,In_257);
and U3274 (N_3274,In_963,In_592);
and U3275 (N_3275,In_486,In_1687);
nand U3276 (N_3276,In_1493,In_1250);
nor U3277 (N_3277,In_862,In_1570);
and U3278 (N_3278,In_1774,In_923);
or U3279 (N_3279,In_1364,In_1357);
and U3280 (N_3280,In_1012,In_1174);
nor U3281 (N_3281,In_1611,In_1536);
nor U3282 (N_3282,In_1901,In_259);
nand U3283 (N_3283,In_596,In_735);
xnor U3284 (N_3284,In_294,In_85);
nand U3285 (N_3285,In_945,In_1529);
and U3286 (N_3286,In_1503,In_1318);
nand U3287 (N_3287,In_559,In_815);
nand U3288 (N_3288,In_732,In_708);
and U3289 (N_3289,In_389,In_922);
and U3290 (N_3290,In_380,In_92);
nand U3291 (N_3291,In_332,In_1528);
and U3292 (N_3292,In_1492,In_83);
nor U3293 (N_3293,In_40,In_1706);
nand U3294 (N_3294,In_140,In_577);
nor U3295 (N_3295,In_1563,In_1995);
and U3296 (N_3296,In_265,In_1432);
nand U3297 (N_3297,In_1013,In_1829);
and U3298 (N_3298,In_1050,In_412);
xnor U3299 (N_3299,In_725,In_1268);
nor U3300 (N_3300,In_298,In_1332);
xnor U3301 (N_3301,In_697,In_1259);
nand U3302 (N_3302,In_1247,In_1403);
xor U3303 (N_3303,In_461,In_460);
or U3304 (N_3304,In_528,In_1873);
nor U3305 (N_3305,In_832,In_595);
xor U3306 (N_3306,In_1446,In_1635);
nand U3307 (N_3307,In_1815,In_1572);
and U3308 (N_3308,In_1699,In_1523);
xor U3309 (N_3309,In_819,In_1922);
nand U3310 (N_3310,In_1101,In_252);
and U3311 (N_3311,In_100,In_258);
and U3312 (N_3312,In_200,In_367);
and U3313 (N_3313,In_581,In_393);
nand U3314 (N_3314,In_1642,In_1413);
and U3315 (N_3315,In_857,In_550);
and U3316 (N_3316,In_1419,In_214);
nor U3317 (N_3317,In_1520,In_689);
and U3318 (N_3318,In_1637,In_855);
and U3319 (N_3319,In_1892,In_500);
xnor U3320 (N_3320,In_62,In_1876);
xor U3321 (N_3321,In_1379,In_774);
nor U3322 (N_3322,In_1169,In_825);
nor U3323 (N_3323,In_294,In_87);
nand U3324 (N_3324,In_253,In_476);
nor U3325 (N_3325,In_1248,In_387);
and U3326 (N_3326,In_1674,In_1394);
and U3327 (N_3327,In_1207,In_1000);
and U3328 (N_3328,In_307,In_567);
nand U3329 (N_3329,In_1248,In_24);
xor U3330 (N_3330,In_938,In_765);
nor U3331 (N_3331,In_952,In_49);
nor U3332 (N_3332,In_1618,In_405);
nand U3333 (N_3333,In_666,In_681);
nor U3334 (N_3334,In_1684,In_1155);
and U3335 (N_3335,In_1626,In_959);
or U3336 (N_3336,In_1522,In_1509);
and U3337 (N_3337,In_738,In_882);
or U3338 (N_3338,In_1518,In_505);
nand U3339 (N_3339,In_293,In_643);
xnor U3340 (N_3340,In_407,In_1038);
nand U3341 (N_3341,In_1744,In_1962);
or U3342 (N_3342,In_1749,In_362);
or U3343 (N_3343,In_1319,In_1850);
and U3344 (N_3344,In_1568,In_1475);
or U3345 (N_3345,In_665,In_1492);
nand U3346 (N_3346,In_41,In_1796);
nor U3347 (N_3347,In_1913,In_388);
or U3348 (N_3348,In_1220,In_1610);
or U3349 (N_3349,In_276,In_1636);
or U3350 (N_3350,In_1417,In_1990);
nand U3351 (N_3351,In_1199,In_608);
nand U3352 (N_3352,In_681,In_802);
nor U3353 (N_3353,In_788,In_824);
xnor U3354 (N_3354,In_285,In_1274);
nand U3355 (N_3355,In_121,In_466);
xor U3356 (N_3356,In_1003,In_1753);
nor U3357 (N_3357,In_206,In_817);
nor U3358 (N_3358,In_306,In_457);
nor U3359 (N_3359,In_1555,In_1513);
xor U3360 (N_3360,In_1672,In_1125);
nand U3361 (N_3361,In_666,In_1780);
or U3362 (N_3362,In_702,In_828);
nand U3363 (N_3363,In_346,In_1262);
xnor U3364 (N_3364,In_1882,In_604);
or U3365 (N_3365,In_1189,In_1385);
nand U3366 (N_3366,In_1361,In_1388);
nand U3367 (N_3367,In_1173,In_1743);
nand U3368 (N_3368,In_299,In_1028);
nor U3369 (N_3369,In_1125,In_729);
and U3370 (N_3370,In_485,In_1802);
nor U3371 (N_3371,In_107,In_880);
nand U3372 (N_3372,In_981,In_827);
and U3373 (N_3373,In_1693,In_1709);
or U3374 (N_3374,In_1712,In_37);
nor U3375 (N_3375,In_1353,In_1034);
nor U3376 (N_3376,In_1240,In_509);
and U3377 (N_3377,In_1471,In_500);
nand U3378 (N_3378,In_657,In_1793);
and U3379 (N_3379,In_1872,In_239);
nor U3380 (N_3380,In_431,In_954);
xor U3381 (N_3381,In_253,In_751);
or U3382 (N_3382,In_1630,In_325);
and U3383 (N_3383,In_14,In_537);
nor U3384 (N_3384,In_1625,In_1510);
or U3385 (N_3385,In_1371,In_1527);
nor U3386 (N_3386,In_670,In_46);
nand U3387 (N_3387,In_1343,In_1281);
or U3388 (N_3388,In_1768,In_934);
nor U3389 (N_3389,In_1203,In_127);
xor U3390 (N_3390,In_647,In_1777);
xnor U3391 (N_3391,In_193,In_1983);
or U3392 (N_3392,In_1268,In_1324);
or U3393 (N_3393,In_138,In_1007);
nor U3394 (N_3394,In_235,In_298);
nand U3395 (N_3395,In_234,In_826);
nand U3396 (N_3396,In_1617,In_117);
and U3397 (N_3397,In_1159,In_1636);
nand U3398 (N_3398,In_1818,In_1205);
nand U3399 (N_3399,In_722,In_1041);
and U3400 (N_3400,In_1870,In_338);
and U3401 (N_3401,In_65,In_1295);
or U3402 (N_3402,In_498,In_12);
xor U3403 (N_3403,In_450,In_634);
nor U3404 (N_3404,In_1807,In_528);
xnor U3405 (N_3405,In_1795,In_691);
and U3406 (N_3406,In_1709,In_1894);
nand U3407 (N_3407,In_26,In_1559);
xor U3408 (N_3408,In_1221,In_1634);
nor U3409 (N_3409,In_1772,In_480);
nand U3410 (N_3410,In_505,In_406);
or U3411 (N_3411,In_693,In_871);
nor U3412 (N_3412,In_1786,In_1174);
and U3413 (N_3413,In_1584,In_698);
or U3414 (N_3414,In_1402,In_1459);
xor U3415 (N_3415,In_559,In_542);
and U3416 (N_3416,In_590,In_1919);
or U3417 (N_3417,In_956,In_289);
nand U3418 (N_3418,In_1638,In_1744);
and U3419 (N_3419,In_1267,In_808);
nor U3420 (N_3420,In_1947,In_1662);
and U3421 (N_3421,In_63,In_1278);
nand U3422 (N_3422,In_1582,In_1748);
and U3423 (N_3423,In_1488,In_465);
and U3424 (N_3424,In_1443,In_41);
nor U3425 (N_3425,In_9,In_715);
nor U3426 (N_3426,In_1720,In_156);
xnor U3427 (N_3427,In_1915,In_181);
nor U3428 (N_3428,In_145,In_1960);
nor U3429 (N_3429,In_410,In_1937);
nand U3430 (N_3430,In_1004,In_1422);
nor U3431 (N_3431,In_1406,In_163);
nor U3432 (N_3432,In_537,In_1779);
or U3433 (N_3433,In_1823,In_1863);
and U3434 (N_3434,In_342,In_279);
nor U3435 (N_3435,In_1367,In_85);
nor U3436 (N_3436,In_1151,In_1653);
or U3437 (N_3437,In_909,In_1748);
xor U3438 (N_3438,In_77,In_1249);
and U3439 (N_3439,In_1834,In_1716);
or U3440 (N_3440,In_911,In_761);
nor U3441 (N_3441,In_1468,In_770);
nand U3442 (N_3442,In_1806,In_437);
nor U3443 (N_3443,In_99,In_1077);
xnor U3444 (N_3444,In_1395,In_1052);
xor U3445 (N_3445,In_1250,In_211);
nand U3446 (N_3446,In_1669,In_533);
nand U3447 (N_3447,In_81,In_906);
or U3448 (N_3448,In_1816,In_1454);
nor U3449 (N_3449,In_1145,In_1939);
nor U3450 (N_3450,In_1330,In_1641);
or U3451 (N_3451,In_293,In_1338);
and U3452 (N_3452,In_1897,In_1945);
and U3453 (N_3453,In_1490,In_448);
nor U3454 (N_3454,In_1849,In_1317);
nor U3455 (N_3455,In_228,In_803);
nor U3456 (N_3456,In_206,In_45);
and U3457 (N_3457,In_807,In_1838);
or U3458 (N_3458,In_941,In_569);
or U3459 (N_3459,In_731,In_97);
xnor U3460 (N_3460,In_1960,In_475);
or U3461 (N_3461,In_301,In_1511);
or U3462 (N_3462,In_749,In_11);
nor U3463 (N_3463,In_121,In_1813);
xor U3464 (N_3464,In_1831,In_1208);
nor U3465 (N_3465,In_1551,In_1025);
nor U3466 (N_3466,In_517,In_1682);
nor U3467 (N_3467,In_1611,In_497);
nand U3468 (N_3468,In_408,In_1611);
xnor U3469 (N_3469,In_889,In_1013);
nor U3470 (N_3470,In_617,In_1068);
and U3471 (N_3471,In_750,In_1308);
or U3472 (N_3472,In_1852,In_1046);
nand U3473 (N_3473,In_1299,In_1952);
and U3474 (N_3474,In_389,In_1058);
nand U3475 (N_3475,In_1157,In_323);
and U3476 (N_3476,In_287,In_1760);
or U3477 (N_3477,In_1170,In_529);
nand U3478 (N_3478,In_1060,In_1985);
or U3479 (N_3479,In_1231,In_1930);
or U3480 (N_3480,In_246,In_723);
or U3481 (N_3481,In_340,In_1211);
nor U3482 (N_3482,In_543,In_1816);
and U3483 (N_3483,In_319,In_635);
and U3484 (N_3484,In_915,In_1843);
nor U3485 (N_3485,In_1830,In_551);
nor U3486 (N_3486,In_38,In_1626);
and U3487 (N_3487,In_1611,In_700);
and U3488 (N_3488,In_793,In_1870);
or U3489 (N_3489,In_734,In_870);
nor U3490 (N_3490,In_1553,In_1299);
xnor U3491 (N_3491,In_1018,In_706);
and U3492 (N_3492,In_1621,In_846);
nor U3493 (N_3493,In_770,In_1526);
or U3494 (N_3494,In_61,In_742);
and U3495 (N_3495,In_662,In_625);
nand U3496 (N_3496,In_401,In_534);
or U3497 (N_3497,In_1040,In_124);
nand U3498 (N_3498,In_1420,In_782);
nor U3499 (N_3499,In_411,In_1581);
nand U3500 (N_3500,In_588,In_1530);
and U3501 (N_3501,In_779,In_371);
nand U3502 (N_3502,In_255,In_307);
and U3503 (N_3503,In_1100,In_1075);
nor U3504 (N_3504,In_0,In_1915);
nand U3505 (N_3505,In_1737,In_1650);
nand U3506 (N_3506,In_965,In_665);
or U3507 (N_3507,In_1185,In_1879);
or U3508 (N_3508,In_1763,In_1510);
or U3509 (N_3509,In_1018,In_1827);
nand U3510 (N_3510,In_1194,In_1266);
and U3511 (N_3511,In_326,In_1087);
xnor U3512 (N_3512,In_1129,In_1738);
and U3513 (N_3513,In_1465,In_1812);
nand U3514 (N_3514,In_948,In_461);
nand U3515 (N_3515,In_89,In_248);
nor U3516 (N_3516,In_1686,In_1691);
and U3517 (N_3517,In_849,In_1121);
and U3518 (N_3518,In_1585,In_1955);
nand U3519 (N_3519,In_1988,In_832);
or U3520 (N_3520,In_1865,In_1825);
nand U3521 (N_3521,In_1362,In_1920);
or U3522 (N_3522,In_1577,In_1826);
nand U3523 (N_3523,In_1479,In_1300);
nand U3524 (N_3524,In_899,In_613);
and U3525 (N_3525,In_500,In_1686);
nor U3526 (N_3526,In_1865,In_1194);
nand U3527 (N_3527,In_716,In_634);
nand U3528 (N_3528,In_1530,In_1971);
nor U3529 (N_3529,In_306,In_308);
xnor U3530 (N_3530,In_988,In_853);
and U3531 (N_3531,In_275,In_1420);
nand U3532 (N_3532,In_67,In_813);
nor U3533 (N_3533,In_188,In_1433);
and U3534 (N_3534,In_1887,In_483);
nor U3535 (N_3535,In_1900,In_495);
nand U3536 (N_3536,In_4,In_243);
nor U3537 (N_3537,In_1911,In_1810);
nand U3538 (N_3538,In_1034,In_1643);
or U3539 (N_3539,In_329,In_1777);
xor U3540 (N_3540,In_694,In_423);
or U3541 (N_3541,In_1389,In_1790);
xor U3542 (N_3542,In_459,In_1226);
nor U3543 (N_3543,In_50,In_1690);
and U3544 (N_3544,In_1571,In_564);
nand U3545 (N_3545,In_1685,In_1673);
or U3546 (N_3546,In_1378,In_276);
nor U3547 (N_3547,In_411,In_1352);
and U3548 (N_3548,In_752,In_1088);
nand U3549 (N_3549,In_188,In_1604);
nor U3550 (N_3550,In_805,In_175);
nand U3551 (N_3551,In_520,In_1583);
nor U3552 (N_3552,In_1400,In_1793);
or U3553 (N_3553,In_1364,In_1688);
nand U3554 (N_3554,In_1174,In_295);
or U3555 (N_3555,In_1413,In_1537);
or U3556 (N_3556,In_140,In_7);
and U3557 (N_3557,In_924,In_1805);
nand U3558 (N_3558,In_1375,In_160);
nand U3559 (N_3559,In_737,In_174);
and U3560 (N_3560,In_1253,In_889);
and U3561 (N_3561,In_1908,In_89);
or U3562 (N_3562,In_624,In_1264);
nand U3563 (N_3563,In_1116,In_384);
nor U3564 (N_3564,In_1117,In_115);
and U3565 (N_3565,In_1311,In_1942);
or U3566 (N_3566,In_1077,In_130);
and U3567 (N_3567,In_1549,In_1453);
and U3568 (N_3568,In_1369,In_71);
and U3569 (N_3569,In_770,In_936);
or U3570 (N_3570,In_222,In_1916);
nand U3571 (N_3571,In_1049,In_227);
and U3572 (N_3572,In_1680,In_946);
and U3573 (N_3573,In_1720,In_1439);
xor U3574 (N_3574,In_1862,In_755);
or U3575 (N_3575,In_1248,In_223);
nor U3576 (N_3576,In_401,In_1003);
xnor U3577 (N_3577,In_1902,In_689);
nand U3578 (N_3578,In_1229,In_586);
or U3579 (N_3579,In_602,In_622);
and U3580 (N_3580,In_1880,In_639);
and U3581 (N_3581,In_1850,In_384);
xor U3582 (N_3582,In_982,In_1272);
nand U3583 (N_3583,In_355,In_1697);
nand U3584 (N_3584,In_1402,In_647);
nor U3585 (N_3585,In_1542,In_926);
xnor U3586 (N_3586,In_938,In_969);
nand U3587 (N_3587,In_1861,In_756);
or U3588 (N_3588,In_323,In_438);
nor U3589 (N_3589,In_667,In_1284);
or U3590 (N_3590,In_284,In_108);
and U3591 (N_3591,In_490,In_1680);
nor U3592 (N_3592,In_1480,In_248);
nor U3593 (N_3593,In_1515,In_1927);
or U3594 (N_3594,In_858,In_1933);
or U3595 (N_3595,In_127,In_1005);
and U3596 (N_3596,In_1169,In_735);
nand U3597 (N_3597,In_393,In_1264);
nor U3598 (N_3598,In_921,In_373);
or U3599 (N_3599,In_774,In_925);
xor U3600 (N_3600,In_204,In_1969);
nand U3601 (N_3601,In_1026,In_502);
xnor U3602 (N_3602,In_429,In_1722);
or U3603 (N_3603,In_1010,In_209);
and U3604 (N_3604,In_1689,In_1774);
nand U3605 (N_3605,In_1031,In_1982);
and U3606 (N_3606,In_266,In_1077);
nand U3607 (N_3607,In_1966,In_1410);
or U3608 (N_3608,In_1288,In_388);
or U3609 (N_3609,In_186,In_903);
or U3610 (N_3610,In_578,In_371);
xor U3611 (N_3611,In_1655,In_313);
and U3612 (N_3612,In_1851,In_1971);
or U3613 (N_3613,In_1876,In_568);
nand U3614 (N_3614,In_729,In_1028);
nor U3615 (N_3615,In_686,In_1403);
xor U3616 (N_3616,In_676,In_115);
nand U3617 (N_3617,In_626,In_136);
nand U3618 (N_3618,In_1356,In_334);
nand U3619 (N_3619,In_574,In_645);
nand U3620 (N_3620,In_698,In_1397);
nand U3621 (N_3621,In_1675,In_1205);
xor U3622 (N_3622,In_1378,In_1067);
nand U3623 (N_3623,In_1536,In_1005);
nor U3624 (N_3624,In_1475,In_554);
nor U3625 (N_3625,In_596,In_1916);
nand U3626 (N_3626,In_1260,In_133);
nor U3627 (N_3627,In_944,In_409);
or U3628 (N_3628,In_86,In_780);
and U3629 (N_3629,In_969,In_926);
xor U3630 (N_3630,In_497,In_1576);
nor U3631 (N_3631,In_1193,In_394);
nor U3632 (N_3632,In_1747,In_1522);
nor U3633 (N_3633,In_321,In_1990);
xor U3634 (N_3634,In_1224,In_1548);
and U3635 (N_3635,In_1853,In_998);
nor U3636 (N_3636,In_1471,In_211);
nor U3637 (N_3637,In_1466,In_295);
nand U3638 (N_3638,In_1095,In_451);
nand U3639 (N_3639,In_593,In_1769);
nand U3640 (N_3640,In_349,In_1729);
nand U3641 (N_3641,In_355,In_1303);
or U3642 (N_3642,In_662,In_1911);
nand U3643 (N_3643,In_693,In_1337);
xnor U3644 (N_3644,In_861,In_1648);
nor U3645 (N_3645,In_874,In_195);
or U3646 (N_3646,In_681,In_1292);
nand U3647 (N_3647,In_1391,In_534);
and U3648 (N_3648,In_1795,In_1885);
xor U3649 (N_3649,In_335,In_1132);
or U3650 (N_3650,In_1560,In_537);
or U3651 (N_3651,In_915,In_903);
and U3652 (N_3652,In_593,In_1343);
or U3653 (N_3653,In_528,In_1787);
and U3654 (N_3654,In_542,In_1534);
and U3655 (N_3655,In_1198,In_632);
and U3656 (N_3656,In_808,In_160);
nand U3657 (N_3657,In_1246,In_159);
or U3658 (N_3658,In_1186,In_1281);
xor U3659 (N_3659,In_1587,In_1698);
xor U3660 (N_3660,In_1968,In_1667);
nand U3661 (N_3661,In_1261,In_1978);
and U3662 (N_3662,In_1426,In_1507);
or U3663 (N_3663,In_448,In_947);
or U3664 (N_3664,In_242,In_226);
or U3665 (N_3665,In_530,In_1235);
nor U3666 (N_3666,In_1294,In_183);
xor U3667 (N_3667,In_640,In_766);
and U3668 (N_3668,In_1510,In_1653);
and U3669 (N_3669,In_766,In_1039);
or U3670 (N_3670,In_1607,In_1659);
xor U3671 (N_3671,In_1298,In_1870);
nand U3672 (N_3672,In_578,In_147);
nor U3673 (N_3673,In_426,In_231);
nor U3674 (N_3674,In_942,In_382);
nand U3675 (N_3675,In_452,In_491);
and U3676 (N_3676,In_1907,In_1579);
or U3677 (N_3677,In_1611,In_1920);
and U3678 (N_3678,In_1172,In_1968);
and U3679 (N_3679,In_1788,In_207);
nand U3680 (N_3680,In_1831,In_1804);
or U3681 (N_3681,In_1605,In_1814);
nand U3682 (N_3682,In_386,In_413);
and U3683 (N_3683,In_566,In_714);
nand U3684 (N_3684,In_1343,In_522);
xnor U3685 (N_3685,In_897,In_1263);
or U3686 (N_3686,In_1083,In_534);
or U3687 (N_3687,In_277,In_1061);
and U3688 (N_3688,In_689,In_1285);
nor U3689 (N_3689,In_1005,In_660);
and U3690 (N_3690,In_1226,In_958);
and U3691 (N_3691,In_655,In_175);
xor U3692 (N_3692,In_1588,In_68);
or U3693 (N_3693,In_1017,In_1498);
nor U3694 (N_3694,In_20,In_1304);
or U3695 (N_3695,In_1587,In_877);
nand U3696 (N_3696,In_174,In_559);
or U3697 (N_3697,In_762,In_552);
nand U3698 (N_3698,In_1446,In_868);
and U3699 (N_3699,In_418,In_1655);
or U3700 (N_3700,In_441,In_992);
and U3701 (N_3701,In_1494,In_15);
or U3702 (N_3702,In_752,In_1100);
xnor U3703 (N_3703,In_1244,In_117);
nand U3704 (N_3704,In_1587,In_956);
and U3705 (N_3705,In_91,In_1336);
and U3706 (N_3706,In_1581,In_267);
xnor U3707 (N_3707,In_1782,In_1858);
nand U3708 (N_3708,In_832,In_1882);
nand U3709 (N_3709,In_1389,In_199);
xnor U3710 (N_3710,In_1983,In_97);
or U3711 (N_3711,In_1095,In_1309);
nor U3712 (N_3712,In_1188,In_1716);
and U3713 (N_3713,In_374,In_1393);
and U3714 (N_3714,In_182,In_764);
nand U3715 (N_3715,In_472,In_255);
and U3716 (N_3716,In_649,In_852);
xnor U3717 (N_3717,In_1468,In_1732);
and U3718 (N_3718,In_810,In_731);
and U3719 (N_3719,In_337,In_122);
nor U3720 (N_3720,In_1861,In_1711);
nor U3721 (N_3721,In_1261,In_299);
or U3722 (N_3722,In_966,In_1211);
xnor U3723 (N_3723,In_42,In_1730);
xnor U3724 (N_3724,In_511,In_521);
nor U3725 (N_3725,In_78,In_1764);
and U3726 (N_3726,In_1476,In_122);
and U3727 (N_3727,In_852,In_95);
nand U3728 (N_3728,In_490,In_356);
nor U3729 (N_3729,In_1606,In_1247);
nand U3730 (N_3730,In_576,In_361);
or U3731 (N_3731,In_998,In_1221);
nand U3732 (N_3732,In_1076,In_49);
or U3733 (N_3733,In_865,In_452);
nor U3734 (N_3734,In_1430,In_443);
or U3735 (N_3735,In_1619,In_144);
nand U3736 (N_3736,In_1751,In_1053);
nor U3737 (N_3737,In_1337,In_878);
xnor U3738 (N_3738,In_1203,In_882);
and U3739 (N_3739,In_1914,In_955);
and U3740 (N_3740,In_641,In_1324);
and U3741 (N_3741,In_1680,In_819);
xnor U3742 (N_3742,In_123,In_1830);
nor U3743 (N_3743,In_107,In_1800);
nand U3744 (N_3744,In_233,In_1283);
and U3745 (N_3745,In_1446,In_1642);
xnor U3746 (N_3746,In_1785,In_136);
nand U3747 (N_3747,In_1780,In_1078);
nand U3748 (N_3748,In_222,In_965);
and U3749 (N_3749,In_44,In_1271);
nand U3750 (N_3750,In_1008,In_288);
nor U3751 (N_3751,In_1892,In_313);
nand U3752 (N_3752,In_1988,In_426);
nor U3753 (N_3753,In_1395,In_260);
and U3754 (N_3754,In_117,In_1010);
nor U3755 (N_3755,In_916,In_1523);
and U3756 (N_3756,In_821,In_740);
nor U3757 (N_3757,In_572,In_252);
and U3758 (N_3758,In_498,In_932);
xor U3759 (N_3759,In_1609,In_1886);
nand U3760 (N_3760,In_1042,In_622);
nor U3761 (N_3761,In_842,In_403);
or U3762 (N_3762,In_244,In_850);
and U3763 (N_3763,In_1981,In_157);
and U3764 (N_3764,In_15,In_117);
nor U3765 (N_3765,In_952,In_1512);
nand U3766 (N_3766,In_363,In_1818);
and U3767 (N_3767,In_1261,In_1384);
xnor U3768 (N_3768,In_1637,In_627);
nor U3769 (N_3769,In_1077,In_366);
and U3770 (N_3770,In_1803,In_1478);
nor U3771 (N_3771,In_176,In_1751);
xnor U3772 (N_3772,In_959,In_156);
and U3773 (N_3773,In_308,In_828);
and U3774 (N_3774,In_223,In_1445);
nand U3775 (N_3775,In_241,In_1161);
or U3776 (N_3776,In_824,In_655);
nand U3777 (N_3777,In_1258,In_632);
xnor U3778 (N_3778,In_1903,In_1478);
and U3779 (N_3779,In_1458,In_1451);
nand U3780 (N_3780,In_1578,In_703);
or U3781 (N_3781,In_1075,In_61);
or U3782 (N_3782,In_1008,In_1203);
nor U3783 (N_3783,In_1043,In_1435);
and U3784 (N_3784,In_1300,In_418);
nor U3785 (N_3785,In_483,In_1450);
and U3786 (N_3786,In_1306,In_1988);
xnor U3787 (N_3787,In_993,In_191);
nor U3788 (N_3788,In_230,In_1959);
nand U3789 (N_3789,In_369,In_1943);
xor U3790 (N_3790,In_865,In_1800);
or U3791 (N_3791,In_923,In_972);
or U3792 (N_3792,In_692,In_567);
and U3793 (N_3793,In_1918,In_1562);
and U3794 (N_3794,In_1356,In_1533);
nor U3795 (N_3795,In_1219,In_792);
nor U3796 (N_3796,In_198,In_1914);
xnor U3797 (N_3797,In_1623,In_423);
or U3798 (N_3798,In_268,In_616);
nand U3799 (N_3799,In_317,In_802);
nand U3800 (N_3800,In_683,In_932);
xor U3801 (N_3801,In_786,In_367);
xor U3802 (N_3802,In_1847,In_800);
or U3803 (N_3803,In_841,In_1930);
or U3804 (N_3804,In_1885,In_1033);
nor U3805 (N_3805,In_1338,In_1444);
xnor U3806 (N_3806,In_1564,In_96);
and U3807 (N_3807,In_554,In_1562);
nor U3808 (N_3808,In_46,In_1567);
nand U3809 (N_3809,In_1916,In_1100);
or U3810 (N_3810,In_817,In_1188);
or U3811 (N_3811,In_304,In_125);
nor U3812 (N_3812,In_1428,In_1561);
and U3813 (N_3813,In_78,In_1485);
or U3814 (N_3814,In_1024,In_754);
and U3815 (N_3815,In_813,In_1437);
and U3816 (N_3816,In_1476,In_1008);
nand U3817 (N_3817,In_1352,In_43);
or U3818 (N_3818,In_419,In_971);
nand U3819 (N_3819,In_1415,In_1364);
nand U3820 (N_3820,In_929,In_1163);
nor U3821 (N_3821,In_1404,In_310);
xor U3822 (N_3822,In_169,In_848);
or U3823 (N_3823,In_997,In_948);
nor U3824 (N_3824,In_148,In_1845);
xor U3825 (N_3825,In_1512,In_1597);
nor U3826 (N_3826,In_1688,In_550);
and U3827 (N_3827,In_1735,In_37);
nand U3828 (N_3828,In_1611,In_908);
nor U3829 (N_3829,In_1474,In_1059);
or U3830 (N_3830,In_194,In_210);
or U3831 (N_3831,In_252,In_1576);
nor U3832 (N_3832,In_1566,In_652);
nand U3833 (N_3833,In_1211,In_1272);
or U3834 (N_3834,In_1190,In_307);
or U3835 (N_3835,In_1031,In_295);
or U3836 (N_3836,In_1692,In_1153);
or U3837 (N_3837,In_1424,In_553);
nor U3838 (N_3838,In_1154,In_1626);
nor U3839 (N_3839,In_1351,In_389);
or U3840 (N_3840,In_1296,In_904);
nand U3841 (N_3841,In_1235,In_28);
nor U3842 (N_3842,In_1685,In_1750);
nand U3843 (N_3843,In_1774,In_435);
or U3844 (N_3844,In_684,In_1336);
nand U3845 (N_3845,In_176,In_1468);
nand U3846 (N_3846,In_145,In_10);
nor U3847 (N_3847,In_960,In_1167);
nand U3848 (N_3848,In_217,In_1153);
nand U3849 (N_3849,In_1509,In_1422);
and U3850 (N_3850,In_1484,In_423);
nand U3851 (N_3851,In_1279,In_412);
nor U3852 (N_3852,In_1602,In_859);
and U3853 (N_3853,In_1156,In_731);
nor U3854 (N_3854,In_1605,In_834);
nor U3855 (N_3855,In_1628,In_1923);
xor U3856 (N_3856,In_1125,In_1674);
and U3857 (N_3857,In_652,In_886);
or U3858 (N_3858,In_908,In_893);
nor U3859 (N_3859,In_1943,In_173);
nor U3860 (N_3860,In_36,In_207);
nand U3861 (N_3861,In_1717,In_1480);
or U3862 (N_3862,In_957,In_1171);
or U3863 (N_3863,In_984,In_985);
nor U3864 (N_3864,In_1436,In_1479);
nand U3865 (N_3865,In_714,In_1091);
or U3866 (N_3866,In_284,In_557);
xnor U3867 (N_3867,In_837,In_1018);
nand U3868 (N_3868,In_1148,In_1548);
nor U3869 (N_3869,In_1846,In_322);
nand U3870 (N_3870,In_521,In_1479);
or U3871 (N_3871,In_620,In_1603);
nand U3872 (N_3872,In_1230,In_1628);
or U3873 (N_3873,In_1736,In_1296);
nand U3874 (N_3874,In_458,In_965);
or U3875 (N_3875,In_1468,In_623);
nand U3876 (N_3876,In_1341,In_1800);
and U3877 (N_3877,In_1036,In_97);
or U3878 (N_3878,In_646,In_1985);
and U3879 (N_3879,In_556,In_1000);
nor U3880 (N_3880,In_909,In_1057);
or U3881 (N_3881,In_1691,In_1094);
nor U3882 (N_3882,In_1346,In_1424);
nor U3883 (N_3883,In_695,In_1330);
xnor U3884 (N_3884,In_1211,In_1464);
nor U3885 (N_3885,In_122,In_1411);
xnor U3886 (N_3886,In_835,In_997);
and U3887 (N_3887,In_1846,In_1888);
and U3888 (N_3888,In_721,In_1925);
xor U3889 (N_3889,In_489,In_799);
nor U3890 (N_3890,In_1758,In_173);
and U3891 (N_3891,In_788,In_403);
and U3892 (N_3892,In_1899,In_1895);
nand U3893 (N_3893,In_1155,In_235);
nor U3894 (N_3894,In_263,In_449);
or U3895 (N_3895,In_1522,In_726);
or U3896 (N_3896,In_303,In_144);
or U3897 (N_3897,In_638,In_625);
nor U3898 (N_3898,In_1899,In_474);
and U3899 (N_3899,In_1658,In_1382);
or U3900 (N_3900,In_1778,In_1453);
nand U3901 (N_3901,In_1614,In_270);
xor U3902 (N_3902,In_870,In_639);
or U3903 (N_3903,In_1696,In_1140);
xor U3904 (N_3904,In_1818,In_397);
nand U3905 (N_3905,In_21,In_684);
nand U3906 (N_3906,In_559,In_1344);
or U3907 (N_3907,In_864,In_1879);
or U3908 (N_3908,In_1890,In_1711);
or U3909 (N_3909,In_1949,In_666);
nor U3910 (N_3910,In_514,In_1242);
nand U3911 (N_3911,In_1904,In_1401);
or U3912 (N_3912,In_1885,In_1993);
nand U3913 (N_3913,In_785,In_810);
xnor U3914 (N_3914,In_1238,In_1973);
or U3915 (N_3915,In_802,In_1284);
and U3916 (N_3916,In_426,In_1335);
and U3917 (N_3917,In_1891,In_1815);
and U3918 (N_3918,In_1050,In_1153);
nor U3919 (N_3919,In_1701,In_1201);
or U3920 (N_3920,In_1578,In_859);
xnor U3921 (N_3921,In_1848,In_1121);
nand U3922 (N_3922,In_1838,In_622);
and U3923 (N_3923,In_664,In_408);
nor U3924 (N_3924,In_1099,In_886);
xor U3925 (N_3925,In_1290,In_1439);
nor U3926 (N_3926,In_967,In_295);
and U3927 (N_3927,In_1614,In_1462);
nand U3928 (N_3928,In_767,In_1387);
xor U3929 (N_3929,In_355,In_1104);
or U3930 (N_3930,In_1709,In_1082);
xnor U3931 (N_3931,In_1096,In_1759);
or U3932 (N_3932,In_1445,In_270);
xor U3933 (N_3933,In_514,In_1504);
nor U3934 (N_3934,In_936,In_1700);
nor U3935 (N_3935,In_298,In_418);
and U3936 (N_3936,In_873,In_1510);
and U3937 (N_3937,In_1756,In_1644);
nand U3938 (N_3938,In_1838,In_1134);
nor U3939 (N_3939,In_692,In_555);
nor U3940 (N_3940,In_1751,In_1042);
and U3941 (N_3941,In_914,In_1745);
nor U3942 (N_3942,In_30,In_1356);
xor U3943 (N_3943,In_813,In_1478);
nor U3944 (N_3944,In_1703,In_830);
xnor U3945 (N_3945,In_1478,In_1574);
and U3946 (N_3946,In_1539,In_1364);
nor U3947 (N_3947,In_167,In_1245);
nand U3948 (N_3948,In_368,In_55);
nand U3949 (N_3949,In_862,In_1538);
nand U3950 (N_3950,In_68,In_1684);
nand U3951 (N_3951,In_17,In_54);
or U3952 (N_3952,In_1220,In_1076);
or U3953 (N_3953,In_397,In_1522);
or U3954 (N_3954,In_626,In_1490);
xnor U3955 (N_3955,In_507,In_1919);
and U3956 (N_3956,In_401,In_99);
or U3957 (N_3957,In_1888,In_1450);
nor U3958 (N_3958,In_1173,In_718);
nor U3959 (N_3959,In_1164,In_1933);
or U3960 (N_3960,In_1569,In_997);
nand U3961 (N_3961,In_1407,In_898);
and U3962 (N_3962,In_1947,In_1916);
or U3963 (N_3963,In_1691,In_1301);
xor U3964 (N_3964,In_307,In_570);
or U3965 (N_3965,In_1385,In_1477);
nor U3966 (N_3966,In_1575,In_1998);
and U3967 (N_3967,In_1093,In_1239);
nand U3968 (N_3968,In_1527,In_98);
xnor U3969 (N_3969,In_1563,In_1885);
nand U3970 (N_3970,In_184,In_1975);
and U3971 (N_3971,In_233,In_1598);
nand U3972 (N_3972,In_515,In_878);
and U3973 (N_3973,In_1505,In_923);
xor U3974 (N_3974,In_1108,In_1046);
nand U3975 (N_3975,In_1065,In_650);
nand U3976 (N_3976,In_231,In_320);
and U3977 (N_3977,In_1962,In_1858);
and U3978 (N_3978,In_230,In_52);
nor U3979 (N_3979,In_904,In_1810);
nor U3980 (N_3980,In_1908,In_1195);
or U3981 (N_3981,In_759,In_1491);
nand U3982 (N_3982,In_558,In_1817);
nor U3983 (N_3983,In_841,In_703);
nand U3984 (N_3984,In_710,In_568);
xnor U3985 (N_3985,In_1765,In_1864);
nand U3986 (N_3986,In_301,In_1989);
and U3987 (N_3987,In_1228,In_815);
or U3988 (N_3988,In_518,In_1190);
or U3989 (N_3989,In_1864,In_697);
xor U3990 (N_3990,In_549,In_914);
xor U3991 (N_3991,In_864,In_1553);
xor U3992 (N_3992,In_734,In_565);
xor U3993 (N_3993,In_282,In_1777);
nor U3994 (N_3994,In_1121,In_742);
or U3995 (N_3995,In_134,In_859);
nor U3996 (N_3996,In_1415,In_1255);
nor U3997 (N_3997,In_302,In_820);
or U3998 (N_3998,In_1690,In_519);
nand U3999 (N_3999,In_1267,In_777);
xor U4000 (N_4000,In_136,In_1338);
nand U4001 (N_4001,In_1212,In_1642);
xnor U4002 (N_4002,In_702,In_1326);
or U4003 (N_4003,In_900,In_898);
and U4004 (N_4004,In_1424,In_705);
or U4005 (N_4005,In_884,In_428);
nand U4006 (N_4006,In_1409,In_1453);
nor U4007 (N_4007,In_1299,In_747);
nor U4008 (N_4008,In_1470,In_171);
nor U4009 (N_4009,In_1809,In_656);
or U4010 (N_4010,In_466,In_1965);
nand U4011 (N_4011,In_104,In_1195);
nand U4012 (N_4012,In_1559,In_1920);
and U4013 (N_4013,In_1313,In_963);
nor U4014 (N_4014,In_1461,In_1412);
nand U4015 (N_4015,In_1258,In_1282);
or U4016 (N_4016,In_1159,In_1998);
or U4017 (N_4017,In_1781,In_1772);
nor U4018 (N_4018,In_1268,In_1126);
nand U4019 (N_4019,In_1705,In_1595);
or U4020 (N_4020,In_1498,In_772);
nor U4021 (N_4021,In_1320,In_907);
nor U4022 (N_4022,In_1294,In_120);
and U4023 (N_4023,In_1477,In_261);
xor U4024 (N_4024,In_1282,In_299);
nand U4025 (N_4025,In_926,In_1686);
and U4026 (N_4026,In_1539,In_557);
or U4027 (N_4027,In_1470,In_1838);
nand U4028 (N_4028,In_56,In_1692);
nand U4029 (N_4029,In_1819,In_1399);
nor U4030 (N_4030,In_265,In_1854);
or U4031 (N_4031,In_737,In_1984);
or U4032 (N_4032,In_807,In_668);
nand U4033 (N_4033,In_1909,In_1449);
xor U4034 (N_4034,In_1038,In_1859);
nand U4035 (N_4035,In_1203,In_883);
or U4036 (N_4036,In_1295,In_783);
or U4037 (N_4037,In_650,In_1288);
and U4038 (N_4038,In_1864,In_662);
or U4039 (N_4039,In_1400,In_328);
and U4040 (N_4040,In_1725,In_1659);
nor U4041 (N_4041,In_468,In_1155);
or U4042 (N_4042,In_523,In_1601);
or U4043 (N_4043,In_1302,In_1192);
and U4044 (N_4044,In_37,In_1948);
or U4045 (N_4045,In_1514,In_1023);
xnor U4046 (N_4046,In_117,In_1874);
and U4047 (N_4047,In_1846,In_1856);
or U4048 (N_4048,In_753,In_713);
or U4049 (N_4049,In_1860,In_465);
nor U4050 (N_4050,In_1144,In_26);
nand U4051 (N_4051,In_372,In_758);
and U4052 (N_4052,In_1615,In_106);
nand U4053 (N_4053,In_1379,In_627);
or U4054 (N_4054,In_93,In_886);
and U4055 (N_4055,In_1704,In_452);
nor U4056 (N_4056,In_272,In_399);
and U4057 (N_4057,In_668,In_1547);
nor U4058 (N_4058,In_62,In_990);
and U4059 (N_4059,In_935,In_1528);
nand U4060 (N_4060,In_1102,In_1387);
or U4061 (N_4061,In_1128,In_1394);
nand U4062 (N_4062,In_893,In_1756);
or U4063 (N_4063,In_1402,In_1670);
xor U4064 (N_4064,In_1653,In_284);
nor U4065 (N_4065,In_198,In_1859);
and U4066 (N_4066,In_1439,In_1658);
xor U4067 (N_4067,In_1446,In_256);
xor U4068 (N_4068,In_921,In_1812);
nor U4069 (N_4069,In_848,In_122);
nand U4070 (N_4070,In_372,In_1551);
nor U4071 (N_4071,In_1233,In_274);
and U4072 (N_4072,In_458,In_1365);
and U4073 (N_4073,In_1757,In_435);
and U4074 (N_4074,In_1305,In_574);
xnor U4075 (N_4075,In_355,In_1942);
and U4076 (N_4076,In_864,In_175);
and U4077 (N_4077,In_1925,In_761);
xor U4078 (N_4078,In_451,In_525);
nand U4079 (N_4079,In_1937,In_706);
and U4080 (N_4080,In_131,In_1601);
nand U4081 (N_4081,In_1951,In_1233);
and U4082 (N_4082,In_28,In_804);
nand U4083 (N_4083,In_269,In_1360);
or U4084 (N_4084,In_795,In_1642);
nor U4085 (N_4085,In_1721,In_45);
or U4086 (N_4086,In_1846,In_1079);
or U4087 (N_4087,In_1957,In_1518);
nand U4088 (N_4088,In_757,In_763);
or U4089 (N_4089,In_10,In_1729);
or U4090 (N_4090,In_1754,In_69);
nor U4091 (N_4091,In_1124,In_1749);
and U4092 (N_4092,In_1782,In_1322);
or U4093 (N_4093,In_314,In_324);
and U4094 (N_4094,In_759,In_1913);
nand U4095 (N_4095,In_890,In_489);
and U4096 (N_4096,In_365,In_357);
nand U4097 (N_4097,In_6,In_1119);
or U4098 (N_4098,In_105,In_686);
and U4099 (N_4099,In_1238,In_157);
or U4100 (N_4100,In_1294,In_536);
nand U4101 (N_4101,In_1240,In_262);
nor U4102 (N_4102,In_195,In_383);
and U4103 (N_4103,In_92,In_565);
or U4104 (N_4104,In_835,In_793);
nor U4105 (N_4105,In_1184,In_808);
nor U4106 (N_4106,In_1349,In_1179);
xor U4107 (N_4107,In_352,In_25);
nand U4108 (N_4108,In_121,In_1749);
xnor U4109 (N_4109,In_576,In_1770);
nand U4110 (N_4110,In_1977,In_198);
or U4111 (N_4111,In_1461,In_824);
and U4112 (N_4112,In_808,In_177);
or U4113 (N_4113,In_392,In_1187);
xor U4114 (N_4114,In_62,In_1296);
nor U4115 (N_4115,In_1514,In_720);
and U4116 (N_4116,In_597,In_1076);
and U4117 (N_4117,In_899,In_1929);
or U4118 (N_4118,In_1973,In_178);
nor U4119 (N_4119,In_910,In_452);
nand U4120 (N_4120,In_497,In_923);
and U4121 (N_4121,In_685,In_246);
and U4122 (N_4122,In_654,In_1917);
or U4123 (N_4123,In_1007,In_249);
and U4124 (N_4124,In_1940,In_796);
xor U4125 (N_4125,In_1701,In_597);
and U4126 (N_4126,In_415,In_1716);
or U4127 (N_4127,In_434,In_438);
or U4128 (N_4128,In_1876,In_1733);
or U4129 (N_4129,In_795,In_921);
xor U4130 (N_4130,In_1674,In_1051);
or U4131 (N_4131,In_1180,In_436);
nor U4132 (N_4132,In_1198,In_1011);
xor U4133 (N_4133,In_1803,In_1119);
nand U4134 (N_4134,In_51,In_1202);
or U4135 (N_4135,In_1017,In_1661);
nor U4136 (N_4136,In_1703,In_1178);
or U4137 (N_4137,In_158,In_506);
xnor U4138 (N_4138,In_246,In_245);
nand U4139 (N_4139,In_1609,In_1115);
or U4140 (N_4140,In_614,In_64);
nor U4141 (N_4141,In_17,In_680);
and U4142 (N_4142,In_778,In_1234);
nand U4143 (N_4143,In_1753,In_1878);
and U4144 (N_4144,In_1647,In_1625);
nand U4145 (N_4145,In_1695,In_116);
and U4146 (N_4146,In_712,In_1954);
and U4147 (N_4147,In_906,In_1843);
xor U4148 (N_4148,In_1769,In_1042);
nor U4149 (N_4149,In_1293,In_1079);
or U4150 (N_4150,In_452,In_818);
or U4151 (N_4151,In_1628,In_983);
and U4152 (N_4152,In_77,In_101);
or U4153 (N_4153,In_1612,In_1883);
and U4154 (N_4154,In_1981,In_628);
xnor U4155 (N_4155,In_505,In_1371);
and U4156 (N_4156,In_1168,In_1155);
nor U4157 (N_4157,In_1690,In_1033);
or U4158 (N_4158,In_798,In_1351);
or U4159 (N_4159,In_1829,In_143);
or U4160 (N_4160,In_1470,In_1870);
nand U4161 (N_4161,In_1774,In_1246);
nand U4162 (N_4162,In_71,In_1005);
and U4163 (N_4163,In_73,In_848);
or U4164 (N_4164,In_192,In_1778);
or U4165 (N_4165,In_732,In_256);
and U4166 (N_4166,In_1225,In_1169);
or U4167 (N_4167,In_872,In_1606);
or U4168 (N_4168,In_121,In_1568);
xnor U4169 (N_4169,In_462,In_958);
nand U4170 (N_4170,In_1888,In_1605);
and U4171 (N_4171,In_1100,In_1675);
nor U4172 (N_4172,In_1910,In_275);
nand U4173 (N_4173,In_875,In_1221);
nand U4174 (N_4174,In_754,In_1553);
or U4175 (N_4175,In_1670,In_107);
and U4176 (N_4176,In_1378,In_263);
xor U4177 (N_4177,In_439,In_774);
xor U4178 (N_4178,In_50,In_731);
nand U4179 (N_4179,In_433,In_1744);
nand U4180 (N_4180,In_377,In_1844);
and U4181 (N_4181,In_723,In_978);
or U4182 (N_4182,In_339,In_469);
and U4183 (N_4183,In_1134,In_1379);
and U4184 (N_4184,In_691,In_674);
nand U4185 (N_4185,In_1117,In_176);
or U4186 (N_4186,In_1221,In_760);
or U4187 (N_4187,In_452,In_840);
nand U4188 (N_4188,In_230,In_805);
xor U4189 (N_4189,In_241,In_1745);
and U4190 (N_4190,In_948,In_1993);
nor U4191 (N_4191,In_370,In_990);
nor U4192 (N_4192,In_1488,In_1108);
or U4193 (N_4193,In_1188,In_717);
or U4194 (N_4194,In_1947,In_227);
xor U4195 (N_4195,In_1022,In_1024);
or U4196 (N_4196,In_569,In_1793);
nor U4197 (N_4197,In_1777,In_449);
or U4198 (N_4198,In_7,In_1543);
nand U4199 (N_4199,In_833,In_888);
nor U4200 (N_4200,In_898,In_354);
nor U4201 (N_4201,In_489,In_983);
and U4202 (N_4202,In_380,In_1384);
nor U4203 (N_4203,In_404,In_1648);
nand U4204 (N_4204,In_67,In_150);
and U4205 (N_4205,In_873,In_869);
xor U4206 (N_4206,In_499,In_1473);
and U4207 (N_4207,In_1522,In_988);
nor U4208 (N_4208,In_563,In_1136);
and U4209 (N_4209,In_119,In_1779);
nor U4210 (N_4210,In_1511,In_1698);
or U4211 (N_4211,In_851,In_764);
and U4212 (N_4212,In_1745,In_895);
nor U4213 (N_4213,In_1947,In_572);
xor U4214 (N_4214,In_35,In_1091);
or U4215 (N_4215,In_119,In_286);
and U4216 (N_4216,In_238,In_533);
xor U4217 (N_4217,In_590,In_1525);
nor U4218 (N_4218,In_309,In_854);
nor U4219 (N_4219,In_1929,In_1683);
or U4220 (N_4220,In_1898,In_647);
nor U4221 (N_4221,In_1493,In_1830);
or U4222 (N_4222,In_888,In_1465);
or U4223 (N_4223,In_1208,In_1203);
and U4224 (N_4224,In_692,In_263);
and U4225 (N_4225,In_1344,In_688);
or U4226 (N_4226,In_1025,In_1717);
nor U4227 (N_4227,In_326,In_1738);
nand U4228 (N_4228,In_1500,In_1747);
nand U4229 (N_4229,In_629,In_1856);
and U4230 (N_4230,In_985,In_957);
or U4231 (N_4231,In_974,In_1583);
nand U4232 (N_4232,In_1144,In_1448);
nand U4233 (N_4233,In_1919,In_1237);
nor U4234 (N_4234,In_172,In_220);
nand U4235 (N_4235,In_77,In_988);
and U4236 (N_4236,In_1974,In_1268);
nor U4237 (N_4237,In_1503,In_632);
xnor U4238 (N_4238,In_537,In_1657);
or U4239 (N_4239,In_1614,In_830);
or U4240 (N_4240,In_1754,In_1305);
nand U4241 (N_4241,In_228,In_1490);
or U4242 (N_4242,In_1845,In_1952);
or U4243 (N_4243,In_767,In_89);
nor U4244 (N_4244,In_1491,In_912);
or U4245 (N_4245,In_889,In_811);
xnor U4246 (N_4246,In_247,In_245);
nand U4247 (N_4247,In_1628,In_1853);
nand U4248 (N_4248,In_640,In_688);
xnor U4249 (N_4249,In_710,In_692);
nand U4250 (N_4250,In_1617,In_1689);
nand U4251 (N_4251,In_410,In_1305);
nor U4252 (N_4252,In_1420,In_1150);
and U4253 (N_4253,In_46,In_1690);
nand U4254 (N_4254,In_1674,In_843);
nor U4255 (N_4255,In_1434,In_1784);
nor U4256 (N_4256,In_1901,In_719);
and U4257 (N_4257,In_1536,In_1264);
and U4258 (N_4258,In_709,In_1851);
nor U4259 (N_4259,In_481,In_461);
and U4260 (N_4260,In_83,In_1066);
and U4261 (N_4261,In_1782,In_1420);
nor U4262 (N_4262,In_319,In_731);
nor U4263 (N_4263,In_716,In_1310);
or U4264 (N_4264,In_1144,In_816);
or U4265 (N_4265,In_701,In_1082);
and U4266 (N_4266,In_667,In_1567);
xnor U4267 (N_4267,In_462,In_1422);
nor U4268 (N_4268,In_515,In_1310);
nand U4269 (N_4269,In_755,In_1441);
and U4270 (N_4270,In_306,In_1092);
and U4271 (N_4271,In_942,In_1268);
nor U4272 (N_4272,In_1232,In_1906);
xnor U4273 (N_4273,In_1225,In_944);
nand U4274 (N_4274,In_879,In_224);
nand U4275 (N_4275,In_1821,In_1993);
or U4276 (N_4276,In_1395,In_1322);
xor U4277 (N_4277,In_197,In_804);
nand U4278 (N_4278,In_501,In_1963);
nor U4279 (N_4279,In_1216,In_961);
nor U4280 (N_4280,In_870,In_1622);
nand U4281 (N_4281,In_785,In_512);
nor U4282 (N_4282,In_1607,In_630);
or U4283 (N_4283,In_230,In_1583);
and U4284 (N_4284,In_691,In_1827);
nand U4285 (N_4285,In_1171,In_722);
nor U4286 (N_4286,In_958,In_1669);
nor U4287 (N_4287,In_1392,In_1020);
nand U4288 (N_4288,In_1689,In_1076);
nor U4289 (N_4289,In_1191,In_501);
xor U4290 (N_4290,In_194,In_1131);
nand U4291 (N_4291,In_838,In_1324);
nand U4292 (N_4292,In_1920,In_230);
nor U4293 (N_4293,In_110,In_383);
nor U4294 (N_4294,In_102,In_964);
nor U4295 (N_4295,In_764,In_215);
or U4296 (N_4296,In_86,In_1552);
or U4297 (N_4297,In_1848,In_200);
and U4298 (N_4298,In_544,In_276);
nor U4299 (N_4299,In_797,In_12);
and U4300 (N_4300,In_181,In_876);
nand U4301 (N_4301,In_701,In_1223);
or U4302 (N_4302,In_1562,In_1701);
xnor U4303 (N_4303,In_532,In_970);
or U4304 (N_4304,In_268,In_1926);
nand U4305 (N_4305,In_1584,In_1604);
or U4306 (N_4306,In_1402,In_1810);
nor U4307 (N_4307,In_950,In_1358);
or U4308 (N_4308,In_595,In_166);
nor U4309 (N_4309,In_1020,In_744);
and U4310 (N_4310,In_1289,In_1138);
and U4311 (N_4311,In_218,In_1526);
and U4312 (N_4312,In_706,In_1582);
nand U4313 (N_4313,In_415,In_568);
or U4314 (N_4314,In_1168,In_462);
and U4315 (N_4315,In_411,In_272);
or U4316 (N_4316,In_1449,In_661);
xor U4317 (N_4317,In_1959,In_1479);
xor U4318 (N_4318,In_1908,In_300);
nand U4319 (N_4319,In_775,In_1855);
or U4320 (N_4320,In_183,In_989);
and U4321 (N_4321,In_1718,In_1119);
and U4322 (N_4322,In_1636,In_718);
nand U4323 (N_4323,In_157,In_1906);
nand U4324 (N_4324,In_1317,In_1778);
nand U4325 (N_4325,In_215,In_1502);
or U4326 (N_4326,In_908,In_1334);
nand U4327 (N_4327,In_670,In_995);
and U4328 (N_4328,In_1506,In_230);
or U4329 (N_4329,In_797,In_1090);
nand U4330 (N_4330,In_1685,In_707);
or U4331 (N_4331,In_506,In_1286);
nor U4332 (N_4332,In_1111,In_677);
and U4333 (N_4333,In_1804,In_212);
nand U4334 (N_4334,In_1872,In_1089);
nor U4335 (N_4335,In_1104,In_179);
nor U4336 (N_4336,In_1847,In_1590);
or U4337 (N_4337,In_1252,In_1597);
xnor U4338 (N_4338,In_210,In_599);
xnor U4339 (N_4339,In_1614,In_1323);
and U4340 (N_4340,In_1311,In_1824);
or U4341 (N_4341,In_1499,In_377);
or U4342 (N_4342,In_602,In_742);
or U4343 (N_4343,In_1283,In_692);
xnor U4344 (N_4344,In_55,In_1608);
nand U4345 (N_4345,In_236,In_420);
nor U4346 (N_4346,In_1708,In_1995);
nand U4347 (N_4347,In_988,In_1329);
nor U4348 (N_4348,In_1787,In_658);
and U4349 (N_4349,In_435,In_1914);
nand U4350 (N_4350,In_1151,In_650);
nand U4351 (N_4351,In_1937,In_332);
xnor U4352 (N_4352,In_1365,In_1086);
xnor U4353 (N_4353,In_964,In_1239);
or U4354 (N_4354,In_808,In_878);
nand U4355 (N_4355,In_1091,In_1303);
or U4356 (N_4356,In_633,In_1066);
nor U4357 (N_4357,In_293,In_1666);
nand U4358 (N_4358,In_555,In_1937);
nand U4359 (N_4359,In_1483,In_163);
and U4360 (N_4360,In_1993,In_399);
nand U4361 (N_4361,In_984,In_33);
xor U4362 (N_4362,In_1715,In_820);
or U4363 (N_4363,In_1739,In_1089);
nor U4364 (N_4364,In_783,In_338);
nand U4365 (N_4365,In_1890,In_967);
or U4366 (N_4366,In_1437,In_1848);
nand U4367 (N_4367,In_866,In_1645);
and U4368 (N_4368,In_1758,In_1698);
or U4369 (N_4369,In_1042,In_913);
and U4370 (N_4370,In_686,In_1521);
or U4371 (N_4371,In_1627,In_579);
or U4372 (N_4372,In_1831,In_42);
or U4373 (N_4373,In_978,In_1536);
or U4374 (N_4374,In_374,In_1217);
nand U4375 (N_4375,In_1510,In_1596);
or U4376 (N_4376,In_1480,In_900);
nor U4377 (N_4377,In_1066,In_453);
and U4378 (N_4378,In_403,In_1642);
and U4379 (N_4379,In_1163,In_722);
or U4380 (N_4380,In_1190,In_1868);
nand U4381 (N_4381,In_75,In_1432);
nor U4382 (N_4382,In_786,In_1582);
and U4383 (N_4383,In_938,In_327);
and U4384 (N_4384,In_680,In_385);
and U4385 (N_4385,In_1327,In_665);
or U4386 (N_4386,In_6,In_1063);
and U4387 (N_4387,In_1239,In_175);
or U4388 (N_4388,In_304,In_1544);
nand U4389 (N_4389,In_770,In_480);
xor U4390 (N_4390,In_1610,In_1583);
and U4391 (N_4391,In_1745,In_879);
nand U4392 (N_4392,In_1367,In_57);
or U4393 (N_4393,In_1443,In_1841);
and U4394 (N_4394,In_181,In_1213);
nand U4395 (N_4395,In_147,In_309);
and U4396 (N_4396,In_1441,In_1075);
xnor U4397 (N_4397,In_668,In_573);
nand U4398 (N_4398,In_0,In_1132);
xnor U4399 (N_4399,In_714,In_1713);
nor U4400 (N_4400,In_1319,In_251);
or U4401 (N_4401,In_417,In_730);
nor U4402 (N_4402,In_173,In_821);
and U4403 (N_4403,In_1637,In_1397);
nor U4404 (N_4404,In_1299,In_705);
nand U4405 (N_4405,In_915,In_1674);
xnor U4406 (N_4406,In_1875,In_1498);
and U4407 (N_4407,In_1186,In_1359);
nor U4408 (N_4408,In_710,In_85);
nor U4409 (N_4409,In_996,In_1511);
or U4410 (N_4410,In_474,In_1500);
nand U4411 (N_4411,In_143,In_829);
or U4412 (N_4412,In_174,In_1690);
nor U4413 (N_4413,In_1865,In_1309);
or U4414 (N_4414,In_237,In_913);
or U4415 (N_4415,In_667,In_1955);
and U4416 (N_4416,In_881,In_1813);
or U4417 (N_4417,In_1901,In_959);
nand U4418 (N_4418,In_489,In_1256);
and U4419 (N_4419,In_1552,In_211);
or U4420 (N_4420,In_1480,In_373);
nand U4421 (N_4421,In_986,In_829);
nand U4422 (N_4422,In_587,In_310);
nand U4423 (N_4423,In_326,In_1483);
nor U4424 (N_4424,In_1218,In_180);
nand U4425 (N_4425,In_1863,In_1602);
or U4426 (N_4426,In_861,In_1503);
nor U4427 (N_4427,In_1560,In_1399);
nand U4428 (N_4428,In_1586,In_1946);
or U4429 (N_4429,In_1927,In_699);
nor U4430 (N_4430,In_804,In_1409);
nor U4431 (N_4431,In_1263,In_193);
and U4432 (N_4432,In_1570,In_1256);
and U4433 (N_4433,In_1220,In_681);
or U4434 (N_4434,In_988,In_1431);
or U4435 (N_4435,In_95,In_1877);
xnor U4436 (N_4436,In_625,In_1572);
nor U4437 (N_4437,In_1547,In_1271);
nand U4438 (N_4438,In_804,In_1000);
nor U4439 (N_4439,In_1171,In_986);
nand U4440 (N_4440,In_1762,In_1275);
nand U4441 (N_4441,In_1368,In_58);
and U4442 (N_4442,In_1725,In_898);
or U4443 (N_4443,In_1771,In_853);
or U4444 (N_4444,In_1672,In_957);
and U4445 (N_4445,In_1913,In_1532);
nor U4446 (N_4446,In_1189,In_616);
nor U4447 (N_4447,In_558,In_1156);
xnor U4448 (N_4448,In_145,In_1055);
nand U4449 (N_4449,In_1056,In_1131);
and U4450 (N_4450,In_1924,In_1154);
nand U4451 (N_4451,In_781,In_1796);
nor U4452 (N_4452,In_390,In_1187);
or U4453 (N_4453,In_835,In_1903);
and U4454 (N_4454,In_1448,In_935);
and U4455 (N_4455,In_1138,In_1207);
and U4456 (N_4456,In_1020,In_995);
or U4457 (N_4457,In_1896,In_1877);
or U4458 (N_4458,In_1253,In_1199);
or U4459 (N_4459,In_1791,In_1471);
and U4460 (N_4460,In_483,In_1863);
or U4461 (N_4461,In_968,In_966);
or U4462 (N_4462,In_1015,In_1451);
nor U4463 (N_4463,In_449,In_594);
nor U4464 (N_4464,In_938,In_390);
and U4465 (N_4465,In_1291,In_725);
nand U4466 (N_4466,In_308,In_660);
or U4467 (N_4467,In_1158,In_1379);
nand U4468 (N_4468,In_975,In_1848);
xor U4469 (N_4469,In_37,In_1460);
nand U4470 (N_4470,In_451,In_1594);
or U4471 (N_4471,In_28,In_847);
nor U4472 (N_4472,In_892,In_926);
nand U4473 (N_4473,In_945,In_874);
or U4474 (N_4474,In_1597,In_134);
or U4475 (N_4475,In_665,In_93);
nor U4476 (N_4476,In_808,In_1480);
xor U4477 (N_4477,In_11,In_210);
or U4478 (N_4478,In_344,In_105);
and U4479 (N_4479,In_1447,In_830);
or U4480 (N_4480,In_1237,In_1957);
nor U4481 (N_4481,In_247,In_1020);
or U4482 (N_4482,In_1294,In_407);
nand U4483 (N_4483,In_1641,In_1427);
or U4484 (N_4484,In_1230,In_405);
xor U4485 (N_4485,In_1885,In_248);
nand U4486 (N_4486,In_1096,In_1938);
or U4487 (N_4487,In_1662,In_924);
and U4488 (N_4488,In_1076,In_1602);
and U4489 (N_4489,In_1851,In_1665);
nand U4490 (N_4490,In_769,In_802);
and U4491 (N_4491,In_957,In_463);
or U4492 (N_4492,In_1013,In_1382);
nand U4493 (N_4493,In_881,In_1075);
and U4494 (N_4494,In_1820,In_1674);
nand U4495 (N_4495,In_444,In_1848);
and U4496 (N_4496,In_1716,In_553);
nand U4497 (N_4497,In_802,In_996);
or U4498 (N_4498,In_1809,In_1636);
nand U4499 (N_4499,In_90,In_1661);
nand U4500 (N_4500,In_1597,In_1884);
nor U4501 (N_4501,In_550,In_558);
or U4502 (N_4502,In_346,In_398);
and U4503 (N_4503,In_187,In_883);
and U4504 (N_4504,In_1,In_372);
nor U4505 (N_4505,In_326,In_1859);
nand U4506 (N_4506,In_102,In_929);
and U4507 (N_4507,In_1387,In_27);
nor U4508 (N_4508,In_1784,In_896);
xnor U4509 (N_4509,In_1112,In_1331);
nand U4510 (N_4510,In_133,In_1206);
nor U4511 (N_4511,In_742,In_777);
or U4512 (N_4512,In_1097,In_954);
nand U4513 (N_4513,In_455,In_1049);
nand U4514 (N_4514,In_1632,In_41);
xor U4515 (N_4515,In_244,In_551);
or U4516 (N_4516,In_1956,In_1664);
nor U4517 (N_4517,In_1019,In_713);
and U4518 (N_4518,In_1443,In_458);
nand U4519 (N_4519,In_1993,In_318);
and U4520 (N_4520,In_1384,In_57);
nor U4521 (N_4521,In_1736,In_1002);
and U4522 (N_4522,In_1831,In_1919);
nand U4523 (N_4523,In_1132,In_772);
xor U4524 (N_4524,In_1940,In_718);
or U4525 (N_4525,In_109,In_774);
nand U4526 (N_4526,In_24,In_1782);
nand U4527 (N_4527,In_19,In_51);
or U4528 (N_4528,In_1717,In_1908);
or U4529 (N_4529,In_1799,In_1494);
nand U4530 (N_4530,In_529,In_1801);
or U4531 (N_4531,In_486,In_215);
nor U4532 (N_4532,In_572,In_971);
and U4533 (N_4533,In_469,In_440);
nor U4534 (N_4534,In_232,In_75);
or U4535 (N_4535,In_1285,In_443);
or U4536 (N_4536,In_325,In_1317);
or U4537 (N_4537,In_635,In_1332);
and U4538 (N_4538,In_881,In_633);
nand U4539 (N_4539,In_333,In_434);
nand U4540 (N_4540,In_1756,In_1424);
and U4541 (N_4541,In_1346,In_659);
and U4542 (N_4542,In_720,In_1063);
nor U4543 (N_4543,In_964,In_230);
and U4544 (N_4544,In_472,In_1272);
nand U4545 (N_4545,In_1714,In_454);
nor U4546 (N_4546,In_1057,In_1727);
nor U4547 (N_4547,In_895,In_686);
and U4548 (N_4548,In_1097,In_1631);
nand U4549 (N_4549,In_1810,In_1264);
or U4550 (N_4550,In_1777,In_488);
and U4551 (N_4551,In_628,In_909);
nor U4552 (N_4552,In_1237,In_1713);
nor U4553 (N_4553,In_296,In_260);
and U4554 (N_4554,In_1878,In_1565);
xor U4555 (N_4555,In_886,In_1259);
xnor U4556 (N_4556,In_1180,In_978);
nand U4557 (N_4557,In_1737,In_581);
nand U4558 (N_4558,In_827,In_1047);
and U4559 (N_4559,In_1592,In_388);
and U4560 (N_4560,In_489,In_832);
or U4561 (N_4561,In_516,In_1071);
nand U4562 (N_4562,In_1968,In_577);
nor U4563 (N_4563,In_1646,In_1530);
nand U4564 (N_4564,In_1204,In_963);
nor U4565 (N_4565,In_1359,In_1586);
and U4566 (N_4566,In_1621,In_1705);
or U4567 (N_4567,In_781,In_1154);
nand U4568 (N_4568,In_1706,In_89);
nand U4569 (N_4569,In_768,In_1958);
nand U4570 (N_4570,In_1304,In_690);
or U4571 (N_4571,In_990,In_115);
or U4572 (N_4572,In_1698,In_1512);
nand U4573 (N_4573,In_1699,In_1573);
or U4574 (N_4574,In_1709,In_121);
nor U4575 (N_4575,In_1887,In_426);
and U4576 (N_4576,In_163,In_64);
nor U4577 (N_4577,In_370,In_1916);
nor U4578 (N_4578,In_1826,In_1418);
or U4579 (N_4579,In_123,In_265);
nand U4580 (N_4580,In_1701,In_638);
and U4581 (N_4581,In_1572,In_479);
xor U4582 (N_4582,In_120,In_849);
or U4583 (N_4583,In_1193,In_1201);
nand U4584 (N_4584,In_1778,In_921);
nand U4585 (N_4585,In_388,In_540);
or U4586 (N_4586,In_531,In_493);
and U4587 (N_4587,In_462,In_182);
and U4588 (N_4588,In_1571,In_690);
and U4589 (N_4589,In_1125,In_1313);
nand U4590 (N_4590,In_1538,In_457);
nand U4591 (N_4591,In_1945,In_859);
nor U4592 (N_4592,In_1588,In_1264);
xor U4593 (N_4593,In_1286,In_1841);
and U4594 (N_4594,In_1985,In_1642);
or U4595 (N_4595,In_450,In_1917);
and U4596 (N_4596,In_711,In_1087);
nor U4597 (N_4597,In_142,In_1214);
nand U4598 (N_4598,In_875,In_1773);
nor U4599 (N_4599,In_1329,In_1765);
nor U4600 (N_4600,In_961,In_308);
nor U4601 (N_4601,In_118,In_1954);
xnor U4602 (N_4602,In_561,In_916);
xor U4603 (N_4603,In_1007,In_564);
and U4604 (N_4604,In_1838,In_1904);
nand U4605 (N_4605,In_1137,In_1457);
nand U4606 (N_4606,In_855,In_876);
xnor U4607 (N_4607,In_1493,In_814);
nor U4608 (N_4608,In_247,In_20);
nor U4609 (N_4609,In_1157,In_858);
and U4610 (N_4610,In_1350,In_753);
and U4611 (N_4611,In_410,In_614);
or U4612 (N_4612,In_471,In_222);
and U4613 (N_4613,In_1058,In_1315);
or U4614 (N_4614,In_1261,In_1435);
or U4615 (N_4615,In_423,In_1620);
nor U4616 (N_4616,In_383,In_545);
nand U4617 (N_4617,In_538,In_1685);
nand U4618 (N_4618,In_207,In_690);
and U4619 (N_4619,In_255,In_158);
nand U4620 (N_4620,In_1740,In_1566);
and U4621 (N_4621,In_75,In_436);
or U4622 (N_4622,In_1262,In_101);
and U4623 (N_4623,In_74,In_562);
or U4624 (N_4624,In_791,In_1548);
or U4625 (N_4625,In_1082,In_1260);
nor U4626 (N_4626,In_942,In_1842);
or U4627 (N_4627,In_1594,In_1222);
and U4628 (N_4628,In_228,In_493);
xor U4629 (N_4629,In_1964,In_1168);
nor U4630 (N_4630,In_1167,In_805);
nor U4631 (N_4631,In_1422,In_1061);
nand U4632 (N_4632,In_407,In_1003);
or U4633 (N_4633,In_316,In_296);
or U4634 (N_4634,In_803,In_588);
nor U4635 (N_4635,In_820,In_459);
nor U4636 (N_4636,In_195,In_1225);
xnor U4637 (N_4637,In_1430,In_1597);
and U4638 (N_4638,In_1981,In_1054);
or U4639 (N_4639,In_1445,In_1);
nand U4640 (N_4640,In_1132,In_1096);
nand U4641 (N_4641,In_970,In_139);
nand U4642 (N_4642,In_1789,In_1050);
and U4643 (N_4643,In_1921,In_97);
or U4644 (N_4644,In_1771,In_1571);
xor U4645 (N_4645,In_699,In_352);
and U4646 (N_4646,In_189,In_567);
nand U4647 (N_4647,In_648,In_1052);
and U4648 (N_4648,In_513,In_129);
or U4649 (N_4649,In_727,In_359);
or U4650 (N_4650,In_1232,In_1704);
or U4651 (N_4651,In_1809,In_975);
nor U4652 (N_4652,In_1646,In_12);
nand U4653 (N_4653,In_998,In_1935);
and U4654 (N_4654,In_1560,In_1673);
and U4655 (N_4655,In_33,In_389);
nor U4656 (N_4656,In_378,In_930);
and U4657 (N_4657,In_1592,In_840);
nor U4658 (N_4658,In_1187,In_45);
nand U4659 (N_4659,In_1572,In_821);
nand U4660 (N_4660,In_1416,In_1648);
or U4661 (N_4661,In_1378,In_1164);
nor U4662 (N_4662,In_827,In_946);
xnor U4663 (N_4663,In_1956,In_253);
or U4664 (N_4664,In_1203,In_1761);
and U4665 (N_4665,In_679,In_1769);
and U4666 (N_4666,In_449,In_1177);
nand U4667 (N_4667,In_722,In_888);
nand U4668 (N_4668,In_1864,In_1487);
nand U4669 (N_4669,In_1017,In_889);
xnor U4670 (N_4670,In_1377,In_1649);
or U4671 (N_4671,In_1306,In_551);
and U4672 (N_4672,In_1649,In_1857);
nor U4673 (N_4673,In_974,In_1007);
nor U4674 (N_4674,In_1228,In_1639);
nor U4675 (N_4675,In_862,In_542);
and U4676 (N_4676,In_1662,In_1852);
or U4677 (N_4677,In_1229,In_762);
nand U4678 (N_4678,In_912,In_725);
nand U4679 (N_4679,In_732,In_309);
xor U4680 (N_4680,In_1387,In_178);
and U4681 (N_4681,In_833,In_1725);
and U4682 (N_4682,In_776,In_1948);
nor U4683 (N_4683,In_123,In_1681);
nor U4684 (N_4684,In_193,In_470);
or U4685 (N_4685,In_1433,In_870);
or U4686 (N_4686,In_1397,In_604);
or U4687 (N_4687,In_739,In_588);
and U4688 (N_4688,In_1517,In_1997);
nand U4689 (N_4689,In_262,In_100);
nand U4690 (N_4690,In_1730,In_490);
nor U4691 (N_4691,In_943,In_1141);
and U4692 (N_4692,In_660,In_174);
nand U4693 (N_4693,In_1932,In_1706);
nor U4694 (N_4694,In_597,In_632);
nand U4695 (N_4695,In_1105,In_1597);
or U4696 (N_4696,In_1155,In_1244);
nor U4697 (N_4697,In_1632,In_250);
nor U4698 (N_4698,In_429,In_1484);
nand U4699 (N_4699,In_1361,In_900);
xor U4700 (N_4700,In_428,In_21);
nand U4701 (N_4701,In_1989,In_328);
nor U4702 (N_4702,In_126,In_133);
nor U4703 (N_4703,In_1168,In_503);
or U4704 (N_4704,In_766,In_686);
or U4705 (N_4705,In_1717,In_1860);
and U4706 (N_4706,In_1732,In_1801);
and U4707 (N_4707,In_1971,In_1208);
or U4708 (N_4708,In_1648,In_1112);
or U4709 (N_4709,In_1330,In_939);
nand U4710 (N_4710,In_1378,In_1434);
nand U4711 (N_4711,In_1537,In_794);
and U4712 (N_4712,In_868,In_1657);
or U4713 (N_4713,In_1962,In_304);
and U4714 (N_4714,In_803,In_510);
or U4715 (N_4715,In_952,In_1132);
nor U4716 (N_4716,In_954,In_974);
nor U4717 (N_4717,In_1975,In_1978);
nor U4718 (N_4718,In_1537,In_563);
nand U4719 (N_4719,In_534,In_1216);
and U4720 (N_4720,In_273,In_185);
nor U4721 (N_4721,In_1235,In_1921);
or U4722 (N_4722,In_340,In_1669);
or U4723 (N_4723,In_1595,In_833);
nand U4724 (N_4724,In_317,In_1828);
nand U4725 (N_4725,In_1821,In_191);
or U4726 (N_4726,In_1384,In_659);
nand U4727 (N_4727,In_1053,In_645);
nand U4728 (N_4728,In_59,In_1019);
or U4729 (N_4729,In_545,In_808);
nor U4730 (N_4730,In_997,In_1470);
and U4731 (N_4731,In_796,In_761);
and U4732 (N_4732,In_889,In_1971);
nor U4733 (N_4733,In_173,In_366);
or U4734 (N_4734,In_1965,In_659);
nand U4735 (N_4735,In_475,In_950);
nor U4736 (N_4736,In_657,In_1054);
and U4737 (N_4737,In_1272,In_103);
nand U4738 (N_4738,In_215,In_1620);
or U4739 (N_4739,In_366,In_1694);
nor U4740 (N_4740,In_522,In_250);
nor U4741 (N_4741,In_280,In_1995);
xor U4742 (N_4742,In_1187,In_897);
nor U4743 (N_4743,In_472,In_1567);
nor U4744 (N_4744,In_1516,In_1148);
or U4745 (N_4745,In_72,In_166);
nand U4746 (N_4746,In_285,In_328);
nand U4747 (N_4747,In_184,In_229);
nand U4748 (N_4748,In_1957,In_803);
nor U4749 (N_4749,In_1703,In_1930);
nand U4750 (N_4750,In_1394,In_321);
nand U4751 (N_4751,In_1847,In_1348);
and U4752 (N_4752,In_400,In_693);
nand U4753 (N_4753,In_1119,In_223);
nand U4754 (N_4754,In_1884,In_1685);
or U4755 (N_4755,In_297,In_1882);
or U4756 (N_4756,In_240,In_217);
xor U4757 (N_4757,In_1507,In_78);
and U4758 (N_4758,In_1616,In_1153);
nand U4759 (N_4759,In_463,In_1591);
nor U4760 (N_4760,In_1644,In_567);
nor U4761 (N_4761,In_1330,In_307);
or U4762 (N_4762,In_1501,In_803);
nor U4763 (N_4763,In_1104,In_1644);
nor U4764 (N_4764,In_1259,In_790);
nand U4765 (N_4765,In_26,In_780);
nand U4766 (N_4766,In_1588,In_458);
xor U4767 (N_4767,In_543,In_1679);
nand U4768 (N_4768,In_43,In_409);
nor U4769 (N_4769,In_502,In_671);
nand U4770 (N_4770,In_1696,In_1545);
nand U4771 (N_4771,In_1828,In_749);
nand U4772 (N_4772,In_653,In_861);
and U4773 (N_4773,In_815,In_1327);
and U4774 (N_4774,In_1221,In_207);
or U4775 (N_4775,In_214,In_502);
nand U4776 (N_4776,In_145,In_1217);
nand U4777 (N_4777,In_1929,In_1408);
nor U4778 (N_4778,In_1917,In_616);
and U4779 (N_4779,In_1385,In_436);
nand U4780 (N_4780,In_1775,In_1359);
and U4781 (N_4781,In_101,In_788);
nor U4782 (N_4782,In_914,In_1668);
nor U4783 (N_4783,In_259,In_538);
nand U4784 (N_4784,In_182,In_1355);
or U4785 (N_4785,In_1866,In_1698);
nor U4786 (N_4786,In_1210,In_1514);
and U4787 (N_4787,In_1324,In_318);
and U4788 (N_4788,In_197,In_730);
or U4789 (N_4789,In_393,In_1761);
nor U4790 (N_4790,In_1345,In_1657);
xnor U4791 (N_4791,In_1630,In_1096);
or U4792 (N_4792,In_1028,In_1642);
or U4793 (N_4793,In_1794,In_378);
and U4794 (N_4794,In_1907,In_1497);
or U4795 (N_4795,In_777,In_1861);
or U4796 (N_4796,In_1880,In_646);
nand U4797 (N_4797,In_1273,In_1114);
nand U4798 (N_4798,In_1479,In_86);
or U4799 (N_4799,In_366,In_1391);
xnor U4800 (N_4800,In_1444,In_1568);
and U4801 (N_4801,In_731,In_1389);
nand U4802 (N_4802,In_765,In_1156);
or U4803 (N_4803,In_1015,In_780);
and U4804 (N_4804,In_635,In_725);
nand U4805 (N_4805,In_259,In_1311);
xor U4806 (N_4806,In_1282,In_27);
nor U4807 (N_4807,In_1259,In_876);
and U4808 (N_4808,In_1721,In_895);
xor U4809 (N_4809,In_1997,In_92);
and U4810 (N_4810,In_284,In_1138);
and U4811 (N_4811,In_1501,In_51);
and U4812 (N_4812,In_722,In_1932);
nor U4813 (N_4813,In_943,In_1513);
nor U4814 (N_4814,In_1595,In_22);
or U4815 (N_4815,In_1429,In_1179);
nor U4816 (N_4816,In_1178,In_796);
nand U4817 (N_4817,In_896,In_217);
nor U4818 (N_4818,In_1444,In_635);
or U4819 (N_4819,In_1766,In_18);
and U4820 (N_4820,In_176,In_762);
or U4821 (N_4821,In_132,In_155);
nand U4822 (N_4822,In_1806,In_1217);
xnor U4823 (N_4823,In_1426,In_1197);
nand U4824 (N_4824,In_1262,In_1449);
and U4825 (N_4825,In_1328,In_1324);
and U4826 (N_4826,In_1239,In_587);
nand U4827 (N_4827,In_938,In_1703);
xnor U4828 (N_4828,In_133,In_49);
and U4829 (N_4829,In_377,In_78);
nor U4830 (N_4830,In_1185,In_1090);
and U4831 (N_4831,In_796,In_1355);
nand U4832 (N_4832,In_1993,In_1066);
nand U4833 (N_4833,In_1209,In_435);
and U4834 (N_4834,In_235,In_1444);
nor U4835 (N_4835,In_1029,In_267);
and U4836 (N_4836,In_1949,In_1409);
or U4837 (N_4837,In_669,In_1018);
and U4838 (N_4838,In_644,In_1995);
and U4839 (N_4839,In_2,In_336);
and U4840 (N_4840,In_1924,In_432);
and U4841 (N_4841,In_633,In_1636);
nor U4842 (N_4842,In_617,In_857);
and U4843 (N_4843,In_1326,In_103);
nand U4844 (N_4844,In_464,In_172);
nand U4845 (N_4845,In_1090,In_830);
or U4846 (N_4846,In_858,In_1007);
or U4847 (N_4847,In_1672,In_1410);
nand U4848 (N_4848,In_713,In_201);
nor U4849 (N_4849,In_1306,In_1315);
nand U4850 (N_4850,In_1815,In_274);
nand U4851 (N_4851,In_1266,In_352);
or U4852 (N_4852,In_1520,In_1438);
nand U4853 (N_4853,In_1503,In_567);
xnor U4854 (N_4854,In_1799,In_1787);
and U4855 (N_4855,In_1691,In_92);
nor U4856 (N_4856,In_432,In_451);
and U4857 (N_4857,In_164,In_293);
or U4858 (N_4858,In_325,In_1801);
nand U4859 (N_4859,In_864,In_348);
or U4860 (N_4860,In_196,In_1207);
and U4861 (N_4861,In_213,In_1640);
and U4862 (N_4862,In_1788,In_76);
nor U4863 (N_4863,In_322,In_310);
or U4864 (N_4864,In_456,In_944);
and U4865 (N_4865,In_1880,In_1174);
and U4866 (N_4866,In_1499,In_513);
or U4867 (N_4867,In_1131,In_1942);
and U4868 (N_4868,In_1566,In_1606);
and U4869 (N_4869,In_1690,In_289);
and U4870 (N_4870,In_1992,In_520);
and U4871 (N_4871,In_783,In_43);
and U4872 (N_4872,In_702,In_1958);
or U4873 (N_4873,In_1552,In_1833);
or U4874 (N_4874,In_1272,In_467);
nand U4875 (N_4875,In_557,In_937);
nor U4876 (N_4876,In_2,In_350);
and U4877 (N_4877,In_1063,In_1192);
xor U4878 (N_4878,In_1478,In_177);
and U4879 (N_4879,In_910,In_586);
and U4880 (N_4880,In_145,In_894);
nor U4881 (N_4881,In_1998,In_1089);
and U4882 (N_4882,In_1205,In_1711);
or U4883 (N_4883,In_46,In_1221);
nor U4884 (N_4884,In_1901,In_494);
and U4885 (N_4885,In_779,In_561);
xnor U4886 (N_4886,In_429,In_35);
or U4887 (N_4887,In_668,In_1904);
nand U4888 (N_4888,In_1801,In_503);
nor U4889 (N_4889,In_111,In_493);
nor U4890 (N_4890,In_582,In_116);
xor U4891 (N_4891,In_866,In_328);
and U4892 (N_4892,In_1680,In_590);
nand U4893 (N_4893,In_1101,In_634);
and U4894 (N_4894,In_1162,In_1691);
and U4895 (N_4895,In_194,In_1105);
nand U4896 (N_4896,In_780,In_1186);
or U4897 (N_4897,In_472,In_785);
and U4898 (N_4898,In_214,In_1327);
or U4899 (N_4899,In_719,In_1396);
nor U4900 (N_4900,In_1708,In_162);
nand U4901 (N_4901,In_1785,In_1322);
nand U4902 (N_4902,In_794,In_175);
nand U4903 (N_4903,In_897,In_928);
nor U4904 (N_4904,In_1417,In_1438);
and U4905 (N_4905,In_1905,In_1999);
nor U4906 (N_4906,In_1449,In_495);
xor U4907 (N_4907,In_1612,In_1087);
or U4908 (N_4908,In_1349,In_819);
or U4909 (N_4909,In_469,In_1290);
and U4910 (N_4910,In_1131,In_1360);
nor U4911 (N_4911,In_1950,In_1999);
and U4912 (N_4912,In_1605,In_1395);
nor U4913 (N_4913,In_1717,In_750);
nor U4914 (N_4914,In_1064,In_887);
nor U4915 (N_4915,In_1307,In_1826);
nor U4916 (N_4916,In_355,In_1902);
nand U4917 (N_4917,In_1259,In_1961);
or U4918 (N_4918,In_120,In_1630);
or U4919 (N_4919,In_783,In_1415);
or U4920 (N_4920,In_1907,In_508);
nand U4921 (N_4921,In_364,In_595);
nand U4922 (N_4922,In_153,In_1016);
and U4923 (N_4923,In_1105,In_109);
and U4924 (N_4924,In_1296,In_881);
xnor U4925 (N_4925,In_1960,In_1024);
xor U4926 (N_4926,In_1839,In_596);
nand U4927 (N_4927,In_297,In_1576);
or U4928 (N_4928,In_1487,In_1740);
or U4929 (N_4929,In_1304,In_636);
or U4930 (N_4930,In_1191,In_1074);
nand U4931 (N_4931,In_1336,In_1223);
xnor U4932 (N_4932,In_561,In_1405);
or U4933 (N_4933,In_1877,In_125);
nand U4934 (N_4934,In_1244,In_327);
nand U4935 (N_4935,In_1413,In_1254);
nand U4936 (N_4936,In_336,In_1938);
nand U4937 (N_4937,In_1130,In_724);
or U4938 (N_4938,In_153,In_204);
nor U4939 (N_4939,In_255,In_1406);
nor U4940 (N_4940,In_634,In_1772);
or U4941 (N_4941,In_1032,In_1981);
nor U4942 (N_4942,In_1050,In_245);
nor U4943 (N_4943,In_1412,In_1924);
xnor U4944 (N_4944,In_488,In_1615);
nor U4945 (N_4945,In_394,In_1190);
nand U4946 (N_4946,In_1312,In_1438);
and U4947 (N_4947,In_244,In_424);
nand U4948 (N_4948,In_430,In_1801);
nand U4949 (N_4949,In_1946,In_1367);
xor U4950 (N_4950,In_1789,In_1586);
and U4951 (N_4951,In_1752,In_816);
or U4952 (N_4952,In_939,In_1071);
nor U4953 (N_4953,In_1571,In_1251);
or U4954 (N_4954,In_1413,In_901);
or U4955 (N_4955,In_1885,In_1903);
and U4956 (N_4956,In_1508,In_1467);
or U4957 (N_4957,In_1125,In_265);
or U4958 (N_4958,In_1751,In_1553);
nor U4959 (N_4959,In_548,In_1979);
and U4960 (N_4960,In_32,In_927);
nand U4961 (N_4961,In_430,In_1502);
or U4962 (N_4962,In_1936,In_1308);
nor U4963 (N_4963,In_714,In_671);
and U4964 (N_4964,In_1072,In_1828);
or U4965 (N_4965,In_146,In_1657);
or U4966 (N_4966,In_1382,In_997);
and U4967 (N_4967,In_944,In_1431);
nand U4968 (N_4968,In_476,In_1523);
nand U4969 (N_4969,In_1035,In_1602);
nor U4970 (N_4970,In_1083,In_1135);
nor U4971 (N_4971,In_1418,In_1821);
nor U4972 (N_4972,In_63,In_1242);
xnor U4973 (N_4973,In_1690,In_492);
nor U4974 (N_4974,In_471,In_435);
or U4975 (N_4975,In_1280,In_1957);
xor U4976 (N_4976,In_1378,In_1850);
nor U4977 (N_4977,In_10,In_668);
xnor U4978 (N_4978,In_1877,In_1869);
and U4979 (N_4979,In_617,In_1530);
nand U4980 (N_4980,In_1246,In_852);
nor U4981 (N_4981,In_988,In_1874);
or U4982 (N_4982,In_787,In_1826);
or U4983 (N_4983,In_458,In_1228);
nor U4984 (N_4984,In_1195,In_1958);
nor U4985 (N_4985,In_564,In_1581);
nor U4986 (N_4986,In_626,In_1817);
xnor U4987 (N_4987,In_550,In_1543);
or U4988 (N_4988,In_1182,In_1303);
and U4989 (N_4989,In_183,In_1407);
nor U4990 (N_4990,In_1225,In_1669);
nor U4991 (N_4991,In_1822,In_605);
nor U4992 (N_4992,In_1743,In_1914);
and U4993 (N_4993,In_257,In_740);
nor U4994 (N_4994,In_1318,In_1099);
and U4995 (N_4995,In_1971,In_1342);
nor U4996 (N_4996,In_1573,In_567);
xnor U4997 (N_4997,In_834,In_1611);
or U4998 (N_4998,In_244,In_1079);
and U4999 (N_4999,In_298,In_1211);
and U5000 (N_5000,N_1752,N_300);
nand U5001 (N_5001,N_2948,N_1037);
or U5002 (N_5002,N_1821,N_1310);
nand U5003 (N_5003,N_2006,N_1942);
or U5004 (N_5004,N_3914,N_3047);
nand U5005 (N_5005,N_3775,N_3796);
xnor U5006 (N_5006,N_1934,N_1580);
nor U5007 (N_5007,N_515,N_880);
nor U5008 (N_5008,N_979,N_2188);
or U5009 (N_5009,N_1237,N_1406);
or U5010 (N_5010,N_4543,N_583);
nor U5011 (N_5011,N_633,N_1043);
and U5012 (N_5012,N_1383,N_1996);
or U5013 (N_5013,N_111,N_3098);
nor U5014 (N_5014,N_2640,N_2865);
nand U5015 (N_5015,N_3686,N_3150);
or U5016 (N_5016,N_2914,N_3334);
nor U5017 (N_5017,N_985,N_4530);
and U5018 (N_5018,N_1687,N_4977);
or U5019 (N_5019,N_1568,N_2126);
xor U5020 (N_5020,N_2412,N_2148);
and U5021 (N_5021,N_744,N_3399);
nor U5022 (N_5022,N_1101,N_231);
nor U5023 (N_5023,N_4152,N_3149);
and U5024 (N_5024,N_390,N_4959);
and U5025 (N_5025,N_3541,N_2060);
or U5026 (N_5026,N_3261,N_2120);
nor U5027 (N_5027,N_198,N_4555);
and U5028 (N_5028,N_4046,N_1407);
nor U5029 (N_5029,N_1901,N_648);
nand U5030 (N_5030,N_146,N_2281);
xor U5031 (N_5031,N_704,N_121);
nor U5032 (N_5032,N_3134,N_1097);
or U5033 (N_5033,N_3614,N_4586);
nor U5034 (N_5034,N_2904,N_1482);
nor U5035 (N_5035,N_1960,N_2354);
nand U5036 (N_5036,N_1065,N_4911);
nand U5037 (N_5037,N_3468,N_3878);
or U5038 (N_5038,N_3429,N_2316);
nand U5039 (N_5039,N_2793,N_82);
xor U5040 (N_5040,N_2759,N_1143);
or U5041 (N_5041,N_4989,N_2703);
nand U5042 (N_5042,N_1606,N_4539);
nand U5043 (N_5043,N_4151,N_4860);
or U5044 (N_5044,N_2272,N_931);
or U5045 (N_5045,N_2372,N_2984);
and U5046 (N_5046,N_1435,N_2743);
xor U5047 (N_5047,N_3644,N_1330);
nor U5048 (N_5048,N_4522,N_3832);
or U5049 (N_5049,N_351,N_2783);
nor U5050 (N_5050,N_2943,N_997);
nand U5051 (N_5051,N_2066,N_1793);
nand U5052 (N_5052,N_4275,N_1259);
nand U5053 (N_5053,N_2061,N_793);
nand U5054 (N_5054,N_3849,N_2645);
nand U5055 (N_5055,N_716,N_3671);
nor U5056 (N_5056,N_16,N_1367);
xor U5057 (N_5057,N_2509,N_2052);
xor U5058 (N_5058,N_2219,N_2920);
or U5059 (N_5059,N_2871,N_968);
xnor U5060 (N_5060,N_508,N_2000);
nand U5061 (N_5061,N_4095,N_4965);
and U5062 (N_5062,N_2994,N_4323);
or U5063 (N_5063,N_4613,N_4225);
nor U5064 (N_5064,N_4643,N_4341);
nand U5065 (N_5065,N_4435,N_4049);
nor U5066 (N_5066,N_3127,N_2970);
nand U5067 (N_5067,N_1211,N_2303);
or U5068 (N_5068,N_3206,N_1356);
nand U5069 (N_5069,N_3940,N_2518);
or U5070 (N_5070,N_2681,N_4150);
and U5071 (N_5071,N_3948,N_542);
nand U5072 (N_5072,N_1648,N_4708);
nor U5073 (N_5073,N_1060,N_3110);
and U5074 (N_5074,N_3576,N_4483);
nor U5075 (N_5075,N_1959,N_2873);
or U5076 (N_5076,N_875,N_714);
nor U5077 (N_5077,N_4388,N_2696);
and U5078 (N_5078,N_2905,N_1739);
nor U5079 (N_5079,N_4358,N_2433);
nor U5080 (N_5080,N_3342,N_4319);
nand U5081 (N_5081,N_682,N_4291);
or U5082 (N_5082,N_1191,N_4104);
nor U5083 (N_5083,N_1714,N_1857);
xnor U5084 (N_5084,N_1472,N_273);
xor U5085 (N_5085,N_4656,N_2773);
nand U5086 (N_5086,N_3091,N_976);
nand U5087 (N_5087,N_750,N_1167);
nor U5088 (N_5088,N_2388,N_1230);
nand U5089 (N_5089,N_1437,N_22);
nor U5090 (N_5090,N_537,N_3709);
nand U5091 (N_5091,N_4966,N_3318);
nor U5092 (N_5092,N_476,N_1339);
nand U5093 (N_5093,N_4187,N_3919);
nor U5094 (N_5094,N_72,N_2860);
and U5095 (N_5095,N_4464,N_4392);
or U5096 (N_5096,N_2157,N_3761);
xnor U5097 (N_5097,N_915,N_3750);
and U5098 (N_5098,N_850,N_895);
xnor U5099 (N_5099,N_4767,N_3771);
or U5100 (N_5100,N_2642,N_1993);
nor U5101 (N_5101,N_4135,N_237);
nand U5102 (N_5102,N_3651,N_993);
nor U5103 (N_5103,N_173,N_1617);
and U5104 (N_5104,N_942,N_230);
nor U5105 (N_5105,N_155,N_2111);
xnor U5106 (N_5106,N_1994,N_2238);
xnor U5107 (N_5107,N_321,N_2532);
and U5108 (N_5108,N_1138,N_3550);
or U5109 (N_5109,N_1907,N_3233);
nand U5110 (N_5110,N_2898,N_952);
nand U5111 (N_5111,N_2715,N_1758);
or U5112 (N_5112,N_3143,N_3662);
nor U5113 (N_5113,N_590,N_1061);
xnor U5114 (N_5114,N_2853,N_3126);
nor U5115 (N_5115,N_4321,N_70);
nor U5116 (N_5116,N_2443,N_4824);
and U5117 (N_5117,N_3743,N_3856);
nand U5118 (N_5118,N_2932,N_2561);
xnor U5119 (N_5119,N_3262,N_4426);
and U5120 (N_5120,N_352,N_1556);
or U5121 (N_5121,N_3284,N_2930);
nand U5122 (N_5122,N_1351,N_177);
xor U5123 (N_5123,N_885,N_3631);
and U5124 (N_5124,N_2494,N_4093);
nand U5125 (N_5125,N_2396,N_1868);
xnor U5126 (N_5126,N_1668,N_4203);
and U5127 (N_5127,N_3257,N_3417);
nand U5128 (N_5128,N_729,N_1995);
or U5129 (N_5129,N_4611,N_4666);
nand U5130 (N_5130,N_3986,N_1627);
nand U5131 (N_5131,N_1346,N_99);
or U5132 (N_5132,N_3546,N_1767);
and U5133 (N_5133,N_2310,N_1615);
and U5134 (N_5134,N_1145,N_40);
and U5135 (N_5135,N_50,N_1587);
nand U5136 (N_5136,N_734,N_792);
nand U5137 (N_5137,N_992,N_1373);
and U5138 (N_5138,N_3868,N_4448);
nand U5139 (N_5139,N_1140,N_3368);
or U5140 (N_5140,N_2840,N_3204);
nand U5141 (N_5141,N_2130,N_677);
nand U5142 (N_5142,N_4159,N_4598);
and U5143 (N_5143,N_4958,N_2549);
nand U5144 (N_5144,N_675,N_4513);
nand U5145 (N_5145,N_4637,N_2809);
and U5146 (N_5146,N_1766,N_4430);
nand U5147 (N_5147,N_3652,N_4905);
xor U5148 (N_5148,N_3305,N_4295);
nor U5149 (N_5149,N_614,N_3747);
or U5150 (N_5150,N_4306,N_4806);
xnor U5151 (N_5151,N_2990,N_4067);
or U5152 (N_5152,N_2530,N_3287);
nand U5153 (N_5153,N_4407,N_4969);
or U5154 (N_5154,N_1799,N_2747);
xor U5155 (N_5155,N_4101,N_3977);
and U5156 (N_5156,N_876,N_1770);
nand U5157 (N_5157,N_3044,N_2401);
xnor U5158 (N_5158,N_4953,N_2967);
nand U5159 (N_5159,N_960,N_4331);
nand U5160 (N_5160,N_1813,N_4444);
and U5161 (N_5161,N_328,N_2191);
nor U5162 (N_5162,N_4970,N_1391);
or U5163 (N_5163,N_651,N_4940);
nor U5164 (N_5164,N_883,N_3441);
nor U5165 (N_5165,N_18,N_2226);
nor U5166 (N_5166,N_3907,N_4029);
and U5167 (N_5167,N_3952,N_4593);
and U5168 (N_5168,N_3934,N_688);
nor U5169 (N_5169,N_4421,N_849);
or U5170 (N_5170,N_2664,N_4785);
nor U5171 (N_5171,N_3202,N_1258);
and U5172 (N_5172,N_4145,N_4719);
nand U5173 (N_5173,N_1011,N_160);
and U5174 (N_5174,N_3293,N_4914);
xnor U5175 (N_5175,N_740,N_3386);
and U5176 (N_5176,N_4147,N_2755);
or U5177 (N_5177,N_721,N_969);
nor U5178 (N_5178,N_5,N_218);
or U5179 (N_5179,N_4610,N_1763);
nand U5180 (N_5180,N_569,N_1871);
nor U5181 (N_5181,N_391,N_3249);
or U5182 (N_5182,N_4237,N_144);
nand U5183 (N_5183,N_2258,N_996);
or U5184 (N_5184,N_832,N_748);
and U5185 (N_5185,N_2260,N_4428);
nand U5186 (N_5186,N_559,N_2545);
and U5187 (N_5187,N_835,N_54);
nor U5188 (N_5188,N_861,N_3697);
xnor U5189 (N_5189,N_776,N_127);
and U5190 (N_5190,N_1120,N_4747);
and U5191 (N_5191,N_1386,N_3398);
nor U5192 (N_5192,N_1914,N_547);
and U5193 (N_5193,N_4238,N_1991);
and U5194 (N_5194,N_4632,N_4776);
nand U5195 (N_5195,N_4654,N_3502);
and U5196 (N_5196,N_3708,N_89);
nor U5197 (N_5197,N_2856,N_2383);
and U5198 (N_5198,N_804,N_1382);
nand U5199 (N_5199,N_4784,N_3496);
or U5200 (N_5200,N_1374,N_3256);
or U5201 (N_5201,N_818,N_4434);
nor U5202 (N_5202,N_1129,N_3620);
and U5203 (N_5203,N_2968,N_1338);
nand U5204 (N_5204,N_836,N_1190);
or U5205 (N_5205,N_1673,N_4329);
xnor U5206 (N_5206,N_1210,N_653);
xnor U5207 (N_5207,N_4916,N_2916);
or U5208 (N_5208,N_2580,N_2496);
nand U5209 (N_5209,N_27,N_2712);
or U5210 (N_5210,N_3933,N_662);
or U5211 (N_5211,N_1173,N_2581);
nand U5212 (N_5212,N_2470,N_529);
xor U5213 (N_5213,N_946,N_3808);
or U5214 (N_5214,N_1912,N_2195);
and U5215 (N_5215,N_4651,N_2169);
nand U5216 (N_5216,N_2381,N_1415);
nand U5217 (N_5217,N_429,N_3029);
xnor U5218 (N_5218,N_2570,N_3749);
or U5219 (N_5219,N_227,N_1042);
or U5220 (N_5220,N_4886,N_178);
nand U5221 (N_5221,N_4597,N_2972);
and U5222 (N_5222,N_596,N_140);
or U5223 (N_5223,N_920,N_4697);
nand U5224 (N_5224,N_4134,N_2056);
and U5225 (N_5225,N_787,N_3894);
nor U5226 (N_5226,N_343,N_3874);
nor U5227 (N_5227,N_3535,N_600);
or U5228 (N_5228,N_3273,N_4142);
or U5229 (N_5229,N_340,N_767);
and U5230 (N_5230,N_1126,N_4762);
nor U5231 (N_5231,N_2467,N_1968);
nand U5232 (N_5232,N_1029,N_2334);
and U5233 (N_5233,N_1711,N_4296);
and U5234 (N_5234,N_1267,N_3279);
and U5235 (N_5235,N_989,N_2838);
and U5236 (N_5236,N_760,N_277);
and U5237 (N_5237,N_986,N_3567);
nand U5238 (N_5238,N_110,N_1581);
nor U5239 (N_5239,N_3325,N_4245);
nor U5240 (N_5240,N_1956,N_195);
nand U5241 (N_5241,N_1908,N_1263);
nor U5242 (N_5242,N_131,N_4128);
or U5243 (N_5243,N_2718,N_2523);
xor U5244 (N_5244,N_2894,N_3158);
xor U5245 (N_5245,N_4962,N_2812);
or U5246 (N_5246,N_2289,N_3391);
nor U5247 (N_5247,N_3676,N_1163);
nor U5248 (N_5248,N_1342,N_3847);
or U5249 (N_5249,N_326,N_680);
nand U5250 (N_5250,N_2446,N_2304);
or U5251 (N_5251,N_404,N_935);
nor U5252 (N_5252,N_2662,N_4172);
xor U5253 (N_5253,N_3632,N_4749);
xor U5254 (N_5254,N_3007,N_48);
xnor U5255 (N_5255,N_2410,N_471);
nor U5256 (N_5256,N_179,N_2674);
or U5257 (N_5257,N_2560,N_3086);
or U5258 (N_5258,N_939,N_1781);
xor U5259 (N_5259,N_4185,N_810);
nor U5260 (N_5260,N_3478,N_3037);
xor U5261 (N_5261,N_3104,N_2734);
nor U5262 (N_5262,N_3053,N_1731);
or U5263 (N_5263,N_2054,N_3359);
or U5264 (N_5264,N_1955,N_4866);
nand U5265 (N_5265,N_4452,N_4362);
nor U5266 (N_5266,N_341,N_1710);
nor U5267 (N_5267,N_3673,N_2697);
or U5268 (N_5268,N_1832,N_13);
nor U5269 (N_5269,N_2824,N_4549);
nor U5270 (N_5270,N_225,N_4960);
or U5271 (N_5271,N_1332,N_3794);
xnor U5272 (N_5272,N_2680,N_2183);
and U5273 (N_5273,N_3175,N_3696);
nand U5274 (N_5274,N_1797,N_3088);
or U5275 (N_5275,N_1574,N_4389);
xnor U5276 (N_5276,N_758,N_3000);
nor U5277 (N_5277,N_1886,N_3635);
nor U5278 (N_5278,N_1474,N_4397);
nor U5279 (N_5279,N_4173,N_3278);
nand U5280 (N_5280,N_3063,N_1679);
and U5281 (N_5281,N_2187,N_248);
xnor U5282 (N_5282,N_3013,N_1814);
and U5283 (N_5283,N_2373,N_3283);
xor U5284 (N_5284,N_3165,N_2101);
nand U5285 (N_5285,N_3473,N_4683);
nand U5286 (N_5286,N_4703,N_1557);
xor U5287 (N_5287,N_794,N_1483);
xnor U5288 (N_5288,N_3485,N_1949);
or U5289 (N_5289,N_4460,N_4222);
nand U5290 (N_5290,N_3804,N_4715);
xnor U5291 (N_5291,N_438,N_2892);
and U5292 (N_5292,N_3394,N_2269);
nand U5293 (N_5293,N_4303,N_655);
and U5294 (N_5294,N_3397,N_2019);
nor U5295 (N_5295,N_3913,N_3595);
xnor U5296 (N_5296,N_2297,N_995);
nor U5297 (N_5297,N_4823,N_2225);
or U5298 (N_5298,N_1108,N_3511);
and U5299 (N_5299,N_4422,N_2139);
and U5300 (N_5300,N_4190,N_3460);
nand U5301 (N_5301,N_1139,N_423);
or U5302 (N_5302,N_4299,N_1780);
or U5303 (N_5303,N_927,N_1262);
and U5304 (N_5304,N_4284,N_2985);
xnor U5305 (N_5305,N_3319,N_1100);
nor U5306 (N_5306,N_3034,N_2806);
nor U5307 (N_5307,N_4164,N_3748);
or U5308 (N_5308,N_2814,N_4809);
nand U5309 (N_5309,N_2579,N_1840);
and U5310 (N_5310,N_2822,N_4277);
xnor U5311 (N_5311,N_998,N_1798);
nor U5312 (N_5312,N_2090,N_1368);
or U5313 (N_5313,N_1461,N_944);
and U5314 (N_5314,N_2369,N_2236);
xor U5315 (N_5315,N_4980,N_4356);
or U5316 (N_5316,N_119,N_557);
or U5317 (N_5317,N_216,N_694);
or U5318 (N_5318,N_4106,N_339);
and U5319 (N_5319,N_1678,N_4605);
xnor U5320 (N_5320,N_4213,N_1327);
or U5321 (N_5321,N_2785,N_4721);
or U5322 (N_5322,N_1031,N_3897);
xor U5323 (N_5323,N_3717,N_4794);
or U5324 (N_5324,N_4402,N_2377);
or U5325 (N_5325,N_2098,N_3813);
and U5326 (N_5326,N_2828,N_1958);
nor U5327 (N_5327,N_2360,N_4459);
and U5328 (N_5328,N_3978,N_676);
or U5329 (N_5329,N_3869,N_4254);
and U5330 (N_5330,N_2729,N_3090);
nor U5331 (N_5331,N_1241,N_1620);
nor U5332 (N_5332,N_4585,N_2908);
nor U5333 (N_5333,N_1089,N_234);
nor U5334 (N_5334,N_2142,N_3375);
xor U5335 (N_5335,N_859,N_3764);
nor U5336 (N_5336,N_2062,N_811);
nand U5337 (N_5337,N_900,N_3809);
and U5338 (N_5338,N_1257,N_309);
xnor U5339 (N_5339,N_673,N_3315);
and U5340 (N_5340,N_1876,N_3976);
nor U5341 (N_5341,N_392,N_3547);
and U5342 (N_5342,N_2278,N_4206);
or U5343 (N_5343,N_1188,N_2163);
and U5344 (N_5344,N_666,N_4207);
and U5345 (N_5345,N_732,N_4639);
nand U5346 (N_5346,N_4451,N_1693);
and U5347 (N_5347,N_1401,N_2843);
and U5348 (N_5348,N_2884,N_4896);
and U5349 (N_5349,N_3757,N_4100);
nand U5350 (N_5350,N_3751,N_428);
nor U5351 (N_5351,N_3639,N_348);
or U5352 (N_5352,N_1791,N_1699);
nand U5353 (N_5353,N_3312,N_1891);
nand U5354 (N_5354,N_3017,N_4236);
nor U5355 (N_5355,N_1283,N_2152);
nand U5356 (N_5356,N_868,N_4034);
and U5357 (N_5357,N_2605,N_3226);
nand U5358 (N_5358,N_58,N_841);
nand U5359 (N_5359,N_2121,N_3211);
nand U5360 (N_5360,N_521,N_2711);
and U5361 (N_5361,N_1535,N_3594);
nand U5362 (N_5362,N_2901,N_4338);
nand U5363 (N_5363,N_4700,N_4913);
nor U5364 (N_5364,N_4900,N_2736);
nand U5365 (N_5365,N_23,N_4230);
xor U5366 (N_5366,N_1228,N_4017);
or U5367 (N_5367,N_604,N_3092);
and U5368 (N_5368,N_1659,N_2237);
nand U5369 (N_5369,N_1526,N_3139);
or U5370 (N_5370,N_3026,N_1625);
and U5371 (N_5371,N_3182,N_3831);
nand U5372 (N_5372,N_4671,N_2848);
nor U5373 (N_5373,N_2543,N_1585);
nand U5374 (N_5374,N_3715,N_4790);
or U5375 (N_5375,N_4045,N_3664);
and U5376 (N_5376,N_4804,N_3393);
or U5377 (N_5377,N_298,N_2285);
or U5378 (N_5378,N_860,N_3536);
xor U5379 (N_5379,N_4871,N_191);
nand U5380 (N_5380,N_2874,N_1005);
nand U5381 (N_5381,N_2691,N_1900);
or U5382 (N_5382,N_2010,N_2105);
or U5383 (N_5383,N_2078,N_2170);
nand U5384 (N_5384,N_501,N_460);
nand U5385 (N_5385,N_2256,N_1085);
or U5386 (N_5386,N_4276,N_2255);
xor U5387 (N_5387,N_4372,N_1986);
and U5388 (N_5388,N_3835,N_4390);
and U5389 (N_5389,N_2673,N_3844);
nand U5390 (N_5390,N_2870,N_1599);
or U5391 (N_5391,N_3077,N_4975);
nand U5392 (N_5392,N_2322,N_4133);
nand U5393 (N_5393,N_3337,N_1296);
and U5394 (N_5394,N_4579,N_1937);
xor U5395 (N_5395,N_2820,N_4878);
nand U5396 (N_5396,N_3285,N_2858);
xnor U5397 (N_5397,N_1183,N_1252);
or U5398 (N_5398,N_3274,N_167);
or U5399 (N_5399,N_4786,N_4509);
or U5400 (N_5400,N_1424,N_588);
and U5401 (N_5401,N_1582,N_2317);
and U5402 (N_5402,N_640,N_544);
xnor U5403 (N_5403,N_1475,N_966);
nor U5404 (N_5404,N_1355,N_3358);
and U5405 (N_5405,N_2244,N_367);
and U5406 (N_5406,N_4746,N_1631);
xnor U5407 (N_5407,N_2155,N_3304);
xor U5408 (N_5408,N_3069,N_1591);
or U5409 (N_5409,N_3670,N_2723);
nor U5410 (N_5410,N_621,N_4355);
or U5411 (N_5411,N_1851,N_1334);
and U5412 (N_5412,N_1450,N_3520);
xnor U5413 (N_5413,N_3828,N_858);
and U5414 (N_5414,N_725,N_4377);
nor U5415 (N_5415,N_467,N_3824);
nand U5416 (N_5416,N_1322,N_162);
or U5417 (N_5417,N_4853,N_2063);
nand U5418 (N_5418,N_2676,N_685);
xor U5419 (N_5419,N_3310,N_3690);
nor U5420 (N_5420,N_3309,N_2328);
xor U5421 (N_5421,N_3028,N_539);
nand U5422 (N_5422,N_2290,N_4116);
xor U5423 (N_5423,N_143,N_1728);
nor U5424 (N_5424,N_1723,N_1842);
or U5425 (N_5425,N_1260,N_1657);
nor U5426 (N_5426,N_416,N_536);
xor U5427 (N_5427,N_3163,N_2732);
xor U5428 (N_5428,N_4760,N_3210);
and U5429 (N_5429,N_586,N_1874);
nand U5430 (N_5430,N_1432,N_2154);
nand U5431 (N_5431,N_364,N_2603);
or U5432 (N_5432,N_645,N_1469);
and U5433 (N_5433,N_1193,N_2082);
nand U5434 (N_5434,N_1047,N_4403);
nor U5435 (N_5435,N_2253,N_1281);
and U5436 (N_5436,N_4630,N_1205);
nor U5437 (N_5437,N_712,N_3138);
nand U5438 (N_5438,N_2131,N_3445);
or U5439 (N_5439,N_132,N_270);
and U5440 (N_5440,N_2533,N_2014);
xor U5441 (N_5441,N_2005,N_2153);
nor U5442 (N_5442,N_3964,N_3011);
nor U5443 (N_5443,N_3787,N_4270);
nor U5444 (N_5444,N_1966,N_1465);
or U5445 (N_5445,N_943,N_4782);
nand U5446 (N_5446,N_1265,N_228);
xnor U5447 (N_5447,N_4305,N_4234);
and U5448 (N_5448,N_2716,N_3132);
nor U5449 (N_5449,N_3850,N_4040);
and U5450 (N_5450,N_454,N_464);
or U5451 (N_5451,N_3649,N_3969);
and U5452 (N_5452,N_157,N_4582);
or U5453 (N_5453,N_3323,N_1292);
nor U5454 (N_5454,N_1529,N_4625);
or U5455 (N_5455,N_1387,N_3626);
nand U5456 (N_5456,N_1936,N_1690);
xnor U5457 (N_5457,N_3338,N_2689);
nand U5458 (N_5458,N_4877,N_4327);
and U5459 (N_5459,N_2162,N_3857);
or U5460 (N_5460,N_4132,N_124);
or U5461 (N_5461,N_602,N_4240);
nor U5462 (N_5462,N_4548,N_3074);
nor U5463 (N_5463,N_4699,N_2181);
nor U5464 (N_5464,N_2086,N_3513);
or U5465 (N_5465,N_4812,N_607);
nor U5466 (N_5466,N_2678,N_159);
and U5467 (N_5467,N_4819,N_2831);
and U5468 (N_5468,N_3612,N_3995);
nand U5469 (N_5469,N_2983,N_2215);
and U5470 (N_5470,N_4153,N_2531);
or U5471 (N_5471,N_749,N_4612);
nor U5472 (N_5472,N_4026,N_1428);
nand U5473 (N_5473,N_4165,N_784);
nand U5474 (N_5474,N_3606,N_4365);
and U5475 (N_5475,N_739,N_2941);
xnor U5476 (N_5476,N_3437,N_2100);
nor U5477 (N_5477,N_1247,N_3954);
and U5478 (N_5478,N_1841,N_3642);
or U5479 (N_5479,N_2522,N_4494);
xnor U5480 (N_5480,N_2677,N_3101);
nand U5481 (N_5481,N_65,N_4366);
nand U5482 (N_5482,N_3871,N_1160);
nor U5483 (N_5483,N_3766,N_213);
and U5484 (N_5484,N_4503,N_104);
and U5485 (N_5485,N_2659,N_450);
or U5486 (N_5486,N_3219,N_4086);
or U5487 (N_5487,N_2817,N_4768);
or U5488 (N_5488,N_896,N_93);
nor U5489 (N_5489,N_532,N_909);
or U5490 (N_5490,N_797,N_2786);
nor U5491 (N_5491,N_2319,N_1946);
nand U5492 (N_5492,N_3842,N_4599);
or U5493 (N_5493,N_2031,N_1048);
or U5494 (N_5494,N_3554,N_4205);
or U5495 (N_5495,N_2210,N_1175);
nor U5496 (N_5496,N_4928,N_452);
nor U5497 (N_5497,N_4438,N_2043);
nand U5498 (N_5498,N_4043,N_623);
or U5499 (N_5499,N_2850,N_2899);
and U5500 (N_5500,N_812,N_135);
nand U5501 (N_5501,N_4525,N_870);
nand U5502 (N_5502,N_1158,N_387);
nand U5503 (N_5503,N_2293,N_1222);
or U5504 (N_5504,N_64,N_1308);
nand U5505 (N_5505,N_299,N_2576);
nor U5506 (N_5506,N_2032,N_4171);
xor U5507 (N_5507,N_2646,N_3753);
nand U5508 (N_5508,N_4385,N_2787);
and U5509 (N_5509,N_3943,N_3930);
xor U5510 (N_5510,N_1273,N_4728);
and U5511 (N_5511,N_2915,N_1419);
nand U5512 (N_5512,N_4742,N_3270);
and U5513 (N_5513,N_2637,N_32);
xor U5514 (N_5514,N_2113,N_689);
nor U5515 (N_5515,N_2452,N_2171);
nor U5516 (N_5516,N_706,N_4440);
or U5517 (N_5517,N_903,N_1704);
nand U5518 (N_5518,N_3941,N_4198);
or U5519 (N_5519,N_632,N_2292);
or U5520 (N_5520,N_2478,N_3744);
xor U5521 (N_5521,N_3590,N_4083);
nand U5522 (N_5522,N_3816,N_4357);
or U5523 (N_5523,N_3531,N_4033);
nand U5524 (N_5524,N_3432,N_887);
or U5525 (N_5525,N_2069,N_499);
and U5526 (N_5526,N_3385,N_2525);
and U5527 (N_5527,N_1982,N_1862);
nand U5528 (N_5528,N_2233,N_3458);
and U5529 (N_5529,N_2857,N_4938);
nand U5530 (N_5530,N_2947,N_3984);
nor U5531 (N_5531,N_1794,N_4955);
nor U5532 (N_5532,N_3275,N_2012);
xnor U5533 (N_5533,N_4710,N_2800);
nor U5534 (N_5534,N_759,N_4396);
and U5535 (N_5535,N_2519,N_3981);
nor U5536 (N_5536,N_2978,N_2627);
nand U5537 (N_5537,N_9,N_4988);
nor U5538 (N_5538,N_1082,N_2168);
and U5539 (N_5539,N_327,N_275);
and U5540 (N_5540,N_1447,N_3518);
nor U5541 (N_5541,N_6,N_3166);
and U5542 (N_5542,N_4813,N_240);
and U5543 (N_5543,N_4791,N_4091);
or U5544 (N_5544,N_936,N_3180);
and U5545 (N_5545,N_779,N_3888);
or U5546 (N_5546,N_626,N_2474);
or U5547 (N_5547,N_2117,N_1052);
nand U5548 (N_5548,N_2422,N_1480);
and U5549 (N_5549,N_3452,N_4808);
or U5550 (N_5550,N_1913,N_874);
and U5551 (N_5551,N_504,N_1306);
or U5552 (N_5552,N_2852,N_2655);
or U5553 (N_5553,N_3030,N_2600);
nor U5554 (N_5554,N_1899,N_4224);
nand U5555 (N_5555,N_381,N_2635);
nor U5556 (N_5556,N_4537,N_1990);
nor U5557 (N_5557,N_2589,N_4879);
or U5558 (N_5558,N_2752,N_35);
and U5559 (N_5559,N_1282,N_4904);
nor U5560 (N_5560,N_1076,N_2832);
or U5561 (N_5561,N_4491,N_3054);
nor U5562 (N_5562,N_518,N_1542);
nor U5563 (N_5563,N_1449,N_863);
and U5564 (N_5564,N_1333,N_629);
nand U5565 (N_5565,N_795,N_3768);
xor U5566 (N_5566,N_4881,N_1579);
nand U5567 (N_5567,N_4758,N_620);
nor U5568 (N_5568,N_4924,N_1411);
nor U5569 (N_5569,N_1553,N_643);
nand U5570 (N_5570,N_446,N_370);
xor U5571 (N_5571,N_3797,N_2287);
nand U5572 (N_5572,N_3018,N_3726);
nand U5573 (N_5573,N_1506,N_2829);
nor U5574 (N_5574,N_1860,N_644);
nand U5575 (N_5575,N_2562,N_2555);
nor U5576 (N_5576,N_3488,N_2628);
and U5577 (N_5577,N_2683,N_4175);
nor U5578 (N_5578,N_2072,N_4925);
and U5579 (N_5579,N_1674,N_3727);
nor U5580 (N_5580,N_2342,N_2623);
nand U5581 (N_5581,N_42,N_4986);
xor U5582 (N_5582,N_3860,N_1083);
or U5583 (N_5583,N_1132,N_1818);
nor U5584 (N_5584,N_3314,N_3401);
and U5585 (N_5585,N_1541,N_4484);
nand U5586 (N_5586,N_284,N_3200);
or U5587 (N_5587,N_2492,N_123);
or U5588 (N_5588,N_4344,N_2748);
nand U5589 (N_5589,N_2073,N_545);
nor U5590 (N_5590,N_4517,N_3533);
nor U5591 (N_5591,N_1970,N_4678);
and U5592 (N_5592,N_530,N_485);
nand U5593 (N_5593,N_152,N_56);
or U5594 (N_5594,N_3553,N_2586);
nor U5595 (N_5595,N_2367,N_1438);
nor U5596 (N_5596,N_2359,N_3701);
nand U5597 (N_5597,N_1676,N_802);
or U5598 (N_5598,N_1989,N_796);
and U5599 (N_5599,N_2479,N_2867);
nand U5600 (N_5600,N_2788,N_2769);
and U5601 (N_5601,N_4156,N_3455);
nand U5602 (N_5602,N_2077,N_219);
nor U5603 (N_5603,N_3131,N_3173);
nand U5604 (N_5604,N_4243,N_4706);
and U5605 (N_5605,N_2704,N_3300);
or U5606 (N_5606,N_2665,N_3793);
xor U5607 (N_5607,N_350,N_2739);
and U5608 (N_5608,N_4265,N_315);
and U5609 (N_5609,N_527,N_631);
or U5610 (N_5610,N_1149,N_2669);
nand U5611 (N_5611,N_386,N_619);
and U5612 (N_5612,N_3362,N_2751);
and U5613 (N_5613,N_149,N_2700);
or U5614 (N_5614,N_1354,N_4951);
or U5615 (N_5615,N_2138,N_2639);
nand U5616 (N_5616,N_4393,N_4814);
nor U5617 (N_5617,N_3663,N_445);
nor U5618 (N_5618,N_4504,N_3827);
or U5619 (N_5619,N_4994,N_3725);
and U5620 (N_5620,N_4227,N_4076);
or U5621 (N_5621,N_456,N_3003);
nand U5622 (N_5622,N_3145,N_4105);
or U5623 (N_5623,N_3582,N_4992);
nor U5624 (N_5624,N_502,N_1514);
or U5625 (N_5625,N_1664,N_2413);
nor U5626 (N_5626,N_3691,N_2742);
nand U5627 (N_5627,N_4155,N_3956);
and U5628 (N_5628,N_3577,N_1055);
nand U5629 (N_5629,N_287,N_2505);
or U5630 (N_5630,N_4734,N_516);
or U5631 (N_5631,N_2140,N_1276);
nor U5632 (N_5632,N_490,N_768);
nand U5633 (N_5633,N_2942,N_1187);
and U5634 (N_5634,N_3355,N_4592);
nand U5635 (N_5635,N_1159,N_4316);
xnor U5636 (N_5636,N_187,N_3080);
nor U5637 (N_5637,N_274,N_4325);
or U5638 (N_5638,N_204,N_2517);
nor U5639 (N_5639,N_2468,N_3089);
nand U5640 (N_5640,N_4314,N_4112);
nor U5641 (N_5641,N_1170,N_260);
or U5642 (N_5642,N_1622,N_426);
nor U5643 (N_5643,N_2430,N_3530);
nor U5644 (N_5644,N_2308,N_1592);
or U5645 (N_5645,N_754,N_4607);
nand U5646 (N_5646,N_4416,N_742);
nor U5647 (N_5647,N_2550,N_973);
nand U5648 (N_5648,N_4594,N_1001);
nand U5649 (N_5649,N_29,N_3289);
or U5650 (N_5650,N_2456,N_2336);
or U5651 (N_5651,N_1018,N_4053);
nand U5652 (N_5652,N_3381,N_4457);
xnor U5653 (N_5653,N_2026,N_3846);
or U5654 (N_5654,N_1727,N_4129);
nand U5655 (N_5655,N_1750,N_840);
nand U5656 (N_5656,N_2976,N_1335);
nand U5657 (N_5657,N_4505,N_696);
nor U5658 (N_5658,N_878,N_399);
or U5659 (N_5659,N_1357,N_4263);
nor U5660 (N_5660,N_657,N_261);
or U5661 (N_5661,N_4113,N_3135);
xor U5662 (N_5662,N_4367,N_494);
nor U5663 (N_5663,N_2477,N_2361);
nor U5664 (N_5664,N_4339,N_453);
or U5665 (N_5665,N_4248,N_1921);
and U5666 (N_5666,N_1567,N_1106);
nor U5667 (N_5667,N_3129,N_3497);
nor U5668 (N_5668,N_1304,N_1870);
nand U5669 (N_5669,N_3414,N_4474);
nor U5670 (N_5670,N_1566,N_672);
nand U5671 (N_5671,N_3041,N_3230);
nand U5672 (N_5672,N_1467,N_929);
or U5673 (N_5673,N_2964,N_2542);
nor U5674 (N_5674,N_1786,N_1724);
or U5675 (N_5675,N_4292,N_4778);
and U5676 (N_5676,N_3361,N_1329);
nor U5677 (N_5677,N_3189,N_1174);
or U5678 (N_5678,N_1398,N_1460);
nor U5679 (N_5679,N_3246,N_1853);
or U5680 (N_5680,N_1720,N_2625);
and U5681 (N_5681,N_2213,N_3482);
nor U5682 (N_5682,N_4720,N_200);
nand U5683 (N_5683,N_4139,N_1516);
or U5684 (N_5684,N_41,N_4765);
nand U5685 (N_5685,N_1941,N_3569);
nor U5686 (N_5686,N_3224,N_3898);
and U5687 (N_5687,N_2485,N_3006);
and U5688 (N_5688,N_3655,N_1044);
nor U5689 (N_5689,N_1481,N_4508);
nand U5690 (N_5690,N_4739,N_2615);
and U5691 (N_5691,N_4577,N_2594);
or U5692 (N_5692,N_4123,N_257);
nor U5693 (N_5693,N_1360,N_4682);
nor U5694 (N_5694,N_4308,N_1695);
nand U5695 (N_5695,N_1177,N_2193);
nand U5696 (N_5696,N_4232,N_2286);
or U5697 (N_5697,N_4861,N_114);
and U5698 (N_5698,N_2949,N_4120);
xor U5699 (N_5699,N_3767,N_4855);
or U5700 (N_5700,N_3688,N_3010);
or U5701 (N_5701,N_4893,N_2107);
nor U5702 (N_5702,N_857,N_3004);
or U5703 (N_5703,N_1007,N_1294);
xor U5704 (N_5704,N_465,N_2437);
or U5705 (N_5705,N_331,N_47);
nor U5706 (N_5706,N_3891,N_1207);
and U5707 (N_5707,N_3779,N_3979);
nor U5708 (N_5708,N_3435,N_3023);
xnor U5709 (N_5709,N_4718,N_182);
nor U5710 (N_5710,N_3422,N_2746);
and U5711 (N_5711,N_4192,N_1078);
and U5712 (N_5712,N_2846,N_755);
and U5713 (N_5713,N_2513,N_1147);
nand U5714 (N_5714,N_511,N_1774);
or U5715 (N_5715,N_637,N_421);
or U5716 (N_5716,N_3936,N_3942);
nand U5717 (N_5717,N_1628,N_1162);
nand U5718 (N_5718,N_4039,N_4466);
nor U5719 (N_5719,N_3780,N_4667);
nand U5720 (N_5720,N_3658,N_3918);
and U5721 (N_5721,N_1390,N_2644);
xor U5722 (N_5722,N_3926,N_2887);
nand U5723 (N_5723,N_202,N_3253);
nand U5724 (N_5724,N_2745,N_417);
and U5725 (N_5725,N_1318,N_2955);
nor U5726 (N_5726,N_2995,N_1828);
or U5727 (N_5727,N_304,N_4502);
nor U5728 (N_5728,N_1347,N_3724);
or U5729 (N_5729,N_3341,N_3805);
and U5730 (N_5730,N_4320,N_2944);
or U5731 (N_5731,N_2547,N_918);
nand U5732 (N_5732,N_279,N_531);
nor U5733 (N_5733,N_362,N_3596);
or U5734 (N_5734,N_221,N_2484);
or U5735 (N_5735,N_3745,N_4271);
and U5736 (N_5736,N_461,N_397);
or U5737 (N_5737,N_3821,N_2571);
nand U5738 (N_5738,N_4603,N_1697);
nor U5739 (N_5739,N_907,N_3556);
or U5740 (N_5740,N_4865,N_1873);
nor U5741 (N_5741,N_2024,N_4617);
and U5742 (N_5742,N_2122,N_1654);
nor U5743 (N_5743,N_3965,N_1311);
nand U5744 (N_5744,N_1399,N_2631);
nor U5745 (N_5745,N_4102,N_4199);
nand U5746 (N_5746,N_1644,N_781);
or U5747 (N_5747,N_430,N_1051);
nand U5748 (N_5748,N_2199,N_1008);
and U5749 (N_5749,N_250,N_4000);
nor U5750 (N_5750,N_890,N_184);
nand U5751 (N_5751,N_2104,N_3350);
or U5752 (N_5752,N_2156,N_1224);
nand U5753 (N_5753,N_4231,N_2536);
nand U5754 (N_5754,N_2501,N_4544);
nand U5755 (N_5755,N_2184,N_161);
or U5756 (N_5756,N_718,N_4077);
nand U5757 (N_5757,N_4501,N_2795);
nand U5758 (N_5758,N_2966,N_2548);
nand U5759 (N_5759,N_4219,N_473);
or U5760 (N_5760,N_3179,N_3900);
nor U5761 (N_5761,N_2537,N_2345);
and U5762 (N_5762,N_565,N_1161);
nand U5763 (N_5763,N_1633,N_3438);
and U5764 (N_5764,N_2866,N_3938);
and U5765 (N_5765,N_3071,N_1819);
and U5766 (N_5766,N_3216,N_3480);
nand U5767 (N_5767,N_3968,N_3661);
or U5768 (N_5768,N_2761,N_4894);
nor U5769 (N_5769,N_2868,N_2490);
and U5770 (N_5770,N_2897,N_1298);
nor U5771 (N_5771,N_1269,N_1379);
nand U5772 (N_5772,N_1069,N_1701);
and U5773 (N_5773,N_3581,N_2900);
xor U5774 (N_5774,N_1184,N_2567);
or U5775 (N_5775,N_3462,N_335);
or U5776 (N_5776,N_3899,N_1102);
nor U5777 (N_5777,N_1858,N_2648);
and U5778 (N_5778,N_3133,N_786);
nand U5779 (N_5779,N_520,N_4712);
or U5780 (N_5780,N_2175,N_1515);
and U5781 (N_5781,N_4471,N_1928);
or U5782 (N_5782,N_4751,N_1696);
nand U5783 (N_5783,N_3601,N_3214);
and U5784 (N_5784,N_751,N_664);
nand U5785 (N_5785,N_4141,N_354);
nor U5786 (N_5786,N_1049,N_1576);
or U5787 (N_5787,N_1457,N_2423);
and U5788 (N_5788,N_4160,N_2638);
nor U5789 (N_5789,N_3870,N_4583);
or U5790 (N_5790,N_2780,N_401);
or U5791 (N_5791,N_4518,N_3223);
or U5792 (N_5792,N_3669,N_2609);
nand U5793 (N_5793,N_2480,N_2987);
and U5794 (N_5794,N_2247,N_2177);
and U5795 (N_5795,N_425,N_634);
or U5796 (N_5796,N_3292,N_705);
nor U5797 (N_5797,N_2575,N_24);
and U5798 (N_5798,N_2160,N_1713);
or U5799 (N_5799,N_432,N_4820);
xor U5800 (N_5800,N_2472,N_965);
xnor U5801 (N_5801,N_2438,N_4695);
and U5802 (N_5802,N_4516,N_2980);
xor U5803 (N_5803,N_1923,N_3106);
nor U5804 (N_5804,N_2684,N_239);
and U5805 (N_5805,N_3637,N_1146);
and U5806 (N_5806,N_3215,N_4658);
nand U5807 (N_5807,N_1195,N_1721);
nor U5808 (N_5808,N_478,N_695);
and U5809 (N_5809,N_2587,N_3406);
or U5810 (N_5810,N_1661,N_3925);
nor U5811 (N_5811,N_963,N_1131);
or U5812 (N_5812,N_3453,N_3861);
nand U5813 (N_5813,N_4482,N_2427);
nand U5814 (N_5814,N_1708,N_1988);
and U5815 (N_5815,N_2309,N_4972);
xor U5816 (N_5816,N_3975,N_1466);
and U5817 (N_5817,N_3762,N_4897);
nor U5818 (N_5818,N_1000,N_3405);
xor U5819 (N_5819,N_949,N_2670);
nor U5820 (N_5820,N_1098,N_3699);
and U5821 (N_5821,N_1831,N_756);
nand U5822 (N_5822,N_1734,N_2234);
or U5823 (N_5823,N_3700,N_78);
nand U5824 (N_5824,N_3484,N_1197);
and U5825 (N_5825,N_3418,N_317);
xor U5826 (N_5826,N_962,N_3040);
nor U5827 (N_5827,N_1393,N_414);
nand U5828 (N_5828,N_3213,N_1537);
nand U5829 (N_5829,N_649,N_4556);
or U5830 (N_5830,N_3495,N_1122);
nor U5831 (N_5831,N_4337,N_4002);
and U5832 (N_5832,N_3162,N_306);
and U5833 (N_5833,N_2733,N_313);
nand U5834 (N_5834,N_3322,N_2151);
and U5835 (N_5835,N_1300,N_2798);
and U5836 (N_5836,N_2305,N_4531);
nor U5837 (N_5837,N_2025,N_2508);
nand U5838 (N_5838,N_3859,N_3705);
nor U5839 (N_5839,N_427,N_2132);
and U5840 (N_5840,N_2776,N_244);
and U5841 (N_5841,N_4670,N_4701);
and U5842 (N_5842,N_4737,N_3944);
xnor U5843 (N_5843,N_3568,N_1254);
or U5844 (N_5844,N_3845,N_4890);
nor U5845 (N_5845,N_4188,N_3410);
or U5846 (N_5846,N_3896,N_2777);
xnor U5847 (N_5847,N_4249,N_1249);
nand U5848 (N_5848,N_4830,N_4361);
or U5849 (N_5849,N_4210,N_1026);
or U5850 (N_5850,N_2167,N_4480);
nand U5851 (N_5851,N_1666,N_3291);
nor U5852 (N_5852,N_2946,N_3065);
xor U5853 (N_5853,N_113,N_3540);
nor U5854 (N_5854,N_4477,N_4876);
or U5855 (N_5855,N_4648,N_3055);
and U5856 (N_5856,N_1665,N_1624);
or U5857 (N_5857,N_2002,N_3108);
and U5858 (N_5858,N_2248,N_4912);
or U5859 (N_5859,N_2591,N_2246);
or U5860 (N_5860,N_1287,N_3387);
and U5861 (N_5861,N_713,N_3910);
xor U5862 (N_5862,N_1528,N_39);
and U5863 (N_5863,N_546,N_3064);
nand U5864 (N_5864,N_3343,N_2928);
and U5865 (N_5865,N_2047,N_3141);
or U5866 (N_5866,N_288,N_1013);
xnor U5867 (N_5867,N_2854,N_3424);
nand U5868 (N_5868,N_2599,N_801);
nand U5869 (N_5869,N_1776,N_4179);
nor U5870 (N_5870,N_3001,N_4822);
or U5871 (N_5871,N_1389,N_553);
or U5872 (N_5872,N_1316,N_3890);
and U5873 (N_5873,N_3263,N_1961);
nand U5874 (N_5874,N_4523,N_2713);
nor U5875 (N_5875,N_1888,N_2996);
xor U5876 (N_5876,N_3377,N_1910);
nand U5877 (N_5877,N_1324,N_4568);
or U5878 (N_5878,N_4752,N_2231);
nand U5879 (N_5879,N_4318,N_628);
xnor U5880 (N_5880,N_4629,N_3773);
nor U5881 (N_5881,N_3380,N_2851);
or U5882 (N_5882,N_1977,N_3675);
nor U5883 (N_5883,N_670,N_2690);
nand U5884 (N_5884,N_2262,N_852);
nand U5885 (N_5885,N_4479,N_1253);
xnor U5886 (N_5886,N_1838,N_3966);
nor U5887 (N_5887,N_2185,N_550);
or U5888 (N_5888,N_3916,N_1094);
and U5889 (N_5889,N_783,N_1608);
and U5890 (N_5890,N_1114,N_830);
nand U5891 (N_5891,N_4829,N_2495);
xor U5892 (N_5892,N_3308,N_4447);
or U5893 (N_5893,N_3024,N_1757);
nand U5894 (N_5894,N_4349,N_106);
and U5895 (N_5895,N_3286,N_1768);
or U5896 (N_5896,N_1019,N_2302);
or U5897 (N_5897,N_2048,N_4799);
or U5898 (N_5898,N_4947,N_4054);
xnor U5899 (N_5899,N_3712,N_1363);
nand U5900 (N_5900,N_1440,N_780);
nor U5901 (N_5901,N_2574,N_3817);
nor U5902 (N_5902,N_2891,N_2462);
nand U5903 (N_5903,N_1881,N_4335);
xor U5904 (N_5904,N_4136,N_1134);
or U5905 (N_5905,N_1922,N_4124);
and U5906 (N_5906,N_981,N_697);
xnor U5907 (N_5907,N_449,N_3464);
or U5908 (N_5908,N_3735,N_4817);
or U5909 (N_5909,N_3839,N_4473);
or U5910 (N_5910,N_4707,N_889);
or U5911 (N_5911,N_1214,N_2064);
xnor U5912 (N_5912,N_1722,N_1063);
nor U5913 (N_5913,N_1551,N_208);
and U5914 (N_5914,N_1623,N_3619);
nor U5915 (N_5915,N_2527,N_2934);
xnor U5916 (N_5916,N_3137,N_958);
xor U5917 (N_5917,N_2165,N_2650);
nand U5918 (N_5918,N_1317,N_2431);
xor U5919 (N_5919,N_4578,N_4589);
xor U5920 (N_5920,N_409,N_587);
nor U5921 (N_5921,N_3172,N_2387);
nor U5922 (N_5922,N_3390,N_4363);
or U5923 (N_5923,N_687,N_2498);
or U5924 (N_5924,N_3885,N_296);
nand U5925 (N_5925,N_3838,N_3302);
nand U5926 (N_5926,N_799,N_735);
or U5927 (N_5927,N_2844,N_1402);
or U5928 (N_5928,N_4115,N_2109);
nand U5929 (N_5929,N_2346,N_1087);
nand U5930 (N_5930,N_3962,N_3012);
and U5931 (N_5931,N_1124,N_3523);
and U5932 (N_5932,N_1869,N_2826);
nor U5933 (N_5933,N_4298,N_2993);
or U5934 (N_5934,N_2766,N_1969);
and U5935 (N_5935,N_1987,N_2872);
or U5936 (N_5936,N_3534,N_3657);
or U5937 (N_5937,N_987,N_1865);
nand U5938 (N_5938,N_4412,N_2242);
nor U5939 (N_5939,N_2753,N_921);
or U5940 (N_5940,N_4056,N_4552);
or U5941 (N_5941,N_4461,N_4126);
xor U5942 (N_5942,N_826,N_1109);
and U5943 (N_5943,N_308,N_3889);
nand U5944 (N_5944,N_1971,N_4411);
xnor U5945 (N_5945,N_1243,N_2039);
or U5946 (N_5946,N_888,N_3425);
and U5947 (N_5947,N_1116,N_4418);
xor U5948 (N_5948,N_3627,N_2924);
nor U5949 (N_5949,N_242,N_3760);
and U5950 (N_5950,N_2460,N_3904);
nand U5951 (N_5951,N_2415,N_2392);
nor U5952 (N_5952,N_3527,N_1980);
nor U5953 (N_5953,N_2925,N_383);
or U5954 (N_5954,N_4193,N_4223);
or U5955 (N_5955,N_4910,N_2886);
and U5956 (N_5956,N_1866,N_1421);
and U5957 (N_5957,N_1738,N_4111);
or U5958 (N_5958,N_4868,N_1088);
or U5959 (N_5959,N_4057,N_3190);
and U5960 (N_5960,N_4626,N_2034);
nand U5961 (N_5961,N_1220,N_4511);
nand U5962 (N_5962,N_1787,N_945);
or U5963 (N_5963,N_3666,N_3983);
xor U5964 (N_5964,N_1802,N_3555);
nand U5965 (N_5965,N_4313,N_3056);
nand U5966 (N_5966,N_3474,N_4680);
nand U5967 (N_5967,N_3051,N_4515);
or U5968 (N_5968,N_2992,N_2882);
or U5969 (N_5969,N_2394,N_636);
nand U5970 (N_5970,N_71,N_1619);
and U5971 (N_5971,N_4687,N_2192);
nand U5972 (N_5972,N_573,N_2911);
xor U5973 (N_5973,N_4404,N_1479);
nand U5974 (N_5974,N_1451,N_2890);
nor U5975 (N_5975,N_2836,N_1545);
nor U5976 (N_5976,N_4441,N_3624);
and U5977 (N_5977,N_762,N_2099);
nor U5978 (N_5978,N_827,N_523);
or U5979 (N_5979,N_1062,N_3920);
and U5980 (N_5980,N_361,N_19);
nand U5981 (N_5981,N_3616,N_822);
or U5982 (N_5982,N_129,N_4908);
nor U5983 (N_5983,N_3384,N_1239);
or U5984 (N_5984,N_2315,N_433);
or U5985 (N_5985,N_4826,N_1898);
or U5986 (N_5986,N_4386,N_4614);
nand U5987 (N_5987,N_3785,N_1040);
or U5988 (N_5988,N_1492,N_1999);
and U5989 (N_5989,N_53,N_585);
nor U5990 (N_5990,N_474,N_2216);
nor U5991 (N_5991,N_4283,N_2379);
nor U5992 (N_5992,N_2596,N_667);
nand U5993 (N_5993,N_1405,N_1743);
or U5994 (N_5994,N_554,N_3027);
nor U5995 (N_5995,N_4167,N_4060);
and U5996 (N_5996,N_495,N_1123);
nor U5997 (N_5997,N_3500,N_2408);
nand U5998 (N_5998,N_4368,N_1609);
nand U5999 (N_5999,N_1429,N_2036);
nor U6000 (N_6000,N_2804,N_3906);
nand U6001 (N_6001,N_3296,N_4653);
nor U6002 (N_6002,N_3854,N_2708);
or U6003 (N_6003,N_1662,N_147);
or U6004 (N_6004,N_773,N_2016);
and U6005 (N_6005,N_2040,N_2614);
nand U6006 (N_6006,N_4660,N_2499);
and U6007 (N_6007,N_91,N_3994);
xnor U6008 (N_6008,N_3471,N_4862);
nor U6009 (N_6009,N_2313,N_4006);
or U6010 (N_6010,N_3477,N_405);
nand U6011 (N_6011,N_3486,N_4326);
nor U6012 (N_6012,N_1691,N_3076);
or U6013 (N_6013,N_782,N_2859);
nor U6014 (N_6014,N_3128,N_4998);
or U6015 (N_6015,N_2731,N_3525);
nor U6016 (N_6016,N_4468,N_1121);
and U6017 (N_6017,N_3660,N_4926);
nand U6018 (N_6018,N_2636,N_90);
nor U6019 (N_6019,N_597,N_567);
and U6020 (N_6020,N_2699,N_2217);
and U6021 (N_6021,N_2268,N_25);
nand U6022 (N_6022,N_4635,N_1905);
xor U6023 (N_6023,N_1413,N_3383);
nor U6024 (N_6024,N_552,N_2945);
nand U6025 (N_6025,N_4560,N_332);
or U6026 (N_6026,N_3611,N_3068);
nand U6027 (N_6027,N_1200,N_1855);
or U6028 (N_6028,N_856,N_138);
and U6029 (N_6029,N_4070,N_4620);
and U6030 (N_6030,N_3046,N_1264);
nand U6031 (N_6031,N_153,N_1133);
nor U6032 (N_6032,N_3271,N_1771);
nor U6033 (N_6033,N_2991,N_916);
or U6034 (N_6034,N_3609,N_4260);
and U6035 (N_6035,N_845,N_2092);
nand U6036 (N_6036,N_2200,N_808);
nor U6037 (N_6037,N_128,N_3993);
nand U6038 (N_6038,N_4647,N_3144);
nand U6039 (N_6039,N_3107,N_622);
and U6040 (N_6040,N_2807,N_3988);
or U6041 (N_6041,N_264,N_2719);
and U6042 (N_6042,N_2660,N_4557);
nor U6043 (N_6043,N_3600,N_4158);
nand U6044 (N_6044,N_3221,N_1125);
xor U6045 (N_6045,N_3142,N_2661);
nand U6046 (N_6046,N_1009,N_2705);
and U6047 (N_6047,N_2312,N_512);
xor U6048 (N_6048,N_1256,N_4838);
nor U6049 (N_6049,N_3400,N_941);
and U6050 (N_6050,N_1105,N_4863);
nor U6051 (N_6051,N_4268,N_1255);
or U6052 (N_6052,N_1307,N_3563);
nor U6053 (N_6053,N_737,N_2182);
nor U6054 (N_6054,N_2981,N_2902);
xnor U6055 (N_6055,N_500,N_3716);
nand U6056 (N_6056,N_3008,N_2393);
xnor U6057 (N_6057,N_1079,N_3299);
xor U6058 (N_6058,N_4993,N_292);
nor U6059 (N_6059,N_2557,N_2962);
nand U6060 (N_6060,N_2554,N_280);
xnor U6061 (N_6061,N_1091,N_4587);
nand U6062 (N_6062,N_2071,N_349);
or U6063 (N_6063,N_4293,N_701);
or U6064 (N_6064,N_4990,N_1602);
nor U6065 (N_6065,N_1059,N_4443);
or U6066 (N_6066,N_1473,N_4740);
nand U6067 (N_6067,N_3719,N_192);
or U6068 (N_6068,N_3049,N_3931);
and U6069 (N_6069,N_1603,N_1749);
nand U6070 (N_6070,N_4035,N_116);
or U6071 (N_6071,N_4999,N_3354);
and U6072 (N_6072,N_2174,N_4109);
and U6073 (N_6073,N_3526,N_4857);
and U6074 (N_6074,N_4769,N_1331);
nor U6075 (N_6075,N_4600,N_568);
nor U6076 (N_6076,N_1824,N_319);
nand U6077 (N_6077,N_4380,N_809);
and U6078 (N_6078,N_2651,N_4566);
or U6079 (N_6079,N_3225,N_2810);
or U6080 (N_6080,N_711,N_719);
nand U6081 (N_6081,N_1050,N_373);
xnor U6082 (N_6082,N_4490,N_4689);
and U6083 (N_6083,N_3640,N_201);
nor U6084 (N_6084,N_3770,N_1362);
or U6085 (N_6085,N_891,N_2203);
nor U6086 (N_6086,N_246,N_2789);
nor U6087 (N_6087,N_2434,N_3326);
and U6088 (N_6088,N_2756,N_1341);
and U6089 (N_6089,N_2487,N_2023);
nor U6090 (N_6090,N_3862,N_4346);
or U6091 (N_6091,N_2938,N_2001);
or U6092 (N_6092,N_3922,N_2218);
nor U6093 (N_6093,N_4027,N_2400);
or U6094 (N_6094,N_3754,N_4487);
nand U6095 (N_6095,N_3290,N_4934);
or U6096 (N_6096,N_4137,N_3115);
or U6097 (N_6097,N_4792,N_2654);
nor U6098 (N_6098,N_3740,N_2325);
and U6099 (N_6099,N_4348,N_52);
xor U6100 (N_6100,N_3588,N_4627);
nand U6101 (N_6101,N_1099,N_1303);
nand U6102 (N_6102,N_3439,N_2469);
nand U6103 (N_6103,N_2558,N_641);
and U6104 (N_6104,N_1221,N_3630);
and U6105 (N_6105,N_4722,N_1165);
nand U6106 (N_6106,N_3371,N_3120);
nand U6107 (N_6107,N_363,N_618);
xor U6108 (N_6108,N_3731,N_1395);
and U6109 (N_6109,N_3416,N_1785);
and U6110 (N_6110,N_3970,N_984);
and U6111 (N_6111,N_902,N_4987);
and U6112 (N_6112,N_3070,N_4883);
xor U6113 (N_6113,N_2391,N_1669);
or U6114 (N_6114,N_3872,N_4979);
and U6115 (N_6115,N_1935,N_2620);
nor U6116 (N_6116,N_4885,N_656);
xor U6117 (N_6117,N_1765,N_4944);
or U6118 (N_6118,N_1015,N_3396);
or U6119 (N_6119,N_1148,N_988);
nor U6120 (N_6120,N_4229,N_4694);
nor U6121 (N_6121,N_4470,N_1973);
or U6122 (N_6122,N_3543,N_4226);
and U6123 (N_6123,N_1951,N_3811);
or U6124 (N_6124,N_4753,N_594);
nand U6125 (N_6125,N_3493,N_4584);
or U6126 (N_6126,N_2371,N_932);
nor U6127 (N_6127,N_3457,N_3073);
or U6128 (N_6128,N_3321,N_4512);
nor U6129 (N_6129,N_4140,N_3061);
or U6130 (N_6130,N_761,N_1204);
nand U6131 (N_6131,N_3544,N_624);
and U6132 (N_6132,N_214,N_1004);
and U6133 (N_6133,N_4084,N_4915);
or U6134 (N_6134,N_3864,N_2055);
and U6135 (N_6135,N_4117,N_1505);
nand U6136 (N_6136,N_2173,N_4370);
nand U6137 (N_6137,N_4553,N_2306);
or U6138 (N_6138,N_3494,N_1361);
or U6139 (N_6139,N_2714,N_4942);
or U6140 (N_6140,N_4731,N_972);
nor U6141 (N_6141,N_37,N_3837);
nor U6142 (N_6142,N_3615,N_2178);
nor U6143 (N_6143,N_3803,N_379);
nand U6144 (N_6144,N_3324,N_839);
nor U6145 (N_6145,N_4957,N_1967);
nand U6146 (N_6146,N_1272,N_4419);
nand U6147 (N_6147,N_3294,N_498);
and U6148 (N_6148,N_3621,N_2332);
xnor U6149 (N_6149,N_4251,N_763);
and U6150 (N_6150,N_3235,N_3687);
nor U6151 (N_6151,N_102,N_3971);
xnor U6152 (N_6152,N_4063,N_1635);
nand U6153 (N_6153,N_671,N_652);
or U6154 (N_6154,N_3095,N_4247);
and U6155 (N_6155,N_4347,N_1792);
nand U6156 (N_6156,N_73,N_3148);
nor U6157 (N_6157,N_4907,N_2294);
and U6158 (N_6158,N_1658,N_3370);
or U6159 (N_6159,N_3038,N_154);
nor U6160 (N_6160,N_1422,N_3633);
nor U6161 (N_6161,N_1889,N_4342);
nor U6162 (N_6162,N_4273,N_117);
nand U6163 (N_6163,N_814,N_4465);
nor U6164 (N_6164,N_1182,N_166);
xor U6165 (N_6165,N_1445,N_871);
xor U6166 (N_6166,N_2075,N_318);
or U6167 (N_6167,N_139,N_3789);
nor U6168 (N_6168,N_2675,N_2629);
and U6169 (N_6169,N_4252,N_2883);
or U6170 (N_6170,N_1647,N_294);
nand U6171 (N_6171,N_1215,N_2421);
or U6172 (N_6172,N_4020,N_486);
nor U6173 (N_6173,N_603,N_4618);
and U6174 (N_6174,N_215,N_2582);
or U6175 (N_6175,N_4078,N_1675);
and U6176 (N_6176,N_679,N_479);
nand U6177 (N_6177,N_3159,N_258);
and U6178 (N_6178,N_4564,N_3470);
and U6179 (N_6179,N_3232,N_4087);
or U6180 (N_6180,N_2841,N_4007);
or U6181 (N_6181,N_1543,N_75);
nor U6182 (N_6182,N_4030,N_4287);
nor U6183 (N_6183,N_3498,N_1448);
nor U6184 (N_6184,N_4759,N_1890);
or U6185 (N_6185,N_551,N_3298);
and U6186 (N_6186,N_4738,N_224);
and U6187 (N_6187,N_4220,N_1611);
nor U6188 (N_6188,N_2762,N_1385);
or U6189 (N_6189,N_3423,N_3584);
xor U6190 (N_6190,N_566,N_4059);
or U6191 (N_6191,N_1242,N_684);
or U6192 (N_6192,N_4445,N_2757);
nor U6193 (N_6193,N_125,N_4301);
nand U6194 (N_6194,N_4843,N_268);
and U6195 (N_6195,N_457,N_4267);
and U6196 (N_6196,N_3937,N_1686);
nor U6197 (N_6197,N_4657,N_109);
and U6198 (N_6198,N_785,N_3636);
or U6199 (N_6199,N_3855,N_3231);
nor U6200 (N_6200,N_803,N_2333);
nand U6201 (N_6201,N_3411,N_233);
nand U6202 (N_6202,N_1939,N_847);
nand U6203 (N_6203,N_164,N_1825);
nor U6204 (N_6204,N_1916,N_1538);
nand U6205 (N_6205,N_1344,N_1983);
xnor U6206 (N_6206,N_975,N_4757);
and U6207 (N_6207,N_4777,N_4274);
nor U6208 (N_6208,N_562,N_3114);
and U6209 (N_6209,N_4685,N_3147);
and U6210 (N_6210,N_1685,N_4723);
and U6211 (N_6211,N_1056,N_959);
nand U6212 (N_6212,N_2796,N_2475);
or U6213 (N_6213,N_269,N_4315);
or U6214 (N_6214,N_4261,N_4495);
and U6215 (N_6215,N_2145,N_4805);
or U6216 (N_6216,N_1232,N_3490);
and U6217 (N_6217,N_2957,N_46);
or U6218 (N_6218,N_3608,N_4943);
nor U6219 (N_6219,N_4570,N_2521);
nor U6220 (N_6220,N_2592,N_2834);
xnor U6221 (N_6221,N_2979,N_3255);
and U6222 (N_6222,N_1155,N_4176);
nor U6223 (N_6223,N_1006,N_1788);
and U6224 (N_6224,N_561,N_360);
or U6225 (N_6225,N_2337,N_1563);
nor U6226 (N_6226,N_100,N_3328);
xnor U6227 (N_6227,N_4732,N_2135);
nor U6228 (N_6228,N_4023,N_805);
and U6229 (N_6229,N_1532,N_1176);
nor U6230 (N_6230,N_3171,N_2307);
nand U6231 (N_6231,N_458,N_1278);
nor U6232 (N_6232,N_4615,N_1297);
and U6233 (N_6233,N_1511,N_3014);
and U6234 (N_6234,N_358,N_3082);
and U6235 (N_6235,N_659,N_3117);
xor U6236 (N_6236,N_4542,N_1038);
and U6237 (N_6237,N_1323,N_1426);
and U6238 (N_6238,N_63,N_2059);
xnor U6239 (N_6239,N_1431,N_3209);
and U6240 (N_6240,N_1442,N_87);
or U6241 (N_6241,N_753,N_151);
and U6242 (N_6242,N_3408,N_3681);
and U6243 (N_6243,N_424,N_86);
xnor U6244 (N_6244,N_1892,N_394);
nand U6245 (N_6245,N_3456,N_1181);
nand U6246 (N_6246,N_435,N_683);
nand U6247 (N_6247,N_4672,N_451);
or U6248 (N_6248,N_3641,N_4197);
nor U6249 (N_6249,N_4665,N_2514);
nor U6250 (N_6250,N_4157,N_3617);
nor U6251 (N_6251,N_2382,N_4010);
nand U6252 (N_6252,N_800,N_4439);
nand U6253 (N_6253,N_772,N_2459);
and U6254 (N_6254,N_4684,N_908);
nor U6255 (N_6255,N_3276,N_1014);
nor U6256 (N_6256,N_1206,N_2538);
nor U6257 (N_6257,N_4,N_3155);
and U6258 (N_6258,N_28,N_3887);
nand U6259 (N_6259,N_1965,N_3087);
and U6260 (N_6260,N_2937,N_455);
and U6261 (N_6261,N_4080,N_1420);
and U6262 (N_6262,N_4282,N_1940);
nor U6263 (N_6263,N_1397,N_3099);
or U6264 (N_6264,N_4409,N_286);
and U6265 (N_6265,N_1135,N_34);
or U6266 (N_6266,N_4429,N_3510);
xor U6267 (N_6267,N_302,N_2808);
and U6268 (N_6268,N_1115,N_3537);
xnor U6269 (N_6269,N_3025,N_1443);
nor U6270 (N_6270,N_2975,N_1064);
nand U6271 (N_6271,N_2204,N_1486);
nor U6272 (N_6272,N_3333,N_917);
nor U6273 (N_6273,N_3472,N_3991);
and U6274 (N_6274,N_2189,N_2956);
nand U6275 (N_6275,N_3197,N_1650);
and U6276 (N_6276,N_2794,N_3507);
and U6277 (N_6277,N_824,N_2147);
xnor U6278 (N_6278,N_4092,N_1275);
nor U6279 (N_6279,N_193,N_4674);
nor U6280 (N_6280,N_4181,N_1887);
or U6281 (N_6281,N_1681,N_4090);
xor U6282 (N_6282,N_2819,N_3169);
nand U6283 (N_6283,N_3264,N_4350);
nor U6284 (N_6284,N_1756,N_4204);
and U6285 (N_6285,N_3181,N_3955);
or U6286 (N_6286,N_4887,N_43);
or U6287 (N_6287,N_1250,N_134);
xnor U6288 (N_6288,N_815,N_1689);
and U6289 (N_6289,N_3783,N_1570);
or U6290 (N_6290,N_2363,N_3509);
nor U6291 (N_6291,N_1632,N_4264);
xnor U6292 (N_6292,N_26,N_1502);
nand U6293 (N_6293,N_1500,N_4250);
nand U6294 (N_6294,N_3800,N_2626);
xnor U6295 (N_6295,N_2827,N_3448);
and U6296 (N_6296,N_3879,N_4851);
nor U6297 (N_6297,N_2503,N_1613);
xor U6298 (N_6298,N_2385,N_420);
nand U6299 (N_6299,N_3479,N_3243);
xor U6300 (N_6300,N_2241,N_1071);
or U6301 (N_6301,N_1285,N_305);
and U6302 (N_6302,N_2821,N_1549);
nand U6303 (N_6303,N_4228,N_1801);
nand U6304 (N_6304,N_668,N_2577);
nor U6305 (N_6305,N_2118,N_4001);
nand U6306 (N_6306,N_999,N_3508);
nor U6307 (N_6307,N_848,N_1251);
and U6308 (N_6308,N_402,N_1845);
xnor U6309 (N_6309,N_1118,N_1352);
xor U6310 (N_6310,N_4352,N_1219);
nand U6311 (N_6311,N_2279,N_4201);
nor U6312 (N_6312,N_788,N_4519);
nor U6313 (N_6313,N_1446,N_271);
nor U6314 (N_6314,N_2374,N_3823);
or U6315 (N_6315,N_741,N_338);
and U6316 (N_6316,N_4664,N_2196);
nor U6317 (N_6317,N_2977,N_1375);
or U6318 (N_6318,N_4244,N_2811);
and U6319 (N_6319,N_1746,N_2186);
and U6320 (N_6320,N_4541,N_1328);
nor U6321 (N_6321,N_3005,N_3413);
and U6322 (N_6322,N_472,N_2335);
or U6323 (N_6323,N_4364,N_1642);
nor U6324 (N_6324,N_4533,N_1231);
or U6325 (N_6325,N_864,N_2931);
or U6326 (N_6326,N_3404,N_3539);
and U6327 (N_6327,N_422,N_1634);
or U6328 (N_6328,N_11,N_4304);
and U6329 (N_6329,N_3836,N_3622);
xor U6330 (N_6330,N_3514,N_1783);
or U6331 (N_6331,N_1045,N_1546);
and U6332 (N_6332,N_2425,N_3160);
and U6333 (N_6333,N_55,N_1510);
nor U6334 (N_6334,N_2277,N_1153);
or U6335 (N_6335,N_3711,N_1933);
nor U6336 (N_6336,N_709,N_3281);
or U6337 (N_6337,N_4588,N_4414);
nor U6338 (N_6338,N_263,N_882);
and U6339 (N_6339,N_3100,N_4954);
nand U6340 (N_6340,N_158,N_4442);
nor U6341 (N_6341,N_3039,N_2418);
nand U6342 (N_6342,N_3788,N_982);
or U6343 (N_6343,N_388,N_1610);
xnor U6344 (N_6344,N_3303,N_4500);
nor U6345 (N_6345,N_1478,N_497);
or U6346 (N_6346,N_3853,N_1534);
xor U6347 (N_6347,N_2271,N_2572);
nor U6348 (N_6348,N_3741,N_1741);
and U6349 (N_6349,N_1370,N_1035);
nor U6350 (N_6350,N_650,N_395);
nor U6351 (N_6351,N_1762,N_4686);
or U6352 (N_6352,N_2694,N_901);
or U6353 (N_6353,N_4256,N_4170);
and U6354 (N_6354,N_2500,N_206);
xnor U6355 (N_6355,N_1199,N_4166);
nand U6356 (N_6356,N_2270,N_3765);
nor U6357 (N_6357,N_2656,N_4103);
xor U6358 (N_6358,N_4836,N_2604);
nor U6359 (N_6359,N_4679,N_1524);
nor U6360 (N_6360,N_1835,N_1573);
or U6361 (N_6361,N_84,N_4903);
or U6362 (N_6362,N_3786,N_2022);
nor U6363 (N_6363,N_4621,N_977);
and U6364 (N_6364,N_2797,N_115);
and U6365 (N_6365,N_3447,N_1718);
and U6366 (N_6366,N_3564,N_1235);
and U6367 (N_6367,N_3227,N_2110);
nand U6368 (N_6368,N_3647,N_928);
xor U6369 (N_6369,N_2687,N_2958);
nand U6370 (N_6370,N_3733,N_1784);
nor U6371 (N_6371,N_2863,N_4218);
nor U6372 (N_6372,N_3668,N_510);
xnor U6373 (N_6373,N_899,N_272);
and U6374 (N_6374,N_1850,N_4216);
and U6375 (N_6375,N_816,N_2833);
nor U6376 (N_6376,N_4514,N_3228);
nor U6377 (N_6377,N_83,N_4576);
nand U6378 (N_6378,N_410,N_3335);
nand U6379 (N_6379,N_2009,N_1726);
or U6380 (N_6380,N_4189,N_2202);
nand U6381 (N_6381,N_4844,N_1493);
or U6382 (N_6382,N_1427,N_301);
or U6383 (N_6383,N_3538,N_4047);
xnor U6384 (N_6384,N_3085,N_4211);
nand U6385 (N_6385,N_1208,N_4162);
or U6386 (N_6386,N_2267,N_3825);
and U6387 (N_6387,N_2176,N_4801);
or U6388 (N_6388,N_170,N_2007);
nor U6389 (N_6389,N_1920,N_67);
or U6390 (N_6390,N_1459,N_2205);
and U6391 (N_6391,N_1864,N_2507);
nor U6392 (N_6392,N_558,N_4449);
or U6393 (N_6393,N_1962,N_2070);
nand U6394 (N_6394,N_336,N_1498);
or U6395 (N_6395,N_4048,N_2439);
nand U6396 (N_6396,N_1773,N_1157);
nor U6397 (N_6397,N_3043,N_60);
or U6398 (N_6398,N_1189,N_1410);
and U6399 (N_6399,N_1929,N_1463);
and U6400 (N_6400,N_4510,N_2411);
xnor U6401 (N_6401,N_4432,N_3351);
or U6402 (N_6402,N_3815,N_3959);
and U6403 (N_6403,N_2227,N_2504);
nor U6404 (N_6404,N_4475,N_3610);
or U6405 (N_6405,N_2068,N_2380);
xor U6406 (N_6406,N_4387,N_1560);
nand U6407 (N_6407,N_2965,N_1861);
or U6408 (N_6408,N_4297,N_3728);
or U6409 (N_6409,N_436,N_2649);
nand U6410 (N_6410,N_2885,N_4807);
nor U6411 (N_6411,N_1425,N_1168);
and U6412 (N_6412,N_1110,N_3066);
and U6413 (N_6413,N_838,N_922);
nand U6414 (N_6414,N_3613,N_1918);
nand U6415 (N_6415,N_4535,N_1503);
nor U6416 (N_6416,N_1637,N_4748);
or U6417 (N_6417,N_398,N_1244);
nand U6418 (N_6418,N_2813,N_4272);
or U6419 (N_6419,N_3332,N_3759);
nand U6420 (N_6420,N_3603,N_3124);
nand U6421 (N_6421,N_4978,N_693);
nor U6422 (N_6422,N_4873,N_33);
nand U6423 (N_6423,N_4169,N_2935);
nand U6424 (N_6424,N_3734,N_893);
and U6425 (N_6425,N_293,N_2988);
and U6426 (N_6426,N_4241,N_2839);
and U6427 (N_6427,N_4072,N_1588);
nand U6428 (N_6428,N_3685,N_2864);
xor U6429 (N_6429,N_4714,N_3376);
nor U6430 (N_6430,N_4693,N_1688);
nor U6431 (N_6431,N_1985,N_4733);
nor U6432 (N_6432,N_2042,N_3443);
and U6433 (N_6433,N_1618,N_97);
nor U6434 (N_6434,N_1663,N_4547);
or U6435 (N_6435,N_440,N_4336);
or U6436 (N_6436,N_3244,N_4775);
and U6437 (N_6437,N_1046,N_4302);
xor U6438 (N_6438,N_2647,N_4842);
xnor U6439 (N_6439,N_820,N_3739);
nor U6440 (N_6440,N_4754,N_2770);
or U6441 (N_6441,N_3459,N_4948);
and U6442 (N_6442,N_2960,N_1540);
nand U6443 (N_6443,N_3002,N_477);
or U6444 (N_6444,N_1203,N_156);
nand U6445 (N_6445,N_2276,N_4450);
nor U6446 (N_6446,N_2085,N_4967);
nor U6447 (N_6447,N_2365,N_4839);
nand U6448 (N_6448,N_3268,N_4016);
nor U6449 (N_6449,N_3575,N_2274);
nand U6450 (N_6450,N_2259,N_506);
nand U6451 (N_6451,N_484,N_3348);
nor U6452 (N_6452,N_2559,N_3237);
or U6453 (N_6453,N_4266,N_4892);
and U6454 (N_6454,N_1683,N_254);
nor U6455 (N_6455,N_4580,N_2737);
nand U6456 (N_6456,N_2951,N_3729);
xnor U6457 (N_6457,N_4936,N_2212);
nor U6458 (N_6458,N_3282,N_4146);
xnor U6459 (N_6459,N_3782,N_548);
nor U6460 (N_6460,N_2849,N_3178);
nand U6461 (N_6461,N_3974,N_2329);
or U6462 (N_6462,N_2349,N_2076);
nand U6463 (N_6463,N_172,N_1997);
or U6464 (N_6464,N_4933,N_4476);
nand U6465 (N_6465,N_1789,N_1290);
nor U6466 (N_6466,N_3592,N_3997);
nor U6467 (N_6467,N_828,N_197);
or U6468 (N_6468,N_1309,N_3694);
nor U6469 (N_6469,N_2907,N_4233);
and U6470 (N_6470,N_3357,N_3431);
nand U6471 (N_6471,N_126,N_1353);
and U6472 (N_6472,N_2658,N_1192);
and U6473 (N_6473,N_2606,N_2818);
nor U6474 (N_6474,N_3288,N_3792);
nand U6475 (N_6475,N_1246,N_4572);
nand U6476 (N_6476,N_1636,N_615);
nor U6477 (N_6477,N_314,N_3113);
xnor U6478 (N_6478,N_2049,N_1684);
nor U6479 (N_6479,N_4376,N_678);
nor U6480 (N_6480,N_1350,N_81);
nand U6481 (N_6481,N_4608,N_3798);
nor U6482 (N_6482,N_4774,N_4891);
nor U6483 (N_6483,N_3996,N_108);
or U6484 (N_6484,N_2257,N_925);
and U6485 (N_6485,N_790,N_3589);
and U6486 (N_6486,N_4677,N_2552);
nor U6487 (N_6487,N_3487,N_2464);
xnor U6488 (N_6488,N_3801,N_3168);
nor U6489 (N_6489,N_3327,N_4378);
nand U6490 (N_6490,N_1600,N_3347);
and U6491 (N_6491,N_369,N_2835);
nand U6492 (N_6492,N_4003,N_4098);
or U6493 (N_6493,N_1834,N_1795);
xnor U6494 (N_6494,N_3360,N_2758);
nor U6495 (N_6495,N_4991,N_3909);
nor U6496 (N_6496,N_660,N_1154);
or U6497 (N_6497,N_4235,N_3915);
and U6498 (N_6498,N_1380,N_283);
or U6499 (N_6499,N_3125,N_1854);
nor U6500 (N_6500,N_4328,N_4406);
or U6501 (N_6501,N_94,N_396);
and U6502 (N_6502,N_4628,N_4815);
or U6503 (N_6503,N_1893,N_4906);
or U6504 (N_6504,N_4856,N_3730);
nand U6505 (N_6505,N_505,N_4569);
and U6506 (N_6506,N_3777,N_1268);
nor U6507 (N_6507,N_7,N_4869);
or U6508 (N_6508,N_4981,N_1963);
and U6509 (N_6509,N_525,N_4066);
or U6510 (N_6510,N_1769,N_730);
nor U6511 (N_6511,N_1521,N_1172);
nor U6512 (N_6512,N_3548,N_2936);
and U6513 (N_6513,N_2051,N_2254);
or U6514 (N_6514,N_577,N_4333);
or U6515 (N_6515,N_2927,N_2386);
nand U6516 (N_6516,N_4859,N_169);
nor U6517 (N_6517,N_4619,N_990);
or U6518 (N_6518,N_1504,N_837);
nand U6519 (N_6519,N_2524,N_3841);
and U6520 (N_6520,N_439,N_2046);
nand U6521 (N_6521,N_3638,N_4212);
nor U6522 (N_6522,N_3822,N_3840);
and U6523 (N_6523,N_4324,N_3469);
or U6524 (N_6524,N_1345,N_2790);
or U6525 (N_6525,N_2573,N_591);
or U6526 (N_6526,N_579,N_2781);
nor U6527 (N_6527,N_3031,N_2397);
and U6528 (N_6528,N_3430,N_3679);
nand U6529 (N_6529,N_3645,N_4114);
nand U6530 (N_6530,N_2324,N_3982);
xor U6531 (N_6531,N_323,N_4622);
nand U6532 (N_6532,N_4691,N_1080);
nand U6533 (N_6533,N_1885,N_3512);
and U6534 (N_6534,N_1621,N_3245);
and U6535 (N_6535,N_3483,N_1067);
or U6536 (N_6536,N_1070,N_3935);
or U6537 (N_6537,N_2143,N_4638);
nor U6538 (N_6538,N_961,N_411);
and U6539 (N_6539,N_1104,N_1883);
and U6540 (N_6540,N_2516,N_1981);
or U6541 (N_6541,N_825,N_4730);
and U6542 (N_6542,N_3297,N_4180);
nor U6543 (N_6543,N_4332,N_2355);
nand U6544 (N_6544,N_4257,N_2123);
or U6545 (N_6545,N_1700,N_3566);
and U6546 (N_6546,N_3883,N_1859);
nor U6547 (N_6547,N_1453,N_1979);
and U6548 (N_6548,N_953,N_4118);
nand U6549 (N_6549,N_77,N_2876);
nand U6550 (N_6550,N_1735,N_1760);
nor U6551 (N_6551,N_2466,N_3252);
and U6552 (N_6552,N_823,N_4486);
nand U6553 (N_6553,N_2115,N_1299);
and U6554 (N_6554,N_4288,N_3659);
nor U6555 (N_6555,N_3951,N_1612);
nor U6556 (N_6556,N_4489,N_3167);
and U6557 (N_6557,N_3419,N_3929);
xnor U6558 (N_6558,N_2595,N_3819);
or U6559 (N_6559,N_1444,N_3265);
nand U6560 (N_6560,N_1906,N_4952);
xnor U6561 (N_6561,N_2506,N_2409);
nor U6562 (N_6562,N_2997,N_2741);
and U6563 (N_6563,N_1127,N_2918);
and U6564 (N_6564,N_1404,N_14);
nand U6565 (N_6565,N_4071,N_940);
nand U6566 (N_6566,N_3119,N_3109);
or U6567 (N_6567,N_1754,N_3057);
nor U6568 (N_6568,N_589,N_101);
xor U6569 (N_6569,N_3515,N_4221);
nor U6570 (N_6570,N_4963,N_4191);
nor U6571 (N_6571,N_1703,N_1777);
nand U6572 (N_6572,N_4616,N_661);
and U6573 (N_6573,N_4481,N_2015);
and U6574 (N_6574,N_1737,N_3212);
or U6575 (N_6575,N_2347,N_266);
and U6576 (N_6576,N_2053,N_3301);
or U6577 (N_6577,N_3505,N_2362);
xor U6578 (N_6578,N_1593,N_663);
and U6579 (N_6579,N_2428,N_4309);
or U6580 (N_6580,N_4025,N_1531);
nand U6581 (N_6581,N_1811,N_316);
nor U6582 (N_6582,N_1274,N_2299);
and U6583 (N_6583,N_2710,N_4383);
or U6584 (N_6584,N_616,N_1433);
or U6585 (N_6585,N_1948,N_3522);
nand U6586 (N_6586,N_503,N_355);
nand U6587 (N_6587,N_3932,N_3203);
or U6588 (N_6588,N_522,N_2764);
nor U6589 (N_6589,N_4538,N_910);
or U6590 (N_6590,N_4540,N_612);
nor U6591 (N_6591,N_3559,N_1584);
nand U6592 (N_6592,N_1555,N_4036);
nor U6593 (N_6593,N_4696,N_3529);
nand U6594 (N_6594,N_2284,N_2353);
and U6595 (N_6595,N_1416,N_1751);
nor U6596 (N_6596,N_919,N_3035);
nand U6597 (N_6597,N_1495,N_4688);
and U6598 (N_6598,N_2515,N_4575);
nor U6599 (N_6599,N_1649,N_1209);
nand U6600 (N_6600,N_1068,N_2065);
xor U6601 (N_6601,N_692,N_833);
nand U6602 (N_6602,N_4424,N_2912);
nor U6603 (N_6603,N_4702,N_1895);
or U6604 (N_6604,N_572,N_617);
nand U6605 (N_6605,N_630,N_4536);
xnor U6606 (N_6606,N_2539,N_2097);
nor U6607 (N_6607,N_1641,N_2730);
or U6608 (N_6608,N_1236,N_2481);
xor U6609 (N_6609,N_4901,N_3545);
nand U6610 (N_6610,N_733,N_722);
or U6611 (N_6611,N_3112,N_1856);
or U6612 (N_6612,N_1812,N_1066);
nand U6613 (N_6613,N_2740,N_2079);
nor U6614 (N_6614,N_3389,N_1705);
and U6615 (N_6615,N_1319,N_2799);
nor U6616 (N_6616,N_2721,N_235);
or U6617 (N_6617,N_4922,N_2881);
nor U6618 (N_6618,N_702,N_2084);
nor U6619 (N_6619,N_3565,N_1884);
nand U6620 (N_6620,N_4478,N_3572);
nor U6621 (N_6621,N_3489,N_2540);
nand U6622 (N_6622,N_2779,N_555);
and U6623 (N_6623,N_2251,N_2909);
nand U6624 (N_6624,N_4330,N_2416);
nand U6625 (N_6625,N_3201,N_2376);
xor U6626 (N_6626,N_3683,N_2435);
xnor U6627 (N_6627,N_3465,N_1919);
and U6628 (N_6628,N_2366,N_3806);
and U6629 (N_6629,N_3999,N_4624);
and U6630 (N_6630,N_2447,N_703);
nor U6631 (N_6631,N_2482,N_1261);
or U6632 (N_6632,N_199,N_1904);
and U6633 (N_6633,N_4075,N_4634);
or U6634 (N_6634,N_1229,N_1394);
nor U6635 (N_6635,N_955,N_3372);
and U6636 (N_6636,N_4974,N_3960);
nand U6637 (N_6637,N_3476,N_252);
nor U6638 (N_6638,N_3672,N_3022);
nor U6639 (N_6639,N_1218,N_4454);
and U6640 (N_6640,N_4148,N_2728);
or U6641 (N_6641,N_168,N_563);
and U6642 (N_6642,N_3234,N_2228);
xor U6643 (N_6643,N_3075,N_1852);
nor U6644 (N_6644,N_4493,N_3961);
or U6645 (N_6645,N_1561,N_3707);
and U6646 (N_6646,N_4019,N_3320);
nand U6647 (N_6647,N_2179,N_4976);
nor U6648 (N_6648,N_3409,N_3059);
and U6649 (N_6649,N_1107,N_2263);
nor U6650 (N_6650,N_4849,N_879);
nand U6651 (N_6651,N_991,N_2250);
and U6652 (N_6652,N_2351,N_2197);
and U6653 (N_6653,N_4797,N_731);
nor U6654 (N_6654,N_3205,N_770);
nand U6655 (N_6655,N_434,N_766);
and U6656 (N_6656,N_699,N_3374);
and U6657 (N_6657,N_2017,N_3395);
or U6658 (N_6658,N_2471,N_1520);
nand U6659 (N_6659,N_4846,N_1033);
xnor U6660 (N_6660,N_186,N_448);
nor U6661 (N_6661,N_4950,N_4498);
and U6662 (N_6662,N_2765,N_3710);
nor U6663 (N_6663,N_2442,N_4246);
nand U6664 (N_6664,N_4127,N_4888);
or U6665 (N_6665,N_2767,N_951);
xor U6666 (N_6666,N_1234,N_278);
nor U6667 (N_6667,N_1320,N_3893);
xnor U6668 (N_6668,N_4138,N_2982);
and U6669 (N_6669,N_1652,N_276);
nand U6670 (N_6670,N_2450,N_1271);
xnor U6671 (N_6671,N_393,N_4929);
and U6672 (N_6672,N_4713,N_4082);
nand U6673 (N_6673,N_2343,N_1651);
xnor U6674 (N_6674,N_4889,N_1194);
and U6675 (N_6675,N_3618,N_1086);
or U6676 (N_6676,N_3532,N_1417);
nor U6677 (N_6677,N_1284,N_1816);
and U6678 (N_6678,N_3454,N_1653);
xnor U6679 (N_6679,N_3140,N_3884);
nor U6680 (N_6680,N_638,N_2134);
nand U6681 (N_6681,N_2265,N_2879);
nor U6682 (N_6682,N_3629,N_1376);
or U6683 (N_6683,N_3504,N_1607);
or U6684 (N_6684,N_1565,N_3118);
nor U6685 (N_6685,N_45,N_2845);
nor U6686 (N_6686,N_4874,N_4750);
and U6687 (N_6687,N_3718,N_353);
nor U6688 (N_6688,N_205,N_4436);
or U6689 (N_6689,N_1020,N_1740);
xor U6690 (N_6690,N_4591,N_4644);
xor U6691 (N_6691,N_2161,N_2816);
nand U6692 (N_6692,N_4149,N_4507);
or U6693 (N_6693,N_1111,N_2320);
and U6694 (N_6694,N_1829,N_608);
nor U6695 (N_6695,N_4024,N_3881);
or U6696 (N_6696,N_970,N_3157);
nor U6697 (N_6697,N_3097,N_2239);
nor U6698 (N_6698,N_674,N_1487);
and U6699 (N_6699,N_103,N_359);
xnor U6700 (N_6700,N_715,N_950);
and U6701 (N_6701,N_1288,N_1957);
or U6702 (N_6702,N_3161,N_4668);
or U6703 (N_6703,N_4183,N_3111);
xnor U6704 (N_6704,N_2201,N_4898);
nand U6705 (N_6705,N_2895,N_2206);
and U6706 (N_6706,N_4307,N_2029);
or U6707 (N_6707,N_1984,N_4400);
nor U6708 (N_6708,N_3269,N_4875);
nor U6709 (N_6709,N_914,N_3238);
nand U6710 (N_6710,N_4744,N_251);
xor U6711 (N_6711,N_1878,N_4704);
nand U6712 (N_6712,N_3693,N_2973);
and U6713 (N_6713,N_210,N_98);
or U6714 (N_6714,N_4300,N_1022);
or U6715 (N_6715,N_1717,N_36);
nand U6716 (N_6716,N_2679,N_4239);
nor U6717 (N_6717,N_1032,N_1725);
xnor U6718 (N_6718,N_3241,N_1186);
and U6719 (N_6719,N_2913,N_1978);
or U6720 (N_6720,N_4178,N_4529);
nor U6721 (N_6721,N_980,N_1790);
and U6722 (N_6722,N_3198,N_2692);
nand U6723 (N_6723,N_1915,N_2534);
nor U6724 (N_6724,N_1513,N_3684);
nor U6725 (N_6725,N_4088,N_978);
nand U6726 (N_6726,N_1130,N_1488);
and U6727 (N_6727,N_376,N_4882);
nand U6728 (N_6728,N_2230,N_3851);
or U6729 (N_6729,N_769,N_757);
nand U6730 (N_6730,N_3239,N_4462);
nand U6731 (N_6731,N_2668,N_1366);
xnor U6732 (N_6732,N_3597,N_2339);
and U6733 (N_6733,N_3248,N_1707);
nor U6734 (N_6734,N_1882,N_1286);
and U6735 (N_6735,N_3170,N_415);
xor U6736 (N_6736,N_1879,N_3772);
nand U6737 (N_6737,N_1489,N_3758);
or U6738 (N_6738,N_708,N_3307);
or U6739 (N_6739,N_2784,N_462);
xor U6740 (N_6740,N_1998,N_15);
or U6741 (N_6741,N_480,N_2722);
nand U6742 (N_6742,N_4334,N_1073);
xor U6743 (N_6743,N_496,N_2602);
nor U6744 (N_6744,N_1733,N_2502);
and U6745 (N_6745,N_4596,N_3755);
nor U6746 (N_6746,N_2815,N_2861);
nor U6747 (N_6747,N_3873,N_2348);
nor U6748 (N_6748,N_3778,N_3586);
nand U6749 (N_6749,N_256,N_1196);
and U6750 (N_6750,N_746,N_3911);
and U6751 (N_6751,N_3407,N_1497);
or U6752 (N_6752,N_4037,N_1820);
nand U6753 (N_6753,N_2221,N_4408);
nand U6754 (N_6754,N_3440,N_538);
nand U6755 (N_6755,N_571,N_366);
nand U6756 (N_6756,N_1558,N_2461);
nor U6757 (N_6757,N_2341,N_4253);
and U6758 (N_6758,N_3561,N_4119);
and U6759 (N_6759,N_866,N_4690);
xnor U6760 (N_6760,N_2688,N_4413);
and U6761 (N_6761,N_2444,N_4918);
or U6762 (N_6762,N_2473,N_2146);
and U6763 (N_6763,N_419,N_2584);
nand U6764 (N_6764,N_4546,N_3183);
nand U6765 (N_6765,N_4956,N_223);
or U6766 (N_6766,N_3972,N_190);
and U6767 (N_6767,N_2136,N_431);
or U6768 (N_6768,N_2451,N_4050);
xor U6769 (N_6769,N_2222,N_4122);
and U6770 (N_6770,N_2283,N_142);
and U6771 (N_6771,N_21,N_1702);
or U6772 (N_6772,N_44,N_1245);
nor U6773 (N_6773,N_1010,N_2544);
nor U6774 (N_6774,N_3587,N_4995);
and U6775 (N_6775,N_3763,N_3123);
nand U6776 (N_6776,N_3146,N_196);
or U6777 (N_6777,N_4089,N_1927);
nor U6778 (N_6778,N_1680,N_971);
or U6779 (N_6779,N_4278,N_3130);
nor U6780 (N_6780,N_3207,N_1894);
and U6781 (N_6781,N_1578,N_1945);
and U6782 (N_6782,N_3313,N_3818);
and U6783 (N_6783,N_1643,N_4847);
nand U6784 (N_6784,N_207,N_3560);
nand U6785 (N_6785,N_3050,N_382);
or U6786 (N_6786,N_2698,N_2370);
or U6787 (N_6787,N_389,N_1179);
nor U6788 (N_6788,N_2094,N_1113);
xnor U6789 (N_6789,N_2106,N_654);
xor U6790 (N_6790,N_1302,N_2211);
and U6791 (N_6791,N_1843,N_819);
nor U6792 (N_6792,N_4391,N_1509);
and U6793 (N_6793,N_2610,N_4745);
nor U6794 (N_6794,N_1837,N_2080);
nand U6795 (N_6795,N_575,N_1764);
nand U6796 (N_6796,N_789,N_2314);
nor U6797 (N_6797,N_3247,N_2709);
nor U6798 (N_6798,N_1672,N_4497);
xor U6799 (N_6799,N_4258,N_829);
or U6800 (N_6800,N_1369,N_212);
nor U6801 (N_6801,N_3036,N_1947);
nand U6802 (N_6802,N_3367,N_3738);
and U6803 (N_6803,N_1150,N_259);
or U6804 (N_6804,N_1742,N_1326);
or U6805 (N_6805,N_1677,N_658);
or U6806 (N_6806,N_4168,N_764);
nor U6807 (N_6807,N_3336,N_4669);
nand U6808 (N_6808,N_576,N_2568);
nor U6809 (N_6809,N_2323,N_1748);
or U6810 (N_6810,N_4021,N_1518);
nor U6811 (N_6811,N_2008,N_222);
nor U6812 (N_6812,N_1844,N_4601);
nor U6813 (N_6813,N_4202,N_2021);
nand U6814 (N_6814,N_2288,N_2643);
and U6815 (N_6815,N_3607,N_1313);
nor U6816 (N_6816,N_2632,N_873);
nand U6817 (N_6817,N_1436,N_2735);
xor U6818 (N_6818,N_524,N_1943);
nor U6819 (N_6819,N_1002,N_189);
nor U6820 (N_6820,N_3191,N_3542);
xor U6821 (N_6821,N_817,N_3340);
or U6822 (N_6822,N_3865,N_475);
nor U6823 (N_6823,N_2249,N_342);
or U6824 (N_6824,N_4163,N_1388);
and U6825 (N_6825,N_1364,N_2954);
nor U6826 (N_6826,N_4094,N_2672);
or U6827 (N_6827,N_3311,N_4781);
nor U6828 (N_6828,N_853,N_4551);
or U6829 (N_6829,N_2119,N_3950);
nor U6830 (N_6830,N_4130,N_194);
nor U6831 (N_6831,N_2702,N_3704);
and U6832 (N_6832,N_2128,N_1358);
nand U6833 (N_6833,N_507,N_923);
or U6834 (N_6834,N_2081,N_4042);
and U6835 (N_6835,N_4269,N_2823);
or U6836 (N_6836,N_1201,N_165);
nand U6837 (N_6837,N_3081,N_3602);
or U6838 (N_6838,N_1418,N_68);
nor U6839 (N_6839,N_1365,N_4780);
nor U6840 (N_6840,N_2291,N_1896);
or U6841 (N_6841,N_599,N_2701);
nand U6842 (N_6842,N_3945,N_3415);
nor U6843 (N_6843,N_1594,N_325);
and U6844 (N_6844,N_4506,N_3992);
and U6845 (N_6845,N_1692,N_4182);
and U6846 (N_6846,N_726,N_4655);
nor U6847 (N_6847,N_4850,N_2497);
nand U6848 (N_6848,N_3877,N_3799);
nand U6849 (N_6849,N_3752,N_4573);
nand U6850 (N_6850,N_3583,N_517);
and U6851 (N_6851,N_1301,N_4312);
or U6852 (N_6852,N_1343,N_898);
or U6853 (N_6853,N_1544,N_1025);
xor U6854 (N_6854,N_4041,N_2896);
nor U6855 (N_6855,N_3067,N_1075);
or U6856 (N_6856,N_3250,N_1604);
nor U6857 (N_6857,N_884,N_1808);
nand U6858 (N_6858,N_4818,N_1185);
nand U6859 (N_6859,N_1336,N_2616);
or U6860 (N_6860,N_3695,N_3450);
or U6861 (N_6861,N_2436,N_185);
nand U6862 (N_6862,N_1779,N_4410);
nor U6863 (N_6863,N_17,N_4902);
nand U6864 (N_6864,N_3019,N_723);
or U6865 (N_6865,N_592,N_3009);
nor U6866 (N_6866,N_534,N_3446);
nor U6867 (N_6867,N_4096,N_2805);
or U6868 (N_6868,N_1458,N_2922);
or U6869 (N_6869,N_4051,N_1877);
nor U6870 (N_6870,N_1412,N_2102);
nor U6871 (N_6871,N_1616,N_3667);
nor U6872 (N_6872,N_862,N_3078);
nand U6873 (N_6873,N_3769,N_2775);
or U6874 (N_6874,N_141,N_3867);
and U6875 (N_6875,N_2424,N_3506);
nor U6876 (N_6876,N_1525,N_2465);
xnor U6877 (N_6877,N_3720,N_188);
nand U6878 (N_6878,N_1090,N_470);
and U6879 (N_6879,N_217,N_1372);
and U6880 (N_6880,N_3880,N_720);
nor U6881 (N_6881,N_4985,N_855);
xor U6882 (N_6882,N_611,N_514);
or U6883 (N_6883,N_3802,N_3365);
nor U6884 (N_6884,N_2018,N_1030);
nand U6885 (N_6885,N_1875,N_2330);
nor U6886 (N_6886,N_1772,N_4004);
nor U6887 (N_6887,N_4716,N_282);
or U6888 (N_6888,N_4463,N_374);
or U6889 (N_6889,N_2613,N_1950);
nand U6890 (N_6890,N_957,N_4011);
and U6891 (N_6891,N_2224,N_2159);
nor U6892 (N_6892,N_133,N_1112);
and U6893 (N_6893,N_2963,N_3466);
nor U6894 (N_6894,N_2417,N_1530);
xnor U6895 (N_6895,N_3048,N_4867);
nand U6896 (N_6896,N_1021,N_2862);
and U6897 (N_6897,N_605,N_3706);
nor U6898 (N_6898,N_377,N_2149);
nor U6899 (N_6899,N_686,N_2940);
and U6900 (N_6900,N_4032,N_4340);
nor U6901 (N_6901,N_4783,N_2921);
nor U6902 (N_6902,N_2045,N_4044);
nand U6903 (N_6903,N_1917,N_1670);
xnor U6904 (N_6904,N_1909,N_775);
and U6905 (N_6905,N_4673,N_2037);
nand U6906 (N_6906,N_1975,N_403);
and U6907 (N_6907,N_724,N_4458);
nand U6908 (N_6908,N_1464,N_3449);
nand U6909 (N_6909,N_3814,N_1054);
and U6910 (N_6910,N_2878,N_1212);
and U6911 (N_6911,N_3174,N_4371);
and U6912 (N_6912,N_930,N_3746);
or U6913 (N_6913,N_3648,N_3980);
nand U6914 (N_6914,N_295,N_3895);
nor U6915 (N_6915,N_4425,N_3251);
nor U6916 (N_6916,N_4833,N_1151);
nor U6917 (N_6917,N_3665,N_10);
or U6918 (N_6918,N_4069,N_3501);
or U6919 (N_6919,N_1117,N_1270);
and U6920 (N_6920,N_4398,N_1348);
nor U6921 (N_6921,N_728,N_3774);
nand U6922 (N_6922,N_344,N_3317);
nand U6923 (N_6923,N_3194,N_4373);
or U6924 (N_6924,N_1848,N_1682);
nand U6925 (N_6925,N_4343,N_2952);
or U6926 (N_6926,N_3461,N_4676);
nor U6927 (N_6927,N_872,N_3451);
nor U6928 (N_6928,N_4642,N_1377);
nand U6929 (N_6929,N_4880,N_463);
or U6930 (N_6930,N_4631,N_2695);
xnor U6931 (N_6931,N_4571,N_1023);
or U6932 (N_6932,N_1815,N_1072);
and U6933 (N_6933,N_3105,N_3032);
nor U6934 (N_6934,N_1491,N_1381);
nand U6935 (N_6935,N_4725,N_291);
or U6936 (N_6936,N_2057,N_1839);
xnor U6937 (N_6937,N_4717,N_38);
nor U6938 (N_6938,N_1095,N_1103);
nand U6939 (N_6939,N_2801,N_253);
nand U6940 (N_6940,N_4143,N_3737);
nand U6941 (N_6941,N_3379,N_122);
xor U6942 (N_6942,N_337,N_3436);
nor U6943 (N_6943,N_365,N_4285);
or U6944 (N_6944,N_4821,N_4563);
nor U6945 (N_6945,N_1403,N_924);
and U6946 (N_6946,N_2593,N_1698);
nor U6947 (N_6947,N_528,N_2020);
or U6948 (N_6948,N_4705,N_4405);
or U6949 (N_6949,N_203,N_307);
nor U6950 (N_6950,N_1938,N_4379);
and U6951 (N_6951,N_2986,N_4692);
nand U6952 (N_6952,N_2893,N_4727);
nand U6953 (N_6953,N_3912,N_2535);
nor U6954 (N_6954,N_2588,N_3570);
nor U6955 (N_6955,N_3650,N_1830);
and U6956 (N_6956,N_2426,N_1499);
and U6957 (N_6957,N_4064,N_543);
nand U6958 (N_6958,N_3062,N_3042);
and U6959 (N_6959,N_4793,N_4013);
nor U6960 (N_6960,N_3503,N_806);
nand U6961 (N_6961,N_1863,N_1096);
or U6962 (N_6962,N_4369,N_4659);
or U6963 (N_6963,N_1074,N_372);
or U6964 (N_6964,N_2368,N_1180);
nor U6965 (N_6965,N_4711,N_964);
and U6966 (N_6966,N_4194,N_1522);
xnor U6967 (N_6967,N_1396,N_2261);
xor U6968 (N_6968,N_4068,N_2906);
nor U6969 (N_6969,N_4899,N_3463);
nor U6970 (N_6970,N_2406,N_1822);
nand U6971 (N_6971,N_0,N_913);
and U6972 (N_6972,N_3093,N_1227);
or U6973 (N_6973,N_66,N_2569);
xnor U6974 (N_6974,N_3196,N_1630);
and U6975 (N_6975,N_4520,N_2356);
nand U6976 (N_6976,N_406,N_1501);
and U6977 (N_6977,N_175,N_4031);
xor U6978 (N_6978,N_2116,N_4795);
nor U6979 (N_6979,N_4374,N_2074);
or U6980 (N_6980,N_2264,N_443);
and U6981 (N_6981,N_4433,N_4646);
nor U6982 (N_6982,N_2318,N_1614);
or U6983 (N_6983,N_3020,N_1954);
nand U6984 (N_6984,N_2058,N_444);
or U6985 (N_6985,N_1595,N_3434);
nor U6986 (N_6986,N_1729,N_4108);
nor U6987 (N_6987,N_1645,N_4971);
nand U6988 (N_6988,N_3388,N_2486);
xnor U6989 (N_6989,N_2144,N_1736);
and U6990 (N_6990,N_2556,N_570);
nand U6991 (N_6991,N_174,N_1517);
nand U6992 (N_6992,N_4996,N_2903);
or U6993 (N_6993,N_906,N_3714);
and U6994 (N_6994,N_85,N_3949);
and U6995 (N_6995,N_1057,N_4065);
or U6996 (N_6996,N_2489,N_2969);
nor U6997 (N_6997,N_1400,N_642);
or U6998 (N_6998,N_4852,N_1470);
nand U6999 (N_6999,N_2389,N_1761);
and U7000 (N_7000,N_1454,N_4864);
nand U7001 (N_7001,N_4107,N_1471);
or U7002 (N_7002,N_1596,N_4290);
and U7003 (N_7003,N_994,N_3222);
and U7004 (N_7004,N_3953,N_778);
and U7005 (N_7005,N_4521,N_4492);
nor U7006 (N_7006,N_1564,N_2553);
xor U7007 (N_7007,N_2888,N_4125);
or U7008 (N_7008,N_3905,N_2768);
nor U7009 (N_7009,N_3830,N_3927);
and U7010 (N_7010,N_1796,N_1414);
nand U7011 (N_7011,N_2445,N_1137);
nor U7012 (N_7012,N_1434,N_4917);
and U7013 (N_7013,N_4310,N_2038);
and U7014 (N_7014,N_1639,N_635);
nand U7015 (N_7015,N_1312,N_4756);
or U7016 (N_7016,N_3467,N_4286);
nor U7017 (N_7017,N_2458,N_4854);
or U7018 (N_7018,N_209,N_4802);
nand U7019 (N_7019,N_1496,N_3923);
nor U7020 (N_7020,N_4196,N_1340);
and U7021 (N_7021,N_4384,N_926);
or U7022 (N_7022,N_1589,N_4281);
or U7023 (N_7023,N_334,N_4214);
xnor U7024 (N_7024,N_4446,N_1081);
nor U7025 (N_7025,N_4453,N_4590);
and U7026 (N_7026,N_2011,N_290);
nand U7027 (N_7027,N_31,N_1667);
nor U7028 (N_7028,N_3444,N_3858);
nor U7029 (N_7029,N_249,N_4131);
nand U7030 (N_7030,N_2243,N_3643);
or U7031 (N_7031,N_3184,N_1706);
and U7032 (N_7032,N_4097,N_1240);
nand U7033 (N_7033,N_1775,N_3258);
and U7034 (N_7034,N_4532,N_1605);
or U7035 (N_7035,N_2825,N_4923);
nor U7036 (N_7036,N_130,N_3784);
and U7037 (N_7037,N_447,N_3426);
and U7038 (N_7038,N_2229,N_330);
or U7039 (N_7039,N_3412,N_717);
nand U7040 (N_7040,N_1539,N_777);
and U7041 (N_7041,N_320,N_2403);
nand U7042 (N_7042,N_2404,N_491);
or U7043 (N_7043,N_4018,N_3677);
and U7044 (N_7044,N_4828,N_897);
nor U7045 (N_7045,N_1640,N_1392);
nor U7046 (N_7046,N_1409,N_2358);
and U7047 (N_7047,N_3475,N_2457);
or U7048 (N_7048,N_681,N_2463);
or U7049 (N_7049,N_2778,N_967);
nor U7050 (N_7050,N_747,N_4949);
and U7051 (N_7051,N_2618,N_2772);
or U7052 (N_7052,N_3990,N_1755);
nor U7053 (N_7053,N_211,N_1548);
nor U7054 (N_7054,N_4154,N_4640);
nand U7055 (N_7055,N_2601,N_609);
nand U7056 (N_7056,N_1655,N_1024);
or U7057 (N_7057,N_1833,N_3866);
or U7058 (N_7058,N_2563,N_613);
nand U7059 (N_7059,N_2398,N_2093);
and U7060 (N_7060,N_2624,N_911);
nor U7061 (N_7061,N_1719,N_983);
and U7062 (N_7062,N_3421,N_1280);
and U7063 (N_7063,N_3682,N_466);
or U7064 (N_7064,N_2266,N_2686);
nand U7065 (N_7065,N_20,N_700);
and U7066 (N_7066,N_2724,N_2802);
nand U7067 (N_7067,N_1569,N_2198);
or U7068 (N_7068,N_4375,N_1626);
nor U7069 (N_7069,N_3236,N_3776);
nor U7070 (N_7070,N_4973,N_1880);
and U7071 (N_7071,N_2528,N_145);
nand U7072 (N_7072,N_1800,N_3353);
and U7073 (N_7073,N_3579,N_1629);
xnor U7074 (N_7074,N_881,N_3963);
and U7075 (N_7075,N_3521,N_2087);
and U7076 (N_7076,N_4360,N_1709);
nor U7077 (N_7077,N_3721,N_1519);
or U7078 (N_7078,N_4005,N_3346);
and U7079 (N_7079,N_2414,N_2919);
xor U7080 (N_7080,N_2331,N_1423);
nor U7081 (N_7081,N_894,N_1238);
and U7082 (N_7082,N_4177,N_745);
nor U7083 (N_7083,N_3240,N_606);
nor U7084 (N_7084,N_1378,N_1827);
or U7085 (N_7085,N_2407,N_1291);
and U7086 (N_7086,N_1902,N_3843);
or U7087 (N_7087,N_2375,N_3605);
and U7088 (N_7088,N_2564,N_1359);
nand U7089 (N_7089,N_956,N_2754);
or U7090 (N_7090,N_4595,N_4028);
nand U7091 (N_7091,N_120,N_2989);
and U7092 (N_7092,N_519,N_2207);
or U7093 (N_7093,N_743,N_4208);
nand U7094 (N_7094,N_954,N_540);
and U7095 (N_7095,N_2917,N_2280);
or U7096 (N_7096,N_1092,N_281);
nor U7097 (N_7097,N_1512,N_513);
xor U7098 (N_7098,N_752,N_3967);
nor U7099 (N_7099,N_2663,N_4528);
and U7100 (N_7100,N_3580,N_1903);
or U7101 (N_7101,N_176,N_80);
and U7102 (N_7102,N_3946,N_4009);
nor U7103 (N_7103,N_2597,N_2298);
or U7104 (N_7104,N_3985,N_4431);
nand U7105 (N_7105,N_3121,N_442);
and U7106 (N_7106,N_2,N_3366);
nand U7107 (N_7107,N_4079,N_4186);
or U7108 (N_7108,N_2717,N_2590);
or U7109 (N_7109,N_1016,N_3220);
and U7110 (N_7110,N_669,N_2114);
nand U7111 (N_7111,N_854,N_4015);
nor U7112 (N_7112,N_4968,N_2720);
and U7113 (N_7113,N_4662,N_1084);
xnor U7114 (N_7114,N_2067,N_2875);
nor U7115 (N_7115,N_3094,N_3598);
xor U7116 (N_7116,N_4761,N_2432);
or U7117 (N_7117,N_2453,N_2164);
nand U7118 (N_7118,N_2630,N_437);
and U7119 (N_7119,N_3742,N_4381);
or U7120 (N_7120,N_2166,N_698);
xor U7121 (N_7121,N_4420,N_892);
nand U7122 (N_7122,N_2384,N_4771);
nand U7123 (N_7123,N_3266,N_3781);
xor U7124 (N_7124,N_3790,N_1586);
nand U7125 (N_7125,N_1164,N_4641);
nand U7126 (N_7126,N_1972,N_3928);
nand U7127 (N_7127,N_4810,N_1058);
nor U7128 (N_7128,N_4675,N_2326);
or U7129 (N_7129,N_57,N_4209);
nor U7130 (N_7130,N_3060,N_2621);
and U7131 (N_7131,N_2301,N_3908);
nand U7132 (N_7132,N_3557,N_1152);
xnor U7133 (N_7133,N_4574,N_3921);
or U7134 (N_7134,N_691,N_12);
and U7135 (N_7135,N_4650,N_3549);
nand U7136 (N_7136,N_3403,N_593);
nor U7137 (N_7137,N_2275,N_1583);
nand U7138 (N_7138,N_1806,N_3939);
nand U7139 (N_7139,N_289,N_4085);
or U7140 (N_7140,N_1547,N_1484);
nor U7141 (N_7141,N_4736,N_1279);
or U7142 (N_7142,N_933,N_2441);
nand U7143 (N_7143,N_3187,N_4606);
xor U7144 (N_7144,N_4526,N_3574);
or U7145 (N_7145,N_4811,N_1136);
xnor U7146 (N_7146,N_3826,N_4858);
xor U7147 (N_7147,N_3193,N_582);
and U7148 (N_7148,N_842,N_578);
nor U7149 (N_7149,N_3176,N_4195);
or U7150 (N_7150,N_1034,N_2028);
nand U7151 (N_7151,N_3481,N_2296);
nor U7152 (N_7152,N_3369,N_4561);
or U7153 (N_7153,N_487,N_2344);
nand U7154 (N_7154,N_2041,N_1872);
nand U7155 (N_7155,N_4770,N_690);
nand U7156 (N_7156,N_1660,N_3277);
xor U7157 (N_7157,N_3947,N_2598);
nand U7158 (N_7158,N_1142,N_2223);
nand U7159 (N_7159,N_1217,N_4835);
or U7160 (N_7160,N_2208,N_1371);
nor U7161 (N_7161,N_947,N_4961);
and U7162 (N_7162,N_1536,N_1455);
nand U7163 (N_7163,N_3625,N_2760);
and U7164 (N_7164,N_3164,N_62);
nor U7165 (N_7165,N_265,N_4661);
xor U7166 (N_7166,N_2910,N_245);
nor U7167 (N_7167,N_4289,N_4984);
or U7168 (N_7168,N_4645,N_3901);
nor U7169 (N_7169,N_2449,N_4764);
or U7170 (N_7170,N_1093,N_905);
nor U7171 (N_7171,N_2088,N_3834);
nor U7172 (N_7172,N_2653,N_3573);
or U7173 (N_7173,N_1202,N_2585);
nand U7174 (N_7174,N_580,N_2565);
and U7175 (N_7175,N_1321,N_2327);
and U7176 (N_7176,N_236,N_285);
and U7177 (N_7177,N_3177,N_3316);
xnor U7178 (N_7178,N_2124,N_4437);
and U7179 (N_7179,N_4930,N_3363);
nand U7180 (N_7180,N_556,N_765);
and U7181 (N_7181,N_4423,N_4567);
nor U7182 (N_7182,N_4698,N_136);
and U7183 (N_7183,N_1747,N_3732);
nand U7184 (N_7184,N_564,N_4562);
nor U7185 (N_7185,N_4012,N_3152);
xor U7186 (N_7186,N_2321,N_4581);
xnor U7187 (N_7187,N_481,N_791);
nand U7188 (N_7188,N_1753,N_1012);
nand U7189 (N_7189,N_4545,N_2706);
nand U7190 (N_7190,N_2125,N_3653);
and U7191 (N_7191,N_4262,N_3329);
and U7192 (N_7192,N_1485,N_4399);
or U7193 (N_7193,N_4322,N_3989);
or U7194 (N_7194,N_574,N_2476);
xor U7195 (N_7195,N_247,N_3646);
nor U7196 (N_7196,N_4649,N_4840);
nand U7197 (N_7197,N_2933,N_4008);
nand U7198 (N_7198,N_2129,N_2232);
and U7199 (N_7199,N_378,N_844);
xnor U7200 (N_7200,N_831,N_2923);
or U7201 (N_7201,N_2252,N_3330);
and U7202 (N_7202,N_2083,N_4837);
or U7203 (N_7203,N_3186,N_627);
nor U7204 (N_7204,N_4255,N_1144);
and U7205 (N_7205,N_4937,N_96);
nand U7206 (N_7206,N_2803,N_4415);
and U7207 (N_7207,N_1598,N_412);
nor U7208 (N_7208,N_2338,N_4602);
xor U7209 (N_7209,N_3689,N_4558);
or U7210 (N_7210,N_2096,N_2749);
xor U7211 (N_7211,N_3924,N_2926);
nand U7212 (N_7212,N_4831,N_3562);
or U7213 (N_7213,N_459,N_813);
nor U7214 (N_7214,N_3058,N_2141);
and U7215 (N_7215,N_238,N_347);
nor U7216 (N_7216,N_2622,N_3392);
and U7217 (N_7217,N_2744,N_1337);
and U7218 (N_7218,N_356,N_4789);
xnor U7219 (N_7219,N_4832,N_4550);
nand U7220 (N_7220,N_3260,N_1953);
nand U7221 (N_7221,N_49,N_51);
and U7222 (N_7222,N_3084,N_2726);
or U7223 (N_7223,N_846,N_408);
nor U7224 (N_7224,N_3692,N_1198);
nor U7225 (N_7225,N_533,N_2004);
nand U7226 (N_7226,N_904,N_4663);
nand U7227 (N_7227,N_3852,N_974);
nand U7228 (N_7228,N_1804,N_4652);
nand U7229 (N_7229,N_1216,N_1590);
xor U7230 (N_7230,N_171,N_886);
or U7231 (N_7231,N_4038,N_4456);
or U7232 (N_7232,N_3722,N_346);
nand U7233 (N_7233,N_3723,N_3713);
nand U7234 (N_7234,N_267,N_3153);
and U7235 (N_7235,N_3876,N_76);
nor U7236 (N_7236,N_2750,N_163);
nand U7237 (N_7237,N_3863,N_4796);
nand U7238 (N_7238,N_4788,N_2880);
nor U7239 (N_7239,N_220,N_4353);
xnor U7240 (N_7240,N_3973,N_2774);
nor U7241 (N_7241,N_2273,N_867);
xor U7242 (N_7242,N_1559,N_4709);
and U7243 (N_7243,N_1554,N_385);
or U7244 (N_7244,N_584,N_3442);
or U7245 (N_7245,N_105,N_2448);
nand U7246 (N_7246,N_3875,N_3136);
nor U7247 (N_7247,N_3052,N_4609);
and U7248 (N_7248,N_1931,N_4499);
or U7249 (N_7249,N_1041,N_1305);
or U7250 (N_7250,N_4763,N_4798);
and U7251 (N_7251,N_1730,N_1476);
and U7252 (N_7252,N_1810,N_1562);
xnor U7253 (N_7253,N_1277,N_1178);
nand U7254 (N_7254,N_2583,N_4280);
nor U7255 (N_7255,N_647,N_3116);
nor U7256 (N_7256,N_3208,N_2612);
nand U7257 (N_7257,N_1550,N_2842);
xnor U7258 (N_7258,N_598,N_375);
and U7259 (N_7259,N_3571,N_3280);
or U7260 (N_7260,N_413,N_2357);
nand U7261 (N_7261,N_74,N_4895);
or U7262 (N_7262,N_1712,N_4841);
and U7263 (N_7263,N_1223,N_3267);
and U7264 (N_7264,N_3229,N_665);
nor U7265 (N_7265,N_2050,N_148);
or U7266 (N_7266,N_1036,N_2300);
nor U7267 (N_7267,N_4982,N_4014);
xnor U7268 (N_7268,N_3736,N_2429);
nand U7269 (N_7269,N_2877,N_3122);
or U7270 (N_7270,N_322,N_2607);
nor U7271 (N_7271,N_1039,N_1523);
nor U7272 (N_7272,N_2108,N_2311);
or U7273 (N_7273,N_2510,N_1003);
nor U7274 (N_7274,N_4729,N_2089);
nor U7275 (N_7275,N_3678,N_3703);
nor U7276 (N_7276,N_407,N_4022);
nor U7277 (N_7277,N_384,N_4743);
nand U7278 (N_7278,N_4055,N_4559);
nor U7279 (N_7279,N_1166,N_1716);
nand U7280 (N_7280,N_1823,N_1053);
nor U7281 (N_7281,N_4174,N_150);
nor U7282 (N_7282,N_2103,N_3185);
nor U7283 (N_7283,N_1,N_2725);
or U7284 (N_7284,N_3987,N_625);
nor U7285 (N_7285,N_3517,N_1897);
and U7286 (N_7286,N_1932,N_4217);
nor U7287 (N_7287,N_4983,N_4724);
nor U7288 (N_7288,N_1964,N_3045);
or U7289 (N_7289,N_371,N_4633);
nand U7290 (N_7290,N_2551,N_2693);
or U7291 (N_7291,N_2566,N_4394);
and U7292 (N_7292,N_69,N_1694);
nand U7293 (N_7293,N_2738,N_1325);
nand U7294 (N_7294,N_774,N_2682);
nor U7295 (N_7295,N_1656,N_1571);
and U7296 (N_7296,N_1533,N_869);
or U7297 (N_7297,N_4351,N_61);
nand U7298 (N_7298,N_2194,N_1944);
and U7299 (N_7299,N_4184,N_3016);
nand U7300 (N_7300,N_1439,N_2454);
or U7301 (N_7301,N_771,N_1156);
xnor U7302 (N_7302,N_843,N_2420);
nand U7303 (N_7303,N_3795,N_4766);
or U7304 (N_7304,N_1732,N_4845);
nor U7305 (N_7305,N_646,N_3272);
nor U7306 (N_7306,N_4485,N_2395);
and U7307 (N_7307,N_1992,N_2611);
or U7308 (N_7308,N_183,N_4081);
xor U7309 (N_7309,N_934,N_3083);
xor U7310 (N_7310,N_2763,N_3217);
or U7311 (N_7311,N_4935,N_59);
nor U7312 (N_7312,N_2666,N_4427);
nand U7313 (N_7313,N_4919,N_4941);
or U7314 (N_7314,N_3886,N_1462);
nand U7315 (N_7315,N_2455,N_2013);
or U7316 (N_7316,N_2837,N_2939);
nand U7317 (N_7317,N_2961,N_1293);
nor U7318 (N_7318,N_1248,N_1452);
nand U7319 (N_7319,N_357,N_4803);
and U7320 (N_7320,N_1349,N_1924);
nor U7321 (N_7321,N_311,N_3102);
xnor U7322 (N_7322,N_1577,N_4359);
nor U7323 (N_7323,N_2529,N_1527);
nor U7324 (N_7324,N_1671,N_441);
nand U7325 (N_7325,N_2707,N_2209);
or U7326 (N_7326,N_4524,N_262);
xor U7327 (N_7327,N_1266,N_3352);
nand U7328 (N_7328,N_4354,N_2617);
and U7329 (N_7329,N_2671,N_1456);
and U7330 (N_7330,N_4946,N_4311);
nor U7331 (N_7331,N_1441,N_4964);
nor U7332 (N_7332,N_3491,N_489);
nand U7333 (N_7333,N_4921,N_1976);
nor U7334 (N_7334,N_4074,N_2791);
nor U7335 (N_7335,N_3331,N_2245);
nor U7336 (N_7336,N_229,N_3810);
nor U7337 (N_7337,N_4604,N_2399);
xor U7338 (N_7338,N_4726,N_4623);
and U7339 (N_7339,N_3345,N_3623);
nand U7340 (N_7340,N_736,N_79);
xnor U7341 (N_7341,N_4200,N_2520);
nor U7342 (N_7342,N_3378,N_4870);
and U7343 (N_7343,N_1384,N_4099);
nor U7344 (N_7344,N_4939,N_1077);
nor U7345 (N_7345,N_2727,N_297);
nor U7346 (N_7346,N_1408,N_3295);
or U7347 (N_7347,N_1128,N_1601);
nand U7348 (N_7348,N_1315,N_2402);
and U7349 (N_7349,N_2929,N_1213);
nor U7350 (N_7350,N_1430,N_1169);
nor U7351 (N_7351,N_137,N_509);
and U7352 (N_7352,N_4317,N_1494);
xnor U7353 (N_7353,N_3103,N_30);
and U7354 (N_7354,N_1745,N_2214);
and U7355 (N_7355,N_4848,N_3558);
nor U7356 (N_7356,N_4259,N_1826);
xnor U7357 (N_7357,N_3917,N_3072);
nand U7358 (N_7358,N_3551,N_1759);
xor U7359 (N_7359,N_1490,N_738);
and U7360 (N_7360,N_3188,N_3306);
and U7361 (N_7361,N_4773,N_2137);
nand U7362 (N_7362,N_1119,N_2830);
or U7363 (N_7363,N_526,N_2091);
or U7364 (N_7364,N_1141,N_2771);
nand U7365 (N_7365,N_241,N_1295);
nor U7366 (N_7366,N_3428,N_2027);
xor U7367 (N_7367,N_1027,N_2220);
nand U7368 (N_7368,N_1809,N_1803);
and U7369 (N_7369,N_937,N_2033);
nor U7370 (N_7370,N_1715,N_560);
and U7371 (N_7371,N_2493,N_2953);
nand U7372 (N_7372,N_4816,N_2657);
nor U7373 (N_7373,N_1233,N_4927);
or U7374 (N_7374,N_3433,N_2792);
nor U7375 (N_7375,N_4772,N_493);
nand U7376 (N_7376,N_3192,N_4554);
nand U7377 (N_7377,N_2095,N_118);
and U7378 (N_7378,N_3259,N_2511);
nand U7379 (N_7379,N_798,N_3998);
and U7380 (N_7380,N_2633,N_4636);
and U7381 (N_7381,N_2998,N_549);
or U7382 (N_7382,N_4920,N_1836);
nor U7383 (N_7383,N_3427,N_1867);
or U7384 (N_7384,N_2340,N_324);
nor U7385 (N_7385,N_2578,N_1805);
nand U7386 (N_7386,N_2641,N_2240);
and U7387 (N_7387,N_1468,N_329);
nand U7388 (N_7388,N_482,N_2971);
nor U7389 (N_7389,N_3151,N_3812);
or U7390 (N_7390,N_938,N_2044);
and U7391 (N_7391,N_1575,N_4382);
nor U7392 (N_7392,N_2483,N_1226);
or U7393 (N_7393,N_4242,N_3154);
or U7394 (N_7394,N_3079,N_3492);
nand U7395 (N_7395,N_2546,N_4565);
and U7396 (N_7396,N_2405,N_1952);
nor U7397 (N_7397,N_3634,N_3591);
nor U7398 (N_7398,N_3654,N_1572);
nand U7399 (N_7399,N_2190,N_727);
or U7400 (N_7400,N_1817,N_3585);
or U7401 (N_7401,N_2295,N_8);
nor U7402 (N_7402,N_3892,N_3254);
nand U7403 (N_7403,N_601,N_3791);
nand U7404 (N_7404,N_2440,N_3528);
or U7405 (N_7405,N_1847,N_535);
nand U7406 (N_7406,N_492,N_3015);
nand U7407 (N_7407,N_3382,N_3628);
xnor U7408 (N_7408,N_1974,N_4884);
nor U7409 (N_7409,N_2127,N_4488);
nand U7410 (N_7410,N_4395,N_4062);
nand U7411 (N_7411,N_851,N_400);
xnor U7412 (N_7412,N_1778,N_3593);
nand U7413 (N_7413,N_3402,N_418);
xor U7414 (N_7414,N_948,N_2491);
and U7415 (N_7415,N_4527,N_2999);
and U7416 (N_7416,N_834,N_710);
nand U7417 (N_7417,N_3903,N_312);
and U7418 (N_7418,N_1744,N_4825);
and U7419 (N_7419,N_3552,N_2282);
and U7420 (N_7420,N_3524,N_95);
nand U7421 (N_7421,N_4469,N_2390);
nor U7422 (N_7422,N_483,N_3199);
and U7423 (N_7423,N_1646,N_2133);
nand U7424 (N_7424,N_1911,N_4121);
or U7425 (N_7425,N_4741,N_1926);
nor U7426 (N_7426,N_1507,N_707);
or U7427 (N_7427,N_2003,N_1017);
nor U7428 (N_7428,N_4345,N_469);
or U7429 (N_7429,N_2235,N_2685);
xor U7430 (N_7430,N_4872,N_3756);
nor U7431 (N_7431,N_4417,N_2180);
and U7432 (N_7432,N_1930,N_3848);
and U7433 (N_7433,N_4496,N_1508);
and U7434 (N_7434,N_2350,N_2172);
and U7435 (N_7435,N_2959,N_3096);
nor U7436 (N_7436,N_1552,N_1925);
nor U7437 (N_7437,N_3519,N_1846);
and U7438 (N_7438,N_181,N_226);
nor U7439 (N_7439,N_3957,N_3656);
and U7440 (N_7440,N_2619,N_1807);
or U7441 (N_7441,N_4931,N_345);
xnor U7442 (N_7442,N_4800,N_3829);
and U7443 (N_7443,N_2667,N_541);
and U7444 (N_7444,N_610,N_3373);
xor U7445 (N_7445,N_2352,N_3218);
and U7446 (N_7446,N_3702,N_1782);
or U7447 (N_7447,N_468,N_3680);
or U7448 (N_7448,N_2782,N_4467);
nand U7449 (N_7449,N_807,N_1597);
or U7450 (N_7450,N_2847,N_2634);
xnor U7451 (N_7451,N_2541,N_3599);
nor U7452 (N_7452,N_3156,N_4061);
xnor U7453 (N_7453,N_88,N_1477);
nor U7454 (N_7454,N_2150,N_4909);
or U7455 (N_7455,N_4681,N_3516);
or U7456 (N_7456,N_2364,N_2869);
or U7457 (N_7457,N_3902,N_333);
and U7458 (N_7458,N_3882,N_1849);
nand U7459 (N_7459,N_380,N_4534);
or U7460 (N_7460,N_2112,N_310);
and U7461 (N_7461,N_4787,N_368);
nand U7462 (N_7462,N_303,N_92);
and U7463 (N_7463,N_877,N_3578);
nand U7464 (N_7464,N_3420,N_4455);
or U7465 (N_7465,N_3356,N_3674);
or U7466 (N_7466,N_821,N_107);
nor U7467 (N_7467,N_1314,N_581);
and U7468 (N_7468,N_4755,N_3958);
nor U7469 (N_7469,N_4215,N_865);
or U7470 (N_7470,N_4052,N_4932);
or U7471 (N_7471,N_4073,N_4294);
and U7472 (N_7472,N_4110,N_595);
nor U7473 (N_7473,N_488,N_2950);
or U7474 (N_7474,N_2608,N_4735);
and U7475 (N_7475,N_3033,N_3698);
or U7476 (N_7476,N_4058,N_2974);
xnor U7477 (N_7477,N_2652,N_3364);
nor U7478 (N_7478,N_1638,N_3);
nand U7479 (N_7479,N_2035,N_2512);
and U7480 (N_7480,N_1225,N_2158);
or U7481 (N_7481,N_3349,N_4144);
xor U7482 (N_7482,N_2378,N_912);
nand U7483 (N_7483,N_180,N_3499);
and U7484 (N_7484,N_4945,N_255);
nor U7485 (N_7485,N_1028,N_1171);
nor U7486 (N_7486,N_2889,N_4997);
and U7487 (N_7487,N_3807,N_243);
nor U7488 (N_7488,N_3604,N_2855);
or U7489 (N_7489,N_4472,N_3195);
nor U7490 (N_7490,N_3021,N_232);
and U7491 (N_7491,N_2030,N_4161);
nand U7492 (N_7492,N_112,N_3820);
xnor U7493 (N_7493,N_3339,N_3242);
or U7494 (N_7494,N_4827,N_4401);
and U7495 (N_7495,N_639,N_4779);
or U7496 (N_7496,N_2488,N_3344);
and U7497 (N_7497,N_2419,N_2526);
or U7498 (N_7498,N_3833,N_4834);
or U7499 (N_7499,N_4279,N_1289);
nor U7500 (N_7500,N_306,N_1055);
and U7501 (N_7501,N_4799,N_1920);
or U7502 (N_7502,N_4698,N_1474);
or U7503 (N_7503,N_4229,N_2896);
and U7504 (N_7504,N_1465,N_483);
and U7505 (N_7505,N_1754,N_4684);
or U7506 (N_7506,N_39,N_3302);
nand U7507 (N_7507,N_2851,N_3528);
and U7508 (N_7508,N_2032,N_1568);
and U7509 (N_7509,N_1021,N_1814);
and U7510 (N_7510,N_4032,N_571);
and U7511 (N_7511,N_3216,N_3629);
nand U7512 (N_7512,N_4574,N_3910);
or U7513 (N_7513,N_3793,N_557);
or U7514 (N_7514,N_4659,N_3506);
xor U7515 (N_7515,N_4777,N_4580);
nor U7516 (N_7516,N_4090,N_4967);
and U7517 (N_7517,N_2443,N_2363);
nand U7518 (N_7518,N_4424,N_1493);
and U7519 (N_7519,N_1372,N_2051);
nand U7520 (N_7520,N_3817,N_1309);
nor U7521 (N_7521,N_4255,N_1331);
nor U7522 (N_7522,N_1889,N_3070);
or U7523 (N_7523,N_2415,N_4899);
or U7524 (N_7524,N_4282,N_3334);
or U7525 (N_7525,N_3054,N_0);
nor U7526 (N_7526,N_122,N_1689);
nand U7527 (N_7527,N_1684,N_1352);
nand U7528 (N_7528,N_1601,N_2150);
xor U7529 (N_7529,N_1560,N_3241);
and U7530 (N_7530,N_3002,N_993);
nor U7531 (N_7531,N_3076,N_794);
nor U7532 (N_7532,N_426,N_4416);
nand U7533 (N_7533,N_146,N_4825);
nand U7534 (N_7534,N_3435,N_752);
or U7535 (N_7535,N_4289,N_1806);
nand U7536 (N_7536,N_4238,N_4318);
and U7537 (N_7537,N_4478,N_1859);
nand U7538 (N_7538,N_2631,N_4367);
and U7539 (N_7539,N_4425,N_1660);
nand U7540 (N_7540,N_2830,N_3015);
xor U7541 (N_7541,N_451,N_3701);
nor U7542 (N_7542,N_1659,N_2535);
nor U7543 (N_7543,N_2691,N_3633);
nand U7544 (N_7544,N_500,N_6);
nor U7545 (N_7545,N_3214,N_2437);
or U7546 (N_7546,N_3765,N_3721);
nor U7547 (N_7547,N_3033,N_3710);
and U7548 (N_7548,N_2334,N_4518);
nor U7549 (N_7549,N_3688,N_4226);
nor U7550 (N_7550,N_2175,N_2960);
nand U7551 (N_7551,N_3219,N_1424);
and U7552 (N_7552,N_3057,N_3871);
nor U7553 (N_7553,N_4887,N_1407);
and U7554 (N_7554,N_4914,N_4106);
nand U7555 (N_7555,N_1999,N_660);
xor U7556 (N_7556,N_4991,N_2437);
and U7557 (N_7557,N_2348,N_3425);
nand U7558 (N_7558,N_501,N_721);
nor U7559 (N_7559,N_2909,N_835);
nor U7560 (N_7560,N_566,N_58);
or U7561 (N_7561,N_3530,N_1444);
and U7562 (N_7562,N_2491,N_375);
or U7563 (N_7563,N_551,N_770);
xor U7564 (N_7564,N_3073,N_1236);
nand U7565 (N_7565,N_1546,N_3860);
xor U7566 (N_7566,N_513,N_778);
nor U7567 (N_7567,N_4527,N_3195);
or U7568 (N_7568,N_4755,N_1020);
nand U7569 (N_7569,N_3263,N_2156);
or U7570 (N_7570,N_3388,N_4841);
xor U7571 (N_7571,N_301,N_3432);
xnor U7572 (N_7572,N_3476,N_2670);
and U7573 (N_7573,N_2044,N_2005);
nor U7574 (N_7574,N_4684,N_4123);
nand U7575 (N_7575,N_449,N_4286);
and U7576 (N_7576,N_961,N_290);
nor U7577 (N_7577,N_4498,N_574);
or U7578 (N_7578,N_1623,N_556);
xor U7579 (N_7579,N_3420,N_1822);
or U7580 (N_7580,N_3921,N_3597);
and U7581 (N_7581,N_3141,N_630);
or U7582 (N_7582,N_4208,N_961);
nand U7583 (N_7583,N_2733,N_1606);
and U7584 (N_7584,N_4701,N_4810);
nor U7585 (N_7585,N_2121,N_32);
and U7586 (N_7586,N_2524,N_3076);
nand U7587 (N_7587,N_4140,N_2743);
nor U7588 (N_7588,N_2832,N_4819);
nand U7589 (N_7589,N_3897,N_1887);
nor U7590 (N_7590,N_762,N_1264);
or U7591 (N_7591,N_2171,N_3094);
xnor U7592 (N_7592,N_4704,N_41);
or U7593 (N_7593,N_3775,N_1120);
nand U7594 (N_7594,N_2454,N_4593);
or U7595 (N_7595,N_3009,N_4408);
or U7596 (N_7596,N_2678,N_2939);
nand U7597 (N_7597,N_1545,N_1724);
nand U7598 (N_7598,N_2435,N_2989);
nor U7599 (N_7599,N_1161,N_1885);
or U7600 (N_7600,N_1014,N_3572);
nand U7601 (N_7601,N_2308,N_2876);
or U7602 (N_7602,N_3100,N_3017);
xor U7603 (N_7603,N_4991,N_3726);
nand U7604 (N_7604,N_2256,N_1795);
and U7605 (N_7605,N_3965,N_3515);
nor U7606 (N_7606,N_4069,N_4277);
or U7607 (N_7607,N_3700,N_3099);
or U7608 (N_7608,N_1357,N_4107);
and U7609 (N_7609,N_3990,N_4730);
nor U7610 (N_7610,N_2032,N_1087);
nand U7611 (N_7611,N_981,N_1652);
nand U7612 (N_7612,N_4041,N_4111);
and U7613 (N_7613,N_392,N_3941);
nor U7614 (N_7614,N_4366,N_1121);
nand U7615 (N_7615,N_1410,N_2063);
and U7616 (N_7616,N_2522,N_2709);
or U7617 (N_7617,N_2436,N_3492);
or U7618 (N_7618,N_3991,N_4983);
xor U7619 (N_7619,N_3230,N_2003);
nor U7620 (N_7620,N_4396,N_3517);
and U7621 (N_7621,N_3811,N_1781);
and U7622 (N_7622,N_4312,N_3319);
nor U7623 (N_7623,N_4574,N_3950);
or U7624 (N_7624,N_3065,N_2013);
and U7625 (N_7625,N_2894,N_1849);
and U7626 (N_7626,N_3243,N_4313);
and U7627 (N_7627,N_1937,N_10);
or U7628 (N_7628,N_4267,N_4711);
and U7629 (N_7629,N_1023,N_224);
and U7630 (N_7630,N_3647,N_2100);
or U7631 (N_7631,N_1835,N_4603);
and U7632 (N_7632,N_3801,N_948);
or U7633 (N_7633,N_4243,N_1054);
or U7634 (N_7634,N_441,N_4445);
and U7635 (N_7635,N_2226,N_1364);
or U7636 (N_7636,N_3659,N_1672);
nand U7637 (N_7637,N_2218,N_2962);
nor U7638 (N_7638,N_4912,N_2616);
nand U7639 (N_7639,N_4850,N_4366);
or U7640 (N_7640,N_449,N_2651);
nor U7641 (N_7641,N_3122,N_4767);
nand U7642 (N_7642,N_156,N_1615);
or U7643 (N_7643,N_623,N_4294);
nor U7644 (N_7644,N_578,N_113);
and U7645 (N_7645,N_1659,N_4467);
and U7646 (N_7646,N_993,N_4970);
xnor U7647 (N_7647,N_3645,N_2018);
and U7648 (N_7648,N_230,N_1628);
or U7649 (N_7649,N_4267,N_760);
nand U7650 (N_7650,N_2748,N_1879);
or U7651 (N_7651,N_2182,N_2718);
and U7652 (N_7652,N_2257,N_4603);
and U7653 (N_7653,N_3469,N_3546);
nor U7654 (N_7654,N_3698,N_1360);
or U7655 (N_7655,N_2470,N_4336);
nor U7656 (N_7656,N_2865,N_968);
or U7657 (N_7657,N_4899,N_1763);
nor U7658 (N_7658,N_4272,N_2996);
and U7659 (N_7659,N_45,N_2863);
nor U7660 (N_7660,N_3172,N_479);
nand U7661 (N_7661,N_1112,N_1828);
nand U7662 (N_7662,N_2916,N_917);
nor U7663 (N_7663,N_1094,N_4506);
nor U7664 (N_7664,N_4733,N_204);
nand U7665 (N_7665,N_3545,N_2778);
nand U7666 (N_7666,N_2044,N_4397);
nor U7667 (N_7667,N_3856,N_1117);
xnor U7668 (N_7668,N_2840,N_2192);
and U7669 (N_7669,N_515,N_1464);
and U7670 (N_7670,N_4372,N_1662);
and U7671 (N_7671,N_4660,N_535);
or U7672 (N_7672,N_218,N_3887);
nand U7673 (N_7673,N_3605,N_1487);
nor U7674 (N_7674,N_1946,N_4923);
nor U7675 (N_7675,N_600,N_348);
xor U7676 (N_7676,N_97,N_2108);
nor U7677 (N_7677,N_2317,N_2753);
and U7678 (N_7678,N_1079,N_4217);
and U7679 (N_7679,N_4420,N_3224);
and U7680 (N_7680,N_2729,N_4370);
nand U7681 (N_7681,N_4170,N_2766);
nand U7682 (N_7682,N_2548,N_4354);
and U7683 (N_7683,N_624,N_3670);
nand U7684 (N_7684,N_1387,N_4255);
or U7685 (N_7685,N_4529,N_1940);
nand U7686 (N_7686,N_3534,N_551);
nor U7687 (N_7687,N_1856,N_799);
nor U7688 (N_7688,N_24,N_4138);
or U7689 (N_7689,N_2847,N_1899);
nor U7690 (N_7690,N_3800,N_900);
xor U7691 (N_7691,N_3829,N_276);
and U7692 (N_7692,N_497,N_2107);
nand U7693 (N_7693,N_1434,N_3213);
or U7694 (N_7694,N_2632,N_2955);
nor U7695 (N_7695,N_1996,N_981);
nand U7696 (N_7696,N_9,N_3425);
xnor U7697 (N_7697,N_1641,N_4492);
nor U7698 (N_7698,N_908,N_2058);
and U7699 (N_7699,N_1211,N_781);
nand U7700 (N_7700,N_877,N_3710);
xor U7701 (N_7701,N_4889,N_893);
or U7702 (N_7702,N_3573,N_583);
nor U7703 (N_7703,N_4115,N_4207);
nor U7704 (N_7704,N_1215,N_2910);
xnor U7705 (N_7705,N_3714,N_960);
and U7706 (N_7706,N_1088,N_3821);
or U7707 (N_7707,N_79,N_4111);
nand U7708 (N_7708,N_173,N_587);
xor U7709 (N_7709,N_2793,N_3394);
nor U7710 (N_7710,N_1759,N_3157);
or U7711 (N_7711,N_4046,N_3297);
or U7712 (N_7712,N_3337,N_993);
and U7713 (N_7713,N_4862,N_3733);
and U7714 (N_7714,N_582,N_899);
or U7715 (N_7715,N_3476,N_1826);
xnor U7716 (N_7716,N_2462,N_1862);
nand U7717 (N_7717,N_3021,N_2956);
nand U7718 (N_7718,N_315,N_3374);
nor U7719 (N_7719,N_955,N_3033);
xor U7720 (N_7720,N_2040,N_1804);
nor U7721 (N_7721,N_4032,N_738);
and U7722 (N_7722,N_4459,N_2330);
nor U7723 (N_7723,N_44,N_2981);
and U7724 (N_7724,N_332,N_4034);
xor U7725 (N_7725,N_1438,N_4000);
or U7726 (N_7726,N_4699,N_2445);
nor U7727 (N_7727,N_417,N_522);
or U7728 (N_7728,N_2192,N_2066);
and U7729 (N_7729,N_2080,N_3742);
or U7730 (N_7730,N_3585,N_1803);
nand U7731 (N_7731,N_630,N_1986);
nand U7732 (N_7732,N_3150,N_3887);
and U7733 (N_7733,N_1058,N_3276);
and U7734 (N_7734,N_2466,N_3004);
nand U7735 (N_7735,N_4063,N_4054);
nor U7736 (N_7736,N_245,N_1914);
xnor U7737 (N_7737,N_1500,N_1173);
nor U7738 (N_7738,N_3147,N_3868);
nor U7739 (N_7739,N_1910,N_2094);
and U7740 (N_7740,N_396,N_4527);
or U7741 (N_7741,N_4141,N_441);
or U7742 (N_7742,N_1229,N_3212);
nand U7743 (N_7743,N_931,N_3078);
nor U7744 (N_7744,N_2511,N_349);
and U7745 (N_7745,N_3470,N_1153);
nand U7746 (N_7746,N_4583,N_1258);
xnor U7747 (N_7747,N_4146,N_2976);
nand U7748 (N_7748,N_3140,N_1422);
or U7749 (N_7749,N_3513,N_3776);
and U7750 (N_7750,N_3788,N_1149);
or U7751 (N_7751,N_782,N_4175);
or U7752 (N_7752,N_254,N_323);
or U7753 (N_7753,N_4847,N_2087);
or U7754 (N_7754,N_998,N_1532);
and U7755 (N_7755,N_1059,N_2404);
and U7756 (N_7756,N_2086,N_4244);
or U7757 (N_7757,N_1552,N_937);
xnor U7758 (N_7758,N_4902,N_3404);
nor U7759 (N_7759,N_1195,N_2283);
nor U7760 (N_7760,N_2704,N_2237);
xor U7761 (N_7761,N_738,N_374);
nor U7762 (N_7762,N_1560,N_4512);
nand U7763 (N_7763,N_3890,N_3013);
or U7764 (N_7764,N_1833,N_2110);
nand U7765 (N_7765,N_2426,N_4433);
or U7766 (N_7766,N_103,N_702);
nand U7767 (N_7767,N_3601,N_3404);
and U7768 (N_7768,N_2104,N_2741);
or U7769 (N_7769,N_3782,N_4783);
xor U7770 (N_7770,N_3451,N_2752);
nor U7771 (N_7771,N_4543,N_4424);
nor U7772 (N_7772,N_1382,N_1185);
or U7773 (N_7773,N_358,N_4552);
nor U7774 (N_7774,N_1077,N_2630);
xnor U7775 (N_7775,N_555,N_4493);
nand U7776 (N_7776,N_2363,N_1347);
and U7777 (N_7777,N_3393,N_3783);
nand U7778 (N_7778,N_6,N_1303);
nand U7779 (N_7779,N_3432,N_829);
nor U7780 (N_7780,N_685,N_4241);
nor U7781 (N_7781,N_4352,N_2110);
and U7782 (N_7782,N_2136,N_152);
nand U7783 (N_7783,N_505,N_2557);
nor U7784 (N_7784,N_2386,N_1830);
nand U7785 (N_7785,N_3258,N_2285);
nand U7786 (N_7786,N_2735,N_3046);
nand U7787 (N_7787,N_2130,N_4561);
nand U7788 (N_7788,N_886,N_2156);
or U7789 (N_7789,N_3743,N_414);
nand U7790 (N_7790,N_4755,N_3427);
nor U7791 (N_7791,N_3741,N_4302);
and U7792 (N_7792,N_4427,N_2650);
and U7793 (N_7793,N_3449,N_41);
and U7794 (N_7794,N_1756,N_673);
nand U7795 (N_7795,N_4547,N_402);
or U7796 (N_7796,N_56,N_4914);
nand U7797 (N_7797,N_2068,N_2715);
and U7798 (N_7798,N_2851,N_1599);
nand U7799 (N_7799,N_713,N_3682);
or U7800 (N_7800,N_4044,N_2172);
nor U7801 (N_7801,N_3127,N_2324);
nand U7802 (N_7802,N_782,N_1305);
nand U7803 (N_7803,N_42,N_1927);
nand U7804 (N_7804,N_3969,N_3775);
nor U7805 (N_7805,N_958,N_212);
or U7806 (N_7806,N_2472,N_2111);
and U7807 (N_7807,N_706,N_4821);
xnor U7808 (N_7808,N_4910,N_703);
and U7809 (N_7809,N_622,N_3813);
nand U7810 (N_7810,N_4945,N_2719);
nand U7811 (N_7811,N_4578,N_2224);
or U7812 (N_7812,N_662,N_2542);
nor U7813 (N_7813,N_1085,N_2502);
or U7814 (N_7814,N_2341,N_3789);
and U7815 (N_7815,N_4963,N_3163);
nand U7816 (N_7816,N_4611,N_1659);
and U7817 (N_7817,N_3335,N_1483);
nand U7818 (N_7818,N_584,N_2325);
nor U7819 (N_7819,N_3886,N_1582);
nand U7820 (N_7820,N_4153,N_1373);
nand U7821 (N_7821,N_3314,N_3429);
nand U7822 (N_7822,N_2330,N_3075);
or U7823 (N_7823,N_2,N_4289);
or U7824 (N_7824,N_3165,N_1312);
nor U7825 (N_7825,N_2959,N_2699);
and U7826 (N_7826,N_80,N_2281);
nand U7827 (N_7827,N_2687,N_2015);
nand U7828 (N_7828,N_528,N_2229);
or U7829 (N_7829,N_2095,N_381);
or U7830 (N_7830,N_2420,N_3119);
and U7831 (N_7831,N_4727,N_4561);
and U7832 (N_7832,N_3155,N_653);
nand U7833 (N_7833,N_4334,N_4546);
nand U7834 (N_7834,N_2517,N_4054);
or U7835 (N_7835,N_2532,N_2845);
xnor U7836 (N_7836,N_3902,N_2617);
xnor U7837 (N_7837,N_4189,N_4721);
and U7838 (N_7838,N_2511,N_1913);
nor U7839 (N_7839,N_1706,N_3258);
nor U7840 (N_7840,N_3189,N_559);
nand U7841 (N_7841,N_4731,N_3477);
xor U7842 (N_7842,N_2710,N_828);
nor U7843 (N_7843,N_2100,N_562);
or U7844 (N_7844,N_3793,N_3219);
and U7845 (N_7845,N_4616,N_3090);
xnor U7846 (N_7846,N_1469,N_2840);
and U7847 (N_7847,N_3925,N_1728);
nor U7848 (N_7848,N_994,N_2695);
or U7849 (N_7849,N_2886,N_1741);
nand U7850 (N_7850,N_2237,N_2760);
nand U7851 (N_7851,N_2472,N_1847);
or U7852 (N_7852,N_1629,N_4818);
nand U7853 (N_7853,N_2427,N_2289);
and U7854 (N_7854,N_2983,N_3350);
xor U7855 (N_7855,N_4299,N_4897);
xor U7856 (N_7856,N_4352,N_1813);
or U7857 (N_7857,N_733,N_4646);
nand U7858 (N_7858,N_2543,N_1231);
or U7859 (N_7859,N_1670,N_3968);
and U7860 (N_7860,N_528,N_1070);
or U7861 (N_7861,N_438,N_1622);
or U7862 (N_7862,N_1178,N_434);
or U7863 (N_7863,N_1727,N_1483);
xor U7864 (N_7864,N_44,N_1307);
xnor U7865 (N_7865,N_4881,N_2866);
nand U7866 (N_7866,N_2325,N_1022);
or U7867 (N_7867,N_2322,N_3277);
or U7868 (N_7868,N_3071,N_501);
and U7869 (N_7869,N_353,N_3646);
and U7870 (N_7870,N_1206,N_270);
and U7871 (N_7871,N_4118,N_4950);
or U7872 (N_7872,N_1752,N_4437);
or U7873 (N_7873,N_3494,N_4741);
or U7874 (N_7874,N_1181,N_354);
xnor U7875 (N_7875,N_463,N_4441);
and U7876 (N_7876,N_2534,N_1513);
and U7877 (N_7877,N_792,N_2071);
nand U7878 (N_7878,N_69,N_1610);
xor U7879 (N_7879,N_1416,N_4746);
nor U7880 (N_7880,N_2265,N_1596);
or U7881 (N_7881,N_392,N_3557);
and U7882 (N_7882,N_4181,N_3682);
nand U7883 (N_7883,N_4179,N_831);
xor U7884 (N_7884,N_4707,N_2730);
and U7885 (N_7885,N_1776,N_470);
xor U7886 (N_7886,N_1651,N_745);
or U7887 (N_7887,N_2767,N_1688);
and U7888 (N_7888,N_829,N_676);
or U7889 (N_7889,N_2393,N_4490);
or U7890 (N_7890,N_3992,N_3655);
xor U7891 (N_7891,N_292,N_2232);
or U7892 (N_7892,N_3511,N_1037);
and U7893 (N_7893,N_1259,N_3677);
or U7894 (N_7894,N_474,N_663);
nand U7895 (N_7895,N_4444,N_3672);
nor U7896 (N_7896,N_1606,N_4055);
or U7897 (N_7897,N_244,N_2923);
nor U7898 (N_7898,N_2551,N_653);
nand U7899 (N_7899,N_1297,N_4073);
nand U7900 (N_7900,N_4636,N_2527);
or U7901 (N_7901,N_589,N_2970);
and U7902 (N_7902,N_3903,N_1722);
and U7903 (N_7903,N_1734,N_3236);
and U7904 (N_7904,N_2972,N_3830);
nor U7905 (N_7905,N_1485,N_2183);
nor U7906 (N_7906,N_2787,N_2079);
nand U7907 (N_7907,N_1485,N_4025);
or U7908 (N_7908,N_1010,N_1839);
nand U7909 (N_7909,N_3663,N_407);
or U7910 (N_7910,N_4012,N_2396);
nand U7911 (N_7911,N_2246,N_3708);
xnor U7912 (N_7912,N_569,N_3941);
or U7913 (N_7913,N_4341,N_979);
nand U7914 (N_7914,N_1808,N_3092);
xor U7915 (N_7915,N_3355,N_1286);
and U7916 (N_7916,N_743,N_1164);
and U7917 (N_7917,N_3952,N_4909);
nor U7918 (N_7918,N_3729,N_3632);
nor U7919 (N_7919,N_3455,N_184);
and U7920 (N_7920,N_3196,N_1016);
and U7921 (N_7921,N_1060,N_2130);
xnor U7922 (N_7922,N_2277,N_3037);
and U7923 (N_7923,N_800,N_4415);
nor U7924 (N_7924,N_822,N_677);
or U7925 (N_7925,N_3577,N_1358);
nand U7926 (N_7926,N_3143,N_1550);
or U7927 (N_7927,N_1059,N_337);
or U7928 (N_7928,N_538,N_2164);
or U7929 (N_7929,N_3316,N_3100);
or U7930 (N_7930,N_1696,N_332);
and U7931 (N_7931,N_1369,N_4955);
nand U7932 (N_7932,N_1082,N_830);
and U7933 (N_7933,N_1994,N_2164);
and U7934 (N_7934,N_168,N_1286);
and U7935 (N_7935,N_4490,N_685);
and U7936 (N_7936,N_4738,N_2431);
nand U7937 (N_7937,N_2302,N_299);
nor U7938 (N_7938,N_1419,N_380);
and U7939 (N_7939,N_964,N_1884);
or U7940 (N_7940,N_869,N_1487);
and U7941 (N_7941,N_1261,N_668);
and U7942 (N_7942,N_4253,N_4132);
and U7943 (N_7943,N_547,N_3508);
nor U7944 (N_7944,N_4666,N_517);
and U7945 (N_7945,N_1438,N_4678);
or U7946 (N_7946,N_555,N_4683);
and U7947 (N_7947,N_1344,N_2366);
nand U7948 (N_7948,N_4180,N_284);
xor U7949 (N_7949,N_4061,N_2187);
and U7950 (N_7950,N_3063,N_66);
nand U7951 (N_7951,N_342,N_1043);
or U7952 (N_7952,N_357,N_68);
and U7953 (N_7953,N_812,N_4332);
nand U7954 (N_7954,N_843,N_4768);
nor U7955 (N_7955,N_4803,N_4917);
nor U7956 (N_7956,N_782,N_3916);
or U7957 (N_7957,N_522,N_2339);
xor U7958 (N_7958,N_3142,N_3379);
and U7959 (N_7959,N_4823,N_2158);
and U7960 (N_7960,N_3205,N_1590);
nand U7961 (N_7961,N_2427,N_4397);
nand U7962 (N_7962,N_1147,N_136);
nand U7963 (N_7963,N_4864,N_2484);
nand U7964 (N_7964,N_2969,N_1965);
nor U7965 (N_7965,N_2410,N_4732);
xor U7966 (N_7966,N_1640,N_285);
or U7967 (N_7967,N_1957,N_3294);
or U7968 (N_7968,N_3335,N_4237);
or U7969 (N_7969,N_4827,N_3412);
nand U7970 (N_7970,N_4621,N_4987);
or U7971 (N_7971,N_1123,N_3178);
nor U7972 (N_7972,N_1745,N_479);
or U7973 (N_7973,N_2416,N_4578);
and U7974 (N_7974,N_1873,N_236);
and U7975 (N_7975,N_841,N_2860);
and U7976 (N_7976,N_3489,N_1089);
and U7977 (N_7977,N_3996,N_4443);
and U7978 (N_7978,N_1956,N_1825);
or U7979 (N_7979,N_4516,N_2268);
and U7980 (N_7980,N_4928,N_1956);
or U7981 (N_7981,N_3156,N_542);
or U7982 (N_7982,N_2157,N_2680);
nor U7983 (N_7983,N_157,N_2480);
and U7984 (N_7984,N_3212,N_2739);
xnor U7985 (N_7985,N_1554,N_688);
nor U7986 (N_7986,N_4420,N_1417);
and U7987 (N_7987,N_3572,N_3481);
nor U7988 (N_7988,N_677,N_4630);
nor U7989 (N_7989,N_12,N_3856);
or U7990 (N_7990,N_2267,N_1824);
nor U7991 (N_7991,N_2042,N_4617);
nand U7992 (N_7992,N_1661,N_4201);
and U7993 (N_7993,N_2119,N_1988);
xnor U7994 (N_7994,N_978,N_2873);
nor U7995 (N_7995,N_4201,N_3352);
and U7996 (N_7996,N_2180,N_4051);
xnor U7997 (N_7997,N_2963,N_4748);
nand U7998 (N_7998,N_4103,N_4601);
nor U7999 (N_7999,N_1502,N_407);
or U8000 (N_8000,N_400,N_2500);
nand U8001 (N_8001,N_428,N_2074);
or U8002 (N_8002,N_2322,N_2816);
or U8003 (N_8003,N_2234,N_2764);
xnor U8004 (N_8004,N_714,N_432);
or U8005 (N_8005,N_2693,N_4472);
or U8006 (N_8006,N_3667,N_354);
and U8007 (N_8007,N_2660,N_2022);
or U8008 (N_8008,N_938,N_4554);
xnor U8009 (N_8009,N_2895,N_3250);
nand U8010 (N_8010,N_4455,N_2704);
nor U8011 (N_8011,N_4619,N_1238);
xnor U8012 (N_8012,N_262,N_2804);
nand U8013 (N_8013,N_4124,N_2954);
xor U8014 (N_8014,N_2779,N_2021);
and U8015 (N_8015,N_2415,N_103);
or U8016 (N_8016,N_2403,N_4736);
nor U8017 (N_8017,N_4743,N_3225);
xnor U8018 (N_8018,N_4727,N_2607);
and U8019 (N_8019,N_4215,N_2697);
or U8020 (N_8020,N_1735,N_586);
or U8021 (N_8021,N_3134,N_586);
or U8022 (N_8022,N_2296,N_893);
or U8023 (N_8023,N_2187,N_3498);
and U8024 (N_8024,N_375,N_4900);
xnor U8025 (N_8025,N_3604,N_4353);
and U8026 (N_8026,N_2528,N_432);
nor U8027 (N_8027,N_998,N_1093);
nor U8028 (N_8028,N_2268,N_1881);
nor U8029 (N_8029,N_211,N_1252);
or U8030 (N_8030,N_2995,N_4036);
xnor U8031 (N_8031,N_1333,N_4804);
nor U8032 (N_8032,N_3513,N_4839);
and U8033 (N_8033,N_3288,N_2092);
and U8034 (N_8034,N_3029,N_1920);
nor U8035 (N_8035,N_47,N_3367);
nand U8036 (N_8036,N_478,N_2899);
nor U8037 (N_8037,N_1183,N_3630);
or U8038 (N_8038,N_2515,N_1181);
nand U8039 (N_8039,N_976,N_1480);
or U8040 (N_8040,N_3205,N_2844);
nand U8041 (N_8041,N_688,N_1858);
nor U8042 (N_8042,N_2610,N_3620);
or U8043 (N_8043,N_3435,N_1473);
and U8044 (N_8044,N_2534,N_4443);
nor U8045 (N_8045,N_4341,N_224);
and U8046 (N_8046,N_3610,N_243);
and U8047 (N_8047,N_937,N_2362);
nor U8048 (N_8048,N_514,N_3527);
nor U8049 (N_8049,N_3184,N_1975);
or U8050 (N_8050,N_623,N_1807);
and U8051 (N_8051,N_2303,N_151);
nor U8052 (N_8052,N_807,N_3678);
nor U8053 (N_8053,N_4187,N_4065);
nand U8054 (N_8054,N_3904,N_3725);
or U8055 (N_8055,N_2850,N_1398);
nor U8056 (N_8056,N_1225,N_4676);
and U8057 (N_8057,N_1957,N_3328);
and U8058 (N_8058,N_1702,N_416);
nor U8059 (N_8059,N_4688,N_3746);
nand U8060 (N_8060,N_635,N_713);
xor U8061 (N_8061,N_491,N_2409);
nor U8062 (N_8062,N_4795,N_731);
or U8063 (N_8063,N_4182,N_1874);
or U8064 (N_8064,N_3865,N_4394);
xor U8065 (N_8065,N_2319,N_851);
xnor U8066 (N_8066,N_2548,N_1495);
nor U8067 (N_8067,N_3656,N_2747);
and U8068 (N_8068,N_3601,N_1925);
xor U8069 (N_8069,N_1450,N_4837);
nor U8070 (N_8070,N_3479,N_1884);
and U8071 (N_8071,N_1138,N_1282);
xor U8072 (N_8072,N_3879,N_1830);
xnor U8073 (N_8073,N_372,N_4610);
nor U8074 (N_8074,N_3988,N_2607);
and U8075 (N_8075,N_4225,N_2349);
nand U8076 (N_8076,N_1109,N_3619);
xnor U8077 (N_8077,N_1868,N_4408);
or U8078 (N_8078,N_3293,N_3831);
nor U8079 (N_8079,N_370,N_3681);
nand U8080 (N_8080,N_2920,N_960);
nor U8081 (N_8081,N_1590,N_2880);
or U8082 (N_8082,N_699,N_4199);
and U8083 (N_8083,N_1536,N_2957);
nand U8084 (N_8084,N_244,N_930);
or U8085 (N_8085,N_1998,N_2638);
nand U8086 (N_8086,N_748,N_4640);
or U8087 (N_8087,N_1471,N_2109);
or U8088 (N_8088,N_331,N_844);
nor U8089 (N_8089,N_143,N_464);
xnor U8090 (N_8090,N_3949,N_970);
xor U8091 (N_8091,N_2809,N_879);
nor U8092 (N_8092,N_4197,N_2781);
or U8093 (N_8093,N_4155,N_4791);
or U8094 (N_8094,N_174,N_3865);
and U8095 (N_8095,N_4249,N_2865);
nand U8096 (N_8096,N_189,N_2092);
and U8097 (N_8097,N_3024,N_4778);
or U8098 (N_8098,N_1359,N_2991);
and U8099 (N_8099,N_1973,N_2366);
or U8100 (N_8100,N_4733,N_11);
and U8101 (N_8101,N_793,N_2552);
nor U8102 (N_8102,N_1726,N_2778);
and U8103 (N_8103,N_2958,N_1329);
nor U8104 (N_8104,N_1201,N_1814);
nand U8105 (N_8105,N_2756,N_2458);
and U8106 (N_8106,N_3327,N_4870);
xnor U8107 (N_8107,N_1205,N_3601);
nor U8108 (N_8108,N_1391,N_1573);
nor U8109 (N_8109,N_884,N_55);
and U8110 (N_8110,N_2467,N_2197);
or U8111 (N_8111,N_1047,N_3742);
nor U8112 (N_8112,N_3212,N_1260);
nand U8113 (N_8113,N_3013,N_4368);
and U8114 (N_8114,N_192,N_715);
and U8115 (N_8115,N_3229,N_1060);
and U8116 (N_8116,N_143,N_223);
or U8117 (N_8117,N_3253,N_1015);
or U8118 (N_8118,N_1976,N_4935);
nand U8119 (N_8119,N_2919,N_1544);
nand U8120 (N_8120,N_26,N_1372);
or U8121 (N_8121,N_3497,N_2781);
nand U8122 (N_8122,N_411,N_3682);
nand U8123 (N_8123,N_1815,N_2826);
and U8124 (N_8124,N_1134,N_1598);
and U8125 (N_8125,N_41,N_2129);
or U8126 (N_8126,N_1249,N_1734);
or U8127 (N_8127,N_2003,N_4725);
nand U8128 (N_8128,N_931,N_2538);
nand U8129 (N_8129,N_844,N_3437);
and U8130 (N_8130,N_4843,N_3102);
or U8131 (N_8131,N_2158,N_4242);
or U8132 (N_8132,N_4850,N_3658);
xnor U8133 (N_8133,N_2248,N_1886);
or U8134 (N_8134,N_4078,N_2435);
nand U8135 (N_8135,N_2946,N_4659);
nand U8136 (N_8136,N_295,N_2171);
nor U8137 (N_8137,N_3938,N_1925);
nand U8138 (N_8138,N_2529,N_1666);
or U8139 (N_8139,N_3525,N_2529);
nand U8140 (N_8140,N_1118,N_2235);
and U8141 (N_8141,N_319,N_4401);
or U8142 (N_8142,N_2356,N_3536);
nor U8143 (N_8143,N_2706,N_590);
nor U8144 (N_8144,N_2286,N_1988);
and U8145 (N_8145,N_29,N_2239);
xnor U8146 (N_8146,N_4254,N_758);
and U8147 (N_8147,N_3691,N_2946);
xnor U8148 (N_8148,N_660,N_4582);
nand U8149 (N_8149,N_2777,N_3073);
nand U8150 (N_8150,N_2578,N_4114);
and U8151 (N_8151,N_2804,N_291);
nand U8152 (N_8152,N_1500,N_3706);
or U8153 (N_8153,N_3426,N_4013);
and U8154 (N_8154,N_1456,N_4087);
nor U8155 (N_8155,N_490,N_2319);
or U8156 (N_8156,N_3160,N_2961);
or U8157 (N_8157,N_1566,N_1773);
xnor U8158 (N_8158,N_2399,N_3410);
or U8159 (N_8159,N_2685,N_4161);
or U8160 (N_8160,N_1734,N_3448);
and U8161 (N_8161,N_4792,N_62);
nor U8162 (N_8162,N_2904,N_2432);
or U8163 (N_8163,N_174,N_2703);
or U8164 (N_8164,N_4117,N_2101);
or U8165 (N_8165,N_636,N_3403);
or U8166 (N_8166,N_1409,N_2811);
or U8167 (N_8167,N_3890,N_2113);
nand U8168 (N_8168,N_4815,N_4991);
xor U8169 (N_8169,N_792,N_3110);
and U8170 (N_8170,N_4998,N_1056);
and U8171 (N_8171,N_1801,N_3267);
nor U8172 (N_8172,N_3835,N_3963);
or U8173 (N_8173,N_4157,N_4356);
nand U8174 (N_8174,N_2556,N_249);
xnor U8175 (N_8175,N_3487,N_4201);
and U8176 (N_8176,N_4388,N_3576);
nor U8177 (N_8177,N_2450,N_1681);
nor U8178 (N_8178,N_3889,N_55);
and U8179 (N_8179,N_3558,N_4602);
or U8180 (N_8180,N_3599,N_2929);
nor U8181 (N_8181,N_1981,N_1658);
and U8182 (N_8182,N_4915,N_3811);
xnor U8183 (N_8183,N_1114,N_265);
nand U8184 (N_8184,N_747,N_1117);
nand U8185 (N_8185,N_295,N_969);
nand U8186 (N_8186,N_526,N_2401);
or U8187 (N_8187,N_271,N_3090);
nand U8188 (N_8188,N_2456,N_4440);
xnor U8189 (N_8189,N_4022,N_1909);
nor U8190 (N_8190,N_4289,N_4586);
nor U8191 (N_8191,N_3750,N_3111);
nand U8192 (N_8192,N_761,N_2075);
nand U8193 (N_8193,N_2248,N_1287);
nand U8194 (N_8194,N_81,N_3845);
nand U8195 (N_8195,N_1425,N_997);
or U8196 (N_8196,N_1087,N_356);
nand U8197 (N_8197,N_3380,N_4496);
xnor U8198 (N_8198,N_2033,N_2848);
and U8199 (N_8199,N_159,N_558);
and U8200 (N_8200,N_240,N_3270);
and U8201 (N_8201,N_1070,N_369);
nor U8202 (N_8202,N_3220,N_4595);
or U8203 (N_8203,N_3774,N_773);
nor U8204 (N_8204,N_684,N_534);
nor U8205 (N_8205,N_2820,N_4061);
or U8206 (N_8206,N_1639,N_3572);
nand U8207 (N_8207,N_2822,N_917);
nor U8208 (N_8208,N_4328,N_4100);
or U8209 (N_8209,N_2703,N_3114);
and U8210 (N_8210,N_1147,N_4616);
nand U8211 (N_8211,N_1367,N_2392);
and U8212 (N_8212,N_3913,N_3614);
nor U8213 (N_8213,N_2371,N_3059);
nor U8214 (N_8214,N_964,N_2615);
and U8215 (N_8215,N_850,N_3226);
nand U8216 (N_8216,N_2498,N_2188);
nand U8217 (N_8217,N_4253,N_2036);
and U8218 (N_8218,N_3688,N_2104);
nand U8219 (N_8219,N_156,N_4837);
xnor U8220 (N_8220,N_4109,N_3771);
and U8221 (N_8221,N_4248,N_1588);
and U8222 (N_8222,N_446,N_2169);
nand U8223 (N_8223,N_71,N_1929);
or U8224 (N_8224,N_2,N_3536);
xnor U8225 (N_8225,N_4063,N_3082);
nand U8226 (N_8226,N_2269,N_4865);
nor U8227 (N_8227,N_2204,N_1511);
xor U8228 (N_8228,N_254,N_2230);
or U8229 (N_8229,N_2543,N_2673);
nand U8230 (N_8230,N_4882,N_4845);
xnor U8231 (N_8231,N_3284,N_1561);
xnor U8232 (N_8232,N_3475,N_1062);
or U8233 (N_8233,N_567,N_2101);
or U8234 (N_8234,N_929,N_1541);
xor U8235 (N_8235,N_1755,N_2298);
and U8236 (N_8236,N_349,N_2579);
xnor U8237 (N_8237,N_2356,N_1539);
nor U8238 (N_8238,N_1879,N_507);
nand U8239 (N_8239,N_2237,N_3404);
nor U8240 (N_8240,N_1634,N_384);
or U8241 (N_8241,N_2403,N_2830);
and U8242 (N_8242,N_1106,N_2713);
or U8243 (N_8243,N_1436,N_3014);
or U8244 (N_8244,N_3409,N_2104);
nor U8245 (N_8245,N_2391,N_1555);
xnor U8246 (N_8246,N_3547,N_517);
nor U8247 (N_8247,N_4463,N_3452);
nand U8248 (N_8248,N_2565,N_199);
nand U8249 (N_8249,N_676,N_2691);
and U8250 (N_8250,N_1552,N_3316);
and U8251 (N_8251,N_1437,N_4838);
nor U8252 (N_8252,N_117,N_1624);
nand U8253 (N_8253,N_1107,N_4590);
and U8254 (N_8254,N_4378,N_1760);
nor U8255 (N_8255,N_3868,N_550);
nand U8256 (N_8256,N_3958,N_412);
nand U8257 (N_8257,N_1769,N_1712);
or U8258 (N_8258,N_3677,N_4522);
and U8259 (N_8259,N_4479,N_1392);
nor U8260 (N_8260,N_3834,N_4904);
and U8261 (N_8261,N_4979,N_3558);
and U8262 (N_8262,N_1902,N_1368);
or U8263 (N_8263,N_3757,N_379);
nand U8264 (N_8264,N_2179,N_406);
or U8265 (N_8265,N_2323,N_428);
nor U8266 (N_8266,N_1510,N_3501);
or U8267 (N_8267,N_1809,N_2476);
xnor U8268 (N_8268,N_509,N_4161);
nand U8269 (N_8269,N_2829,N_3841);
nor U8270 (N_8270,N_3779,N_4908);
and U8271 (N_8271,N_2048,N_220);
nand U8272 (N_8272,N_461,N_4278);
and U8273 (N_8273,N_2412,N_4909);
and U8274 (N_8274,N_1384,N_2923);
or U8275 (N_8275,N_3554,N_1047);
nand U8276 (N_8276,N_3949,N_629);
and U8277 (N_8277,N_1990,N_2098);
nand U8278 (N_8278,N_1146,N_1365);
or U8279 (N_8279,N_2148,N_2431);
nor U8280 (N_8280,N_1269,N_3538);
xor U8281 (N_8281,N_3704,N_178);
and U8282 (N_8282,N_3916,N_3822);
nand U8283 (N_8283,N_2947,N_2830);
nand U8284 (N_8284,N_1172,N_4912);
xor U8285 (N_8285,N_4420,N_842);
nand U8286 (N_8286,N_237,N_4928);
and U8287 (N_8287,N_1583,N_4406);
or U8288 (N_8288,N_4648,N_4240);
and U8289 (N_8289,N_2966,N_4659);
nand U8290 (N_8290,N_444,N_3651);
nand U8291 (N_8291,N_1121,N_1590);
nand U8292 (N_8292,N_2837,N_4057);
or U8293 (N_8293,N_4721,N_785);
nor U8294 (N_8294,N_345,N_2041);
and U8295 (N_8295,N_3423,N_2543);
and U8296 (N_8296,N_2775,N_773);
xnor U8297 (N_8297,N_2621,N_920);
xor U8298 (N_8298,N_2572,N_3753);
and U8299 (N_8299,N_142,N_3585);
and U8300 (N_8300,N_4152,N_3863);
and U8301 (N_8301,N_2160,N_2740);
nor U8302 (N_8302,N_1411,N_2189);
or U8303 (N_8303,N_3016,N_4100);
or U8304 (N_8304,N_1194,N_655);
nor U8305 (N_8305,N_3209,N_4186);
nand U8306 (N_8306,N_1982,N_762);
nand U8307 (N_8307,N_3091,N_2819);
nor U8308 (N_8308,N_4950,N_3534);
nand U8309 (N_8309,N_2660,N_1156);
nand U8310 (N_8310,N_846,N_257);
nor U8311 (N_8311,N_3919,N_1253);
nand U8312 (N_8312,N_2976,N_4292);
and U8313 (N_8313,N_1187,N_1258);
or U8314 (N_8314,N_3561,N_2333);
or U8315 (N_8315,N_3296,N_3743);
and U8316 (N_8316,N_4305,N_2073);
or U8317 (N_8317,N_88,N_2935);
or U8318 (N_8318,N_512,N_1319);
xnor U8319 (N_8319,N_3672,N_4857);
nand U8320 (N_8320,N_3486,N_3976);
nand U8321 (N_8321,N_4573,N_3726);
or U8322 (N_8322,N_2841,N_4822);
or U8323 (N_8323,N_1599,N_2733);
nand U8324 (N_8324,N_4325,N_3415);
nor U8325 (N_8325,N_2108,N_1674);
and U8326 (N_8326,N_2497,N_4908);
and U8327 (N_8327,N_3702,N_3399);
xnor U8328 (N_8328,N_4801,N_1418);
or U8329 (N_8329,N_4240,N_1098);
xor U8330 (N_8330,N_2213,N_2082);
and U8331 (N_8331,N_4780,N_3092);
and U8332 (N_8332,N_2141,N_4647);
and U8333 (N_8333,N_571,N_2189);
nand U8334 (N_8334,N_2198,N_2003);
nand U8335 (N_8335,N_2277,N_1191);
xor U8336 (N_8336,N_85,N_904);
xnor U8337 (N_8337,N_1614,N_2787);
or U8338 (N_8338,N_2682,N_1042);
or U8339 (N_8339,N_1624,N_2189);
and U8340 (N_8340,N_2247,N_1930);
and U8341 (N_8341,N_1349,N_4996);
or U8342 (N_8342,N_2857,N_118);
or U8343 (N_8343,N_3551,N_462);
nor U8344 (N_8344,N_1796,N_952);
nor U8345 (N_8345,N_3086,N_827);
nor U8346 (N_8346,N_1126,N_2664);
and U8347 (N_8347,N_4122,N_967);
nor U8348 (N_8348,N_4532,N_1175);
or U8349 (N_8349,N_1443,N_1606);
nand U8350 (N_8350,N_4664,N_563);
nand U8351 (N_8351,N_1531,N_1769);
and U8352 (N_8352,N_1885,N_3730);
nor U8353 (N_8353,N_4387,N_1514);
xor U8354 (N_8354,N_2349,N_600);
xnor U8355 (N_8355,N_1848,N_811);
nand U8356 (N_8356,N_3888,N_3681);
xor U8357 (N_8357,N_3969,N_3311);
nand U8358 (N_8358,N_3739,N_4698);
nor U8359 (N_8359,N_3842,N_4277);
nor U8360 (N_8360,N_3948,N_4515);
and U8361 (N_8361,N_2053,N_324);
nor U8362 (N_8362,N_4369,N_3277);
or U8363 (N_8363,N_918,N_4653);
xnor U8364 (N_8364,N_4438,N_2935);
and U8365 (N_8365,N_104,N_2672);
nor U8366 (N_8366,N_3384,N_79);
xor U8367 (N_8367,N_1566,N_1798);
and U8368 (N_8368,N_2716,N_804);
nor U8369 (N_8369,N_3740,N_920);
or U8370 (N_8370,N_1410,N_1288);
or U8371 (N_8371,N_1782,N_2930);
and U8372 (N_8372,N_150,N_2201);
or U8373 (N_8373,N_4486,N_4925);
nor U8374 (N_8374,N_4709,N_679);
nor U8375 (N_8375,N_2396,N_1958);
and U8376 (N_8376,N_882,N_4273);
and U8377 (N_8377,N_1962,N_4751);
nand U8378 (N_8378,N_2432,N_4648);
nand U8379 (N_8379,N_2974,N_2728);
nand U8380 (N_8380,N_4462,N_3958);
nor U8381 (N_8381,N_347,N_3743);
and U8382 (N_8382,N_2857,N_3580);
or U8383 (N_8383,N_3366,N_4824);
nand U8384 (N_8384,N_3012,N_2703);
nand U8385 (N_8385,N_2309,N_3835);
and U8386 (N_8386,N_4064,N_2969);
or U8387 (N_8387,N_1689,N_4101);
nand U8388 (N_8388,N_4932,N_875);
nand U8389 (N_8389,N_2656,N_896);
or U8390 (N_8390,N_4732,N_3346);
nand U8391 (N_8391,N_101,N_4301);
and U8392 (N_8392,N_3667,N_4331);
or U8393 (N_8393,N_3295,N_758);
or U8394 (N_8394,N_4000,N_4986);
and U8395 (N_8395,N_1736,N_380);
and U8396 (N_8396,N_47,N_4086);
xnor U8397 (N_8397,N_1053,N_1258);
and U8398 (N_8398,N_1062,N_291);
nor U8399 (N_8399,N_4617,N_4787);
and U8400 (N_8400,N_2243,N_4256);
and U8401 (N_8401,N_4793,N_4800);
or U8402 (N_8402,N_4742,N_3576);
nand U8403 (N_8403,N_1014,N_3803);
nand U8404 (N_8404,N_3480,N_3242);
and U8405 (N_8405,N_2224,N_585);
nand U8406 (N_8406,N_3484,N_1159);
nor U8407 (N_8407,N_940,N_3821);
or U8408 (N_8408,N_1166,N_1837);
nor U8409 (N_8409,N_1749,N_2510);
nor U8410 (N_8410,N_3543,N_1817);
or U8411 (N_8411,N_4562,N_215);
nand U8412 (N_8412,N_2088,N_1942);
nor U8413 (N_8413,N_1401,N_2480);
and U8414 (N_8414,N_4987,N_3872);
xor U8415 (N_8415,N_4039,N_2815);
xnor U8416 (N_8416,N_3411,N_906);
nor U8417 (N_8417,N_865,N_3845);
nand U8418 (N_8418,N_2239,N_404);
nor U8419 (N_8419,N_2665,N_2860);
or U8420 (N_8420,N_3645,N_2995);
nand U8421 (N_8421,N_2508,N_4505);
xor U8422 (N_8422,N_3459,N_2191);
nand U8423 (N_8423,N_744,N_1688);
nand U8424 (N_8424,N_1510,N_1024);
nor U8425 (N_8425,N_253,N_1090);
or U8426 (N_8426,N_4921,N_4288);
nand U8427 (N_8427,N_1930,N_4198);
nand U8428 (N_8428,N_1201,N_917);
and U8429 (N_8429,N_2692,N_3749);
or U8430 (N_8430,N_3864,N_2581);
xor U8431 (N_8431,N_3606,N_4792);
or U8432 (N_8432,N_212,N_3063);
nor U8433 (N_8433,N_3345,N_4961);
xnor U8434 (N_8434,N_1293,N_4162);
or U8435 (N_8435,N_4288,N_1415);
and U8436 (N_8436,N_3056,N_2607);
nor U8437 (N_8437,N_4602,N_4503);
and U8438 (N_8438,N_4831,N_1223);
nand U8439 (N_8439,N_2451,N_2477);
or U8440 (N_8440,N_4192,N_1013);
nand U8441 (N_8441,N_2744,N_2997);
nand U8442 (N_8442,N_2036,N_4236);
nor U8443 (N_8443,N_819,N_2307);
and U8444 (N_8444,N_4364,N_2571);
and U8445 (N_8445,N_2046,N_949);
or U8446 (N_8446,N_3769,N_1056);
nor U8447 (N_8447,N_3508,N_3998);
and U8448 (N_8448,N_1649,N_2948);
xnor U8449 (N_8449,N_4485,N_3045);
and U8450 (N_8450,N_30,N_1516);
nor U8451 (N_8451,N_2264,N_1543);
or U8452 (N_8452,N_396,N_662);
and U8453 (N_8453,N_2411,N_2913);
nor U8454 (N_8454,N_1970,N_695);
or U8455 (N_8455,N_3033,N_1187);
nand U8456 (N_8456,N_3294,N_4592);
nor U8457 (N_8457,N_2320,N_4327);
nand U8458 (N_8458,N_385,N_4343);
nand U8459 (N_8459,N_4246,N_1503);
or U8460 (N_8460,N_1469,N_4069);
nor U8461 (N_8461,N_3240,N_4598);
nor U8462 (N_8462,N_2819,N_3738);
nand U8463 (N_8463,N_1380,N_4616);
nand U8464 (N_8464,N_4599,N_4305);
and U8465 (N_8465,N_490,N_2522);
nor U8466 (N_8466,N_4453,N_1301);
or U8467 (N_8467,N_264,N_325);
nand U8468 (N_8468,N_4337,N_2449);
or U8469 (N_8469,N_660,N_1786);
or U8470 (N_8470,N_1082,N_3331);
nor U8471 (N_8471,N_1016,N_4827);
nor U8472 (N_8472,N_1149,N_2332);
nor U8473 (N_8473,N_4928,N_4292);
or U8474 (N_8474,N_2249,N_3030);
and U8475 (N_8475,N_2320,N_759);
or U8476 (N_8476,N_2314,N_2956);
or U8477 (N_8477,N_3813,N_4777);
nand U8478 (N_8478,N_236,N_481);
or U8479 (N_8479,N_3559,N_619);
nor U8480 (N_8480,N_4341,N_3159);
and U8481 (N_8481,N_2285,N_3822);
or U8482 (N_8482,N_4611,N_33);
nor U8483 (N_8483,N_1761,N_47);
and U8484 (N_8484,N_113,N_1457);
nor U8485 (N_8485,N_3925,N_3825);
or U8486 (N_8486,N_998,N_4015);
or U8487 (N_8487,N_4264,N_935);
nand U8488 (N_8488,N_1044,N_1715);
and U8489 (N_8489,N_186,N_4253);
xnor U8490 (N_8490,N_617,N_1015);
xnor U8491 (N_8491,N_2487,N_2658);
nor U8492 (N_8492,N_4785,N_1700);
and U8493 (N_8493,N_4752,N_1312);
and U8494 (N_8494,N_530,N_4847);
and U8495 (N_8495,N_2437,N_792);
or U8496 (N_8496,N_2198,N_1974);
and U8497 (N_8497,N_3727,N_2918);
nand U8498 (N_8498,N_1304,N_1158);
nand U8499 (N_8499,N_2028,N_1484);
nor U8500 (N_8500,N_1874,N_216);
nand U8501 (N_8501,N_691,N_898);
nand U8502 (N_8502,N_2534,N_4141);
and U8503 (N_8503,N_288,N_3516);
nand U8504 (N_8504,N_2363,N_78);
nor U8505 (N_8505,N_3218,N_1494);
xnor U8506 (N_8506,N_2798,N_2866);
or U8507 (N_8507,N_1280,N_1541);
nand U8508 (N_8508,N_791,N_2541);
nor U8509 (N_8509,N_1195,N_3657);
and U8510 (N_8510,N_2816,N_2039);
or U8511 (N_8511,N_772,N_722);
nor U8512 (N_8512,N_2414,N_144);
or U8513 (N_8513,N_1763,N_875);
and U8514 (N_8514,N_2635,N_633);
or U8515 (N_8515,N_593,N_2067);
xnor U8516 (N_8516,N_2366,N_2158);
nor U8517 (N_8517,N_3187,N_2548);
or U8518 (N_8518,N_1793,N_4395);
nor U8519 (N_8519,N_2156,N_1812);
xnor U8520 (N_8520,N_3598,N_3653);
nand U8521 (N_8521,N_1599,N_4543);
and U8522 (N_8522,N_427,N_4795);
nand U8523 (N_8523,N_339,N_1317);
or U8524 (N_8524,N_1060,N_2173);
nand U8525 (N_8525,N_2821,N_883);
and U8526 (N_8526,N_2025,N_4247);
or U8527 (N_8527,N_2797,N_63);
nor U8528 (N_8528,N_4425,N_1370);
xnor U8529 (N_8529,N_4464,N_2966);
xnor U8530 (N_8530,N_708,N_3965);
xor U8531 (N_8531,N_961,N_1345);
or U8532 (N_8532,N_3764,N_3457);
and U8533 (N_8533,N_3984,N_3116);
and U8534 (N_8534,N_1815,N_3593);
or U8535 (N_8535,N_2457,N_833);
xnor U8536 (N_8536,N_3678,N_853);
and U8537 (N_8537,N_328,N_1101);
nand U8538 (N_8538,N_3698,N_1080);
nand U8539 (N_8539,N_3403,N_4497);
or U8540 (N_8540,N_1189,N_4360);
nor U8541 (N_8541,N_4447,N_2209);
xnor U8542 (N_8542,N_1625,N_210);
and U8543 (N_8543,N_1818,N_399);
or U8544 (N_8544,N_668,N_3153);
nor U8545 (N_8545,N_1878,N_1622);
xnor U8546 (N_8546,N_4894,N_1240);
or U8547 (N_8547,N_1542,N_3369);
or U8548 (N_8548,N_4179,N_2777);
or U8549 (N_8549,N_3642,N_773);
xor U8550 (N_8550,N_3,N_3260);
xor U8551 (N_8551,N_3603,N_2820);
or U8552 (N_8552,N_4108,N_84);
and U8553 (N_8553,N_3403,N_3113);
xnor U8554 (N_8554,N_3719,N_702);
nand U8555 (N_8555,N_1451,N_3182);
or U8556 (N_8556,N_4106,N_3537);
nor U8557 (N_8557,N_1776,N_975);
or U8558 (N_8558,N_1306,N_647);
nor U8559 (N_8559,N_1953,N_193);
nor U8560 (N_8560,N_4668,N_1319);
and U8561 (N_8561,N_47,N_796);
or U8562 (N_8562,N_3555,N_2539);
or U8563 (N_8563,N_1308,N_4509);
and U8564 (N_8564,N_562,N_2194);
or U8565 (N_8565,N_4859,N_1281);
or U8566 (N_8566,N_4082,N_2964);
or U8567 (N_8567,N_3152,N_1187);
xor U8568 (N_8568,N_4492,N_2613);
nand U8569 (N_8569,N_184,N_3115);
and U8570 (N_8570,N_2026,N_4115);
nor U8571 (N_8571,N_4307,N_941);
and U8572 (N_8572,N_4123,N_4647);
nand U8573 (N_8573,N_4233,N_3542);
nand U8574 (N_8574,N_930,N_628);
or U8575 (N_8575,N_851,N_4780);
nand U8576 (N_8576,N_1444,N_4442);
or U8577 (N_8577,N_1050,N_4479);
and U8578 (N_8578,N_914,N_4560);
nand U8579 (N_8579,N_3515,N_2933);
or U8580 (N_8580,N_2406,N_3031);
nand U8581 (N_8581,N_4926,N_4540);
nor U8582 (N_8582,N_3887,N_3811);
nand U8583 (N_8583,N_1392,N_1705);
and U8584 (N_8584,N_4150,N_1448);
and U8585 (N_8585,N_838,N_1616);
and U8586 (N_8586,N_502,N_4621);
nor U8587 (N_8587,N_3566,N_3298);
nand U8588 (N_8588,N_989,N_1857);
xnor U8589 (N_8589,N_4253,N_3765);
nor U8590 (N_8590,N_107,N_3647);
nor U8591 (N_8591,N_972,N_433);
and U8592 (N_8592,N_536,N_2809);
nor U8593 (N_8593,N_4065,N_328);
nor U8594 (N_8594,N_3124,N_3208);
xnor U8595 (N_8595,N_2088,N_2786);
or U8596 (N_8596,N_1067,N_3241);
or U8597 (N_8597,N_1007,N_586);
and U8598 (N_8598,N_4855,N_2949);
nor U8599 (N_8599,N_1176,N_2084);
nor U8600 (N_8600,N_2312,N_10);
nor U8601 (N_8601,N_676,N_1766);
and U8602 (N_8602,N_934,N_4386);
or U8603 (N_8603,N_2567,N_4108);
nor U8604 (N_8604,N_3744,N_1680);
or U8605 (N_8605,N_1984,N_1958);
nand U8606 (N_8606,N_2642,N_4333);
or U8607 (N_8607,N_2849,N_2148);
or U8608 (N_8608,N_1170,N_1705);
nand U8609 (N_8609,N_3290,N_4907);
nand U8610 (N_8610,N_1979,N_4522);
nor U8611 (N_8611,N_222,N_3659);
nand U8612 (N_8612,N_554,N_4630);
nor U8613 (N_8613,N_4177,N_790);
nor U8614 (N_8614,N_2943,N_311);
nor U8615 (N_8615,N_3274,N_2144);
nand U8616 (N_8616,N_3139,N_3361);
and U8617 (N_8617,N_2879,N_3213);
or U8618 (N_8618,N_4651,N_2435);
and U8619 (N_8619,N_2638,N_931);
nor U8620 (N_8620,N_1991,N_4049);
or U8621 (N_8621,N_2937,N_2029);
and U8622 (N_8622,N_3078,N_2314);
or U8623 (N_8623,N_1800,N_482);
and U8624 (N_8624,N_1731,N_2175);
nand U8625 (N_8625,N_1033,N_3669);
and U8626 (N_8626,N_1203,N_168);
and U8627 (N_8627,N_973,N_1439);
nand U8628 (N_8628,N_2632,N_1504);
nand U8629 (N_8629,N_206,N_4592);
xor U8630 (N_8630,N_4036,N_972);
or U8631 (N_8631,N_4371,N_1170);
nor U8632 (N_8632,N_3769,N_4461);
or U8633 (N_8633,N_872,N_4203);
xor U8634 (N_8634,N_1162,N_750);
nor U8635 (N_8635,N_1502,N_1483);
or U8636 (N_8636,N_3453,N_1963);
nor U8637 (N_8637,N_3687,N_71);
nor U8638 (N_8638,N_432,N_1174);
xor U8639 (N_8639,N_629,N_1988);
xnor U8640 (N_8640,N_81,N_1009);
or U8641 (N_8641,N_3081,N_4232);
nor U8642 (N_8642,N_4784,N_2203);
nand U8643 (N_8643,N_753,N_4769);
and U8644 (N_8644,N_1875,N_4622);
nand U8645 (N_8645,N_4139,N_1624);
nand U8646 (N_8646,N_1426,N_4049);
nor U8647 (N_8647,N_4761,N_574);
or U8648 (N_8648,N_3587,N_544);
nand U8649 (N_8649,N_153,N_3445);
nor U8650 (N_8650,N_1171,N_1633);
nand U8651 (N_8651,N_2741,N_954);
xor U8652 (N_8652,N_3640,N_3052);
nand U8653 (N_8653,N_2205,N_169);
nor U8654 (N_8654,N_2063,N_3127);
nor U8655 (N_8655,N_2314,N_3878);
or U8656 (N_8656,N_667,N_2064);
nor U8657 (N_8657,N_4160,N_3092);
or U8658 (N_8658,N_743,N_2343);
nor U8659 (N_8659,N_3402,N_1564);
and U8660 (N_8660,N_2249,N_3681);
and U8661 (N_8661,N_2088,N_952);
and U8662 (N_8662,N_2768,N_152);
nor U8663 (N_8663,N_4381,N_350);
nand U8664 (N_8664,N_1959,N_1630);
xor U8665 (N_8665,N_1737,N_4099);
or U8666 (N_8666,N_2404,N_1995);
and U8667 (N_8667,N_1596,N_3388);
or U8668 (N_8668,N_3317,N_3806);
or U8669 (N_8669,N_1599,N_4711);
nand U8670 (N_8670,N_2212,N_3105);
or U8671 (N_8671,N_99,N_3271);
and U8672 (N_8672,N_4460,N_1143);
nand U8673 (N_8673,N_2715,N_4302);
nand U8674 (N_8674,N_3878,N_586);
and U8675 (N_8675,N_1645,N_3834);
nor U8676 (N_8676,N_929,N_2979);
or U8677 (N_8677,N_4694,N_4148);
nor U8678 (N_8678,N_2316,N_459);
nand U8679 (N_8679,N_4149,N_2803);
or U8680 (N_8680,N_4118,N_496);
nor U8681 (N_8681,N_4908,N_168);
xor U8682 (N_8682,N_1426,N_2923);
nand U8683 (N_8683,N_830,N_2743);
or U8684 (N_8684,N_2384,N_2679);
and U8685 (N_8685,N_3453,N_3570);
or U8686 (N_8686,N_3344,N_3678);
and U8687 (N_8687,N_3378,N_3344);
and U8688 (N_8688,N_4101,N_4081);
xor U8689 (N_8689,N_3313,N_4504);
nor U8690 (N_8690,N_767,N_3983);
xnor U8691 (N_8691,N_2579,N_4715);
nor U8692 (N_8692,N_2353,N_4389);
nor U8693 (N_8693,N_3393,N_3080);
or U8694 (N_8694,N_1226,N_2749);
or U8695 (N_8695,N_2966,N_3824);
nand U8696 (N_8696,N_2829,N_2013);
nor U8697 (N_8697,N_4493,N_4999);
or U8698 (N_8698,N_234,N_3578);
nor U8699 (N_8699,N_3588,N_845);
nor U8700 (N_8700,N_2138,N_1879);
nand U8701 (N_8701,N_2669,N_4152);
xor U8702 (N_8702,N_913,N_4611);
nor U8703 (N_8703,N_814,N_2211);
or U8704 (N_8704,N_1143,N_874);
and U8705 (N_8705,N_130,N_3488);
nor U8706 (N_8706,N_489,N_2706);
nor U8707 (N_8707,N_4905,N_1277);
nor U8708 (N_8708,N_3420,N_383);
xnor U8709 (N_8709,N_2696,N_636);
and U8710 (N_8710,N_822,N_1481);
or U8711 (N_8711,N_1110,N_3398);
xor U8712 (N_8712,N_4550,N_4849);
nand U8713 (N_8713,N_1536,N_633);
nand U8714 (N_8714,N_4549,N_360);
nand U8715 (N_8715,N_2263,N_288);
nand U8716 (N_8716,N_3222,N_3727);
and U8717 (N_8717,N_3234,N_4016);
nor U8718 (N_8718,N_4261,N_3775);
xor U8719 (N_8719,N_3484,N_934);
xor U8720 (N_8720,N_2618,N_459);
xnor U8721 (N_8721,N_1571,N_4203);
nor U8722 (N_8722,N_2458,N_4913);
nand U8723 (N_8723,N_223,N_933);
xor U8724 (N_8724,N_4808,N_1870);
xor U8725 (N_8725,N_2023,N_2841);
nor U8726 (N_8726,N_829,N_1318);
nor U8727 (N_8727,N_691,N_1906);
nand U8728 (N_8728,N_2617,N_3689);
nor U8729 (N_8729,N_640,N_1111);
or U8730 (N_8730,N_2512,N_3555);
xor U8731 (N_8731,N_2292,N_1198);
or U8732 (N_8732,N_4385,N_4031);
nor U8733 (N_8733,N_4496,N_2324);
xor U8734 (N_8734,N_392,N_3067);
and U8735 (N_8735,N_1706,N_4240);
nand U8736 (N_8736,N_1501,N_561);
or U8737 (N_8737,N_2469,N_4544);
or U8738 (N_8738,N_794,N_3498);
or U8739 (N_8739,N_4396,N_3150);
and U8740 (N_8740,N_1773,N_40);
and U8741 (N_8741,N_1548,N_4914);
and U8742 (N_8742,N_2289,N_1832);
or U8743 (N_8743,N_330,N_3361);
and U8744 (N_8744,N_3250,N_2075);
or U8745 (N_8745,N_965,N_1907);
nand U8746 (N_8746,N_1857,N_2196);
and U8747 (N_8747,N_1170,N_4376);
or U8748 (N_8748,N_3259,N_1284);
nor U8749 (N_8749,N_3764,N_3048);
nor U8750 (N_8750,N_620,N_3565);
nand U8751 (N_8751,N_2060,N_4446);
xnor U8752 (N_8752,N_1126,N_4734);
or U8753 (N_8753,N_103,N_2102);
or U8754 (N_8754,N_2329,N_262);
nor U8755 (N_8755,N_2821,N_1814);
nor U8756 (N_8756,N_3293,N_3869);
nand U8757 (N_8757,N_652,N_819);
or U8758 (N_8758,N_3941,N_4131);
and U8759 (N_8759,N_4497,N_4103);
or U8760 (N_8760,N_4826,N_4624);
nor U8761 (N_8761,N_4520,N_3165);
and U8762 (N_8762,N_1510,N_1191);
and U8763 (N_8763,N_4165,N_735);
nand U8764 (N_8764,N_4734,N_2227);
xnor U8765 (N_8765,N_3276,N_4568);
nand U8766 (N_8766,N_1948,N_1309);
or U8767 (N_8767,N_3656,N_2898);
nand U8768 (N_8768,N_3946,N_2223);
nand U8769 (N_8769,N_823,N_2772);
nand U8770 (N_8770,N_962,N_2418);
or U8771 (N_8771,N_432,N_818);
nor U8772 (N_8772,N_4651,N_130);
and U8773 (N_8773,N_492,N_3632);
or U8774 (N_8774,N_3524,N_3131);
or U8775 (N_8775,N_2220,N_3332);
nand U8776 (N_8776,N_1525,N_4169);
or U8777 (N_8777,N_4141,N_56);
nor U8778 (N_8778,N_964,N_1146);
nor U8779 (N_8779,N_4677,N_498);
and U8780 (N_8780,N_1428,N_3643);
or U8781 (N_8781,N_972,N_2536);
nor U8782 (N_8782,N_2664,N_1630);
nor U8783 (N_8783,N_2249,N_4435);
or U8784 (N_8784,N_4350,N_167);
nand U8785 (N_8785,N_4645,N_4722);
and U8786 (N_8786,N_3433,N_2894);
or U8787 (N_8787,N_275,N_2974);
nand U8788 (N_8788,N_3867,N_51);
and U8789 (N_8789,N_325,N_4635);
nor U8790 (N_8790,N_3043,N_3075);
nand U8791 (N_8791,N_3243,N_1959);
and U8792 (N_8792,N_4723,N_3752);
or U8793 (N_8793,N_2,N_3764);
nor U8794 (N_8794,N_4284,N_4489);
and U8795 (N_8795,N_4622,N_3590);
or U8796 (N_8796,N_1520,N_1529);
or U8797 (N_8797,N_1229,N_1765);
nor U8798 (N_8798,N_4653,N_15);
nor U8799 (N_8799,N_3337,N_93);
or U8800 (N_8800,N_1551,N_3580);
nor U8801 (N_8801,N_647,N_2394);
and U8802 (N_8802,N_3002,N_584);
nor U8803 (N_8803,N_4647,N_4861);
nand U8804 (N_8804,N_372,N_2726);
or U8805 (N_8805,N_3904,N_922);
xnor U8806 (N_8806,N_1486,N_1769);
xnor U8807 (N_8807,N_4211,N_248);
or U8808 (N_8808,N_4015,N_1582);
xnor U8809 (N_8809,N_1707,N_1023);
and U8810 (N_8810,N_4633,N_2636);
xor U8811 (N_8811,N_371,N_638);
nor U8812 (N_8812,N_2337,N_1351);
or U8813 (N_8813,N_1390,N_2677);
and U8814 (N_8814,N_24,N_2270);
nor U8815 (N_8815,N_2433,N_233);
nor U8816 (N_8816,N_2848,N_3284);
and U8817 (N_8817,N_3626,N_3062);
and U8818 (N_8818,N_146,N_2414);
and U8819 (N_8819,N_2786,N_1067);
nor U8820 (N_8820,N_4906,N_1277);
or U8821 (N_8821,N_2764,N_4848);
nand U8822 (N_8822,N_1470,N_487);
nand U8823 (N_8823,N_2152,N_3877);
and U8824 (N_8824,N_3597,N_3968);
or U8825 (N_8825,N_4582,N_4618);
or U8826 (N_8826,N_4170,N_4071);
nand U8827 (N_8827,N_1983,N_3990);
nand U8828 (N_8828,N_1110,N_277);
and U8829 (N_8829,N_1359,N_3165);
and U8830 (N_8830,N_697,N_2062);
nor U8831 (N_8831,N_4905,N_4303);
nand U8832 (N_8832,N_3483,N_2532);
nor U8833 (N_8833,N_2225,N_2144);
nand U8834 (N_8834,N_4639,N_960);
xor U8835 (N_8835,N_4401,N_4270);
nand U8836 (N_8836,N_2756,N_4631);
and U8837 (N_8837,N_3485,N_3477);
nor U8838 (N_8838,N_1637,N_2006);
or U8839 (N_8839,N_1133,N_4297);
and U8840 (N_8840,N_1084,N_4403);
and U8841 (N_8841,N_3659,N_4022);
and U8842 (N_8842,N_2441,N_4132);
nand U8843 (N_8843,N_3906,N_1212);
nand U8844 (N_8844,N_2586,N_2871);
or U8845 (N_8845,N_3656,N_2011);
or U8846 (N_8846,N_142,N_1392);
nor U8847 (N_8847,N_3815,N_3910);
and U8848 (N_8848,N_2825,N_4432);
nand U8849 (N_8849,N_155,N_1323);
and U8850 (N_8850,N_2832,N_1191);
nor U8851 (N_8851,N_3797,N_3867);
or U8852 (N_8852,N_2001,N_2089);
nor U8853 (N_8853,N_3323,N_4842);
nor U8854 (N_8854,N_195,N_4393);
nand U8855 (N_8855,N_2992,N_806);
nand U8856 (N_8856,N_4342,N_3657);
and U8857 (N_8857,N_4759,N_770);
nor U8858 (N_8858,N_2783,N_3161);
or U8859 (N_8859,N_941,N_2906);
xor U8860 (N_8860,N_4255,N_3319);
nand U8861 (N_8861,N_2586,N_604);
nor U8862 (N_8862,N_2933,N_3201);
and U8863 (N_8863,N_698,N_3633);
xor U8864 (N_8864,N_204,N_764);
nor U8865 (N_8865,N_3641,N_1244);
nand U8866 (N_8866,N_4804,N_4444);
nand U8867 (N_8867,N_3964,N_910);
xor U8868 (N_8868,N_1868,N_4575);
xnor U8869 (N_8869,N_2918,N_4197);
and U8870 (N_8870,N_1292,N_2281);
nand U8871 (N_8871,N_2464,N_3566);
nand U8872 (N_8872,N_974,N_4891);
and U8873 (N_8873,N_4478,N_3022);
and U8874 (N_8874,N_2146,N_3163);
nand U8875 (N_8875,N_4294,N_991);
and U8876 (N_8876,N_1745,N_4233);
or U8877 (N_8877,N_1173,N_4675);
and U8878 (N_8878,N_1691,N_1454);
nand U8879 (N_8879,N_1272,N_1261);
or U8880 (N_8880,N_3340,N_2116);
xnor U8881 (N_8881,N_764,N_662);
or U8882 (N_8882,N_791,N_4964);
and U8883 (N_8883,N_818,N_3619);
and U8884 (N_8884,N_1539,N_1827);
or U8885 (N_8885,N_2595,N_4734);
and U8886 (N_8886,N_4073,N_1388);
nand U8887 (N_8887,N_4488,N_2338);
xor U8888 (N_8888,N_3543,N_3392);
nor U8889 (N_8889,N_4907,N_1369);
or U8890 (N_8890,N_2866,N_4968);
nand U8891 (N_8891,N_4719,N_2002);
nand U8892 (N_8892,N_2551,N_1288);
and U8893 (N_8893,N_647,N_293);
nand U8894 (N_8894,N_2124,N_1936);
and U8895 (N_8895,N_778,N_3689);
xnor U8896 (N_8896,N_3738,N_2742);
and U8897 (N_8897,N_267,N_1298);
and U8898 (N_8898,N_4496,N_2856);
or U8899 (N_8899,N_709,N_570);
nor U8900 (N_8900,N_311,N_86);
or U8901 (N_8901,N_2125,N_1169);
nor U8902 (N_8902,N_3735,N_3473);
nand U8903 (N_8903,N_1776,N_759);
or U8904 (N_8904,N_3983,N_1835);
nor U8905 (N_8905,N_2016,N_1521);
nand U8906 (N_8906,N_1484,N_3903);
or U8907 (N_8907,N_3013,N_3685);
and U8908 (N_8908,N_1324,N_2195);
nor U8909 (N_8909,N_3129,N_965);
xnor U8910 (N_8910,N_3956,N_1438);
nand U8911 (N_8911,N_2898,N_1366);
nor U8912 (N_8912,N_1082,N_401);
nor U8913 (N_8913,N_1287,N_2927);
or U8914 (N_8914,N_215,N_3371);
and U8915 (N_8915,N_1392,N_848);
or U8916 (N_8916,N_706,N_3458);
and U8917 (N_8917,N_4375,N_1113);
nand U8918 (N_8918,N_2106,N_1203);
and U8919 (N_8919,N_2264,N_4546);
or U8920 (N_8920,N_4865,N_1105);
or U8921 (N_8921,N_2213,N_658);
nand U8922 (N_8922,N_3714,N_570);
or U8923 (N_8923,N_1731,N_3675);
and U8924 (N_8924,N_654,N_3991);
or U8925 (N_8925,N_1052,N_47);
xor U8926 (N_8926,N_4700,N_3401);
xnor U8927 (N_8927,N_866,N_1566);
and U8928 (N_8928,N_241,N_3772);
nor U8929 (N_8929,N_4528,N_3498);
and U8930 (N_8930,N_2576,N_4142);
xor U8931 (N_8931,N_3658,N_495);
nand U8932 (N_8932,N_3763,N_592);
or U8933 (N_8933,N_1368,N_2120);
and U8934 (N_8934,N_1177,N_3738);
or U8935 (N_8935,N_420,N_4836);
and U8936 (N_8936,N_2391,N_2320);
and U8937 (N_8937,N_763,N_324);
and U8938 (N_8938,N_2014,N_1164);
nand U8939 (N_8939,N_189,N_730);
nand U8940 (N_8940,N_2037,N_4881);
or U8941 (N_8941,N_3608,N_1712);
or U8942 (N_8942,N_3483,N_1438);
and U8943 (N_8943,N_1421,N_3694);
xor U8944 (N_8944,N_458,N_3696);
xor U8945 (N_8945,N_2096,N_1415);
or U8946 (N_8946,N_4545,N_2718);
nand U8947 (N_8947,N_2854,N_4849);
and U8948 (N_8948,N_4378,N_4214);
nand U8949 (N_8949,N_3749,N_1362);
nand U8950 (N_8950,N_1807,N_4207);
and U8951 (N_8951,N_1177,N_3827);
nor U8952 (N_8952,N_3142,N_3357);
or U8953 (N_8953,N_629,N_1792);
nand U8954 (N_8954,N_1183,N_4432);
and U8955 (N_8955,N_3512,N_3467);
and U8956 (N_8956,N_876,N_4501);
xnor U8957 (N_8957,N_4490,N_2916);
or U8958 (N_8958,N_3067,N_2924);
and U8959 (N_8959,N_3496,N_4624);
or U8960 (N_8960,N_795,N_3906);
nand U8961 (N_8961,N_3103,N_2611);
or U8962 (N_8962,N_4717,N_1406);
nor U8963 (N_8963,N_2466,N_977);
nor U8964 (N_8964,N_4854,N_3063);
nand U8965 (N_8965,N_994,N_4650);
xor U8966 (N_8966,N_2592,N_3417);
or U8967 (N_8967,N_3759,N_3055);
and U8968 (N_8968,N_4559,N_1065);
nand U8969 (N_8969,N_3887,N_1736);
and U8970 (N_8970,N_537,N_1800);
or U8971 (N_8971,N_2939,N_1465);
or U8972 (N_8972,N_676,N_2045);
or U8973 (N_8973,N_4140,N_2209);
nand U8974 (N_8974,N_4815,N_1927);
nand U8975 (N_8975,N_3971,N_2389);
nor U8976 (N_8976,N_3334,N_4785);
nor U8977 (N_8977,N_3978,N_2623);
and U8978 (N_8978,N_1416,N_4887);
or U8979 (N_8979,N_3409,N_656);
nand U8980 (N_8980,N_1794,N_1818);
or U8981 (N_8981,N_4796,N_3910);
and U8982 (N_8982,N_4803,N_972);
and U8983 (N_8983,N_4164,N_3441);
and U8984 (N_8984,N_4472,N_1003);
nand U8985 (N_8985,N_1229,N_642);
or U8986 (N_8986,N_1757,N_1848);
nand U8987 (N_8987,N_3318,N_4045);
and U8988 (N_8988,N_1128,N_924);
nor U8989 (N_8989,N_2345,N_3592);
nor U8990 (N_8990,N_2381,N_1579);
or U8991 (N_8991,N_3760,N_1268);
xnor U8992 (N_8992,N_391,N_2786);
and U8993 (N_8993,N_685,N_2228);
nand U8994 (N_8994,N_1685,N_3229);
nand U8995 (N_8995,N_1084,N_137);
nand U8996 (N_8996,N_1661,N_1537);
xor U8997 (N_8997,N_1494,N_999);
and U8998 (N_8998,N_3003,N_4632);
nand U8999 (N_8999,N_1938,N_4311);
nor U9000 (N_9000,N_4405,N_2619);
or U9001 (N_9001,N_312,N_3952);
nand U9002 (N_9002,N_2024,N_1377);
nand U9003 (N_9003,N_3625,N_572);
or U9004 (N_9004,N_1234,N_4612);
nor U9005 (N_9005,N_1949,N_923);
and U9006 (N_9006,N_1608,N_2939);
xor U9007 (N_9007,N_2365,N_2548);
and U9008 (N_9008,N_3379,N_2625);
nand U9009 (N_9009,N_4390,N_3824);
and U9010 (N_9010,N_1577,N_415);
nor U9011 (N_9011,N_2974,N_1468);
and U9012 (N_9012,N_4448,N_1141);
and U9013 (N_9013,N_2551,N_2326);
xor U9014 (N_9014,N_2926,N_2905);
nand U9015 (N_9015,N_1517,N_1883);
nor U9016 (N_9016,N_679,N_1013);
nand U9017 (N_9017,N_3948,N_3055);
or U9018 (N_9018,N_3203,N_2840);
and U9019 (N_9019,N_879,N_1198);
xor U9020 (N_9020,N_608,N_1176);
or U9021 (N_9021,N_2043,N_1935);
or U9022 (N_9022,N_49,N_1285);
nor U9023 (N_9023,N_3167,N_4822);
or U9024 (N_9024,N_78,N_4519);
nand U9025 (N_9025,N_4714,N_3254);
and U9026 (N_9026,N_2820,N_702);
nor U9027 (N_9027,N_1717,N_497);
and U9028 (N_9028,N_4442,N_729);
and U9029 (N_9029,N_3957,N_1445);
xnor U9030 (N_9030,N_264,N_1884);
or U9031 (N_9031,N_1281,N_2740);
and U9032 (N_9032,N_32,N_4159);
xor U9033 (N_9033,N_1470,N_4334);
nor U9034 (N_9034,N_3148,N_106);
and U9035 (N_9035,N_4509,N_3247);
nand U9036 (N_9036,N_1188,N_2188);
or U9037 (N_9037,N_1816,N_1772);
and U9038 (N_9038,N_4499,N_1521);
nand U9039 (N_9039,N_1663,N_145);
and U9040 (N_9040,N_4891,N_1946);
and U9041 (N_9041,N_1340,N_3973);
or U9042 (N_9042,N_1448,N_3560);
and U9043 (N_9043,N_1036,N_4013);
nand U9044 (N_9044,N_1846,N_1884);
nand U9045 (N_9045,N_1233,N_2139);
and U9046 (N_9046,N_3702,N_308);
xnor U9047 (N_9047,N_2763,N_1814);
nand U9048 (N_9048,N_4147,N_99);
or U9049 (N_9049,N_1041,N_3414);
and U9050 (N_9050,N_546,N_3164);
nor U9051 (N_9051,N_3964,N_3796);
nand U9052 (N_9052,N_4762,N_1437);
nor U9053 (N_9053,N_3188,N_713);
nor U9054 (N_9054,N_2910,N_4134);
or U9055 (N_9055,N_2943,N_4068);
nor U9056 (N_9056,N_3729,N_1798);
nor U9057 (N_9057,N_718,N_2986);
xor U9058 (N_9058,N_2359,N_3032);
xnor U9059 (N_9059,N_1782,N_4882);
or U9060 (N_9060,N_2643,N_297);
and U9061 (N_9061,N_3736,N_410);
nand U9062 (N_9062,N_3922,N_2998);
nand U9063 (N_9063,N_1155,N_4064);
or U9064 (N_9064,N_169,N_3662);
xor U9065 (N_9065,N_2513,N_894);
nand U9066 (N_9066,N_2856,N_196);
nor U9067 (N_9067,N_3704,N_2330);
and U9068 (N_9068,N_3534,N_2059);
or U9069 (N_9069,N_384,N_3983);
nand U9070 (N_9070,N_3733,N_2846);
or U9071 (N_9071,N_1059,N_3158);
nand U9072 (N_9072,N_3924,N_1224);
and U9073 (N_9073,N_2674,N_4517);
and U9074 (N_9074,N_4228,N_1012);
or U9075 (N_9075,N_3143,N_3630);
and U9076 (N_9076,N_2760,N_394);
and U9077 (N_9077,N_1547,N_1205);
nand U9078 (N_9078,N_2574,N_3374);
nor U9079 (N_9079,N_4862,N_2521);
xor U9080 (N_9080,N_4980,N_4412);
nand U9081 (N_9081,N_3737,N_2865);
and U9082 (N_9082,N_4750,N_3487);
xnor U9083 (N_9083,N_4631,N_4581);
nor U9084 (N_9084,N_2007,N_3820);
nor U9085 (N_9085,N_0,N_825);
or U9086 (N_9086,N_2434,N_4951);
nor U9087 (N_9087,N_2339,N_3840);
nand U9088 (N_9088,N_2413,N_2704);
nand U9089 (N_9089,N_3878,N_1773);
and U9090 (N_9090,N_2005,N_256);
nor U9091 (N_9091,N_3548,N_3206);
or U9092 (N_9092,N_3116,N_3114);
xnor U9093 (N_9093,N_4422,N_2012);
nor U9094 (N_9094,N_925,N_302);
nor U9095 (N_9095,N_4565,N_1078);
nand U9096 (N_9096,N_1842,N_715);
nand U9097 (N_9097,N_1476,N_362);
nor U9098 (N_9098,N_1119,N_2558);
and U9099 (N_9099,N_4089,N_4926);
nor U9100 (N_9100,N_68,N_2705);
nor U9101 (N_9101,N_1165,N_2650);
or U9102 (N_9102,N_709,N_3888);
or U9103 (N_9103,N_4269,N_3966);
nor U9104 (N_9104,N_1503,N_1995);
and U9105 (N_9105,N_830,N_4640);
or U9106 (N_9106,N_2479,N_4547);
and U9107 (N_9107,N_766,N_2392);
nand U9108 (N_9108,N_3163,N_3850);
or U9109 (N_9109,N_450,N_3494);
nor U9110 (N_9110,N_1864,N_346);
nor U9111 (N_9111,N_2627,N_3645);
nor U9112 (N_9112,N_3161,N_3189);
or U9113 (N_9113,N_2509,N_3614);
and U9114 (N_9114,N_2182,N_3539);
xnor U9115 (N_9115,N_1136,N_1505);
and U9116 (N_9116,N_1838,N_1435);
nand U9117 (N_9117,N_1658,N_3779);
or U9118 (N_9118,N_4147,N_2258);
nand U9119 (N_9119,N_3095,N_159);
nand U9120 (N_9120,N_1621,N_4306);
nor U9121 (N_9121,N_3757,N_3792);
and U9122 (N_9122,N_3344,N_2349);
and U9123 (N_9123,N_1900,N_271);
or U9124 (N_9124,N_344,N_2190);
nand U9125 (N_9125,N_3285,N_3894);
or U9126 (N_9126,N_2148,N_3376);
or U9127 (N_9127,N_1573,N_3446);
or U9128 (N_9128,N_3851,N_2100);
or U9129 (N_9129,N_3683,N_910);
or U9130 (N_9130,N_3721,N_3677);
and U9131 (N_9131,N_1879,N_4378);
nor U9132 (N_9132,N_640,N_2803);
and U9133 (N_9133,N_933,N_3625);
nor U9134 (N_9134,N_2029,N_3860);
or U9135 (N_9135,N_3982,N_1966);
nor U9136 (N_9136,N_2026,N_1516);
nand U9137 (N_9137,N_4871,N_2527);
nor U9138 (N_9138,N_294,N_4673);
or U9139 (N_9139,N_2463,N_1502);
and U9140 (N_9140,N_4232,N_2771);
nor U9141 (N_9141,N_3934,N_531);
nor U9142 (N_9142,N_652,N_843);
nand U9143 (N_9143,N_4169,N_2171);
and U9144 (N_9144,N_1889,N_647);
nand U9145 (N_9145,N_4508,N_2199);
nand U9146 (N_9146,N_1540,N_4313);
and U9147 (N_9147,N_3133,N_1204);
xnor U9148 (N_9148,N_2674,N_2749);
and U9149 (N_9149,N_4108,N_2886);
nor U9150 (N_9150,N_4108,N_1245);
and U9151 (N_9151,N_913,N_734);
and U9152 (N_9152,N_4875,N_4217);
and U9153 (N_9153,N_4045,N_898);
and U9154 (N_9154,N_3400,N_1754);
nand U9155 (N_9155,N_1293,N_4987);
nor U9156 (N_9156,N_4676,N_2062);
or U9157 (N_9157,N_769,N_2762);
nor U9158 (N_9158,N_2258,N_2393);
nor U9159 (N_9159,N_2892,N_1368);
and U9160 (N_9160,N_4831,N_3019);
nor U9161 (N_9161,N_479,N_3650);
nor U9162 (N_9162,N_405,N_1510);
nand U9163 (N_9163,N_337,N_2444);
and U9164 (N_9164,N_3625,N_4115);
xor U9165 (N_9165,N_498,N_786);
and U9166 (N_9166,N_314,N_116);
nor U9167 (N_9167,N_1034,N_1385);
xnor U9168 (N_9168,N_3438,N_3366);
nand U9169 (N_9169,N_1767,N_2929);
nor U9170 (N_9170,N_956,N_1790);
xnor U9171 (N_9171,N_4534,N_3492);
nor U9172 (N_9172,N_4667,N_458);
nor U9173 (N_9173,N_3107,N_753);
or U9174 (N_9174,N_1073,N_245);
or U9175 (N_9175,N_910,N_3615);
or U9176 (N_9176,N_3043,N_4428);
xor U9177 (N_9177,N_778,N_4909);
nand U9178 (N_9178,N_3206,N_4062);
nor U9179 (N_9179,N_2777,N_3740);
nand U9180 (N_9180,N_1055,N_2933);
nand U9181 (N_9181,N_2498,N_2559);
and U9182 (N_9182,N_3376,N_4748);
xor U9183 (N_9183,N_1034,N_1040);
nor U9184 (N_9184,N_3380,N_218);
or U9185 (N_9185,N_908,N_2956);
nand U9186 (N_9186,N_4084,N_585);
nor U9187 (N_9187,N_535,N_3245);
and U9188 (N_9188,N_4713,N_576);
nor U9189 (N_9189,N_1602,N_1985);
nand U9190 (N_9190,N_2412,N_3348);
and U9191 (N_9191,N_2479,N_2014);
nand U9192 (N_9192,N_3166,N_3132);
and U9193 (N_9193,N_967,N_3718);
and U9194 (N_9194,N_1078,N_1489);
nand U9195 (N_9195,N_2379,N_3603);
nand U9196 (N_9196,N_3615,N_519);
or U9197 (N_9197,N_3675,N_1653);
nor U9198 (N_9198,N_2565,N_1657);
nor U9199 (N_9199,N_3077,N_4239);
or U9200 (N_9200,N_763,N_3842);
nand U9201 (N_9201,N_3022,N_2912);
or U9202 (N_9202,N_234,N_1133);
or U9203 (N_9203,N_2785,N_3832);
nor U9204 (N_9204,N_470,N_2978);
nor U9205 (N_9205,N_4134,N_2454);
xor U9206 (N_9206,N_4348,N_2599);
and U9207 (N_9207,N_1649,N_303);
nor U9208 (N_9208,N_3870,N_1688);
nand U9209 (N_9209,N_1012,N_3842);
nor U9210 (N_9210,N_4926,N_4851);
and U9211 (N_9211,N_2904,N_1902);
nand U9212 (N_9212,N_4544,N_1435);
or U9213 (N_9213,N_3858,N_3714);
or U9214 (N_9214,N_4719,N_4331);
nand U9215 (N_9215,N_2723,N_3613);
nand U9216 (N_9216,N_939,N_1121);
xnor U9217 (N_9217,N_4345,N_3294);
or U9218 (N_9218,N_3550,N_13);
xnor U9219 (N_9219,N_4553,N_2576);
nor U9220 (N_9220,N_3941,N_1171);
xnor U9221 (N_9221,N_930,N_2750);
nor U9222 (N_9222,N_99,N_587);
and U9223 (N_9223,N_2193,N_3207);
or U9224 (N_9224,N_3770,N_2121);
nand U9225 (N_9225,N_3002,N_954);
nor U9226 (N_9226,N_4336,N_3795);
nand U9227 (N_9227,N_2147,N_1450);
nor U9228 (N_9228,N_578,N_4988);
nor U9229 (N_9229,N_4841,N_4573);
nor U9230 (N_9230,N_3244,N_2231);
xor U9231 (N_9231,N_4709,N_4565);
or U9232 (N_9232,N_1109,N_3485);
and U9233 (N_9233,N_566,N_859);
and U9234 (N_9234,N_21,N_1404);
or U9235 (N_9235,N_4307,N_3328);
or U9236 (N_9236,N_848,N_249);
nand U9237 (N_9237,N_173,N_3483);
or U9238 (N_9238,N_822,N_2191);
and U9239 (N_9239,N_942,N_740);
xor U9240 (N_9240,N_3788,N_4853);
and U9241 (N_9241,N_4704,N_3141);
xnor U9242 (N_9242,N_4821,N_399);
nand U9243 (N_9243,N_1666,N_3011);
or U9244 (N_9244,N_1318,N_3239);
nand U9245 (N_9245,N_883,N_1405);
xor U9246 (N_9246,N_1147,N_2971);
nor U9247 (N_9247,N_3057,N_2873);
or U9248 (N_9248,N_4954,N_4151);
and U9249 (N_9249,N_70,N_4816);
nand U9250 (N_9250,N_3790,N_1753);
nand U9251 (N_9251,N_4840,N_3593);
nand U9252 (N_9252,N_2942,N_992);
and U9253 (N_9253,N_1211,N_3041);
or U9254 (N_9254,N_3059,N_1447);
nor U9255 (N_9255,N_121,N_3150);
or U9256 (N_9256,N_3050,N_3999);
nand U9257 (N_9257,N_1702,N_3066);
nand U9258 (N_9258,N_2454,N_3551);
or U9259 (N_9259,N_4744,N_920);
and U9260 (N_9260,N_3877,N_41);
nor U9261 (N_9261,N_4815,N_2822);
and U9262 (N_9262,N_2882,N_2164);
nor U9263 (N_9263,N_4660,N_3002);
nand U9264 (N_9264,N_4330,N_1392);
or U9265 (N_9265,N_1428,N_1010);
nand U9266 (N_9266,N_3277,N_3496);
nor U9267 (N_9267,N_267,N_3738);
nor U9268 (N_9268,N_658,N_3652);
nor U9269 (N_9269,N_2046,N_4770);
nand U9270 (N_9270,N_4032,N_1932);
or U9271 (N_9271,N_4293,N_2019);
nor U9272 (N_9272,N_748,N_806);
and U9273 (N_9273,N_4490,N_1443);
or U9274 (N_9274,N_4596,N_4321);
nor U9275 (N_9275,N_848,N_3724);
nand U9276 (N_9276,N_3432,N_583);
or U9277 (N_9277,N_3538,N_402);
nor U9278 (N_9278,N_4062,N_3126);
or U9279 (N_9279,N_1564,N_1146);
or U9280 (N_9280,N_4848,N_1501);
nand U9281 (N_9281,N_4034,N_2355);
nor U9282 (N_9282,N_3429,N_3387);
nor U9283 (N_9283,N_4557,N_4834);
or U9284 (N_9284,N_1302,N_2286);
or U9285 (N_9285,N_3710,N_4990);
and U9286 (N_9286,N_4473,N_64);
nor U9287 (N_9287,N_1277,N_1820);
nand U9288 (N_9288,N_1219,N_2088);
nor U9289 (N_9289,N_3962,N_732);
nand U9290 (N_9290,N_781,N_2451);
or U9291 (N_9291,N_3057,N_3526);
or U9292 (N_9292,N_243,N_3216);
nand U9293 (N_9293,N_3241,N_4683);
nand U9294 (N_9294,N_2562,N_2602);
nand U9295 (N_9295,N_602,N_3121);
and U9296 (N_9296,N_2877,N_2868);
nor U9297 (N_9297,N_3647,N_4187);
nor U9298 (N_9298,N_4350,N_3818);
and U9299 (N_9299,N_3251,N_2926);
and U9300 (N_9300,N_3507,N_2697);
or U9301 (N_9301,N_784,N_4266);
or U9302 (N_9302,N_3094,N_1941);
or U9303 (N_9303,N_3480,N_4284);
nand U9304 (N_9304,N_4278,N_3081);
xnor U9305 (N_9305,N_4419,N_1716);
or U9306 (N_9306,N_3080,N_1903);
nand U9307 (N_9307,N_362,N_3192);
and U9308 (N_9308,N_533,N_3267);
or U9309 (N_9309,N_4305,N_1851);
nand U9310 (N_9310,N_3284,N_3662);
or U9311 (N_9311,N_4834,N_2644);
nand U9312 (N_9312,N_4706,N_2062);
nor U9313 (N_9313,N_1729,N_616);
and U9314 (N_9314,N_2001,N_2016);
xnor U9315 (N_9315,N_2929,N_4237);
or U9316 (N_9316,N_1972,N_4378);
nand U9317 (N_9317,N_868,N_2195);
or U9318 (N_9318,N_4756,N_2072);
or U9319 (N_9319,N_3375,N_863);
xnor U9320 (N_9320,N_3442,N_1483);
nor U9321 (N_9321,N_2388,N_2370);
and U9322 (N_9322,N_4241,N_453);
nand U9323 (N_9323,N_2668,N_3616);
or U9324 (N_9324,N_147,N_2196);
or U9325 (N_9325,N_2231,N_3328);
nor U9326 (N_9326,N_2124,N_527);
xnor U9327 (N_9327,N_575,N_763);
nand U9328 (N_9328,N_1183,N_3368);
and U9329 (N_9329,N_4853,N_4062);
or U9330 (N_9330,N_1681,N_1153);
or U9331 (N_9331,N_4682,N_1127);
nor U9332 (N_9332,N_4809,N_1874);
and U9333 (N_9333,N_3573,N_436);
or U9334 (N_9334,N_257,N_1110);
or U9335 (N_9335,N_4055,N_4292);
nor U9336 (N_9336,N_3510,N_4583);
nor U9337 (N_9337,N_3117,N_3664);
and U9338 (N_9338,N_3539,N_1883);
and U9339 (N_9339,N_3341,N_2544);
or U9340 (N_9340,N_1052,N_4334);
nand U9341 (N_9341,N_3158,N_2768);
and U9342 (N_9342,N_708,N_1780);
and U9343 (N_9343,N_1337,N_2328);
xor U9344 (N_9344,N_2969,N_726);
nor U9345 (N_9345,N_1459,N_2215);
nor U9346 (N_9346,N_3464,N_4454);
and U9347 (N_9347,N_15,N_312);
and U9348 (N_9348,N_3049,N_2471);
nand U9349 (N_9349,N_1315,N_4447);
nor U9350 (N_9350,N_3808,N_1998);
and U9351 (N_9351,N_3576,N_1604);
nor U9352 (N_9352,N_1425,N_1490);
and U9353 (N_9353,N_2867,N_3706);
nor U9354 (N_9354,N_1896,N_2203);
nor U9355 (N_9355,N_1721,N_1767);
and U9356 (N_9356,N_3799,N_3006);
and U9357 (N_9357,N_947,N_4276);
nand U9358 (N_9358,N_3020,N_931);
nor U9359 (N_9359,N_2939,N_4707);
xnor U9360 (N_9360,N_3522,N_3706);
nor U9361 (N_9361,N_2192,N_721);
nand U9362 (N_9362,N_2425,N_832);
nand U9363 (N_9363,N_4952,N_2431);
nand U9364 (N_9364,N_1777,N_122);
and U9365 (N_9365,N_1151,N_2161);
xor U9366 (N_9366,N_2312,N_1818);
and U9367 (N_9367,N_4438,N_2287);
and U9368 (N_9368,N_4462,N_98);
nor U9369 (N_9369,N_3824,N_3867);
and U9370 (N_9370,N_3774,N_2901);
or U9371 (N_9371,N_4071,N_4210);
xnor U9372 (N_9372,N_4457,N_2131);
nand U9373 (N_9373,N_2882,N_1934);
nor U9374 (N_9374,N_3208,N_260);
nor U9375 (N_9375,N_4936,N_3994);
nor U9376 (N_9376,N_4772,N_565);
or U9377 (N_9377,N_2714,N_2728);
xor U9378 (N_9378,N_3462,N_187);
or U9379 (N_9379,N_4470,N_2786);
nor U9380 (N_9380,N_3109,N_1483);
nand U9381 (N_9381,N_183,N_4992);
nor U9382 (N_9382,N_4018,N_1624);
nand U9383 (N_9383,N_3050,N_3930);
nor U9384 (N_9384,N_3431,N_1320);
or U9385 (N_9385,N_2940,N_2008);
nand U9386 (N_9386,N_3707,N_3918);
nor U9387 (N_9387,N_4184,N_829);
nand U9388 (N_9388,N_480,N_3242);
and U9389 (N_9389,N_4842,N_4102);
nand U9390 (N_9390,N_219,N_770);
nand U9391 (N_9391,N_232,N_574);
nor U9392 (N_9392,N_2949,N_282);
nand U9393 (N_9393,N_2858,N_460);
and U9394 (N_9394,N_1864,N_3751);
or U9395 (N_9395,N_2810,N_4103);
or U9396 (N_9396,N_4629,N_1350);
nor U9397 (N_9397,N_4129,N_4501);
nand U9398 (N_9398,N_628,N_4922);
and U9399 (N_9399,N_2047,N_3495);
nand U9400 (N_9400,N_3213,N_1279);
or U9401 (N_9401,N_59,N_2664);
nand U9402 (N_9402,N_2240,N_3852);
xnor U9403 (N_9403,N_3461,N_4105);
or U9404 (N_9404,N_2309,N_2484);
nor U9405 (N_9405,N_256,N_4002);
and U9406 (N_9406,N_2154,N_3818);
and U9407 (N_9407,N_1372,N_2460);
nand U9408 (N_9408,N_2426,N_2605);
nand U9409 (N_9409,N_4845,N_1036);
and U9410 (N_9410,N_4788,N_1739);
xnor U9411 (N_9411,N_1603,N_4955);
nand U9412 (N_9412,N_2209,N_4446);
and U9413 (N_9413,N_3672,N_4485);
nand U9414 (N_9414,N_4959,N_4580);
or U9415 (N_9415,N_3523,N_3502);
and U9416 (N_9416,N_72,N_4931);
and U9417 (N_9417,N_3256,N_1455);
xnor U9418 (N_9418,N_4300,N_3834);
nor U9419 (N_9419,N_2078,N_1173);
nor U9420 (N_9420,N_1406,N_3662);
nor U9421 (N_9421,N_1838,N_963);
nand U9422 (N_9422,N_3934,N_4527);
nand U9423 (N_9423,N_4000,N_2858);
nor U9424 (N_9424,N_836,N_3477);
nand U9425 (N_9425,N_4764,N_3436);
nand U9426 (N_9426,N_3740,N_756);
nand U9427 (N_9427,N_3298,N_1628);
or U9428 (N_9428,N_2732,N_4835);
nand U9429 (N_9429,N_846,N_4298);
nor U9430 (N_9430,N_1941,N_322);
nor U9431 (N_9431,N_1896,N_3147);
xor U9432 (N_9432,N_1053,N_507);
or U9433 (N_9433,N_2651,N_3542);
or U9434 (N_9434,N_1393,N_2517);
and U9435 (N_9435,N_625,N_618);
nand U9436 (N_9436,N_2844,N_3405);
and U9437 (N_9437,N_2378,N_676);
or U9438 (N_9438,N_523,N_3758);
or U9439 (N_9439,N_3671,N_2662);
nor U9440 (N_9440,N_1735,N_2417);
and U9441 (N_9441,N_3918,N_1231);
and U9442 (N_9442,N_1983,N_1816);
and U9443 (N_9443,N_4857,N_132);
nor U9444 (N_9444,N_2806,N_3991);
or U9445 (N_9445,N_2136,N_4391);
and U9446 (N_9446,N_2285,N_246);
and U9447 (N_9447,N_309,N_2106);
or U9448 (N_9448,N_900,N_3743);
nor U9449 (N_9449,N_4760,N_799);
nand U9450 (N_9450,N_252,N_4954);
nand U9451 (N_9451,N_2386,N_2580);
nor U9452 (N_9452,N_4750,N_798);
nand U9453 (N_9453,N_2980,N_2816);
nand U9454 (N_9454,N_36,N_3990);
or U9455 (N_9455,N_4272,N_1799);
nor U9456 (N_9456,N_492,N_757);
nand U9457 (N_9457,N_3880,N_2528);
and U9458 (N_9458,N_3451,N_820);
nor U9459 (N_9459,N_4412,N_4451);
or U9460 (N_9460,N_3299,N_549);
or U9461 (N_9461,N_3026,N_3650);
nor U9462 (N_9462,N_1694,N_3715);
nand U9463 (N_9463,N_524,N_1314);
nor U9464 (N_9464,N_579,N_2316);
nand U9465 (N_9465,N_734,N_2673);
or U9466 (N_9466,N_2886,N_373);
nor U9467 (N_9467,N_4311,N_3118);
and U9468 (N_9468,N_490,N_1143);
or U9469 (N_9469,N_431,N_188);
nor U9470 (N_9470,N_1658,N_2443);
nand U9471 (N_9471,N_3061,N_3324);
nand U9472 (N_9472,N_91,N_906);
and U9473 (N_9473,N_4961,N_3018);
xnor U9474 (N_9474,N_3231,N_637);
xor U9475 (N_9475,N_1764,N_129);
nand U9476 (N_9476,N_567,N_2088);
and U9477 (N_9477,N_1297,N_370);
xnor U9478 (N_9478,N_684,N_2260);
nor U9479 (N_9479,N_1074,N_3384);
or U9480 (N_9480,N_411,N_4770);
nor U9481 (N_9481,N_4459,N_1585);
or U9482 (N_9482,N_4810,N_3375);
nand U9483 (N_9483,N_176,N_500);
or U9484 (N_9484,N_637,N_2379);
nand U9485 (N_9485,N_4418,N_3612);
or U9486 (N_9486,N_2698,N_39);
or U9487 (N_9487,N_1848,N_3125);
nand U9488 (N_9488,N_1770,N_4586);
nor U9489 (N_9489,N_4855,N_2952);
and U9490 (N_9490,N_294,N_414);
and U9491 (N_9491,N_1230,N_208);
and U9492 (N_9492,N_3223,N_826);
and U9493 (N_9493,N_2872,N_176);
or U9494 (N_9494,N_1152,N_4545);
nor U9495 (N_9495,N_1189,N_3404);
and U9496 (N_9496,N_2153,N_2946);
or U9497 (N_9497,N_3274,N_3731);
nor U9498 (N_9498,N_669,N_2528);
nand U9499 (N_9499,N_3984,N_3207);
nor U9500 (N_9500,N_3682,N_1098);
and U9501 (N_9501,N_2016,N_2840);
or U9502 (N_9502,N_73,N_2006);
xor U9503 (N_9503,N_111,N_1500);
nand U9504 (N_9504,N_15,N_3358);
or U9505 (N_9505,N_76,N_601);
or U9506 (N_9506,N_2484,N_326);
nor U9507 (N_9507,N_3058,N_462);
nor U9508 (N_9508,N_3320,N_4930);
nand U9509 (N_9509,N_4058,N_4370);
nor U9510 (N_9510,N_1864,N_1254);
or U9511 (N_9511,N_184,N_653);
nor U9512 (N_9512,N_4856,N_1955);
nand U9513 (N_9513,N_2822,N_3104);
nor U9514 (N_9514,N_3136,N_8);
nand U9515 (N_9515,N_3408,N_2468);
xnor U9516 (N_9516,N_1910,N_539);
nor U9517 (N_9517,N_4352,N_3449);
nor U9518 (N_9518,N_2756,N_2749);
and U9519 (N_9519,N_1411,N_518);
nor U9520 (N_9520,N_4615,N_1332);
xor U9521 (N_9521,N_4972,N_1005);
nor U9522 (N_9522,N_3310,N_1539);
nor U9523 (N_9523,N_4012,N_1836);
nand U9524 (N_9524,N_3409,N_896);
and U9525 (N_9525,N_2148,N_1462);
and U9526 (N_9526,N_1014,N_70);
and U9527 (N_9527,N_4629,N_4486);
and U9528 (N_9528,N_4645,N_1641);
and U9529 (N_9529,N_1885,N_4056);
nand U9530 (N_9530,N_3449,N_2663);
and U9531 (N_9531,N_402,N_154);
nand U9532 (N_9532,N_3378,N_4906);
nand U9533 (N_9533,N_2481,N_968);
nand U9534 (N_9534,N_4525,N_4644);
xor U9535 (N_9535,N_2398,N_3631);
and U9536 (N_9536,N_2448,N_611);
xor U9537 (N_9537,N_4883,N_4047);
or U9538 (N_9538,N_3099,N_2612);
and U9539 (N_9539,N_3707,N_4304);
nor U9540 (N_9540,N_363,N_1451);
and U9541 (N_9541,N_4756,N_3589);
and U9542 (N_9542,N_1597,N_3941);
xor U9543 (N_9543,N_2148,N_4711);
nand U9544 (N_9544,N_1649,N_4032);
nor U9545 (N_9545,N_3559,N_1100);
and U9546 (N_9546,N_4311,N_4604);
and U9547 (N_9547,N_3468,N_2815);
and U9548 (N_9548,N_3304,N_1130);
and U9549 (N_9549,N_1658,N_1152);
and U9550 (N_9550,N_4578,N_1634);
or U9551 (N_9551,N_957,N_4731);
xnor U9552 (N_9552,N_2370,N_350);
nor U9553 (N_9553,N_1941,N_3663);
and U9554 (N_9554,N_1358,N_1570);
nand U9555 (N_9555,N_4755,N_4892);
nor U9556 (N_9556,N_260,N_432);
nand U9557 (N_9557,N_2305,N_1016);
or U9558 (N_9558,N_2658,N_3818);
nand U9559 (N_9559,N_746,N_4122);
nand U9560 (N_9560,N_3330,N_3545);
xor U9561 (N_9561,N_4668,N_2293);
and U9562 (N_9562,N_1674,N_4436);
xor U9563 (N_9563,N_3482,N_1003);
or U9564 (N_9564,N_2962,N_1418);
or U9565 (N_9565,N_183,N_4887);
nor U9566 (N_9566,N_1292,N_3366);
or U9567 (N_9567,N_2726,N_4293);
nand U9568 (N_9568,N_1718,N_4587);
nand U9569 (N_9569,N_2393,N_123);
or U9570 (N_9570,N_4646,N_4518);
and U9571 (N_9571,N_2642,N_2796);
nor U9572 (N_9572,N_2377,N_3605);
or U9573 (N_9573,N_4955,N_1679);
or U9574 (N_9574,N_3553,N_2511);
nor U9575 (N_9575,N_247,N_994);
nand U9576 (N_9576,N_783,N_4308);
or U9577 (N_9577,N_3881,N_3164);
xor U9578 (N_9578,N_4483,N_1930);
nand U9579 (N_9579,N_1922,N_1010);
and U9580 (N_9580,N_2078,N_4556);
xnor U9581 (N_9581,N_1546,N_1506);
and U9582 (N_9582,N_1908,N_2587);
or U9583 (N_9583,N_4272,N_2161);
xnor U9584 (N_9584,N_4922,N_2210);
nor U9585 (N_9585,N_2326,N_4231);
or U9586 (N_9586,N_4847,N_4463);
and U9587 (N_9587,N_4746,N_1754);
nor U9588 (N_9588,N_2152,N_1417);
nand U9589 (N_9589,N_778,N_3549);
or U9590 (N_9590,N_4945,N_3737);
nor U9591 (N_9591,N_3212,N_881);
or U9592 (N_9592,N_4327,N_323);
or U9593 (N_9593,N_2327,N_4544);
and U9594 (N_9594,N_3261,N_3008);
or U9595 (N_9595,N_1868,N_1580);
nand U9596 (N_9596,N_2543,N_4660);
nor U9597 (N_9597,N_1531,N_4748);
nand U9598 (N_9598,N_3498,N_4643);
or U9599 (N_9599,N_3492,N_534);
or U9600 (N_9600,N_1672,N_3752);
nand U9601 (N_9601,N_4587,N_4352);
and U9602 (N_9602,N_4456,N_2454);
or U9603 (N_9603,N_1356,N_4557);
nor U9604 (N_9604,N_3535,N_108);
nor U9605 (N_9605,N_1488,N_214);
nand U9606 (N_9606,N_2170,N_4720);
nand U9607 (N_9607,N_2032,N_2296);
nor U9608 (N_9608,N_2603,N_4727);
nor U9609 (N_9609,N_1285,N_4667);
nor U9610 (N_9610,N_2632,N_32);
nand U9611 (N_9611,N_4184,N_1811);
nor U9612 (N_9612,N_1330,N_2358);
nand U9613 (N_9613,N_1848,N_1967);
or U9614 (N_9614,N_1406,N_2392);
nand U9615 (N_9615,N_4245,N_4878);
or U9616 (N_9616,N_4244,N_1125);
and U9617 (N_9617,N_505,N_51);
and U9618 (N_9618,N_4149,N_51);
or U9619 (N_9619,N_1674,N_1333);
nor U9620 (N_9620,N_2937,N_3004);
nor U9621 (N_9621,N_498,N_3884);
nor U9622 (N_9622,N_2585,N_3662);
nor U9623 (N_9623,N_2892,N_2417);
nand U9624 (N_9624,N_742,N_2650);
xnor U9625 (N_9625,N_2456,N_4827);
or U9626 (N_9626,N_2009,N_2546);
nand U9627 (N_9627,N_560,N_4350);
nor U9628 (N_9628,N_3994,N_332);
xnor U9629 (N_9629,N_853,N_2337);
xnor U9630 (N_9630,N_3034,N_1959);
xor U9631 (N_9631,N_4423,N_283);
nor U9632 (N_9632,N_3631,N_3377);
nand U9633 (N_9633,N_810,N_4295);
or U9634 (N_9634,N_816,N_285);
nand U9635 (N_9635,N_54,N_3507);
nand U9636 (N_9636,N_782,N_2475);
xor U9637 (N_9637,N_876,N_424);
and U9638 (N_9638,N_1945,N_2166);
and U9639 (N_9639,N_699,N_4546);
and U9640 (N_9640,N_1749,N_3605);
nand U9641 (N_9641,N_1932,N_3366);
xnor U9642 (N_9642,N_4665,N_953);
and U9643 (N_9643,N_3973,N_4918);
nor U9644 (N_9644,N_611,N_1222);
and U9645 (N_9645,N_637,N_2370);
and U9646 (N_9646,N_930,N_2713);
nand U9647 (N_9647,N_3874,N_3032);
nor U9648 (N_9648,N_3085,N_2937);
and U9649 (N_9649,N_3674,N_457);
nor U9650 (N_9650,N_1048,N_2188);
xor U9651 (N_9651,N_4028,N_3859);
and U9652 (N_9652,N_2416,N_4907);
nand U9653 (N_9653,N_411,N_3728);
nor U9654 (N_9654,N_3956,N_374);
or U9655 (N_9655,N_3456,N_2096);
nor U9656 (N_9656,N_2150,N_1422);
xnor U9657 (N_9657,N_647,N_225);
or U9658 (N_9658,N_273,N_385);
nor U9659 (N_9659,N_3501,N_4589);
and U9660 (N_9660,N_4575,N_4454);
and U9661 (N_9661,N_4886,N_3068);
and U9662 (N_9662,N_3810,N_1347);
and U9663 (N_9663,N_3599,N_4346);
and U9664 (N_9664,N_1826,N_4321);
or U9665 (N_9665,N_4974,N_2194);
and U9666 (N_9666,N_2578,N_1860);
nor U9667 (N_9667,N_1104,N_1876);
or U9668 (N_9668,N_3715,N_2694);
nand U9669 (N_9669,N_1098,N_1614);
nor U9670 (N_9670,N_4338,N_2315);
nand U9671 (N_9671,N_4986,N_2233);
xor U9672 (N_9672,N_2777,N_2649);
nand U9673 (N_9673,N_1010,N_495);
and U9674 (N_9674,N_4309,N_322);
nand U9675 (N_9675,N_3586,N_3846);
nand U9676 (N_9676,N_345,N_4966);
and U9677 (N_9677,N_3127,N_4585);
or U9678 (N_9678,N_1046,N_144);
or U9679 (N_9679,N_265,N_3525);
and U9680 (N_9680,N_2420,N_3877);
xnor U9681 (N_9681,N_441,N_422);
and U9682 (N_9682,N_4000,N_63);
nand U9683 (N_9683,N_1930,N_4165);
xnor U9684 (N_9684,N_4763,N_3842);
and U9685 (N_9685,N_4112,N_2346);
nor U9686 (N_9686,N_3981,N_4827);
nand U9687 (N_9687,N_4816,N_1037);
nor U9688 (N_9688,N_1022,N_3386);
and U9689 (N_9689,N_204,N_4633);
nor U9690 (N_9690,N_1697,N_1680);
and U9691 (N_9691,N_2980,N_3312);
or U9692 (N_9692,N_3906,N_2108);
and U9693 (N_9693,N_2132,N_65);
and U9694 (N_9694,N_3192,N_2830);
nor U9695 (N_9695,N_3416,N_1672);
nor U9696 (N_9696,N_3953,N_1966);
nor U9697 (N_9697,N_380,N_1556);
and U9698 (N_9698,N_3449,N_2096);
nand U9699 (N_9699,N_3617,N_3419);
or U9700 (N_9700,N_594,N_1109);
nand U9701 (N_9701,N_1459,N_3355);
or U9702 (N_9702,N_4264,N_1668);
or U9703 (N_9703,N_2452,N_2403);
or U9704 (N_9704,N_1638,N_4237);
or U9705 (N_9705,N_4186,N_2841);
or U9706 (N_9706,N_2832,N_4829);
and U9707 (N_9707,N_914,N_4497);
and U9708 (N_9708,N_1915,N_2437);
nor U9709 (N_9709,N_4048,N_1846);
or U9710 (N_9710,N_2784,N_1791);
or U9711 (N_9711,N_2092,N_1882);
or U9712 (N_9712,N_2707,N_1997);
nor U9713 (N_9713,N_3405,N_1185);
nor U9714 (N_9714,N_3820,N_2113);
or U9715 (N_9715,N_4089,N_2423);
nand U9716 (N_9716,N_2134,N_2676);
and U9717 (N_9717,N_3440,N_2134);
or U9718 (N_9718,N_958,N_1064);
nor U9719 (N_9719,N_639,N_292);
or U9720 (N_9720,N_2705,N_282);
and U9721 (N_9721,N_3390,N_2526);
or U9722 (N_9722,N_2399,N_4179);
and U9723 (N_9723,N_4048,N_3475);
nand U9724 (N_9724,N_2549,N_2793);
xor U9725 (N_9725,N_4254,N_4687);
xnor U9726 (N_9726,N_4375,N_3523);
nor U9727 (N_9727,N_2501,N_2488);
and U9728 (N_9728,N_4500,N_1185);
and U9729 (N_9729,N_1584,N_2006);
nand U9730 (N_9730,N_512,N_391);
nand U9731 (N_9731,N_162,N_3650);
and U9732 (N_9732,N_3547,N_376);
and U9733 (N_9733,N_4952,N_160);
and U9734 (N_9734,N_2247,N_2547);
nand U9735 (N_9735,N_1744,N_1304);
or U9736 (N_9736,N_3333,N_132);
or U9737 (N_9737,N_644,N_4929);
nor U9738 (N_9738,N_1832,N_991);
nand U9739 (N_9739,N_4080,N_27);
nor U9740 (N_9740,N_3877,N_2371);
xor U9741 (N_9741,N_1837,N_1522);
or U9742 (N_9742,N_3889,N_244);
nand U9743 (N_9743,N_2004,N_2168);
nor U9744 (N_9744,N_2006,N_4468);
nand U9745 (N_9745,N_1151,N_3903);
nand U9746 (N_9746,N_434,N_4505);
or U9747 (N_9747,N_1864,N_4838);
and U9748 (N_9748,N_2380,N_4920);
nor U9749 (N_9749,N_577,N_252);
and U9750 (N_9750,N_403,N_2148);
xor U9751 (N_9751,N_73,N_3153);
nand U9752 (N_9752,N_154,N_3548);
or U9753 (N_9753,N_4082,N_3805);
and U9754 (N_9754,N_1115,N_1156);
or U9755 (N_9755,N_3006,N_2883);
and U9756 (N_9756,N_2129,N_1881);
nor U9757 (N_9757,N_4033,N_460);
nand U9758 (N_9758,N_3309,N_429);
and U9759 (N_9759,N_3504,N_3572);
or U9760 (N_9760,N_2837,N_1854);
or U9761 (N_9761,N_650,N_1166);
nor U9762 (N_9762,N_838,N_4524);
nor U9763 (N_9763,N_1767,N_3466);
and U9764 (N_9764,N_4423,N_512);
nor U9765 (N_9765,N_1870,N_3846);
nor U9766 (N_9766,N_2648,N_3944);
nor U9767 (N_9767,N_1206,N_3815);
or U9768 (N_9768,N_1898,N_4111);
or U9769 (N_9769,N_1392,N_3556);
nor U9770 (N_9770,N_1970,N_2846);
or U9771 (N_9771,N_1918,N_1105);
or U9772 (N_9772,N_3188,N_725);
or U9773 (N_9773,N_2978,N_2393);
and U9774 (N_9774,N_2244,N_956);
nand U9775 (N_9775,N_2615,N_3977);
xor U9776 (N_9776,N_2071,N_659);
nand U9777 (N_9777,N_2429,N_4378);
and U9778 (N_9778,N_4328,N_4149);
xor U9779 (N_9779,N_3997,N_2303);
xor U9780 (N_9780,N_1458,N_210);
or U9781 (N_9781,N_3735,N_3363);
or U9782 (N_9782,N_1860,N_4814);
nor U9783 (N_9783,N_2843,N_318);
nand U9784 (N_9784,N_505,N_2733);
or U9785 (N_9785,N_1351,N_1998);
nand U9786 (N_9786,N_1981,N_2719);
or U9787 (N_9787,N_154,N_4828);
xnor U9788 (N_9788,N_1403,N_2880);
nand U9789 (N_9789,N_906,N_1826);
nand U9790 (N_9790,N_639,N_1786);
nor U9791 (N_9791,N_3680,N_804);
nand U9792 (N_9792,N_3684,N_419);
or U9793 (N_9793,N_1201,N_4339);
nor U9794 (N_9794,N_4223,N_3190);
nand U9795 (N_9795,N_1598,N_3792);
or U9796 (N_9796,N_594,N_3155);
nor U9797 (N_9797,N_3444,N_4394);
or U9798 (N_9798,N_2103,N_3678);
nand U9799 (N_9799,N_2955,N_1015);
nand U9800 (N_9800,N_4935,N_4866);
xnor U9801 (N_9801,N_2916,N_710);
nor U9802 (N_9802,N_4275,N_4590);
nor U9803 (N_9803,N_3980,N_1487);
nor U9804 (N_9804,N_346,N_4412);
nand U9805 (N_9805,N_328,N_863);
nand U9806 (N_9806,N_2577,N_4072);
nand U9807 (N_9807,N_4650,N_1556);
nor U9808 (N_9808,N_4295,N_107);
or U9809 (N_9809,N_2626,N_2258);
and U9810 (N_9810,N_1403,N_4914);
and U9811 (N_9811,N_1169,N_2578);
and U9812 (N_9812,N_2375,N_3775);
or U9813 (N_9813,N_3477,N_3544);
nor U9814 (N_9814,N_4399,N_125);
nand U9815 (N_9815,N_4214,N_4419);
or U9816 (N_9816,N_3530,N_3735);
nor U9817 (N_9817,N_3051,N_1881);
or U9818 (N_9818,N_1429,N_51);
nand U9819 (N_9819,N_1484,N_4819);
nor U9820 (N_9820,N_564,N_3103);
and U9821 (N_9821,N_2391,N_1662);
or U9822 (N_9822,N_2490,N_4345);
nor U9823 (N_9823,N_1812,N_4884);
nor U9824 (N_9824,N_3778,N_1282);
nand U9825 (N_9825,N_3445,N_3092);
nand U9826 (N_9826,N_1451,N_2257);
nor U9827 (N_9827,N_1106,N_2093);
xor U9828 (N_9828,N_437,N_4591);
nand U9829 (N_9829,N_4049,N_565);
and U9830 (N_9830,N_3155,N_977);
nand U9831 (N_9831,N_3592,N_2056);
nand U9832 (N_9832,N_2132,N_994);
or U9833 (N_9833,N_2354,N_4136);
nor U9834 (N_9834,N_2396,N_3649);
xnor U9835 (N_9835,N_2434,N_2907);
and U9836 (N_9836,N_3077,N_2054);
or U9837 (N_9837,N_3392,N_1194);
or U9838 (N_9838,N_55,N_4925);
and U9839 (N_9839,N_1657,N_3623);
xnor U9840 (N_9840,N_4596,N_2524);
xnor U9841 (N_9841,N_2978,N_4923);
nor U9842 (N_9842,N_2077,N_3275);
nor U9843 (N_9843,N_4058,N_1041);
nand U9844 (N_9844,N_1504,N_3109);
or U9845 (N_9845,N_509,N_3405);
or U9846 (N_9846,N_212,N_4802);
nand U9847 (N_9847,N_168,N_4015);
or U9848 (N_9848,N_699,N_439);
nand U9849 (N_9849,N_4092,N_380);
nand U9850 (N_9850,N_4542,N_4728);
or U9851 (N_9851,N_3810,N_2263);
nand U9852 (N_9852,N_413,N_3093);
nand U9853 (N_9853,N_3468,N_3184);
nor U9854 (N_9854,N_3197,N_4840);
or U9855 (N_9855,N_2771,N_1119);
nor U9856 (N_9856,N_2928,N_2272);
and U9857 (N_9857,N_3752,N_4428);
or U9858 (N_9858,N_3039,N_2909);
or U9859 (N_9859,N_3315,N_4958);
and U9860 (N_9860,N_4310,N_2712);
and U9861 (N_9861,N_4364,N_2099);
or U9862 (N_9862,N_2728,N_2453);
or U9863 (N_9863,N_1461,N_1165);
nor U9864 (N_9864,N_2238,N_341);
and U9865 (N_9865,N_95,N_3595);
nand U9866 (N_9866,N_3201,N_1298);
nor U9867 (N_9867,N_4980,N_3934);
and U9868 (N_9868,N_2419,N_2624);
nand U9869 (N_9869,N_2314,N_4244);
xor U9870 (N_9870,N_2198,N_3300);
or U9871 (N_9871,N_3015,N_4678);
or U9872 (N_9872,N_1855,N_1743);
or U9873 (N_9873,N_2570,N_2172);
or U9874 (N_9874,N_4728,N_2032);
nor U9875 (N_9875,N_3792,N_3990);
nand U9876 (N_9876,N_3863,N_4652);
xnor U9877 (N_9877,N_1265,N_3268);
nand U9878 (N_9878,N_3924,N_2631);
nor U9879 (N_9879,N_1082,N_2110);
or U9880 (N_9880,N_204,N_3762);
or U9881 (N_9881,N_4699,N_2275);
nor U9882 (N_9882,N_4599,N_1965);
nand U9883 (N_9883,N_1866,N_1325);
or U9884 (N_9884,N_2881,N_1563);
nor U9885 (N_9885,N_633,N_2708);
nor U9886 (N_9886,N_3639,N_2960);
nor U9887 (N_9887,N_3951,N_4880);
nand U9888 (N_9888,N_1713,N_4298);
nor U9889 (N_9889,N_977,N_1576);
nor U9890 (N_9890,N_4241,N_4672);
nor U9891 (N_9891,N_4459,N_4229);
nor U9892 (N_9892,N_4758,N_3561);
or U9893 (N_9893,N_4783,N_2080);
or U9894 (N_9894,N_867,N_2060);
xnor U9895 (N_9895,N_3294,N_4807);
nor U9896 (N_9896,N_364,N_1546);
nor U9897 (N_9897,N_405,N_4889);
nand U9898 (N_9898,N_3541,N_4099);
or U9899 (N_9899,N_4780,N_3415);
or U9900 (N_9900,N_2024,N_913);
nand U9901 (N_9901,N_4972,N_696);
and U9902 (N_9902,N_1943,N_4374);
and U9903 (N_9903,N_3319,N_4931);
nand U9904 (N_9904,N_1899,N_3105);
nor U9905 (N_9905,N_68,N_4918);
and U9906 (N_9906,N_2633,N_1882);
nor U9907 (N_9907,N_4736,N_4794);
or U9908 (N_9908,N_2010,N_2112);
nor U9909 (N_9909,N_4255,N_2971);
and U9910 (N_9910,N_2415,N_3366);
and U9911 (N_9911,N_3824,N_3213);
nand U9912 (N_9912,N_2632,N_2327);
nand U9913 (N_9913,N_507,N_2058);
xnor U9914 (N_9914,N_2565,N_2391);
or U9915 (N_9915,N_2263,N_4666);
xor U9916 (N_9916,N_1918,N_3468);
nor U9917 (N_9917,N_173,N_1782);
nor U9918 (N_9918,N_3728,N_4343);
nor U9919 (N_9919,N_615,N_1649);
nor U9920 (N_9920,N_2750,N_575);
and U9921 (N_9921,N_2346,N_2105);
nand U9922 (N_9922,N_3672,N_1891);
nand U9923 (N_9923,N_4880,N_1239);
nand U9924 (N_9924,N_4001,N_3631);
or U9925 (N_9925,N_3897,N_4616);
and U9926 (N_9926,N_2529,N_837);
nor U9927 (N_9927,N_4754,N_1874);
nor U9928 (N_9928,N_2800,N_1534);
nor U9929 (N_9929,N_3742,N_4931);
nand U9930 (N_9930,N_1824,N_304);
and U9931 (N_9931,N_4541,N_4070);
nand U9932 (N_9932,N_4366,N_3658);
nand U9933 (N_9933,N_3701,N_736);
and U9934 (N_9934,N_3901,N_1260);
and U9935 (N_9935,N_3996,N_4401);
and U9936 (N_9936,N_3345,N_4528);
nand U9937 (N_9937,N_899,N_149);
or U9938 (N_9938,N_600,N_674);
xor U9939 (N_9939,N_2183,N_3632);
or U9940 (N_9940,N_1403,N_1475);
nor U9941 (N_9941,N_3301,N_4483);
xor U9942 (N_9942,N_966,N_2737);
nand U9943 (N_9943,N_295,N_4051);
nand U9944 (N_9944,N_284,N_872);
or U9945 (N_9945,N_1548,N_3711);
nand U9946 (N_9946,N_4592,N_2021);
or U9947 (N_9947,N_4653,N_978);
or U9948 (N_9948,N_57,N_1937);
nand U9949 (N_9949,N_1579,N_3231);
or U9950 (N_9950,N_662,N_1348);
and U9951 (N_9951,N_2411,N_3037);
nand U9952 (N_9952,N_2375,N_4276);
nor U9953 (N_9953,N_2399,N_4181);
or U9954 (N_9954,N_4274,N_3608);
or U9955 (N_9955,N_1021,N_3644);
nor U9956 (N_9956,N_994,N_809);
and U9957 (N_9957,N_1417,N_2467);
or U9958 (N_9958,N_4830,N_4739);
or U9959 (N_9959,N_1497,N_1787);
and U9960 (N_9960,N_606,N_66);
and U9961 (N_9961,N_2691,N_3267);
and U9962 (N_9962,N_1006,N_3166);
nand U9963 (N_9963,N_1998,N_4471);
xnor U9964 (N_9964,N_2341,N_4133);
nand U9965 (N_9965,N_1804,N_1638);
xor U9966 (N_9966,N_2318,N_413);
xnor U9967 (N_9967,N_298,N_793);
or U9968 (N_9968,N_2516,N_2911);
nand U9969 (N_9969,N_2334,N_2822);
or U9970 (N_9970,N_111,N_2095);
nand U9971 (N_9971,N_4298,N_3137);
nor U9972 (N_9972,N_660,N_3053);
and U9973 (N_9973,N_3313,N_1200);
nand U9974 (N_9974,N_4623,N_986);
or U9975 (N_9975,N_3887,N_2774);
and U9976 (N_9976,N_3711,N_4750);
nand U9977 (N_9977,N_236,N_4370);
and U9978 (N_9978,N_4166,N_3082);
xor U9979 (N_9979,N_1219,N_1324);
xor U9980 (N_9980,N_4564,N_3015);
and U9981 (N_9981,N_4262,N_2446);
xnor U9982 (N_9982,N_3518,N_481);
and U9983 (N_9983,N_185,N_3343);
or U9984 (N_9984,N_3996,N_1089);
nand U9985 (N_9985,N_4762,N_28);
or U9986 (N_9986,N_2460,N_4485);
nor U9987 (N_9987,N_2901,N_1916);
nand U9988 (N_9988,N_58,N_502);
nand U9989 (N_9989,N_4778,N_2291);
or U9990 (N_9990,N_2325,N_1645);
nor U9991 (N_9991,N_2760,N_2752);
nand U9992 (N_9992,N_1475,N_1331);
nor U9993 (N_9993,N_4837,N_2571);
xnor U9994 (N_9994,N_1505,N_4194);
and U9995 (N_9995,N_4535,N_2643);
or U9996 (N_9996,N_4497,N_999);
or U9997 (N_9997,N_4328,N_2844);
nand U9998 (N_9998,N_905,N_1005);
nor U9999 (N_9999,N_1711,N_2427);
and U10000 (N_10000,N_7553,N_7233);
and U10001 (N_10001,N_8665,N_6665);
nor U10002 (N_10002,N_8003,N_6975);
xor U10003 (N_10003,N_9587,N_6547);
or U10004 (N_10004,N_6143,N_9571);
and U10005 (N_10005,N_7745,N_8105);
and U10006 (N_10006,N_8161,N_8765);
and U10007 (N_10007,N_9973,N_5689);
and U10008 (N_10008,N_8044,N_8096);
or U10009 (N_10009,N_6062,N_9225);
nor U10010 (N_10010,N_9492,N_8602);
or U10011 (N_10011,N_5981,N_6429);
xnor U10012 (N_10012,N_7965,N_7242);
and U10013 (N_10013,N_8787,N_9490);
nand U10014 (N_10014,N_5439,N_5279);
nor U10015 (N_10015,N_6255,N_5743);
and U10016 (N_10016,N_7825,N_6059);
or U10017 (N_10017,N_9299,N_7260);
nand U10018 (N_10018,N_6057,N_6859);
nand U10019 (N_10019,N_8842,N_9643);
xnor U10020 (N_10020,N_8738,N_6477);
and U10021 (N_10021,N_8658,N_7528);
nand U10022 (N_10022,N_7775,N_5301);
or U10023 (N_10023,N_5566,N_7299);
xnor U10024 (N_10024,N_9155,N_7157);
nor U10025 (N_10025,N_9339,N_8009);
or U10026 (N_10026,N_7339,N_5309);
and U10027 (N_10027,N_9873,N_5433);
nor U10028 (N_10028,N_9807,N_7283);
and U10029 (N_10029,N_9043,N_7262);
or U10030 (N_10030,N_9397,N_9217);
nand U10031 (N_10031,N_7342,N_6948);
nand U10032 (N_10032,N_6878,N_9906);
nor U10033 (N_10033,N_9250,N_9683);
or U10034 (N_10034,N_7420,N_7143);
or U10035 (N_10035,N_6371,N_7959);
nor U10036 (N_10036,N_6598,N_8021);
nand U10037 (N_10037,N_7802,N_7888);
xor U10038 (N_10038,N_7414,N_5174);
nor U10039 (N_10039,N_7987,N_7990);
and U10040 (N_10040,N_5485,N_7708);
or U10041 (N_10041,N_8501,N_8784);
nand U10042 (N_10042,N_5907,N_7798);
nor U10043 (N_10043,N_9540,N_9083);
nand U10044 (N_10044,N_5809,N_9495);
or U10045 (N_10045,N_9528,N_7711);
nand U10046 (N_10046,N_8715,N_5274);
nand U10047 (N_10047,N_6799,N_5448);
or U10048 (N_10048,N_7218,N_6289);
xnor U10049 (N_10049,N_7874,N_7464);
nor U10050 (N_10050,N_6258,N_9939);
and U10051 (N_10051,N_9150,N_7063);
nor U10052 (N_10052,N_9201,N_7939);
and U10053 (N_10053,N_8213,N_6712);
or U10054 (N_10054,N_9343,N_5357);
nor U10055 (N_10055,N_7899,N_7168);
xnor U10056 (N_10056,N_6783,N_6296);
or U10057 (N_10057,N_9669,N_5685);
xnor U10058 (N_10058,N_9472,N_7633);
and U10059 (N_10059,N_9538,N_9197);
nand U10060 (N_10060,N_9936,N_9519);
or U10061 (N_10061,N_5478,N_5952);
and U10062 (N_10062,N_9488,N_6067);
nand U10063 (N_10063,N_9967,N_8831);
nand U10064 (N_10064,N_5782,N_8557);
nor U10065 (N_10065,N_7497,N_8865);
nor U10066 (N_10066,N_8091,N_5479);
or U10067 (N_10067,N_5970,N_8795);
nor U10068 (N_10068,N_8004,N_6071);
nor U10069 (N_10069,N_5994,N_6733);
nor U10070 (N_10070,N_8996,N_5386);
or U10071 (N_10071,N_8440,N_5823);
or U10072 (N_10072,N_9458,N_8500);
nor U10073 (N_10073,N_5169,N_6807);
and U10074 (N_10074,N_9626,N_5781);
nor U10075 (N_10075,N_8172,N_8099);
and U10076 (N_10076,N_9696,N_8456);
nand U10077 (N_10077,N_6877,N_8809);
or U10078 (N_10078,N_6624,N_8546);
nand U10079 (N_10079,N_6595,N_9286);
and U10080 (N_10080,N_7270,N_9752);
and U10081 (N_10081,N_6747,N_6970);
or U10082 (N_10082,N_6374,N_5061);
and U10083 (N_10083,N_8540,N_9303);
nor U10084 (N_10084,N_7183,N_9029);
and U10085 (N_10085,N_6239,N_5855);
and U10086 (N_10086,N_8821,N_5385);
nand U10087 (N_10087,N_9118,N_7125);
or U10088 (N_10088,N_7228,N_5872);
nand U10089 (N_10089,N_9822,N_9287);
xor U10090 (N_10090,N_5260,N_9269);
and U10091 (N_10091,N_9414,N_5463);
nand U10092 (N_10092,N_9819,N_9653);
nand U10093 (N_10093,N_7510,N_5741);
nand U10094 (N_10094,N_9642,N_5161);
nor U10095 (N_10095,N_9173,N_7467);
nor U10096 (N_10096,N_5567,N_9985);
and U10097 (N_10097,N_8010,N_7118);
nor U10098 (N_10098,N_8428,N_8049);
nor U10099 (N_10099,N_8116,N_5103);
xnor U10100 (N_10100,N_8683,N_5012);
nand U10101 (N_10101,N_8356,N_9417);
xnor U10102 (N_10102,N_7127,N_7541);
or U10103 (N_10103,N_8164,N_8539);
nor U10104 (N_10104,N_9026,N_5793);
nand U10105 (N_10105,N_7818,N_6197);
nand U10106 (N_10106,N_6999,N_5946);
nor U10107 (N_10107,N_7855,N_5514);
nand U10108 (N_10108,N_7515,N_9394);
and U10109 (N_10109,N_6209,N_8047);
and U10110 (N_10110,N_9534,N_7456);
and U10111 (N_10111,N_5575,N_9360);
and U10112 (N_10112,N_8297,N_6698);
nand U10113 (N_10113,N_9881,N_7132);
nand U10114 (N_10114,N_7694,N_5461);
nand U10115 (N_10115,N_9570,N_5978);
xnor U10116 (N_10116,N_8930,N_6885);
nand U10117 (N_10117,N_5421,N_8413);
and U10118 (N_10118,N_8818,N_5954);
xor U10119 (N_10119,N_5966,N_8200);
and U10120 (N_10120,N_6927,N_6512);
and U10121 (N_10121,N_5602,N_9236);
nor U10122 (N_10122,N_6575,N_8187);
nand U10123 (N_10123,N_5430,N_8774);
xor U10124 (N_10124,N_9659,N_5960);
xor U10125 (N_10125,N_6757,N_6043);
xnor U10126 (N_10126,N_8945,N_8654);
nand U10127 (N_10127,N_8574,N_6623);
nand U10128 (N_10128,N_6250,N_7814);
xnor U10129 (N_10129,N_8701,N_8534);
nor U10130 (N_10130,N_9148,N_6246);
nor U10131 (N_10131,N_9410,N_6883);
and U10132 (N_10132,N_7116,N_7551);
nand U10133 (N_10133,N_7376,N_7101);
nand U10134 (N_10134,N_5880,N_7423);
nor U10135 (N_10135,N_8670,N_9905);
nor U10136 (N_10136,N_9529,N_7377);
xor U10137 (N_10137,N_8875,N_5917);
nor U10138 (N_10138,N_8035,N_5121);
or U10139 (N_10139,N_5024,N_6338);
and U10140 (N_10140,N_5064,N_9419);
and U10141 (N_10141,N_9937,N_8320);
nor U10142 (N_10142,N_8901,N_5411);
and U10143 (N_10143,N_9176,N_8580);
and U10144 (N_10144,N_8008,N_8569);
nand U10145 (N_10145,N_8823,N_8472);
nand U10146 (N_10146,N_7369,N_8314);
or U10147 (N_10147,N_8308,N_7120);
or U10148 (N_10148,N_8438,N_9969);
and U10149 (N_10149,N_8754,N_5246);
or U10150 (N_10150,N_6847,N_5520);
and U10151 (N_10151,N_9992,N_9221);
and U10152 (N_10152,N_9087,N_5340);
nand U10153 (N_10153,N_9787,N_5480);
nand U10154 (N_10154,N_7506,N_6987);
nand U10155 (N_10155,N_8951,N_9063);
nor U10156 (N_10156,N_7858,N_6179);
nor U10157 (N_10157,N_5863,N_9849);
or U10158 (N_10158,N_6039,N_8169);
and U10159 (N_10159,N_5968,N_5539);
or U10160 (N_10160,N_7252,N_7220);
nand U10161 (N_10161,N_9756,N_7668);
and U10162 (N_10162,N_7549,N_7759);
or U10163 (N_10163,N_9632,N_7454);
nand U10164 (N_10164,N_8327,N_8730);
or U10165 (N_10165,N_5353,N_5808);
nor U10166 (N_10166,N_6169,N_7636);
nand U10167 (N_10167,N_8081,N_5194);
nor U10168 (N_10168,N_6633,N_7623);
and U10169 (N_10169,N_6366,N_8118);
nand U10170 (N_10170,N_9815,N_6928);
xnor U10171 (N_10171,N_6639,N_6774);
nor U10172 (N_10172,N_8202,N_7459);
and U10173 (N_10173,N_5010,N_5755);
nand U10174 (N_10174,N_9098,N_5687);
xor U10175 (N_10175,N_7209,N_9987);
nand U10176 (N_10176,N_7196,N_9412);
or U10177 (N_10177,N_6777,N_9172);
or U10178 (N_10178,N_9651,N_6666);
or U10179 (N_10179,N_9550,N_7854);
and U10180 (N_10180,N_9341,N_7882);
and U10181 (N_10181,N_6470,N_7169);
and U10182 (N_10182,N_9837,N_9091);
nand U10183 (N_10183,N_8043,N_9289);
nand U10184 (N_10184,N_5344,N_7630);
nor U10185 (N_10185,N_7522,N_6709);
or U10186 (N_10186,N_6044,N_6051);
or U10187 (N_10187,N_8289,N_6533);
or U10188 (N_10188,N_6714,N_5071);
xor U10189 (N_10189,N_8903,N_5066);
nand U10190 (N_10190,N_9180,N_8847);
or U10191 (N_10191,N_6858,N_5920);
nor U10192 (N_10192,N_9437,N_8068);
nor U10193 (N_10193,N_5720,N_9588);
xor U10194 (N_10194,N_8231,N_7883);
xnor U10195 (N_10195,N_6327,N_6375);
and U10196 (N_10196,N_5371,N_9629);
nor U10197 (N_10197,N_5653,N_6861);
and U10198 (N_10198,N_5556,N_5234);
nor U10199 (N_10199,N_9797,N_7500);
nand U10200 (N_10200,N_9102,N_7960);
nor U10201 (N_10201,N_6579,N_7344);
and U10202 (N_10202,N_5155,N_7792);
nand U10203 (N_10203,N_8732,N_5664);
and U10204 (N_10204,N_9989,N_9486);
nor U10205 (N_10205,N_8175,N_8562);
nor U10206 (N_10206,N_7834,N_9684);
nand U10207 (N_10207,N_5098,N_9230);
and U10208 (N_10208,N_9443,N_7057);
or U10209 (N_10209,N_7128,N_9609);
nor U10210 (N_10210,N_5454,N_5762);
nand U10211 (N_10211,N_7455,N_7554);
nor U10212 (N_10212,N_7019,N_9170);
or U10213 (N_10213,N_5495,N_8245);
or U10214 (N_10214,N_5402,N_6136);
and U10215 (N_10215,N_5395,N_8740);
nand U10216 (N_10216,N_6577,N_9578);
nand U10217 (N_10217,N_7176,N_6290);
and U10218 (N_10218,N_8958,N_5891);
or U10219 (N_10219,N_9845,N_7383);
nand U10220 (N_10220,N_7017,N_5325);
and U10221 (N_10221,N_5468,N_9135);
and U10222 (N_10222,N_7331,N_9457);
nor U10223 (N_10223,N_5204,N_6850);
xnor U10224 (N_10224,N_5362,N_6875);
and U10225 (N_10225,N_8249,N_6362);
and U10226 (N_10226,N_6114,N_9060);
nand U10227 (N_10227,N_8931,N_8643);
and U10228 (N_10228,N_5936,N_9882);
nand U10229 (N_10229,N_8535,N_9853);
nand U10230 (N_10230,N_5022,N_8444);
nor U10231 (N_10231,N_9470,N_6393);
and U10232 (N_10232,N_8114,N_8647);
nor U10233 (N_10233,N_8728,N_6347);
nand U10234 (N_10234,N_5959,N_9335);
or U10235 (N_10235,N_9715,N_9884);
nor U10236 (N_10236,N_7763,N_6635);
nand U10237 (N_10237,N_8817,N_9071);
and U10238 (N_10238,N_8712,N_9446);
nand U10239 (N_10239,N_5216,N_9051);
or U10240 (N_10240,N_7167,N_9961);
and U10241 (N_10241,N_8642,N_5899);
xor U10242 (N_10242,N_8064,N_8837);
xor U10243 (N_10243,N_5323,N_5562);
nor U10244 (N_10244,N_9056,N_8461);
nor U10245 (N_10245,N_9163,N_9793);
nand U10246 (N_10246,N_8625,N_7483);
nor U10247 (N_10247,N_7947,N_6590);
nand U10248 (N_10248,N_6520,N_7698);
or U10249 (N_10249,N_7654,N_6700);
or U10250 (N_10250,N_8007,N_7583);
and U10251 (N_10251,N_5987,N_5571);
nor U10252 (N_10252,N_7637,N_6430);
nor U10253 (N_10253,N_5504,N_6804);
and U10254 (N_10254,N_9292,N_8352);
xor U10255 (N_10255,N_5476,N_9976);
nor U10256 (N_10256,N_7096,N_6205);
xor U10257 (N_10257,N_6616,N_9031);
and U10258 (N_10258,N_7393,N_9551);
nand U10259 (N_10259,N_7389,N_8362);
nand U10260 (N_10260,N_8229,N_7785);
nand U10261 (N_10261,N_7461,N_9321);
or U10262 (N_10262,N_8190,N_7417);
and U10263 (N_10263,N_9547,N_6415);
nand U10264 (N_10264,N_8361,N_8707);
nor U10265 (N_10265,N_7392,N_8056);
nand U10266 (N_10266,N_7829,N_6103);
and U10267 (N_10267,N_8688,N_7719);
or U10268 (N_10268,N_5841,N_5700);
nand U10269 (N_10269,N_9982,N_9034);
nor U10270 (N_10270,N_9999,N_8347);
nor U10271 (N_10271,N_8490,N_5735);
nor U10272 (N_10272,N_5014,N_9861);
and U10273 (N_10273,N_8640,N_5488);
nor U10274 (N_10274,N_5135,N_5815);
nand U10275 (N_10275,N_6706,N_6284);
nand U10276 (N_10276,N_5063,N_5701);
and U10277 (N_10277,N_9154,N_9352);
and U10278 (N_10278,N_7511,N_8988);
nor U10279 (N_10279,N_9010,N_6066);
or U10280 (N_10280,N_6405,N_6110);
and U10281 (N_10281,N_9854,N_6125);
and U10282 (N_10282,N_6278,N_5965);
and U10283 (N_10283,N_7879,N_6846);
and U10284 (N_10284,N_8702,N_5189);
nand U10285 (N_10285,N_5242,N_8078);
nor U10286 (N_10286,N_6560,N_9650);
nand U10287 (N_10287,N_6176,N_5472);
nor U10288 (N_10288,N_9070,N_6812);
and U10289 (N_10289,N_7893,N_9549);
nand U10290 (N_10290,N_9582,N_7475);
and U10291 (N_10291,N_9860,N_7535);
nor U10292 (N_10292,N_5695,N_6619);
nand U10293 (N_10293,N_7673,N_5572);
or U10294 (N_10294,N_6550,N_6569);
nand U10295 (N_10295,N_5890,N_5541);
and U10296 (N_10296,N_9189,N_5941);
xnor U10297 (N_10297,N_8354,N_6450);
or U10298 (N_10298,N_8850,N_5453);
nand U10299 (N_10299,N_8946,N_8504);
or U10300 (N_10300,N_9466,N_5606);
nor U10301 (N_10301,N_5191,N_6782);
and U10302 (N_10302,N_5142,N_6283);
or U10303 (N_10303,N_8492,N_7146);
xor U10304 (N_10304,N_5412,N_9991);
nor U10305 (N_10305,N_6187,N_5914);
nor U10306 (N_10306,N_5069,N_7737);
and U10307 (N_10307,N_6391,N_5903);
nand U10308 (N_10308,N_8416,N_5766);
nor U10309 (N_10309,N_5122,N_9656);
and U10310 (N_10310,N_9479,N_5141);
and U10311 (N_10311,N_5982,N_5086);
or U10312 (N_10312,N_5679,N_9315);
nor U10313 (N_10313,N_7486,N_5087);
nor U10314 (N_10314,N_5106,N_5549);
and U10315 (N_10315,N_7022,N_8090);
nor U10316 (N_10316,N_9398,N_6135);
and U10317 (N_10317,N_9400,N_6823);
nand U10318 (N_10318,N_6944,N_6832);
xor U10319 (N_10319,N_5585,N_5662);
and U10320 (N_10320,N_8531,N_6126);
nand U10321 (N_10321,N_9366,N_6682);
nand U10322 (N_10322,N_9762,N_5996);
or U10323 (N_10323,N_8247,N_9858);
nand U10324 (N_10324,N_9866,N_9776);
nand U10325 (N_10325,N_5202,N_7624);
nand U10326 (N_10326,N_8267,N_8209);
nand U10327 (N_10327,N_5600,N_7170);
nor U10328 (N_10328,N_7838,N_9838);
or U10329 (N_10329,N_5916,N_9726);
and U10330 (N_10330,N_7223,N_8384);
or U10331 (N_10331,N_6012,N_7171);
or U10332 (N_10332,N_5338,N_5082);
and U10333 (N_10333,N_7532,N_7325);
nand U10334 (N_10334,N_6662,N_8620);
or U10335 (N_10335,N_5108,N_9892);
nor U10336 (N_10336,N_5257,N_9260);
and U10337 (N_10337,N_6215,N_5641);
xor U10338 (N_10338,N_6701,N_6626);
or U10339 (N_10339,N_6552,N_5032);
and U10340 (N_10340,N_7362,N_6089);
or U10341 (N_10341,N_9962,N_7150);
nor U10342 (N_10342,N_6522,N_8893);
or U10343 (N_10343,N_5302,N_8756);
or U10344 (N_10344,N_8139,N_9137);
nand U10345 (N_10345,N_7920,N_6177);
nor U10346 (N_10346,N_9140,N_7064);
or U10347 (N_10347,N_8537,N_5898);
and U10348 (N_10348,N_9688,N_6383);
nor U10349 (N_10349,N_8855,N_9621);
or U10350 (N_10350,N_7749,N_5991);
and U10351 (N_10351,N_8884,N_7867);
and U10352 (N_10352,N_9872,N_8826);
or U10353 (N_10353,N_8455,N_6922);
or U10354 (N_10354,N_6266,N_5626);
and U10355 (N_10355,N_7786,N_9298);
or U10356 (N_10356,N_8019,N_6866);
nor U10357 (N_10357,N_9978,N_9218);
nand U10358 (N_10358,N_9660,N_7027);
nor U10359 (N_10359,N_6868,N_6485);
nor U10360 (N_10360,N_9062,N_5530);
nand U10361 (N_10361,N_6449,N_9789);
nor U10362 (N_10362,N_7876,N_9790);
nor U10363 (N_10363,N_9532,N_6815);
and U10364 (N_10364,N_5774,N_9206);
xor U10365 (N_10365,N_8879,N_8508);
or U10366 (N_10366,N_9891,N_5151);
nand U10367 (N_10367,N_7021,N_9947);
and U10368 (N_10368,N_7738,N_9001);
nand U10369 (N_10369,N_5055,N_9243);
nand U10370 (N_10370,N_8374,N_6335);
and U10371 (N_10371,N_6705,N_6459);
or U10372 (N_10372,N_6913,N_9259);
or U10373 (N_10373,N_8517,N_7665);
xnor U10374 (N_10374,N_6687,N_7296);
or U10375 (N_10375,N_6149,N_7783);
nor U10376 (N_10376,N_5699,N_5772);
or U10377 (N_10377,N_7887,N_7368);
and U10378 (N_10378,N_9003,N_7353);
or U10379 (N_10379,N_5243,N_6504);
nand U10380 (N_10380,N_6117,N_5788);
nor U10381 (N_10381,N_5590,N_8813);
nand U10382 (N_10382,N_5578,N_9317);
nand U10383 (N_10383,N_7762,N_6989);
or U10384 (N_10384,N_6995,N_6910);
nand U10385 (N_10385,N_8952,N_5975);
nand U10386 (N_10386,N_6498,N_6033);
nand U10387 (N_10387,N_8146,N_7330);
xor U10388 (N_10388,N_5401,N_7797);
xor U10389 (N_10389,N_6958,N_8564);
nand U10390 (N_10390,N_8572,N_7134);
nor U10391 (N_10391,N_8418,N_9313);
nand U10392 (N_10392,N_5080,N_5310);
xor U10393 (N_10393,N_5535,N_8991);
nand U10394 (N_10394,N_7370,N_5526);
nand U10395 (N_10395,N_7687,N_5640);
nand U10396 (N_10396,N_6088,N_7787);
and U10397 (N_10397,N_7225,N_8538);
nand U10398 (N_10398,N_7133,N_9302);
and U10399 (N_10399,N_8196,N_5674);
nand U10400 (N_10400,N_6792,N_6882);
and U10401 (N_10401,N_7030,N_7755);
nand U10402 (N_10402,N_9624,N_8167);
and U10403 (N_10403,N_7277,N_9145);
nor U10404 (N_10404,N_7560,N_6681);
nand U10405 (N_10405,N_9052,N_6399);
and U10406 (N_10406,N_8124,N_7436);
nand U10407 (N_10407,N_6786,N_7255);
and U10408 (N_10408,N_8706,N_6082);
and U10409 (N_10409,N_6896,N_6940);
xor U10410 (N_10410,N_6398,N_5584);
xor U10411 (N_10411,N_5493,N_9185);
or U10412 (N_10412,N_8197,N_8807);
nand U10413 (N_10413,N_5949,N_7943);
and U10414 (N_10414,N_7265,N_9627);
nand U10415 (N_10415,N_8601,N_8790);
or U10416 (N_10416,N_5611,N_9657);
and U10417 (N_10417,N_7499,N_5555);
xor U10418 (N_10418,N_5587,N_8864);
nor U10419 (N_10419,N_8017,N_8275);
nand U10420 (N_10420,N_8210,N_9648);
nand U10421 (N_10421,N_5784,N_5643);
and U10422 (N_10422,N_7219,N_7906);
nand U10423 (N_10423,N_9103,N_8668);
and U10424 (N_10424,N_5612,N_6241);
nand U10425 (N_10425,N_5967,N_7081);
and U10426 (N_10426,N_6343,N_6613);
nor U10427 (N_10427,N_5477,N_6422);
or U10428 (N_10428,N_9164,N_5175);
nand U10429 (N_10429,N_6261,N_8899);
xnor U10430 (N_10430,N_8020,N_6000);
nor U10431 (N_10431,N_5305,N_6601);
xnor U10432 (N_10432,N_5510,N_9589);
and U10433 (N_10433,N_5356,N_6490);
or U10434 (N_10434,N_7453,N_9246);
nand U10435 (N_10435,N_5844,N_7190);
and U10436 (N_10436,N_7736,N_5756);
nor U10437 (N_10437,N_5482,N_7774);
nand U10438 (N_10438,N_8329,N_9902);
or U10439 (N_10439,N_7789,N_6424);
nor U10440 (N_10440,N_8423,N_5413);
xor U10441 (N_10441,N_6996,N_5328);
or U10442 (N_10442,N_7251,N_6876);
nand U10443 (N_10443,N_9126,N_6814);
and U10444 (N_10444,N_5599,N_8457);
and U10445 (N_10445,N_6447,N_6240);
nand U10446 (N_10446,N_5450,N_8311);
or U10447 (N_10447,N_8030,N_8731);
and U10448 (N_10448,N_5837,N_8264);
nand U10449 (N_10449,N_9717,N_7379);
and U10450 (N_10450,N_8458,N_5307);
or U10451 (N_10451,N_6760,N_9054);
or U10452 (N_10452,N_5199,N_9687);
nor U10453 (N_10453,N_9265,N_7718);
and U10454 (N_10454,N_8571,N_7995);
nor U10455 (N_10455,N_6129,N_5104);
and U10456 (N_10456,N_9968,N_9593);
and U10457 (N_10457,N_6981,N_6065);
xnor U10458 (N_10458,N_5840,N_7725);
nand U10459 (N_10459,N_8934,N_5984);
nand U10460 (N_10460,N_7817,N_8744);
or U10461 (N_10461,N_7836,N_7268);
nand U10462 (N_10462,N_7285,N_7112);
and U10463 (N_10463,N_8723,N_9035);
nor U10464 (N_10464,N_6372,N_7878);
or U10465 (N_10465,N_8881,N_6862);
and U10466 (N_10466,N_9637,N_7447);
or U10467 (N_10467,N_5832,N_7426);
or U10468 (N_10468,N_7715,N_9107);
nor U10469 (N_10469,N_8026,N_7215);
and U10470 (N_10470,N_9195,N_5558);
or U10471 (N_10471,N_8959,N_8059);
nor U10472 (N_10472,N_8365,N_8248);
xor U10473 (N_10473,N_7562,N_9471);
nor U10474 (N_10474,N_6969,N_5275);
or U10475 (N_10475,N_8322,N_5429);
or U10476 (N_10476,N_8749,N_7682);
nor U10477 (N_10477,N_7570,N_8006);
and U10478 (N_10478,N_8257,N_7469);
nor U10479 (N_10479,N_7723,N_7484);
and U10480 (N_10480,N_5217,N_8699);
nor U10481 (N_10481,N_6194,N_5637);
or U10482 (N_10482,N_8331,N_9552);
nor U10483 (N_10483,N_5331,N_7020);
and U10484 (N_10484,N_7358,N_6548);
nand U10485 (N_10485,N_9191,N_9878);
and U10486 (N_10486,N_5909,N_5546);
nand U10487 (N_10487,N_6578,N_9938);
nor U10488 (N_10488,N_6659,N_8639);
or U10489 (N_10489,N_6937,N_5375);
and U10490 (N_10490,N_7246,N_7032);
and U10491 (N_10491,N_7490,N_6654);
nor U10492 (N_10492,N_9830,N_7068);
nand U10493 (N_10493,N_7764,N_7075);
nor U10494 (N_10494,N_5138,N_7320);
nor U10495 (N_10495,N_8812,N_7576);
nand U10496 (N_10496,N_9465,N_9385);
nor U10497 (N_10497,N_7380,N_8632);
nor U10498 (N_10498,N_9401,N_9505);
nor U10499 (N_10499,N_6482,N_7741);
nand U10500 (N_10500,N_9271,N_6824);
nor U10501 (N_10501,N_7962,N_5659);
or U10502 (N_10502,N_6454,N_5418);
nor U10503 (N_10503,N_6069,N_9557);
or U10504 (N_10504,N_6419,N_8390);
and U10505 (N_10505,N_5597,N_6472);
or U10506 (N_10506,N_6174,N_9454);
nor U10507 (N_10507,N_5026,N_5047);
or U10508 (N_10508,N_7471,N_7097);
nand U10509 (N_10509,N_8401,N_6765);
nor U10510 (N_10510,N_6219,N_5111);
or U10511 (N_10511,N_8393,N_6873);
or U10512 (N_10512,N_8936,N_7078);
nor U10513 (N_10513,N_5277,N_5859);
nor U10514 (N_10514,N_9546,N_5505);
nor U10515 (N_10515,N_8147,N_8760);
nor U10516 (N_10516,N_5399,N_9809);
nand U10517 (N_10517,N_7158,N_9614);
nor U10518 (N_10518,N_8814,N_5715);
and U10519 (N_10519,N_5369,N_9934);
and U10520 (N_10520,N_9018,N_8145);
and U10521 (N_10521,N_8134,N_7772);
or U10522 (N_10522,N_8404,N_6006);
and U10523 (N_10523,N_9732,N_7868);
or U10524 (N_10524,N_9821,N_7942);
or U10525 (N_10525,N_9100,N_7831);
nor U10526 (N_10526,N_5775,N_8559);
xnor U10527 (N_10527,N_7643,N_9734);
nor U10528 (N_10528,N_6445,N_9678);
nand U10529 (N_10529,N_8672,N_9751);
or U10530 (N_10530,N_5349,N_9738);
nand U10531 (N_10531,N_7847,N_5608);
nand U10532 (N_10532,N_6887,N_8675);
nor U10533 (N_10533,N_9024,N_5846);
nor U10534 (N_10534,N_9174,N_7381);
xor U10535 (N_10535,N_6572,N_6007);
nand U10536 (N_10536,N_7514,N_9257);
nand U10537 (N_10537,N_8898,N_9718);
nand U10538 (N_10538,N_9452,N_5425);
xnor U10539 (N_10539,N_9580,N_8761);
nand U10540 (N_10540,N_7492,N_8725);
nand U10541 (N_10541,N_5223,N_9262);
nor U10542 (N_10542,N_6243,N_8979);
or U10543 (N_10543,N_9707,N_9149);
xor U10544 (N_10544,N_8181,N_6003);
or U10545 (N_10545,N_9988,N_7345);
and U10546 (N_10546,N_9094,N_8166);
nand U10547 (N_10547,N_7808,N_8713);
or U10548 (N_10548,N_7573,N_8062);
or U10549 (N_10549,N_8285,N_9285);
and U10550 (N_10550,N_9607,N_5249);
and U10551 (N_10551,N_5431,N_7830);
nand U10552 (N_10552,N_7746,N_9372);
nor U10553 (N_10553,N_9795,N_6617);
or U10554 (N_10554,N_5168,N_9710);
or U10555 (N_10555,N_6605,N_5613);
nor U10556 (N_10556,N_6740,N_6667);
xnor U10557 (N_10557,N_6138,N_6941);
nand U10558 (N_10558,N_5971,N_5085);
nand U10559 (N_10559,N_7588,N_9771);
xnor U10560 (N_10560,N_9663,N_7589);
nor U10561 (N_10561,N_6954,N_5661);
or U10562 (N_10562,N_8597,N_8470);
or U10563 (N_10563,N_7065,N_6156);
and U10564 (N_10564,N_6736,N_7744);
or U10565 (N_10565,N_6476,N_7581);
or U10566 (N_10566,N_6992,N_8985);
nor U10567 (N_10567,N_7846,N_5417);
nand U10568 (N_10568,N_6257,N_7287);
and U10569 (N_10569,N_7066,N_5262);
nor U10570 (N_10570,N_8700,N_8415);
nand U10571 (N_10571,N_6475,N_9918);
nand U10572 (N_10572,N_9668,N_9625);
or U10573 (N_10573,N_6741,N_8905);
xor U10574 (N_10574,N_8443,N_6152);
and U10575 (N_10575,N_5790,N_6462);
nor U10576 (N_10576,N_7948,N_8610);
or U10577 (N_10577,N_7210,N_8506);
nand U10578 (N_10578,N_8364,N_7513);
or U10579 (N_10579,N_5144,N_5258);
or U10580 (N_10580,N_5292,N_8204);
nand U10581 (N_10581,N_9565,N_7984);
and U10582 (N_10582,N_7073,N_5156);
nor U10583 (N_10583,N_5459,N_9498);
nand U10584 (N_10584,N_9058,N_8271);
nor U10585 (N_10585,N_8290,N_8466);
or U10586 (N_10586,N_8845,N_7341);
or U10587 (N_10587,N_6793,N_8929);
nand U10588 (N_10588,N_7336,N_5806);
and U10589 (N_10589,N_5915,N_9055);
or U10590 (N_10590,N_7051,N_5830);
nand U10591 (N_10591,N_8092,N_7616);
nor U10592 (N_10592,N_7597,N_5706);
nand U10593 (N_10593,N_6116,N_5728);
nor U10594 (N_10594,N_7095,N_9086);
or U10595 (N_10595,N_8974,N_5528);
or U10596 (N_10596,N_7351,N_9158);
and U10597 (N_10597,N_8874,N_8488);
and U10598 (N_10598,N_9768,N_6831);
or U10599 (N_10599,N_8298,N_5215);
nand U10600 (N_10600,N_9782,N_8360);
and U10601 (N_10601,N_9117,N_6721);
nand U10602 (N_10602,N_8788,N_5496);
xnor U10603 (N_10603,N_7701,N_6945);
nor U10604 (N_10604,N_8560,N_8407);
xnor U10605 (N_10605,N_5938,N_6348);
xor U10606 (N_10606,N_6268,N_7024);
and U10607 (N_10607,N_6926,N_8392);
nor U10608 (N_10608,N_8001,N_8346);
or U10609 (N_10609,N_5019,N_8694);
nand U10610 (N_10610,N_7572,N_9560);
and U10611 (N_10611,N_9152,N_9336);
nor U10612 (N_10612,N_9233,N_9727);
xor U10613 (N_10613,N_9161,N_8408);
xnor U10614 (N_10614,N_6788,N_8077);
xnor U10615 (N_10615,N_7534,N_5725);
nand U10616 (N_10616,N_9227,N_7776);
and U10617 (N_10617,N_7709,N_7076);
or U10618 (N_10618,N_5035,N_5752);
nor U10619 (N_10619,N_6660,N_5449);
xor U10620 (N_10620,N_8523,N_6610);
nand U10621 (N_10621,N_7410,N_9096);
nor U10622 (N_10622,N_8151,N_6802);
or U10623 (N_10623,N_5293,N_9983);
nor U10624 (N_10624,N_8355,N_6565);
nand U10625 (N_10625,N_8465,N_5604);
nor U10626 (N_10626,N_8193,N_9672);
and U10627 (N_10627,N_8636,N_5434);
nor U10628 (N_10628,N_5716,N_8716);
nand U10629 (N_10629,N_9638,N_5540);
nand U10630 (N_10630,N_8332,N_7617);
or U10631 (N_10631,N_7237,N_8487);
and U10632 (N_10632,N_6267,N_7372);
xor U10633 (N_10633,N_6281,N_7023);
nand U10634 (N_10634,N_8094,N_9730);
or U10635 (N_10635,N_7197,N_9464);
nor U10636 (N_10636,N_7470,N_6078);
xor U10637 (N_10637,N_9512,N_9530);
and U10638 (N_10638,N_6413,N_7298);
nor U10639 (N_10639,N_5011,N_5004);
or U10640 (N_10640,N_8246,N_8207);
nand U10641 (N_10641,N_7648,N_5722);
xnor U10642 (N_10642,N_5861,N_7093);
and U10643 (N_10643,N_8645,N_7509);
nand U10644 (N_10644,N_8782,N_8093);
nor U10645 (N_10645,N_8611,N_7185);
xor U10646 (N_10646,N_7288,N_8046);
and U10647 (N_10647,N_5939,N_9633);
and U10648 (N_10648,N_5927,N_6918);
or U10649 (N_10649,N_5273,N_7234);
nand U10650 (N_10650,N_7644,N_9857);
nor U10651 (N_10651,N_7155,N_8316);
and U10652 (N_10652,N_5229,N_5314);
or U10653 (N_10653,N_6892,N_9507);
or U10654 (N_10654,N_6112,N_8425);
and U10655 (N_10655,N_7517,N_9645);
and U10656 (N_10656,N_5484,N_9240);
or U10657 (N_10657,N_6536,N_5831);
or U10658 (N_10658,N_9196,N_5116);
nand U10659 (N_10659,N_6872,N_7172);
nor U10660 (N_10660,N_7761,N_7915);
nor U10661 (N_10661,N_8155,N_5383);
or U10662 (N_10662,N_7924,N_8857);
nand U10663 (N_10663,N_9818,N_9208);
and U10664 (N_10664,N_6060,N_5714);
and U10665 (N_10665,N_6048,N_8833);
or U10666 (N_10666,N_5218,N_9931);
xor U10667 (N_10667,N_5276,N_9090);
nand U10668 (N_10668,N_9735,N_9222);
nand U10669 (N_10669,N_9508,N_6469);
nand U10670 (N_10670,N_6189,N_8241);
and U10671 (N_10671,N_5134,N_6592);
nor U10672 (N_10672,N_8615,N_6019);
or U10673 (N_10673,N_6836,N_6392);
xnor U10674 (N_10674,N_6155,N_9577);
or U10675 (N_10675,N_5698,N_9205);
and U10676 (N_10676,N_5290,N_7010);
nand U10677 (N_10677,N_5095,N_8803);
and U10678 (N_10678,N_9133,N_8674);
nor U10679 (N_10679,N_8750,N_5056);
nor U10680 (N_10680,N_5561,N_6916);
nor U10681 (N_10681,N_5836,N_7645);
or U10682 (N_10682,N_8778,N_6924);
nand U10683 (N_10683,N_9569,N_6265);
nor U10684 (N_10684,N_6537,N_5081);
nand U10685 (N_10685,N_8900,N_6618);
and U10686 (N_10686,N_8550,N_5077);
nand U10687 (N_10687,N_6213,N_7047);
xor U10688 (N_10688,N_8921,N_6978);
nor U10689 (N_10689,N_9750,N_8173);
nand U10690 (N_10690,N_7928,N_8963);
nor U10691 (N_10691,N_7564,N_7318);
xnor U10692 (N_10692,N_7793,N_6964);
nor U10693 (N_10693,N_9545,N_5207);
or U10694 (N_10694,N_7337,N_9820);
nand U10695 (N_10695,N_8964,N_9733);
and U10696 (N_10696,N_8174,N_7332);
or U10697 (N_10697,N_7894,N_6559);
nand U10698 (N_10698,N_9760,N_8324);
and U10699 (N_10699,N_8781,N_9017);
nor U10700 (N_10700,N_9712,N_6917);
nor U10701 (N_10701,N_9109,N_8442);
nand U10702 (N_10702,N_8066,N_9436);
or U10703 (N_10703,N_6523,N_8772);
nand U10704 (N_10704,N_7773,N_9615);
nor U10705 (N_10705,N_8098,N_9829);
or U10706 (N_10706,N_7944,N_8612);
nand U10707 (N_10707,N_9942,N_5498);
nand U10708 (N_10708,N_8274,N_5568);
or U10709 (N_10709,N_5464,N_6484);
or U10710 (N_10710,N_9012,N_5391);
nand U10711 (N_10711,N_8395,N_5569);
nor U10712 (N_10712,N_5000,N_7437);
and U10713 (N_10713,N_5744,N_6604);
nand U10714 (N_10714,N_6857,N_6646);
and U10715 (N_10715,N_9484,N_9404);
and U10716 (N_10716,N_8800,N_9324);
nor U10717 (N_10717,N_6540,N_7994);
nor U10718 (N_10718,N_5839,N_7578);
and U10719 (N_10719,N_8766,N_8820);
or U10720 (N_10720,N_5944,N_8621);
nand U10721 (N_10721,N_9929,N_5871);
and U10722 (N_10722,N_5733,N_7695);
xor U10723 (N_10723,N_5983,N_7850);
nand U10724 (N_10724,N_6608,N_7932);
and U10725 (N_10725,N_6983,N_5538);
and U10726 (N_10726,N_7114,N_6784);
xor U10727 (N_10727,N_7756,N_8698);
nor U10728 (N_10728,N_8097,N_6768);
or U10729 (N_10729,N_5119,N_9680);
nand U10730 (N_10730,N_6526,N_7079);
nor U10731 (N_10731,N_8130,N_8033);
xnor U10732 (N_10732,N_8811,N_7267);
and U10733 (N_10733,N_5601,N_5627);
or U10734 (N_10734,N_5542,N_7374);
xor U10735 (N_10735,N_9093,N_6772);
nor U10736 (N_10736,N_6446,N_6132);
nor U10737 (N_10737,N_5521,N_5379);
nor U10738 (N_10738,N_9690,N_7395);
nand U10739 (N_10739,N_7224,N_7865);
nand U10740 (N_10740,N_8448,N_9312);
nand U10741 (N_10741,N_9574,N_6516);
or U10742 (N_10742,N_7651,N_8967);
or U10743 (N_10743,N_6201,N_7324);
nand U10744 (N_10744,N_9801,N_8110);
nor U10745 (N_10745,N_8624,N_5550);
nor U10746 (N_10746,N_5016,N_5548);
nor U10747 (N_10747,N_7460,N_5885);
nor U10748 (N_10748,N_9365,N_8977);
and U10749 (N_10749,N_9778,N_5255);
nand U10750 (N_10750,N_8074,N_9159);
nand U10751 (N_10751,N_8453,N_6538);
nor U10752 (N_10752,N_8858,N_7028);
or U10753 (N_10753,N_8272,N_7936);
nand U10754 (N_10754,N_6403,N_6723);
or U10755 (N_10755,N_7151,N_9116);
nand U10756 (N_10756,N_9157,N_5188);
nand U10757 (N_10757,N_9214,N_8583);
nor U10758 (N_10758,N_8184,N_8478);
nor U10759 (N_10759,N_8031,N_8050);
or U10760 (N_10760,N_6769,N_9393);
and U10761 (N_10761,N_5536,N_7873);
and U10762 (N_10762,N_8536,N_5271);
nand U10763 (N_10763,N_7303,N_6703);
nor U10764 (N_10764,N_9316,N_9527);
xor U10765 (N_10765,N_9047,N_7226);
nor U10766 (N_10766,N_6318,N_8661);
xnor U10767 (N_10767,N_6600,N_5090);
nand U10768 (N_10768,N_9802,N_8543);
and U10769 (N_10769,N_7013,N_5039);
and U10770 (N_10770,N_8927,N_9068);
nand U10771 (N_10771,N_8182,N_7555);
xor U10772 (N_10772,N_7355,N_7031);
and U10773 (N_10773,N_9606,N_7502);
nand U10774 (N_10774,N_7300,N_8547);
xnor U10775 (N_10775,N_9224,N_7390);
or U10776 (N_10776,N_5455,N_7664);
and U10777 (N_10777,N_7991,N_5989);
nand U10778 (N_10778,N_9943,N_5074);
or U10779 (N_10779,N_5748,N_5947);
or U10780 (N_10780,N_7275,N_9039);
or U10781 (N_10781,N_6585,N_9345);
nor U10782 (N_10782,N_7388,N_6781);
nand U10783 (N_10783,N_5381,N_7851);
xor U10784 (N_10784,N_5233,N_7083);
nand U10785 (N_10785,N_5506,N_5930);
xnor U10786 (N_10786,N_9368,N_9876);
or U10787 (N_10787,N_7778,N_7790);
nand U10788 (N_10788,N_5393,N_7164);
and U10789 (N_10789,N_7347,N_7729);
nor U10790 (N_10790,N_7699,N_9449);
or U10791 (N_10791,N_6407,N_9141);
or U10792 (N_10792,N_9253,N_8616);
nor U10793 (N_10793,N_7805,N_8844);
xnor U10794 (N_10794,N_9714,N_7008);
nand U10795 (N_10795,N_5669,N_9390);
or U10796 (N_10796,N_7439,N_7156);
or U10797 (N_10797,N_9612,N_7811);
nor U10798 (N_10798,N_9188,N_5091);
or U10799 (N_10799,N_5878,N_7473);
or U10800 (N_10800,N_8460,N_9956);
and U10801 (N_10801,N_6596,N_5723);
and U10802 (N_10802,N_5432,N_9504);
and U10803 (N_10803,N_6704,N_9908);
xor U10804 (N_10804,N_7683,N_5059);
or U10805 (N_10805,N_6332,N_6730);
nor U10806 (N_10806,N_8512,N_5663);
or U10807 (N_10807,N_9941,N_6031);
and U10808 (N_10808,N_8711,N_9867);
nand U10809 (N_10809,N_5995,N_9831);
nand U10810 (N_10810,N_8370,N_5303);
xor U10811 (N_10811,N_6014,N_6642);
nand U10812 (N_10812,N_8468,N_5422);
nor U10813 (N_10813,N_8315,N_6122);
nand U10814 (N_10814,N_6047,N_7852);
nand U10815 (N_10815,N_6496,N_8497);
nand U10816 (N_10816,N_5642,N_7679);
nor U10817 (N_10817,N_8947,N_9814);
nor U10818 (N_10818,N_9074,N_8303);
nand U10819 (N_10819,N_6672,N_5312);
nand U10820 (N_10820,N_5771,N_6513);
nand U10821 (N_10821,N_7537,N_7833);
or U10822 (N_10822,N_9111,N_8254);
nor U10823 (N_10823,N_9330,N_6607);
nand U10824 (N_10824,N_6955,N_5849);
xor U10825 (N_10825,N_5672,N_7279);
nor U10826 (N_10826,N_7702,N_9515);
and U10827 (N_10827,N_9781,N_5322);
or U10828 (N_10828,N_8753,N_5140);
nor U10829 (N_10829,N_7304,N_6380);
or U10830 (N_10830,N_6220,N_9255);
or U10831 (N_10831,N_7521,N_8038);
and U10832 (N_10832,N_8709,N_9347);
nor U10833 (N_10833,N_6742,N_9700);
nand U10834 (N_10834,N_6074,N_7231);
nor U10835 (N_10835,N_8948,N_9922);
or U10836 (N_10836,N_7124,N_9491);
xnor U10837 (N_10837,N_9291,N_5980);
nor U10838 (N_10838,N_5084,N_9812);
or U10839 (N_10839,N_9720,N_5497);
nor U10840 (N_10840,N_5251,N_7740);
or U10841 (N_10841,N_9895,N_9270);
or U10842 (N_10842,N_6563,N_8325);
nand U10843 (N_10843,N_5605,N_8679);
or U10844 (N_10844,N_5284,N_8449);
or U10845 (N_10845,N_5105,N_6797);
nand U10846 (N_10846,N_6423,N_6022);
nor U10847 (N_10847,N_9112,N_9030);
or U10848 (N_10848,N_6154,N_7110);
nand U10849 (N_10849,N_8317,N_7387);
nand U10850 (N_10850,N_8920,N_5544);
or U10851 (N_10851,N_8111,N_8065);
xor U10852 (N_10852,N_9723,N_7263);
and U10853 (N_10853,N_9392,N_5018);
and U10854 (N_10854,N_5183,N_6505);
nand U10855 (N_10855,N_6166,N_7769);
or U10856 (N_10856,N_8510,N_6897);
or U10857 (N_10857,N_5804,N_9628);
nor U10858 (N_10858,N_8757,N_9211);
and U10859 (N_10859,N_7969,N_7412);
and U10860 (N_10860,N_6079,N_5171);
xnor U10861 (N_10861,N_8148,N_7474);
nor U10862 (N_10862,N_7925,N_7147);
and U10863 (N_10863,N_5692,N_6615);
nor U10864 (N_10864,N_6647,N_6968);
or U10865 (N_10865,N_7670,N_5596);
nor U10866 (N_10866,N_9900,N_8323);
nor U10867 (N_10867,N_6160,N_8153);
and U10868 (N_10868,N_7411,N_9509);
or U10869 (N_10869,N_6310,N_9272);
and U10870 (N_10870,N_5208,N_9072);
nor U10871 (N_10871,N_9827,N_6821);
nand U10872 (N_10872,N_9932,N_5582);
nor U10873 (N_10873,N_9796,N_8194);
nor U10874 (N_10874,N_7996,N_7964);
or U10875 (N_10875,N_6570,N_8867);
nor U10876 (N_10876,N_8319,N_7592);
or U10877 (N_10877,N_8133,N_6719);
nor U10878 (N_10878,N_8459,N_8909);
or U10879 (N_10879,N_6695,N_8524);
or U10880 (N_10880,N_6693,N_9850);
nor U10881 (N_10881,N_9382,N_7927);
nor U10882 (N_10882,N_7009,N_8337);
nor U10883 (N_10883,N_6854,N_7107);
nand U10884 (N_10884,N_8704,N_8034);
nand U10885 (N_10885,N_8873,N_8676);
nand U10886 (N_10886,N_9834,N_6689);
nand U10887 (N_10887,N_9194,N_9237);
and U10888 (N_10888,N_5791,N_6178);
and U10889 (N_10889,N_5149,N_9970);
nand U10890 (N_10890,N_9489,N_7771);
or U10891 (N_10891,N_9590,N_5818);
or U10892 (N_10892,N_7054,N_7354);
nor U10893 (N_10893,N_9666,N_7860);
xnor U10894 (N_10894,N_8013,N_5129);
xnor U10895 (N_10895,N_9424,N_8419);
nor U10896 (N_10896,N_7640,N_7429);
and U10897 (N_10897,N_6196,N_7911);
and U10898 (N_10898,N_9946,N_6478);
and U10899 (N_10899,N_8897,N_5245);
nand U10900 (N_10900,N_6364,N_6440);
nor U10901 (N_10901,N_8023,N_8265);
and U10902 (N_10902,N_9661,N_5825);
nand U10903 (N_10903,N_6436,N_9944);
and U10904 (N_10904,N_6801,N_5058);
xnor U10905 (N_10905,N_9252,N_6956);
xor U10906 (N_10906,N_6185,N_5598);
nor U10907 (N_10907,N_9911,N_6843);
nand U10908 (N_10908,N_5405,N_5281);
or U10909 (N_10909,N_5296,N_9554);
and U10910 (N_10910,N_6080,N_8195);
nand U10911 (N_10911,N_8693,N_6716);
or U10912 (N_10912,N_9682,N_7765);
nand U10913 (N_10913,N_8708,N_7828);
nand U10914 (N_10914,N_9219,N_9245);
nand U10915 (N_10915,N_7751,N_7937);
or U10916 (N_10916,N_8086,N_5563);
nor U10917 (N_10917,N_7005,N_7311);
nor U10918 (N_10918,N_5625,N_5153);
and U10919 (N_10919,N_5170,N_6810);
nor U10920 (N_10920,N_6853,N_8565);
nand U10921 (N_10921,N_5652,N_9568);
and U10922 (N_10922,N_7696,N_9306);
or U10923 (N_10923,N_9605,N_5732);
and U10924 (N_10924,N_8287,N_8328);
and U10925 (N_10925,N_8529,N_6808);
nand U10926 (N_10926,N_6562,N_9618);
or U10927 (N_10927,N_7971,N_9543);
nor U10928 (N_10928,N_9602,N_6755);
and U10929 (N_10929,N_8495,N_6370);
nand U10930 (N_10930,N_9215,N_5254);
nor U10931 (N_10931,N_8581,N_9474);
or U10932 (N_10932,N_8379,N_9516);
nor U10933 (N_10933,N_6840,N_7194);
and U10934 (N_10934,N_6161,N_7735);
nor U10935 (N_10935,N_9694,N_7804);
nand U10936 (N_10936,N_5200,N_9127);
nand U10937 (N_10937,N_6834,N_8618);
nor U10938 (N_10938,N_6054,N_6076);
nand U10939 (N_10939,N_9708,N_8886);
and U10940 (N_10940,N_8424,N_5221);
nor U10941 (N_10941,N_5718,N_7113);
nand U10942 (N_10942,N_8846,N_8775);
or U10943 (N_10943,N_7478,N_5677);
and U10944 (N_10944,N_9779,N_7444);
or U10945 (N_10945,N_7596,N_8891);
nor U10946 (N_10946,N_8486,N_7739);
or U10947 (N_10947,N_9667,N_7266);
or U10948 (N_10948,N_5709,N_9496);
nor U10949 (N_10949,N_5146,N_9566);
xnor U10950 (N_10950,N_8783,N_6297);
nand U10951 (N_10951,N_8593,N_5437);
or U10952 (N_10952,N_9559,N_7750);
and U10953 (N_10953,N_9351,N_5992);
nand U10954 (N_10954,N_5564,N_9179);
nand U10955 (N_10955,N_9428,N_8887);
xnor U10956 (N_10956,N_7861,N_8270);
or U10957 (N_10957,N_6457,N_8941);
and U10958 (N_10958,N_9451,N_5214);
or U10959 (N_10959,N_8984,N_7690);
and U10960 (N_10960,N_5154,N_5509);
and U10961 (N_10961,N_8982,N_9711);
nand U10962 (N_10962,N_6787,N_9979);
and U10963 (N_10963,N_5717,N_6771);
nand U10964 (N_10964,N_8859,N_8326);
and U10965 (N_10965,N_8171,N_8530);
nor U10966 (N_10966,N_6725,N_6170);
nand U10967 (N_10967,N_8777,N_9297);
nor U10968 (N_10968,N_5988,N_7077);
or U10969 (N_10969,N_8069,N_5746);
and U10970 (N_10970,N_8344,N_8667);
and U10971 (N_10971,N_9816,N_6990);
or U10972 (N_10972,N_9573,N_7734);
nand U10973 (N_10973,N_5688,N_8848);
and U10974 (N_10974,N_5583,N_8815);
nor U10975 (N_10975,N_8061,N_6641);
or U10976 (N_10976,N_8341,N_9765);
nand U10977 (N_10977,N_8998,N_9958);
nor U10978 (N_10978,N_5187,N_8135);
nor U10979 (N_10979,N_7981,N_6218);
nor U10980 (N_10980,N_6779,N_5474);
or U10981 (N_10981,N_6507,N_7328);
or U10982 (N_10982,N_8978,N_6165);
xor U10983 (N_10983,N_6751,N_6603);
nand U10984 (N_10984,N_7935,N_6295);
or U10985 (N_10985,N_5673,N_5935);
nor U10986 (N_10986,N_9473,N_5348);
and U10987 (N_10987,N_9113,N_7386);
and U10988 (N_10988,N_9409,N_7538);
or U10989 (N_10989,N_8002,N_8348);
or U10990 (N_10990,N_5350,N_7129);
nand U10991 (N_10991,N_9120,N_9810);
and U10992 (N_10992,N_5319,N_9425);
and U10993 (N_10993,N_7346,N_8568);
or U10994 (N_10994,N_8932,N_5853);
nor U10995 (N_10995,N_8793,N_7993);
or U10996 (N_10996,N_7405,N_7089);
or U10997 (N_10997,N_7949,N_8983);
nand U10998 (N_10998,N_5486,N_8343);
nor U10999 (N_10999,N_8735,N_9431);
nand U11000 (N_11000,N_8794,N_5893);
or U11001 (N_11001,N_6911,N_6743);
nor U11002 (N_11002,N_5368,N_7918);
nand U11003 (N_11003,N_6480,N_8206);
nor U11004 (N_11004,N_8312,N_7014);
or U11005 (N_11005,N_9808,N_8131);
and U11006 (N_11006,N_6418,N_8868);
nand U11007 (N_11007,N_9533,N_7653);
nand U11008 (N_11008,N_9608,N_5136);
and U11009 (N_11009,N_9702,N_6365);
nand U11010 (N_11010,N_8600,N_6571);
and U11011 (N_11011,N_6107,N_9901);
nor U11012 (N_11012,N_7978,N_8222);
nand U11013 (N_11013,N_5529,N_6325);
nor U11014 (N_11014,N_9319,N_5739);
nand U11015 (N_11015,N_6688,N_9177);
or U11016 (N_11016,N_9691,N_5633);
nor U11017 (N_11017,N_8156,N_7145);
xor U11018 (N_11018,N_8382,N_8714);
nor U11019 (N_11019,N_5236,N_9965);
nor U11020 (N_11020,N_7001,N_8253);
and U11021 (N_11021,N_5594,N_7329);
nor U11022 (N_11022,N_9769,N_5435);
nor U11023 (N_11023,N_5372,N_6387);
or U11024 (N_11024,N_5736,N_9362);
nand U11025 (N_11025,N_6302,N_7087);
nor U11026 (N_11026,N_8016,N_9388);
nor U11027 (N_11027,N_6953,N_8961);
or U11028 (N_11028,N_5457,N_9925);
nand U11029 (N_11029,N_7256,N_6588);
or U11030 (N_11030,N_7884,N_6101);
nand U11031 (N_11031,N_6627,N_8689);
nor U11032 (N_11032,N_7348,N_9933);
nand U11033 (N_11033,N_6256,N_6464);
nor U11034 (N_11034,N_8745,N_7100);
xnor U11035 (N_11035,N_9251,N_8350);
or U11036 (N_11036,N_7302,N_8862);
and U11037 (N_11037,N_8662,N_5332);
nor U11038 (N_11038,N_6567,N_6848);
and U11039 (N_11039,N_6262,N_9169);
and U11040 (N_11040,N_9384,N_7289);
nand U11041 (N_11041,N_5492,N_6830);
or U11042 (N_11042,N_7523,N_9293);
xor U11043 (N_11043,N_9888,N_6041);
nor U11044 (N_11044,N_5850,N_8545);
or U11045 (N_11045,N_7768,N_8970);
nor U11046 (N_11046,N_7316,N_9463);
nor U11047 (N_11047,N_8747,N_6002);
nor U11048 (N_11048,N_9304,N_8032);
and U11049 (N_11049,N_6369,N_7241);
nor U11050 (N_11050,N_9128,N_6204);
nand U11051 (N_11051,N_6244,N_9101);
or U11052 (N_11052,N_9402,N_5678);
and U11053 (N_11053,N_9879,N_7872);
or U11054 (N_11054,N_9521,N_5828);
nor U11055 (N_11055,N_8664,N_9079);
nand U11056 (N_11056,N_7914,N_9940);
nor U11057 (N_11057,N_6860,N_5315);
and U11058 (N_11058,N_9841,N_9482);
nand U11059 (N_11059,N_5889,N_7476);
or U11060 (N_11060,N_7586,N_5374);
nand U11061 (N_11061,N_9737,N_5458);
nor U11062 (N_11062,N_6865,N_5220);
nand U11063 (N_11063,N_8870,N_8214);
nor U11064 (N_11064,N_6734,N_8773);
and U11065 (N_11065,N_6648,N_7820);
nand U11066 (N_11066,N_6506,N_6109);
nand U11067 (N_11067,N_7638,N_7434);
or U11068 (N_11068,N_6502,N_6935);
and U11069 (N_11069,N_5345,N_9561);
nor U11070 (N_11070,N_5925,N_5924);
and U11071 (N_11071,N_8349,N_8690);
and U11072 (N_11072,N_5336,N_6467);
nor U11073 (N_11073,N_9974,N_6050);
nor U11074 (N_11074,N_8301,N_5428);
nand U11075 (N_11075,N_5648,N_7601);
or U11076 (N_11076,N_5093,N_8024);
nor U11077 (N_11077,N_5190,N_8876);
and U11078 (N_11078,N_6053,N_8678);
nand U11079 (N_11079,N_7657,N_8157);
xnor U11080 (N_11080,N_6748,N_9132);
or U11081 (N_11081,N_5195,N_9346);
or U11082 (N_11082,N_6396,N_9544);
nor U11083 (N_11083,N_7477,N_9380);
xnor U11084 (N_11084,N_6481,N_6130);
or U11085 (N_11085,N_8302,N_9020);
nor U11086 (N_11086,N_8394,N_7366);
and U11087 (N_11087,N_9411,N_8353);
nor U11088 (N_11088,N_9002,N_5342);
or U11089 (N_11089,N_9806,N_5592);
nor U11090 (N_11090,N_5657,N_8573);
and U11091 (N_11091,N_6349,N_9146);
nand U11092 (N_11092,N_5876,N_9904);
nor U11093 (N_11093,N_8957,N_6891);
or U11094 (N_11094,N_7985,N_9485);
nor U11095 (N_11095,N_9282,N_8368);
or U11096 (N_11096,N_5157,N_9483);
or U11097 (N_11097,N_6479,N_8446);
or U11098 (N_11098,N_5139,N_8626);
and U11099 (N_11099,N_6722,N_7966);
nor U11100 (N_11100,N_7812,N_6997);
or U11101 (N_11101,N_7823,N_6188);
nor U11102 (N_11102,N_7693,N_7264);
nand U11103 (N_11103,N_6867,N_7466);
and U11104 (N_11104,N_7126,N_7485);
nand U11105 (N_11105,N_5686,N_8221);
and U11106 (N_11106,N_7015,N_9462);
nor U11107 (N_11107,N_7152,N_8036);
nor U11108 (N_11108,N_8406,N_8885);
and U11109 (N_11109,N_5770,N_5339);
and U11110 (N_11110,N_8861,N_6527);
or U11111 (N_11111,N_5852,N_5330);
or U11112 (N_11112,N_9427,N_7641);
nor U11113 (N_11113,N_6382,N_8426);
or U11114 (N_11114,N_6238,N_9877);
or U11115 (N_11115,N_9740,N_8053);
nand U11116 (N_11116,N_9268,N_6034);
nor U11117 (N_11117,N_6546,N_8907);
or U11118 (N_11118,N_5580,N_7162);
nor U11119 (N_11119,N_6167,N_8617);
nor U11120 (N_11120,N_5031,N_6345);
xnor U11121 (N_11121,N_8280,N_8755);
or U11122 (N_11122,N_8089,N_8894);
nand U11123 (N_11123,N_7025,N_5423);
nor U11124 (N_11124,N_6217,N_7250);
and U11125 (N_11125,N_7067,N_5416);
and U11126 (N_11126,N_9187,N_5237);
nor U11127 (N_11127,N_5410,N_6385);
xor U11128 (N_11128,N_9061,N_7491);
and U11129 (N_11129,N_9450,N_7394);
and U11130 (N_11130,N_7552,N_9784);
nor U11131 (N_11131,N_7367,N_6312);
and U11132 (N_11132,N_8398,N_7002);
nand U11133 (N_11133,N_6874,N_7422);
xor U11134 (N_11134,N_7910,N_7642);
xor U11135 (N_11135,N_6299,N_5668);
or U11136 (N_11136,N_8429,N_6432);
nor U11137 (N_11137,N_8586,N_5803);
xnor U11138 (N_11138,N_8888,N_7239);
or U11139 (N_11139,N_8878,N_5167);
nand U11140 (N_11140,N_8041,N_6702);
xnor U11141 (N_11141,N_9585,N_8829);
nor U11142 (N_11142,N_9556,N_9288);
nand U11143 (N_11143,N_9963,N_6386);
or U11144 (N_11144,N_8233,N_9216);
nor U11145 (N_11145,N_9239,N_8717);
nor U11146 (N_11146,N_6282,N_8992);
and U11147 (N_11147,N_7607,N_5858);
or U11148 (N_11148,N_5570,N_6972);
nand U11149 (N_11149,N_6580,N_7312);
or U11150 (N_11150,N_5239,N_9745);
or U11151 (N_11151,N_5101,N_7837);
and U11152 (N_11152,N_7091,N_5445);
and U11153 (N_11153,N_6497,N_8011);
and U11154 (N_11154,N_6833,N_7088);
or U11155 (N_11155,N_6993,N_6542);
and U11156 (N_11156,N_8284,N_7122);
nand U11157 (N_11157,N_9596,N_5053);
nor U11158 (N_11158,N_7752,N_8129);
or U11159 (N_11159,N_8141,N_7986);
nand U11160 (N_11160,N_5738,N_7929);
or U11161 (N_11161,N_8336,N_9136);
and U11162 (N_11162,N_9889,N_6182);
xor U11163 (N_11163,N_5067,N_8576);
and U11164 (N_11164,N_7340,N_6141);
or U11165 (N_11165,N_6521,N_7189);
nand U11166 (N_11166,N_8541,N_9279);
xnor U11167 (N_11167,N_5388,N_6455);
and U11168 (N_11168,N_5517,N_9459);
and U11169 (N_11169,N_9281,N_8479);
or U11170 (N_11170,N_9444,N_6291);
and U11171 (N_11171,N_8825,N_6461);
and U11172 (N_11172,N_8939,N_6692);
or U11173 (N_11173,N_7628,N_5358);
or U11174 (N_11174,N_6021,N_7550);
and U11175 (N_11175,N_5130,N_7205);
nand U11176 (N_11176,N_5523,N_8276);
or U11177 (N_11177,N_8819,N_5976);
nand U11178 (N_11178,N_6566,N_7137);
or U11179 (N_11179,N_6171,N_7148);
or U11180 (N_11180,N_8473,N_9583);
nand U11181 (N_11181,N_7619,N_7232);
nor U11182 (N_11182,N_8451,N_6230);
or U11183 (N_11183,N_9598,N_9701);
and U11184 (N_11184,N_5078,N_6753);
or U11185 (N_11185,N_7048,N_9405);
xor U11186 (N_11186,N_9826,N_9000);
nand U11187 (N_11187,N_9310,N_6173);
nand U11188 (N_11188,N_8763,N_5380);
nand U11189 (N_11189,N_5588,N_8505);
and U11190 (N_11190,N_6491,N_6406);
and U11191 (N_11191,N_5038,N_8882);
and U11192 (N_11192,N_9332,N_9619);
nand U11193 (N_11193,N_7059,N_7717);
nand U11194 (N_11194,N_6274,N_9746);
xor U11195 (N_11195,N_6534,N_9775);
or U11196 (N_11196,N_6530,N_5419);
and U11197 (N_11197,N_5176,N_5833);
and U11198 (N_11198,N_6735,N_9518);
and U11199 (N_11199,N_8071,N_9824);
and U11200 (N_11200,N_7721,N_7663);
nand U11201 (N_11201,N_7743,N_6849);
nor U11202 (N_11202,N_8528,N_7382);
xnor U11203 (N_11203,N_9006,N_7807);
or U11204 (N_11204,N_7254,N_8083);
and U11205 (N_11205,N_5869,N_7946);
or U11206 (N_11206,N_8863,N_8737);
nand U11207 (N_11207,N_8692,N_9813);
nor U11208 (N_11208,N_6920,N_5392);
nor U11209 (N_11209,N_6144,N_5868);
nor U11210 (N_11210,N_5123,N_8989);
nor U11211 (N_11211,N_6625,N_8192);
nor U11212 (N_11212,N_6886,N_8304);
or U11213 (N_11213,N_8122,N_8269);
nand U11214 (N_11214,N_6713,N_5964);
or U11215 (N_11215,N_8786,N_7885);
nand U11216 (N_11216,N_5912,N_9910);
xor U11217 (N_11217,N_6754,N_9220);
nand U11218 (N_11218,N_9108,N_7397);
and U11219 (N_11219,N_5502,N_5042);
or U11220 (N_11220,N_8554,N_7481);
or U11221 (N_11221,N_7507,N_8039);
nor U11222 (N_11222,N_6314,N_9783);
or U11223 (N_11223,N_8591,N_9370);
xor U11224 (N_11224,N_7571,N_5905);
or U11225 (N_11225,N_8067,N_6086);
or U11226 (N_11226,N_8385,N_8366);
nand U11227 (N_11227,N_5634,N_9757);
and U11228 (N_11228,N_9134,N_9344);
nand U11229 (N_11229,N_5117,N_7487);
nor U11230 (N_11230,N_7108,N_8880);
nor U11231 (N_11231,N_9964,N_8313);
or U11232 (N_11232,N_9665,N_5182);
and U11233 (N_11233,N_6015,N_6895);
and U11234 (N_11234,N_6168,N_5649);
or U11235 (N_11235,N_5088,N_7809);
nand U11236 (N_11236,N_8125,N_7240);
nor U11237 (N_11237,N_6744,N_6717);
or U11238 (N_11238,N_8969,N_6181);
nand U11239 (N_11239,N_9349,N_9617);
xnor U11240 (N_11240,N_5800,N_6324);
and U11241 (N_11241,N_6621,N_9950);
nand U11242 (N_11242,N_5874,N_7819);
nand U11243 (N_11243,N_7281,N_5267);
xnor U11244 (N_11244,N_9644,N_6306);
and U11245 (N_11245,N_7099,N_8638);
and U11246 (N_11246,N_8872,N_5888);
and U11247 (N_11247,N_6919,N_8474);
or U11248 (N_11248,N_9926,N_8427);
or U11249 (N_11249,N_7647,N_6226);
nor U11250 (N_11250,N_5919,N_7615);
and U11251 (N_11251,N_6223,N_6207);
and U11252 (N_11252,N_7880,N_7204);
and U11253 (N_11253,N_9248,N_6435);
or U11254 (N_11254,N_7635,N_7214);
and U11255 (N_11255,N_7084,N_9228);
and U11256 (N_11256,N_8295,N_9975);
nand U11257 (N_11257,N_7245,N_9193);
nor U11258 (N_11258,N_9478,N_8677);
nand U11259 (N_11259,N_7191,N_9966);
nor U11260 (N_11260,N_6098,N_8256);
nand U11261 (N_11261,N_5922,N_8511);
nor U11262 (N_11262,N_6389,N_9276);
or U11263 (N_11263,N_7430,N_6018);
or U11264 (N_11264,N_6611,N_8734);
nor U11265 (N_11265,N_5647,N_7371);
nor U11266 (N_11266,N_5904,N_5986);
nor U11267 (N_11267,N_6984,N_7230);
nand U11268 (N_11268,N_5635,N_6489);
and U11269 (N_11269,N_8680,N_5860);
nor U11270 (N_11270,N_9453,N_7173);
or U11271 (N_11271,N_5742,N_8310);
nor U11272 (N_11272,N_5977,N_6950);
or U11273 (N_11273,N_7016,N_6063);
nand U11274 (N_11274,N_8113,N_6106);
nor U11275 (N_11275,N_5178,N_7621);
and U11276 (N_11276,N_5910,N_6817);
and U11277 (N_11277,N_9719,N_5628);
nor U11278 (N_11278,N_8480,N_6614);
nand U11279 (N_11279,N_7049,N_9600);
nor U11280 (N_11280,N_8288,N_5658);
and U11281 (N_11281,N_7940,N_6738);
or U11282 (N_11282,N_9121,N_5283);
xnor U11283 (N_11283,N_5631,N_6696);
or U11284 (N_11284,N_8801,N_8260);
nor U11285 (N_11285,N_6805,N_6708);
nand U11286 (N_11286,N_9014,N_8759);
nor U11287 (N_11287,N_8827,N_7501);
nor U11288 (N_11288,N_6947,N_6024);
or U11289 (N_11289,N_8656,N_8112);
and U11290 (N_11290,N_9558,N_9468);
or U11291 (N_11291,N_5240,N_8128);
nand U11292 (N_11292,N_5854,N_8993);
nor U11293 (N_11293,N_5999,N_5802);
or U11294 (N_11294,N_8926,N_8189);
or U11295 (N_11295,N_5953,N_7293);
and U11296 (N_11296,N_7448,N_7086);
and U11297 (N_11297,N_7308,N_8721);
nor U11298 (N_11298,N_7689,N_5670);
nand U11299 (N_11299,N_9156,N_5227);
and U11300 (N_11300,N_7174,N_6656);
and U11301 (N_11301,N_5033,N_8578);
or U11302 (N_11302,N_6408,N_8296);
nand U11303 (N_11303,N_5819,N_7999);
and U11304 (N_11304,N_6378,N_7676);
nand U11305 (N_11305,N_9416,N_7732);
nor U11306 (N_11306,N_8496,N_5654);
nand U11307 (N_11307,N_6500,N_5882);
nand U11308 (N_11308,N_5451,N_8048);
or U11309 (N_11309,N_7800,N_9865);
nor U11310 (N_11310,N_6118,N_6192);
xor U11311 (N_11311,N_8629,N_8525);
or U11312 (N_11312,N_5681,N_5886);
and U11313 (N_11313,N_7034,N_9803);
and U11314 (N_11314,N_7753,N_9327);
and U11315 (N_11315,N_6245,N_5745);
xnor U11316 (N_11316,N_7323,N_7666);
nor U11317 (N_11317,N_9994,N_6001);
and U11318 (N_11318,N_5377,N_6525);
nand U11319 (N_11319,N_7945,N_7121);
and U11320 (N_11320,N_8860,N_6899);
or U11321 (N_11321,N_8908,N_6745);
nand U11322 (N_11322,N_7391,N_7766);
nand U11323 (N_11323,N_8177,N_5552);
or U11324 (N_11324,N_6305,N_6404);
nand U11325 (N_11325,N_6068,N_5928);
nor U11326 (N_11326,N_9915,N_9679);
or U11327 (N_11327,N_5326,N_5511);
xnor U11328 (N_11328,N_5705,N_8910);
or U11329 (N_11329,N_9371,N_5798);
nand U11330 (N_11330,N_9616,N_9242);
and U11331 (N_11331,N_6541,N_5589);
and U11332 (N_11332,N_6100,N_5203);
nand U11333 (N_11333,N_8389,N_9399);
nand U11334 (N_11334,N_7813,N_9673);
or U11335 (N_11335,N_8613,N_7085);
nor U11336 (N_11336,N_9305,N_7671);
nand U11337 (N_11337,N_8666,N_5973);
and U11338 (N_11338,N_5280,N_7396);
nor U11339 (N_11339,N_9537,N_9104);
nand U11340 (N_11340,N_6083,N_5027);
nand U11341 (N_11341,N_9984,N_7102);
or U11342 (N_11342,N_8835,N_7848);
nand U11343 (N_11343,N_6514,N_5740);
nor U11344 (N_11344,N_7435,N_6838);
or U11345 (N_11345,N_8158,N_7594);
and U11346 (N_11346,N_5475,N_8383);
nand U11347 (N_11347,N_7142,N_6634);
and U11348 (N_11348,N_6234,N_6870);
xor U11349 (N_11349,N_7109,N_7103);
and U11350 (N_11350,N_5209,N_6589);
and U11351 (N_11351,N_5682,N_6638);
or U11352 (N_11352,N_8950,N_6685);
nor U11353 (N_11353,N_8121,N_9069);
and U11354 (N_11354,N_6421,N_7018);
and U11355 (N_11355,N_9125,N_8375);
and U11356 (N_11356,N_8623,N_9119);
nor U11357 (N_11357,N_9766,N_9234);
nand U11358 (N_11358,N_9264,N_6690);
nand U11359 (N_11359,N_7926,N_8585);
nor U11360 (N_11360,N_5554,N_8736);
and U11361 (N_11361,N_7443,N_7933);
or U11362 (N_11362,N_6444,N_7130);
or U11363 (N_11363,N_7988,N_6967);
and U11364 (N_11364,N_9328,N_6558);
nand U11365 (N_11365,N_5460,N_7892);
and U11366 (N_11366,N_9909,N_6184);
nand U11367 (N_11367,N_7806,N_8463);
and U11368 (N_11368,N_6251,N_8232);
or U11369 (N_11369,N_5263,N_8300);
and U11370 (N_11370,N_6674,N_7011);
nor U11371 (N_11371,N_5758,N_7620);
or U11372 (N_11372,N_6852,N_8822);
and U11373 (N_11373,N_7794,N_9280);
or U11374 (N_11374,N_7199,N_7533);
nor U11375 (N_11375,N_7686,N_8719);
and U11376 (N_11376,N_9990,N_8592);
and U11377 (N_11377,N_6142,N_7863);
nor U11378 (N_11378,N_6409,N_9258);
nand U11379 (N_11379,N_9073,N_6903);
or U11380 (N_11380,N_6148,N_6583);
xor U11381 (N_11381,N_8278,N_6092);
and U11382 (N_11382,N_6511,N_6115);
nand U11383 (N_11383,N_7692,N_6237);
nand U11384 (N_11384,N_5591,N_5164);
nand U11385 (N_11385,N_5902,N_6058);
nor U11386 (N_11386,N_8681,N_6495);
and U11387 (N_11387,N_5001,N_8144);
nand U11388 (N_11388,N_5269,N_6963);
or U11389 (N_11389,N_9705,N_6806);
or U11390 (N_11390,N_8080,N_8558);
and U11391 (N_11391,N_5707,N_7591);
or U11392 (N_11392,N_7418,N_5197);
nor U11393 (N_11393,N_6040,N_5030);
nand U11394 (N_11394,N_5335,N_7972);
and U11395 (N_11395,N_9455,N_7898);
and U11396 (N_11396,N_7135,N_8980);
nor U11397 (N_11397,N_6029,N_6652);
or U11398 (N_11398,N_6976,N_8420);
nand U11399 (N_11399,N_7306,N_9692);
nor U11400 (N_11400,N_7593,N_5115);
and U11401 (N_11401,N_6888,N_5807);
nor U11402 (N_11402,N_5767,N_8108);
nor U11403 (N_11403,N_7967,N_5089);
or U11404 (N_11404,N_8381,N_6096);
nand U11405 (N_11405,N_9883,N_7037);
and U11406 (N_11406,N_9338,N_8160);
nand U11407 (N_11407,N_5734,N_8954);
and U11408 (N_11408,N_8376,N_6880);
nor U11409 (N_11409,N_7104,N_6344);
nand U11410 (N_11410,N_8663,N_6008);
nor U11411 (N_11411,N_6233,N_7222);
nor U11412 (N_11412,N_6798,N_7516);
or U11413 (N_11413,N_9526,N_7646);
or U11414 (N_11414,N_8168,N_5145);
nand U11415 (N_11415,N_8682,N_7413);
and U11416 (N_11416,N_7203,N_9232);
or U11417 (N_11417,N_7198,N_5957);
nor U11418 (N_11418,N_6599,N_9716);
or U11419 (N_11419,N_8622,N_6221);
nor U11420 (N_11420,N_6539,N_7577);
or U11421 (N_11421,N_8060,N_8937);
and U11422 (N_11422,N_8770,N_7512);
nor U11423 (N_11423,N_6673,N_5918);
or U11424 (N_11424,N_6253,N_8203);
and U11425 (N_11425,N_6515,N_7598);
nor U11426 (N_11426,N_9015,N_7409);
and U11427 (N_11427,N_7229,N_9952);
xor U11428 (N_11428,N_9322,N_9948);
xnor U11429 (N_11429,N_6235,N_7442);
nand U11430 (N_11430,N_5367,N_8140);
and U11431 (N_11431,N_7697,N_8371);
and U11432 (N_11432,N_6264,N_7916);
or U11433 (N_11433,N_9181,N_7856);
and U11434 (N_11434,N_6653,N_5816);
xor U11435 (N_11435,N_5062,N_6037);
nor U11436 (N_11436,N_8489,N_8724);
nor U11437 (N_11437,N_9295,N_5159);
nor U11438 (N_11438,N_9130,N_6901);
nand U11439 (N_11439,N_7656,N_9930);
nor U11440 (N_11440,N_9314,N_5341);
nor U11441 (N_11441,N_5969,N_6576);
or U11442 (N_11442,N_7451,N_5690);
or U11443 (N_11443,N_8684,N_9997);
or U11444 (N_11444,N_8072,N_5414);
and U11445 (N_11445,N_7799,N_6508);
nand U11446 (N_11446,N_5205,N_9256);
nor U11447 (N_11447,N_9432,N_6139);
and U11448 (N_11448,N_9036,N_8695);
and U11449 (N_11449,N_5693,N_5862);
or U11450 (N_11450,N_6871,N_9320);
nor U11451 (N_11451,N_5879,N_8527);
and U11452 (N_11452,N_9099,N_8513);
and U11453 (N_11453,N_6355,N_5843);
xnor U11454 (N_11454,N_9755,N_9772);
nor U11455 (N_11455,N_7796,N_8481);
nand U11456 (N_11456,N_5160,N_6146);
nor U11457 (N_11457,N_8839,N_5013);
xor U11458 (N_11458,N_9277,N_8587);
nand U11459 (N_11459,N_7243,N_7886);
nor U11460 (N_11460,N_5845,N_7930);
nand U11461 (N_11461,N_9896,N_7338);
nor U11462 (N_11462,N_5265,N_9729);
and U11463 (N_11463,N_9868,N_6818);
and U11464 (N_11464,N_7139,N_9124);
and U11465 (N_11465,N_7810,N_9622);
or U11466 (N_11466,N_7269,N_7317);
nor U11467 (N_11467,N_8045,N_9378);
or U11468 (N_11468,N_6350,N_5948);
and U11469 (N_11469,N_8798,N_8439);
or U11470 (N_11470,N_6319,N_6661);
and U11471 (N_11471,N_7631,N_5212);
nand U11472 (N_11472,N_7599,N_6300);
nand U11473 (N_11473,N_9044,N_7069);
or U11474 (N_11474,N_6694,N_9611);
nor U11475 (N_11475,N_5810,N_8273);
nor U11476 (N_11476,N_7700,N_6017);
nand U11477 (N_11477,N_9949,N_8150);
xor U11478 (N_11478,N_6845,N_5378);
and U11479 (N_11479,N_6474,N_7976);
or U11480 (N_11480,N_8849,N_7667);
or U11481 (N_11481,N_5180,N_5711);
xor U11482 (N_11482,N_6183,N_5607);
and U11483 (N_11483,N_5586,N_9923);
or U11484 (N_11484,N_5534,N_5444);
nor U11485 (N_11485,N_7006,N_8037);
or U11486 (N_11486,N_9323,N_6084);
nor U11487 (N_11487,N_7310,N_5865);
nor U11488 (N_11488,N_5527,N_5792);
or U11489 (N_11489,N_8335,N_6637);
and U11490 (N_11490,N_9426,N_9996);
nand U11491 (N_11491,N_5500,N_7257);
xor U11492 (N_11492,N_8103,N_5851);
nor U11493 (N_11493,N_6236,N_6356);
nor U11494 (N_11494,N_6780,N_5581);
and U11495 (N_11495,N_7608,N_8178);
nand U11496 (N_11496,N_5436,N_7688);
nand U11497 (N_11497,N_7315,N_5616);
nor U11498 (N_11498,N_7244,N_7544);
or U11499 (N_11499,N_7463,N_5666);
nand U11500 (N_11500,N_5943,N_8359);
xnor U11501 (N_11501,N_6200,N_6487);
or U11502 (N_11502,N_9743,N_7934);
and U11503 (N_11503,N_6961,N_7622);
xor U11504 (N_11504,N_8519,N_9448);
and U11505 (N_11505,N_8132,N_5956);
or U11506 (N_11506,N_6224,N_8633);
nand U11507 (N_11507,N_7072,N_5206);
nand U11508 (N_11508,N_5440,N_9805);
or U11509 (N_11509,N_5193,N_7153);
nor U11510 (N_11510,N_5201,N_8691);
and U11511 (N_11511,N_9674,N_9415);
nor U11512 (N_11512,N_7452,N_6671);
and U11513 (N_11513,N_8614,N_5408);
or U11514 (N_11514,N_7111,N_8025);
and U11515 (N_11515,N_9460,N_7159);
and U11516 (N_11516,N_5043,N_6333);
or U11517 (N_11517,N_5244,N_5173);
nand U11518 (N_11518,N_8082,N_9579);
and U11519 (N_11519,N_6531,N_5856);
or U11520 (N_11520,N_6353,N_6651);
nand U11521 (N_11521,N_9871,N_7425);
and U11522 (N_11522,N_7681,N_8768);
xor U11523 (N_11523,N_6811,N_6352);
nor U11524 (N_11524,N_8960,N_5226);
nand U11525 (N_11525,N_8743,N_5503);
xnor U11526 (N_11526,N_7181,N_9836);
and U11527 (N_11527,N_7438,N_5072);
nand U11528 (N_11528,N_5041,N_7235);
nand U11529 (N_11529,N_9438,N_8119);
nand U11530 (N_11530,N_9192,N_5867);
or U11531 (N_11531,N_5768,N_6010);
and U11532 (N_11532,N_6287,N_6691);
xnor U11533 (N_11533,N_8236,N_7042);
nor U11534 (N_11534,N_5911,N_5787);
nand U11535 (N_11535,N_5667,N_9497);
and U11536 (N_11536,N_6270,N_5131);
nor U11537 (N_11537,N_5282,N_6728);
nor U11538 (N_11538,N_8990,N_5826);
or U11539 (N_11539,N_5366,N_9377);
nor U11540 (N_11540,N_6341,N_9212);
nor U11541 (N_11541,N_9284,N_7360);
and U11542 (N_11542,N_7206,N_7963);
or U11543 (N_11543,N_8598,N_5522);
nor U11544 (N_11544,N_9342,N_9981);
xor U11545 (N_11545,N_9442,N_9407);
xor U11546 (N_11546,N_7877,N_8607);
nand U11547 (N_11547,N_7465,N_7923);
nand U11548 (N_11548,N_9977,N_7503);
or U11549 (N_11549,N_8477,N_7870);
and U11550 (N_11550,N_8482,N_5184);
and U11551 (N_11551,N_9709,N_7595);
nand U11552 (N_11552,N_7952,N_9536);
and U11553 (N_11553,N_6752,N_7056);
or U11554 (N_11554,N_8856,N_7525);
and U11555 (N_11555,N_8218,N_9631);
nor U11556 (N_11556,N_6759,N_9993);
xor U11557 (N_11557,N_8070,N_6727);
nor U11558 (N_11558,N_6657,N_9364);
or U11559 (N_11559,N_9689,N_6414);
xnor U11560 (N_11560,N_9131,N_9951);
nor U11561 (N_11561,N_6930,N_6822);
or U11562 (N_11562,N_8619,N_9340);
and U11563 (N_11563,N_6113,N_9050);
xor U11564 (N_11564,N_7519,N_6518);
nor U11565 (N_11565,N_7272,N_6046);
nor U11566 (N_11566,N_7060,N_9263);
nor U11567 (N_11567,N_5256,N_6586);
nor U11568 (N_11568,N_9671,N_7705);
nor U11569 (N_11569,N_8830,N_6655);
nor U11570 (N_11570,N_9899,N_9754);
and U11571 (N_11571,N_6025,N_5238);
and U11572 (N_11572,N_6150,N_9649);
and U11573 (N_11573,N_7071,N_6456);
nor U11574 (N_11574,N_7357,N_9851);
and U11575 (N_11575,N_6027,N_6368);
or U11576 (N_11576,N_5998,N_7402);
and U11577 (N_11577,N_7909,N_7685);
xor U11578 (N_11578,N_5225,N_5516);
xor U11579 (N_11579,N_7557,N_6612);
and U11580 (N_11580,N_5761,N_9209);
and U11581 (N_11581,N_9761,N_6669);
and U11582 (N_11582,N_5447,N_7428);
and U11583 (N_11583,N_7033,N_7433);
nor U11584 (N_11584,N_6842,N_8242);
nor U11585 (N_11585,N_7843,N_6381);
nor U11586 (N_11586,N_7450,N_9503);
xnor U11587 (N_11587,N_7117,N_8883);
or U11588 (N_11588,N_8515,N_9275);
nand U11589 (N_11589,N_5150,N_8567);
nor U11590 (N_11590,N_6232,N_5884);
nor U11591 (N_11591,N_9791,N_6826);
nor U11592 (N_11592,N_8729,N_6553);
or U11593 (N_11593,N_6650,N_9728);
or U11594 (N_11594,N_7482,N_5926);
nor U11595 (N_11595,N_6816,N_6767);
nand U11596 (N_11596,N_7334,N_9620);
nand U11597 (N_11597,N_7131,N_7053);
and U11598 (N_11598,N_7195,N_7871);
and U11599 (N_11599,N_7043,N_7707);
nor U11600 (N_11600,N_7587,N_8447);
nand U11601 (N_11601,N_7610,N_5525);
nand U11602 (N_11602,N_6869,N_7154);
nor U11603 (N_11603,N_8170,N_6795);
nand U11604 (N_11604,N_9833,N_8104);
and U11605 (N_11605,N_9774,N_7177);
xnor U11606 (N_11606,N_7542,N_7286);
and U11607 (N_11607,N_5397,N_9924);
nor U11608 (N_11608,N_9706,N_6277);
or U11609 (N_11609,N_7781,N_5298);
or U11610 (N_11610,N_6923,N_7842);
nor U11611 (N_11611,N_8005,N_7760);
nor U11612 (N_11612,N_8973,N_7958);
nand U11613 (N_11613,N_8853,N_8655);
or U11614 (N_11614,N_8432,N_8250);
or U11615 (N_11615,N_6158,N_8521);
nor U11616 (N_11616,N_5934,N_9433);
nor U11617 (N_11617,N_8255,N_9021);
and U11618 (N_11618,N_9564,N_9178);
nand U11619 (N_11619,N_9309,N_8292);
and U11620 (N_11620,N_5143,N_8263);
nor U11621 (N_11621,N_6337,N_7401);
or U11622 (N_11622,N_5034,N_9917);
nor U11623 (N_11623,N_9998,N_8464);
xor U11624 (N_11624,N_9207,N_6959);
nand U11625 (N_11625,N_9301,N_8120);
and U11626 (N_11626,N_5406,N_5704);
nor U11627 (N_11627,N_9013,N_8802);
and U11628 (N_11628,N_8758,N_7896);
nor U11629 (N_11629,N_5036,N_5443);
and U11630 (N_11630,N_9844,N_6309);
nand U11631 (N_11631,N_7982,N_6134);
nor U11632 (N_11632,N_7161,N_8040);
nor U11633 (N_11633,N_7907,N_9885);
nand U11634 (N_11634,N_5764,N_6863);
xnor U11635 (N_11635,N_8238,N_7403);
or U11636 (N_11636,N_5501,N_6620);
xnor U11637 (N_11637,N_5407,N_7187);
nand U11638 (N_11638,N_5650,N_5972);
nand U11639 (N_11639,N_5308,N_5894);
nand U11640 (N_11640,N_8956,N_8421);
nor U11641 (N_11641,N_7992,N_6658);
nor U11642 (N_11642,N_6554,N_6072);
or U11643 (N_11643,N_5481,N_5864);
nand U11644 (N_11644,N_7649,N_9435);
nand U11645 (N_11645,N_7384,N_8896);
and U11646 (N_11646,N_7788,N_8767);
and U11647 (N_11647,N_6416,N_7361);
xor U11648 (N_11648,N_9759,N_8201);
or U11649 (N_11649,N_7508,N_9067);
and U11650 (N_11650,N_7859,N_8542);
nor U11651 (N_11651,N_6453,N_7691);
nor U11652 (N_11652,N_7180,N_5680);
or U11653 (N_11653,N_6715,N_9038);
nor U11654 (N_11654,N_6906,N_7165);
or U11655 (N_11655,N_9420,N_6943);
and U11656 (N_11656,N_8516,N_5632);
and U11657 (N_11657,N_7970,N_6316);
nor U11658 (N_11658,N_8076,N_5289);
nand U11659 (N_11659,N_8251,N_6151);
and U11660 (N_11660,N_5125,N_5102);
or U11661 (N_11661,N_9640,N_5390);
nor U11662 (N_11662,N_9241,N_5892);
and U11663 (N_11663,N_8012,N_6222);
nor U11664 (N_11664,N_8417,N_7824);
and U11665 (N_11665,N_5724,N_9972);
xor U11666 (N_11666,N_6762,N_9501);
or U11667 (N_11667,N_7613,N_7609);
and U11668 (N_11668,N_8309,N_7722);
nand U11669 (N_11669,N_8851,N_7951);
xor U11670 (N_11670,N_6208,N_7565);
or U11671 (N_11671,N_5021,N_7258);
nor U11672 (N_11672,N_7399,N_8237);
or U11673 (N_11673,N_8503,N_5524);
xor U11674 (N_11674,N_7791,N_7494);
or U11675 (N_11675,N_5092,N_8084);
or U11676 (N_11676,N_6439,N_6358);
and U11677 (N_11677,N_8938,N_9913);
or U11678 (N_11678,N_7343,N_5822);
xnor U11679 (N_11679,N_8277,N_9358);
or U11680 (N_11680,N_5545,N_8372);
and U11681 (N_11681,N_5373,N_8286);
or U11682 (N_11682,N_5219,N_5691);
nand U11683 (N_11683,N_5128,N_7777);
or U11684 (N_11684,N_5186,N_7954);
and U11685 (N_11685,N_5900,N_9893);
or U11686 (N_11686,N_5629,N_6889);
nor U11687 (N_11687,N_5241,N_6005);
nor U11688 (N_11688,N_7758,N_8928);
and U11689 (N_11689,N_9887,N_5729);
and U11690 (N_11690,N_8727,N_5518);
nand U11691 (N_11691,N_5834,N_6966);
or U11692 (N_11692,N_6331,N_5993);
nand U11693 (N_11693,N_6172,N_9089);
and U11694 (N_11694,N_6631,N_7629);
or U11695 (N_11695,N_5210,N_7567);
or U11696 (N_11696,N_6991,N_7747);
or U11697 (N_11697,N_6011,N_5291);
xnor U11698 (N_11698,N_5513,N_6544);
or U11699 (N_11699,N_6809,N_9166);
nand U11700 (N_11700,N_6433,N_9894);
nor U11701 (N_11701,N_8318,N_7980);
nand U11702 (N_11702,N_6026,N_6932);
and U11703 (N_11703,N_7864,N_6212);
or U11704 (N_11704,N_6707,N_6473);
or U11705 (N_11705,N_5537,N_8595);
nor U11706 (N_11706,N_9334,N_7524);
nand U11707 (N_11707,N_5675,N_5908);
and U11708 (N_11708,N_6761,N_8650);
or U11709 (N_11709,N_7349,N_8741);
or U11710 (N_11710,N_9266,N_6279);
nand U11711 (N_11711,N_7035,N_9553);
nor U11712 (N_11712,N_8388,N_5945);
nor U11713 (N_11713,N_8162,N_9927);
or U11714 (N_11714,N_6038,N_6739);
and U11715 (N_11715,N_6680,N_5794);
and U11716 (N_11716,N_8588,N_5786);
or U11717 (N_11717,N_5895,N_6304);
and U11718 (N_11718,N_6379,N_5547);
nor U11719 (N_11719,N_8995,N_8437);
and U11720 (N_11720,N_9456,N_6420);
nand U11721 (N_11721,N_7207,N_9875);
nand U11722 (N_11722,N_7090,N_7543);
or U11723 (N_11723,N_7314,N_7424);
or U11724 (N_11724,N_9576,N_9847);
and U11725 (N_11725,N_6425,N_5531);
or U11726 (N_11726,N_7036,N_5337);
and U11727 (N_11727,N_5820,N_5286);
or U11728 (N_11728,N_7192,N_6750);
or U11729 (N_11729,N_5370,N_6032);
nor U11730 (N_11730,N_6731,N_5921);
or U11731 (N_11731,N_7294,N_5473);
or U11732 (N_11732,N_6488,N_6030);
or U11733 (N_11733,N_9106,N_5466);
or U11734 (N_11734,N_8671,N_7662);
nand U11735 (N_11735,N_9898,N_6293);
nand U11736 (N_11736,N_9110,N_8604);
nand U11737 (N_11737,N_7282,N_7957);
and U11738 (N_11738,N_6448,N_6912);
or U11739 (N_11739,N_6545,N_8216);
nor U11740 (N_11740,N_7728,N_7479);
or U11741 (N_11741,N_6494,N_8015);
and U11742 (N_11742,N_9788,N_7866);
or U11743 (N_11743,N_7661,N_6517);
and U11744 (N_11744,N_9434,N_7271);
or U11745 (N_11745,N_5222,N_9542);
and U11746 (N_11746,N_7007,N_5765);
nand U11747 (N_11747,N_6133,N_6075);
xor U11748 (N_11748,N_9513,N_7835);
xor U11749 (N_11749,N_8152,N_5623);
and U11750 (N_11750,N_5779,N_6519);
nor U11751 (N_11751,N_5665,N_7912);
nand U11752 (N_11752,N_9506,N_9028);
and U11753 (N_11753,N_8653,N_8106);
or U11754 (N_11754,N_6214,N_5324);
xor U11755 (N_11755,N_9777,N_6820);
nor U11756 (N_11756,N_9722,N_7352);
and U11757 (N_11757,N_8363,N_6388);
nand U11758 (N_11758,N_9046,N_6164);
nand U11759 (N_11759,N_5610,N_5198);
nor U11760 (N_11760,N_9477,N_5424);
and U11761 (N_11761,N_9862,N_5703);
or U11762 (N_11762,N_6259,N_8476);
xor U11763 (N_11763,N_7639,N_6336);
nand U11764 (N_11764,N_5008,N_7105);
nor U11765 (N_11765,N_9855,N_5318);
nand U11766 (N_11766,N_7446,N_5270);
nand U11767 (N_11767,N_6778,N_6373);
and U11768 (N_11768,N_8752,N_6357);
nand U11769 (N_11769,N_9957,N_6790);
or U11770 (N_11770,N_9333,N_8940);
or U11771 (N_11771,N_8975,N_5264);
and U11772 (N_11772,N_6330,N_6376);
or U11773 (N_11773,N_7730,N_5557);
xor U11774 (N_11774,N_9523,N_9510);
nand U11775 (N_11775,N_9575,N_8687);
and U11776 (N_11776,N_6837,N_8579);
or U11777 (N_11777,N_9749,N_9092);
and U11778 (N_11778,N_8462,N_5441);
nor U11779 (N_11779,N_9023,N_9736);
or U11780 (N_11780,N_5044,N_8191);
nand U11781 (N_11781,N_7291,N_8779);
nor U11782 (N_11782,N_5404,N_8972);
xor U11783 (N_11783,N_5515,N_7975);
and U11784 (N_11784,N_9367,N_8685);
and U11785 (N_11785,N_9082,N_9481);
nor U11786 (N_11786,N_8965,N_9591);
and U11787 (N_11787,N_6153,N_5165);
nor U11788 (N_11788,N_7625,N_7895);
nor U11789 (N_11789,N_6902,N_6131);
or U11790 (N_11790,N_8185,N_7385);
or U11791 (N_11791,N_6121,N_9753);
and U11792 (N_11792,N_8919,N_8966);
nor U11793 (N_11793,N_6556,N_6683);
and U11794 (N_11794,N_5866,N_7536);
or U11795 (N_11795,N_9676,N_6198);
nand U11796 (N_11796,N_6678,N_5624);
and U11797 (N_11797,N_7166,N_8976);
or U11798 (N_11798,N_8627,N_8509);
xnor U11799 (N_11799,N_8696,N_6939);
and U11800 (N_11800,N_7326,N_9374);
or U11801 (N_11801,N_5361,N_8657);
nor U11802 (N_11802,N_5278,N_7449);
and U11803 (N_11803,N_5577,N_8357);
or U11804 (N_11804,N_8115,N_9361);
or U11805 (N_11805,N_6925,N_6632);
and U11806 (N_11806,N_8208,N_8918);
or U11807 (N_11807,N_8000,N_7527);
nand U11808 (N_11808,N_7378,N_8330);
nand U11809 (N_11809,N_6628,N_9859);
and U11810 (N_11810,N_9907,N_5483);
nor U11811 (N_11811,N_8922,N_7733);
and U11812 (N_11812,N_5107,N_7767);
xor U11813 (N_11813,N_8594,N_7938);
or U11814 (N_11814,N_8933,N_7742);
xnor U11815 (N_11815,N_6609,N_5958);
xor U11816 (N_11816,N_7674,N_5352);
nand U11817 (N_11817,N_9267,N_6315);
nor U11818 (N_11818,N_9203,N_5017);
nand U11819 (N_11819,N_8838,N_8483);
nand U11820 (N_11820,N_8686,N_9662);
nor U11821 (N_11821,N_5285,N_6340);
nand U11822 (N_11822,N_7441,N_6974);
or U11823 (N_11823,N_8126,N_6841);
nand U11824 (N_11824,N_8987,N_5737);
nand U11825 (N_11825,N_7261,N_9048);
xor U11826 (N_11826,N_8824,N_6049);
and U11827 (N_11827,N_6998,N_9199);
and U11828 (N_11828,N_6402,N_5456);
xor U11829 (N_11829,N_6549,N_9403);
nor U11830 (N_11830,N_6137,N_6108);
and U11831 (N_11831,N_6856,N_9165);
and U11832 (N_11832,N_6091,N_8107);
and U11833 (N_11833,N_7462,N_6061);
nand U11834 (N_11834,N_8434,N_8399);
xnor U11835 (N_11835,N_7046,N_7844);
nor U11836 (N_11836,N_5442,N_8220);
xnor U11837 (N_11837,N_6898,N_5747);
or U11838 (N_11838,N_7584,N_6770);
nor U11839 (N_11839,N_5253,N_5776);
or U11840 (N_11840,N_9832,N_6466);
nor U11841 (N_11841,N_6329,N_6813);
nand U11842 (N_11842,N_6328,N_8652);
nor U11843 (N_11843,N_7950,N_7253);
or U11844 (N_11844,N_8805,N_8179);
or U11845 (N_11845,N_5321,N_8526);
nor U11846 (N_11846,N_9200,N_7273);
nor U11847 (N_11847,N_5519,N_5780);
or U11848 (N_11848,N_8396,N_6951);
and U11849 (N_11849,N_8400,N_7284);
nand U11850 (N_11850,N_9066,N_8911);
and U11851 (N_11851,N_7115,N_9151);
nor U11852 (N_11852,N_6758,N_6229);
and U11853 (N_11853,N_5446,N_9081);
or U11854 (N_11854,N_8127,N_6004);
and U11855 (N_11855,N_9160,N_8553);
nor U11856 (N_11856,N_5565,N_7526);
or U11857 (N_11857,N_5532,N_7274);
nand U11858 (N_11858,N_8345,N_6686);
xnor U11859 (N_11859,N_5355,N_8913);
xnor U11860 (N_11860,N_7175,N_6307);
or U11861 (N_11861,N_9601,N_7801);
nand U11862 (N_11862,N_5462,N_7039);
and U11863 (N_11863,N_7236,N_7004);
and U11864 (N_11864,N_5754,N_9247);
nor U11865 (N_11865,N_5873,N_7897);
and U11866 (N_11866,N_9798,N_9959);
and U11867 (N_11867,N_9238,N_5694);
or U11868 (N_11868,N_7770,N_8769);
xor U11869 (N_11869,N_8748,N_8402);
nor U11870 (N_11870,N_7498,N_6909);
nand U11871 (N_11871,N_5213,N_5651);
and U11872 (N_11872,N_8548,N_7445);
or U11873 (N_11873,N_8834,N_7821);
nor U11874 (N_11874,N_9823,N_7227);
or U11875 (N_11875,N_6800,N_5719);
nand U11876 (N_11876,N_7605,N_6803);
or U11877 (N_11877,N_5817,N_6776);
xor U11878 (N_11878,N_7998,N_7956);
or U11879 (N_11879,N_8705,N_6904);
xor U11880 (N_11880,N_8079,N_6124);
and U11881 (N_11881,N_6028,N_5877);
nor U11882 (N_11882,N_8136,N_7973);
or U11883 (N_11883,N_5710,N_8430);
and U11884 (N_11884,N_9811,N_9848);
nor U11885 (N_11885,N_7472,N_6789);
or U11886 (N_11886,N_6400,N_8789);
nor U11887 (N_11887,N_9337,N_9476);
or U11888 (N_11888,N_5211,N_8435);
nor U11889 (N_11889,N_9630,N_9080);
nor U11890 (N_11890,N_6248,N_9037);
xor U11891 (N_11891,N_5796,N_9114);
nand U11892 (N_11892,N_6499,N_8268);
or U11893 (N_11893,N_8239,N_5683);
and U11894 (N_11894,N_5075,N_9785);
or U11895 (N_11895,N_6225,N_7333);
nand U11896 (N_11896,N_9326,N_6271);
nand U11897 (N_11897,N_8075,N_9311);
and U11898 (N_11898,N_7655,N_9685);
or U11899 (N_11899,N_7026,N_8828);
nand U11900 (N_11900,N_8566,N_5712);
or U11901 (N_11901,N_7913,N_6908);
or U11902 (N_11902,N_9175,N_6791);
and U11903 (N_11903,N_5471,N_5316);
nand U11904 (N_11904,N_5359,N_8994);
nand U11905 (N_11905,N_8889,N_8333);
xor U11906 (N_11906,N_5313,N_6438);
nand U11907 (N_11907,N_5559,N_8063);
or U11908 (N_11908,N_9664,N_5985);
xor U11909 (N_11909,N_7082,N_8414);
nor U11910 (N_11910,N_8142,N_5881);
nand U11911 (N_11911,N_9586,N_9115);
nor U11912 (N_11912,N_9870,N_8912);
and U11913 (N_11913,N_7080,N_6093);
nand U11914 (N_11914,N_9487,N_9076);
nand U11915 (N_11915,N_6035,N_5252);
nand U11916 (N_11916,N_9520,N_7182);
and U11917 (N_11917,N_6228,N_9525);
or U11918 (N_11918,N_5046,N_7055);
nor U11919 (N_11919,N_9721,N_7238);
nor U11920 (N_11920,N_5560,N_7050);
nand U11921 (N_11921,N_5622,N_6195);
and U11922 (N_11922,N_7212,N_9139);
and U11923 (N_11923,N_7600,N_7052);
or U11924 (N_11924,N_9226,N_5054);
and U11925 (N_11925,N_8532,N_5609);
or U11926 (N_11926,N_8234,N_8514);
nor U11927 (N_11927,N_5923,N_8307);
and U11928 (N_11928,N_6231,N_7582);
nand U11929 (N_11929,N_6555,N_6394);
nand U11930 (N_11930,N_6573,N_8450);
or U11931 (N_11931,N_9376,N_7431);
nand U11932 (N_11932,N_5961,N_5950);
xor U11933 (N_11933,N_7098,N_6442);
or U11934 (N_11934,N_8742,N_5835);
nor U11935 (N_11935,N_8259,N_7217);
or U11936 (N_11936,N_7558,N_7074);
nand U11937 (N_11937,N_5619,N_6190);
nor U11938 (N_11938,N_5099,N_7903);
or U11939 (N_11939,N_9283,N_7712);
xnor U11940 (N_11940,N_6584,N_6864);
and U11941 (N_11941,N_9842,N_6679);
or U11942 (N_11942,N_9514,N_9864);
or U11943 (N_11943,N_9592,N_6210);
or U11944 (N_11944,N_8154,N_6468);
or U11945 (N_11945,N_6829,N_5329);
nor U11946 (N_11946,N_7862,N_9817);
or U11947 (N_11947,N_5382,N_5660);
xor U11948 (N_11948,N_9863,N_6145);
nor U11949 (N_11949,N_6191,N_7188);
nand U11950 (N_11950,N_9223,N_5185);
and U11951 (N_11951,N_9713,N_7276);
nand U11952 (N_11952,N_5801,N_5360);
or U11953 (N_11953,N_5494,N_5068);
nor U11954 (N_11954,N_9541,N_7044);
and U11955 (N_11955,N_6252,N_8916);
or U11956 (N_11956,N_6825,N_5487);
xor U11957 (N_11957,N_6979,N_6710);
xor U11958 (N_11958,N_6339,N_9960);
nand U11959 (N_11959,N_8673,N_7365);
nor U11960 (N_11960,N_6272,N_6835);
or U11961 (N_11961,N_9387,N_5294);
nand U11962 (N_11962,N_8291,N_6095);
nand U11963 (N_11963,N_8028,N_7356);
nor U11964 (N_11964,N_7917,N_6247);
and U11965 (N_11965,N_6263,N_7136);
and U11966 (N_11966,N_8866,N_7660);
nand U11967 (N_11967,N_8646,N_7149);
nand U11968 (N_11968,N_6326,N_8852);
and U11969 (N_11969,N_9494,N_8266);
nand U11970 (N_11970,N_5645,N_5387);
and U11971 (N_11971,N_6844,N_8871);
or U11972 (N_11972,N_6510,N_5618);
nor U11973 (N_11973,N_5137,N_5696);
xor U11974 (N_11974,N_9009,N_5896);
xor U11975 (N_11975,N_8042,N_5166);
nor U11976 (N_11976,N_7857,N_8109);
or U11977 (N_11977,N_6643,N_8895);
and U11978 (N_11978,N_6668,N_9945);
and U11979 (N_11979,N_5630,N_8018);
nor U11980 (N_11980,N_6988,N_8410);
nor U11981 (N_11981,N_9604,N_8997);
nand U11982 (N_11982,N_6346,N_9646);
or U11983 (N_11983,N_6361,N_7359);
nand U11984 (N_11984,N_5452,N_7710);
and U11985 (N_11985,N_5133,N_7003);
or U11986 (N_11986,N_5974,N_8262);
or U11987 (N_11987,N_6568,N_7561);
and U11988 (N_11988,N_8338,N_9548);
or U11989 (N_11989,N_8906,N_5094);
nor U11990 (N_11990,N_7720,N_6982);
nand U11991 (N_11991,N_7540,N_8258);
xor U11992 (N_11992,N_6052,N_6729);
nand U11993 (N_11993,N_5990,N_7138);
nor U11994 (N_11994,N_9567,N_5364);
or U11995 (N_11995,N_7989,N_7248);
nor U11996 (N_11996,N_8431,N_7724);
or U11997 (N_11997,N_8923,N_6952);
nand U11998 (N_11998,N_5327,N_9792);
and U11999 (N_11999,N_9059,N_5028);
nand U12000 (N_12000,N_6013,N_7575);
or U12001 (N_12001,N_6921,N_8596);
nor U12002 (N_12002,N_9040,N_6211);
or U12003 (N_12003,N_7144,N_8475);
nand U12004 (N_12004,N_8582,N_6929);
or U12005 (N_12005,N_9699,N_7375);
nand U12006 (N_12006,N_8556,N_8606);
nand U12007 (N_12007,N_8608,N_5636);
or U12008 (N_12008,N_9502,N_5177);
nor U12009 (N_12009,N_9695,N_6501);
nand U12010 (N_12010,N_9563,N_5231);
and U12011 (N_12011,N_9406,N_9085);
nand U12012 (N_12012,N_8212,N_7546);
and U12013 (N_12013,N_6180,N_9652);
nand U12014 (N_12014,N_8143,N_6452);
nor U12015 (N_12015,N_7901,N_6288);
nand U12016 (N_12016,N_9381,N_7179);
nand U12017 (N_12017,N_8293,N_5469);
nor U12018 (N_12018,N_5073,N_6907);
or U12019 (N_12019,N_9008,N_6186);
nand U12020 (N_12020,N_9318,N_9499);
and U12021 (N_12021,N_8433,N_5015);
and U12022 (N_12022,N_9903,N_5490);
and U12023 (N_12023,N_7295,N_5351);
or U12024 (N_12024,N_7440,N_7795);
nand U12025 (N_12025,N_8102,N_6973);
or U12026 (N_12026,N_5702,N_8299);
or U12027 (N_12027,N_7495,N_6763);
nor U12028 (N_12028,N_9445,N_7221);
and U12029 (N_12029,N_5721,N_6794);
nand U12030 (N_12030,N_7531,N_8223);
and U12031 (N_12031,N_5751,N_6020);
nand U12032 (N_12032,N_7160,N_6881);
and U12033 (N_12033,N_9129,N_7979);
xnor U12034 (N_12034,N_6377,N_9846);
or U12035 (N_12035,N_8669,N_8294);
nor U12036 (N_12036,N_9261,N_6677);
nor U12037 (N_12037,N_6111,N_9840);
nor U12038 (N_12038,N_7398,N_8391);
and U12039 (N_12039,N_8022,N_5783);
nand U12040 (N_12040,N_6938,N_7726);
or U12041 (N_12041,N_9767,N_5931);
xnor U12042 (N_12042,N_8369,N_5065);
or U12043 (N_12043,N_7313,N_7319);
and U12044 (N_12044,N_5857,N_9786);
and U12045 (N_12045,N_8029,N_7669);
or U12046 (N_12046,N_8551,N_8841);
or U12047 (N_12047,N_9300,N_9182);
nor U12048 (N_12048,N_7247,N_6147);
nand U12049 (N_12049,N_5162,N_7556);
or U12050 (N_12050,N_5420,N_6276);
or U12051 (N_12051,N_7259,N_7961);
and U12052 (N_12052,N_8561,N_8914);
nor U12053 (N_12053,N_6561,N_6395);
nand U12054 (N_12054,N_6023,N_5112);
nand U12055 (N_12055,N_9886,N_6936);
and U12056 (N_12056,N_7574,N_8739);
and U12057 (N_12057,N_7606,N_8412);
nand U12058 (N_12058,N_5795,N_7029);
xnor U12059 (N_12059,N_7213,N_9852);
nand U12060 (N_12060,N_6317,N_9461);
xnor U12061 (N_12061,N_7530,N_8282);
and U12062 (N_12062,N_5671,N_6557);
nor U12063 (N_12063,N_5365,N_7505);
nor U12064 (N_12064,N_9122,N_7731);
nor U12065 (N_12065,N_5304,N_5334);
nor U12066 (N_12066,N_5070,N_9986);
nor U12067 (N_12067,N_9095,N_8955);
xnor U12068 (N_12068,N_9353,N_7309);
xnor U12069 (N_12069,N_7997,N_9202);
and U12070 (N_12070,N_6960,N_8634);
or U12071 (N_12071,N_7000,N_7400);
and U12072 (N_12072,N_9007,N_9647);
nand U12073 (N_12073,N_5196,N_5799);
or U12074 (N_12074,N_5079,N_9539);
nor U12075 (N_12075,N_8925,N_5777);
nand U12076 (N_12076,N_7547,N_9430);
nor U12077 (N_12077,N_8726,N_6323);
nor U12078 (N_12078,N_7590,N_6980);
nor U12079 (N_12079,N_5113,N_5749);
and U12080 (N_12080,N_6942,N_7404);
and U12081 (N_12081,N_6756,N_8810);
or U12082 (N_12082,N_9773,N_7321);
xor U12083 (N_12083,N_5913,N_9955);
nor U12084 (N_12084,N_8058,N_6227);
and U12085 (N_12085,N_9869,N_9804);
and U12086 (N_12086,N_6427,N_7201);
nor U12087 (N_12087,N_5343,N_8637);
or U12088 (N_12088,N_8243,N_6764);
xor U12089 (N_12089,N_5040,N_7094);
or U12090 (N_12090,N_9016,N_9153);
or U12091 (N_12091,N_8073,N_7779);
nor U12092 (N_12092,N_6193,N_7327);
and U12093 (N_12093,N_6644,N_6591);
nand U12094 (N_12094,N_5003,N_8780);
nor U12095 (N_12095,N_6354,N_5805);
nand U12096 (N_12096,N_7780,N_6564);
and U12097 (N_12097,N_8986,N_8340);
nand U12098 (N_12098,N_8225,N_6206);
or U12099 (N_12099,N_8057,N_9697);
nand U12100 (N_12100,N_8441,N_6663);
or U12101 (N_12101,N_7045,N_9613);
xnor U12102 (N_12102,N_6081,N_6321);
or U12103 (N_12103,N_6630,N_8836);
and U12104 (N_12104,N_5347,N_9389);
nand U12105 (N_12105,N_9290,N_5593);
nand U12106 (N_12106,N_5118,N_9467);
or U12107 (N_12107,N_8235,N_8380);
and U12108 (N_12108,N_6649,N_9097);
and U12109 (N_12109,N_8279,N_5603);
nand U12110 (N_12110,N_7427,N_8943);
nand U12111 (N_12111,N_7832,N_6994);
and U12112 (N_12112,N_8165,N_5750);
and U12113 (N_12113,N_6587,N_8334);
nand U12114 (N_12114,N_7493,N_6492);
nand U12115 (N_12115,N_7559,N_5394);
and U12116 (N_12116,N_8339,N_9535);
xor U12117 (N_12117,N_8630,N_6313);
nand U12118 (N_12118,N_8843,N_7840);
and U12119 (N_12119,N_8397,N_8522);
xor U12120 (N_12120,N_8599,N_8796);
or U12121 (N_12121,N_5224,N_5389);
nand U12122 (N_12122,N_6509,N_7634);
nor U12123 (N_12123,N_8869,N_9480);
nand U12124 (N_12124,N_5489,N_7012);
nand U12125 (N_12125,N_6064,N_5951);
nand U12126 (N_12126,N_9249,N_7713);
xor U12127 (N_12127,N_7297,N_8806);
and U12128 (N_12128,N_8648,N_6493);
nor U12129 (N_12129,N_8791,N_5470);
nand U12130 (N_12130,N_6463,N_5409);
nand U12131 (N_12131,N_5639,N_5060);
nor U12132 (N_12132,N_7714,N_5620);
nand U12133 (N_12133,N_9348,N_6426);
nor U12134 (N_12134,N_8533,N_6073);
and U12135 (N_12135,N_8808,N_9843);
and U12136 (N_12136,N_9874,N_9770);
and U12137 (N_12137,N_7675,N_7974);
or U12138 (N_12138,N_5726,N_8226);
and U12139 (N_12139,N_6827,N_6597);
or U12140 (N_12140,N_8877,N_9396);
or U12141 (N_12141,N_7618,N_9980);
nand U12142 (N_12142,N_7612,N_9386);
and U12143 (N_12143,N_8409,N_6551);
and U12144 (N_12144,N_7305,N_8306);
or U12145 (N_12145,N_8520,N_5821);
nand U12146 (N_12146,N_7322,N_7585);
nor U12147 (N_12147,N_8228,N_6216);
nor U12148 (N_12148,N_7193,N_6839);
nand U12149 (N_12149,N_8445,N_6102);
nand U12150 (N_12150,N_6157,N_7364);
or U12151 (N_12151,N_6384,N_9511);
or U12152 (N_12152,N_8471,N_8452);
or U12153 (N_12153,N_6676,N_5838);
and U12154 (N_12154,N_8603,N_5757);
nand U12155 (N_12155,N_9296,N_5615);
nand U12156 (N_12156,N_9357,N_8944);
or U12157 (N_12157,N_6104,N_5333);
nor U12158 (N_12158,N_8552,N_8641);
or U12159 (N_12159,N_7853,N_7603);
nor U12160 (N_12160,N_5465,N_5842);
nor U12161 (N_12161,N_8117,N_7202);
nand U12162 (N_12162,N_7184,N_8159);
nand U12163 (N_12163,N_5962,N_9500);
or U12164 (N_12164,N_8176,N_7408);
nand U12165 (N_12165,N_5543,N_5266);
nor U12166 (N_12166,N_9423,N_5363);
xnor U12167 (N_12167,N_6957,N_8149);
or U12168 (N_12168,N_9493,N_6090);
nor U12169 (N_12169,N_7684,N_5491);
nor U12170 (N_12170,N_6582,N_6934);
or U12171 (N_12171,N_8493,N_5181);
nand U12172 (N_12172,N_5179,N_5963);
or U12173 (N_12173,N_6460,N_5760);
nor U12174 (N_12174,N_9354,N_8342);
or U12175 (N_12175,N_8137,N_5887);
or U12176 (N_12176,N_8953,N_7782);
and U12177 (N_12177,N_7548,N_6412);
and U12178 (N_12178,N_6127,N_9057);
xor U12179 (N_12179,N_6749,N_9429);
or U12180 (N_12180,N_5697,N_6292);
nand U12181 (N_12181,N_8917,N_7432);
nor U12182 (N_12182,N_7480,N_6401);
nand U12183 (N_12183,N_7058,N_5250);
or U12184 (N_12184,N_5400,N_6775);
xnor U12185 (N_12185,N_7875,N_8138);
nor U12186 (N_12186,N_9686,N_6298);
and U12187 (N_12187,N_7363,N_9634);
nand U12188 (N_12188,N_6914,N_6602);
nand U12189 (N_12189,N_6202,N_6119);
or U12190 (N_12190,N_6428,N_9581);
xor U12191 (N_12191,N_8697,N_5120);
or U12192 (N_12192,N_6606,N_9278);
or U12193 (N_12193,N_7904,N_8217);
nand U12194 (N_12194,N_7922,N_5901);
nor U12195 (N_12195,N_6486,N_8085);
and U12196 (N_12196,N_6056,N_9041);
nand U12197 (N_12197,N_7890,N_9610);
nor U12198 (N_12198,N_6593,N_6360);
nor U12199 (N_12199,N_9995,N_6532);
or U12200 (N_12200,N_6675,N_7458);
and U12201 (N_12201,N_7658,N_5789);
and U12202 (N_12202,N_6851,N_8635);
or U12203 (N_12203,N_6087,N_5300);
or U12204 (N_12204,N_5929,N_6720);
nor U12205 (N_12205,N_5124,N_6737);
or U12206 (N_12206,N_9379,N_9599);
or U12207 (N_12207,N_8799,N_8577);
and U12208 (N_12208,N_7757,N_9636);
nand U12209 (N_12209,N_6410,N_9422);
and U12210 (N_12210,N_9331,N_6458);
or U12211 (N_12211,N_5052,N_5656);
nor U12212 (N_12212,N_5396,N_9954);
nand U12213 (N_12213,N_8962,N_8101);
or U12214 (N_12214,N_5002,N_8904);
or U12215 (N_12215,N_9421,N_5076);
or U12216 (N_12216,N_9744,N_5576);
nand U12217 (N_12217,N_8411,N_7677);
or U12218 (N_12218,N_6732,N_5376);
nand U12219 (N_12219,N_8422,N_7539);
or U12220 (N_12220,N_5812,N_7881);
nor U12221 (N_12221,N_9171,N_6159);
or U12222 (N_12222,N_5023,N_5295);
nand U12223 (N_12223,N_9764,N_5979);
and U12224 (N_12224,N_9897,N_8892);
or U12225 (N_12225,N_8840,N_7208);
or U12226 (N_12226,N_7716,N_5997);
nand U12227 (N_12227,N_6905,N_9075);
and U12228 (N_12228,N_6640,N_6977);
nand U12229 (N_12229,N_7941,N_8405);
or U12230 (N_12230,N_9229,N_8631);
nor U12231 (N_12231,N_6260,N_6009);
nand U12232 (N_12232,N_6879,N_5763);
xnor U12233 (N_12233,N_9825,N_6933);
and U12234 (N_12234,N_7520,N_6434);
xor U12235 (N_12235,N_5192,N_6664);
and U12236 (N_12236,N_5730,N_9555);
nand U12237 (N_12237,N_7827,N_5897);
nor U12238 (N_12238,N_8902,N_5551);
nand U12239 (N_12239,N_6417,N_5247);
xnor U12240 (N_12240,N_9635,N_5261);
nor U12241 (N_12241,N_7335,N_9033);
and U12242 (N_12242,N_6684,N_6275);
and U12243 (N_12243,N_8100,N_7849);
or U12244 (N_12244,N_8227,N_8188);
and U12245 (N_12245,N_7632,N_8762);
xor U12246 (N_12246,N_6581,N_9880);
nand U12247 (N_12247,N_5426,N_6045);
and U12248 (N_12248,N_9308,N_7680);
or U12249 (N_12249,N_5906,N_8211);
nand U12250 (N_12250,N_6303,N_5870);
nor U12251 (N_12251,N_6971,N_5940);
or U12252 (N_12252,N_6120,N_9928);
or U12253 (N_12253,N_5114,N_5955);
or U12254 (N_12254,N_8052,N_7092);
nor U12255 (N_12255,N_9144,N_9294);
nor U12256 (N_12256,N_9562,N_8054);
or U12257 (N_12257,N_5813,N_8832);
nor U12258 (N_12258,N_9739,N_9921);
or U12259 (N_12259,N_9654,N_6085);
nor U12260 (N_12260,N_8710,N_9049);
nand U12261 (N_12261,N_6311,N_6894);
nand U12262 (N_12262,N_8454,N_8373);
and U12263 (N_12263,N_9703,N_6471);
and U12264 (N_12264,N_6629,N_6322);
or U12265 (N_12265,N_9077,N_7163);
or U12266 (N_12266,N_6443,N_9204);
and U12267 (N_12267,N_7841,N_7822);
and U12268 (N_12268,N_5829,N_5009);
nor U12269 (N_12269,N_8224,N_9441);
or U12270 (N_12270,N_8469,N_5100);
nand U12271 (N_12271,N_9693,N_7626);
xnor U12272 (N_12272,N_8283,N_6123);
or U12273 (N_12273,N_7038,N_5354);
nand U12274 (N_12274,N_8570,N_5933);
nor U12275 (N_12275,N_8055,N_8722);
nor U12276 (N_12276,N_6199,N_7140);
and U12277 (N_12277,N_9916,N_9027);
and U12278 (N_12278,N_5573,N_6965);
nor U12279 (N_12279,N_9531,N_5676);
nand U12280 (N_12280,N_7415,N_5049);
or U12281 (N_12281,N_5731,N_6451);
nand U12282 (N_12282,N_5403,N_7566);
nor U12283 (N_12283,N_8854,N_8494);
nor U12284 (N_12284,N_5163,N_6308);
and U12285 (N_12285,N_6016,N_7977);
or U12286 (N_12286,N_7545,N_8733);
or U12287 (N_12287,N_8087,N_5467);
and U12288 (N_12288,N_7889,N_7604);
nand U12289 (N_12289,N_8281,N_6915);
and U12290 (N_12290,N_7784,N_7839);
nand U12291 (N_12291,N_8518,N_8386);
nor U12292 (N_12292,N_7350,N_5684);
and U12293 (N_12293,N_6724,N_7489);
nor U12294 (N_12294,N_7580,N_5248);
nand U12295 (N_12295,N_6670,N_6363);
xor U12296 (N_12296,N_6390,N_6483);
and U12297 (N_12297,N_8198,N_9213);
or U12298 (N_12298,N_8563,N_5020);
and U12299 (N_12299,N_7488,N_9183);
xnor U12300 (N_12300,N_9780,N_7816);
nand U12301 (N_12301,N_8751,N_8764);
xnor U12302 (N_12302,N_8890,N_6796);
nand U12303 (N_12303,N_5048,N_9123);
xnor U12304 (N_12304,N_6334,N_8804);
nor U12305 (N_12305,N_6294,N_7529);
nor U12306 (N_12306,N_6249,N_5005);
nand U12307 (N_12307,N_9373,N_9355);
and U12308 (N_12308,N_5096,N_9383);
nand U12309 (N_12309,N_8215,N_7200);
nand U12310 (N_12310,N_7955,N_8163);
nand U12311 (N_12311,N_6359,N_5438);
or U12312 (N_12312,N_9641,N_8924);
and U12313 (N_12313,N_7672,N_8771);
nand U12314 (N_12314,N_8792,N_9418);
nand U12315 (N_12315,N_8549,N_6622);
nand U12316 (N_12316,N_7704,N_8186);
nand U12317 (N_12317,N_5533,N_8351);
nor U12318 (N_12318,N_7650,N_9447);
nand U12319 (N_12319,N_9681,N_7826);
and U12320 (N_12320,N_6828,N_9912);
or U12321 (N_12321,N_7249,N_6254);
and U12322 (N_12322,N_8491,N_6893);
xnor U12323 (N_12323,N_8205,N_6785);
nor U12324 (N_12324,N_7652,N_5127);
nor U12325 (N_12325,N_8305,N_9350);
nand U12326 (N_12326,N_7568,N_9655);
or U12327 (N_12327,N_9105,N_5109);
or U12328 (N_12328,N_9623,N_9307);
and U12329 (N_12329,N_8660,N_6070);
xor U12330 (N_12330,N_9914,N_8590);
or U12331 (N_12331,N_6535,N_9244);
nand U12332 (N_12332,N_8605,N_9475);
xor U12333 (N_12333,N_7953,N_8659);
and U12334 (N_12334,N_9704,N_5848);
and U12335 (N_12335,N_6528,N_5655);
nand U12336 (N_12336,N_5051,N_6055);
nand U12337 (N_12337,N_9025,N_9231);
nor U12338 (N_12338,N_8252,N_6397);
or U12339 (N_12339,N_6367,N_5753);
nand U12340 (N_12340,N_8484,N_5638);
and U12341 (N_12341,N_5317,N_8321);
and U12342 (N_12342,N_5759,N_9595);
and U12343 (N_12343,N_7123,N_7211);
or U12344 (N_12344,N_6718,N_8718);
nor U12345 (N_12345,N_5769,N_9045);
nor U12346 (N_12346,N_8981,N_9469);
or U12347 (N_12347,N_9147,N_8644);
and U12348 (N_12348,N_9065,N_9799);
nor U12349 (N_12349,N_5172,N_7062);
nor U12350 (N_12350,N_5299,N_6746);
or U12351 (N_12351,N_9953,N_7900);
or U12352 (N_12352,N_7627,N_9670);
and U12353 (N_12353,N_5272,N_8014);
nor U12354 (N_12354,N_8797,N_6042);
or U12355 (N_12355,N_9920,N_8358);
and U12356 (N_12356,N_9439,N_5942);
xnor U12357 (N_12357,N_7178,N_5727);
xor U12358 (N_12358,N_6900,N_8544);
nor U12359 (N_12359,N_7611,N_7419);
and U12360 (N_12360,N_9363,N_8436);
xor U12361 (N_12361,N_6773,N_8499);
nor U12362 (N_12362,N_5148,N_9142);
xnor U12363 (N_12363,N_5773,N_6503);
nand U12364 (N_12364,N_8502,N_9731);
or U12365 (N_12365,N_5384,N_8942);
nor U12366 (N_12366,N_5508,N_7706);
xnor U12367 (N_12367,N_7040,N_9143);
xnor U12368 (N_12368,N_5232,N_8485);
nand U12369 (N_12369,N_5297,N_8651);
nand U12370 (N_12370,N_9828,N_5595);
and U12371 (N_12371,N_7659,N_8949);
and U12372 (N_12372,N_8628,N_8199);
or U12373 (N_12373,N_9603,N_9168);
and U12374 (N_12374,N_6162,N_6699);
and U12375 (N_12375,N_8649,N_6351);
or U12376 (N_12376,N_9019,N_9594);
or U12377 (N_12377,N_5617,N_5713);
or U12378 (N_12378,N_9042,N_7496);
nand U12379 (N_12379,N_6855,N_7891);
nor U12380 (N_12380,N_6890,N_9572);
nand U12381 (N_12381,N_5937,N_5311);
or U12382 (N_12382,N_5778,N_7919);
xor U12383 (N_12383,N_7186,N_7468);
nand U12384 (N_12384,N_5037,N_5614);
nor U12385 (N_12385,N_8785,N_9839);
nor U12386 (N_12386,N_9391,N_7290);
or U12387 (N_12387,N_7301,N_9763);
and U12388 (N_12388,N_5132,N_8507);
xnor U12389 (N_12389,N_9748,N_5025);
nand U12390 (N_12390,N_5346,N_6949);
nor U12391 (N_12391,N_6465,N_9138);
and U12392 (N_12392,N_9794,N_6986);
nand U12393 (N_12393,N_7727,N_8183);
nor U12394 (N_12394,N_7748,N_8720);
nor U12395 (N_12395,N_7307,N_6105);
xor U12396 (N_12396,N_9741,N_7678);
or U12397 (N_12397,N_5708,N_6962);
nor U12398 (N_12398,N_7869,N_5883);
or U12399 (N_12399,N_5259,N_5152);
nand U12400 (N_12400,N_7921,N_6529);
nand U12401 (N_12401,N_6574,N_9005);
and U12402 (N_12402,N_7070,N_9184);
and U12403 (N_12403,N_9524,N_5147);
nand U12404 (N_12404,N_7845,N_6097);
nand U12405 (N_12405,N_9210,N_7905);
xor U12406 (N_12406,N_9971,N_5235);
nor U12407 (N_12407,N_6099,N_9375);
nand U12408 (N_12408,N_7908,N_9395);
xnor U12409 (N_12409,N_8575,N_6269);
or U12410 (N_12410,N_6128,N_6094);
nand U12411 (N_12411,N_7931,N_6175);
or U12412 (N_12412,N_8555,N_6524);
nor U12413 (N_12413,N_5875,N_6645);
nor U12414 (N_12414,N_7407,N_6036);
nor U12415 (N_12415,N_7421,N_8123);
xnor U12416 (N_12416,N_6594,N_6242);
nor U12417 (N_12417,N_5553,N_5083);
nand U12418 (N_12418,N_6441,N_8467);
nor U12419 (N_12419,N_8589,N_5932);
nor U12420 (N_12420,N_9658,N_5029);
xnor U12421 (N_12421,N_5398,N_5824);
and U12422 (N_12422,N_8027,N_9235);
or U12423 (N_12423,N_5045,N_7106);
nand U12424 (N_12424,N_5827,N_5415);
and U12425 (N_12425,N_9725,N_8244);
xor U12426 (N_12426,N_7902,N_7983);
nand U12427 (N_12427,N_8935,N_8180);
and U12428 (N_12428,N_6431,N_8261);
nand U12429 (N_12429,N_7518,N_9639);
nor U12430 (N_12430,N_9522,N_7703);
or U12431 (N_12431,N_9800,N_8378);
nand U12432 (N_12432,N_5797,N_7563);
nor U12433 (N_12433,N_6342,N_8088);
nand U12434 (N_12434,N_6411,N_5268);
or U12435 (N_12435,N_9369,N_5785);
nand U12436 (N_12436,N_7119,N_9254);
or U12437 (N_12437,N_7141,N_7602);
and U12438 (N_12438,N_5427,N_8703);
nand U12439 (N_12439,N_7061,N_5050);
or U12440 (N_12440,N_6286,N_8584);
and U12441 (N_12441,N_9747,N_8219);
nor U12442 (N_12442,N_9186,N_5287);
or U12443 (N_12443,N_5057,N_7569);
or U12444 (N_12444,N_6819,N_9198);
nor U12445 (N_12445,N_5621,N_8387);
nor U12446 (N_12446,N_9359,N_6884);
nand U12447 (N_12447,N_8367,N_9084);
xnor U12448 (N_12448,N_9440,N_9022);
and U12449 (N_12449,N_7815,N_8999);
nand U12450 (N_12450,N_6163,N_9758);
nor U12451 (N_12451,N_9517,N_8915);
xnor U12452 (N_12452,N_6543,N_9078);
nand U12453 (N_12453,N_9935,N_6280);
nand U12454 (N_12454,N_9004,N_8816);
nor U12455 (N_12455,N_9053,N_7968);
nand U12456 (N_12456,N_6320,N_8051);
nor U12457 (N_12457,N_6636,N_8240);
nor U12458 (N_12458,N_5006,N_9408);
nor U12459 (N_12459,N_6697,N_9325);
and U12460 (N_12460,N_6140,N_7416);
nor U12461 (N_12461,N_7292,N_5097);
or U12462 (N_12462,N_6273,N_7579);
nor U12463 (N_12463,N_5811,N_9413);
nor U12464 (N_12464,N_9890,N_9835);
and U12465 (N_12465,N_9677,N_5110);
nor U12466 (N_12466,N_5507,N_8095);
nor U12467 (N_12467,N_6946,N_6203);
or U12468 (N_12468,N_6301,N_6711);
xnor U12469 (N_12469,N_6931,N_7373);
nand U12470 (N_12470,N_8498,N_9724);
and U12471 (N_12471,N_6437,N_9032);
or U12472 (N_12472,N_5158,N_5306);
or U12473 (N_12473,N_8230,N_9064);
xor U12474 (N_12474,N_8746,N_9742);
nor U12475 (N_12475,N_9273,N_5230);
or U12476 (N_12476,N_5007,N_6726);
or U12477 (N_12477,N_5646,N_9162);
and U12478 (N_12478,N_8609,N_7406);
and U12479 (N_12479,N_5814,N_7278);
nor U12480 (N_12480,N_5288,N_7803);
nand U12481 (N_12481,N_9597,N_7041);
or U12482 (N_12482,N_7457,N_6766);
xnor U12483 (N_12483,N_8971,N_9088);
nor U12484 (N_12484,N_5574,N_6285);
nor U12485 (N_12485,N_8403,N_9329);
and U12486 (N_12486,N_7504,N_8377);
or U12487 (N_12487,N_7280,N_5228);
and U12488 (N_12488,N_5579,N_9584);
nor U12489 (N_12489,N_5126,N_5320);
or U12490 (N_12490,N_9356,N_9274);
nand U12491 (N_12491,N_5512,N_9856);
and U12492 (N_12492,N_7754,N_9698);
or U12493 (N_12493,N_6985,N_8776);
nor U12494 (N_12494,N_9919,N_9011);
and U12495 (N_12495,N_6077,N_5499);
nor U12496 (N_12496,N_7614,N_9167);
nand U12497 (N_12497,N_5644,N_8968);
nand U12498 (N_12498,N_9190,N_7216);
nor U12499 (N_12499,N_9675,N_5847);
or U12500 (N_12500,N_6011,N_9327);
or U12501 (N_12501,N_6083,N_9131);
or U12502 (N_12502,N_8562,N_7835);
nand U12503 (N_12503,N_5209,N_6778);
and U12504 (N_12504,N_8842,N_7828);
or U12505 (N_12505,N_7556,N_5293);
or U12506 (N_12506,N_7416,N_6040);
nor U12507 (N_12507,N_7582,N_8786);
xor U12508 (N_12508,N_8188,N_7913);
nand U12509 (N_12509,N_5950,N_6166);
and U12510 (N_12510,N_8854,N_7286);
and U12511 (N_12511,N_7802,N_7523);
and U12512 (N_12512,N_5732,N_5988);
nand U12513 (N_12513,N_6975,N_5684);
and U12514 (N_12514,N_5607,N_5974);
or U12515 (N_12515,N_5166,N_5356);
xor U12516 (N_12516,N_6686,N_9231);
and U12517 (N_12517,N_6126,N_7615);
or U12518 (N_12518,N_6443,N_5183);
nand U12519 (N_12519,N_6812,N_9841);
and U12520 (N_12520,N_6163,N_9392);
and U12521 (N_12521,N_5271,N_7461);
xor U12522 (N_12522,N_8589,N_5386);
or U12523 (N_12523,N_9403,N_7674);
and U12524 (N_12524,N_7411,N_5191);
nor U12525 (N_12525,N_7462,N_7820);
nor U12526 (N_12526,N_7494,N_6904);
nand U12527 (N_12527,N_7644,N_6606);
and U12528 (N_12528,N_8456,N_6958);
xnor U12529 (N_12529,N_6514,N_6447);
nand U12530 (N_12530,N_7710,N_9755);
nand U12531 (N_12531,N_6205,N_8956);
or U12532 (N_12532,N_5781,N_5531);
or U12533 (N_12533,N_7381,N_9353);
and U12534 (N_12534,N_8966,N_9067);
or U12535 (N_12535,N_9649,N_7587);
nand U12536 (N_12536,N_5881,N_9819);
nand U12537 (N_12537,N_5905,N_9566);
nand U12538 (N_12538,N_5637,N_5153);
or U12539 (N_12539,N_8601,N_5550);
and U12540 (N_12540,N_7108,N_6799);
nand U12541 (N_12541,N_8624,N_7946);
xnor U12542 (N_12542,N_9977,N_8645);
nand U12543 (N_12543,N_9382,N_5389);
or U12544 (N_12544,N_6240,N_9997);
or U12545 (N_12545,N_5176,N_7060);
nor U12546 (N_12546,N_6445,N_7650);
and U12547 (N_12547,N_9262,N_5787);
or U12548 (N_12548,N_5084,N_7151);
and U12549 (N_12549,N_6832,N_7649);
nor U12550 (N_12550,N_8719,N_9740);
and U12551 (N_12551,N_5766,N_8878);
and U12552 (N_12552,N_9741,N_8314);
and U12553 (N_12553,N_7239,N_8243);
nand U12554 (N_12554,N_8185,N_5916);
or U12555 (N_12555,N_6529,N_9005);
nor U12556 (N_12556,N_9884,N_5481);
or U12557 (N_12557,N_5311,N_5535);
or U12558 (N_12558,N_7717,N_9242);
nand U12559 (N_12559,N_9221,N_8266);
nor U12560 (N_12560,N_7340,N_9195);
xor U12561 (N_12561,N_6708,N_8124);
and U12562 (N_12562,N_7374,N_7710);
and U12563 (N_12563,N_6515,N_6054);
or U12564 (N_12564,N_7823,N_5998);
nor U12565 (N_12565,N_7250,N_9867);
nand U12566 (N_12566,N_8520,N_5296);
or U12567 (N_12567,N_6076,N_6549);
or U12568 (N_12568,N_9445,N_9052);
or U12569 (N_12569,N_7995,N_9091);
or U12570 (N_12570,N_7895,N_6623);
or U12571 (N_12571,N_5459,N_7699);
and U12572 (N_12572,N_5631,N_8345);
and U12573 (N_12573,N_5316,N_7554);
and U12574 (N_12574,N_9596,N_5606);
nor U12575 (N_12575,N_8903,N_8005);
and U12576 (N_12576,N_8795,N_9358);
nand U12577 (N_12577,N_9937,N_6319);
nand U12578 (N_12578,N_7517,N_5606);
nand U12579 (N_12579,N_9597,N_9020);
or U12580 (N_12580,N_5732,N_7475);
nand U12581 (N_12581,N_6651,N_7886);
and U12582 (N_12582,N_8069,N_5223);
nor U12583 (N_12583,N_8705,N_6632);
or U12584 (N_12584,N_7965,N_6775);
nor U12585 (N_12585,N_7510,N_7558);
xnor U12586 (N_12586,N_5438,N_7680);
nor U12587 (N_12587,N_6944,N_5054);
xnor U12588 (N_12588,N_8684,N_7322);
or U12589 (N_12589,N_8154,N_7750);
nand U12590 (N_12590,N_6977,N_8629);
nor U12591 (N_12591,N_9775,N_7757);
and U12592 (N_12592,N_9002,N_5323);
or U12593 (N_12593,N_7857,N_6706);
nor U12594 (N_12594,N_6253,N_6975);
and U12595 (N_12595,N_5930,N_5794);
nor U12596 (N_12596,N_7349,N_7083);
nor U12597 (N_12597,N_9466,N_8604);
nand U12598 (N_12598,N_9526,N_5478);
nand U12599 (N_12599,N_8094,N_5808);
nand U12600 (N_12600,N_8330,N_7194);
nor U12601 (N_12601,N_5282,N_8087);
or U12602 (N_12602,N_7076,N_6902);
nand U12603 (N_12603,N_9747,N_8066);
and U12604 (N_12604,N_7361,N_5483);
xnor U12605 (N_12605,N_7576,N_8877);
or U12606 (N_12606,N_8383,N_7852);
or U12607 (N_12607,N_8772,N_5255);
nand U12608 (N_12608,N_7073,N_5761);
nand U12609 (N_12609,N_7021,N_9469);
nor U12610 (N_12610,N_5965,N_8267);
and U12611 (N_12611,N_6626,N_5765);
nor U12612 (N_12612,N_7076,N_5641);
and U12613 (N_12613,N_8489,N_7905);
or U12614 (N_12614,N_9268,N_5474);
nor U12615 (N_12615,N_7536,N_5137);
and U12616 (N_12616,N_9604,N_6845);
and U12617 (N_12617,N_5382,N_8252);
nand U12618 (N_12618,N_8883,N_6996);
or U12619 (N_12619,N_9308,N_6740);
and U12620 (N_12620,N_5233,N_5931);
nand U12621 (N_12621,N_8979,N_6547);
and U12622 (N_12622,N_6786,N_8852);
nand U12623 (N_12623,N_9919,N_8215);
or U12624 (N_12624,N_9752,N_6417);
nand U12625 (N_12625,N_8166,N_8052);
nor U12626 (N_12626,N_7531,N_7467);
nor U12627 (N_12627,N_8076,N_8122);
nor U12628 (N_12628,N_5439,N_7612);
and U12629 (N_12629,N_6248,N_9270);
nand U12630 (N_12630,N_8841,N_6023);
and U12631 (N_12631,N_8396,N_9036);
nor U12632 (N_12632,N_5005,N_9317);
or U12633 (N_12633,N_7492,N_6598);
nand U12634 (N_12634,N_7637,N_5967);
nor U12635 (N_12635,N_9686,N_8105);
or U12636 (N_12636,N_8064,N_8852);
or U12637 (N_12637,N_8843,N_7950);
nor U12638 (N_12638,N_8756,N_7756);
and U12639 (N_12639,N_5227,N_7821);
nor U12640 (N_12640,N_9525,N_8869);
and U12641 (N_12641,N_7491,N_6864);
or U12642 (N_12642,N_5245,N_5181);
nand U12643 (N_12643,N_8088,N_8677);
nor U12644 (N_12644,N_9344,N_7741);
nor U12645 (N_12645,N_8022,N_5654);
or U12646 (N_12646,N_7723,N_6691);
or U12647 (N_12647,N_9617,N_7627);
nand U12648 (N_12648,N_5044,N_5146);
nor U12649 (N_12649,N_8285,N_7834);
xor U12650 (N_12650,N_9434,N_5507);
or U12651 (N_12651,N_6669,N_7643);
or U12652 (N_12652,N_8521,N_7795);
nor U12653 (N_12653,N_5534,N_9131);
or U12654 (N_12654,N_8583,N_8490);
and U12655 (N_12655,N_7694,N_9753);
xnor U12656 (N_12656,N_9393,N_9397);
or U12657 (N_12657,N_7928,N_8416);
or U12658 (N_12658,N_5180,N_9390);
and U12659 (N_12659,N_9723,N_9253);
or U12660 (N_12660,N_6167,N_7917);
nand U12661 (N_12661,N_8932,N_8969);
nor U12662 (N_12662,N_8251,N_9715);
nand U12663 (N_12663,N_9673,N_7338);
and U12664 (N_12664,N_8258,N_8262);
nand U12665 (N_12665,N_6388,N_7670);
and U12666 (N_12666,N_6403,N_9995);
nand U12667 (N_12667,N_7134,N_5038);
nand U12668 (N_12668,N_7660,N_6462);
nand U12669 (N_12669,N_6283,N_7521);
and U12670 (N_12670,N_7551,N_9409);
or U12671 (N_12671,N_6288,N_5133);
and U12672 (N_12672,N_6572,N_9288);
or U12673 (N_12673,N_7726,N_7419);
and U12674 (N_12674,N_6241,N_7093);
nand U12675 (N_12675,N_6919,N_9925);
nand U12676 (N_12676,N_5020,N_6503);
or U12677 (N_12677,N_9016,N_5678);
or U12678 (N_12678,N_5615,N_5767);
or U12679 (N_12679,N_6471,N_9707);
or U12680 (N_12680,N_5690,N_8998);
and U12681 (N_12681,N_9368,N_6561);
nand U12682 (N_12682,N_7564,N_5308);
and U12683 (N_12683,N_6759,N_7503);
xnor U12684 (N_12684,N_5650,N_6677);
or U12685 (N_12685,N_9450,N_8398);
and U12686 (N_12686,N_8254,N_7737);
nor U12687 (N_12687,N_8248,N_9324);
and U12688 (N_12688,N_7425,N_9265);
or U12689 (N_12689,N_5744,N_6070);
nor U12690 (N_12690,N_6947,N_5908);
and U12691 (N_12691,N_6079,N_9562);
or U12692 (N_12692,N_6956,N_9746);
xnor U12693 (N_12693,N_5202,N_8848);
or U12694 (N_12694,N_5036,N_5990);
or U12695 (N_12695,N_7184,N_8356);
nand U12696 (N_12696,N_7653,N_9442);
xor U12697 (N_12697,N_6864,N_6044);
or U12698 (N_12698,N_8147,N_9947);
and U12699 (N_12699,N_9003,N_5585);
nand U12700 (N_12700,N_6977,N_8713);
and U12701 (N_12701,N_8640,N_5226);
nand U12702 (N_12702,N_9965,N_7586);
or U12703 (N_12703,N_7588,N_9049);
nor U12704 (N_12704,N_7716,N_6883);
nor U12705 (N_12705,N_7505,N_9155);
or U12706 (N_12706,N_7375,N_9073);
and U12707 (N_12707,N_8604,N_6554);
nand U12708 (N_12708,N_6525,N_8285);
nor U12709 (N_12709,N_8574,N_6621);
or U12710 (N_12710,N_5270,N_6644);
or U12711 (N_12711,N_9674,N_7665);
xor U12712 (N_12712,N_6323,N_7250);
xor U12713 (N_12713,N_8539,N_7996);
and U12714 (N_12714,N_8663,N_7837);
nor U12715 (N_12715,N_6001,N_9834);
nor U12716 (N_12716,N_7766,N_5050);
and U12717 (N_12717,N_6729,N_9953);
nor U12718 (N_12718,N_5388,N_7029);
or U12719 (N_12719,N_8114,N_9091);
and U12720 (N_12720,N_9546,N_9968);
nor U12721 (N_12721,N_8331,N_5981);
and U12722 (N_12722,N_9121,N_6472);
nor U12723 (N_12723,N_8386,N_5951);
nand U12724 (N_12724,N_5092,N_6952);
or U12725 (N_12725,N_9487,N_9951);
nor U12726 (N_12726,N_7489,N_8862);
xnor U12727 (N_12727,N_8959,N_5130);
xnor U12728 (N_12728,N_7015,N_5228);
or U12729 (N_12729,N_8461,N_8228);
and U12730 (N_12730,N_7213,N_7137);
or U12731 (N_12731,N_7683,N_8091);
and U12732 (N_12732,N_9404,N_7133);
xnor U12733 (N_12733,N_8309,N_6360);
xor U12734 (N_12734,N_9210,N_7133);
or U12735 (N_12735,N_7613,N_7132);
nand U12736 (N_12736,N_6136,N_6145);
or U12737 (N_12737,N_8385,N_7023);
and U12738 (N_12738,N_8394,N_5787);
xor U12739 (N_12739,N_6440,N_5344);
and U12740 (N_12740,N_7663,N_7603);
and U12741 (N_12741,N_9831,N_5063);
nand U12742 (N_12742,N_6538,N_9723);
or U12743 (N_12743,N_6638,N_9094);
nand U12744 (N_12744,N_9670,N_6963);
nor U12745 (N_12745,N_8353,N_8057);
nand U12746 (N_12746,N_7010,N_8707);
and U12747 (N_12747,N_8982,N_9475);
nand U12748 (N_12748,N_5223,N_7591);
and U12749 (N_12749,N_9952,N_9667);
and U12750 (N_12750,N_6013,N_6030);
nand U12751 (N_12751,N_8496,N_8548);
nand U12752 (N_12752,N_8634,N_5663);
nand U12753 (N_12753,N_7832,N_5829);
nand U12754 (N_12754,N_5415,N_8580);
or U12755 (N_12755,N_5741,N_6155);
xor U12756 (N_12756,N_9308,N_8212);
nor U12757 (N_12757,N_7919,N_6936);
nand U12758 (N_12758,N_7383,N_7159);
or U12759 (N_12759,N_7895,N_6229);
and U12760 (N_12760,N_8392,N_5612);
and U12761 (N_12761,N_5429,N_5281);
and U12762 (N_12762,N_6581,N_6877);
or U12763 (N_12763,N_8635,N_8764);
nand U12764 (N_12764,N_6284,N_8132);
and U12765 (N_12765,N_9825,N_5606);
or U12766 (N_12766,N_8097,N_9185);
or U12767 (N_12767,N_7736,N_8542);
or U12768 (N_12768,N_6895,N_9268);
nor U12769 (N_12769,N_6591,N_9834);
xnor U12770 (N_12770,N_7819,N_7260);
and U12771 (N_12771,N_6900,N_7591);
or U12772 (N_12772,N_7351,N_9607);
and U12773 (N_12773,N_8242,N_7213);
nor U12774 (N_12774,N_6650,N_5004);
nor U12775 (N_12775,N_9836,N_7191);
nor U12776 (N_12776,N_5826,N_7837);
or U12777 (N_12777,N_6292,N_7752);
xor U12778 (N_12778,N_7423,N_8042);
nand U12779 (N_12779,N_9957,N_8178);
nand U12780 (N_12780,N_9704,N_8251);
nand U12781 (N_12781,N_8730,N_5839);
and U12782 (N_12782,N_8775,N_7289);
nand U12783 (N_12783,N_9266,N_5756);
nand U12784 (N_12784,N_7721,N_6569);
nor U12785 (N_12785,N_7266,N_5257);
and U12786 (N_12786,N_7721,N_6395);
or U12787 (N_12787,N_9262,N_8412);
and U12788 (N_12788,N_7084,N_6072);
nand U12789 (N_12789,N_6304,N_9318);
or U12790 (N_12790,N_5656,N_7930);
nor U12791 (N_12791,N_6403,N_5214);
nor U12792 (N_12792,N_6576,N_5388);
nor U12793 (N_12793,N_5331,N_6133);
nor U12794 (N_12794,N_7504,N_6045);
or U12795 (N_12795,N_8534,N_9176);
or U12796 (N_12796,N_7856,N_9333);
nand U12797 (N_12797,N_7130,N_7279);
nor U12798 (N_12798,N_8790,N_8618);
nor U12799 (N_12799,N_5194,N_5493);
nor U12800 (N_12800,N_5397,N_5420);
nand U12801 (N_12801,N_9301,N_8180);
or U12802 (N_12802,N_5808,N_6168);
and U12803 (N_12803,N_7645,N_7632);
nor U12804 (N_12804,N_8850,N_9513);
and U12805 (N_12805,N_9752,N_9540);
xnor U12806 (N_12806,N_8010,N_5808);
and U12807 (N_12807,N_6266,N_6158);
or U12808 (N_12808,N_7004,N_9363);
and U12809 (N_12809,N_8945,N_7399);
nor U12810 (N_12810,N_7445,N_8390);
or U12811 (N_12811,N_9526,N_7127);
and U12812 (N_12812,N_7680,N_6953);
nand U12813 (N_12813,N_7697,N_9769);
nor U12814 (N_12814,N_5953,N_6406);
or U12815 (N_12815,N_9304,N_6129);
nand U12816 (N_12816,N_5093,N_8378);
nor U12817 (N_12817,N_7895,N_5756);
or U12818 (N_12818,N_5723,N_7520);
and U12819 (N_12819,N_9357,N_5804);
nand U12820 (N_12820,N_8665,N_7405);
nand U12821 (N_12821,N_9154,N_6427);
or U12822 (N_12822,N_8951,N_8477);
nor U12823 (N_12823,N_9693,N_9765);
or U12824 (N_12824,N_9399,N_5682);
xnor U12825 (N_12825,N_5556,N_7700);
nor U12826 (N_12826,N_6887,N_8267);
nand U12827 (N_12827,N_7136,N_8104);
or U12828 (N_12828,N_6515,N_6746);
and U12829 (N_12829,N_8614,N_5185);
nor U12830 (N_12830,N_6669,N_8583);
nand U12831 (N_12831,N_7072,N_5679);
or U12832 (N_12832,N_7983,N_9800);
nand U12833 (N_12833,N_7632,N_6132);
and U12834 (N_12834,N_8665,N_9624);
nor U12835 (N_12835,N_5381,N_9600);
or U12836 (N_12836,N_8757,N_5153);
or U12837 (N_12837,N_8110,N_7504);
and U12838 (N_12838,N_5556,N_6737);
and U12839 (N_12839,N_8977,N_5780);
nand U12840 (N_12840,N_5505,N_5935);
nor U12841 (N_12841,N_5188,N_7453);
or U12842 (N_12842,N_6036,N_8782);
and U12843 (N_12843,N_9650,N_6413);
xnor U12844 (N_12844,N_5488,N_5022);
and U12845 (N_12845,N_8190,N_6008);
nor U12846 (N_12846,N_7855,N_8766);
nor U12847 (N_12847,N_8331,N_8592);
or U12848 (N_12848,N_9905,N_6655);
or U12849 (N_12849,N_8738,N_7658);
nor U12850 (N_12850,N_5384,N_9661);
nand U12851 (N_12851,N_5572,N_5953);
or U12852 (N_12852,N_7647,N_5206);
nand U12853 (N_12853,N_9555,N_6343);
nor U12854 (N_12854,N_5592,N_6076);
nand U12855 (N_12855,N_7907,N_6137);
nor U12856 (N_12856,N_8934,N_7618);
nor U12857 (N_12857,N_7109,N_6269);
nor U12858 (N_12858,N_9512,N_6045);
nand U12859 (N_12859,N_5910,N_8859);
nor U12860 (N_12860,N_8931,N_6176);
nor U12861 (N_12861,N_8344,N_7123);
nor U12862 (N_12862,N_9896,N_9336);
and U12863 (N_12863,N_5512,N_8716);
nor U12864 (N_12864,N_8551,N_8740);
nor U12865 (N_12865,N_6842,N_5092);
or U12866 (N_12866,N_6176,N_8749);
nor U12867 (N_12867,N_5479,N_5463);
nor U12868 (N_12868,N_6569,N_5739);
nor U12869 (N_12869,N_9199,N_6769);
and U12870 (N_12870,N_5210,N_7831);
or U12871 (N_12871,N_8586,N_9227);
nand U12872 (N_12872,N_9875,N_8764);
or U12873 (N_12873,N_8212,N_5319);
xnor U12874 (N_12874,N_6132,N_9802);
nand U12875 (N_12875,N_8326,N_7791);
or U12876 (N_12876,N_9940,N_8243);
or U12877 (N_12877,N_9533,N_7683);
or U12878 (N_12878,N_7941,N_6223);
nor U12879 (N_12879,N_7324,N_5729);
or U12880 (N_12880,N_8981,N_5039);
or U12881 (N_12881,N_7232,N_7309);
and U12882 (N_12882,N_9690,N_8871);
nor U12883 (N_12883,N_9712,N_5620);
nand U12884 (N_12884,N_5618,N_6920);
or U12885 (N_12885,N_5174,N_5739);
nand U12886 (N_12886,N_9071,N_5327);
and U12887 (N_12887,N_8607,N_5245);
and U12888 (N_12888,N_7025,N_7274);
nand U12889 (N_12889,N_8924,N_9700);
nor U12890 (N_12890,N_6422,N_6191);
and U12891 (N_12891,N_8421,N_7655);
and U12892 (N_12892,N_7290,N_8823);
nand U12893 (N_12893,N_8473,N_7026);
nor U12894 (N_12894,N_6102,N_5493);
or U12895 (N_12895,N_6433,N_5540);
xor U12896 (N_12896,N_9892,N_8758);
and U12897 (N_12897,N_5452,N_8986);
nand U12898 (N_12898,N_7473,N_6087);
and U12899 (N_12899,N_6996,N_6008);
or U12900 (N_12900,N_8671,N_6950);
nand U12901 (N_12901,N_8349,N_6777);
nor U12902 (N_12902,N_5732,N_9348);
nand U12903 (N_12903,N_8700,N_8291);
and U12904 (N_12904,N_7192,N_8241);
and U12905 (N_12905,N_8986,N_5136);
and U12906 (N_12906,N_7301,N_9875);
nand U12907 (N_12907,N_8233,N_7333);
nor U12908 (N_12908,N_6511,N_9148);
and U12909 (N_12909,N_9011,N_8692);
nor U12910 (N_12910,N_5384,N_8133);
nor U12911 (N_12911,N_6852,N_9994);
nand U12912 (N_12912,N_6513,N_8063);
nand U12913 (N_12913,N_5574,N_9362);
nand U12914 (N_12914,N_5554,N_6202);
or U12915 (N_12915,N_8640,N_5221);
nand U12916 (N_12916,N_6848,N_5234);
nand U12917 (N_12917,N_6752,N_8156);
and U12918 (N_12918,N_5266,N_9125);
nand U12919 (N_12919,N_8904,N_9969);
nor U12920 (N_12920,N_6896,N_5984);
or U12921 (N_12921,N_9830,N_9986);
and U12922 (N_12922,N_6294,N_8952);
xnor U12923 (N_12923,N_8256,N_5555);
nor U12924 (N_12924,N_8759,N_6818);
nand U12925 (N_12925,N_5820,N_5979);
nand U12926 (N_12926,N_5943,N_7292);
nor U12927 (N_12927,N_7744,N_8300);
nand U12928 (N_12928,N_9361,N_6178);
or U12929 (N_12929,N_7119,N_9790);
nand U12930 (N_12930,N_5343,N_6584);
or U12931 (N_12931,N_5884,N_9599);
nor U12932 (N_12932,N_5551,N_8602);
nand U12933 (N_12933,N_8148,N_7939);
and U12934 (N_12934,N_8840,N_6154);
nand U12935 (N_12935,N_6703,N_5715);
nor U12936 (N_12936,N_9807,N_5513);
nand U12937 (N_12937,N_5906,N_5066);
nand U12938 (N_12938,N_9379,N_8672);
nor U12939 (N_12939,N_7663,N_7094);
nor U12940 (N_12940,N_6734,N_9870);
nand U12941 (N_12941,N_5932,N_8152);
nand U12942 (N_12942,N_8837,N_6876);
nand U12943 (N_12943,N_8144,N_7424);
and U12944 (N_12944,N_5353,N_7961);
nand U12945 (N_12945,N_9173,N_8248);
and U12946 (N_12946,N_5975,N_5881);
or U12947 (N_12947,N_8932,N_6135);
or U12948 (N_12948,N_6891,N_8964);
and U12949 (N_12949,N_9302,N_5281);
or U12950 (N_12950,N_8698,N_7495);
xor U12951 (N_12951,N_9172,N_5157);
or U12952 (N_12952,N_7195,N_8537);
nand U12953 (N_12953,N_7759,N_5320);
xor U12954 (N_12954,N_6168,N_8442);
and U12955 (N_12955,N_5346,N_5231);
or U12956 (N_12956,N_7232,N_6912);
nor U12957 (N_12957,N_7238,N_8339);
and U12958 (N_12958,N_7121,N_5837);
nor U12959 (N_12959,N_5544,N_9470);
or U12960 (N_12960,N_5193,N_6332);
nor U12961 (N_12961,N_5451,N_8550);
nand U12962 (N_12962,N_7034,N_9633);
or U12963 (N_12963,N_8502,N_9446);
nand U12964 (N_12964,N_5486,N_7280);
and U12965 (N_12965,N_9462,N_5303);
or U12966 (N_12966,N_6750,N_9887);
or U12967 (N_12967,N_8578,N_8723);
nand U12968 (N_12968,N_9164,N_7068);
nor U12969 (N_12969,N_8112,N_9950);
and U12970 (N_12970,N_8168,N_8312);
nor U12971 (N_12971,N_6846,N_8364);
or U12972 (N_12972,N_5454,N_9094);
or U12973 (N_12973,N_5779,N_7078);
nand U12974 (N_12974,N_9547,N_6319);
or U12975 (N_12975,N_6767,N_9127);
and U12976 (N_12976,N_9402,N_6774);
nand U12977 (N_12977,N_7887,N_6385);
and U12978 (N_12978,N_8868,N_7744);
and U12979 (N_12979,N_5819,N_5137);
nor U12980 (N_12980,N_8610,N_9557);
xor U12981 (N_12981,N_9747,N_8834);
nand U12982 (N_12982,N_6267,N_8471);
nor U12983 (N_12983,N_7033,N_6908);
nand U12984 (N_12984,N_5263,N_6856);
or U12985 (N_12985,N_9036,N_5582);
or U12986 (N_12986,N_8224,N_5821);
nor U12987 (N_12987,N_6559,N_9628);
and U12988 (N_12988,N_8435,N_9841);
or U12989 (N_12989,N_8337,N_8341);
or U12990 (N_12990,N_8824,N_6321);
nor U12991 (N_12991,N_5960,N_7669);
and U12992 (N_12992,N_6457,N_7511);
or U12993 (N_12993,N_9941,N_8587);
nand U12994 (N_12994,N_7327,N_6774);
nor U12995 (N_12995,N_8231,N_6202);
nand U12996 (N_12996,N_9100,N_8837);
and U12997 (N_12997,N_5108,N_9173);
nor U12998 (N_12998,N_8446,N_9683);
or U12999 (N_12999,N_6631,N_6941);
or U13000 (N_13000,N_8712,N_7789);
nand U13001 (N_13001,N_9219,N_9896);
and U13002 (N_13002,N_8412,N_9217);
or U13003 (N_13003,N_5758,N_6096);
nor U13004 (N_13004,N_6897,N_7742);
or U13005 (N_13005,N_6526,N_9715);
nor U13006 (N_13006,N_7843,N_6331);
or U13007 (N_13007,N_8623,N_6861);
and U13008 (N_13008,N_5609,N_9465);
xor U13009 (N_13009,N_8488,N_9249);
or U13010 (N_13010,N_6800,N_7393);
xor U13011 (N_13011,N_8535,N_7443);
or U13012 (N_13012,N_8400,N_5067);
nand U13013 (N_13013,N_6094,N_5306);
or U13014 (N_13014,N_7550,N_8523);
nand U13015 (N_13015,N_8527,N_8841);
or U13016 (N_13016,N_8213,N_6072);
or U13017 (N_13017,N_9146,N_5258);
nand U13018 (N_13018,N_9408,N_9946);
nand U13019 (N_13019,N_5726,N_7601);
and U13020 (N_13020,N_8869,N_6039);
or U13021 (N_13021,N_6301,N_8117);
or U13022 (N_13022,N_6956,N_9925);
nor U13023 (N_13023,N_5862,N_6450);
and U13024 (N_13024,N_9211,N_8487);
or U13025 (N_13025,N_8231,N_6184);
or U13026 (N_13026,N_6663,N_6740);
nand U13027 (N_13027,N_5557,N_6172);
and U13028 (N_13028,N_7920,N_5758);
or U13029 (N_13029,N_6022,N_6308);
and U13030 (N_13030,N_7622,N_8046);
nor U13031 (N_13031,N_5875,N_6120);
and U13032 (N_13032,N_5934,N_6797);
and U13033 (N_13033,N_5674,N_8241);
or U13034 (N_13034,N_9749,N_8547);
and U13035 (N_13035,N_9419,N_8392);
nand U13036 (N_13036,N_9685,N_8285);
or U13037 (N_13037,N_6490,N_6447);
xnor U13038 (N_13038,N_9446,N_6690);
or U13039 (N_13039,N_8929,N_7534);
or U13040 (N_13040,N_9711,N_9128);
nor U13041 (N_13041,N_6845,N_8725);
and U13042 (N_13042,N_6962,N_7638);
nor U13043 (N_13043,N_8223,N_8998);
or U13044 (N_13044,N_5375,N_7179);
nor U13045 (N_13045,N_8228,N_8098);
xnor U13046 (N_13046,N_8699,N_9023);
nand U13047 (N_13047,N_5865,N_6488);
nor U13048 (N_13048,N_7894,N_8673);
or U13049 (N_13049,N_6662,N_7088);
or U13050 (N_13050,N_6267,N_6622);
and U13051 (N_13051,N_8376,N_8727);
and U13052 (N_13052,N_5538,N_9194);
nor U13053 (N_13053,N_6375,N_6558);
nor U13054 (N_13054,N_8815,N_7081);
and U13055 (N_13055,N_8949,N_6655);
or U13056 (N_13056,N_6963,N_9015);
and U13057 (N_13057,N_5089,N_5461);
and U13058 (N_13058,N_7025,N_6350);
nand U13059 (N_13059,N_7957,N_7762);
nand U13060 (N_13060,N_5131,N_7890);
xor U13061 (N_13061,N_9928,N_6728);
or U13062 (N_13062,N_9556,N_7261);
and U13063 (N_13063,N_5518,N_7942);
nor U13064 (N_13064,N_8941,N_5898);
nor U13065 (N_13065,N_5962,N_9252);
and U13066 (N_13066,N_5262,N_6902);
nor U13067 (N_13067,N_6269,N_6795);
nor U13068 (N_13068,N_6287,N_8478);
nand U13069 (N_13069,N_9892,N_5382);
and U13070 (N_13070,N_5928,N_7291);
and U13071 (N_13071,N_9267,N_5131);
xor U13072 (N_13072,N_6596,N_5706);
nand U13073 (N_13073,N_5052,N_7762);
or U13074 (N_13074,N_8967,N_7027);
and U13075 (N_13075,N_9318,N_9849);
and U13076 (N_13076,N_6975,N_8749);
and U13077 (N_13077,N_7632,N_9283);
or U13078 (N_13078,N_7925,N_7155);
nand U13079 (N_13079,N_5412,N_8041);
nand U13080 (N_13080,N_9178,N_7151);
nor U13081 (N_13081,N_7815,N_6511);
nor U13082 (N_13082,N_7355,N_7813);
and U13083 (N_13083,N_9126,N_7864);
nand U13084 (N_13084,N_9733,N_6783);
nand U13085 (N_13085,N_6284,N_7888);
or U13086 (N_13086,N_8184,N_8129);
nor U13087 (N_13087,N_6661,N_8795);
and U13088 (N_13088,N_7991,N_6320);
or U13089 (N_13089,N_6901,N_9748);
and U13090 (N_13090,N_7723,N_6299);
nor U13091 (N_13091,N_7804,N_5672);
xnor U13092 (N_13092,N_6188,N_6993);
nor U13093 (N_13093,N_6684,N_7105);
nor U13094 (N_13094,N_5184,N_7526);
nand U13095 (N_13095,N_9505,N_5297);
or U13096 (N_13096,N_7213,N_7420);
nor U13097 (N_13097,N_9442,N_7747);
and U13098 (N_13098,N_7737,N_7786);
nand U13099 (N_13099,N_5206,N_9465);
and U13100 (N_13100,N_9495,N_8124);
and U13101 (N_13101,N_8455,N_6956);
and U13102 (N_13102,N_7888,N_8051);
nand U13103 (N_13103,N_7285,N_9798);
and U13104 (N_13104,N_9876,N_5757);
and U13105 (N_13105,N_8564,N_7015);
nand U13106 (N_13106,N_9623,N_8193);
nand U13107 (N_13107,N_6761,N_5711);
xnor U13108 (N_13108,N_8068,N_5049);
nand U13109 (N_13109,N_6159,N_5143);
nand U13110 (N_13110,N_9238,N_7353);
nor U13111 (N_13111,N_6437,N_9511);
or U13112 (N_13112,N_8436,N_5787);
nor U13113 (N_13113,N_8400,N_8011);
and U13114 (N_13114,N_5449,N_7882);
and U13115 (N_13115,N_8295,N_5839);
nand U13116 (N_13116,N_6300,N_7360);
and U13117 (N_13117,N_5614,N_7418);
and U13118 (N_13118,N_8564,N_6597);
xnor U13119 (N_13119,N_8098,N_5974);
nand U13120 (N_13120,N_7421,N_7880);
or U13121 (N_13121,N_7910,N_5714);
xnor U13122 (N_13122,N_8116,N_8028);
or U13123 (N_13123,N_5857,N_7300);
xnor U13124 (N_13124,N_8983,N_7007);
nor U13125 (N_13125,N_7293,N_8862);
or U13126 (N_13126,N_6242,N_7982);
nand U13127 (N_13127,N_8567,N_9890);
nand U13128 (N_13128,N_9910,N_5159);
nor U13129 (N_13129,N_5284,N_5050);
or U13130 (N_13130,N_8334,N_9694);
and U13131 (N_13131,N_8956,N_8521);
nand U13132 (N_13132,N_6419,N_8188);
nor U13133 (N_13133,N_9653,N_7243);
or U13134 (N_13134,N_9567,N_7741);
nor U13135 (N_13135,N_9163,N_6717);
or U13136 (N_13136,N_9271,N_6765);
and U13137 (N_13137,N_9167,N_8877);
and U13138 (N_13138,N_9591,N_8738);
and U13139 (N_13139,N_8626,N_8176);
and U13140 (N_13140,N_8976,N_7834);
nand U13141 (N_13141,N_8350,N_9741);
nand U13142 (N_13142,N_9206,N_9200);
and U13143 (N_13143,N_7613,N_9124);
or U13144 (N_13144,N_7904,N_9484);
and U13145 (N_13145,N_5609,N_9346);
nand U13146 (N_13146,N_5447,N_9126);
xor U13147 (N_13147,N_7263,N_7232);
and U13148 (N_13148,N_9334,N_5532);
nor U13149 (N_13149,N_5195,N_5641);
nand U13150 (N_13150,N_9441,N_6345);
nor U13151 (N_13151,N_6298,N_8744);
nand U13152 (N_13152,N_9992,N_9893);
or U13153 (N_13153,N_9450,N_6518);
and U13154 (N_13154,N_8619,N_9294);
or U13155 (N_13155,N_8515,N_5587);
nor U13156 (N_13156,N_9373,N_6002);
or U13157 (N_13157,N_5794,N_6935);
xor U13158 (N_13158,N_7854,N_7068);
nor U13159 (N_13159,N_9084,N_7713);
nor U13160 (N_13160,N_9479,N_7734);
nand U13161 (N_13161,N_5899,N_7437);
nand U13162 (N_13162,N_7503,N_7269);
xor U13163 (N_13163,N_7310,N_7339);
and U13164 (N_13164,N_8048,N_7894);
and U13165 (N_13165,N_5856,N_8970);
nand U13166 (N_13166,N_7989,N_8813);
and U13167 (N_13167,N_8986,N_8872);
nand U13168 (N_13168,N_6412,N_8380);
nand U13169 (N_13169,N_7009,N_8568);
xor U13170 (N_13170,N_6679,N_5072);
nand U13171 (N_13171,N_9548,N_6227);
xnor U13172 (N_13172,N_8188,N_6275);
nand U13173 (N_13173,N_5120,N_8799);
and U13174 (N_13174,N_6900,N_8620);
xor U13175 (N_13175,N_9304,N_7997);
nand U13176 (N_13176,N_5011,N_8484);
nand U13177 (N_13177,N_5527,N_9316);
nor U13178 (N_13178,N_8798,N_5219);
nor U13179 (N_13179,N_5184,N_7534);
nand U13180 (N_13180,N_5707,N_8692);
nand U13181 (N_13181,N_7920,N_6604);
nor U13182 (N_13182,N_7806,N_8551);
or U13183 (N_13183,N_8421,N_7255);
nor U13184 (N_13184,N_8940,N_9175);
and U13185 (N_13185,N_5715,N_5800);
xor U13186 (N_13186,N_5099,N_8323);
or U13187 (N_13187,N_6405,N_6659);
or U13188 (N_13188,N_8520,N_7380);
or U13189 (N_13189,N_8546,N_9999);
nand U13190 (N_13190,N_7289,N_8587);
nand U13191 (N_13191,N_5124,N_5411);
or U13192 (N_13192,N_5470,N_9719);
nand U13193 (N_13193,N_5516,N_5043);
nor U13194 (N_13194,N_6971,N_8177);
xor U13195 (N_13195,N_7786,N_8092);
xor U13196 (N_13196,N_5773,N_9820);
or U13197 (N_13197,N_6342,N_7356);
and U13198 (N_13198,N_5085,N_6782);
xor U13199 (N_13199,N_8764,N_8216);
or U13200 (N_13200,N_9227,N_5327);
or U13201 (N_13201,N_8747,N_6530);
nand U13202 (N_13202,N_8846,N_5757);
and U13203 (N_13203,N_9486,N_8630);
nor U13204 (N_13204,N_6518,N_9110);
nor U13205 (N_13205,N_7130,N_9713);
or U13206 (N_13206,N_7505,N_8745);
nand U13207 (N_13207,N_5769,N_9168);
xnor U13208 (N_13208,N_6460,N_6917);
xor U13209 (N_13209,N_5049,N_6987);
xor U13210 (N_13210,N_8927,N_7091);
nand U13211 (N_13211,N_6042,N_5617);
or U13212 (N_13212,N_7059,N_6104);
or U13213 (N_13213,N_6267,N_7732);
xnor U13214 (N_13214,N_7132,N_6334);
nand U13215 (N_13215,N_5605,N_5018);
and U13216 (N_13216,N_9098,N_7445);
or U13217 (N_13217,N_7684,N_7710);
or U13218 (N_13218,N_5544,N_5209);
or U13219 (N_13219,N_5276,N_5051);
nand U13220 (N_13220,N_7384,N_9385);
and U13221 (N_13221,N_9740,N_5108);
nand U13222 (N_13222,N_7508,N_8929);
nor U13223 (N_13223,N_7188,N_9106);
xnor U13224 (N_13224,N_6466,N_5127);
and U13225 (N_13225,N_7912,N_6792);
nor U13226 (N_13226,N_8325,N_5439);
xnor U13227 (N_13227,N_6585,N_8511);
or U13228 (N_13228,N_9041,N_7923);
nor U13229 (N_13229,N_5188,N_9432);
xnor U13230 (N_13230,N_7094,N_7393);
xnor U13231 (N_13231,N_5643,N_9976);
nor U13232 (N_13232,N_7859,N_6107);
nand U13233 (N_13233,N_9762,N_8237);
nor U13234 (N_13234,N_7958,N_9592);
and U13235 (N_13235,N_6395,N_5099);
nor U13236 (N_13236,N_7607,N_8341);
or U13237 (N_13237,N_8168,N_9833);
and U13238 (N_13238,N_5400,N_8871);
nand U13239 (N_13239,N_6159,N_5783);
or U13240 (N_13240,N_5976,N_5353);
nand U13241 (N_13241,N_8392,N_6485);
nor U13242 (N_13242,N_8377,N_5667);
xnor U13243 (N_13243,N_7857,N_5080);
xnor U13244 (N_13244,N_8043,N_6967);
nand U13245 (N_13245,N_8666,N_9902);
xor U13246 (N_13246,N_5824,N_6662);
nand U13247 (N_13247,N_9653,N_5046);
nor U13248 (N_13248,N_5311,N_9973);
xnor U13249 (N_13249,N_5215,N_6133);
and U13250 (N_13250,N_6336,N_7748);
nand U13251 (N_13251,N_6795,N_5630);
and U13252 (N_13252,N_5032,N_5974);
nor U13253 (N_13253,N_9806,N_9194);
and U13254 (N_13254,N_7381,N_6864);
nor U13255 (N_13255,N_9730,N_6342);
or U13256 (N_13256,N_5733,N_5450);
or U13257 (N_13257,N_7183,N_7307);
nand U13258 (N_13258,N_8242,N_6888);
and U13259 (N_13259,N_7225,N_5178);
nor U13260 (N_13260,N_5147,N_6803);
xnor U13261 (N_13261,N_8048,N_8296);
xor U13262 (N_13262,N_7243,N_5120);
and U13263 (N_13263,N_8268,N_9903);
nand U13264 (N_13264,N_9472,N_8522);
nor U13265 (N_13265,N_6336,N_8466);
nor U13266 (N_13266,N_9854,N_8541);
xnor U13267 (N_13267,N_5382,N_5581);
nor U13268 (N_13268,N_9479,N_6472);
and U13269 (N_13269,N_6505,N_9580);
or U13270 (N_13270,N_5214,N_5879);
and U13271 (N_13271,N_6328,N_5779);
and U13272 (N_13272,N_9255,N_6574);
nand U13273 (N_13273,N_7613,N_9732);
nor U13274 (N_13274,N_9802,N_8190);
and U13275 (N_13275,N_9763,N_5469);
nand U13276 (N_13276,N_7162,N_6933);
and U13277 (N_13277,N_7762,N_7107);
or U13278 (N_13278,N_8567,N_9917);
or U13279 (N_13279,N_6282,N_5500);
nor U13280 (N_13280,N_8244,N_9085);
xnor U13281 (N_13281,N_8686,N_7776);
nand U13282 (N_13282,N_7480,N_7902);
nand U13283 (N_13283,N_9485,N_7185);
nor U13284 (N_13284,N_8178,N_8916);
xor U13285 (N_13285,N_8920,N_8774);
and U13286 (N_13286,N_7857,N_5585);
and U13287 (N_13287,N_5528,N_7711);
or U13288 (N_13288,N_8710,N_6920);
nand U13289 (N_13289,N_5728,N_5763);
and U13290 (N_13290,N_6602,N_9417);
nor U13291 (N_13291,N_9892,N_6727);
nor U13292 (N_13292,N_6324,N_9193);
nor U13293 (N_13293,N_7150,N_6230);
nor U13294 (N_13294,N_6533,N_5927);
nand U13295 (N_13295,N_9496,N_8084);
and U13296 (N_13296,N_7097,N_9112);
nand U13297 (N_13297,N_8787,N_5478);
nor U13298 (N_13298,N_6856,N_8745);
or U13299 (N_13299,N_9345,N_5255);
and U13300 (N_13300,N_6468,N_9916);
or U13301 (N_13301,N_8486,N_9357);
nand U13302 (N_13302,N_9351,N_8845);
and U13303 (N_13303,N_6306,N_5123);
nand U13304 (N_13304,N_7696,N_7764);
and U13305 (N_13305,N_9890,N_8520);
or U13306 (N_13306,N_5298,N_7352);
nand U13307 (N_13307,N_9466,N_8598);
xnor U13308 (N_13308,N_7705,N_8620);
or U13309 (N_13309,N_6235,N_7579);
nor U13310 (N_13310,N_6187,N_5808);
and U13311 (N_13311,N_9606,N_9809);
nor U13312 (N_13312,N_8168,N_8868);
and U13313 (N_13313,N_7060,N_8863);
or U13314 (N_13314,N_9930,N_9035);
nor U13315 (N_13315,N_5354,N_9685);
nand U13316 (N_13316,N_5832,N_5778);
nor U13317 (N_13317,N_5034,N_9547);
or U13318 (N_13318,N_5801,N_6051);
or U13319 (N_13319,N_5434,N_9030);
and U13320 (N_13320,N_7337,N_8781);
and U13321 (N_13321,N_6892,N_5961);
nand U13322 (N_13322,N_6349,N_7688);
or U13323 (N_13323,N_5513,N_9665);
nand U13324 (N_13324,N_8012,N_8403);
nor U13325 (N_13325,N_7721,N_5233);
and U13326 (N_13326,N_7676,N_7242);
and U13327 (N_13327,N_7897,N_5801);
and U13328 (N_13328,N_5389,N_5152);
or U13329 (N_13329,N_8835,N_6200);
nand U13330 (N_13330,N_5904,N_5006);
nand U13331 (N_13331,N_8260,N_9221);
nor U13332 (N_13332,N_7194,N_5040);
nor U13333 (N_13333,N_9271,N_6748);
or U13334 (N_13334,N_7430,N_5635);
nor U13335 (N_13335,N_8077,N_9135);
or U13336 (N_13336,N_9157,N_7878);
or U13337 (N_13337,N_5658,N_9640);
and U13338 (N_13338,N_8288,N_5842);
and U13339 (N_13339,N_9117,N_8171);
nor U13340 (N_13340,N_9986,N_7670);
nor U13341 (N_13341,N_7696,N_6640);
or U13342 (N_13342,N_7452,N_5446);
xor U13343 (N_13343,N_8954,N_7960);
xnor U13344 (N_13344,N_8132,N_8765);
nand U13345 (N_13345,N_6365,N_7349);
nor U13346 (N_13346,N_9014,N_5799);
nor U13347 (N_13347,N_9208,N_6432);
nor U13348 (N_13348,N_5464,N_8318);
or U13349 (N_13349,N_9001,N_9936);
and U13350 (N_13350,N_5953,N_6495);
nand U13351 (N_13351,N_6566,N_9394);
or U13352 (N_13352,N_7286,N_6717);
nor U13353 (N_13353,N_7802,N_7198);
xor U13354 (N_13354,N_7032,N_7604);
nand U13355 (N_13355,N_9418,N_7343);
xor U13356 (N_13356,N_8501,N_9455);
nand U13357 (N_13357,N_6379,N_6371);
or U13358 (N_13358,N_6172,N_8291);
or U13359 (N_13359,N_5492,N_8402);
or U13360 (N_13360,N_6549,N_6407);
and U13361 (N_13361,N_6032,N_8488);
nor U13362 (N_13362,N_6349,N_6089);
or U13363 (N_13363,N_5510,N_9886);
nand U13364 (N_13364,N_9042,N_8670);
or U13365 (N_13365,N_9782,N_8993);
nor U13366 (N_13366,N_5186,N_6807);
or U13367 (N_13367,N_7787,N_5061);
or U13368 (N_13368,N_9996,N_8837);
nor U13369 (N_13369,N_7607,N_7417);
and U13370 (N_13370,N_5627,N_9946);
or U13371 (N_13371,N_8348,N_7494);
nor U13372 (N_13372,N_5413,N_6647);
xor U13373 (N_13373,N_5753,N_5277);
or U13374 (N_13374,N_6586,N_8749);
nand U13375 (N_13375,N_7221,N_9085);
xnor U13376 (N_13376,N_9190,N_9264);
and U13377 (N_13377,N_8105,N_6494);
nand U13378 (N_13378,N_8717,N_6471);
or U13379 (N_13379,N_6436,N_8568);
and U13380 (N_13380,N_9687,N_9369);
xnor U13381 (N_13381,N_8459,N_8940);
nand U13382 (N_13382,N_5017,N_6721);
nand U13383 (N_13383,N_5974,N_7603);
and U13384 (N_13384,N_7819,N_7888);
nor U13385 (N_13385,N_8447,N_9863);
nand U13386 (N_13386,N_9743,N_6751);
and U13387 (N_13387,N_6164,N_6952);
nor U13388 (N_13388,N_7418,N_9088);
nand U13389 (N_13389,N_7434,N_7546);
nand U13390 (N_13390,N_6236,N_9320);
nand U13391 (N_13391,N_7529,N_5812);
nor U13392 (N_13392,N_9045,N_8598);
or U13393 (N_13393,N_6705,N_6907);
and U13394 (N_13394,N_9030,N_8142);
nand U13395 (N_13395,N_9775,N_6450);
nand U13396 (N_13396,N_6285,N_5318);
and U13397 (N_13397,N_5781,N_9523);
nor U13398 (N_13398,N_6129,N_7470);
or U13399 (N_13399,N_8502,N_6315);
nand U13400 (N_13400,N_5359,N_5268);
xor U13401 (N_13401,N_5036,N_5446);
nand U13402 (N_13402,N_9334,N_7101);
xor U13403 (N_13403,N_9836,N_7506);
or U13404 (N_13404,N_8858,N_8941);
nor U13405 (N_13405,N_9331,N_9096);
nand U13406 (N_13406,N_5576,N_8583);
and U13407 (N_13407,N_5535,N_9503);
nand U13408 (N_13408,N_5386,N_9904);
and U13409 (N_13409,N_9450,N_8592);
nand U13410 (N_13410,N_6431,N_9991);
or U13411 (N_13411,N_6303,N_8908);
nor U13412 (N_13412,N_7763,N_8697);
nand U13413 (N_13413,N_6851,N_6717);
xnor U13414 (N_13414,N_7347,N_6600);
nor U13415 (N_13415,N_6291,N_5043);
or U13416 (N_13416,N_8842,N_8074);
nor U13417 (N_13417,N_7663,N_9472);
or U13418 (N_13418,N_9169,N_5842);
xor U13419 (N_13419,N_8398,N_5048);
nand U13420 (N_13420,N_9527,N_8202);
and U13421 (N_13421,N_6271,N_6615);
and U13422 (N_13422,N_7047,N_8564);
nand U13423 (N_13423,N_7643,N_5952);
or U13424 (N_13424,N_7532,N_8649);
or U13425 (N_13425,N_5430,N_7366);
nor U13426 (N_13426,N_7626,N_6624);
and U13427 (N_13427,N_7889,N_6807);
or U13428 (N_13428,N_7632,N_8644);
or U13429 (N_13429,N_7850,N_9907);
and U13430 (N_13430,N_9074,N_9438);
nor U13431 (N_13431,N_8923,N_7167);
nand U13432 (N_13432,N_6032,N_8168);
nand U13433 (N_13433,N_5316,N_6180);
nor U13434 (N_13434,N_7599,N_6329);
nand U13435 (N_13435,N_9101,N_7099);
nor U13436 (N_13436,N_7079,N_6643);
nand U13437 (N_13437,N_8985,N_9913);
nor U13438 (N_13438,N_9178,N_6678);
and U13439 (N_13439,N_5736,N_6037);
nand U13440 (N_13440,N_6979,N_5303);
or U13441 (N_13441,N_7581,N_8202);
nor U13442 (N_13442,N_8149,N_9978);
or U13443 (N_13443,N_8296,N_9176);
nand U13444 (N_13444,N_5073,N_6924);
and U13445 (N_13445,N_7896,N_8845);
nor U13446 (N_13446,N_6005,N_9751);
and U13447 (N_13447,N_6564,N_7236);
or U13448 (N_13448,N_6297,N_6769);
nor U13449 (N_13449,N_5935,N_9524);
nand U13450 (N_13450,N_5660,N_7188);
and U13451 (N_13451,N_8842,N_5824);
nand U13452 (N_13452,N_8030,N_5123);
or U13453 (N_13453,N_8899,N_8163);
nor U13454 (N_13454,N_5595,N_7859);
and U13455 (N_13455,N_8030,N_6762);
nand U13456 (N_13456,N_6393,N_7174);
nand U13457 (N_13457,N_7640,N_5189);
nand U13458 (N_13458,N_7162,N_5274);
or U13459 (N_13459,N_5435,N_8728);
xor U13460 (N_13460,N_5748,N_5626);
and U13461 (N_13461,N_5244,N_9861);
nand U13462 (N_13462,N_8706,N_9477);
or U13463 (N_13463,N_5204,N_5727);
and U13464 (N_13464,N_5924,N_6912);
nand U13465 (N_13465,N_8112,N_6434);
xor U13466 (N_13466,N_5347,N_5737);
nor U13467 (N_13467,N_5591,N_5840);
nor U13468 (N_13468,N_8344,N_8002);
nor U13469 (N_13469,N_5749,N_9972);
nor U13470 (N_13470,N_8610,N_5029);
nand U13471 (N_13471,N_8737,N_8211);
and U13472 (N_13472,N_7033,N_6155);
and U13473 (N_13473,N_6155,N_8629);
or U13474 (N_13474,N_6411,N_6097);
nand U13475 (N_13475,N_8743,N_5365);
or U13476 (N_13476,N_5805,N_7695);
xnor U13477 (N_13477,N_5792,N_6697);
nand U13478 (N_13478,N_7119,N_7246);
or U13479 (N_13479,N_5560,N_6017);
or U13480 (N_13480,N_9250,N_6517);
and U13481 (N_13481,N_5472,N_9708);
or U13482 (N_13482,N_5581,N_9370);
and U13483 (N_13483,N_8431,N_8170);
xnor U13484 (N_13484,N_5941,N_6510);
or U13485 (N_13485,N_5405,N_5820);
and U13486 (N_13486,N_5052,N_8023);
and U13487 (N_13487,N_9561,N_6790);
or U13488 (N_13488,N_5416,N_8503);
or U13489 (N_13489,N_6281,N_6428);
or U13490 (N_13490,N_8198,N_7003);
nor U13491 (N_13491,N_6271,N_6184);
xor U13492 (N_13492,N_9030,N_8059);
and U13493 (N_13493,N_8565,N_6074);
and U13494 (N_13494,N_9368,N_6685);
nand U13495 (N_13495,N_5249,N_7122);
nor U13496 (N_13496,N_5339,N_5930);
and U13497 (N_13497,N_7892,N_6570);
or U13498 (N_13498,N_7865,N_7600);
nand U13499 (N_13499,N_8531,N_6282);
nor U13500 (N_13500,N_9810,N_6302);
nand U13501 (N_13501,N_5312,N_8596);
nor U13502 (N_13502,N_7161,N_8801);
and U13503 (N_13503,N_6437,N_9727);
or U13504 (N_13504,N_8398,N_7841);
nand U13505 (N_13505,N_6827,N_8081);
xor U13506 (N_13506,N_6753,N_5082);
nand U13507 (N_13507,N_5838,N_8458);
nand U13508 (N_13508,N_5658,N_7831);
or U13509 (N_13509,N_7064,N_9332);
nand U13510 (N_13510,N_8445,N_8539);
and U13511 (N_13511,N_5538,N_9769);
nand U13512 (N_13512,N_5089,N_9051);
nand U13513 (N_13513,N_6208,N_9702);
and U13514 (N_13514,N_7823,N_6129);
nor U13515 (N_13515,N_5719,N_7015);
nor U13516 (N_13516,N_6397,N_9573);
nor U13517 (N_13517,N_6537,N_6945);
nand U13518 (N_13518,N_6914,N_6355);
nor U13519 (N_13519,N_6187,N_6036);
nor U13520 (N_13520,N_5023,N_7085);
or U13521 (N_13521,N_6227,N_9815);
xor U13522 (N_13522,N_7950,N_9579);
and U13523 (N_13523,N_5517,N_7027);
nor U13524 (N_13524,N_5259,N_9196);
or U13525 (N_13525,N_6231,N_9423);
xor U13526 (N_13526,N_5235,N_8568);
nor U13527 (N_13527,N_8174,N_7585);
nand U13528 (N_13528,N_6166,N_9702);
and U13529 (N_13529,N_6196,N_8358);
and U13530 (N_13530,N_6371,N_9123);
nand U13531 (N_13531,N_5130,N_6301);
nand U13532 (N_13532,N_5959,N_8460);
nand U13533 (N_13533,N_5143,N_5098);
nor U13534 (N_13534,N_8903,N_7758);
and U13535 (N_13535,N_5276,N_8687);
and U13536 (N_13536,N_7760,N_8101);
xnor U13537 (N_13537,N_8574,N_8560);
and U13538 (N_13538,N_5070,N_7597);
nor U13539 (N_13539,N_7713,N_9773);
nand U13540 (N_13540,N_8086,N_5207);
nand U13541 (N_13541,N_5711,N_6181);
xnor U13542 (N_13542,N_8803,N_7791);
nand U13543 (N_13543,N_6927,N_9207);
and U13544 (N_13544,N_6421,N_9761);
nand U13545 (N_13545,N_5900,N_9319);
nand U13546 (N_13546,N_7083,N_5293);
and U13547 (N_13547,N_6924,N_6384);
nand U13548 (N_13548,N_5105,N_7720);
or U13549 (N_13549,N_6602,N_9601);
or U13550 (N_13550,N_8370,N_8115);
and U13551 (N_13551,N_6287,N_8852);
nand U13552 (N_13552,N_9546,N_7408);
nor U13553 (N_13553,N_7561,N_7167);
or U13554 (N_13554,N_5285,N_8997);
xnor U13555 (N_13555,N_5926,N_7535);
nor U13556 (N_13556,N_5861,N_8312);
nor U13557 (N_13557,N_8193,N_9937);
nor U13558 (N_13558,N_8799,N_6043);
nand U13559 (N_13559,N_7150,N_7650);
nand U13560 (N_13560,N_9624,N_8350);
nand U13561 (N_13561,N_9242,N_5774);
and U13562 (N_13562,N_6321,N_8694);
and U13563 (N_13563,N_9580,N_5504);
nor U13564 (N_13564,N_7882,N_8293);
nand U13565 (N_13565,N_9522,N_8860);
nand U13566 (N_13566,N_5847,N_6724);
xnor U13567 (N_13567,N_5237,N_5951);
xor U13568 (N_13568,N_5470,N_9557);
and U13569 (N_13569,N_7769,N_9476);
or U13570 (N_13570,N_8173,N_9206);
nor U13571 (N_13571,N_8157,N_7554);
or U13572 (N_13572,N_8226,N_5785);
or U13573 (N_13573,N_6624,N_8011);
and U13574 (N_13574,N_8825,N_9349);
nor U13575 (N_13575,N_7561,N_5587);
xnor U13576 (N_13576,N_6614,N_8122);
and U13577 (N_13577,N_9364,N_6878);
or U13578 (N_13578,N_7206,N_5986);
and U13579 (N_13579,N_7447,N_7528);
or U13580 (N_13580,N_7465,N_7819);
and U13581 (N_13581,N_5772,N_5863);
and U13582 (N_13582,N_8588,N_6225);
or U13583 (N_13583,N_6760,N_5767);
nor U13584 (N_13584,N_8555,N_7192);
xor U13585 (N_13585,N_8628,N_6900);
nor U13586 (N_13586,N_8959,N_8786);
nor U13587 (N_13587,N_9598,N_8552);
or U13588 (N_13588,N_8142,N_8995);
or U13589 (N_13589,N_7663,N_8731);
nor U13590 (N_13590,N_5767,N_5257);
or U13591 (N_13591,N_5272,N_8775);
nor U13592 (N_13592,N_7453,N_7161);
or U13593 (N_13593,N_5176,N_6412);
nand U13594 (N_13594,N_8614,N_7322);
nor U13595 (N_13595,N_6589,N_7241);
xnor U13596 (N_13596,N_6904,N_9980);
nor U13597 (N_13597,N_6032,N_5641);
or U13598 (N_13598,N_7881,N_5567);
or U13599 (N_13599,N_9596,N_8287);
nor U13600 (N_13600,N_5745,N_6486);
and U13601 (N_13601,N_9379,N_7952);
and U13602 (N_13602,N_8252,N_7794);
nor U13603 (N_13603,N_9258,N_6110);
nand U13604 (N_13604,N_9250,N_6934);
and U13605 (N_13605,N_7890,N_7327);
nand U13606 (N_13606,N_7391,N_6680);
or U13607 (N_13607,N_8243,N_5401);
nor U13608 (N_13608,N_5142,N_9615);
nor U13609 (N_13609,N_9185,N_5292);
or U13610 (N_13610,N_5367,N_8931);
nand U13611 (N_13611,N_9117,N_7461);
or U13612 (N_13612,N_7848,N_9490);
and U13613 (N_13613,N_9831,N_8937);
or U13614 (N_13614,N_9366,N_7301);
and U13615 (N_13615,N_6812,N_7669);
and U13616 (N_13616,N_6772,N_5866);
or U13617 (N_13617,N_5333,N_6452);
nand U13618 (N_13618,N_7059,N_7863);
or U13619 (N_13619,N_8757,N_6231);
nor U13620 (N_13620,N_8269,N_9777);
nor U13621 (N_13621,N_9125,N_8548);
nand U13622 (N_13622,N_6037,N_7236);
or U13623 (N_13623,N_9116,N_8715);
xor U13624 (N_13624,N_9556,N_8857);
or U13625 (N_13625,N_9892,N_7359);
nor U13626 (N_13626,N_9791,N_9323);
and U13627 (N_13627,N_9307,N_8883);
nand U13628 (N_13628,N_6443,N_9898);
and U13629 (N_13629,N_6339,N_5462);
and U13630 (N_13630,N_5809,N_8453);
or U13631 (N_13631,N_7482,N_8190);
or U13632 (N_13632,N_5354,N_9650);
or U13633 (N_13633,N_8555,N_6253);
and U13634 (N_13634,N_7257,N_8944);
nand U13635 (N_13635,N_9573,N_5593);
nor U13636 (N_13636,N_6331,N_8138);
nor U13637 (N_13637,N_8666,N_8911);
nand U13638 (N_13638,N_6240,N_5130);
or U13639 (N_13639,N_7496,N_5396);
and U13640 (N_13640,N_8628,N_6549);
or U13641 (N_13641,N_6242,N_9663);
or U13642 (N_13642,N_9880,N_8039);
and U13643 (N_13643,N_5731,N_5662);
and U13644 (N_13644,N_7331,N_7176);
and U13645 (N_13645,N_9057,N_5053);
or U13646 (N_13646,N_6289,N_7983);
nand U13647 (N_13647,N_9918,N_5198);
or U13648 (N_13648,N_6134,N_6153);
nor U13649 (N_13649,N_5982,N_9022);
or U13650 (N_13650,N_6245,N_7476);
nand U13651 (N_13651,N_8730,N_9834);
nor U13652 (N_13652,N_9205,N_8100);
and U13653 (N_13653,N_9175,N_7877);
nand U13654 (N_13654,N_5785,N_8273);
or U13655 (N_13655,N_8425,N_9520);
nand U13656 (N_13656,N_6356,N_9645);
nor U13657 (N_13657,N_9761,N_9612);
nor U13658 (N_13658,N_7786,N_9169);
xnor U13659 (N_13659,N_9074,N_9143);
nor U13660 (N_13660,N_8605,N_5502);
nand U13661 (N_13661,N_9010,N_5316);
or U13662 (N_13662,N_8314,N_5202);
nor U13663 (N_13663,N_5931,N_5939);
xnor U13664 (N_13664,N_8919,N_5799);
and U13665 (N_13665,N_6860,N_7307);
or U13666 (N_13666,N_6210,N_5406);
nand U13667 (N_13667,N_8788,N_6613);
and U13668 (N_13668,N_9739,N_5220);
nand U13669 (N_13669,N_8896,N_5023);
nor U13670 (N_13670,N_5508,N_6592);
or U13671 (N_13671,N_8757,N_5137);
nand U13672 (N_13672,N_7342,N_5335);
or U13673 (N_13673,N_7918,N_6308);
or U13674 (N_13674,N_6931,N_6089);
or U13675 (N_13675,N_7771,N_5381);
nand U13676 (N_13676,N_8179,N_7809);
and U13677 (N_13677,N_8145,N_6886);
and U13678 (N_13678,N_7317,N_9869);
nor U13679 (N_13679,N_8383,N_7635);
nor U13680 (N_13680,N_8791,N_6819);
and U13681 (N_13681,N_9960,N_8603);
xor U13682 (N_13682,N_9428,N_9665);
nor U13683 (N_13683,N_7990,N_8995);
xor U13684 (N_13684,N_7785,N_9031);
nand U13685 (N_13685,N_5625,N_5275);
and U13686 (N_13686,N_7214,N_6917);
and U13687 (N_13687,N_7572,N_6788);
or U13688 (N_13688,N_6970,N_7331);
or U13689 (N_13689,N_9868,N_8529);
nor U13690 (N_13690,N_9022,N_6154);
and U13691 (N_13691,N_7942,N_9212);
xnor U13692 (N_13692,N_7829,N_5704);
or U13693 (N_13693,N_5230,N_5877);
and U13694 (N_13694,N_6477,N_5877);
nor U13695 (N_13695,N_6672,N_6666);
nand U13696 (N_13696,N_6774,N_8226);
nor U13697 (N_13697,N_8000,N_7858);
nand U13698 (N_13698,N_6263,N_7450);
nand U13699 (N_13699,N_6910,N_8504);
nand U13700 (N_13700,N_7837,N_8544);
nand U13701 (N_13701,N_7015,N_9440);
or U13702 (N_13702,N_6455,N_6360);
nor U13703 (N_13703,N_8051,N_8283);
and U13704 (N_13704,N_6762,N_7239);
or U13705 (N_13705,N_9489,N_5757);
nand U13706 (N_13706,N_8760,N_8843);
nand U13707 (N_13707,N_5941,N_5058);
nor U13708 (N_13708,N_6256,N_5000);
nor U13709 (N_13709,N_9231,N_7933);
or U13710 (N_13710,N_5237,N_9216);
xnor U13711 (N_13711,N_9789,N_6459);
or U13712 (N_13712,N_5656,N_9556);
nand U13713 (N_13713,N_5016,N_5538);
nand U13714 (N_13714,N_7154,N_8172);
nor U13715 (N_13715,N_8377,N_7795);
and U13716 (N_13716,N_7059,N_6434);
or U13717 (N_13717,N_8712,N_5731);
nand U13718 (N_13718,N_6061,N_6739);
nand U13719 (N_13719,N_6927,N_5059);
nor U13720 (N_13720,N_9781,N_7112);
and U13721 (N_13721,N_5375,N_8162);
and U13722 (N_13722,N_5251,N_6552);
and U13723 (N_13723,N_9994,N_7142);
nand U13724 (N_13724,N_6823,N_9877);
nand U13725 (N_13725,N_5754,N_7845);
and U13726 (N_13726,N_7359,N_9492);
nor U13727 (N_13727,N_5930,N_6483);
nand U13728 (N_13728,N_8395,N_9221);
nand U13729 (N_13729,N_8285,N_6346);
and U13730 (N_13730,N_9405,N_8430);
and U13731 (N_13731,N_8759,N_9083);
nand U13732 (N_13732,N_9276,N_5772);
nor U13733 (N_13733,N_9098,N_7926);
nor U13734 (N_13734,N_9556,N_5801);
nand U13735 (N_13735,N_5724,N_9906);
and U13736 (N_13736,N_7071,N_5031);
nor U13737 (N_13737,N_6028,N_5345);
nand U13738 (N_13738,N_5123,N_8414);
nand U13739 (N_13739,N_5777,N_5259);
or U13740 (N_13740,N_5273,N_7183);
and U13741 (N_13741,N_5010,N_6889);
xor U13742 (N_13742,N_9116,N_6623);
or U13743 (N_13743,N_5848,N_8042);
nand U13744 (N_13744,N_6553,N_7077);
and U13745 (N_13745,N_9333,N_7360);
nor U13746 (N_13746,N_7791,N_6568);
xor U13747 (N_13747,N_5845,N_5934);
and U13748 (N_13748,N_9485,N_6436);
nor U13749 (N_13749,N_7878,N_7501);
nand U13750 (N_13750,N_9157,N_9110);
and U13751 (N_13751,N_5664,N_6056);
nor U13752 (N_13752,N_5790,N_5508);
or U13753 (N_13753,N_7109,N_9948);
or U13754 (N_13754,N_5643,N_9470);
or U13755 (N_13755,N_6090,N_5233);
nor U13756 (N_13756,N_6476,N_8039);
and U13757 (N_13757,N_8041,N_5284);
nand U13758 (N_13758,N_9883,N_6981);
nor U13759 (N_13759,N_7962,N_5442);
xnor U13760 (N_13760,N_7282,N_5474);
nand U13761 (N_13761,N_9994,N_7631);
nor U13762 (N_13762,N_7714,N_8596);
or U13763 (N_13763,N_5600,N_8508);
and U13764 (N_13764,N_7089,N_9628);
and U13765 (N_13765,N_7895,N_8754);
or U13766 (N_13766,N_8602,N_6874);
nand U13767 (N_13767,N_9707,N_6941);
nand U13768 (N_13768,N_8409,N_7431);
nor U13769 (N_13769,N_8799,N_7825);
or U13770 (N_13770,N_9247,N_8626);
nor U13771 (N_13771,N_7052,N_6080);
nand U13772 (N_13772,N_7431,N_5583);
xnor U13773 (N_13773,N_8820,N_6101);
and U13774 (N_13774,N_6123,N_9063);
nand U13775 (N_13775,N_6520,N_6287);
or U13776 (N_13776,N_9182,N_9060);
nand U13777 (N_13777,N_8120,N_7916);
or U13778 (N_13778,N_9400,N_7009);
and U13779 (N_13779,N_9689,N_6686);
xor U13780 (N_13780,N_7451,N_6089);
xnor U13781 (N_13781,N_8927,N_6819);
or U13782 (N_13782,N_9107,N_6843);
or U13783 (N_13783,N_8917,N_9257);
nor U13784 (N_13784,N_7819,N_5006);
nand U13785 (N_13785,N_5040,N_7752);
xnor U13786 (N_13786,N_6767,N_6271);
and U13787 (N_13787,N_6082,N_6233);
or U13788 (N_13788,N_6954,N_8302);
or U13789 (N_13789,N_9100,N_8853);
xor U13790 (N_13790,N_5535,N_9826);
nand U13791 (N_13791,N_7064,N_7082);
or U13792 (N_13792,N_6292,N_9320);
nor U13793 (N_13793,N_5746,N_6364);
and U13794 (N_13794,N_7437,N_5658);
nor U13795 (N_13795,N_6161,N_7460);
nor U13796 (N_13796,N_7520,N_7105);
nor U13797 (N_13797,N_7866,N_6131);
nand U13798 (N_13798,N_5687,N_6962);
nor U13799 (N_13799,N_8580,N_6763);
nand U13800 (N_13800,N_9422,N_8273);
and U13801 (N_13801,N_7270,N_8839);
or U13802 (N_13802,N_7907,N_6326);
and U13803 (N_13803,N_7385,N_5585);
nand U13804 (N_13804,N_7673,N_9277);
and U13805 (N_13805,N_5661,N_7510);
nor U13806 (N_13806,N_9158,N_7769);
or U13807 (N_13807,N_7783,N_6770);
nor U13808 (N_13808,N_9763,N_9328);
and U13809 (N_13809,N_9449,N_7179);
nor U13810 (N_13810,N_6766,N_6485);
and U13811 (N_13811,N_8421,N_6203);
nand U13812 (N_13812,N_5282,N_9949);
or U13813 (N_13813,N_5186,N_7403);
nor U13814 (N_13814,N_7845,N_6575);
nor U13815 (N_13815,N_9712,N_5883);
and U13816 (N_13816,N_9349,N_7071);
nand U13817 (N_13817,N_6394,N_8817);
or U13818 (N_13818,N_5363,N_9756);
nor U13819 (N_13819,N_9902,N_9451);
xnor U13820 (N_13820,N_9313,N_5575);
nand U13821 (N_13821,N_5734,N_8219);
and U13822 (N_13822,N_9462,N_8321);
and U13823 (N_13823,N_5201,N_5758);
nor U13824 (N_13824,N_6134,N_9943);
nand U13825 (N_13825,N_8233,N_7342);
nand U13826 (N_13826,N_5893,N_7089);
nor U13827 (N_13827,N_5566,N_5671);
nor U13828 (N_13828,N_6452,N_5918);
and U13829 (N_13829,N_9137,N_9544);
nand U13830 (N_13830,N_9823,N_8195);
nor U13831 (N_13831,N_8479,N_8730);
xor U13832 (N_13832,N_7681,N_9473);
or U13833 (N_13833,N_9377,N_6215);
or U13834 (N_13834,N_6086,N_5651);
or U13835 (N_13835,N_7150,N_7017);
nand U13836 (N_13836,N_7312,N_5133);
nor U13837 (N_13837,N_8782,N_7077);
and U13838 (N_13838,N_7063,N_6933);
nand U13839 (N_13839,N_6500,N_7875);
nor U13840 (N_13840,N_9112,N_7398);
and U13841 (N_13841,N_5460,N_5981);
nand U13842 (N_13842,N_5731,N_8024);
and U13843 (N_13843,N_8845,N_8660);
nor U13844 (N_13844,N_7090,N_5951);
nor U13845 (N_13845,N_7560,N_6624);
or U13846 (N_13846,N_5253,N_8076);
nor U13847 (N_13847,N_7928,N_6713);
xor U13848 (N_13848,N_9531,N_7989);
and U13849 (N_13849,N_9665,N_7876);
and U13850 (N_13850,N_5472,N_8582);
nor U13851 (N_13851,N_6931,N_9464);
nand U13852 (N_13852,N_8152,N_7163);
xnor U13853 (N_13853,N_9407,N_6794);
or U13854 (N_13854,N_5310,N_8995);
nand U13855 (N_13855,N_7419,N_8414);
or U13856 (N_13856,N_8187,N_8768);
nor U13857 (N_13857,N_7041,N_6857);
and U13858 (N_13858,N_7888,N_8118);
or U13859 (N_13859,N_7852,N_5318);
nand U13860 (N_13860,N_7581,N_5943);
and U13861 (N_13861,N_5246,N_6598);
nand U13862 (N_13862,N_5070,N_8753);
xor U13863 (N_13863,N_8553,N_7375);
xor U13864 (N_13864,N_7249,N_8996);
nand U13865 (N_13865,N_7273,N_9993);
nor U13866 (N_13866,N_6622,N_7279);
nand U13867 (N_13867,N_5398,N_6038);
or U13868 (N_13868,N_5308,N_6885);
or U13869 (N_13869,N_7375,N_5750);
nand U13870 (N_13870,N_8033,N_9304);
nand U13871 (N_13871,N_8167,N_9620);
and U13872 (N_13872,N_6866,N_7462);
nand U13873 (N_13873,N_7821,N_8660);
and U13874 (N_13874,N_9778,N_8702);
nand U13875 (N_13875,N_5891,N_5864);
or U13876 (N_13876,N_8902,N_7006);
xor U13877 (N_13877,N_8223,N_5438);
nand U13878 (N_13878,N_6709,N_6066);
nand U13879 (N_13879,N_5312,N_6173);
nand U13880 (N_13880,N_6451,N_7903);
nand U13881 (N_13881,N_9324,N_8688);
nand U13882 (N_13882,N_8698,N_8151);
xnor U13883 (N_13883,N_9465,N_5811);
and U13884 (N_13884,N_5605,N_9015);
nand U13885 (N_13885,N_8078,N_6971);
nand U13886 (N_13886,N_6605,N_8817);
xnor U13887 (N_13887,N_9026,N_9002);
nand U13888 (N_13888,N_6400,N_7249);
and U13889 (N_13889,N_6477,N_7554);
and U13890 (N_13890,N_6877,N_8419);
or U13891 (N_13891,N_7966,N_7022);
or U13892 (N_13892,N_9706,N_8777);
and U13893 (N_13893,N_5926,N_5764);
or U13894 (N_13894,N_5956,N_6594);
and U13895 (N_13895,N_8348,N_9438);
nand U13896 (N_13896,N_8380,N_6669);
nand U13897 (N_13897,N_9348,N_9573);
and U13898 (N_13898,N_9125,N_7300);
nand U13899 (N_13899,N_7562,N_5631);
nand U13900 (N_13900,N_9355,N_9154);
or U13901 (N_13901,N_5915,N_6948);
nand U13902 (N_13902,N_9744,N_7275);
nor U13903 (N_13903,N_7848,N_5462);
nor U13904 (N_13904,N_9351,N_6897);
nor U13905 (N_13905,N_9426,N_7827);
nor U13906 (N_13906,N_9738,N_5125);
or U13907 (N_13907,N_9847,N_5270);
or U13908 (N_13908,N_8007,N_8425);
nand U13909 (N_13909,N_8296,N_8300);
nor U13910 (N_13910,N_6964,N_5338);
and U13911 (N_13911,N_5564,N_6537);
nor U13912 (N_13912,N_9125,N_8993);
nand U13913 (N_13913,N_8830,N_7516);
nor U13914 (N_13914,N_5935,N_5665);
or U13915 (N_13915,N_8349,N_8926);
or U13916 (N_13916,N_9851,N_9975);
and U13917 (N_13917,N_5711,N_5523);
or U13918 (N_13918,N_7183,N_7268);
and U13919 (N_13919,N_5817,N_9533);
and U13920 (N_13920,N_9805,N_8563);
nor U13921 (N_13921,N_6529,N_7249);
nand U13922 (N_13922,N_9197,N_8564);
and U13923 (N_13923,N_5267,N_7935);
xor U13924 (N_13924,N_9137,N_8552);
nor U13925 (N_13925,N_5384,N_9722);
or U13926 (N_13926,N_5020,N_7329);
nand U13927 (N_13927,N_8379,N_8786);
or U13928 (N_13928,N_9796,N_5012);
xor U13929 (N_13929,N_8775,N_7493);
xor U13930 (N_13930,N_7040,N_8572);
xor U13931 (N_13931,N_6086,N_7703);
nor U13932 (N_13932,N_9120,N_5700);
nor U13933 (N_13933,N_8942,N_5190);
or U13934 (N_13934,N_8951,N_6536);
and U13935 (N_13935,N_8058,N_7617);
and U13936 (N_13936,N_5849,N_7663);
or U13937 (N_13937,N_9070,N_9251);
nor U13938 (N_13938,N_5395,N_6041);
xnor U13939 (N_13939,N_8901,N_8476);
or U13940 (N_13940,N_5163,N_8161);
nor U13941 (N_13941,N_9021,N_6801);
or U13942 (N_13942,N_5994,N_5723);
and U13943 (N_13943,N_5213,N_7873);
nor U13944 (N_13944,N_8033,N_8383);
and U13945 (N_13945,N_7570,N_7597);
or U13946 (N_13946,N_5396,N_5533);
nor U13947 (N_13947,N_8965,N_6687);
nand U13948 (N_13948,N_9175,N_7634);
nand U13949 (N_13949,N_5779,N_9560);
nor U13950 (N_13950,N_9706,N_5027);
nor U13951 (N_13951,N_8671,N_7042);
or U13952 (N_13952,N_5248,N_5975);
nor U13953 (N_13953,N_5859,N_8913);
or U13954 (N_13954,N_7180,N_8410);
and U13955 (N_13955,N_7011,N_8364);
or U13956 (N_13956,N_8088,N_7223);
nor U13957 (N_13957,N_8246,N_9021);
or U13958 (N_13958,N_6172,N_8304);
nand U13959 (N_13959,N_9794,N_7604);
or U13960 (N_13960,N_5979,N_5008);
nor U13961 (N_13961,N_8368,N_9832);
nor U13962 (N_13962,N_8163,N_9015);
xor U13963 (N_13963,N_9508,N_7411);
or U13964 (N_13964,N_8916,N_5522);
xor U13965 (N_13965,N_5613,N_5124);
xnor U13966 (N_13966,N_9577,N_6073);
nand U13967 (N_13967,N_9678,N_7264);
nand U13968 (N_13968,N_7341,N_5938);
and U13969 (N_13969,N_6285,N_5564);
nand U13970 (N_13970,N_9328,N_8888);
xor U13971 (N_13971,N_5422,N_8148);
nand U13972 (N_13972,N_7412,N_9263);
nor U13973 (N_13973,N_6732,N_8745);
nor U13974 (N_13974,N_5985,N_9857);
nand U13975 (N_13975,N_8085,N_7973);
or U13976 (N_13976,N_9167,N_9568);
nor U13977 (N_13977,N_9213,N_9017);
nor U13978 (N_13978,N_9109,N_7374);
and U13979 (N_13979,N_9057,N_5645);
or U13980 (N_13980,N_8841,N_9803);
xor U13981 (N_13981,N_5228,N_5326);
nand U13982 (N_13982,N_6277,N_9055);
or U13983 (N_13983,N_6569,N_5101);
and U13984 (N_13984,N_6414,N_7497);
and U13985 (N_13985,N_8309,N_6644);
and U13986 (N_13986,N_5840,N_7897);
nor U13987 (N_13987,N_7772,N_9006);
or U13988 (N_13988,N_8546,N_7736);
nand U13989 (N_13989,N_6227,N_7514);
or U13990 (N_13990,N_7881,N_8854);
or U13991 (N_13991,N_8352,N_8993);
or U13992 (N_13992,N_5453,N_5135);
or U13993 (N_13993,N_9998,N_9776);
nor U13994 (N_13994,N_5232,N_6558);
nor U13995 (N_13995,N_9509,N_7902);
nand U13996 (N_13996,N_5921,N_5643);
nand U13997 (N_13997,N_8430,N_7462);
nand U13998 (N_13998,N_8297,N_6709);
xor U13999 (N_13999,N_7753,N_8586);
or U14000 (N_14000,N_9931,N_9042);
nand U14001 (N_14001,N_8947,N_7611);
and U14002 (N_14002,N_8611,N_7609);
nand U14003 (N_14003,N_6282,N_5189);
xnor U14004 (N_14004,N_8289,N_9206);
nor U14005 (N_14005,N_8549,N_9447);
xor U14006 (N_14006,N_5581,N_5696);
or U14007 (N_14007,N_7832,N_8832);
nand U14008 (N_14008,N_8754,N_8309);
nor U14009 (N_14009,N_8986,N_8377);
xor U14010 (N_14010,N_8145,N_9970);
nor U14011 (N_14011,N_5177,N_5682);
and U14012 (N_14012,N_8352,N_8615);
and U14013 (N_14013,N_9756,N_8857);
or U14014 (N_14014,N_6010,N_5422);
nor U14015 (N_14015,N_8789,N_8696);
nand U14016 (N_14016,N_7810,N_7207);
or U14017 (N_14017,N_5998,N_9858);
or U14018 (N_14018,N_6030,N_9161);
nand U14019 (N_14019,N_7242,N_8916);
or U14020 (N_14020,N_9043,N_9493);
nand U14021 (N_14021,N_7632,N_7007);
and U14022 (N_14022,N_9949,N_6043);
or U14023 (N_14023,N_6662,N_8749);
or U14024 (N_14024,N_8213,N_5103);
nor U14025 (N_14025,N_9654,N_7278);
nor U14026 (N_14026,N_9656,N_7957);
and U14027 (N_14027,N_7811,N_8221);
nor U14028 (N_14028,N_6123,N_8459);
nand U14029 (N_14029,N_6641,N_9485);
nand U14030 (N_14030,N_8732,N_8784);
or U14031 (N_14031,N_9314,N_5599);
nand U14032 (N_14032,N_9279,N_6016);
and U14033 (N_14033,N_9190,N_7815);
nor U14034 (N_14034,N_7129,N_5086);
nand U14035 (N_14035,N_8534,N_5339);
xor U14036 (N_14036,N_8951,N_6899);
or U14037 (N_14037,N_6791,N_6057);
nor U14038 (N_14038,N_9026,N_9896);
xor U14039 (N_14039,N_5246,N_5431);
xor U14040 (N_14040,N_6847,N_6089);
nand U14041 (N_14041,N_6606,N_7435);
and U14042 (N_14042,N_9593,N_9377);
and U14043 (N_14043,N_6477,N_6830);
xnor U14044 (N_14044,N_6558,N_6852);
and U14045 (N_14045,N_8120,N_7726);
or U14046 (N_14046,N_9862,N_5163);
or U14047 (N_14047,N_9313,N_6801);
and U14048 (N_14048,N_8054,N_6448);
or U14049 (N_14049,N_5291,N_8144);
nand U14050 (N_14050,N_6801,N_7758);
xnor U14051 (N_14051,N_7090,N_7425);
xnor U14052 (N_14052,N_8697,N_7465);
xnor U14053 (N_14053,N_5536,N_9106);
and U14054 (N_14054,N_8677,N_7099);
and U14055 (N_14055,N_5582,N_8617);
nor U14056 (N_14056,N_7441,N_8387);
and U14057 (N_14057,N_9141,N_5512);
xnor U14058 (N_14058,N_6354,N_7537);
and U14059 (N_14059,N_6391,N_5224);
nor U14060 (N_14060,N_9392,N_6634);
nand U14061 (N_14061,N_5289,N_7997);
nand U14062 (N_14062,N_9027,N_7451);
xnor U14063 (N_14063,N_9616,N_8499);
nand U14064 (N_14064,N_9173,N_8822);
nor U14065 (N_14065,N_7781,N_5564);
or U14066 (N_14066,N_8922,N_6351);
and U14067 (N_14067,N_9503,N_6533);
and U14068 (N_14068,N_8661,N_5559);
and U14069 (N_14069,N_6946,N_8949);
xor U14070 (N_14070,N_5175,N_6237);
nor U14071 (N_14071,N_5151,N_8159);
xor U14072 (N_14072,N_6900,N_8214);
nor U14073 (N_14073,N_5329,N_9455);
nand U14074 (N_14074,N_6449,N_8688);
and U14075 (N_14075,N_6009,N_8897);
or U14076 (N_14076,N_8311,N_6635);
and U14077 (N_14077,N_9545,N_9980);
and U14078 (N_14078,N_6010,N_7322);
nand U14079 (N_14079,N_9380,N_8928);
or U14080 (N_14080,N_7278,N_6334);
or U14081 (N_14081,N_5931,N_8476);
xor U14082 (N_14082,N_6618,N_5093);
and U14083 (N_14083,N_6362,N_8808);
nor U14084 (N_14084,N_8167,N_6811);
nand U14085 (N_14085,N_9812,N_5629);
or U14086 (N_14086,N_6937,N_5180);
nand U14087 (N_14087,N_9686,N_8011);
nor U14088 (N_14088,N_7087,N_7324);
and U14089 (N_14089,N_7078,N_9709);
or U14090 (N_14090,N_6847,N_9814);
and U14091 (N_14091,N_7569,N_9833);
nor U14092 (N_14092,N_5348,N_9062);
nor U14093 (N_14093,N_9521,N_9639);
nor U14094 (N_14094,N_7347,N_5671);
or U14095 (N_14095,N_5246,N_7906);
nor U14096 (N_14096,N_5133,N_5149);
and U14097 (N_14097,N_7560,N_7185);
nor U14098 (N_14098,N_5462,N_6588);
nand U14099 (N_14099,N_7210,N_6784);
nor U14100 (N_14100,N_9269,N_5036);
nand U14101 (N_14101,N_6623,N_7059);
or U14102 (N_14102,N_8660,N_5331);
nor U14103 (N_14103,N_9737,N_5612);
nor U14104 (N_14104,N_7100,N_6887);
nand U14105 (N_14105,N_7209,N_5415);
nor U14106 (N_14106,N_5180,N_9286);
and U14107 (N_14107,N_5506,N_7686);
nand U14108 (N_14108,N_7360,N_5865);
nand U14109 (N_14109,N_7253,N_7387);
nor U14110 (N_14110,N_7249,N_9768);
xnor U14111 (N_14111,N_7922,N_6984);
nor U14112 (N_14112,N_9146,N_8221);
nand U14113 (N_14113,N_7352,N_8503);
and U14114 (N_14114,N_7618,N_5483);
nor U14115 (N_14115,N_7411,N_7265);
or U14116 (N_14116,N_9098,N_7427);
or U14117 (N_14117,N_7177,N_8299);
or U14118 (N_14118,N_8629,N_8837);
nand U14119 (N_14119,N_6836,N_9061);
and U14120 (N_14120,N_5824,N_6113);
nor U14121 (N_14121,N_7064,N_9544);
nor U14122 (N_14122,N_9517,N_6293);
nand U14123 (N_14123,N_9781,N_5364);
nand U14124 (N_14124,N_8266,N_7396);
and U14125 (N_14125,N_8869,N_5452);
nor U14126 (N_14126,N_6494,N_5421);
nand U14127 (N_14127,N_7408,N_7434);
nand U14128 (N_14128,N_5911,N_6100);
and U14129 (N_14129,N_6446,N_8720);
xor U14130 (N_14130,N_9118,N_7596);
or U14131 (N_14131,N_8502,N_8659);
nand U14132 (N_14132,N_9444,N_9080);
nand U14133 (N_14133,N_5982,N_5294);
or U14134 (N_14134,N_5375,N_9062);
or U14135 (N_14135,N_5891,N_9020);
or U14136 (N_14136,N_6391,N_6049);
and U14137 (N_14137,N_9085,N_6612);
and U14138 (N_14138,N_5585,N_6452);
nand U14139 (N_14139,N_9520,N_6048);
and U14140 (N_14140,N_8476,N_5554);
and U14141 (N_14141,N_8653,N_7515);
and U14142 (N_14142,N_6014,N_8296);
xor U14143 (N_14143,N_6499,N_7763);
nand U14144 (N_14144,N_8640,N_8737);
and U14145 (N_14145,N_6940,N_5130);
nand U14146 (N_14146,N_8478,N_7895);
nand U14147 (N_14147,N_7951,N_5342);
or U14148 (N_14148,N_5294,N_7889);
nand U14149 (N_14149,N_8990,N_8359);
nand U14150 (N_14150,N_6564,N_6783);
and U14151 (N_14151,N_7879,N_7201);
or U14152 (N_14152,N_7394,N_8373);
nor U14153 (N_14153,N_7820,N_6238);
and U14154 (N_14154,N_8729,N_9021);
nand U14155 (N_14155,N_6332,N_5822);
or U14156 (N_14156,N_5749,N_9970);
or U14157 (N_14157,N_9584,N_8943);
and U14158 (N_14158,N_6692,N_5138);
and U14159 (N_14159,N_9068,N_7718);
or U14160 (N_14160,N_6383,N_7855);
nand U14161 (N_14161,N_8085,N_6383);
nor U14162 (N_14162,N_6525,N_6627);
and U14163 (N_14163,N_5893,N_5614);
nand U14164 (N_14164,N_8842,N_8698);
nand U14165 (N_14165,N_5728,N_8024);
or U14166 (N_14166,N_5656,N_7010);
and U14167 (N_14167,N_7465,N_5312);
or U14168 (N_14168,N_5273,N_9791);
or U14169 (N_14169,N_9839,N_7122);
or U14170 (N_14170,N_6865,N_7181);
nand U14171 (N_14171,N_5132,N_9036);
nor U14172 (N_14172,N_6832,N_6245);
and U14173 (N_14173,N_8106,N_7426);
and U14174 (N_14174,N_6075,N_7594);
or U14175 (N_14175,N_7779,N_6457);
nand U14176 (N_14176,N_5404,N_8052);
and U14177 (N_14177,N_6666,N_9056);
nor U14178 (N_14178,N_7475,N_6044);
or U14179 (N_14179,N_5105,N_8252);
xor U14180 (N_14180,N_5704,N_5791);
or U14181 (N_14181,N_5934,N_7872);
or U14182 (N_14182,N_9503,N_6295);
nor U14183 (N_14183,N_6061,N_6098);
nand U14184 (N_14184,N_9129,N_7639);
or U14185 (N_14185,N_6465,N_7796);
nor U14186 (N_14186,N_9047,N_7113);
nor U14187 (N_14187,N_7437,N_5688);
nor U14188 (N_14188,N_9246,N_7760);
xor U14189 (N_14189,N_7980,N_8454);
or U14190 (N_14190,N_7903,N_6960);
and U14191 (N_14191,N_6604,N_5194);
or U14192 (N_14192,N_7419,N_7663);
or U14193 (N_14193,N_6161,N_9706);
or U14194 (N_14194,N_7236,N_6830);
nor U14195 (N_14195,N_8007,N_7705);
and U14196 (N_14196,N_8420,N_7458);
xnor U14197 (N_14197,N_5673,N_5916);
nand U14198 (N_14198,N_9916,N_6369);
or U14199 (N_14199,N_6631,N_5108);
or U14200 (N_14200,N_9772,N_9959);
nand U14201 (N_14201,N_5639,N_5188);
nand U14202 (N_14202,N_5491,N_9847);
and U14203 (N_14203,N_8699,N_5341);
or U14204 (N_14204,N_7055,N_6864);
nor U14205 (N_14205,N_7625,N_6164);
or U14206 (N_14206,N_7332,N_8166);
or U14207 (N_14207,N_8712,N_8636);
and U14208 (N_14208,N_7496,N_9771);
or U14209 (N_14209,N_6988,N_6421);
or U14210 (N_14210,N_7885,N_5065);
or U14211 (N_14211,N_8055,N_8320);
nor U14212 (N_14212,N_7597,N_9620);
xor U14213 (N_14213,N_9068,N_6749);
or U14214 (N_14214,N_9475,N_8503);
or U14215 (N_14215,N_6015,N_8320);
nand U14216 (N_14216,N_5633,N_9236);
nand U14217 (N_14217,N_9712,N_7815);
or U14218 (N_14218,N_9008,N_9383);
nand U14219 (N_14219,N_5075,N_9824);
and U14220 (N_14220,N_8583,N_5294);
and U14221 (N_14221,N_5590,N_7569);
or U14222 (N_14222,N_6554,N_5971);
nand U14223 (N_14223,N_8555,N_7580);
or U14224 (N_14224,N_8725,N_9522);
and U14225 (N_14225,N_9987,N_9994);
nor U14226 (N_14226,N_7276,N_9703);
nor U14227 (N_14227,N_7200,N_5810);
and U14228 (N_14228,N_6122,N_6843);
xnor U14229 (N_14229,N_8578,N_8979);
and U14230 (N_14230,N_9672,N_6322);
nor U14231 (N_14231,N_8961,N_8770);
xor U14232 (N_14232,N_6751,N_7690);
xor U14233 (N_14233,N_9053,N_5243);
xor U14234 (N_14234,N_6629,N_7273);
nor U14235 (N_14235,N_5946,N_8565);
nand U14236 (N_14236,N_9400,N_5596);
or U14237 (N_14237,N_8410,N_7136);
nor U14238 (N_14238,N_8091,N_8621);
nor U14239 (N_14239,N_7543,N_7033);
or U14240 (N_14240,N_6061,N_9748);
nand U14241 (N_14241,N_5130,N_5383);
and U14242 (N_14242,N_8359,N_7422);
xor U14243 (N_14243,N_8861,N_8621);
nand U14244 (N_14244,N_8361,N_5885);
xor U14245 (N_14245,N_9725,N_9651);
nor U14246 (N_14246,N_9891,N_8678);
nand U14247 (N_14247,N_9429,N_7242);
and U14248 (N_14248,N_6556,N_8030);
and U14249 (N_14249,N_9209,N_9556);
nand U14250 (N_14250,N_5246,N_9251);
and U14251 (N_14251,N_7382,N_8848);
and U14252 (N_14252,N_8721,N_9968);
or U14253 (N_14253,N_8406,N_8833);
and U14254 (N_14254,N_8307,N_9750);
nand U14255 (N_14255,N_5657,N_6645);
or U14256 (N_14256,N_8049,N_5522);
or U14257 (N_14257,N_9656,N_7069);
nor U14258 (N_14258,N_6619,N_8834);
or U14259 (N_14259,N_8434,N_6008);
or U14260 (N_14260,N_8650,N_7056);
or U14261 (N_14261,N_8369,N_7087);
nand U14262 (N_14262,N_7498,N_7777);
and U14263 (N_14263,N_6611,N_6836);
nand U14264 (N_14264,N_8281,N_9723);
nor U14265 (N_14265,N_9961,N_9201);
nor U14266 (N_14266,N_5433,N_9088);
nand U14267 (N_14267,N_7327,N_9553);
xor U14268 (N_14268,N_9813,N_7249);
nor U14269 (N_14269,N_7522,N_7700);
xor U14270 (N_14270,N_9392,N_5251);
nand U14271 (N_14271,N_7707,N_8369);
nor U14272 (N_14272,N_7543,N_8793);
and U14273 (N_14273,N_7332,N_8772);
nand U14274 (N_14274,N_6775,N_7003);
nand U14275 (N_14275,N_8904,N_7815);
nand U14276 (N_14276,N_8726,N_6672);
and U14277 (N_14277,N_7404,N_7645);
nor U14278 (N_14278,N_5636,N_8548);
nand U14279 (N_14279,N_8389,N_5840);
nand U14280 (N_14280,N_8262,N_7190);
and U14281 (N_14281,N_5306,N_9975);
and U14282 (N_14282,N_5718,N_8077);
nor U14283 (N_14283,N_8140,N_5923);
nor U14284 (N_14284,N_8848,N_8130);
or U14285 (N_14285,N_5526,N_5438);
or U14286 (N_14286,N_6254,N_8462);
and U14287 (N_14287,N_8666,N_5450);
nor U14288 (N_14288,N_8896,N_5710);
and U14289 (N_14289,N_8591,N_7063);
nor U14290 (N_14290,N_9596,N_8266);
or U14291 (N_14291,N_8286,N_7000);
nor U14292 (N_14292,N_8615,N_7281);
xor U14293 (N_14293,N_7282,N_5534);
and U14294 (N_14294,N_7410,N_8326);
and U14295 (N_14295,N_7813,N_5421);
xor U14296 (N_14296,N_7408,N_8956);
xnor U14297 (N_14297,N_5101,N_6891);
or U14298 (N_14298,N_5545,N_7228);
nor U14299 (N_14299,N_5230,N_8728);
nand U14300 (N_14300,N_9797,N_7991);
nand U14301 (N_14301,N_7252,N_6393);
or U14302 (N_14302,N_5275,N_6191);
or U14303 (N_14303,N_5685,N_7714);
and U14304 (N_14304,N_5609,N_7213);
or U14305 (N_14305,N_5724,N_7898);
or U14306 (N_14306,N_9225,N_9743);
xnor U14307 (N_14307,N_8386,N_9034);
or U14308 (N_14308,N_9551,N_6532);
and U14309 (N_14309,N_9584,N_9641);
and U14310 (N_14310,N_6587,N_5796);
and U14311 (N_14311,N_6589,N_8926);
and U14312 (N_14312,N_5061,N_6277);
nor U14313 (N_14313,N_5950,N_6978);
and U14314 (N_14314,N_5169,N_9007);
xor U14315 (N_14315,N_6952,N_8676);
or U14316 (N_14316,N_6218,N_6716);
and U14317 (N_14317,N_5154,N_7103);
or U14318 (N_14318,N_6009,N_8577);
and U14319 (N_14319,N_6095,N_6069);
nor U14320 (N_14320,N_9205,N_5282);
or U14321 (N_14321,N_8991,N_8517);
or U14322 (N_14322,N_6140,N_9508);
or U14323 (N_14323,N_9533,N_9327);
nor U14324 (N_14324,N_7232,N_9118);
nand U14325 (N_14325,N_9383,N_7967);
nor U14326 (N_14326,N_8669,N_6499);
or U14327 (N_14327,N_5722,N_8550);
and U14328 (N_14328,N_5677,N_7265);
or U14329 (N_14329,N_8591,N_8270);
or U14330 (N_14330,N_7466,N_9831);
nand U14331 (N_14331,N_5337,N_6663);
xor U14332 (N_14332,N_6253,N_5480);
and U14333 (N_14333,N_9006,N_7210);
nand U14334 (N_14334,N_8999,N_5953);
or U14335 (N_14335,N_9451,N_6593);
or U14336 (N_14336,N_8769,N_6836);
and U14337 (N_14337,N_6185,N_9043);
nand U14338 (N_14338,N_6668,N_9860);
or U14339 (N_14339,N_5685,N_7891);
and U14340 (N_14340,N_8140,N_7593);
or U14341 (N_14341,N_5819,N_7882);
or U14342 (N_14342,N_7688,N_6354);
nor U14343 (N_14343,N_5144,N_5686);
and U14344 (N_14344,N_5795,N_6490);
xnor U14345 (N_14345,N_8120,N_7582);
nor U14346 (N_14346,N_8461,N_8323);
or U14347 (N_14347,N_6963,N_6331);
nor U14348 (N_14348,N_9785,N_7333);
xor U14349 (N_14349,N_7971,N_8722);
nor U14350 (N_14350,N_5767,N_6490);
nor U14351 (N_14351,N_9536,N_5813);
nand U14352 (N_14352,N_8070,N_6599);
and U14353 (N_14353,N_9910,N_7191);
or U14354 (N_14354,N_8193,N_5902);
and U14355 (N_14355,N_5129,N_6596);
and U14356 (N_14356,N_9747,N_9405);
nand U14357 (N_14357,N_5169,N_7784);
and U14358 (N_14358,N_5105,N_6045);
xor U14359 (N_14359,N_8040,N_9709);
or U14360 (N_14360,N_9807,N_6692);
or U14361 (N_14361,N_5028,N_5662);
or U14362 (N_14362,N_6841,N_6152);
xnor U14363 (N_14363,N_6977,N_5135);
and U14364 (N_14364,N_6722,N_6491);
or U14365 (N_14365,N_7224,N_6440);
and U14366 (N_14366,N_6284,N_6358);
nor U14367 (N_14367,N_7232,N_7163);
nand U14368 (N_14368,N_5056,N_6375);
and U14369 (N_14369,N_9512,N_5405);
or U14370 (N_14370,N_8199,N_5735);
nand U14371 (N_14371,N_6526,N_7102);
nand U14372 (N_14372,N_7732,N_5710);
nand U14373 (N_14373,N_9396,N_9823);
or U14374 (N_14374,N_5734,N_7128);
or U14375 (N_14375,N_7702,N_6300);
nor U14376 (N_14376,N_8527,N_9964);
nor U14377 (N_14377,N_9719,N_7122);
and U14378 (N_14378,N_9875,N_5635);
or U14379 (N_14379,N_7284,N_8233);
xor U14380 (N_14380,N_5622,N_6916);
xor U14381 (N_14381,N_8353,N_9061);
and U14382 (N_14382,N_6434,N_5477);
nor U14383 (N_14383,N_6468,N_5179);
or U14384 (N_14384,N_6534,N_9656);
nor U14385 (N_14385,N_5105,N_5903);
or U14386 (N_14386,N_5592,N_9179);
nor U14387 (N_14387,N_9490,N_5575);
nor U14388 (N_14388,N_7043,N_6632);
or U14389 (N_14389,N_5918,N_7579);
or U14390 (N_14390,N_7921,N_8163);
nand U14391 (N_14391,N_8336,N_5110);
nor U14392 (N_14392,N_9312,N_5118);
nand U14393 (N_14393,N_8196,N_6892);
nand U14394 (N_14394,N_8574,N_5352);
nor U14395 (N_14395,N_5299,N_7071);
nor U14396 (N_14396,N_5589,N_9646);
nor U14397 (N_14397,N_8403,N_6632);
and U14398 (N_14398,N_9984,N_8202);
nand U14399 (N_14399,N_5470,N_6431);
xor U14400 (N_14400,N_9098,N_5402);
or U14401 (N_14401,N_5240,N_6284);
nand U14402 (N_14402,N_8422,N_9526);
nand U14403 (N_14403,N_6692,N_9477);
and U14404 (N_14404,N_6952,N_7145);
and U14405 (N_14405,N_7793,N_8588);
and U14406 (N_14406,N_7870,N_5621);
nor U14407 (N_14407,N_8460,N_6755);
xor U14408 (N_14408,N_5691,N_8749);
or U14409 (N_14409,N_6038,N_8019);
nand U14410 (N_14410,N_6333,N_5116);
and U14411 (N_14411,N_8261,N_6256);
or U14412 (N_14412,N_8795,N_9813);
nand U14413 (N_14413,N_6215,N_7984);
nor U14414 (N_14414,N_7062,N_9939);
or U14415 (N_14415,N_7681,N_9658);
nand U14416 (N_14416,N_6921,N_6048);
nor U14417 (N_14417,N_9970,N_9250);
nand U14418 (N_14418,N_5586,N_7015);
or U14419 (N_14419,N_5260,N_7400);
nor U14420 (N_14420,N_6124,N_7835);
or U14421 (N_14421,N_7234,N_9072);
nand U14422 (N_14422,N_5709,N_7881);
and U14423 (N_14423,N_6774,N_8429);
and U14424 (N_14424,N_9926,N_8778);
or U14425 (N_14425,N_5054,N_8910);
or U14426 (N_14426,N_7084,N_6024);
or U14427 (N_14427,N_9956,N_6846);
nand U14428 (N_14428,N_9438,N_9383);
and U14429 (N_14429,N_5702,N_8501);
and U14430 (N_14430,N_9931,N_9359);
nor U14431 (N_14431,N_7207,N_8410);
nor U14432 (N_14432,N_6330,N_9260);
or U14433 (N_14433,N_8224,N_6598);
and U14434 (N_14434,N_9037,N_6094);
and U14435 (N_14435,N_6519,N_7870);
nor U14436 (N_14436,N_7419,N_5875);
and U14437 (N_14437,N_5388,N_7069);
nor U14438 (N_14438,N_7675,N_5234);
nor U14439 (N_14439,N_6898,N_8294);
or U14440 (N_14440,N_6621,N_5625);
and U14441 (N_14441,N_7625,N_8538);
and U14442 (N_14442,N_7770,N_8746);
or U14443 (N_14443,N_8072,N_9085);
xor U14444 (N_14444,N_5525,N_7095);
nand U14445 (N_14445,N_8364,N_9582);
or U14446 (N_14446,N_6144,N_9953);
nand U14447 (N_14447,N_5300,N_6893);
nor U14448 (N_14448,N_6758,N_8736);
and U14449 (N_14449,N_9511,N_6171);
and U14450 (N_14450,N_8928,N_8864);
nor U14451 (N_14451,N_5821,N_5021);
and U14452 (N_14452,N_9824,N_6447);
or U14453 (N_14453,N_5193,N_5139);
and U14454 (N_14454,N_5283,N_7470);
or U14455 (N_14455,N_8921,N_5245);
or U14456 (N_14456,N_5782,N_7543);
or U14457 (N_14457,N_6110,N_8784);
nor U14458 (N_14458,N_7251,N_8973);
and U14459 (N_14459,N_6128,N_9919);
or U14460 (N_14460,N_6730,N_6614);
xor U14461 (N_14461,N_9464,N_8264);
and U14462 (N_14462,N_5360,N_7189);
or U14463 (N_14463,N_9268,N_8456);
or U14464 (N_14464,N_7578,N_5375);
nand U14465 (N_14465,N_8516,N_7813);
or U14466 (N_14466,N_8665,N_7067);
or U14467 (N_14467,N_8270,N_9109);
nand U14468 (N_14468,N_7831,N_5111);
xor U14469 (N_14469,N_7653,N_8143);
nand U14470 (N_14470,N_6878,N_7548);
nand U14471 (N_14471,N_9657,N_7458);
and U14472 (N_14472,N_6080,N_8091);
and U14473 (N_14473,N_5875,N_5934);
nor U14474 (N_14474,N_6028,N_7402);
or U14475 (N_14475,N_9690,N_8286);
nand U14476 (N_14476,N_5297,N_5788);
nor U14477 (N_14477,N_5419,N_9691);
and U14478 (N_14478,N_9597,N_9659);
xor U14479 (N_14479,N_7590,N_6277);
and U14480 (N_14480,N_8285,N_5376);
or U14481 (N_14481,N_9111,N_9586);
and U14482 (N_14482,N_7305,N_6328);
nor U14483 (N_14483,N_7401,N_6169);
nor U14484 (N_14484,N_8940,N_6770);
nor U14485 (N_14485,N_6316,N_5865);
nor U14486 (N_14486,N_8127,N_8446);
and U14487 (N_14487,N_9675,N_7728);
and U14488 (N_14488,N_6554,N_6621);
nor U14489 (N_14489,N_7246,N_9907);
or U14490 (N_14490,N_5542,N_9348);
nor U14491 (N_14491,N_7884,N_6105);
and U14492 (N_14492,N_5511,N_6503);
and U14493 (N_14493,N_6527,N_8863);
and U14494 (N_14494,N_9415,N_5908);
or U14495 (N_14495,N_7981,N_9440);
or U14496 (N_14496,N_8785,N_9076);
nand U14497 (N_14497,N_5392,N_6006);
and U14498 (N_14498,N_9273,N_5704);
nor U14499 (N_14499,N_7150,N_9972);
and U14500 (N_14500,N_6241,N_7785);
or U14501 (N_14501,N_9699,N_9174);
and U14502 (N_14502,N_8996,N_6211);
or U14503 (N_14503,N_8315,N_7881);
and U14504 (N_14504,N_8083,N_9729);
nor U14505 (N_14505,N_8702,N_6129);
and U14506 (N_14506,N_9802,N_5467);
nand U14507 (N_14507,N_5645,N_7186);
xnor U14508 (N_14508,N_9571,N_8655);
or U14509 (N_14509,N_6646,N_9248);
xnor U14510 (N_14510,N_8992,N_8358);
nor U14511 (N_14511,N_7427,N_8581);
and U14512 (N_14512,N_8198,N_7279);
nor U14513 (N_14513,N_8652,N_8175);
or U14514 (N_14514,N_6670,N_6237);
nor U14515 (N_14515,N_9800,N_6190);
or U14516 (N_14516,N_5939,N_6837);
xnor U14517 (N_14517,N_6248,N_8354);
xor U14518 (N_14518,N_9962,N_9855);
nand U14519 (N_14519,N_9446,N_8019);
or U14520 (N_14520,N_5737,N_8756);
and U14521 (N_14521,N_9401,N_7401);
nand U14522 (N_14522,N_6057,N_7660);
nand U14523 (N_14523,N_7534,N_7300);
nor U14524 (N_14524,N_5900,N_7180);
or U14525 (N_14525,N_6753,N_9860);
nor U14526 (N_14526,N_6594,N_7819);
and U14527 (N_14527,N_8602,N_5683);
nor U14528 (N_14528,N_6807,N_6193);
nand U14529 (N_14529,N_8037,N_5512);
or U14530 (N_14530,N_5495,N_9199);
nand U14531 (N_14531,N_6588,N_6394);
or U14532 (N_14532,N_5660,N_6767);
and U14533 (N_14533,N_5970,N_9925);
and U14534 (N_14534,N_9703,N_5733);
nor U14535 (N_14535,N_5937,N_9766);
nor U14536 (N_14536,N_9491,N_7816);
nand U14537 (N_14537,N_6123,N_5881);
nand U14538 (N_14538,N_5679,N_7982);
nor U14539 (N_14539,N_8931,N_7490);
nor U14540 (N_14540,N_7878,N_6917);
and U14541 (N_14541,N_7689,N_9353);
or U14542 (N_14542,N_8658,N_9961);
nand U14543 (N_14543,N_9994,N_7216);
and U14544 (N_14544,N_8531,N_8966);
or U14545 (N_14545,N_5119,N_5734);
nand U14546 (N_14546,N_6847,N_7384);
and U14547 (N_14547,N_5068,N_6056);
nand U14548 (N_14548,N_7483,N_7060);
or U14549 (N_14549,N_7387,N_7866);
and U14550 (N_14550,N_5286,N_5279);
and U14551 (N_14551,N_9339,N_7716);
and U14552 (N_14552,N_5281,N_5271);
xor U14553 (N_14553,N_7195,N_5685);
nand U14554 (N_14554,N_6591,N_5227);
or U14555 (N_14555,N_6397,N_6025);
and U14556 (N_14556,N_5444,N_6130);
xnor U14557 (N_14557,N_9069,N_6878);
or U14558 (N_14558,N_7973,N_5195);
nor U14559 (N_14559,N_8549,N_8188);
and U14560 (N_14560,N_7199,N_7214);
or U14561 (N_14561,N_7584,N_8527);
or U14562 (N_14562,N_6684,N_8562);
and U14563 (N_14563,N_7910,N_6938);
and U14564 (N_14564,N_9578,N_8246);
or U14565 (N_14565,N_8888,N_7068);
and U14566 (N_14566,N_5763,N_7288);
nand U14567 (N_14567,N_6371,N_8798);
nand U14568 (N_14568,N_6021,N_6432);
and U14569 (N_14569,N_6994,N_8119);
or U14570 (N_14570,N_5136,N_8941);
and U14571 (N_14571,N_5834,N_6787);
nor U14572 (N_14572,N_9550,N_7576);
or U14573 (N_14573,N_7370,N_8558);
and U14574 (N_14574,N_8436,N_8408);
or U14575 (N_14575,N_8638,N_7850);
nor U14576 (N_14576,N_5600,N_7569);
nand U14577 (N_14577,N_5198,N_9254);
or U14578 (N_14578,N_8835,N_7657);
nor U14579 (N_14579,N_7026,N_9202);
or U14580 (N_14580,N_5464,N_9988);
xnor U14581 (N_14581,N_5546,N_5793);
and U14582 (N_14582,N_9651,N_8773);
nor U14583 (N_14583,N_8990,N_6979);
and U14584 (N_14584,N_6829,N_6211);
nor U14585 (N_14585,N_9232,N_5256);
nor U14586 (N_14586,N_9035,N_8547);
or U14587 (N_14587,N_9247,N_8280);
or U14588 (N_14588,N_7569,N_6315);
xnor U14589 (N_14589,N_8846,N_6809);
nor U14590 (N_14590,N_6087,N_9834);
xor U14591 (N_14591,N_6838,N_5819);
nor U14592 (N_14592,N_6181,N_9431);
nand U14593 (N_14593,N_5959,N_9505);
or U14594 (N_14594,N_5423,N_5210);
and U14595 (N_14595,N_5765,N_6926);
nor U14596 (N_14596,N_5084,N_6129);
nor U14597 (N_14597,N_6034,N_8701);
xnor U14598 (N_14598,N_7547,N_5744);
or U14599 (N_14599,N_5248,N_5294);
nand U14600 (N_14600,N_8130,N_8969);
nand U14601 (N_14601,N_6038,N_5782);
or U14602 (N_14602,N_6103,N_7477);
and U14603 (N_14603,N_6621,N_5765);
nor U14604 (N_14604,N_5299,N_7584);
and U14605 (N_14605,N_6089,N_7846);
nor U14606 (N_14606,N_6939,N_8537);
xor U14607 (N_14607,N_9116,N_7714);
xor U14608 (N_14608,N_5781,N_8423);
or U14609 (N_14609,N_6481,N_7509);
xnor U14610 (N_14610,N_9860,N_8035);
xnor U14611 (N_14611,N_8997,N_9750);
nor U14612 (N_14612,N_9870,N_7882);
nor U14613 (N_14613,N_9136,N_7186);
xnor U14614 (N_14614,N_6002,N_5760);
and U14615 (N_14615,N_8236,N_8927);
and U14616 (N_14616,N_6677,N_8345);
or U14617 (N_14617,N_7355,N_8177);
nand U14618 (N_14618,N_7814,N_7733);
nor U14619 (N_14619,N_5687,N_7129);
or U14620 (N_14620,N_5327,N_9487);
and U14621 (N_14621,N_6325,N_6187);
and U14622 (N_14622,N_5742,N_6425);
xor U14623 (N_14623,N_7599,N_9038);
nand U14624 (N_14624,N_5948,N_7097);
or U14625 (N_14625,N_7855,N_9407);
nor U14626 (N_14626,N_7681,N_5320);
nand U14627 (N_14627,N_7757,N_7643);
or U14628 (N_14628,N_7315,N_5423);
nand U14629 (N_14629,N_6124,N_8310);
nand U14630 (N_14630,N_7180,N_5807);
nor U14631 (N_14631,N_9762,N_9348);
or U14632 (N_14632,N_9535,N_8751);
or U14633 (N_14633,N_6455,N_8125);
and U14634 (N_14634,N_6512,N_6857);
xor U14635 (N_14635,N_9894,N_6583);
or U14636 (N_14636,N_5612,N_7505);
nor U14637 (N_14637,N_9376,N_8311);
or U14638 (N_14638,N_5659,N_5362);
nor U14639 (N_14639,N_9595,N_5436);
and U14640 (N_14640,N_6948,N_6175);
or U14641 (N_14641,N_7978,N_6466);
nor U14642 (N_14642,N_8985,N_9740);
or U14643 (N_14643,N_8019,N_7845);
xnor U14644 (N_14644,N_6746,N_7955);
or U14645 (N_14645,N_5114,N_8524);
nand U14646 (N_14646,N_9199,N_8150);
nor U14647 (N_14647,N_7278,N_8786);
nor U14648 (N_14648,N_5257,N_9001);
and U14649 (N_14649,N_7081,N_9968);
and U14650 (N_14650,N_7099,N_6241);
or U14651 (N_14651,N_7424,N_9900);
and U14652 (N_14652,N_9900,N_9901);
nand U14653 (N_14653,N_6981,N_5622);
nand U14654 (N_14654,N_5020,N_6438);
nor U14655 (N_14655,N_9289,N_6019);
nand U14656 (N_14656,N_5852,N_7501);
nor U14657 (N_14657,N_5793,N_9492);
or U14658 (N_14658,N_9350,N_5242);
or U14659 (N_14659,N_8618,N_9985);
nand U14660 (N_14660,N_6460,N_9743);
nand U14661 (N_14661,N_6859,N_7532);
nand U14662 (N_14662,N_8443,N_6352);
or U14663 (N_14663,N_5021,N_8052);
and U14664 (N_14664,N_6274,N_7292);
or U14665 (N_14665,N_6447,N_5512);
nor U14666 (N_14666,N_7689,N_6766);
nor U14667 (N_14667,N_9825,N_5905);
nand U14668 (N_14668,N_9975,N_8563);
nand U14669 (N_14669,N_8991,N_5120);
nand U14670 (N_14670,N_5677,N_9472);
nand U14671 (N_14671,N_7415,N_5310);
and U14672 (N_14672,N_9660,N_9895);
and U14673 (N_14673,N_6204,N_6134);
nor U14674 (N_14674,N_5263,N_8234);
xnor U14675 (N_14675,N_5660,N_7640);
nor U14676 (N_14676,N_8262,N_5931);
nand U14677 (N_14677,N_7197,N_6443);
and U14678 (N_14678,N_9213,N_8124);
and U14679 (N_14679,N_9730,N_5208);
and U14680 (N_14680,N_7939,N_9441);
and U14681 (N_14681,N_8623,N_9774);
nor U14682 (N_14682,N_6571,N_8084);
or U14683 (N_14683,N_9130,N_6203);
nand U14684 (N_14684,N_5637,N_5722);
or U14685 (N_14685,N_8334,N_9842);
or U14686 (N_14686,N_7323,N_7489);
and U14687 (N_14687,N_8138,N_8716);
nand U14688 (N_14688,N_6759,N_8737);
or U14689 (N_14689,N_7674,N_9993);
xor U14690 (N_14690,N_8890,N_5738);
and U14691 (N_14691,N_9129,N_9122);
nor U14692 (N_14692,N_5807,N_7941);
or U14693 (N_14693,N_5197,N_5744);
and U14694 (N_14694,N_5201,N_5192);
nor U14695 (N_14695,N_5062,N_8733);
nand U14696 (N_14696,N_9017,N_8974);
nand U14697 (N_14697,N_5689,N_8864);
and U14698 (N_14698,N_5458,N_5737);
nor U14699 (N_14699,N_5389,N_8231);
and U14700 (N_14700,N_6677,N_9614);
nor U14701 (N_14701,N_7700,N_8537);
nor U14702 (N_14702,N_6739,N_9182);
nand U14703 (N_14703,N_6935,N_9812);
nor U14704 (N_14704,N_9695,N_8149);
nand U14705 (N_14705,N_5422,N_6856);
nor U14706 (N_14706,N_9290,N_7324);
nand U14707 (N_14707,N_9431,N_8937);
nor U14708 (N_14708,N_8455,N_8826);
nor U14709 (N_14709,N_5782,N_7441);
and U14710 (N_14710,N_7733,N_5835);
or U14711 (N_14711,N_5411,N_5122);
xnor U14712 (N_14712,N_5537,N_8048);
and U14713 (N_14713,N_8188,N_5615);
nor U14714 (N_14714,N_9142,N_6525);
nand U14715 (N_14715,N_6542,N_8370);
nor U14716 (N_14716,N_7694,N_9903);
or U14717 (N_14717,N_8404,N_8647);
xnor U14718 (N_14718,N_7691,N_9162);
nand U14719 (N_14719,N_5340,N_8206);
and U14720 (N_14720,N_9770,N_5621);
nor U14721 (N_14721,N_8129,N_8603);
nor U14722 (N_14722,N_5483,N_6841);
nand U14723 (N_14723,N_8576,N_8437);
nand U14724 (N_14724,N_8443,N_9303);
nand U14725 (N_14725,N_9200,N_8226);
nand U14726 (N_14726,N_6987,N_6483);
nand U14727 (N_14727,N_5752,N_9465);
or U14728 (N_14728,N_5230,N_7804);
and U14729 (N_14729,N_5582,N_9731);
nand U14730 (N_14730,N_5418,N_5611);
nor U14731 (N_14731,N_9041,N_6685);
nand U14732 (N_14732,N_8673,N_9356);
or U14733 (N_14733,N_7196,N_8648);
and U14734 (N_14734,N_7309,N_7847);
nor U14735 (N_14735,N_7337,N_9048);
and U14736 (N_14736,N_8145,N_9853);
nand U14737 (N_14737,N_8601,N_6340);
nand U14738 (N_14738,N_5634,N_6451);
nor U14739 (N_14739,N_9542,N_9719);
nor U14740 (N_14740,N_7434,N_6438);
nor U14741 (N_14741,N_6232,N_9092);
nor U14742 (N_14742,N_9003,N_7016);
or U14743 (N_14743,N_6571,N_5375);
nand U14744 (N_14744,N_8220,N_9977);
nor U14745 (N_14745,N_6177,N_6501);
or U14746 (N_14746,N_5308,N_6611);
and U14747 (N_14747,N_8082,N_7688);
nor U14748 (N_14748,N_6531,N_5811);
or U14749 (N_14749,N_8104,N_6614);
nand U14750 (N_14750,N_8155,N_8275);
and U14751 (N_14751,N_9449,N_9486);
or U14752 (N_14752,N_6101,N_7678);
or U14753 (N_14753,N_8685,N_9688);
nand U14754 (N_14754,N_9138,N_5887);
and U14755 (N_14755,N_6646,N_9154);
or U14756 (N_14756,N_6210,N_9743);
and U14757 (N_14757,N_7995,N_5175);
or U14758 (N_14758,N_7823,N_9050);
or U14759 (N_14759,N_6749,N_9376);
or U14760 (N_14760,N_7528,N_6651);
nand U14761 (N_14761,N_9965,N_7523);
and U14762 (N_14762,N_8331,N_6275);
nor U14763 (N_14763,N_9086,N_6717);
nor U14764 (N_14764,N_8901,N_8989);
nand U14765 (N_14765,N_5016,N_5286);
and U14766 (N_14766,N_8842,N_8433);
and U14767 (N_14767,N_8025,N_5072);
nand U14768 (N_14768,N_7434,N_6538);
nor U14769 (N_14769,N_9781,N_7610);
and U14770 (N_14770,N_5318,N_6411);
nor U14771 (N_14771,N_7920,N_7141);
xnor U14772 (N_14772,N_8609,N_9192);
or U14773 (N_14773,N_8427,N_6918);
nand U14774 (N_14774,N_6821,N_7094);
and U14775 (N_14775,N_8421,N_7540);
or U14776 (N_14776,N_6573,N_8174);
xnor U14777 (N_14777,N_5564,N_6329);
and U14778 (N_14778,N_7097,N_5899);
or U14779 (N_14779,N_7026,N_9620);
nor U14780 (N_14780,N_8005,N_9854);
or U14781 (N_14781,N_5324,N_6015);
and U14782 (N_14782,N_9110,N_5519);
and U14783 (N_14783,N_8914,N_7688);
xnor U14784 (N_14784,N_7395,N_5495);
and U14785 (N_14785,N_8452,N_6453);
and U14786 (N_14786,N_5394,N_5868);
or U14787 (N_14787,N_8284,N_6634);
nand U14788 (N_14788,N_7973,N_5867);
nor U14789 (N_14789,N_6531,N_7383);
or U14790 (N_14790,N_5996,N_5444);
and U14791 (N_14791,N_7546,N_9798);
nor U14792 (N_14792,N_6250,N_5940);
or U14793 (N_14793,N_8045,N_7061);
or U14794 (N_14794,N_6530,N_9271);
or U14795 (N_14795,N_8095,N_7592);
nand U14796 (N_14796,N_7158,N_5156);
nand U14797 (N_14797,N_9507,N_8517);
nand U14798 (N_14798,N_8112,N_8687);
nor U14799 (N_14799,N_8099,N_6949);
nand U14800 (N_14800,N_8174,N_7559);
xnor U14801 (N_14801,N_9630,N_6607);
and U14802 (N_14802,N_5277,N_8743);
xnor U14803 (N_14803,N_9657,N_7771);
and U14804 (N_14804,N_6387,N_5791);
nand U14805 (N_14805,N_7647,N_9253);
nand U14806 (N_14806,N_6653,N_8095);
and U14807 (N_14807,N_9651,N_5515);
or U14808 (N_14808,N_6250,N_5757);
or U14809 (N_14809,N_6436,N_5073);
nor U14810 (N_14810,N_7087,N_5341);
nor U14811 (N_14811,N_8072,N_5389);
and U14812 (N_14812,N_9336,N_6352);
and U14813 (N_14813,N_8766,N_5291);
and U14814 (N_14814,N_7009,N_5112);
and U14815 (N_14815,N_7997,N_8701);
nor U14816 (N_14816,N_9639,N_8474);
and U14817 (N_14817,N_5045,N_5373);
and U14818 (N_14818,N_8553,N_5390);
and U14819 (N_14819,N_9123,N_8238);
or U14820 (N_14820,N_8454,N_9855);
and U14821 (N_14821,N_6331,N_5742);
nor U14822 (N_14822,N_8072,N_5630);
or U14823 (N_14823,N_7346,N_9691);
and U14824 (N_14824,N_6714,N_9298);
nand U14825 (N_14825,N_8963,N_9174);
and U14826 (N_14826,N_8950,N_7594);
or U14827 (N_14827,N_8157,N_8753);
nor U14828 (N_14828,N_8597,N_8253);
and U14829 (N_14829,N_9637,N_8828);
nor U14830 (N_14830,N_5367,N_6302);
and U14831 (N_14831,N_5565,N_6511);
or U14832 (N_14832,N_6270,N_5062);
nor U14833 (N_14833,N_9796,N_5047);
nand U14834 (N_14834,N_5237,N_8826);
or U14835 (N_14835,N_6682,N_9047);
and U14836 (N_14836,N_8299,N_8767);
or U14837 (N_14837,N_5621,N_9019);
nand U14838 (N_14838,N_7007,N_5250);
or U14839 (N_14839,N_6888,N_7452);
nor U14840 (N_14840,N_6467,N_9950);
xor U14841 (N_14841,N_9577,N_5385);
xnor U14842 (N_14842,N_5957,N_6427);
nor U14843 (N_14843,N_9384,N_5063);
or U14844 (N_14844,N_9663,N_9590);
or U14845 (N_14845,N_8532,N_5338);
or U14846 (N_14846,N_8395,N_9046);
nor U14847 (N_14847,N_9257,N_7649);
nor U14848 (N_14848,N_8402,N_9949);
nor U14849 (N_14849,N_5761,N_9477);
or U14850 (N_14850,N_7580,N_6814);
xor U14851 (N_14851,N_8572,N_6545);
nor U14852 (N_14852,N_8051,N_5888);
nor U14853 (N_14853,N_8375,N_5814);
or U14854 (N_14854,N_8354,N_5460);
nor U14855 (N_14855,N_5891,N_6543);
and U14856 (N_14856,N_6578,N_7231);
nor U14857 (N_14857,N_9254,N_6554);
nor U14858 (N_14858,N_5732,N_8960);
and U14859 (N_14859,N_8548,N_9739);
or U14860 (N_14860,N_6636,N_6736);
or U14861 (N_14861,N_7614,N_7080);
or U14862 (N_14862,N_9618,N_5635);
nand U14863 (N_14863,N_6459,N_6014);
nor U14864 (N_14864,N_6790,N_8461);
or U14865 (N_14865,N_9201,N_8839);
nand U14866 (N_14866,N_8721,N_6943);
and U14867 (N_14867,N_6026,N_5962);
nand U14868 (N_14868,N_6993,N_7480);
and U14869 (N_14869,N_5597,N_5327);
or U14870 (N_14870,N_6383,N_5743);
or U14871 (N_14871,N_9122,N_9528);
and U14872 (N_14872,N_7652,N_6188);
and U14873 (N_14873,N_6147,N_5121);
or U14874 (N_14874,N_7117,N_6449);
nand U14875 (N_14875,N_9333,N_7751);
or U14876 (N_14876,N_8535,N_6627);
nand U14877 (N_14877,N_5959,N_6654);
nand U14878 (N_14878,N_8111,N_7981);
nand U14879 (N_14879,N_9078,N_6500);
nor U14880 (N_14880,N_7444,N_7534);
xor U14881 (N_14881,N_8272,N_7723);
or U14882 (N_14882,N_7512,N_7642);
nor U14883 (N_14883,N_8255,N_9786);
xnor U14884 (N_14884,N_7771,N_5195);
and U14885 (N_14885,N_7539,N_8012);
nor U14886 (N_14886,N_8057,N_7122);
nor U14887 (N_14887,N_6911,N_5631);
or U14888 (N_14888,N_5430,N_5053);
nand U14889 (N_14889,N_9524,N_8734);
nand U14890 (N_14890,N_7977,N_8575);
nand U14891 (N_14891,N_6531,N_9969);
nand U14892 (N_14892,N_9660,N_6890);
nand U14893 (N_14893,N_5102,N_6745);
nor U14894 (N_14894,N_7958,N_9270);
nor U14895 (N_14895,N_6032,N_9275);
nor U14896 (N_14896,N_7563,N_7564);
nand U14897 (N_14897,N_8432,N_6780);
nand U14898 (N_14898,N_7398,N_7438);
nor U14899 (N_14899,N_5843,N_9904);
and U14900 (N_14900,N_5779,N_5038);
or U14901 (N_14901,N_9387,N_5569);
and U14902 (N_14902,N_5270,N_6615);
nand U14903 (N_14903,N_5850,N_5152);
and U14904 (N_14904,N_9943,N_7559);
xnor U14905 (N_14905,N_8394,N_8402);
nor U14906 (N_14906,N_6007,N_5570);
nor U14907 (N_14907,N_5549,N_7188);
nor U14908 (N_14908,N_8420,N_7386);
or U14909 (N_14909,N_6035,N_9371);
and U14910 (N_14910,N_8448,N_6862);
or U14911 (N_14911,N_8625,N_9789);
and U14912 (N_14912,N_5740,N_6202);
or U14913 (N_14913,N_8238,N_8150);
or U14914 (N_14914,N_6567,N_7922);
nand U14915 (N_14915,N_6504,N_5425);
nand U14916 (N_14916,N_7948,N_9509);
and U14917 (N_14917,N_8597,N_7481);
xor U14918 (N_14918,N_7791,N_6126);
or U14919 (N_14919,N_7684,N_7017);
nor U14920 (N_14920,N_7828,N_9246);
nand U14921 (N_14921,N_5638,N_8536);
nand U14922 (N_14922,N_9182,N_5277);
nand U14923 (N_14923,N_6022,N_8222);
xor U14924 (N_14924,N_7752,N_6828);
nand U14925 (N_14925,N_7124,N_8201);
and U14926 (N_14926,N_6350,N_5304);
xor U14927 (N_14927,N_9495,N_5819);
nor U14928 (N_14928,N_7638,N_9336);
or U14929 (N_14929,N_6618,N_7817);
and U14930 (N_14930,N_7094,N_7282);
or U14931 (N_14931,N_9766,N_6540);
and U14932 (N_14932,N_8051,N_7822);
nand U14933 (N_14933,N_7372,N_7319);
nand U14934 (N_14934,N_6365,N_8883);
nand U14935 (N_14935,N_7822,N_5936);
nor U14936 (N_14936,N_9907,N_6116);
nor U14937 (N_14937,N_6228,N_9809);
or U14938 (N_14938,N_8714,N_7146);
or U14939 (N_14939,N_5399,N_8579);
and U14940 (N_14940,N_9224,N_9819);
nor U14941 (N_14941,N_7646,N_6194);
or U14942 (N_14942,N_6966,N_5612);
and U14943 (N_14943,N_8981,N_7702);
or U14944 (N_14944,N_5940,N_5865);
nand U14945 (N_14945,N_8667,N_6966);
and U14946 (N_14946,N_5866,N_7908);
xor U14947 (N_14947,N_9751,N_5641);
nand U14948 (N_14948,N_8255,N_9498);
nor U14949 (N_14949,N_6164,N_8372);
and U14950 (N_14950,N_6684,N_5635);
nor U14951 (N_14951,N_8966,N_6381);
and U14952 (N_14952,N_7700,N_7574);
or U14953 (N_14953,N_7852,N_5449);
nand U14954 (N_14954,N_7318,N_9882);
nor U14955 (N_14955,N_5942,N_7839);
or U14956 (N_14956,N_7174,N_6338);
nand U14957 (N_14957,N_8104,N_9078);
and U14958 (N_14958,N_9310,N_6437);
nor U14959 (N_14959,N_7940,N_8175);
nand U14960 (N_14960,N_8722,N_9343);
nor U14961 (N_14961,N_5816,N_8854);
nor U14962 (N_14962,N_5122,N_6740);
and U14963 (N_14963,N_8266,N_5146);
nor U14964 (N_14964,N_8332,N_9309);
nor U14965 (N_14965,N_6118,N_6468);
xor U14966 (N_14966,N_8671,N_9845);
nand U14967 (N_14967,N_6356,N_5588);
xor U14968 (N_14968,N_7417,N_7292);
or U14969 (N_14969,N_9724,N_8386);
nor U14970 (N_14970,N_9971,N_9619);
and U14971 (N_14971,N_9830,N_9036);
and U14972 (N_14972,N_5776,N_8980);
nor U14973 (N_14973,N_9389,N_8226);
and U14974 (N_14974,N_9195,N_8997);
or U14975 (N_14975,N_5057,N_7927);
nand U14976 (N_14976,N_5396,N_6373);
or U14977 (N_14977,N_7450,N_5441);
nor U14978 (N_14978,N_5438,N_6662);
nand U14979 (N_14979,N_8248,N_6619);
nand U14980 (N_14980,N_9321,N_6900);
xnor U14981 (N_14981,N_7910,N_6975);
nand U14982 (N_14982,N_7671,N_5367);
xor U14983 (N_14983,N_9913,N_9880);
nor U14984 (N_14984,N_6875,N_8244);
or U14985 (N_14985,N_7544,N_6195);
nor U14986 (N_14986,N_6042,N_5606);
nor U14987 (N_14987,N_8642,N_7673);
and U14988 (N_14988,N_8726,N_6627);
and U14989 (N_14989,N_7460,N_7983);
xnor U14990 (N_14990,N_8588,N_5037);
nor U14991 (N_14991,N_6074,N_9230);
nor U14992 (N_14992,N_9385,N_8681);
or U14993 (N_14993,N_7255,N_9595);
nor U14994 (N_14994,N_5027,N_5310);
and U14995 (N_14995,N_6333,N_9649);
nor U14996 (N_14996,N_5786,N_7969);
nand U14997 (N_14997,N_9987,N_7492);
nor U14998 (N_14998,N_8762,N_8676);
nor U14999 (N_14999,N_7316,N_7695);
xnor U15000 (N_15000,N_13510,N_14855);
nor U15001 (N_15001,N_10635,N_13951);
nand U15002 (N_15002,N_14947,N_10501);
and U15003 (N_15003,N_11862,N_13345);
nand U15004 (N_15004,N_10560,N_10283);
nand U15005 (N_15005,N_10348,N_10448);
and U15006 (N_15006,N_14473,N_12503);
xor U15007 (N_15007,N_14000,N_12092);
nand U15008 (N_15008,N_10985,N_14668);
nor U15009 (N_15009,N_14512,N_10157);
nor U15010 (N_15010,N_14130,N_13112);
nand U15011 (N_15011,N_12280,N_12000);
nand U15012 (N_15012,N_11603,N_10138);
xnor U15013 (N_15013,N_13597,N_12712);
and U15014 (N_15014,N_14238,N_11759);
nand U15015 (N_15015,N_10023,N_14915);
nand U15016 (N_15016,N_11812,N_14450);
or U15017 (N_15017,N_10551,N_11465);
nand U15018 (N_15018,N_13950,N_10204);
and U15019 (N_15019,N_11439,N_10994);
and U15020 (N_15020,N_13586,N_10774);
nand U15021 (N_15021,N_10946,N_14418);
nor U15022 (N_15022,N_12592,N_13116);
and U15023 (N_15023,N_14296,N_13973);
nor U15024 (N_15024,N_12424,N_12049);
nor U15025 (N_15025,N_11770,N_12153);
nor U15026 (N_15026,N_12593,N_14825);
or U15027 (N_15027,N_11123,N_10103);
nand U15028 (N_15028,N_10073,N_14592);
nor U15029 (N_15029,N_10993,N_14550);
nand U15030 (N_15030,N_12668,N_10207);
and U15031 (N_15031,N_13857,N_12998);
or U15032 (N_15032,N_10285,N_13039);
or U15033 (N_15033,N_10528,N_12744);
nand U15034 (N_15034,N_11941,N_14613);
nand U15035 (N_15035,N_14342,N_10469);
xnor U15036 (N_15036,N_12850,N_14294);
nor U15037 (N_15037,N_10851,N_14015);
nor U15038 (N_15038,N_12577,N_10415);
nand U15039 (N_15039,N_14928,N_10789);
nand U15040 (N_15040,N_10158,N_14498);
nand U15041 (N_15041,N_14924,N_12058);
or U15042 (N_15042,N_12071,N_11779);
nor U15043 (N_15043,N_11607,N_12772);
nor U15044 (N_15044,N_14288,N_11416);
and U15045 (N_15045,N_14791,N_10180);
nor U15046 (N_15046,N_13372,N_12108);
and U15047 (N_15047,N_10060,N_13732);
xnor U15048 (N_15048,N_12711,N_10386);
nand U15049 (N_15049,N_14610,N_10772);
nor U15050 (N_15050,N_10403,N_14862);
xor U15051 (N_15051,N_11578,N_10570);
nor U15052 (N_15052,N_13226,N_11846);
or U15053 (N_15053,N_10788,N_14898);
nand U15054 (N_15054,N_10588,N_13984);
nor U15055 (N_15055,N_14198,N_13686);
and U15056 (N_15056,N_14303,N_12670);
nand U15057 (N_15057,N_11494,N_14360);
or U15058 (N_15058,N_12272,N_13759);
nand U15059 (N_15059,N_14606,N_11271);
xnor U15060 (N_15060,N_13336,N_13204);
and U15061 (N_15061,N_11196,N_13040);
xor U15062 (N_15062,N_13472,N_10547);
nor U15063 (N_15063,N_14931,N_11815);
nor U15064 (N_15064,N_10798,N_13632);
and U15065 (N_15065,N_10384,N_10540);
and U15066 (N_15066,N_10886,N_12131);
nor U15067 (N_15067,N_10456,N_11042);
xnor U15068 (N_15068,N_10730,N_12716);
xnor U15069 (N_15069,N_11476,N_12404);
and U15070 (N_15070,N_11143,N_10077);
or U15071 (N_15071,N_12410,N_14093);
nor U15072 (N_15072,N_14828,N_12030);
or U15073 (N_15073,N_10858,N_12776);
xor U15074 (N_15074,N_11313,N_13488);
nor U15075 (N_15075,N_14467,N_14654);
nor U15076 (N_15076,N_13971,N_11972);
nand U15077 (N_15077,N_13952,N_14322);
or U15078 (N_15078,N_11139,N_10380);
nor U15079 (N_15079,N_14234,N_13918);
and U15080 (N_15080,N_12556,N_13388);
and U15081 (N_15081,N_12804,N_12706);
nor U15082 (N_15082,N_14203,N_10099);
xor U15083 (N_15083,N_12758,N_13694);
or U15084 (N_15084,N_10184,N_13313);
and U15085 (N_15085,N_14797,N_13095);
nand U15086 (N_15086,N_12888,N_12165);
and U15087 (N_15087,N_14332,N_11024);
and U15088 (N_15088,N_12393,N_11626);
xnor U15089 (N_15089,N_14653,N_10010);
nor U15090 (N_15090,N_14736,N_14359);
nand U15091 (N_15091,N_12650,N_14035);
nand U15092 (N_15092,N_13363,N_12797);
or U15093 (N_15093,N_12036,N_10022);
nand U15094 (N_15094,N_14516,N_13707);
and U15095 (N_15095,N_11899,N_12295);
nor U15096 (N_15096,N_11702,N_13786);
and U15097 (N_15097,N_10559,N_11664);
and U15098 (N_15098,N_13411,N_14306);
nor U15099 (N_15099,N_10988,N_14064);
nor U15100 (N_15100,N_13937,N_12193);
nand U15101 (N_15101,N_10997,N_12047);
or U15102 (N_15102,N_10032,N_14741);
and U15103 (N_15103,N_13470,N_11793);
nor U15104 (N_15104,N_12315,N_12430);
xor U15105 (N_15105,N_14701,N_11566);
nor U15106 (N_15106,N_11946,N_14054);
or U15107 (N_15107,N_12061,N_11673);
nor U15108 (N_15108,N_14546,N_10967);
and U15109 (N_15109,N_14826,N_10233);
or U15110 (N_15110,N_10741,N_12113);
nor U15111 (N_15111,N_10136,N_11776);
xor U15112 (N_15112,N_12226,N_14199);
xnor U15113 (N_15113,N_11025,N_11484);
and U15114 (N_15114,N_14852,N_14709);
nand U15115 (N_15115,N_13281,N_14095);
nand U15116 (N_15116,N_13268,N_10038);
and U15117 (N_15117,N_14352,N_10148);
or U15118 (N_15118,N_10008,N_11799);
nand U15119 (N_15119,N_11341,N_10497);
and U15120 (N_15120,N_10612,N_12903);
and U15121 (N_15121,N_10290,N_13946);
nand U15122 (N_15122,N_12261,N_14247);
or U15123 (N_15123,N_13282,N_12245);
xnor U15124 (N_15124,N_10553,N_10471);
or U15125 (N_15125,N_11914,N_10583);
or U15126 (N_15126,N_13060,N_10930);
nand U15127 (N_15127,N_12137,N_11022);
or U15128 (N_15128,N_14495,N_13800);
nor U15129 (N_15129,N_12001,N_14047);
and U15130 (N_15130,N_13691,N_10841);
nor U15131 (N_15131,N_10240,N_13748);
nand U15132 (N_15132,N_10241,N_12987);
and U15133 (N_15133,N_11384,N_12639);
nor U15134 (N_15134,N_14887,N_13839);
or U15135 (N_15135,N_10777,N_13464);
and U15136 (N_15136,N_11178,N_14993);
nor U15137 (N_15137,N_13297,N_13585);
nand U15138 (N_15138,N_11882,N_13794);
or U15139 (N_15139,N_10410,N_10688);
nor U15140 (N_15140,N_12100,N_13762);
nand U15141 (N_15141,N_13427,N_10899);
nor U15142 (N_15142,N_11761,N_13574);
nor U15143 (N_15143,N_10272,N_11102);
nor U15144 (N_15144,N_12331,N_11058);
nor U15145 (N_15145,N_10607,N_11550);
or U15146 (N_15146,N_10030,N_14411);
xnor U15147 (N_15147,N_11757,N_14477);
and U15148 (N_15148,N_14397,N_13624);
or U15149 (N_15149,N_10866,N_14201);
nor U15150 (N_15150,N_11834,N_10373);
nor U15151 (N_15151,N_10832,N_14770);
and U15152 (N_15152,N_11093,N_11694);
and U15153 (N_15153,N_12627,N_12297);
nand U15154 (N_15154,N_10467,N_12451);
and U15155 (N_15155,N_13016,N_10938);
or U15156 (N_15156,N_14765,N_10826);
nor U15157 (N_15157,N_12629,N_14548);
and U15158 (N_15158,N_12926,N_10773);
and U15159 (N_15159,N_13399,N_10428);
and U15160 (N_15160,N_11720,N_14399);
and U15161 (N_15161,N_11273,N_12363);
nor U15162 (N_15162,N_14591,N_10481);
nor U15163 (N_15163,N_10557,N_10696);
nand U15164 (N_15164,N_14390,N_14036);
or U15165 (N_15165,N_14070,N_14402);
nor U15166 (N_15166,N_10161,N_11016);
xnor U15167 (N_15167,N_11451,N_12805);
nand U15168 (N_15168,N_11149,N_11639);
and U15169 (N_15169,N_10532,N_10383);
nor U15170 (N_15170,N_14599,N_12962);
or U15171 (N_15171,N_13768,N_11721);
nand U15172 (N_15172,N_10813,N_11863);
nand U15173 (N_15173,N_11806,N_11382);
xnor U15174 (N_15174,N_11684,N_12228);
and U15175 (N_15175,N_12879,N_13658);
nor U15176 (N_15176,N_12464,N_13305);
or U15177 (N_15177,N_10854,N_13481);
nand U15178 (N_15178,N_13214,N_12275);
xnor U15179 (N_15179,N_10662,N_12220);
xnor U15180 (N_15180,N_10418,N_12999);
nor U15181 (N_15181,N_14496,N_11150);
xnor U15182 (N_15182,N_12109,N_11224);
and U15183 (N_15183,N_13067,N_14929);
and U15184 (N_15184,N_13101,N_10794);
xor U15185 (N_15185,N_13247,N_12892);
xnor U15186 (N_15186,N_13178,N_12687);
and U15187 (N_15187,N_11839,N_13660);
and U15188 (N_15188,N_11453,N_10550);
or U15189 (N_15189,N_13432,N_11415);
or U15190 (N_15190,N_10968,N_13107);
nand U15191 (N_15191,N_13493,N_10232);
and U15192 (N_15192,N_11873,N_14018);
or U15193 (N_15193,N_14807,N_10527);
nor U15194 (N_15194,N_14998,N_14953);
or U15195 (N_15195,N_14588,N_14499);
and U15196 (N_15196,N_12619,N_11199);
nand U15197 (N_15197,N_13706,N_12886);
and U15198 (N_15198,N_11127,N_14661);
and U15199 (N_15199,N_10438,N_10529);
nand U15200 (N_15200,N_10931,N_14253);
and U15201 (N_15201,N_10745,N_11810);
nor U15202 (N_15202,N_11750,N_12831);
or U15203 (N_15203,N_12548,N_13054);
or U15204 (N_15204,N_14539,N_11924);
or U15205 (N_15205,N_14721,N_14270);
xor U15206 (N_15206,N_14514,N_13299);
xnor U15207 (N_15207,N_11174,N_12320);
nor U15208 (N_15208,N_12009,N_13514);
or U15209 (N_15209,N_13128,N_11852);
nand U15210 (N_15210,N_14367,N_13277);
nand U15211 (N_15211,N_11619,N_14124);
or U15212 (N_15212,N_13939,N_10883);
nor U15213 (N_15213,N_13303,N_12027);
and U15214 (N_15214,N_11867,N_13661);
nor U15215 (N_15215,N_13530,N_10932);
nand U15216 (N_15216,N_11755,N_12209);
or U15217 (N_15217,N_11786,N_10133);
xor U15218 (N_15218,N_10606,N_13004);
and U15219 (N_15219,N_10024,N_14478);
xnor U15220 (N_15220,N_14281,N_14380);
and U15221 (N_15221,N_10127,N_12042);
and U15222 (N_15222,N_11589,N_11039);
or U15223 (N_15223,N_10096,N_14401);
and U15224 (N_15224,N_12172,N_11577);
and U15225 (N_15225,N_11335,N_14747);
and U15226 (N_15226,N_12858,N_14959);
nor U15227 (N_15227,N_14967,N_11175);
nor U15228 (N_15228,N_11712,N_12943);
or U15229 (N_15229,N_14774,N_14318);
xnor U15230 (N_15230,N_10189,N_12395);
or U15231 (N_15231,N_14347,N_14176);
xor U15232 (N_15232,N_11671,N_12074);
and U15233 (N_15233,N_13958,N_13217);
or U15234 (N_15234,N_11256,N_12221);
nand U15235 (N_15235,N_13743,N_12972);
or U15236 (N_15236,N_13075,N_12814);
and U15237 (N_15237,N_11238,N_13292);
nor U15238 (N_15238,N_11134,N_13288);
or U15239 (N_15239,N_12572,N_13199);
and U15240 (N_15240,N_11710,N_11269);
and U15241 (N_15241,N_14594,N_14614);
or U15242 (N_15242,N_12002,N_11165);
nor U15243 (N_15243,N_13249,N_10039);
and U15244 (N_15244,N_10785,N_10359);
nor U15245 (N_15245,N_12928,N_12021);
nor U15246 (N_15246,N_11825,N_10581);
nor U15247 (N_15247,N_11816,N_11686);
and U15248 (N_15248,N_13190,N_12095);
xnor U15249 (N_15249,N_12422,N_12440);
and U15250 (N_15250,N_10442,N_12233);
xor U15251 (N_15251,N_10677,N_14188);
nand U15252 (N_15252,N_12124,N_10421);
xnor U15253 (N_15253,N_13989,N_14366);
or U15254 (N_15254,N_13494,N_14143);
nor U15255 (N_15255,N_13244,N_12833);
nand U15256 (N_15256,N_10712,N_12082);
or U15257 (N_15257,N_12159,N_10939);
nor U15258 (N_15258,N_14532,N_10728);
or U15259 (N_15259,N_12466,N_12586);
nor U15260 (N_15260,N_12685,N_14687);
nor U15261 (N_15261,N_11172,N_13877);
and U15262 (N_15262,N_10050,N_13122);
nand U15263 (N_15263,N_11186,N_10424);
or U15264 (N_15264,N_12116,N_10273);
nor U15265 (N_15265,N_11192,N_13780);
or U15266 (N_15266,N_10895,N_13499);
or U15267 (N_15267,N_13591,N_10731);
nor U15268 (N_15268,N_13572,N_10166);
or U15269 (N_15269,N_13925,N_13182);
and U15270 (N_15270,N_14519,N_14547);
or U15271 (N_15271,N_14507,N_13327);
nand U15272 (N_15272,N_12876,N_11448);
nand U15273 (N_15273,N_12816,N_11412);
nand U15274 (N_15274,N_12256,N_14046);
nand U15275 (N_15275,N_13923,N_12319);
or U15276 (N_15276,N_12278,N_14739);
nand U15277 (N_15277,N_10372,N_10294);
nor U15278 (N_15278,N_13695,N_11975);
nor U15279 (N_15279,N_13964,N_11742);
and U15280 (N_15280,N_13955,N_11983);
xnor U15281 (N_15281,N_12849,N_10909);
nand U15282 (N_15282,N_10561,N_14415);
and U15283 (N_15283,N_13023,N_10164);
or U15284 (N_15284,N_13310,N_10811);
nand U15285 (N_15285,N_10873,N_11754);
nor U15286 (N_15286,N_13053,N_12733);
and U15287 (N_15287,N_14982,N_13015);
nand U15288 (N_15288,N_14878,N_13522);
or U15289 (N_15289,N_13814,N_13259);
nand U15290 (N_15290,N_12514,N_14564);
or U15291 (N_15291,N_12832,N_13169);
or U15292 (N_15292,N_11969,N_13334);
and U15293 (N_15293,N_11414,N_10847);
nor U15294 (N_15294,N_13570,N_10107);
or U15295 (N_15295,N_10258,N_14902);
or U15296 (N_15296,N_14986,N_11140);
and U15297 (N_15297,N_14321,N_12625);
nand U15298 (N_15298,N_13717,N_12622);
nor U15299 (N_15299,N_10036,N_12559);
xor U15300 (N_15300,N_11278,N_12371);
and U15301 (N_15301,N_13698,N_13202);
or U15302 (N_15302,N_12800,N_14008);
nor U15303 (N_15303,N_12249,N_14920);
and U15304 (N_15304,N_12346,N_14034);
nand U15305 (N_15305,N_11680,N_13999);
or U15306 (N_15306,N_13631,N_11602);
xor U15307 (N_15307,N_14671,N_14102);
or U15308 (N_15308,N_12325,N_10709);
nand U15309 (N_15309,N_13225,N_12142);
or U15310 (N_15310,N_13507,N_12755);
xnor U15311 (N_15311,N_14596,N_10262);
nor U15312 (N_15312,N_14842,N_10964);
xor U15313 (N_15313,N_10948,N_11843);
nor U15314 (N_15314,N_10076,N_13393);
nand U15315 (N_15315,N_12232,N_11803);
and U15316 (N_15316,N_12538,N_13492);
nand U15317 (N_15317,N_12475,N_12223);
xnor U15318 (N_15318,N_13189,N_13068);
nand U15319 (N_15319,N_11253,N_14424);
and U15320 (N_15320,N_11753,N_12033);
nand U15321 (N_15321,N_10009,N_12667);
nor U15322 (N_15322,N_13934,N_10223);
or U15323 (N_15323,N_12553,N_12683);
nor U15324 (N_15324,N_11660,N_14118);
nand U15325 (N_15325,N_12219,N_12678);
nor U15326 (N_15326,N_14704,N_13765);
or U15327 (N_15327,N_10393,N_10183);
nor U15328 (N_15328,N_12923,N_10308);
nand U15329 (N_15329,N_12413,N_14573);
nor U15330 (N_15330,N_13823,N_12182);
or U15331 (N_15331,N_14077,N_11728);
and U15332 (N_15332,N_11512,N_13688);
nor U15333 (N_15333,N_12300,N_12782);
nor U15334 (N_15334,N_14438,N_14699);
and U15335 (N_15335,N_11670,N_13761);
and U15336 (N_15336,N_10427,N_10436);
nand U15337 (N_15337,N_14137,N_12840);
or U15338 (N_15338,N_14927,N_11001);
or U15339 (N_15339,N_11301,N_10515);
xor U15340 (N_15340,N_11109,N_13298);
and U15341 (N_15341,N_10548,N_10005);
nor U15342 (N_15342,N_11356,N_11966);
xnor U15343 (N_15343,N_12296,N_14702);
xor U15344 (N_15344,N_12358,N_12313);
and U15345 (N_15345,N_11961,N_10818);
and U15346 (N_15346,N_13617,N_11203);
or U15347 (N_15347,N_13087,N_10454);
and U15348 (N_15348,N_13469,N_10605);
and U15349 (N_15349,N_13014,N_12271);
and U15350 (N_15350,N_13519,N_11044);
nor U15351 (N_15351,N_12705,N_11145);
and U15352 (N_15352,N_13001,N_13733);
nor U15353 (N_15353,N_12872,N_11866);
and U15354 (N_15354,N_12736,N_13098);
nand U15355 (N_15355,N_11040,N_14462);
nand U15356 (N_15356,N_10848,N_11171);
nor U15357 (N_15357,N_11677,N_10235);
nand U15358 (N_15358,N_10889,N_11299);
nand U15359 (N_15359,N_10770,N_11324);
or U15360 (N_15360,N_13207,N_13440);
nor U15361 (N_15361,N_10500,N_11691);
nor U15362 (N_15362,N_11420,N_10679);
nand U15363 (N_15363,N_12243,N_10823);
nor U15364 (N_15364,N_12050,N_12195);
xnor U15365 (N_15365,N_12427,N_10014);
and U15366 (N_15366,N_11887,N_10535);
or U15367 (N_15367,N_12255,N_10920);
and U15368 (N_15368,N_11855,N_10095);
and U15369 (N_15369,N_10460,N_11170);
and U15370 (N_15370,N_11387,N_14955);
or U15371 (N_15371,N_12248,N_11344);
nor U15372 (N_15372,N_14187,N_13394);
nand U15373 (N_15373,N_14793,N_10914);
or U15374 (N_15374,N_11153,N_10863);
xor U15375 (N_15375,N_13455,N_11478);
xnor U15376 (N_15376,N_10695,N_14043);
or U15377 (N_15377,N_11413,N_13398);
nand U15378 (N_15378,N_13516,N_12884);
or U15379 (N_15379,N_10324,N_14572);
and U15380 (N_15380,N_10354,N_13943);
and U15381 (N_15381,N_10657,N_11369);
and U15382 (N_15382,N_12873,N_11185);
nand U15383 (N_15383,N_11830,N_11556);
xnor U15384 (N_15384,N_14363,N_14628);
xor U15385 (N_15385,N_10724,N_12495);
xnor U15386 (N_15386,N_12561,N_12380);
nor U15387 (N_15387,N_11459,N_10057);
nand U15388 (N_15388,N_11479,N_13708);
or U15389 (N_15389,N_14503,N_11361);
and U15390 (N_15390,N_14700,N_12337);
nand U15391 (N_15391,N_13020,N_11560);
and U15392 (N_15392,N_12088,N_14232);
nand U15393 (N_15393,N_14189,N_12516);
or U15394 (N_15394,N_10664,N_11108);
nor U15395 (N_15395,N_11938,N_12183);
xnor U15396 (N_15396,N_11426,N_10865);
and U15397 (N_15397,N_14108,N_10905);
and U15398 (N_15398,N_13049,N_11934);
nand U15399 (N_15399,N_10182,N_11661);
and U15400 (N_15400,N_10408,N_14427);
nor U15401 (N_15401,N_11083,N_13667);
nor U15402 (N_15402,N_10170,N_11408);
nand U15403 (N_15403,N_10167,N_11101);
nand U15404 (N_15404,N_12607,N_14895);
or U15405 (N_15405,N_12575,N_11762);
or U15406 (N_15406,N_14973,N_12590);
and U15407 (N_15407,N_10042,N_13656);
nand U15408 (N_15408,N_13302,N_11687);
and U15409 (N_15409,N_13562,N_12633);
nor U15410 (N_15410,N_14492,N_12551);
or U15411 (N_15411,N_13414,N_10970);
and U15412 (N_15412,N_10213,N_10470);
nand U15413 (N_15413,N_12789,N_13361);
nor U15414 (N_15414,N_13969,N_10817);
nand U15415 (N_15415,N_12354,N_14975);
and U15416 (N_15416,N_12127,N_13273);
and U15417 (N_15417,N_14755,N_11999);
nand U15418 (N_15418,N_12930,N_14286);
nand U15419 (N_15419,N_14313,N_10526);
or U15420 (N_15420,N_11137,N_14241);
and U15421 (N_15421,N_11425,N_13272);
nor U15422 (N_15422,N_14864,N_13752);
nand U15423 (N_15423,N_10649,N_11122);
and U15424 (N_15424,N_13265,N_14529);
and U15425 (N_15425,N_12834,N_14814);
nand U15426 (N_15426,N_14589,N_11620);
or U15427 (N_15427,N_13364,N_12947);
nand U15428 (N_15428,N_11698,N_14375);
and U15429 (N_15429,N_13161,N_11539);
nand U15430 (N_15430,N_14555,N_10545);
and U15431 (N_15431,N_12084,N_11031);
nand U15432 (N_15432,N_12155,N_12026);
or U15433 (N_15433,N_13828,N_11049);
nand U15434 (N_15434,N_11537,N_12734);
nor U15435 (N_15435,N_14212,N_14940);
and U15436 (N_15436,N_14263,N_12569);
and U15437 (N_15437,N_11628,N_14307);
and U15438 (N_15438,N_10986,N_10725);
or U15439 (N_15439,N_10726,N_12138);
or U15440 (N_15440,N_14673,N_13865);
or U15441 (N_15441,N_12680,N_11454);
nand U15442 (N_15442,N_10414,N_12645);
or U15443 (N_15443,N_11404,N_13536);
or U15444 (N_15444,N_10463,N_12485);
nand U15445 (N_15445,N_10435,N_12502);
and U15446 (N_15446,N_14480,N_11717);
or U15447 (N_15447,N_12383,N_10027);
xnor U15448 (N_15448,N_13612,N_13228);
nor U15449 (N_15449,N_11505,N_10844);
nand U15450 (N_15450,N_13367,N_14521);
nor U15451 (N_15451,N_13319,N_11474);
nor U15452 (N_15452,N_13389,N_10703);
and U15453 (N_15453,N_13383,N_13858);
nand U15454 (N_15454,N_13847,N_11032);
and U15455 (N_15455,N_10302,N_11239);
nand U15456 (N_15456,N_11504,N_11875);
or U15457 (N_15457,N_11591,N_13235);
xnor U15458 (N_15458,N_10434,N_13033);
or U15459 (N_15459,N_11115,N_14984);
xnor U15460 (N_15460,N_12925,N_11460);
or U15461 (N_15461,N_13252,N_14436);
xnor U15462 (N_15462,N_11284,N_14131);
xor U15463 (N_15463,N_10655,N_10714);
or U15464 (N_15464,N_10202,N_14487);
and U15465 (N_15465,N_11160,N_10768);
and U15466 (N_15466,N_11015,N_13370);
and U15467 (N_15467,N_14966,N_10831);
nor U15468 (N_15468,N_13255,N_13554);
and U15469 (N_15469,N_11877,N_10861);
nor U15470 (N_15470,N_10510,N_14013);
nor U15471 (N_15471,N_12937,N_11265);
nor U15472 (N_15472,N_10626,N_12902);
or U15473 (N_15473,N_13135,N_14756);
nand U15474 (N_15474,N_14361,N_12311);
xor U15475 (N_15475,N_11385,N_13106);
nand U15476 (N_15476,N_10162,N_13931);
and U15477 (N_15477,N_12406,N_12274);
xor U15478 (N_15478,N_11007,N_11871);
or U15479 (N_15479,N_12669,N_10398);
nand U15480 (N_15480,N_13719,N_10052);
nor U15481 (N_15481,N_12157,N_10867);
or U15482 (N_15482,N_13730,N_10694);
xor U15483 (N_15483,N_14935,N_14060);
nor U15484 (N_15484,N_14751,N_14264);
and U15485 (N_15485,N_12339,N_10020);
nor U15486 (N_15486,N_10622,N_11989);
nor U15487 (N_15487,N_13876,N_11821);
or U15488 (N_15488,N_11864,N_11388);
xor U15489 (N_15489,N_10576,N_12149);
and U15490 (N_15490,N_14847,N_10297);
and U15491 (N_15491,N_13967,N_14441);
or U15492 (N_15492,N_10852,N_14162);
nor U15493 (N_15493,N_13788,N_14491);
or U15494 (N_15494,N_12842,N_12614);
nand U15495 (N_15495,N_14630,N_12072);
nand U15496 (N_15496,N_13861,N_13728);
and U15497 (N_15497,N_14713,N_13099);
or U15498 (N_15498,N_14204,N_12162);
and U15499 (N_15499,N_12709,N_14048);
xor U15500 (N_15500,N_12321,N_14871);
and U15501 (N_15501,N_14430,N_10402);
or U15502 (N_15502,N_10019,N_12521);
nor U15503 (N_15503,N_14084,N_13309);
nand U15504 (N_15504,N_10585,N_12231);
xnor U15505 (N_15505,N_10321,N_12034);
nor U15506 (N_15506,N_10305,N_10109);
nand U15507 (N_15507,N_12342,N_10681);
nand U15508 (N_15508,N_10417,N_14537);
nand U15509 (N_15509,N_14784,N_13197);
and U15510 (N_15510,N_11587,N_12103);
or U15511 (N_15511,N_11200,N_12490);
nor U15512 (N_15512,N_12520,N_12343);
and U15513 (N_15513,N_13474,N_14886);
or U15514 (N_15514,N_13286,N_14261);
nand U15515 (N_15515,N_11189,N_12438);
or U15516 (N_15516,N_10544,N_10225);
nor U15517 (N_15517,N_12006,N_11772);
nand U15518 (N_15518,N_11407,N_12971);
nand U15519 (N_15519,N_10563,N_12004);
nor U15520 (N_15520,N_11151,N_10053);
or U15521 (N_15521,N_10644,N_12580);
nand U15522 (N_15522,N_11167,N_13995);
nand U15523 (N_15523,N_11051,N_12803);
nand U15524 (N_15524,N_13219,N_10836);
or U15525 (N_15525,N_12398,N_11142);
nor U15526 (N_15526,N_10758,N_12106);
and U15527 (N_15527,N_13483,N_12436);
xnor U15528 (N_15528,N_11209,N_14652);
nor U15529 (N_15529,N_12511,N_13052);
or U15530 (N_15530,N_10450,N_14896);
nand U15531 (N_15531,N_11461,N_10680);
nand U15532 (N_15532,N_12156,N_12953);
and U15533 (N_15533,N_13433,N_11738);
or U15534 (N_15534,N_13571,N_10879);
or U15535 (N_15535,N_11807,N_13172);
nand U15536 (N_15536,N_14180,N_11883);
nor U15537 (N_15537,N_13579,N_11976);
xnor U15538 (N_15538,N_10723,N_14722);
or U15539 (N_15539,N_11586,N_13760);
nand U15540 (N_15540,N_12180,N_11748);
nor U15541 (N_15541,N_10891,N_14945);
nand U15542 (N_15542,N_10830,N_10565);
or U15543 (N_15543,N_11154,N_13245);
or U15544 (N_15544,N_14951,N_11350);
nor U15545 (N_15545,N_12423,N_14149);
nor U15546 (N_15546,N_12381,N_11767);
nand U15547 (N_15547,N_13956,N_12396);
and U15548 (N_15548,N_11509,N_14609);
or U15549 (N_15549,N_13168,N_11813);
xor U15550 (N_15550,N_13030,N_12277);
or U15551 (N_15551,N_11105,N_11943);
xor U15552 (N_15552,N_10792,N_14466);
and U15553 (N_15553,N_10819,N_12164);
and U15554 (N_15554,N_13232,N_10295);
or U15555 (N_15555,N_13086,N_13236);
xnor U15556 (N_15556,N_13230,N_12871);
nor U15557 (N_15557,N_13439,N_11645);
or U15558 (N_15558,N_11900,N_14746);
and U15559 (N_15559,N_12416,N_11700);
or U15560 (N_15560,N_14685,N_14773);
or U15561 (N_15561,N_13606,N_10115);
or U15562 (N_15562,N_11784,N_11874);
and U15563 (N_15563,N_12461,N_12038);
nor U15564 (N_15564,N_14033,N_10686);
nand U15565 (N_15565,N_12839,N_14683);
or U15566 (N_15566,N_11611,N_10683);
or U15567 (N_15567,N_13495,N_13634);
nor U15568 (N_15568,N_11314,N_11320);
nand U15569 (N_15569,N_12299,N_12679);
nor U15570 (N_15570,N_10803,N_11094);
xnor U15571 (N_15571,N_11971,N_12390);
nand U15572 (N_15572,N_13789,N_11630);
and U15573 (N_15573,N_13349,N_11547);
and U15574 (N_15574,N_12129,N_12005);
nand U15575 (N_15575,N_12236,N_14963);
nand U15576 (N_15576,N_13032,N_12985);
or U15577 (N_15577,N_11464,N_14349);
or U15578 (N_15578,N_11087,N_11879);
nand U15579 (N_15579,N_14827,N_12012);
nand U15580 (N_15580,N_11397,N_11402);
and U15581 (N_15581,N_10685,N_11741);
nor U15582 (N_15582,N_13945,N_11681);
nand U15583 (N_15583,N_14718,N_13758);
xor U15584 (N_15584,N_12967,N_11099);
and U15585 (N_15585,N_14273,N_13954);
or U15586 (N_15586,N_13712,N_14090);
and U15587 (N_15587,N_14501,N_11695);
or U15588 (N_15588,N_13156,N_10592);
xnor U15589 (N_15589,N_12146,N_10996);
or U15590 (N_15590,N_13021,N_13976);
or U15591 (N_15591,N_11184,N_12563);
xor U15592 (N_15592,N_11013,N_14804);
nand U15593 (N_15593,N_11522,N_11510);
or U15594 (N_15594,N_12719,N_10080);
or U15595 (N_15595,N_12112,N_12114);
nor U15596 (N_15596,N_12023,N_14298);
nor U15597 (N_15597,N_10894,N_13287);
nor U15598 (N_15598,N_14910,N_10656);
or U15599 (N_15599,N_13435,N_14992);
nand U15600 (N_15600,N_11181,N_13250);
nor U15601 (N_15601,N_13801,N_10089);
and U15602 (N_15602,N_14062,N_13485);
or U15603 (N_15603,N_10678,N_14447);
and U15604 (N_15604,N_11456,N_13140);
nand U15605 (N_15605,N_14937,N_13831);
nor U15606 (N_15606,N_13234,N_14824);
and U15607 (N_15607,N_11090,N_10211);
and U15608 (N_15608,N_12718,N_11230);
or U15609 (N_15609,N_11658,N_13625);
and U15610 (N_15610,N_10468,N_12096);
or U15611 (N_15611,N_10074,N_13314);
or U15612 (N_15612,N_14806,N_14482);
or U15613 (N_15613,N_13509,N_12039);
xor U15614 (N_15614,N_11618,N_14971);
nand U15615 (N_15615,N_10834,N_14374);
and U15616 (N_15616,N_12702,N_13248);
or U15617 (N_15617,N_10864,N_14003);
nand U15618 (N_15618,N_11377,N_12062);
xor U15619 (N_15619,N_10494,N_14063);
and U15620 (N_15620,N_13317,N_12980);
and U15621 (N_15621,N_10495,N_11318);
nor U15622 (N_15622,N_10266,N_10575);
xnor U15623 (N_15623,N_10318,N_14239);
and U15624 (N_15624,N_14250,N_10114);
nand U15625 (N_15625,N_10749,N_12811);
and U15626 (N_15626,N_11796,N_13137);
nor U15627 (N_15627,N_10111,N_13409);
and U15628 (N_15628,N_10849,N_13491);
xor U15629 (N_15629,N_11466,N_13038);
nor U15630 (N_15630,N_12582,N_12990);
and U15631 (N_15631,N_14873,N_11084);
nand U15632 (N_15632,N_14672,N_12933);
xnor U15633 (N_15633,N_11555,N_12699);
or U15634 (N_15634,N_13919,N_10522);
nor U15635 (N_15635,N_13149,N_10667);
nand U15636 (N_15636,N_14860,N_12509);
nor U15637 (N_15637,N_11517,N_12905);
nand U15638 (N_15638,N_12877,N_10693);
xnor U15639 (N_15639,N_12426,N_14811);
or U15640 (N_15640,N_14259,N_14178);
and U15641 (N_15641,N_13147,N_14730);
or U15642 (N_15642,N_11627,N_13838);
nand U15643 (N_15643,N_12978,N_14074);
nor U15644 (N_15644,N_10268,N_13410);
or U15645 (N_15645,N_13549,N_10573);
nor U15646 (N_15646,N_12628,N_10382);
and U15647 (N_15647,N_14423,N_13556);
and U15648 (N_15648,N_14370,N_13256);
nand U15649 (N_15649,N_10094,N_12316);
and U15650 (N_15650,N_12135,N_14777);
and U15651 (N_15651,N_10331,N_12016);
or U15652 (N_15652,N_14780,N_13845);
or U15653 (N_15653,N_13103,N_13048);
or U15654 (N_15654,N_12965,N_11352);
or U15655 (N_15655,N_14843,N_10490);
or U15656 (N_15656,N_13643,N_14612);
or U15657 (N_15657,N_10775,N_12573);
nand U15658 (N_15658,N_10542,N_13329);
or U15659 (N_15659,N_13921,N_13051);
or U15660 (N_15660,N_14340,N_13035);
or U15661 (N_15661,N_12500,N_10280);
or U15662 (N_15662,N_11251,N_12666);
nor U15663 (N_15663,N_12636,N_11292);
or U15664 (N_15664,N_10720,N_14205);
nor U15665 (N_15665,N_14566,N_12769);
nor U15666 (N_15666,N_14011,N_13907);
nand U15667 (N_15667,N_10228,N_13194);
nand U15668 (N_15668,N_10992,N_13927);
nand U15669 (N_15669,N_10193,N_13423);
xnor U15670 (N_15670,N_10732,N_11405);
nand U15671 (N_15671,N_10533,N_11706);
nor U15672 (N_15672,N_12507,N_13825);
or U15673 (N_15673,N_10098,N_10660);
nor U15674 (N_15674,N_14752,N_11854);
nand U15675 (N_15675,N_14989,N_14136);
nand U15676 (N_15676,N_10156,N_10461);
and U15677 (N_15677,N_14454,N_13963);
or U15678 (N_15678,N_13443,N_12979);
or U15679 (N_15679,N_12856,N_14448);
or U15680 (N_15680,N_13872,N_12085);
and U15681 (N_15681,N_11100,N_11657);
nor U15682 (N_15682,N_12764,N_10227);
or U15683 (N_15683,N_13767,N_14169);
and U15684 (N_15684,N_11243,N_14511);
and U15685 (N_15685,N_14839,N_10610);
nand U15686 (N_15686,N_12830,N_14735);
nand U15687 (N_15687,N_12497,N_12753);
nand U15688 (N_15688,N_11915,N_12265);
nor U15689 (N_15689,N_11919,N_10721);
or U15690 (N_15690,N_12494,N_12684);
and U15691 (N_15691,N_12428,N_10287);
and U15692 (N_15692,N_14651,N_14578);
xnor U15693 (N_15693,N_10360,N_11814);
xor U15694 (N_15694,N_12080,N_14894);
or U15695 (N_15695,N_14643,N_12653);
xnor U15696 (N_15696,N_10739,N_10025);
and U15697 (N_15697,N_12094,N_14874);
nand U15698 (N_15698,N_14891,N_10595);
or U15699 (N_15699,N_14944,N_14163);
and U15700 (N_15700,N_13774,N_10590);
nor U15701 (N_15701,N_14088,N_10807);
and U15702 (N_15702,N_13843,N_12289);
nor U15703 (N_15703,N_12608,N_11788);
or U15704 (N_15704,N_14236,N_12958);
and U15705 (N_15705,N_13498,N_14880);
and U15706 (N_15706,N_12779,N_11308);
and U15707 (N_15707,N_14087,N_14502);
nor U15708 (N_15708,N_13110,N_13124);
nor U15709 (N_15709,N_11354,N_13867);
nand U15710 (N_15710,N_14517,N_14422);
xor U15711 (N_15711,N_12986,N_14794);
nor U15712 (N_15712,N_13347,N_10346);
or U15713 (N_15713,N_12432,N_10253);
nor U15714 (N_15714,N_10137,N_14508);
xor U15715 (N_15715,N_10625,N_13741);
or U15716 (N_15716,N_12493,N_14939);
xor U15717 (N_15717,N_12823,N_11467);
or U15718 (N_15718,N_14042,N_13775);
nor U15719 (N_15719,N_10314,N_11434);
nor U15720 (N_15720,N_13262,N_11506);
or U15721 (N_15721,N_10796,N_11124);
and U15722 (N_15722,N_13704,N_12492);
or U15723 (N_15723,N_14908,N_12752);
and U15724 (N_15724,N_11390,N_11339);
xor U15725 (N_15725,N_14428,N_12983);
and U15726 (N_15726,N_10972,N_10088);
nand U15727 (N_15727,N_10399,N_13848);
nand U15728 (N_15728,N_10962,N_12796);
or U15729 (N_15729,N_11368,N_14115);
nor U15730 (N_15730,N_14289,N_13630);
nor U15731 (N_15731,N_12724,N_14039);
nor U15732 (N_15732,N_10928,N_14484);
and U15733 (N_15733,N_13258,N_13076);
nand U15734 (N_15734,N_14055,N_12056);
xor U15735 (N_15735,N_12533,N_12565);
nand U15736 (N_15736,N_11218,N_10049);
xor U15737 (N_15737,N_13502,N_11158);
xnor U15738 (N_15738,N_12117,N_13192);
xnor U15739 (N_15739,N_14160,N_12412);
xor U15740 (N_15740,N_12869,N_12324);
and U15741 (N_15741,N_14829,N_11820);
nor U15742 (N_15742,N_10707,N_10484);
or U15743 (N_15743,N_10653,N_13211);
nand U15744 (N_15744,N_14969,N_14867);
nand U15745 (N_15745,N_11632,N_14650);
nor U15746 (N_15746,N_11764,N_10507);
xnor U15747 (N_15747,N_14522,N_11840);
or U15748 (N_15748,N_11861,N_12644);
nand U15749 (N_15749,N_10328,N_10842);
or U15750 (N_15750,N_14579,N_13368);
nor U15751 (N_15751,N_13987,N_13079);
nand U15752 (N_15752,N_14684,N_11483);
and U15753 (N_15753,N_13224,N_13009);
nor U15754 (N_15754,N_13864,N_13824);
and U15755 (N_15755,N_11069,N_10719);
nand U15756 (N_15756,N_12471,N_12051);
or U15757 (N_15757,N_14688,N_11274);
nand U15758 (N_15758,N_12328,N_11849);
nand U15759 (N_15759,N_14304,N_10430);
and U15760 (N_15760,N_13155,N_13560);
nor U15761 (N_15761,N_13567,N_14429);
or U15762 (N_15762,N_11781,N_13866);
nand U15763 (N_15763,N_12686,N_11227);
nand U15764 (N_15764,N_14242,N_11870);
nor U15765 (N_15765,N_10191,N_10840);
nor U15766 (N_15766,N_12244,N_10449);
nor U15767 (N_15767,N_11832,N_10199);
nand U15768 (N_15768,N_11532,N_13895);
nor U15769 (N_15769,N_14526,N_12907);
nor U15770 (N_15770,N_14666,N_10718);
or U15771 (N_15771,N_12123,N_11472);
nand U15772 (N_15772,N_11121,N_12266);
nor U15773 (N_15773,N_11190,N_11008);
nand U15774 (N_15774,N_12602,N_12418);
or U15775 (N_15775,N_13335,N_10284);
and U15776 (N_15776,N_13915,N_14338);
nor U15777 (N_15777,N_11237,N_12472);
nand U15778 (N_15778,N_12140,N_12911);
nand U15779 (N_15779,N_11856,N_10369);
or U15780 (N_15780,N_10300,N_13713);
or U15781 (N_15781,N_14145,N_12927);
nand U15782 (N_15782,N_13716,N_14575);
nand U15783 (N_15783,N_10673,N_13091);
nor U15784 (N_15784,N_14875,N_13384);
nor U15785 (N_15785,N_11876,N_11869);
or U15786 (N_15786,N_10558,N_13682);
and U15787 (N_15787,N_12098,N_12454);
nand U15788 (N_15788,N_11080,N_11316);
nor U15789 (N_15789,N_13690,N_12460);
and U15790 (N_15790,N_11254,N_10058);
or U15791 (N_15791,N_14226,N_10129);
or U15792 (N_15792,N_10927,N_13284);
nand U15793 (N_15793,N_11903,N_13216);
nand U15794 (N_15794,N_10394,N_12453);
and U15795 (N_15795,N_11208,N_14767);
nor U15796 (N_15796,N_12882,N_10850);
or U15797 (N_15797,N_13901,N_11944);
nor U15798 (N_15798,N_12043,N_12480);
or U15799 (N_15799,N_13646,N_11307);
or U15800 (N_15800,N_13077,N_10108);
xor U15801 (N_15801,N_14598,N_10222);
or U15802 (N_15802,N_13993,N_13933);
and U15803 (N_15803,N_14020,N_12641);
nand U15804 (N_15804,N_11642,N_13027);
or U15805 (N_15805,N_12078,N_10648);
nor U15806 (N_15806,N_12385,N_13856);
and U15807 (N_15807,N_12007,N_10234);
nor U15808 (N_15808,N_10855,N_12931);
nor U15809 (N_15809,N_10037,N_12865);
or U15810 (N_15810,N_10665,N_14941);
xnor U15811 (N_15811,N_13701,N_13813);
and U15812 (N_15812,N_13118,N_13365);
or U15813 (N_15813,N_10958,N_11447);
or U15814 (N_15814,N_12483,N_12576);
nand U15815 (N_15815,N_12604,N_11559);
and U15816 (N_15816,N_12809,N_12025);
and U15817 (N_15817,N_11910,N_12040);
xnor U15818 (N_15818,N_11366,N_10641);
and U15819 (N_15819,N_14227,N_13868);
nor U15820 (N_15820,N_10578,N_11046);
xnor U15821 (N_15821,N_12110,N_10041);
or U15822 (N_15822,N_11948,N_12045);
nand U15823 (N_15823,N_13322,N_12929);
nand U15824 (N_15824,N_12708,N_11068);
nor U15825 (N_15825,N_11562,N_10046);
nor U15826 (N_15826,N_10556,N_11678);
and U15827 (N_15827,N_14622,N_13929);
nor U15828 (N_15828,N_11010,N_12400);
nand U15829 (N_15829,N_12194,N_14607);
nor U15830 (N_15830,N_13283,N_13260);
xnor U15831 (N_15831,N_11654,N_13157);
nand U15832 (N_15832,N_11631,N_11475);
or U15833 (N_15833,N_13911,N_12912);
or U15834 (N_15834,N_13576,N_13648);
nor U15835 (N_15835,N_11111,N_10900);
nand U15836 (N_15836,N_13799,N_13807);
nor U15837 (N_15837,N_14823,N_14580);
nand U15838 (N_15838,N_13677,N_13885);
or U15839 (N_15839,N_10846,N_10121);
and U15840 (N_15840,N_12204,N_13390);
nor U15841 (N_15841,N_12024,N_11701);
and U15842 (N_15842,N_12738,N_13424);
xnor U15843 (N_15843,N_14656,N_13962);
nand U15844 (N_15844,N_10684,N_12196);
and U15845 (N_15845,N_12510,N_13090);
nor U15846 (N_15846,N_11629,N_13702);
nor U15847 (N_15847,N_13601,N_14272);
and U15848 (N_15848,N_14369,N_12722);
and U15849 (N_15849,N_13293,N_11898);
and U15850 (N_15850,N_14445,N_14132);
nor U15851 (N_15851,N_10951,N_10120);
or U15852 (N_15852,N_11279,N_13773);
nor U15853 (N_15853,N_12658,N_12474);
nand U15854 (N_15854,N_10257,N_14625);
and U15855 (N_15855,N_14800,N_14412);
and U15856 (N_15856,N_13180,N_12918);
nor U15857 (N_15857,N_11255,N_14834);
nor U15858 (N_15858,N_14626,N_13022);
xnor U15859 (N_15859,N_12771,N_14761);
nor U15860 (N_15860,N_12065,N_12382);
or U15861 (N_15861,N_13994,N_13640);
and U15862 (N_15862,N_13829,N_12044);
nand U15863 (N_15863,N_14392,N_11928);
nand U15864 (N_15864,N_10956,N_12022);
and U15865 (N_15865,N_12306,N_13842);
or U15866 (N_15866,N_14876,N_11163);
nand U15867 (N_15867,N_14435,N_11957);
nand U15868 (N_15868,N_13121,N_12340);
nor U15869 (N_15869,N_14440,N_12963);
nand U15870 (N_15870,N_11266,N_10659);
nand U15871 (N_15871,N_10420,N_12158);
nand U15872 (N_15872,N_10999,N_13869);
nand U15873 (N_15873,N_11519,N_14616);
nand U15874 (N_15874,N_12285,N_11338);
or U15875 (N_15875,N_14717,N_10853);
nor U15876 (N_15876,N_14356,N_12356);
nor U15877 (N_15877,N_11794,N_11666);
nand U15878 (N_15878,N_10619,N_11217);
and U15879 (N_15879,N_13436,N_14726);
nand U15880 (N_15880,N_11703,N_11551);
and U15881 (N_15881,N_10276,N_13878);
nor U15882 (N_15882,N_13378,N_14759);
nand U15883 (N_15883,N_10174,N_12906);
and U15884 (N_15884,N_11396,N_11797);
nor U15885 (N_15885,N_10169,N_13577);
nor U15886 (N_15886,N_12855,N_14490);
nor U15887 (N_15887,N_14720,N_13797);
xor U15888 (N_15888,N_11782,N_10690);
nand U15889 (N_15889,N_14452,N_14419);
or U15890 (N_15890,N_14442,N_14328);
nand U15891 (N_15891,N_13476,N_14988);
or U15892 (N_15892,N_13749,N_11980);
nor U15893 (N_15893,N_13276,N_14870);
or U15894 (N_15894,N_13104,N_13463);
and U15895 (N_15895,N_10637,N_13715);
nand U15896 (N_15896,N_11889,N_13082);
or U15897 (N_15897,N_14890,N_13111);
and U15898 (N_15898,N_14049,N_13796);
nor U15899 (N_15899,N_14956,N_12139);
nand U15900 (N_15900,N_10296,N_14934);
and U15901 (N_15901,N_13763,N_12799);
or U15902 (N_15902,N_11836,N_12546);
nor U15903 (N_15903,N_13468,N_12167);
xor U15904 (N_15904,N_12822,N_13628);
nand U15905 (N_15905,N_14667,N_10800);
and U15906 (N_15906,N_10672,N_14235);
nor U15907 (N_15907,N_14792,N_13988);
nand U15908 (N_15908,N_12145,N_13914);
nand U15909 (N_15909,N_12397,N_11497);
or U15910 (N_15910,N_13587,N_12018);
or U15911 (N_15911,N_11897,N_13669);
nand U15912 (N_15912,N_12345,N_14151);
or U15913 (N_15913,N_11394,N_13011);
and U15914 (N_15914,N_10483,N_13531);
nor U15915 (N_15915,N_11988,N_14488);
or U15916 (N_15916,N_10620,N_10001);
or U15917 (N_15917,N_12938,N_11252);
and U15918 (N_15918,N_10629,N_10973);
nor U15919 (N_15919,N_10144,N_11375);
or U15920 (N_15920,N_13784,N_13325);
nor U15921 (N_15921,N_11079,N_10298);
and U15922 (N_15922,N_13375,N_10409);
or U15923 (N_15923,N_12742,N_13213);
nand U15924 (N_15924,N_14660,N_12365);
nor U15925 (N_15925,N_10989,N_12890);
or U15926 (N_15926,N_11991,N_11372);
nor U15927 (N_15927,N_10897,N_11378);
and U15928 (N_15928,N_12660,N_10140);
and U15929 (N_15929,N_12847,N_13271);
or U15930 (N_15930,N_10125,N_10190);
nand U15931 (N_15931,N_11362,N_10734);
nand U15932 (N_15932,N_12469,N_12003);
nand U15933 (N_15933,N_14883,N_14067);
and U15934 (N_15934,N_14587,N_13366);
nor U15935 (N_15935,N_11059,N_12425);
xnor U15936 (N_15936,N_13627,N_10012);
and U15937 (N_15937,N_12247,N_10476);
and U15938 (N_15938,N_11891,N_10913);
and U15939 (N_15939,N_12863,N_11330);
or U15940 (N_15940,N_10816,N_12336);
nand U15941 (N_15941,N_10639,N_11398);
and U15942 (N_15942,N_11711,N_12120);
nand U15943 (N_15943,N_11146,N_14549);
nand U15944 (N_15944,N_10594,N_10780);
or U15945 (N_15945,N_13590,N_13066);
and U15946 (N_15946,N_10790,N_10922);
and U15947 (N_15947,N_11530,N_10525);
nand U15948 (N_15948,N_12770,N_13274);
or U15949 (N_15949,N_12960,N_12281);
nor U15950 (N_15950,N_12817,N_12222);
and U15951 (N_15951,N_13412,N_14368);
xor U15952 (N_15952,N_11668,N_14414);
nor U15953 (N_15953,N_14559,N_14892);
xnor U15954 (N_15954,N_11612,N_10026);
nor U15955 (N_15955,N_13242,N_10181);
xor U15956 (N_15956,N_11043,N_12350);
nor U15957 (N_15957,N_13544,N_13836);
xnor U15958 (N_15958,N_13391,N_13608);
nor U15959 (N_15959,N_11367,N_14504);
and U15960 (N_15960,N_12874,N_14278);
nor U15961 (N_15961,N_11193,N_13243);
and U15962 (N_15962,N_14099,N_14576);
nand U15963 (N_15963,N_12909,N_11901);
or U15964 (N_15964,N_14165,N_13220);
xor U15965 (N_15965,N_14856,N_13018);
nand U15966 (N_15966,N_13680,N_13722);
or U15967 (N_15967,N_13605,N_12989);
xnor U15968 (N_15968,N_12555,N_13237);
xor U15969 (N_15969,N_12035,N_12060);
nor U15970 (N_15970,N_13136,N_14911);
or U15971 (N_15971,N_12185,N_14284);
or U15972 (N_15972,N_13922,N_14565);
nand U15973 (N_15973,N_12739,N_14728);
and U15974 (N_15974,N_12974,N_13210);
nor U15975 (N_15975,N_11525,N_10779);
nor U15976 (N_15976,N_10671,N_14353);
and U15977 (N_15977,N_10856,N_13871);
nor U15978 (N_15978,N_14073,N_11743);
and U15979 (N_15979,N_10224,N_14329);
and U15980 (N_15980,N_14096,N_14185);
nor U15981 (N_15981,N_10496,N_10474);
nand U15982 (N_15982,N_10782,N_14657);
nand U15983 (N_15983,N_14648,N_10271);
nor U15984 (N_15984,N_14218,N_12727);
xnor U15985 (N_15985,N_10093,N_14775);
or U15986 (N_15986,N_14305,N_10885);
xnor U15987 (N_15987,N_13985,N_12173);
nand U15988 (N_15988,N_13792,N_11103);
nor U15989 (N_15989,N_13024,N_12603);
xnor U15990 (N_15990,N_14119,N_13655);
xor U15991 (N_15991,N_12889,N_11859);
nor U15992 (N_15992,N_13108,N_14351);
nor U15993 (N_15993,N_13487,N_12326);
nor U15994 (N_15994,N_13482,N_10139);
xor U15995 (N_15995,N_10531,N_13705);
nand U15996 (N_15996,N_12441,N_12743);
nor U15997 (N_15997,N_14193,N_12861);
nand U15998 (N_15998,N_14954,N_12542);
xor U15999 (N_15999,N_13756,N_11746);
xor U16000 (N_16000,N_12191,N_10669);
nand U16001 (N_16001,N_13870,N_14838);
and U16002 (N_16002,N_11258,N_12969);
nand U16003 (N_16003,N_14343,N_14243);
nor U16004 (N_16004,N_13405,N_12786);
nand U16005 (N_16005,N_13642,N_11868);
and U16006 (N_16006,N_10843,N_14357);
or U16007 (N_16007,N_12375,N_10512);
nand U16008 (N_16008,N_13408,N_13875);
nor U16009 (N_16009,N_14027,N_11708);
nor U16010 (N_16010,N_11091,N_14655);
and U16011 (N_16011,N_14471,N_10437);
nand U16012 (N_16012,N_12169,N_11360);
and U16013 (N_16013,N_13471,N_14680);
nor U16014 (N_16014,N_12760,N_10194);
nand U16015 (N_16015,N_14383,N_12854);
nand U16016 (N_16016,N_10933,N_11918);
or U16017 (N_16017,N_14802,N_10361);
xnor U16018 (N_16018,N_14072,N_14738);
xnor U16019 (N_16019,N_10200,N_12399);
or U16020 (N_16020,N_14964,N_14279);
nor U16021 (N_16021,N_11878,N_10633);
or U16022 (N_16022,N_13898,N_14696);
or U16023 (N_16023,N_12632,N_11235);
xor U16024 (N_16024,N_10159,N_13451);
nand U16025 (N_16025,N_13899,N_12883);
or U16026 (N_16026,N_12643,N_12444);
or U16027 (N_16027,N_11724,N_12330);
nor U16028 (N_16028,N_14267,N_10344);
and U16029 (N_16029,N_11739,N_11336);
or U16030 (N_16030,N_13300,N_14798);
and U16031 (N_16031,N_10357,N_10069);
xnor U16032 (N_16032,N_13097,N_10310);
and U16033 (N_16033,N_13602,N_13905);
and U16034 (N_16034,N_13356,N_13385);
or U16035 (N_16035,N_11643,N_12052);
and U16036 (N_16036,N_10492,N_10636);
nand U16037 (N_16037,N_14645,N_11038);
or U16038 (N_16038,N_10152,N_10646);
nand U16039 (N_16039,N_14949,N_13873);
nand U16040 (N_16040,N_10950,N_12675);
nand U16041 (N_16041,N_13184,N_10457);
xor U16042 (N_16042,N_12160,N_12184);
or U16043 (N_16043,N_11228,N_14509);
and U16044 (N_16044,N_14946,N_13152);
xor U16045 (N_16045,N_10937,N_13187);
or U16046 (N_16046,N_13511,N_14796);
or U16047 (N_16047,N_14900,N_10888);
nor U16048 (N_16048,N_14405,N_14907);
or U16049 (N_16049,N_10979,N_14069);
nand U16050 (N_16050,N_11656,N_12837);
or U16051 (N_16051,N_11063,N_11523);
or U16052 (N_16052,N_10045,N_13637);
and U16053 (N_16053,N_14965,N_11455);
and U16054 (N_16054,N_10248,N_14979);
and U16055 (N_16055,N_12420,N_12567);
and U16056 (N_16056,N_13037,N_13803);
and U16057 (N_16057,N_13636,N_14106);
nand U16058 (N_16058,N_12655,N_13113);
nor U16059 (N_16059,N_10062,N_13665);
and U16060 (N_16060,N_11207,N_14601);
nand U16061 (N_16061,N_13539,N_13115);
nand U16062 (N_16062,N_14771,N_13527);
and U16063 (N_16063,N_11411,N_11696);
nand U16064 (N_16064,N_11225,N_14582);
or U16065 (N_16065,N_14059,N_10087);
and U16066 (N_16066,N_11644,N_11471);
nor U16067 (N_16067,N_13675,N_14520);
nand U16068 (N_16068,N_10043,N_10197);
nor U16069 (N_16069,N_14515,N_11865);
nor U16070 (N_16070,N_13693,N_14523);
nand U16071 (N_16071,N_13240,N_13304);
nand U16072 (N_16072,N_12732,N_14009);
and U16073 (N_16073,N_11649,N_12462);
or U16074 (N_16074,N_11481,N_12344);
nand U16075 (N_16075,N_11911,N_10982);
nor U16076 (N_16076,N_14708,N_11319);
or U16077 (N_16077,N_13295,N_14568);
or U16078 (N_16078,N_12037,N_11508);
nor U16079 (N_16079,N_10265,N_10643);
and U16080 (N_16080,N_12489,N_10801);
or U16081 (N_16081,N_10815,N_11197);
nor U16082 (N_16082,N_12213,N_13045);
or U16083 (N_16083,N_10903,N_14293);
nand U16084 (N_16084,N_10908,N_11400);
nor U16085 (N_16085,N_12970,N_10371);
or U16086 (N_16086,N_13932,N_11960);
or U16087 (N_16087,N_14692,N_13966);
and U16088 (N_16088,N_11722,N_12672);
nand U16089 (N_16089,N_10086,N_14943);
and U16090 (N_16090,N_12225,N_13747);
and U16091 (N_16091,N_11489,N_11729);
or U16092 (N_16092,N_11482,N_13445);
or U16093 (N_16093,N_11098,N_10960);
nor U16094 (N_16094,N_10487,N_12616);
xnor U16095 (N_16095,N_11826,N_10890);
and U16096 (N_16096,N_14695,N_13312);
nand U16097 (N_16097,N_10998,N_10282);
and U16098 (N_16098,N_11634,N_11731);
and U16099 (N_16099,N_11526,N_12870);
and U16100 (N_16100,N_11949,N_12778);
or U16101 (N_16101,N_10983,N_11159);
or U16102 (N_16102,N_10747,N_10814);
and U16103 (N_16103,N_11418,N_11682);
or U16104 (N_16104,N_14148,N_13461);
nand U16105 (N_16105,N_12450,N_14153);
nor U16106 (N_16106,N_14319,N_14972);
nor U16107 (N_16107,N_14619,N_11348);
nand U16108 (N_16108,N_12263,N_14697);
and U16109 (N_16109,N_14675,N_14344);
nor U16110 (N_16110,N_13891,N_10543);
and U16111 (N_16111,N_14208,N_11260);
nor U16112 (N_16112,N_10413,N_10367);
nand U16113 (N_16113,N_13183,N_13791);
or U16114 (N_16114,N_13267,N_12945);
xnor U16115 (N_16115,N_13269,N_12759);
or U16116 (N_16116,N_10552,N_10031);
or U16117 (N_16117,N_13344,N_12107);
and U16118 (N_16118,N_10446,N_13034);
nor U16119 (N_16119,N_13674,N_13231);
or U16120 (N_16120,N_11535,N_10769);
or U16121 (N_16121,N_14346,N_10591);
xor U16122 (N_16122,N_14663,N_12991);
and U16123 (N_16123,N_14608,N_11104);
and U16124 (N_16124,N_12401,N_11148);
nor U16125 (N_16125,N_13822,N_13545);
or U16126 (N_16126,N_12795,N_11132);
nand U16127 (N_16127,N_13311,N_10279);
and U16128 (N_16128,N_14849,N_14128);
nor U16129 (N_16129,N_11293,N_11593);
nand U16130 (N_16130,N_12163,N_12914);
nand U16131 (N_16131,N_12994,N_13696);
nor U16132 (N_16132,N_13785,N_14213);
nand U16133 (N_16133,N_14562,N_11441);
or U16134 (N_16134,N_10631,N_13176);
nand U16135 (N_16135,N_11304,N_12372);
or U16136 (N_16136,N_12488,N_12366);
and U16137 (N_16137,N_10727,N_14228);
xnor U16138 (N_16138,N_12762,N_12448);
and U16139 (N_16139,N_11688,N_11872);
nor U16140 (N_16140,N_10616,N_10966);
or U16141 (N_16141,N_11531,N_11380);
xor U16142 (N_16142,N_14350,N_12237);
nand U16143 (N_16143,N_13403,N_11979);
nor U16144 (N_16144,N_10238,N_13096);
nand U16145 (N_16145,N_13308,N_14600);
nor U16146 (N_16146,N_13917,N_14078);
nand U16147 (N_16147,N_13484,N_14215);
nor U16148 (N_16148,N_12506,N_12919);
nor U16149 (N_16149,N_11147,N_11205);
nand U16150 (N_16150,N_12332,N_10288);
nor U16151 (N_16151,N_11707,N_11985);
or U16152 (N_16152,N_11493,N_12031);
nor U16153 (N_16153,N_14527,N_14552);
and U16154 (N_16154,N_12287,N_11272);
or U16155 (N_16155,N_11740,N_12558);
and U16156 (N_16156,N_11514,N_11638);
nand U16157 (N_16157,N_10249,N_10134);
nand U16158 (N_16158,N_12177,N_12202);
or U16159 (N_16159,N_11744,N_13936);
nor U16160 (N_16160,N_14538,N_14431);
nor U16161 (N_16161,N_12552,N_10862);
and U16162 (N_16162,N_11590,N_12370);
xnor U16163 (N_16163,N_13721,N_10762);
xnor U16164 (N_16164,N_14101,N_10051);
and U16165 (N_16165,N_10198,N_11735);
or U16166 (N_16166,N_12700,N_11355);
nor U16167 (N_16167,N_14994,N_12361);
nand U16168 (N_16168,N_14745,N_13757);
and U16169 (N_16169,N_14925,N_11808);
nand U16170 (N_16170,N_10701,N_11594);
and U16171 (N_16171,N_10961,N_10201);
nand U16172 (N_16172,N_13837,N_13017);
nor U16173 (N_16173,N_14336,N_14214);
nor U16174 (N_16174,N_13206,N_10187);
nor U16175 (N_16175,N_13331,N_10186);
or U16176 (N_16176,N_12200,N_12528);
nor U16177 (N_16177,N_14493,N_14832);
xnor U16178 (N_16178,N_10307,N_13342);
or U16179 (N_16179,N_14376,N_14952);
or U16180 (N_16180,N_14995,N_12917);
xor U16181 (N_16181,N_11326,N_10220);
and U16182 (N_16182,N_14260,N_14385);
nor U16183 (N_16183,N_10013,N_12134);
or U16184 (N_16184,N_10462,N_10822);
nor U16185 (N_16185,N_12757,N_10582);
or U16186 (N_16186,N_13737,N_12186);
xor U16187 (N_16187,N_13143,N_14602);
or U16188 (N_16188,N_14071,N_11386);
nor U16189 (N_16189,N_12792,N_11383);
nand U16190 (N_16190,N_12417,N_12252);
nor U16191 (N_16191,N_14542,N_10597);
or U16192 (N_16192,N_12597,N_13094);
or U16193 (N_16193,N_10579,N_13431);
or U16194 (N_16194,N_13146,N_11311);
nor U16195 (N_16195,N_14324,N_14689);
or U16196 (N_16196,N_14123,N_12691);
or U16197 (N_16197,N_12443,N_14381);
nor U16198 (N_16198,N_11288,N_11119);
or U16199 (N_16199,N_13573,N_10101);
and U16200 (N_16200,N_13029,N_14330);
nor U16201 (N_16201,N_11726,N_13986);
or U16202 (N_16202,N_14641,N_12463);
xnor U16203 (N_16203,N_12079,N_11730);
and U16204 (N_16204,N_11220,N_13687);
and U16205 (N_16205,N_11012,N_11276);
nor U16206 (N_16206,N_14916,N_11597);
or U16207 (N_16207,N_10274,N_14772);
or U16208 (N_16208,N_11609,N_13351);
nand U16209 (N_16209,N_12618,N_11860);
and U16210 (N_16210,N_10486,N_11908);
and U16211 (N_16211,N_12467,N_14617);
or U16212 (N_16212,N_11241,N_10110);
or U16213 (N_16213,N_14453,N_10118);
nand U16214 (N_16214,N_13456,N_13341);
or U16215 (N_16215,N_10124,N_13318);
nand U16216 (N_16216,N_12334,N_12470);
nand U16217 (N_16217,N_11685,N_14481);
nor U16218 (N_16218,N_13863,N_12013);
or U16219 (N_16219,N_10217,N_11592);
nand U16220 (N_16220,N_13827,N_11734);
nor U16221 (N_16221,N_11845,N_14024);
or U16222 (N_16222,N_11403,N_13916);
nor U16223 (N_16223,N_11693,N_13739);
or U16224 (N_16224,N_13810,N_12564);
or U16225 (N_16225,N_11655,N_14202);
or U16226 (N_16226,N_12308,N_11520);
nor U16227 (N_16227,N_12199,N_11214);
or U16228 (N_16228,N_11226,N_12258);
nand U16229 (N_16229,N_11125,N_10054);
nand U16230 (N_16230,N_11773,N_14879);
nor U16231 (N_16231,N_14021,N_10267);
or U16232 (N_16232,N_11389,N_14282);
and U16233 (N_16233,N_12887,N_13910);
and U16234 (N_16234,N_12499,N_14211);
nor U16235 (N_16235,N_14841,N_12218);
nor U16236 (N_16236,N_13735,N_13772);
xor U16237 (N_16237,N_11614,N_12624);
nor U16238 (N_16238,N_11393,N_14525);
nand U16239 (N_16239,N_14642,N_14459);
and U16240 (N_16240,N_12808,N_10875);
or U16241 (N_16241,N_13751,N_14544);
nor U16242 (N_16242,N_10799,N_13490);
nand U16243 (N_16243,N_10231,N_13338);
nand U16244 (N_16244,N_14732,N_10574);
nand U16245 (N_16245,N_14583,N_10562);
or U16246 (N_16246,N_11580,N_11082);
or U16247 (N_16247,N_10388,N_10188);
and U16248 (N_16248,N_12961,N_10128);
nand U16249 (N_16249,N_12504,N_13395);
nand U16250 (N_16250,N_14698,N_14217);
and U16251 (N_16251,N_13938,N_14275);
or U16252 (N_16252,N_11126,N_11516);
nor U16253 (N_16253,N_11838,N_12866);
and U16254 (N_16254,N_11954,N_14846);
nand U16255 (N_16255,N_13139,N_14229);
or U16256 (N_16256,N_13460,N_12654);
or U16257 (N_16257,N_10401,N_14733);
and U16258 (N_16258,N_14413,N_12102);
or U16259 (N_16259,N_14141,N_12067);
nand U16260 (N_16260,N_11215,N_13459);
and U16261 (N_16261,N_14364,N_11295);
nor U16262 (N_16262,N_12192,N_10651);
or U16263 (N_16263,N_12181,N_10941);
nand U16264 (N_16264,N_10389,N_10748);
and U16265 (N_16265,N_13724,N_14574);
nor U16266 (N_16266,N_14271,N_10898);
nand U16267 (N_16267,N_13673,N_12446);
xor U16268 (N_16268,N_12205,N_14505);
and U16269 (N_16269,N_11769,N_14192);
nor U16270 (N_16270,N_11736,N_11443);
nand U16271 (N_16271,N_12349,N_13428);
or U16272 (N_16272,N_10286,N_11204);
xnor U16273 (N_16273,N_13979,N_13069);
nand U16274 (N_16274,N_10106,N_11927);
and U16275 (N_16275,N_13315,N_13198);
nand U16276 (N_16276,N_12838,N_10306);
nand U16277 (N_16277,N_10325,N_13616);
nor U16278 (N_16278,N_13555,N_13065);
and U16279 (N_16279,N_14570,N_12501);
nor U16280 (N_16280,N_12750,N_12996);
nor U16281 (N_16281,N_12775,N_10882);
and U16282 (N_16282,N_10293,N_13821);
xnor U16283 (N_16283,N_10944,N_12747);
or U16284 (N_16284,N_10426,N_12293);
or U16285 (N_16285,N_12777,N_13808);
or U16286 (N_16286,N_10433,N_14593);
xor U16287 (N_16287,N_13671,N_11294);
xor U16288 (N_16288,N_11473,N_10776);
nand U16289 (N_16289,N_14711,N_10059);
nor U16290 (N_16290,N_14597,N_13689);
nand U16291 (N_16291,N_11557,N_14590);
nor U16292 (N_16292,N_10613,N_13346);
or U16293 (N_16293,N_14223,N_14302);
or U16294 (N_16294,N_14085,N_14094);
or U16295 (N_16295,N_12439,N_13421);
nor U16296 (N_16296,N_10638,N_12692);
nand U16297 (N_16297,N_13725,N_11070);
and U16298 (N_16298,N_12126,N_12785);
nand U16299 (N_16299,N_14320,N_11349);
and U16300 (N_16300,N_14882,N_10987);
or U16301 (N_16301,N_13854,N_13275);
nor U16302 (N_16302,N_10342,N_13416);
xor U16303 (N_16303,N_11841,N_13600);
nor U16304 (N_16304,N_10423,N_10698);
and U16305 (N_16305,N_12327,N_13019);
nor U16306 (N_16306,N_11575,N_12421);
nand U16307 (N_16307,N_11713,N_11081);
and U16308 (N_16308,N_10901,N_10154);
xnor U16309 (N_16309,N_12403,N_14068);
and U16310 (N_16310,N_13533,N_12115);
and U16311 (N_16311,N_12055,N_11242);
and U16312 (N_16312,N_11322,N_13246);
nand U16313 (N_16313,N_13402,N_11842);
and U16314 (N_16314,N_13816,N_10015);
or U16315 (N_16315,N_14703,N_13497);
nand U16316 (N_16316,N_12900,N_14981);
nand U16317 (N_16317,N_12977,N_10736);
and U16318 (N_16318,N_14458,N_11947);
or U16319 (N_16319,N_12609,N_10151);
or U16320 (N_16320,N_10006,N_10925);
or U16321 (N_16321,N_12161,N_11567);
and U16322 (N_16322,N_11828,N_12093);
nand U16323 (N_16323,N_10252,N_12452);
nand U16324 (N_16324,N_11399,N_14460);
nor U16325 (N_16325,N_14129,N_11364);
or U16326 (N_16326,N_14465,N_14316);
nand U16327 (N_16327,N_11732,N_11527);
nand U16328 (N_16328,N_12189,N_10316);
and U16329 (N_16329,N_13201,N_11499);
xor U16330 (N_16330,N_13766,N_13990);
nor U16331 (N_16331,N_13815,N_10676);
xnor U16332 (N_16332,N_14586,N_10033);
xor U16333 (N_16333,N_12767,N_10219);
or U16334 (N_16334,N_13148,N_11329);
nor U16335 (N_16335,N_10918,N_12373);
or U16336 (N_16336,N_14866,N_12081);
nor U16337 (N_16337,N_13894,N_13477);
nand U16338 (N_16338,N_11141,N_14056);
nand U16339 (N_16339,N_13830,N_12203);
nand U16340 (N_16340,N_13061,N_10517);
and U16341 (N_16341,N_14788,N_14561);
and U16342 (N_16342,N_14437,N_14269);
or U16343 (N_16343,N_10537,N_11719);
nand U16344 (N_16344,N_13138,N_11379);
nand U16345 (N_16345,N_11353,N_10256);
nand U16346 (N_16346,N_11468,N_12894);
nand U16347 (N_16347,N_11990,N_10757);
and U16348 (N_16348,N_14299,N_14533);
nor U16349 (N_16349,N_10004,N_13465);
nor U16350 (N_16350,N_14345,N_14076);
and U16351 (N_16351,N_10275,N_12329);
nor U16352 (N_16352,N_13320,N_11853);
and U16353 (N_16353,N_14743,N_14536);
and U16354 (N_16354,N_13880,N_12587);
or U16355 (N_16355,N_12836,N_10337);
xor U16356 (N_16356,N_11912,N_13010);
nand U16357 (N_16357,N_10835,N_10255);
nor U16358 (N_16358,N_14494,N_13132);
or U16359 (N_16359,N_10185,N_14919);
or U16360 (N_16360,N_10347,N_12431);
and U16361 (N_16361,N_11431,N_13158);
nor U16362 (N_16362,N_11438,N_14323);
or U16363 (N_16363,N_13419,N_13874);
or U16364 (N_16364,N_11804,N_10705);
nand U16365 (N_16365,N_10142,N_10244);
and U16366 (N_16366,N_10569,N_10521);
or U16367 (N_16367,N_12821,N_14075);
nand U16368 (N_16368,N_13164,N_11659);
or U16369 (N_16369,N_14820,N_12599);
nor U16370 (N_16370,N_11637,N_14348);
nor U16371 (N_16371,N_12815,N_14335);
and U16372 (N_16372,N_13438,N_13526);
xor U16373 (N_16373,N_10917,N_14803);
nor U16374 (N_16374,N_13170,N_14152);
nand U16375 (N_16375,N_11071,N_12364);
nand U16376 (N_16376,N_11502,N_10085);
or U16377 (N_16377,N_10513,N_13771);
nand U16378 (N_16378,N_14836,N_12008);
nor U16379 (N_16379,N_14970,N_12878);
xnor U16380 (N_16380,N_12477,N_13598);
nor U16381 (N_16381,N_12032,N_13050);
xor U16382 (N_16382,N_12539,N_11727);
nand U16383 (N_16383,N_14135,N_14463);
nor U16384 (N_16384,N_11206,N_10729);
nand U16385 (N_16385,N_11345,N_11585);
nor U16386 (N_16386,N_14822,N_10700);
and U16387 (N_16387,N_12508,N_13462);
nand U16388 (N_16388,N_10829,N_12290);
or U16389 (N_16389,N_13996,N_13089);
nor U16390 (N_16390,N_11212,N_14629);
nand U16391 (N_16391,N_10760,N_11264);
and U16392 (N_16392,N_12318,N_12288);
nor U16393 (N_16393,N_14869,N_11737);
or U16394 (N_16394,N_11725,N_12956);
nor U16395 (N_16395,N_11588,N_11890);
nor U16396 (N_16396,N_10247,N_10615);
nor U16397 (N_16397,N_11581,N_11180);
nand U16398 (N_16398,N_12818,N_14179);
nand U16399 (N_16399,N_14404,N_12435);
nand U16400 (N_16400,N_12717,N_14038);
or U16401 (N_16401,N_10311,N_12105);
nor U16402 (N_16402,N_14425,N_13859);
and U16403 (N_16403,N_11002,N_13548);
nor U16404 (N_16404,N_12369,N_11667);
or U16405 (N_16405,N_13740,N_10689);
or U16406 (N_16406,N_14112,N_11110);
nor U16407 (N_16407,N_11833,N_10884);
nor U16408 (N_16408,N_14948,N_10345);
nor U16409 (N_16409,N_12647,N_11953);
or U16410 (N_16410,N_10208,N_11822);
nand U16411 (N_16411,N_13454,N_14790);
xnor U16412 (N_16412,N_10809,N_12913);
nor U16413 (N_16413,N_14451,N_14310);
nor U16414 (N_16414,N_14694,N_11371);
and U16415 (N_16415,N_12824,N_12988);
and U16416 (N_16416,N_14647,N_11406);
or U16417 (N_16417,N_12352,N_11328);
xor U16418 (N_16418,N_14764,N_11951);
nor U16419 (N_16419,N_11978,N_10910);
nand U16420 (N_16420,N_11675,N_13222);
nand U16421 (N_16421,N_11033,N_14932);
or U16422 (N_16422,N_14379,N_11576);
nor U16423 (N_16423,N_10260,N_14150);
nand U16424 (N_16424,N_13754,N_12845);
or U16425 (N_16425,N_10604,N_10259);
nor U16426 (N_16426,N_11290,N_14416);
and U16427 (N_16427,N_14050,N_11429);
nand U16428 (N_16428,N_13444,N_11428);
nand U16429 (N_16429,N_12130,N_11624);
nand U16430 (N_16430,N_13620,N_12531);
nor U16431 (N_16431,N_12714,N_11950);
and U16432 (N_16432,N_12239,N_14789);
and U16433 (N_16433,N_10784,N_10906);
nor U16434 (N_16434,N_14976,N_11281);
or U16435 (N_16435,N_12801,N_13543);
and U16436 (N_16436,N_10160,N_12652);
or U16437 (N_16437,N_11285,N_14669);
nand U16438 (N_16438,N_12661,N_11075);
and U16439 (N_16439,N_10534,N_11536);
and U16440 (N_16440,N_13770,N_11747);
nand U16441 (N_16441,N_10902,N_11538);
and U16442 (N_16442,N_10564,N_12086);
and U16443 (N_16443,N_12068,N_13819);
nor U16444 (N_16444,N_11450,N_10035);
nor U16445 (N_16445,N_14121,N_14734);
xor U16446 (N_16446,N_13805,N_10704);
nor U16447 (N_16447,N_14691,N_12895);
or U16448 (N_16448,N_14848,N_14674);
and U16449 (N_16449,N_11442,N_11173);
and U16450 (N_16450,N_13947,N_11540);
nor U16451 (N_16451,N_12391,N_13982);
or U16452 (N_16452,N_14958,N_10977);
or U16453 (N_16453,N_13744,N_13663);
or U16454 (N_16454,N_13141,N_12626);
and U16455 (N_16455,N_12179,N_11790);
nand U16456 (N_16456,N_14831,N_13254);
and U16457 (N_16457,N_11622,N_14156);
and U16458 (N_16458,N_13697,N_13977);
nand U16459 (N_16459,N_13339,N_14611);
or U16460 (N_16460,N_10261,N_12541);
or U16461 (N_16461,N_14245,N_10584);
or U16462 (N_16462,N_11275,N_12314);
nor U16463 (N_16463,N_10017,N_12781);
nand U16464 (N_16464,N_11449,N_12920);
or U16465 (N_16465,N_14434,N_11036);
and U16466 (N_16466,N_11023,N_13179);
and U16467 (N_16467,N_13750,N_13557);
nor U16468 (N_16468,N_13133,N_13904);
nor U16469 (N_16469,N_14749,N_14089);
nand U16470 (N_16470,N_10336,N_10405);
nor U16471 (N_16471,N_10165,N_11495);
nand U16472 (N_16472,N_11974,N_14904);
nand U16473 (N_16473,N_14002,N_10381);
nor U16474 (N_16474,N_12229,N_10327);
or U16475 (N_16475,N_13779,N_14742);
nor U16476 (N_16476,N_12445,N_14513);
xor U16477 (N_16477,N_13997,N_10892);
and U16478 (N_16478,N_11922,N_13354);
and U16479 (N_16479,N_10313,N_10126);
nand U16480 (N_16480,N_12523,N_12136);
nor U16481 (N_16481,N_13047,N_14224);
and U16482 (N_16482,N_14665,N_11582);
nand U16483 (N_16483,N_14426,N_14821);
nand U16484 (N_16484,N_14815,N_14872);
and U16485 (N_16485,N_10387,N_13392);
nand U16486 (N_16486,N_11325,N_11162);
and U16487 (N_16487,N_12825,N_14210);
and U16488 (N_16488,N_10292,N_12810);
nand U16489 (N_16489,N_11391,N_14170);
nand U16490 (N_16490,N_12707,N_14019);
and U16491 (N_16491,N_14103,N_14200);
or U16492 (N_16492,N_13552,N_10911);
nor U16493 (N_16493,N_14446,N_14818);
nand U16494 (N_16494,N_11881,N_12241);
or U16495 (N_16495,N_13812,N_12317);
nand U16496 (N_16496,N_14164,N_12429);
or U16497 (N_16497,N_14769,N_12648);
or U16498 (N_16498,N_14810,N_13418);
and U16499 (N_16499,N_11327,N_14181);
nand U16500 (N_16500,N_10940,N_12740);
nor U16501 (N_16501,N_12982,N_12015);
nor U16502 (N_16502,N_10838,N_14083);
or U16503 (N_16503,N_10746,N_14677);
nor U16504 (N_16504,N_14635,N_14853);
or U16505 (N_16505,N_10825,N_12698);
nor U16506 (N_16506,N_10459,N_14813);
or U16507 (N_16507,N_12638,N_11521);
and U16508 (N_16508,N_11888,N_11477);
and U16509 (N_16509,N_14805,N_14240);
xnor U16510 (N_16510,N_11935,N_12457);
nor U16511 (N_16511,N_10153,N_12482);
nand U16512 (N_16512,N_13257,N_14154);
or U16513 (N_16513,N_11500,N_14173);
and U16514 (N_16514,N_13003,N_12264);
nor U16515 (N_16515,N_11334,N_10499);
nand U16516 (N_16516,N_12170,N_14809);
nor U16517 (N_16517,N_13592,N_13524);
nand U16518 (N_16518,N_12583,N_11652);
or U16519 (N_16519,N_13710,N_10119);
nand U16520 (N_16520,N_11229,N_11463);
or U16521 (N_16521,N_11317,N_11026);
nor U16522 (N_16522,N_13251,N_13127);
or U16523 (N_16523,N_14712,N_13289);
and U16524 (N_16524,N_13475,N_14186);
nor U16525 (N_16525,N_13348,N_10554);
or U16526 (N_16526,N_13727,N_11824);
nor U16527 (N_16527,N_12589,N_14545);
and U16528 (N_16528,N_13114,N_11357);
or U16529 (N_16529,N_12897,N_11819);
nor U16530 (N_16530,N_12885,N_12240);
or U16531 (N_16531,N_12083,N_13229);
xnor U16532 (N_16532,N_14760,N_14980);
nor U16533 (N_16533,N_10400,N_12826);
xor U16534 (N_16534,N_13518,N_14195);
nor U16535 (N_16535,N_14744,N_11177);
nand U16536 (N_16536,N_13442,N_11342);
or U16537 (N_16537,N_12302,N_11097);
nand U16538 (N_16538,N_13888,N_14133);
nor U16539 (N_16539,N_13105,N_14585);
or U16540 (N_16540,N_10466,N_13093);
nand U16541 (N_16541,N_13058,N_11435);
or U16542 (N_16542,N_11213,N_13420);
or U16543 (N_16543,N_13448,N_11905);
and U16544 (N_16544,N_12763,N_12376);
nand U16545 (N_16545,N_10874,N_10379);
nand U16546 (N_16546,N_11528,N_12725);
nor U16547 (N_16547,N_13559,N_12066);
nor U16548 (N_16548,N_11440,N_14355);
nor U16549 (N_16549,N_13886,N_14365);
and U16550 (N_16550,N_11568,N_11020);
nor U16551 (N_16551,N_14125,N_13264);
nand U16552 (N_16552,N_10172,N_10624);
and U16553 (N_16553,N_14389,N_12515);
or U16554 (N_16554,N_11992,N_13337);
or U16555 (N_16555,N_14378,N_13447);
and U16556 (N_16556,N_11263,N_13850);
and U16557 (N_16557,N_14960,N_13882);
nand U16558 (N_16558,N_13215,N_11662);
nor U16559 (N_16559,N_12578,N_10587);
nor U16560 (N_16560,N_14518,N_11679);
and U16561 (N_16561,N_10945,N_11683);
and U16562 (N_16562,N_11287,N_10439);
nand U16563 (N_16563,N_12519,N_12166);
or U16564 (N_16564,N_12260,N_13672);
nor U16565 (N_16565,N_10821,N_12802);
and U16566 (N_16566,N_11558,N_13266);
or U16567 (N_16567,N_14197,N_14785);
nor U16568 (N_16568,N_14999,N_12020);
nand U16569 (N_16569,N_14506,N_12574);
and U16570 (N_16570,N_13159,N_13083);
nand U16571 (N_16571,N_14750,N_11250);
nand U16572 (N_16572,N_10978,N_11138);
or U16573 (N_16573,N_12064,N_10210);
and U16574 (N_16574,N_12737,N_13185);
and U16575 (N_16575,N_12353,N_11480);
and U16576 (N_16576,N_10980,N_11895);
nand U16577 (N_16577,N_14987,N_11995);
and U16578 (N_16578,N_12046,N_11965);
or U16579 (N_16579,N_10810,N_11723);
nor U16580 (N_16580,N_10329,N_10934);
or U16581 (N_16581,N_11765,N_12857);
nand U16582 (N_16582,N_13769,N_12613);
nand U16583 (N_16583,N_12125,N_13434);
and U16584 (N_16584,N_10205,N_11981);
nor U16585 (N_16585,N_13564,N_11433);
xnor U16586 (N_16586,N_12875,N_14762);
nand U16587 (N_16587,N_10955,N_10786);
nand U16588 (N_16588,N_14903,N_11191);
and U16589 (N_16589,N_12844,N_14830);
nand U16590 (N_16590,N_14126,N_14476);
xnor U16591 (N_16591,N_12952,N_12623);
or U16592 (N_16592,N_13046,N_13957);
and U16593 (N_16593,N_12227,N_14748);
or U16594 (N_16594,N_13291,N_13505);
xor U16595 (N_16595,N_11085,N_14921);
or U16596 (N_16596,N_12659,N_12529);
nor U16597 (N_16597,N_13753,N_13002);
nand U16598 (N_16598,N_13373,N_14926);
nor U16599 (N_16599,N_12761,N_11359);
nand U16600 (N_16600,N_13466,N_12262);
nor U16601 (N_16601,N_14833,N_14930);
nor U16602 (N_16602,N_12721,N_10503);
nand U16603 (N_16603,N_10959,N_14104);
or U16604 (N_16604,N_14120,N_12368);
nor U16605 (N_16605,N_11775,N_13793);
or U16606 (N_16606,N_12099,N_14678);
or U16607 (N_16607,N_11351,N_14707);
nand U16608 (N_16608,N_14845,N_13860);
nand U16609 (N_16609,N_11774,N_14620);
or U16610 (N_16610,N_10628,N_11529);
nor U16611 (N_16611,N_11152,N_13301);
xnor U16612 (N_16612,N_14395,N_10092);
nor U16613 (N_16613,N_12512,N_13426);
nand U16614 (N_16614,N_11169,N_13594);
nor U16615 (N_16615,N_14044,N_13629);
and U16616 (N_16616,N_10479,N_10609);
nand U16617 (N_16617,N_10488,N_11096);
nand U16618 (N_16618,N_11374,N_10312);
and U16619 (N_16619,N_13818,N_14410);
or U16620 (N_16620,N_12286,N_14725);
nand U16621 (N_16621,N_12347,N_14812);
or U16622 (N_16622,N_11114,N_10524);
and U16623 (N_16623,N_11601,N_11669);
and U16624 (N_16624,N_13166,N_11346);
and U16625 (N_16625,N_12765,N_14014);
nor U16626 (N_16626,N_14991,N_11297);
nand U16627 (N_16627,N_13352,N_13676);
or U16628 (N_16628,N_14012,N_11604);
or U16629 (N_16629,N_11616,N_13806);
nor U16630 (N_16630,N_13528,N_12915);
nor U16631 (N_16631,N_10916,N_13849);
or U16632 (N_16632,N_11831,N_11486);
or U16633 (N_16633,N_10869,N_12536);
or U16634 (N_16634,N_14449,N_12455);
or U16635 (N_16635,N_10320,N_12476);
xor U16636 (N_16636,N_12357,N_14023);
nand U16637 (N_16637,N_10002,N_14778);
nand U16638 (N_16638,N_12676,N_10396);
and U16639 (N_16639,N_10411,N_14605);
and U16640 (N_16640,N_10921,N_11053);
or U16641 (N_16641,N_13449,N_11886);
or U16642 (N_16642,N_14801,N_11401);
nor U16643 (N_16643,N_10067,N_12936);
or U16644 (N_16644,N_14309,N_13745);
nor U16645 (N_16645,N_10452,N_12063);
and U16646 (N_16646,N_13610,N_10105);
or U16647 (N_16647,N_10715,N_12518);
nor U16648 (N_16648,N_13981,N_12075);
nor U16649 (N_16649,N_14016,N_14191);
nor U16650 (N_16650,N_11202,N_12748);
and U16651 (N_16651,N_11923,N_12754);
and U16652 (N_16652,N_11034,N_10965);
nor U16653 (N_16653,N_10839,N_13078);
or U16654 (N_16654,N_10877,N_13887);
nor U16655 (N_16655,N_12550,N_10242);
nor U16656 (N_16656,N_12611,N_10149);
nand U16657 (N_16657,N_12029,N_10935);
nand U16658 (N_16658,N_13333,N_11305);
nand U16659 (N_16659,N_13726,N_10340);
or U16660 (N_16660,N_14373,N_14786);
or U16661 (N_16661,N_11462,N_13881);
xor U16662 (N_16662,N_13279,N_12323);
nand U16663 (N_16663,N_12696,N_12791);
and U16664 (N_16664,N_13036,N_12338);
xor U16665 (N_16665,N_12954,N_13223);
and U16666 (N_16666,N_13457,N_11133);
nor U16667 (N_16667,N_12881,N_12073);
nor U16668 (N_16668,N_14850,N_12695);
nor U16669 (N_16669,N_11422,N_13056);
xor U16670 (N_16670,N_12207,N_10301);
nor U16671 (N_16671,N_11035,N_11088);
and U16672 (N_16672,N_11283,N_13174);
nand U16673 (N_16673,N_10538,N_12333);
and U16674 (N_16674,N_13568,N_11758);
and U16675 (N_16675,N_14334,N_11240);
xnor U16676 (N_16676,N_12646,N_11646);
nor U16677 (N_16677,N_13826,N_12591);
and U16678 (N_16678,N_12843,N_10480);
nand U16679 (N_16679,N_12934,N_12662);
nand U16680 (N_16680,N_11332,N_13949);
and U16681 (N_16681,N_11791,N_12995);
or U16682 (N_16682,N_13380,N_10778);
and U16683 (N_16683,N_11247,N_10263);
or U16684 (N_16684,N_13195,N_12487);
nand U16685 (N_16685,N_13353,N_10751);
nor U16686 (N_16686,N_14877,N_13992);
xnor U16687 (N_16687,N_12392,N_12028);
nor U16688 (N_16688,N_12014,N_11381);
nor U16689 (N_16689,N_12188,N_10912);
or U16690 (N_16690,N_14475,N_14543);
or U16691 (N_16691,N_11792,N_12726);
nor U16692 (N_16692,N_10872,N_13782);
or U16693 (N_16693,N_13328,N_14406);
or U16694 (N_16694,N_12713,N_12588);
or U16695 (N_16695,N_13900,N_10061);
or U16696 (N_16696,N_11113,N_14109);
nor U16697 (N_16697,N_14633,N_13833);
nand U16698 (N_16698,N_10682,N_12807);
nand U16699 (N_16699,N_12442,N_11028);
or U16700 (N_16700,N_11286,N_11608);
and U16701 (N_16701,N_11689,N_10236);
or U16702 (N_16702,N_10566,N_11916);
nand U16703 (N_16703,N_13102,N_13109);
nand U16704 (N_16704,N_12484,N_13208);
or U16705 (N_16705,N_11850,N_12415);
nand U16706 (N_16706,N_10953,N_12407);
or U16707 (N_16707,N_12690,N_11994);
and U16708 (N_16708,N_11745,N_13343);
or U16709 (N_16709,N_10697,N_14331);
or U16710 (N_16710,N_12891,N_13692);
or U16711 (N_16711,N_13064,N_13892);
xnor U16712 (N_16712,N_11699,N_13241);
nand U16713 (N_16713,N_12367,N_10546);
xnor U16714 (N_16714,N_12351,N_11962);
nor U16715 (N_16715,N_11236,N_13776);
and U16716 (N_16716,N_12496,N_14097);
and U16717 (N_16717,N_14007,N_10445);
and U16718 (N_16718,N_14222,N_12828);
and U16719 (N_16719,N_10315,N_11340);
or U16720 (N_16720,N_13553,N_11663);
and U16721 (N_16721,N_14391,N_12545);
and U16722 (N_16722,N_13025,N_10708);
nand U16723 (N_16723,N_14207,N_13703);
xor U16724 (N_16724,N_10919,N_11716);
and U16725 (N_16725,N_12387,N_12701);
nor U16726 (N_16726,N_14086,N_14938);
xnor U16727 (N_16727,N_14177,N_14854);
nor U16728 (N_16728,N_13840,N_12720);
or U16729 (N_16729,N_13387,N_14001);
xor U16730 (N_16730,N_10349,N_10177);
xnor U16731 (N_16731,N_12409,N_13817);
nor U16732 (N_16732,N_11998,N_14029);
xnor U16733 (N_16733,N_11848,N_10797);
and U16734 (N_16734,N_14066,N_12554);
or U16735 (N_16735,N_12132,N_10334);
nand U16736 (N_16736,N_10071,N_12269);
or U16737 (N_16737,N_10963,N_11893);
and U16738 (N_16738,N_10078,N_11061);
nor U16739 (N_16739,N_14584,N_14577);
and U16740 (N_16740,N_13777,N_14194);
or U16741 (N_16741,N_14312,N_14551);
and U16742 (N_16742,N_12579,N_12437);
nand U16743 (N_16743,N_10755,N_11107);
and U16744 (N_16744,N_11756,N_11470);
or U16745 (N_16745,N_10756,N_11780);
nand U16746 (N_16746,N_14729,N_12651);
nor U16747 (N_16747,N_14631,N_12341);
nand U16748 (N_16748,N_12434,N_12689);
nand U16749 (N_16749,N_10733,N_10072);
and U16750 (N_16750,N_13920,N_12242);
and U16751 (N_16751,N_10355,N_10995);
nand U16752 (N_16752,N_13783,N_12790);
nor U16753 (N_16753,N_11847,N_10011);
and U16754 (N_16754,N_12171,N_13651);
nor U16755 (N_16755,N_13961,N_10254);
nor U16756 (N_16756,N_10974,N_10055);
or U16757 (N_16757,N_12820,N_14138);
nand U16758 (N_16758,N_12946,N_14256);
nand U16759 (N_16759,N_10176,N_11337);
nor U16760 (N_16760,N_11749,N_11907);
nor U16761 (N_16761,N_13641,N_13546);
nand U16762 (N_16762,N_10412,N_13970);
and U16763 (N_16763,N_10212,N_14251);
nand U16764 (N_16764,N_13633,N_12904);
and U16765 (N_16765,N_12766,N_13802);
xnor U16766 (N_16766,N_10451,N_11503);
nand U16767 (N_16767,N_13062,N_11545);
nor U16768 (N_16768,N_11595,N_12731);
or U16769 (N_16769,N_13835,N_12693);
and U16770 (N_16770,N_13131,N_11458);
or U16771 (N_16771,N_12525,N_10441);
nor U16772 (N_16772,N_13145,N_14909);
nand U16773 (N_16773,N_14384,N_12751);
nand U16774 (N_16774,N_12335,N_13512);
xor U16775 (N_16775,N_12411,N_13261);
and U16776 (N_16776,N_12940,N_13382);
and U16777 (N_16777,N_10942,N_13173);
or U16778 (N_16778,N_14157,N_12677);
xor U16779 (N_16779,N_13978,N_13326);
nor U16780 (N_16780,N_13928,N_12948);
xnor U16781 (N_16781,N_14957,N_13683);
nor U16782 (N_16782,N_13175,N_14567);
xnor U16783 (N_16783,N_13538,N_12812);
nand U16784 (N_16784,N_11818,N_11289);
and U16785 (N_16785,N_10716,N_12284);
or U16786 (N_16786,N_13417,N_10122);
nor U16787 (N_16787,N_14757,N_10364);
nand U16788 (N_16788,N_13975,N_13080);
nor U16789 (N_16789,N_12517,N_10618);
nor U16790 (N_16790,N_14417,N_13649);
nor U16791 (N_16791,N_13177,N_14421);
and U16792 (N_16792,N_10245,N_11760);
or U16793 (N_16793,N_14558,N_10752);
nand U16794 (N_16794,N_11086,N_14974);
nand U16795 (N_16795,N_10498,N_13968);
nand U16796 (N_16796,N_13972,N_13959);
nor U16797 (N_16797,N_14409,N_14901);
or U16798 (N_16798,N_14923,N_14560);
nand U16799 (N_16799,N_11945,N_13316);
and U16800 (N_16800,N_12543,N_14977);
and U16801 (N_16801,N_13504,N_12089);
and U16802 (N_16802,N_12312,N_10065);
and U16803 (N_16803,N_13092,N_12215);
and U16804 (N_16804,N_14300,N_11309);
nor U16805 (N_16805,N_14337,N_14479);
or U16806 (N_16806,N_12788,N_13566);
nand U16807 (N_16807,N_14534,N_14783);
or U16808 (N_16808,N_12309,N_13239);
and U16809 (N_16809,N_14433,N_10520);
or U16810 (N_16810,N_13503,N_10143);
and U16811 (N_16811,N_10000,N_14556);
nand U16812 (N_16812,N_13913,N_13296);
nand U16813 (N_16813,N_13290,N_13647);
nand U16814 (N_16814,N_12997,N_14041);
nand U16815 (N_16815,N_14394,N_10113);
nor U16816 (N_16816,N_13974,N_10091);
nand U16817 (N_16817,N_11323,N_11373);
and U16818 (N_16818,N_12144,N_12526);
nand U16819 (N_16819,N_12964,N_13684);
nor U16820 (N_16820,N_14753,N_11030);
nor U16821 (N_16821,N_14297,N_13044);
nor U16822 (N_16822,N_12944,N_14285);
or U16823 (N_16823,N_10598,N_10478);
nand U16824 (N_16824,N_11851,N_14161);
nand U16825 (N_16825,N_12957,N_10221);
nor U16826 (N_16826,N_12119,N_13853);
or U16827 (N_16827,N_10218,N_14682);
and U16828 (N_16828,N_12498,N_10163);
nor U16829 (N_16829,N_11533,N_13607);
nor U16830 (N_16830,N_11885,N_12017);
and U16831 (N_16831,N_14372,N_14676);
and U16832 (N_16832,N_14339,N_13618);
nand U16833 (N_16833,N_12048,N_10717);
and U16834 (N_16834,N_10952,N_11223);
or U16835 (N_16835,N_11417,N_14569);
and U16836 (N_16836,N_14301,N_14268);
and U16837 (N_16837,N_10787,N_13561);
or U16838 (N_16838,N_10621,N_10600);
or U16839 (N_16839,N_10632,N_12090);
nand U16840 (N_16840,N_10491,N_12053);
nor U16841 (N_16841,N_10100,N_13238);
or U16842 (N_16842,N_11963,N_13679);
xnor U16843 (N_16843,N_10021,N_12405);
and U16844 (N_16844,N_11310,N_11583);
nor U16845 (N_16845,N_10845,N_11120);
and U16846 (N_16846,N_14040,N_13578);
nand U16847 (N_16847,N_12208,N_12143);
and U16848 (N_16848,N_10112,N_11800);
xor U16849 (N_16849,N_14387,N_13415);
xnor U16850 (N_16850,N_10737,N_14486);
or U16851 (N_16851,N_11964,N_10150);
nand U16852 (N_16852,N_11333,N_11917);
nand U16853 (N_16853,N_12057,N_10358);
and U16854 (N_16854,N_13188,N_14530);
nor U16855 (N_16855,N_14107,N_12704);
nor U16856 (N_16856,N_14913,N_10596);
and U16857 (N_16857,N_14325,N_13662);
and U16858 (N_16858,N_11549,N_12976);
or U16859 (N_16859,N_12746,N_10404);
and U16860 (N_16860,N_10687,N_13144);
or U16861 (N_16861,N_13589,N_10577);
or U16862 (N_16862,N_11939,N_14248);
or U16863 (N_16863,N_14037,N_13820);
or U16864 (N_16864,N_13407,N_11959);
nor U16865 (N_16865,N_11977,N_10390);
nand U16866 (N_16866,N_10330,N_13381);
or U16867 (N_16867,N_12975,N_11697);
or U16868 (N_16868,N_11931,N_13358);
nor U16869 (N_16869,N_10539,N_14081);
nor U16870 (N_16870,N_12250,N_12362);
or U16871 (N_16871,N_12276,N_14918);
xor U16872 (N_16872,N_14649,N_13070);
nor U16873 (N_16873,N_11210,N_13369);
nor U16874 (N_16874,N_13323,N_10440);
nor U16875 (N_16875,N_12924,N_11858);
and U16876 (N_16876,N_10363,N_10237);
nand U16877 (N_16877,N_14382,N_11835);
and U16878 (N_16878,N_10130,N_12447);
nor U16879 (N_16879,N_10432,N_13263);
and U16880 (N_16880,N_14483,N_14528);
and U16881 (N_16881,N_14341,N_10168);
and U16882 (N_16882,N_14362,N_12596);
xnor U16883 (N_16883,N_10395,N_14659);
and U16884 (N_16884,N_10617,N_12922);
xor U16885 (N_16885,N_14553,N_14127);
nand U16886 (N_16886,N_11613,N_11041);
nor U16887 (N_16887,N_14615,N_13203);
xnor U16888 (N_16888,N_12176,N_11956);
nor U16889 (N_16889,N_10668,N_13026);
nand U16890 (N_16890,N_11617,N_12087);
nor U16891 (N_16891,N_13521,N_10465);
or U16892 (N_16892,N_11561,N_12665);
xnor U16893 (N_16893,N_14621,N_12568);
and U16894 (N_16894,N_14265,N_13855);
and U16895 (N_16895,N_10692,N_14190);
and U16896 (N_16896,N_14258,N_10075);
and U16897 (N_16897,N_14174,N_14917);
nor U16898 (N_16898,N_10833,N_13478);
nor U16899 (N_16899,N_12530,N_13781);
nand U16900 (N_16900,N_10366,N_10464);
xnor U16901 (N_16901,N_11219,N_13718);
and U16902 (N_16902,N_10647,N_11052);
or U16903 (N_16903,N_14116,N_10192);
and U16904 (N_16904,N_10146,N_13535);
nor U16905 (N_16905,N_11409,N_11543);
and U16906 (N_16906,N_12544,N_12070);
or U16907 (N_16907,N_14983,N_10350);
nor U16908 (N_16908,N_10509,N_11277);
nor U16909 (N_16909,N_13623,N_13125);
nor U16910 (N_16910,N_11584,N_13467);
xor U16911 (N_16911,N_10203,N_10519);
or U16912 (N_16912,N_14010,N_11296);
and U16913 (N_16913,N_11615,N_13540);
or U16914 (N_16914,N_13041,N_11128);
or U16915 (N_16915,N_12723,N_12581);
and U16916 (N_16916,N_12019,N_14358);
nand U16917 (N_16917,N_13965,N_11940);
nor U16918 (N_16918,N_13437,N_10422);
and U16919 (N_16919,N_12235,N_14489);
nand U16920 (N_16920,N_11211,N_12910);
nand U16921 (N_16921,N_13604,N_14632);
nand U16922 (N_16922,N_13846,N_10447);
nand U16923 (N_16923,N_14246,N_11987);
and U16924 (N_16924,N_10365,N_13657);
nand U16925 (N_16925,N_13280,N_10123);
or U16926 (N_16926,N_13664,N_11315);
nand U16927 (N_16927,N_12168,N_12908);
nand U16928 (N_16928,N_13401,N_10028);
or U16929 (N_16929,N_11623,N_12547);
xor U16930 (N_16930,N_13008,N_14985);
and U16931 (N_16931,N_13930,N_12458);
nor U16932 (N_16932,N_11166,N_13386);
or U16933 (N_16933,N_10102,N_13221);
and U16934 (N_16934,N_14781,N_12600);
nand U16935 (N_16935,N_12993,N_11937);
nor U16936 (N_16936,N_13340,N_12257);
or U16937 (N_16937,N_12773,N_11906);
xor U16938 (N_16938,N_10250,N_10586);
or U16939 (N_16939,N_14808,N_11072);
or U16940 (N_16940,N_11358,N_12674);
and U16941 (N_16941,N_11641,N_10991);
or U16942 (N_16942,N_11574,N_12522);
nand U16943 (N_16943,N_13422,N_14950);
and U16944 (N_16944,N_12851,N_13377);
nor U16945 (N_16945,N_13852,N_14317);
xnor U16946 (N_16946,N_10429,N_10976);
or U16947 (N_16947,N_12601,N_11488);
or U16948 (N_16948,N_14280,N_10981);
and U16949 (N_16949,N_10630,N_14061);
nand U16950 (N_16950,N_11798,N_12784);
nand U16951 (N_16951,N_12631,N_11805);
xnor U16952 (N_16952,N_14031,N_14311);
nand U16953 (N_16953,N_10508,N_13532);
nor U16954 (N_16954,N_11055,N_14100);
nor U16955 (N_16955,N_12234,N_10603);
or U16956 (N_16956,N_11298,N_13541);
and U16957 (N_16957,N_10735,N_11300);
or U16958 (N_16958,N_13191,N_12829);
and U16959 (N_16959,N_13611,N_13486);
nand U16960 (N_16960,N_14799,N_12305);
nand U16961 (N_16961,N_13357,N_13057);
xnor U16962 (N_16962,N_13163,N_10602);
and U16963 (N_16963,N_11596,N_12360);
nand U16964 (N_16964,N_11541,N_12378);
xnor U16965 (N_16965,N_12267,N_10239);
or U16966 (N_16966,N_12584,N_11573);
and U16967 (N_16967,N_11570,N_10808);
nor U16968 (N_16968,N_14723,N_12813);
and U16969 (N_16969,N_10870,N_13537);
or U16970 (N_16970,N_11552,N_12259);
and U16971 (N_16971,N_14398,N_13729);
and U16972 (N_16972,N_11970,N_14400);
xnor U16973 (N_16973,N_11982,N_11507);
or U16974 (N_16974,N_10706,N_10493);
xor U16975 (N_16975,N_11045,N_14053);
nand U16976 (N_16976,N_10195,N_10827);
nand U16977 (N_16977,N_14581,N_10304);
nor U16978 (N_16978,N_11306,N_13063);
nor U16979 (N_16979,N_12939,N_11829);
and U16980 (N_16980,N_10868,N_12787);
nor U16981 (N_16981,N_11270,N_10289);
nor U16982 (N_16982,N_10319,N_13450);
xor U16983 (N_16983,N_10229,N_10406);
or U16984 (N_16984,N_10514,N_11003);
or U16985 (N_16985,N_12966,N_11343);
and U16986 (N_16986,N_11376,N_11076);
and U16987 (N_16987,N_12273,N_11809);
nor U16988 (N_16988,N_12664,N_13942);
and U16989 (N_16989,N_13013,N_10675);
nand U16990 (N_16990,N_14535,N_10650);
and U16991 (N_16991,N_14079,N_13551);
nand U16992 (N_16992,N_14782,N_12389);
and U16993 (N_16993,N_11195,N_12901);
and U16994 (N_16994,N_10323,N_14962);
nand U16995 (N_16995,N_13520,N_13924);
or U16996 (N_16996,N_10326,N_12768);
xnor U16997 (N_16997,N_13941,N_13072);
and U16998 (N_16998,N_11282,N_13171);
nand U16999 (N_16999,N_10173,N_12187);
or U17000 (N_17000,N_14058,N_10505);
nor U17001 (N_17001,N_10589,N_11019);
and U17002 (N_17002,N_13134,N_11194);
nor U17003 (N_17003,N_12151,N_10443);
or U17004 (N_17004,N_13120,N_14758);
nor U17005 (N_17005,N_10230,N_10765);
nor U17006 (N_17006,N_12617,N_11395);
nand U17007 (N_17007,N_10206,N_10048);
nand U17008 (N_17008,N_10214,N_10608);
or U17009 (N_17009,N_12635,N_11092);
and U17010 (N_17010,N_13862,N_13429);
xor U17011 (N_17011,N_11984,N_10599);
and U17012 (N_17012,N_10485,N_10003);
nand U17013 (N_17013,N_10781,N_11811);
nor U17014 (N_17014,N_10805,N_14899);
nand U17015 (N_17015,N_10652,N_14393);
nor U17016 (N_17016,N_11554,N_12097);
or U17017 (N_17017,N_12465,N_10473);
xnor U17018 (N_17018,N_13746,N_14857);
xor U17019 (N_17019,N_11176,N_13453);
nor U17020 (N_17020,N_10303,N_12992);
nand U17021 (N_17021,N_11896,N_14257);
xor U17022 (N_17022,N_14326,N_11156);
nand U17023 (N_17023,N_14724,N_14237);
nand U17024 (N_17024,N_14146,N_10090);
nand U17025 (N_17025,N_11027,N_13668);
or U17026 (N_17026,N_10971,N_11565);
and U17027 (N_17027,N_14644,N_13742);
or U17028 (N_17028,N_12896,N_12741);
and U17029 (N_17029,N_14175,N_13714);
or U17030 (N_17030,N_10209,N_10453);
or U17031 (N_17031,N_10601,N_10132);
and U17032 (N_17032,N_13515,N_12212);
and U17033 (N_17033,N_10504,N_14225);
nor U17034 (N_17034,N_10339,N_14868);
and U17035 (N_17035,N_13513,N_14914);
nand U17036 (N_17036,N_10291,N_12621);
nor U17037 (N_17037,N_13935,N_11909);
nor U17038 (N_17038,N_13795,N_11692);
nand U17039 (N_17039,N_12846,N_14209);
nor U17040 (N_17040,N_11095,N_11777);
nor U17041 (N_17041,N_11648,N_11245);
nand U17042 (N_17042,N_12148,N_14030);
nand U17043 (N_17043,N_12594,N_10878);
or U17044 (N_17044,N_13253,N_12524);
or U17045 (N_17045,N_11892,N_12077);
nand U17046 (N_17046,N_12301,N_14978);
nand U17047 (N_17047,N_12637,N_11967);
and U17048 (N_17048,N_11161,N_11321);
nand U17049 (N_17049,N_11787,N_10530);
or U17050 (N_17050,N_13580,N_11801);
and U17051 (N_17051,N_13896,N_11913);
nand U17052 (N_17052,N_12634,N_13736);
nand U17053 (N_17053,N_12728,N_13897);
or U17054 (N_17054,N_10555,N_10431);
nand U17055 (N_17055,N_13088,N_13278);
and U17056 (N_17056,N_13678,N_12649);
xor U17057 (N_17057,N_14885,N_14859);
xor U17058 (N_17058,N_13129,N_12282);
or U17059 (N_17059,N_10407,N_10458);
nor U17060 (N_17060,N_12640,N_12230);
nand U17061 (N_17061,N_12657,N_11553);
or U17062 (N_17062,N_11485,N_13650);
nand U17063 (N_17063,N_10362,N_12348);
nand U17064 (N_17064,N_11795,N_14113);
nor U17065 (N_17065,N_10926,N_10767);
nor U17066 (N_17066,N_13596,N_10580);
nand U17067 (N_17067,N_13355,N_11733);
and U17068 (N_17068,N_14142,N_13798);
and U17069 (N_17069,N_13960,N_11248);
nand U17070 (N_17070,N_11048,N_14500);
or U17071 (N_17071,N_11135,N_13906);
and U17072 (N_17072,N_12091,N_13071);
nand U17073 (N_17073,N_11653,N_13130);
and U17074 (N_17074,N_12307,N_11021);
and U17075 (N_17075,N_13621,N_13059);
or U17076 (N_17076,N_12174,N_10332);
nand U17077 (N_17077,N_13043,N_13007);
or U17078 (N_17078,N_12268,N_13000);
nand U17079 (N_17079,N_13790,N_10370);
and U17080 (N_17080,N_10081,N_14006);
or U17081 (N_17081,N_14819,N_11579);
or U17082 (N_17082,N_12069,N_14439);
nand U17083 (N_17083,N_14716,N_14897);
nor U17084 (N_17084,N_10368,N_14595);
nand U17085 (N_17085,N_10541,N_11060);
or U17086 (N_17086,N_10518,N_14768);
xor U17087 (N_17087,N_14727,N_13441);
or U17088 (N_17088,N_14715,N_11423);
or U17089 (N_17089,N_14557,N_13841);
and U17090 (N_17090,N_12468,N_12133);
nor U17091 (N_17091,N_12386,N_11932);
xor U17092 (N_17092,N_12694,N_13851);
or U17093 (N_17093,N_10277,N_14315);
and U17094 (N_17094,N_14221,N_11542);
or U17095 (N_17095,N_10568,N_11546);
xnor U17096 (N_17096,N_10044,N_14693);
nor U17097 (N_17097,N_14117,N_14474);
nor U17098 (N_17098,N_13609,N_11766);
nor U17099 (N_17099,N_11392,N_11410);
nor U17100 (N_17100,N_10710,N_11621);
xor U17101 (N_17101,N_13723,N_11365);
nor U17102 (N_17102,N_14737,N_12916);
nand U17103 (N_17103,N_12560,N_13575);
and U17104 (N_17104,N_10750,N_12473);
and U17105 (N_17105,N_11259,N_11564);
or U17106 (N_17106,N_12612,N_12491);
nand U17107 (N_17107,N_14639,N_11789);
nor U17108 (N_17108,N_10947,N_13186);
or U17109 (N_17109,N_13517,N_10871);
or U17110 (N_17110,N_11118,N_13720);
nand U17111 (N_17111,N_12682,N_14004);
or U17112 (N_17112,N_10887,N_11432);
nand U17113 (N_17113,N_10196,N_12595);
nand U17114 (N_17114,N_13700,N_10171);
and U17115 (N_17115,N_14167,N_14354);
or U17116 (N_17116,N_14134,N_10766);
or U17117 (N_17117,N_13681,N_14216);
nor U17118 (N_17118,N_12921,N_10744);
and U17119 (N_17119,N_10740,N_14618);
and U17120 (N_17120,N_14603,N_13084);
nand U17121 (N_17121,N_11050,N_12294);
and U17122 (N_17122,N_11188,N_10246);
nor U17123 (N_17123,N_14407,N_12059);
and U17124 (N_17124,N_11106,N_11436);
nand U17125 (N_17125,N_14266,N_13005);
or U17126 (N_17126,N_13584,N_11066);
nor U17127 (N_17127,N_13903,N_12147);
nor U17128 (N_17128,N_11752,N_11183);
and U17129 (N_17129,N_12835,N_14456);
nand U17130 (N_17130,N_10482,N_12570);
xnor U17131 (N_17131,N_14893,N_13360);
nand U17132 (N_17132,N_11650,N_10391);
nand U17133 (N_17133,N_10397,N_13400);
and U17134 (N_17134,N_11303,N_13595);
or U17135 (N_17135,N_14140,N_12535);
nor U17136 (N_17136,N_10791,N_10516);
nor U17137 (N_17137,N_14763,N_10343);
and U17138 (N_17138,N_12549,N_11929);
or U17139 (N_17139,N_11004,N_12101);
xor U17140 (N_17140,N_10761,N_12749);
nor U17141 (N_17141,N_11062,N_10356);
xor U17142 (N_17142,N_10634,N_10795);
nor U17143 (N_17143,N_12729,N_13731);
and U17144 (N_17144,N_10881,N_10771);
or U17145 (N_17145,N_13151,N_14295);
or U17146 (N_17146,N_13711,N_14766);
xor U17147 (N_17147,N_11312,N_10084);
nand U17148 (N_17148,N_14844,N_14098);
nor U17149 (N_17149,N_14554,N_13734);
and U17150 (N_17150,N_14005,N_10341);
or U17151 (N_17151,N_10536,N_13074);
and U17152 (N_17152,N_13879,N_10975);
and U17153 (N_17153,N_14420,N_14032);
xnor U17154 (N_17154,N_12374,N_13991);
nand U17155 (N_17155,N_12585,N_12478);
nand U17156 (N_17156,N_11074,N_11942);
nor U17157 (N_17157,N_11718,N_10567);
nand U17158 (N_17158,N_13350,N_14740);
or U17159 (N_17159,N_13307,N_11187);
xor U17160 (N_17160,N_14444,N_12419);
nor U17161 (N_17161,N_11544,N_10178);
and U17162 (N_17162,N_11065,N_14710);
nor U17163 (N_17163,N_10425,N_11921);
or U17164 (N_17164,N_13162,N_14166);
and U17165 (N_17165,N_10477,N_10226);
or U17166 (N_17166,N_11018,N_10924);
nand U17167 (N_17167,N_14906,N_10627);
or U17168 (N_17168,N_13652,N_11534);
nand U17169 (N_17169,N_10475,N_14497);
and U17170 (N_17170,N_13167,N_13893);
nand U17171 (N_17171,N_10645,N_13153);
nand U17172 (N_17172,N_14623,N_12216);
or U17173 (N_17173,N_12688,N_14333);
nand U17174 (N_17174,N_14754,N_11029);
or U17175 (N_17175,N_14065,N_14840);
nor U17176 (N_17176,N_14865,N_11952);
nand U17177 (N_17177,N_13055,N_14706);
nand U17178 (N_17178,N_12238,N_12292);
xor U17179 (N_17179,N_12121,N_13599);
nor U17180 (N_17180,N_14249,N_11600);
and U17181 (N_17181,N_13073,N_14776);
nand U17182 (N_17182,N_14634,N_13479);
nor U17183 (N_17183,N_10640,N_11257);
and U17184 (N_17184,N_11131,N_14111);
nor U17185 (N_17185,N_12898,N_13670);
nand U17186 (N_17186,N_13446,N_10802);
nand U17187 (N_17187,N_12246,N_10824);
nand U17188 (N_17188,N_12841,N_11651);
and U17189 (N_17189,N_11894,N_14291);
or U17190 (N_17190,N_12537,N_13884);
nand U17191 (N_17191,N_12852,N_13150);
or U17192 (N_17192,N_14388,N_11421);
xor U17193 (N_17193,N_10175,N_13834);
nand U17194 (N_17194,N_10068,N_14022);
nor U17195 (N_17195,N_13413,N_10896);
xnor U17196 (N_17196,N_13653,N_12557);
nand U17197 (N_17197,N_10907,N_10385);
and U17198 (N_17198,N_12201,N_11491);
xor U17199 (N_17199,N_10029,N_13622);
xor U17200 (N_17200,N_13212,N_11823);
nor U17201 (N_17201,N_11955,N_12253);
nor U17202 (N_17202,N_11056,N_11997);
and U17203 (N_17203,N_10338,N_13912);
or U17204 (N_17204,N_11605,N_10352);
nand U17205 (N_17205,N_13523,N_14905);
and U17206 (N_17206,N_11244,N_10117);
xor U17207 (N_17207,N_12384,N_12735);
nand U17208 (N_17208,N_10419,N_12128);
or U17209 (N_17209,N_12481,N_10264);
nor U17210 (N_17210,N_12303,N_11705);
nand U17211 (N_17211,N_10857,N_14233);
nor U17212 (N_17212,N_11958,N_10141);
xor U17213 (N_17213,N_11268,N_13508);
nor U17214 (N_17214,N_14690,N_10661);
or U17215 (N_17215,N_12981,N_13615);
nor U17216 (N_17216,N_12756,N_12955);
nand U17217 (N_17217,N_14640,N_14196);
or U17218 (N_17218,N_13294,N_13396);
or U17219 (N_17219,N_14968,N_11130);
nand U17220 (N_17220,N_11457,N_13953);
or U17221 (N_17221,N_14779,N_13270);
nand U17222 (N_17222,N_10056,N_13374);
nor U17223 (N_17223,N_10804,N_13126);
nand U17224 (N_17224,N_14122,N_13764);
xnor U17225 (N_17225,N_10691,N_11569);
xor U17226 (N_17226,N_10063,N_12254);
xor U17227 (N_17227,N_13371,N_12532);
nor U17228 (N_17228,N_12932,N_10251);
nand U17229 (N_17229,N_11201,N_12848);
and U17230 (N_17230,N_12899,N_14158);
nor U17231 (N_17231,N_12283,N_11571);
nand U17232 (N_17232,N_13285,N_10738);
nand U17233 (N_17233,N_12279,N_11427);
or U17234 (N_17234,N_13193,N_14795);
or U17235 (N_17235,N_10392,N_12642);
nor U17236 (N_17236,N_11817,N_14816);
nor U17237 (N_17237,N_14461,N_12010);
and U17238 (N_17238,N_11116,N_10376);
nor U17239 (N_17239,N_11078,N_13755);
and U17240 (N_17240,N_14091,N_12868);
and U17241 (N_17241,N_10763,N_13645);
or U17242 (N_17242,N_12197,N_10179);
nand U17243 (N_17243,N_12206,N_12298);
nor U17244 (N_17244,N_11636,N_11280);
nor U17245 (N_17245,N_12304,N_11179);
or U17246 (N_17246,N_10969,N_14171);
or U17247 (N_17247,N_10658,N_14540);
nor U17248 (N_17248,N_10642,N_13227);
nor U17249 (N_17249,N_14817,N_13458);
nand U17250 (N_17250,N_11234,N_12402);
nand U17251 (N_17251,N_13028,N_12175);
or U17252 (N_17252,N_11771,N_10549);
nor U17253 (N_17253,N_11331,N_13709);
nand U17254 (N_17254,N_11884,N_13205);
nor U17255 (N_17255,N_12459,N_11751);
nor U17256 (N_17256,N_12076,N_13324);
and U17257 (N_17257,N_11077,N_11778);
or U17258 (N_17258,N_14714,N_13406);
nor U17259 (N_17259,N_14283,N_13635);
or U17260 (N_17260,N_12210,N_11424);
and U17261 (N_17261,N_10793,N_12745);
and U17262 (N_17262,N_12562,N_10954);
or U17263 (N_17263,N_13890,N_10375);
nand U17264 (N_17264,N_10116,N_11768);
and U17265 (N_17265,N_14144,N_14646);
nand U17266 (N_17266,N_11444,N_12377);
nand U17267 (N_17267,N_12178,N_14455);
nor U17268 (N_17268,N_12534,N_11073);
nor U17269 (N_17269,N_13489,N_14443);
or U17270 (N_17270,N_12656,N_13909);
nor U17271 (N_17271,N_10990,N_11904);
or U17272 (N_17272,N_13031,N_14541);
and U17273 (N_17273,N_11674,N_10281);
nor U17274 (N_17274,N_10416,N_11155);
nand U17275 (N_17275,N_11704,N_12730);
and U17276 (N_17276,N_13588,N_14408);
nand U17277 (N_17277,N_12198,N_11261);
or U17278 (N_17278,N_13998,N_10743);
or U17279 (N_17279,N_10309,N_14627);
or U17280 (N_17280,N_10335,N_10007);
and U17281 (N_17281,N_10216,N_12949);
and U17282 (N_17282,N_14262,N_14837);
or U17283 (N_17283,N_13563,N_10502);
or U17284 (N_17284,N_13809,N_13944);
and U17285 (N_17285,N_12959,N_10472);
nand U17286 (N_17286,N_14681,N_14922);
and U17287 (N_17287,N_10876,N_13613);
nand U17288 (N_17288,N_12388,N_12794);
and U17289 (N_17289,N_12673,N_14080);
nor U17290 (N_17290,N_14531,N_12150);
or U17291 (N_17291,N_11902,N_14670);
or U17292 (N_17292,N_10837,N_11548);
nand U17293 (N_17293,N_12540,N_12819);
and U17294 (N_17294,N_11221,N_14664);
nor U17295 (N_17295,N_13119,N_11599);
or U17296 (N_17296,N_13778,N_13200);
and U17297 (N_17297,N_11157,N_12571);
or U17298 (N_17298,N_13006,N_11676);
nor U17299 (N_17299,N_12793,N_14464);
nand U17300 (N_17300,N_10097,N_10523);
nor U17301 (N_17301,N_10299,N_11802);
and U17302 (N_17302,N_12449,N_11490);
nor U17303 (N_17303,N_10353,N_12893);
nand U17304 (N_17304,N_11492,N_10377);
or U17305 (N_17305,N_11067,N_11112);
nand U17306 (N_17306,N_12973,N_14996);
xnor U17307 (N_17307,N_11291,N_13811);
and U17308 (N_17308,N_14432,N_14105);
and U17309 (N_17309,N_12054,N_10764);
nand U17310 (N_17310,N_10860,N_11672);
or U17311 (N_17311,N_11640,N_14219);
nor U17312 (N_17312,N_12774,N_12152);
xor U17313 (N_17313,N_14731,N_13154);
or U17314 (N_17314,N_11598,N_11267);
nand U17315 (N_17315,N_10034,N_14524);
and U17316 (N_17316,N_10759,N_11232);
nor U17317 (N_17317,N_12606,N_11064);
nor U17318 (N_17318,N_11837,N_10820);
nor U17319 (N_17319,N_12486,N_14184);
nand U17320 (N_17320,N_13948,N_11496);
and U17321 (N_17321,N_14045,N_14051);
and U17322 (N_17322,N_11563,N_13100);
nand U17323 (N_17323,N_11347,N_10674);
nor U17324 (N_17324,N_11168,N_12408);
nor U17325 (N_17325,N_10915,N_13332);
or U17326 (N_17326,N_12566,N_12984);
or U17327 (N_17327,N_11515,N_11880);
nand U17328 (N_17328,N_13501,N_11182);
nor U17329 (N_17329,N_14472,N_14933);
nor U17330 (N_17330,N_12456,N_12433);
xnor U17331 (N_17331,N_11625,N_10806);
nand U17332 (N_17332,N_10742,N_12310);
nand U17333 (N_17333,N_14851,N_14287);
and U17334 (N_17334,N_11054,N_14230);
and U17335 (N_17335,N_13500,N_13940);
or U17336 (N_17336,N_14182,N_12880);
nor U17337 (N_17337,N_14159,N_13012);
nand U17338 (N_17338,N_10351,N_11715);
nor U17339 (N_17339,N_12950,N_13362);
nand U17340 (N_17340,N_10083,N_10374);
nand U17341 (N_17341,N_13787,N_12605);
and U17342 (N_17342,N_11009,N_11501);
nand U17343 (N_17343,N_13209,N_12798);
nand U17344 (N_17344,N_12118,N_10018);
xor U17345 (N_17345,N_13321,N_13582);
nor U17346 (N_17346,N_14679,N_11518);
xnor U17347 (N_17347,N_14403,N_13506);
or U17348 (N_17348,N_10670,N_11011);
and U17349 (N_17349,N_12862,N_13902);
and U17350 (N_17350,N_13123,N_12867);
or U17351 (N_17351,N_14114,N_13666);
and U17352 (N_17352,N_11973,N_10572);
nor U17353 (N_17353,N_12860,N_12154);
nand U17354 (N_17354,N_11089,N_11827);
or U17355 (N_17355,N_12783,N_12968);
nor U17356 (N_17356,N_12630,N_10489);
nand U17357 (N_17357,N_10828,N_11037);
and U17358 (N_17358,N_13883,N_13685);
nand U17359 (N_17359,N_11920,N_11014);
nand U17360 (N_17360,N_14277,N_13452);
nand U17361 (N_17361,N_12620,N_10278);
or U17362 (N_17362,N_14571,N_11930);
nor U17363 (N_17363,N_14206,N_10904);
or U17364 (N_17364,N_11144,N_13558);
and U17365 (N_17365,N_11017,N_14110);
nand U17366 (N_17366,N_13359,N_10506);
nand U17367 (N_17367,N_11216,N_11005);
and U17368 (N_17368,N_11665,N_12270);
xnor U17369 (N_17369,N_11446,N_12780);
nor U17370 (N_17370,N_13196,N_14637);
nand U17371 (N_17371,N_10066,N_10135);
nand U17372 (N_17372,N_13542,N_10943);
nand U17373 (N_17373,N_14314,N_14624);
nand U17374 (N_17374,N_11302,N_12355);
nand U17375 (N_17375,N_10623,N_12011);
or U17376 (N_17376,N_10444,N_14254);
or U17377 (N_17377,N_10131,N_11513);
or U17378 (N_17378,N_13160,N_12806);
or U17379 (N_17379,N_13425,N_11249);
and U17380 (N_17380,N_12935,N_13397);
and U17381 (N_17381,N_14604,N_11933);
xnor U17382 (N_17382,N_13529,N_14244);
and U17383 (N_17383,N_10984,N_13983);
nand U17384 (N_17384,N_13233,N_14255);
or U17385 (N_17385,N_11783,N_10923);
xor U17386 (N_17386,N_11006,N_13081);
xnor U17387 (N_17387,N_10611,N_11925);
nor U17388 (N_17388,N_12598,N_12291);
nand U17389 (N_17389,N_12359,N_10333);
xor U17390 (N_17390,N_11572,N_12941);
nand U17391 (N_17391,N_11986,N_14028);
nand U17392 (N_17392,N_13639,N_10666);
nand U17393 (N_17393,N_11709,N_12214);
or U17394 (N_17394,N_14057,N_14469);
xor U17395 (N_17395,N_11047,N_11606);
and U17396 (N_17396,N_11633,N_10614);
or U17397 (N_17397,N_11136,N_14386);
or U17398 (N_17398,N_10880,N_12211);
xor U17399 (N_17399,N_10654,N_11363);
or U17400 (N_17400,N_14172,N_13565);
or U17401 (N_17401,N_14468,N_13181);
xnor U17402 (N_17402,N_10711,N_13496);
nand U17403 (N_17403,N_12681,N_14026);
nand U17404 (N_17404,N_10812,N_13581);
or U17405 (N_17405,N_13550,N_14082);
and U17406 (N_17406,N_12141,N_10511);
nand U17407 (N_17407,N_10571,N_11936);
nand U17408 (N_17408,N_13699,N_12615);
and U17409 (N_17409,N_13142,N_11445);
or U17410 (N_17410,N_14997,N_12951);
or U17411 (N_17411,N_10957,N_14231);
and U17412 (N_17412,N_14858,N_10929);
nor U17413 (N_17413,N_10859,N_14835);
and U17414 (N_17414,N_14863,N_13547);
and U17415 (N_17415,N_12697,N_14052);
nor U17416 (N_17416,N_13844,N_12663);
nand U17417 (N_17417,N_14705,N_11498);
xor U17418 (N_17418,N_11233,N_11198);
or U17419 (N_17419,N_13638,N_13376);
and U17420 (N_17420,N_11246,N_11968);
nor U17421 (N_17421,N_10016,N_11635);
or U17422 (N_17422,N_11419,N_11524);
or U17423 (N_17423,N_12379,N_13534);
and U17424 (N_17424,N_11647,N_14942);
nor U17425 (N_17425,N_12513,N_11452);
or U17426 (N_17426,N_13619,N_10699);
xor U17427 (N_17427,N_14276,N_14308);
xor U17428 (N_17428,N_13889,N_10215);
or U17429 (N_17429,N_12864,N_10064);
nand U17430 (N_17430,N_14457,N_12224);
or U17431 (N_17431,N_13218,N_11487);
and U17432 (N_17432,N_10047,N_13480);
and U17433 (N_17433,N_11926,N_13654);
nor U17434 (N_17434,N_13330,N_11993);
xnor U17435 (N_17435,N_14638,N_14686);
nor U17436 (N_17436,N_14719,N_11785);
and U17437 (N_17437,N_10243,N_10663);
nand U17438 (N_17438,N_13603,N_14470);
nor U17439 (N_17439,N_14377,N_14220);
xnor U17440 (N_17440,N_10040,N_10147);
nor U17441 (N_17441,N_10104,N_11057);
nor U17442 (N_17442,N_11231,N_13738);
xor U17443 (N_17443,N_14252,N_14017);
or U17444 (N_17444,N_13644,N_11714);
or U17445 (N_17445,N_10082,N_10783);
nand U17446 (N_17446,N_14888,N_12853);
nand U17447 (N_17447,N_10593,N_10079);
nand U17448 (N_17448,N_12942,N_13593);
nor U17449 (N_17449,N_14371,N_14147);
and U17450 (N_17450,N_10713,N_10322);
and U17451 (N_17451,N_14327,N_12859);
nand U17452 (N_17452,N_10378,N_10753);
or U17453 (N_17453,N_13804,N_12217);
and U17454 (N_17454,N_14861,N_12710);
nor U17455 (N_17455,N_11610,N_14881);
and U17456 (N_17456,N_12111,N_13306);
nand U17457 (N_17457,N_10269,N_14168);
or U17458 (N_17458,N_13404,N_11857);
nor U17459 (N_17459,N_12122,N_12041);
xor U17460 (N_17460,N_10155,N_11690);
nand U17461 (N_17461,N_11164,N_10145);
xnor U17462 (N_17462,N_14889,N_10722);
and U17463 (N_17463,N_14884,N_14510);
or U17464 (N_17464,N_13908,N_11763);
or U17465 (N_17465,N_13085,N_11129);
and U17466 (N_17466,N_13525,N_13926);
nor U17467 (N_17467,N_13980,N_10070);
and U17468 (N_17468,N_10936,N_13614);
nor U17469 (N_17469,N_14662,N_10893);
xnor U17470 (N_17470,N_13430,N_14485);
nor U17471 (N_17471,N_12104,N_14658);
nand U17472 (N_17472,N_12671,N_12715);
nand U17473 (N_17473,N_13117,N_12703);
and U17474 (N_17474,N_13379,N_11000);
nor U17475 (N_17475,N_10702,N_11117);
nor U17476 (N_17476,N_12190,N_14912);
nor U17477 (N_17477,N_14290,N_12414);
and U17478 (N_17478,N_11222,N_12610);
nor U17479 (N_17479,N_11469,N_12527);
and U17480 (N_17480,N_13473,N_11996);
nand U17481 (N_17481,N_13832,N_13569);
nor U17482 (N_17482,N_12479,N_14139);
or U17483 (N_17483,N_10949,N_10317);
nand U17484 (N_17484,N_10270,N_14183);
or U17485 (N_17485,N_14787,N_11262);
nand U17486 (N_17486,N_11437,N_14092);
and U17487 (N_17487,N_10754,N_11511);
and U17488 (N_17488,N_14636,N_12505);
or U17489 (N_17489,N_14025,N_14563);
and U17490 (N_17490,N_11370,N_12394);
nand U17491 (N_17491,N_10455,N_11844);
nor U17492 (N_17492,N_14292,N_13165);
or U17493 (N_17493,N_14936,N_12827);
and U17494 (N_17494,N_14396,N_14990);
nor U17495 (N_17495,N_14274,N_12322);
nand U17496 (N_17496,N_13583,N_14961);
nand U17497 (N_17497,N_13042,N_13659);
and U17498 (N_17498,N_11430,N_13626);
or U17499 (N_17499,N_12251,N_14155);
or U17500 (N_17500,N_11783,N_10478);
nor U17501 (N_17501,N_11034,N_12838);
xnor U17502 (N_17502,N_11535,N_13649);
nand U17503 (N_17503,N_14235,N_12117);
nor U17504 (N_17504,N_10737,N_12597);
xnor U17505 (N_17505,N_11257,N_14962);
xor U17506 (N_17506,N_10126,N_14872);
and U17507 (N_17507,N_12751,N_10844);
xor U17508 (N_17508,N_10150,N_11365);
and U17509 (N_17509,N_10651,N_11552);
xor U17510 (N_17510,N_11146,N_14133);
or U17511 (N_17511,N_12142,N_14871);
nand U17512 (N_17512,N_14607,N_13812);
nor U17513 (N_17513,N_12788,N_13718);
nor U17514 (N_17514,N_12049,N_14697);
xor U17515 (N_17515,N_12932,N_13253);
and U17516 (N_17516,N_11614,N_14394);
nand U17517 (N_17517,N_13106,N_14558);
and U17518 (N_17518,N_12846,N_14563);
nor U17519 (N_17519,N_13888,N_14902);
nor U17520 (N_17520,N_13180,N_10665);
or U17521 (N_17521,N_10648,N_11968);
and U17522 (N_17522,N_10074,N_13995);
nand U17523 (N_17523,N_13177,N_12542);
nor U17524 (N_17524,N_11650,N_12011);
and U17525 (N_17525,N_10736,N_10921);
nand U17526 (N_17526,N_14195,N_14618);
nor U17527 (N_17527,N_13650,N_10439);
nand U17528 (N_17528,N_11617,N_13281);
and U17529 (N_17529,N_10610,N_14033);
nor U17530 (N_17530,N_14558,N_13906);
and U17531 (N_17531,N_13476,N_12352);
nor U17532 (N_17532,N_12248,N_14523);
and U17533 (N_17533,N_14046,N_14064);
nand U17534 (N_17534,N_10379,N_14955);
or U17535 (N_17535,N_10611,N_11747);
and U17536 (N_17536,N_12263,N_13970);
nor U17537 (N_17537,N_13536,N_12718);
nor U17538 (N_17538,N_13651,N_13387);
nand U17539 (N_17539,N_10463,N_11741);
or U17540 (N_17540,N_14824,N_14039);
xor U17541 (N_17541,N_11311,N_12493);
or U17542 (N_17542,N_10505,N_14091);
xor U17543 (N_17543,N_11931,N_10989);
and U17544 (N_17544,N_10040,N_13713);
and U17545 (N_17545,N_10493,N_12237);
nor U17546 (N_17546,N_13924,N_13786);
xor U17547 (N_17547,N_14078,N_14498);
or U17548 (N_17548,N_11171,N_12291);
nand U17549 (N_17549,N_12805,N_10390);
xnor U17550 (N_17550,N_14926,N_13162);
or U17551 (N_17551,N_10385,N_10679);
xnor U17552 (N_17552,N_10357,N_12997);
xnor U17553 (N_17553,N_10938,N_14602);
and U17554 (N_17554,N_13573,N_13992);
nand U17555 (N_17555,N_13963,N_10251);
nor U17556 (N_17556,N_12473,N_12177);
and U17557 (N_17557,N_11423,N_11355);
nand U17558 (N_17558,N_10124,N_12255);
nand U17559 (N_17559,N_14946,N_13599);
nand U17560 (N_17560,N_14378,N_10858);
nor U17561 (N_17561,N_12310,N_14060);
and U17562 (N_17562,N_14375,N_10847);
nor U17563 (N_17563,N_14050,N_13544);
nor U17564 (N_17564,N_13912,N_10472);
or U17565 (N_17565,N_12161,N_14121);
xnor U17566 (N_17566,N_14295,N_12397);
nand U17567 (N_17567,N_11148,N_12540);
and U17568 (N_17568,N_11118,N_11348);
nor U17569 (N_17569,N_14885,N_11977);
xor U17570 (N_17570,N_12239,N_12791);
and U17571 (N_17571,N_12274,N_10204);
and U17572 (N_17572,N_13131,N_14289);
nor U17573 (N_17573,N_11843,N_12597);
or U17574 (N_17574,N_12676,N_13810);
or U17575 (N_17575,N_11512,N_10022);
and U17576 (N_17576,N_14959,N_13209);
nor U17577 (N_17577,N_12741,N_10003);
nand U17578 (N_17578,N_12519,N_14133);
nor U17579 (N_17579,N_14651,N_12909);
nand U17580 (N_17580,N_12448,N_14747);
nor U17581 (N_17581,N_14187,N_14339);
nand U17582 (N_17582,N_11422,N_11462);
or U17583 (N_17583,N_13482,N_11708);
nand U17584 (N_17584,N_14317,N_12479);
and U17585 (N_17585,N_10816,N_12603);
nand U17586 (N_17586,N_14963,N_13206);
nand U17587 (N_17587,N_14921,N_10747);
nor U17588 (N_17588,N_10769,N_12170);
nor U17589 (N_17589,N_14650,N_13283);
nor U17590 (N_17590,N_10437,N_11256);
and U17591 (N_17591,N_10949,N_14037);
nand U17592 (N_17592,N_11505,N_12566);
nand U17593 (N_17593,N_10056,N_12584);
nand U17594 (N_17594,N_14137,N_12946);
and U17595 (N_17595,N_13120,N_14942);
or U17596 (N_17596,N_10361,N_14959);
xor U17597 (N_17597,N_13293,N_14104);
nor U17598 (N_17598,N_11691,N_14203);
nor U17599 (N_17599,N_14677,N_12207);
nand U17600 (N_17600,N_14427,N_14750);
or U17601 (N_17601,N_12447,N_13640);
xnor U17602 (N_17602,N_14362,N_11580);
or U17603 (N_17603,N_11823,N_11545);
and U17604 (N_17604,N_14634,N_12419);
xnor U17605 (N_17605,N_11171,N_10660);
nor U17606 (N_17606,N_14047,N_14220);
or U17607 (N_17607,N_14911,N_13205);
nor U17608 (N_17608,N_13868,N_10004);
or U17609 (N_17609,N_10118,N_11489);
nor U17610 (N_17610,N_10554,N_13387);
nor U17611 (N_17611,N_14150,N_12578);
or U17612 (N_17612,N_14955,N_12333);
nor U17613 (N_17613,N_10325,N_11438);
nand U17614 (N_17614,N_11463,N_14698);
and U17615 (N_17615,N_11836,N_13360);
or U17616 (N_17616,N_14692,N_14361);
or U17617 (N_17617,N_11081,N_13978);
nor U17618 (N_17618,N_14070,N_11525);
and U17619 (N_17619,N_11557,N_13086);
nand U17620 (N_17620,N_13903,N_12382);
nand U17621 (N_17621,N_12952,N_14990);
nand U17622 (N_17622,N_13500,N_14913);
or U17623 (N_17623,N_14517,N_10904);
and U17624 (N_17624,N_10635,N_13698);
xor U17625 (N_17625,N_11121,N_14488);
nand U17626 (N_17626,N_11696,N_13286);
and U17627 (N_17627,N_10493,N_10374);
and U17628 (N_17628,N_10204,N_10642);
and U17629 (N_17629,N_11656,N_13979);
nor U17630 (N_17630,N_14505,N_12100);
nor U17631 (N_17631,N_12159,N_14709);
xor U17632 (N_17632,N_11224,N_14601);
and U17633 (N_17633,N_11173,N_11396);
or U17634 (N_17634,N_14862,N_14957);
xnor U17635 (N_17635,N_10275,N_12465);
nor U17636 (N_17636,N_10482,N_11654);
and U17637 (N_17637,N_14660,N_10749);
nand U17638 (N_17638,N_10401,N_13047);
nand U17639 (N_17639,N_14636,N_13085);
nand U17640 (N_17640,N_10044,N_11432);
or U17641 (N_17641,N_13679,N_12486);
nand U17642 (N_17642,N_10045,N_12260);
or U17643 (N_17643,N_13173,N_10451);
and U17644 (N_17644,N_14471,N_10983);
nor U17645 (N_17645,N_10951,N_13573);
and U17646 (N_17646,N_10357,N_10374);
nor U17647 (N_17647,N_12483,N_11405);
or U17648 (N_17648,N_11976,N_12218);
nand U17649 (N_17649,N_13328,N_12776);
nand U17650 (N_17650,N_10299,N_13574);
xnor U17651 (N_17651,N_11635,N_10617);
nand U17652 (N_17652,N_10417,N_14148);
nand U17653 (N_17653,N_13511,N_11750);
xor U17654 (N_17654,N_11386,N_10495);
or U17655 (N_17655,N_14109,N_14846);
xnor U17656 (N_17656,N_11072,N_14210);
nand U17657 (N_17657,N_12370,N_12693);
and U17658 (N_17658,N_11138,N_11872);
and U17659 (N_17659,N_14994,N_12391);
nand U17660 (N_17660,N_14371,N_10641);
nand U17661 (N_17661,N_11549,N_13027);
nand U17662 (N_17662,N_12926,N_13844);
nand U17663 (N_17663,N_11524,N_13550);
and U17664 (N_17664,N_10060,N_13222);
or U17665 (N_17665,N_14097,N_12308);
and U17666 (N_17666,N_11663,N_14944);
xor U17667 (N_17667,N_14561,N_14515);
nand U17668 (N_17668,N_13617,N_10447);
nand U17669 (N_17669,N_13420,N_10475);
or U17670 (N_17670,N_12735,N_13256);
nand U17671 (N_17671,N_10661,N_13579);
nor U17672 (N_17672,N_10413,N_13052);
xnor U17673 (N_17673,N_10724,N_11574);
xnor U17674 (N_17674,N_14274,N_14511);
nand U17675 (N_17675,N_11712,N_10682);
nor U17676 (N_17676,N_10771,N_14509);
or U17677 (N_17677,N_14276,N_10612);
and U17678 (N_17678,N_12717,N_14676);
and U17679 (N_17679,N_12737,N_10793);
or U17680 (N_17680,N_12012,N_14594);
nand U17681 (N_17681,N_10702,N_12752);
nand U17682 (N_17682,N_10650,N_14883);
or U17683 (N_17683,N_11886,N_10257);
nor U17684 (N_17684,N_11354,N_14925);
nor U17685 (N_17685,N_11353,N_13260);
nor U17686 (N_17686,N_14000,N_14547);
nand U17687 (N_17687,N_11915,N_10382);
nor U17688 (N_17688,N_13181,N_13772);
nor U17689 (N_17689,N_11591,N_14607);
or U17690 (N_17690,N_14618,N_12555);
and U17691 (N_17691,N_12145,N_14582);
or U17692 (N_17692,N_13406,N_14254);
and U17693 (N_17693,N_13369,N_13642);
nand U17694 (N_17694,N_12914,N_14573);
and U17695 (N_17695,N_11763,N_11853);
and U17696 (N_17696,N_13342,N_13145);
or U17697 (N_17697,N_13490,N_13815);
nor U17698 (N_17698,N_13006,N_10608);
nor U17699 (N_17699,N_12506,N_14883);
nor U17700 (N_17700,N_11346,N_11590);
nand U17701 (N_17701,N_10626,N_13511);
nand U17702 (N_17702,N_12011,N_10075);
nand U17703 (N_17703,N_12572,N_12864);
nor U17704 (N_17704,N_14935,N_12161);
and U17705 (N_17705,N_14892,N_12293);
or U17706 (N_17706,N_14684,N_10727);
nand U17707 (N_17707,N_10558,N_11741);
and U17708 (N_17708,N_10248,N_12137);
nand U17709 (N_17709,N_14992,N_14188);
nor U17710 (N_17710,N_10365,N_12398);
or U17711 (N_17711,N_12088,N_11445);
nor U17712 (N_17712,N_14880,N_10836);
nor U17713 (N_17713,N_13417,N_12930);
nand U17714 (N_17714,N_11037,N_11420);
nand U17715 (N_17715,N_13183,N_11583);
or U17716 (N_17716,N_14397,N_12341);
nand U17717 (N_17717,N_13942,N_12341);
nand U17718 (N_17718,N_14477,N_13756);
xor U17719 (N_17719,N_12186,N_10013);
nand U17720 (N_17720,N_10376,N_12652);
nand U17721 (N_17721,N_14833,N_11037);
nand U17722 (N_17722,N_14741,N_14259);
and U17723 (N_17723,N_11961,N_10549);
nor U17724 (N_17724,N_14454,N_12134);
nand U17725 (N_17725,N_10117,N_13351);
nand U17726 (N_17726,N_12356,N_13249);
and U17727 (N_17727,N_13867,N_11103);
or U17728 (N_17728,N_12808,N_10766);
nor U17729 (N_17729,N_14983,N_13512);
nor U17730 (N_17730,N_12690,N_13725);
nand U17731 (N_17731,N_12988,N_12876);
nand U17732 (N_17732,N_10016,N_13955);
and U17733 (N_17733,N_11387,N_14904);
nor U17734 (N_17734,N_10863,N_10154);
xnor U17735 (N_17735,N_11606,N_10883);
xor U17736 (N_17736,N_12245,N_10623);
nor U17737 (N_17737,N_12921,N_14062);
nor U17738 (N_17738,N_13598,N_11257);
or U17739 (N_17739,N_11452,N_13161);
xor U17740 (N_17740,N_13376,N_10890);
nor U17741 (N_17741,N_11686,N_12992);
nand U17742 (N_17742,N_12735,N_12517);
nand U17743 (N_17743,N_14555,N_10103);
nor U17744 (N_17744,N_14668,N_11646);
nand U17745 (N_17745,N_13182,N_10410);
and U17746 (N_17746,N_13461,N_11059);
nor U17747 (N_17747,N_14014,N_14702);
and U17748 (N_17748,N_14858,N_10351);
or U17749 (N_17749,N_14369,N_11959);
nand U17750 (N_17750,N_12241,N_14573);
and U17751 (N_17751,N_10562,N_13044);
nand U17752 (N_17752,N_14276,N_13477);
and U17753 (N_17753,N_13004,N_14187);
nand U17754 (N_17754,N_10847,N_11329);
nor U17755 (N_17755,N_13620,N_12657);
or U17756 (N_17756,N_10843,N_14845);
nor U17757 (N_17757,N_13967,N_13108);
and U17758 (N_17758,N_11344,N_13682);
or U17759 (N_17759,N_14514,N_12260);
nand U17760 (N_17760,N_14825,N_14878);
nand U17761 (N_17761,N_12202,N_12230);
nor U17762 (N_17762,N_10727,N_11611);
nor U17763 (N_17763,N_13746,N_13352);
and U17764 (N_17764,N_10068,N_14638);
nand U17765 (N_17765,N_14753,N_10346);
nand U17766 (N_17766,N_11991,N_10033);
and U17767 (N_17767,N_11594,N_13397);
nand U17768 (N_17768,N_11854,N_10471);
nand U17769 (N_17769,N_14433,N_12184);
nor U17770 (N_17770,N_12004,N_11599);
nor U17771 (N_17771,N_11526,N_12412);
xor U17772 (N_17772,N_11244,N_14504);
and U17773 (N_17773,N_14665,N_10977);
nor U17774 (N_17774,N_10325,N_14275);
and U17775 (N_17775,N_11797,N_13825);
or U17776 (N_17776,N_14305,N_14721);
xor U17777 (N_17777,N_12644,N_12122);
nand U17778 (N_17778,N_13623,N_12688);
xor U17779 (N_17779,N_12468,N_13874);
and U17780 (N_17780,N_11088,N_13826);
or U17781 (N_17781,N_10040,N_14485);
or U17782 (N_17782,N_11249,N_11400);
nor U17783 (N_17783,N_10439,N_10213);
and U17784 (N_17784,N_10369,N_14821);
or U17785 (N_17785,N_11701,N_14622);
and U17786 (N_17786,N_11498,N_10628);
nand U17787 (N_17787,N_13958,N_11471);
and U17788 (N_17788,N_14700,N_11623);
nor U17789 (N_17789,N_11195,N_13052);
nand U17790 (N_17790,N_11475,N_11449);
xor U17791 (N_17791,N_10117,N_12903);
nor U17792 (N_17792,N_12929,N_11512);
or U17793 (N_17793,N_10183,N_14541);
nor U17794 (N_17794,N_14955,N_12066);
and U17795 (N_17795,N_11459,N_13456);
nand U17796 (N_17796,N_13538,N_12142);
nand U17797 (N_17797,N_11406,N_11876);
xor U17798 (N_17798,N_14670,N_12947);
nand U17799 (N_17799,N_10801,N_11747);
nand U17800 (N_17800,N_14834,N_11603);
and U17801 (N_17801,N_14078,N_12046);
nor U17802 (N_17802,N_13359,N_14056);
or U17803 (N_17803,N_10244,N_12578);
xnor U17804 (N_17804,N_14971,N_13918);
nand U17805 (N_17805,N_10713,N_14197);
and U17806 (N_17806,N_14305,N_10880);
or U17807 (N_17807,N_11899,N_14684);
and U17808 (N_17808,N_13642,N_13017);
or U17809 (N_17809,N_13465,N_13726);
nor U17810 (N_17810,N_10941,N_11991);
nor U17811 (N_17811,N_10321,N_12183);
or U17812 (N_17812,N_13313,N_11597);
xnor U17813 (N_17813,N_14479,N_10271);
nor U17814 (N_17814,N_13553,N_12717);
or U17815 (N_17815,N_10232,N_10655);
or U17816 (N_17816,N_11043,N_12887);
and U17817 (N_17817,N_11083,N_11477);
and U17818 (N_17818,N_12186,N_14685);
nor U17819 (N_17819,N_10510,N_10044);
and U17820 (N_17820,N_14404,N_14511);
or U17821 (N_17821,N_14537,N_10761);
nor U17822 (N_17822,N_14367,N_10886);
nor U17823 (N_17823,N_14343,N_13864);
nand U17824 (N_17824,N_12229,N_12198);
xor U17825 (N_17825,N_14741,N_13213);
nor U17826 (N_17826,N_11625,N_10032);
and U17827 (N_17827,N_14378,N_10810);
nor U17828 (N_17828,N_10016,N_14552);
xor U17829 (N_17829,N_14211,N_11401);
and U17830 (N_17830,N_10734,N_12183);
nor U17831 (N_17831,N_11707,N_12847);
nand U17832 (N_17832,N_12382,N_14080);
and U17833 (N_17833,N_11869,N_13007);
nor U17834 (N_17834,N_12085,N_13282);
and U17835 (N_17835,N_11093,N_12244);
or U17836 (N_17836,N_12159,N_12545);
nand U17837 (N_17837,N_11115,N_10563);
nor U17838 (N_17838,N_11808,N_12636);
nand U17839 (N_17839,N_12214,N_13387);
nor U17840 (N_17840,N_13632,N_14877);
and U17841 (N_17841,N_11282,N_11023);
or U17842 (N_17842,N_13020,N_13400);
and U17843 (N_17843,N_12392,N_11095);
or U17844 (N_17844,N_12199,N_13057);
nand U17845 (N_17845,N_12673,N_12679);
or U17846 (N_17846,N_13317,N_13000);
xor U17847 (N_17847,N_10363,N_13906);
or U17848 (N_17848,N_10289,N_12622);
and U17849 (N_17849,N_12431,N_14434);
nor U17850 (N_17850,N_11447,N_12890);
nand U17851 (N_17851,N_10056,N_12826);
nor U17852 (N_17852,N_14867,N_12747);
nor U17853 (N_17853,N_14431,N_10824);
and U17854 (N_17854,N_11267,N_11640);
xnor U17855 (N_17855,N_14448,N_10963);
nor U17856 (N_17856,N_12984,N_12391);
xor U17857 (N_17857,N_10164,N_13924);
and U17858 (N_17858,N_12000,N_10286);
nor U17859 (N_17859,N_10227,N_12467);
nand U17860 (N_17860,N_12877,N_13497);
nand U17861 (N_17861,N_12658,N_10048);
or U17862 (N_17862,N_14978,N_12980);
or U17863 (N_17863,N_10622,N_11978);
nor U17864 (N_17864,N_14133,N_13678);
nand U17865 (N_17865,N_13690,N_13883);
nand U17866 (N_17866,N_12134,N_14774);
and U17867 (N_17867,N_14626,N_13065);
or U17868 (N_17868,N_14950,N_14597);
or U17869 (N_17869,N_14236,N_14107);
nand U17870 (N_17870,N_10985,N_13364);
nand U17871 (N_17871,N_13845,N_13715);
nand U17872 (N_17872,N_10074,N_14171);
nor U17873 (N_17873,N_14233,N_12699);
nand U17874 (N_17874,N_11999,N_12927);
and U17875 (N_17875,N_13710,N_14338);
or U17876 (N_17876,N_13412,N_11352);
nor U17877 (N_17877,N_12617,N_11876);
or U17878 (N_17878,N_10903,N_10212);
or U17879 (N_17879,N_12514,N_10035);
xor U17880 (N_17880,N_10948,N_12060);
nor U17881 (N_17881,N_11904,N_11336);
nand U17882 (N_17882,N_11494,N_11242);
nor U17883 (N_17883,N_10974,N_13883);
xnor U17884 (N_17884,N_12336,N_11248);
nor U17885 (N_17885,N_10662,N_11905);
or U17886 (N_17886,N_12846,N_10739);
and U17887 (N_17887,N_14782,N_12589);
nand U17888 (N_17888,N_12512,N_10770);
nor U17889 (N_17889,N_10865,N_12871);
nor U17890 (N_17890,N_12313,N_12919);
and U17891 (N_17891,N_13569,N_10135);
nor U17892 (N_17892,N_11154,N_14920);
nor U17893 (N_17893,N_13056,N_11428);
nor U17894 (N_17894,N_11704,N_12367);
or U17895 (N_17895,N_13233,N_10287);
or U17896 (N_17896,N_13162,N_13827);
nand U17897 (N_17897,N_14292,N_13193);
or U17898 (N_17898,N_11960,N_12860);
and U17899 (N_17899,N_10442,N_11529);
nor U17900 (N_17900,N_13087,N_13458);
or U17901 (N_17901,N_12375,N_12551);
or U17902 (N_17902,N_12740,N_11797);
and U17903 (N_17903,N_10019,N_14794);
nor U17904 (N_17904,N_12007,N_13486);
or U17905 (N_17905,N_11635,N_10998);
nand U17906 (N_17906,N_14733,N_14517);
nor U17907 (N_17907,N_12711,N_12152);
or U17908 (N_17908,N_13150,N_12974);
nor U17909 (N_17909,N_11794,N_12498);
or U17910 (N_17910,N_12979,N_14825);
nand U17911 (N_17911,N_12481,N_11643);
nand U17912 (N_17912,N_12734,N_10900);
or U17913 (N_17913,N_10003,N_13665);
nand U17914 (N_17914,N_14956,N_11055);
or U17915 (N_17915,N_11115,N_13757);
or U17916 (N_17916,N_10828,N_13957);
nand U17917 (N_17917,N_11844,N_12204);
or U17918 (N_17918,N_13888,N_11175);
nor U17919 (N_17919,N_14096,N_10773);
nor U17920 (N_17920,N_11631,N_13648);
nand U17921 (N_17921,N_14089,N_10740);
nor U17922 (N_17922,N_13991,N_10080);
and U17923 (N_17923,N_10796,N_14665);
or U17924 (N_17924,N_10713,N_11739);
or U17925 (N_17925,N_12926,N_10237);
nor U17926 (N_17926,N_10358,N_14990);
and U17927 (N_17927,N_12455,N_11873);
nor U17928 (N_17928,N_11802,N_13904);
nand U17929 (N_17929,N_13075,N_10471);
nand U17930 (N_17930,N_14371,N_10919);
and U17931 (N_17931,N_10126,N_12158);
nor U17932 (N_17932,N_11663,N_14050);
or U17933 (N_17933,N_12173,N_13247);
xor U17934 (N_17934,N_14533,N_13137);
and U17935 (N_17935,N_14232,N_14201);
nor U17936 (N_17936,N_14374,N_11562);
and U17937 (N_17937,N_10615,N_11108);
or U17938 (N_17938,N_13847,N_12939);
and U17939 (N_17939,N_10679,N_13788);
or U17940 (N_17940,N_11706,N_11433);
nand U17941 (N_17941,N_11153,N_13722);
and U17942 (N_17942,N_14866,N_10681);
or U17943 (N_17943,N_11851,N_12797);
nand U17944 (N_17944,N_11883,N_11063);
and U17945 (N_17945,N_14118,N_13137);
xnor U17946 (N_17946,N_10932,N_11992);
nor U17947 (N_17947,N_13404,N_14689);
nand U17948 (N_17948,N_10576,N_14543);
nand U17949 (N_17949,N_11748,N_13880);
and U17950 (N_17950,N_13650,N_14251);
nor U17951 (N_17951,N_14732,N_14579);
nand U17952 (N_17952,N_13419,N_10679);
or U17953 (N_17953,N_14468,N_10196);
nor U17954 (N_17954,N_11339,N_12035);
nor U17955 (N_17955,N_12427,N_13429);
nor U17956 (N_17956,N_13001,N_14532);
nor U17957 (N_17957,N_11819,N_13551);
nand U17958 (N_17958,N_10799,N_14896);
nand U17959 (N_17959,N_14178,N_10537);
nor U17960 (N_17960,N_14669,N_14157);
nand U17961 (N_17961,N_10906,N_10088);
nor U17962 (N_17962,N_12853,N_10318);
and U17963 (N_17963,N_13499,N_10622);
xor U17964 (N_17964,N_14189,N_13328);
nor U17965 (N_17965,N_11029,N_10134);
and U17966 (N_17966,N_14467,N_14601);
nor U17967 (N_17967,N_11196,N_10023);
xor U17968 (N_17968,N_13483,N_13245);
nor U17969 (N_17969,N_12651,N_13794);
xnor U17970 (N_17970,N_14372,N_12692);
nor U17971 (N_17971,N_14426,N_13239);
and U17972 (N_17972,N_11313,N_13771);
nor U17973 (N_17973,N_13388,N_11221);
and U17974 (N_17974,N_11915,N_13855);
xor U17975 (N_17975,N_14098,N_11213);
nand U17976 (N_17976,N_10765,N_13937);
xor U17977 (N_17977,N_13289,N_12542);
nand U17978 (N_17978,N_12918,N_13948);
or U17979 (N_17979,N_14173,N_10957);
or U17980 (N_17980,N_11065,N_12967);
nand U17981 (N_17981,N_14295,N_14584);
nand U17982 (N_17982,N_13579,N_14061);
xor U17983 (N_17983,N_10328,N_12287);
and U17984 (N_17984,N_11693,N_12719);
nand U17985 (N_17985,N_13956,N_12122);
nand U17986 (N_17986,N_10844,N_12624);
nand U17987 (N_17987,N_14696,N_12519);
xor U17988 (N_17988,N_13015,N_13619);
and U17989 (N_17989,N_14871,N_14700);
nor U17990 (N_17990,N_13988,N_14106);
xor U17991 (N_17991,N_13056,N_11348);
xnor U17992 (N_17992,N_11826,N_12714);
nand U17993 (N_17993,N_14991,N_14047);
nand U17994 (N_17994,N_14901,N_12977);
and U17995 (N_17995,N_13463,N_14105);
nor U17996 (N_17996,N_10872,N_14744);
nor U17997 (N_17997,N_12673,N_14671);
xor U17998 (N_17998,N_13122,N_14132);
and U17999 (N_17999,N_13820,N_12609);
and U18000 (N_18000,N_13914,N_14410);
nor U18001 (N_18001,N_11789,N_14536);
nor U18002 (N_18002,N_12902,N_14263);
nand U18003 (N_18003,N_12747,N_14053);
nand U18004 (N_18004,N_13047,N_12142);
or U18005 (N_18005,N_14425,N_12925);
xor U18006 (N_18006,N_11045,N_13115);
and U18007 (N_18007,N_14533,N_10058);
nand U18008 (N_18008,N_12729,N_11550);
and U18009 (N_18009,N_12133,N_11565);
nor U18010 (N_18010,N_12048,N_14907);
or U18011 (N_18011,N_10239,N_10851);
xnor U18012 (N_18012,N_14759,N_13723);
xor U18013 (N_18013,N_13903,N_12286);
or U18014 (N_18014,N_12575,N_14914);
and U18015 (N_18015,N_12177,N_13203);
xnor U18016 (N_18016,N_13363,N_12738);
nand U18017 (N_18017,N_14977,N_13039);
or U18018 (N_18018,N_10826,N_13520);
or U18019 (N_18019,N_12403,N_13660);
and U18020 (N_18020,N_12965,N_14387);
nor U18021 (N_18021,N_11542,N_13934);
and U18022 (N_18022,N_14055,N_14968);
xor U18023 (N_18023,N_12052,N_10594);
or U18024 (N_18024,N_13682,N_10113);
nor U18025 (N_18025,N_13949,N_11924);
nand U18026 (N_18026,N_14804,N_10769);
nand U18027 (N_18027,N_10839,N_10671);
nor U18028 (N_18028,N_11436,N_13849);
nor U18029 (N_18029,N_12048,N_13090);
and U18030 (N_18030,N_13567,N_14315);
or U18031 (N_18031,N_11942,N_11999);
nand U18032 (N_18032,N_13150,N_12960);
and U18033 (N_18033,N_13914,N_14777);
or U18034 (N_18034,N_14400,N_12657);
or U18035 (N_18035,N_13149,N_10586);
nand U18036 (N_18036,N_12479,N_10641);
and U18037 (N_18037,N_13677,N_14135);
or U18038 (N_18038,N_12084,N_10370);
nor U18039 (N_18039,N_11602,N_12454);
or U18040 (N_18040,N_10325,N_13889);
nand U18041 (N_18041,N_13181,N_12055);
xnor U18042 (N_18042,N_12784,N_11616);
nor U18043 (N_18043,N_13124,N_10183);
or U18044 (N_18044,N_10247,N_10791);
nand U18045 (N_18045,N_14232,N_14619);
nand U18046 (N_18046,N_11903,N_13790);
nor U18047 (N_18047,N_12635,N_10549);
xnor U18048 (N_18048,N_13750,N_12280);
and U18049 (N_18049,N_13325,N_11270);
and U18050 (N_18050,N_11035,N_11640);
nor U18051 (N_18051,N_13465,N_14841);
xnor U18052 (N_18052,N_12572,N_11439);
or U18053 (N_18053,N_10623,N_11108);
or U18054 (N_18054,N_12558,N_11414);
nand U18055 (N_18055,N_11540,N_12949);
and U18056 (N_18056,N_14375,N_11875);
nor U18057 (N_18057,N_11532,N_10020);
and U18058 (N_18058,N_10526,N_11718);
nor U18059 (N_18059,N_10024,N_11962);
nand U18060 (N_18060,N_11198,N_13332);
and U18061 (N_18061,N_13072,N_13091);
and U18062 (N_18062,N_10677,N_14961);
nand U18063 (N_18063,N_14760,N_10618);
nor U18064 (N_18064,N_13166,N_14301);
nand U18065 (N_18065,N_13666,N_12652);
and U18066 (N_18066,N_12189,N_11809);
nor U18067 (N_18067,N_11575,N_13484);
or U18068 (N_18068,N_10677,N_12355);
and U18069 (N_18069,N_12518,N_12408);
or U18070 (N_18070,N_14242,N_12876);
or U18071 (N_18071,N_10546,N_11607);
xor U18072 (N_18072,N_10068,N_13238);
or U18073 (N_18073,N_10070,N_12156);
nand U18074 (N_18074,N_14575,N_11486);
xor U18075 (N_18075,N_11578,N_12378);
nand U18076 (N_18076,N_11342,N_10360);
or U18077 (N_18077,N_12600,N_13988);
or U18078 (N_18078,N_10081,N_11989);
nor U18079 (N_18079,N_14445,N_10069);
or U18080 (N_18080,N_14426,N_11227);
and U18081 (N_18081,N_13356,N_10864);
or U18082 (N_18082,N_10378,N_14367);
nor U18083 (N_18083,N_14430,N_10645);
and U18084 (N_18084,N_14288,N_14868);
nand U18085 (N_18085,N_13999,N_10305);
xnor U18086 (N_18086,N_12289,N_14424);
or U18087 (N_18087,N_11131,N_11856);
and U18088 (N_18088,N_12696,N_13514);
and U18089 (N_18089,N_10168,N_13732);
xor U18090 (N_18090,N_13600,N_12797);
nor U18091 (N_18091,N_13582,N_13567);
nand U18092 (N_18092,N_14196,N_14898);
xnor U18093 (N_18093,N_10466,N_12712);
nand U18094 (N_18094,N_10346,N_13217);
nand U18095 (N_18095,N_12442,N_11092);
nand U18096 (N_18096,N_13141,N_13628);
nand U18097 (N_18097,N_14625,N_10864);
and U18098 (N_18098,N_13104,N_10580);
and U18099 (N_18099,N_10890,N_14941);
or U18100 (N_18100,N_14644,N_13668);
and U18101 (N_18101,N_10963,N_10783);
nand U18102 (N_18102,N_13988,N_12754);
nor U18103 (N_18103,N_12224,N_12835);
and U18104 (N_18104,N_12554,N_11722);
nor U18105 (N_18105,N_14304,N_12275);
or U18106 (N_18106,N_12556,N_12851);
and U18107 (N_18107,N_10186,N_14868);
or U18108 (N_18108,N_12812,N_13669);
or U18109 (N_18109,N_14089,N_10452);
or U18110 (N_18110,N_14512,N_14624);
and U18111 (N_18111,N_10103,N_14138);
nor U18112 (N_18112,N_12696,N_14977);
and U18113 (N_18113,N_12548,N_11149);
nand U18114 (N_18114,N_14400,N_10066);
or U18115 (N_18115,N_10906,N_12229);
nand U18116 (N_18116,N_11256,N_13668);
and U18117 (N_18117,N_10545,N_13478);
and U18118 (N_18118,N_13884,N_12574);
xor U18119 (N_18119,N_11695,N_13706);
or U18120 (N_18120,N_13418,N_13477);
and U18121 (N_18121,N_14992,N_12021);
or U18122 (N_18122,N_14514,N_12855);
and U18123 (N_18123,N_13728,N_13656);
nor U18124 (N_18124,N_12541,N_12937);
xnor U18125 (N_18125,N_11883,N_10851);
and U18126 (N_18126,N_10941,N_13892);
nand U18127 (N_18127,N_11633,N_10505);
nor U18128 (N_18128,N_11002,N_13093);
and U18129 (N_18129,N_14298,N_11598);
nand U18130 (N_18130,N_10722,N_13438);
nand U18131 (N_18131,N_13281,N_10591);
and U18132 (N_18132,N_12107,N_10251);
or U18133 (N_18133,N_11584,N_13301);
and U18134 (N_18134,N_10100,N_13487);
nor U18135 (N_18135,N_10805,N_12265);
nor U18136 (N_18136,N_14634,N_12744);
nand U18137 (N_18137,N_12564,N_14891);
or U18138 (N_18138,N_10757,N_12171);
nand U18139 (N_18139,N_11991,N_12955);
or U18140 (N_18140,N_14243,N_10383);
nor U18141 (N_18141,N_13686,N_12244);
and U18142 (N_18142,N_10568,N_14357);
and U18143 (N_18143,N_11122,N_12696);
xnor U18144 (N_18144,N_14707,N_12543);
and U18145 (N_18145,N_13680,N_10241);
or U18146 (N_18146,N_12328,N_12661);
and U18147 (N_18147,N_14143,N_12187);
nand U18148 (N_18148,N_11514,N_10099);
nor U18149 (N_18149,N_11167,N_12957);
nand U18150 (N_18150,N_11551,N_13932);
or U18151 (N_18151,N_11236,N_12653);
nor U18152 (N_18152,N_12718,N_12581);
nand U18153 (N_18153,N_14264,N_10531);
and U18154 (N_18154,N_12939,N_13777);
or U18155 (N_18155,N_12089,N_14374);
nand U18156 (N_18156,N_11382,N_12355);
nor U18157 (N_18157,N_11145,N_13445);
nand U18158 (N_18158,N_10530,N_10137);
and U18159 (N_18159,N_13291,N_10424);
xor U18160 (N_18160,N_13983,N_12489);
xor U18161 (N_18161,N_13138,N_10393);
or U18162 (N_18162,N_12494,N_14002);
or U18163 (N_18163,N_14965,N_12354);
nand U18164 (N_18164,N_11620,N_13922);
nand U18165 (N_18165,N_11169,N_11046);
and U18166 (N_18166,N_12375,N_13287);
and U18167 (N_18167,N_10582,N_12356);
xor U18168 (N_18168,N_11819,N_14412);
xnor U18169 (N_18169,N_12445,N_10415);
nand U18170 (N_18170,N_13274,N_13800);
nand U18171 (N_18171,N_14099,N_11704);
xnor U18172 (N_18172,N_11707,N_11221);
nand U18173 (N_18173,N_10798,N_10272);
or U18174 (N_18174,N_10336,N_14752);
nor U18175 (N_18175,N_14438,N_12386);
nand U18176 (N_18176,N_14260,N_14276);
and U18177 (N_18177,N_12939,N_12679);
nor U18178 (N_18178,N_13498,N_12257);
and U18179 (N_18179,N_13658,N_14550);
or U18180 (N_18180,N_12167,N_12100);
nand U18181 (N_18181,N_12394,N_11762);
nor U18182 (N_18182,N_11228,N_11552);
nand U18183 (N_18183,N_13078,N_12401);
nand U18184 (N_18184,N_13870,N_13016);
or U18185 (N_18185,N_13078,N_13280);
nor U18186 (N_18186,N_13397,N_14290);
nor U18187 (N_18187,N_13861,N_10558);
xnor U18188 (N_18188,N_10992,N_12183);
nor U18189 (N_18189,N_10245,N_11229);
nor U18190 (N_18190,N_11400,N_10531);
or U18191 (N_18191,N_11059,N_12684);
and U18192 (N_18192,N_14441,N_14411);
or U18193 (N_18193,N_11948,N_14323);
nand U18194 (N_18194,N_12652,N_14194);
nand U18195 (N_18195,N_10941,N_12061);
nand U18196 (N_18196,N_10689,N_10003);
xor U18197 (N_18197,N_13840,N_11325);
or U18198 (N_18198,N_12743,N_13453);
or U18199 (N_18199,N_13429,N_11870);
or U18200 (N_18200,N_10629,N_12450);
nand U18201 (N_18201,N_14481,N_13217);
xor U18202 (N_18202,N_13045,N_12624);
and U18203 (N_18203,N_12254,N_12299);
and U18204 (N_18204,N_14408,N_14700);
and U18205 (N_18205,N_14801,N_14489);
and U18206 (N_18206,N_10631,N_13024);
or U18207 (N_18207,N_12402,N_12941);
and U18208 (N_18208,N_10044,N_10681);
nor U18209 (N_18209,N_10552,N_11048);
and U18210 (N_18210,N_13227,N_12315);
nand U18211 (N_18211,N_14061,N_11627);
xnor U18212 (N_18212,N_10742,N_11691);
or U18213 (N_18213,N_13524,N_14565);
or U18214 (N_18214,N_12680,N_10217);
nor U18215 (N_18215,N_10342,N_11362);
nand U18216 (N_18216,N_13314,N_12639);
nor U18217 (N_18217,N_10801,N_13934);
nand U18218 (N_18218,N_10682,N_13851);
xor U18219 (N_18219,N_13195,N_10771);
or U18220 (N_18220,N_14123,N_13372);
and U18221 (N_18221,N_11367,N_10425);
or U18222 (N_18222,N_12431,N_10448);
nand U18223 (N_18223,N_13919,N_13764);
xnor U18224 (N_18224,N_12618,N_11803);
nand U18225 (N_18225,N_10337,N_11805);
and U18226 (N_18226,N_13785,N_14919);
xnor U18227 (N_18227,N_14790,N_11528);
and U18228 (N_18228,N_14419,N_11196);
xnor U18229 (N_18229,N_13194,N_14743);
and U18230 (N_18230,N_11976,N_10467);
nand U18231 (N_18231,N_12309,N_14609);
nor U18232 (N_18232,N_11489,N_12223);
and U18233 (N_18233,N_12512,N_14324);
and U18234 (N_18234,N_11026,N_14050);
or U18235 (N_18235,N_12265,N_13444);
and U18236 (N_18236,N_11270,N_12223);
nor U18237 (N_18237,N_12012,N_13918);
and U18238 (N_18238,N_11956,N_12306);
or U18239 (N_18239,N_11795,N_10035);
nand U18240 (N_18240,N_14397,N_11592);
nor U18241 (N_18241,N_10910,N_11889);
nand U18242 (N_18242,N_13228,N_11619);
or U18243 (N_18243,N_10715,N_12838);
nor U18244 (N_18244,N_11239,N_12452);
nor U18245 (N_18245,N_11046,N_13454);
or U18246 (N_18246,N_12783,N_13845);
and U18247 (N_18247,N_12754,N_13216);
nand U18248 (N_18248,N_13930,N_11556);
nor U18249 (N_18249,N_10940,N_14048);
nand U18250 (N_18250,N_13131,N_14479);
or U18251 (N_18251,N_12468,N_14202);
or U18252 (N_18252,N_13623,N_14647);
and U18253 (N_18253,N_10390,N_12961);
or U18254 (N_18254,N_12497,N_10318);
or U18255 (N_18255,N_12472,N_11642);
or U18256 (N_18256,N_11931,N_10865);
or U18257 (N_18257,N_14165,N_10057);
and U18258 (N_18258,N_11467,N_10679);
and U18259 (N_18259,N_13873,N_14338);
and U18260 (N_18260,N_10129,N_11089);
or U18261 (N_18261,N_11449,N_12352);
nor U18262 (N_18262,N_10478,N_10851);
nor U18263 (N_18263,N_14840,N_11633);
or U18264 (N_18264,N_10877,N_13905);
nor U18265 (N_18265,N_12693,N_11695);
and U18266 (N_18266,N_13596,N_12498);
nor U18267 (N_18267,N_11632,N_14046);
and U18268 (N_18268,N_10862,N_13015);
xnor U18269 (N_18269,N_11351,N_12178);
nor U18270 (N_18270,N_12158,N_13807);
and U18271 (N_18271,N_14477,N_13142);
nand U18272 (N_18272,N_12104,N_13269);
nor U18273 (N_18273,N_10643,N_12161);
and U18274 (N_18274,N_11684,N_10771);
nand U18275 (N_18275,N_11114,N_12900);
and U18276 (N_18276,N_14222,N_14512);
nand U18277 (N_18277,N_12846,N_14473);
and U18278 (N_18278,N_10031,N_14369);
and U18279 (N_18279,N_11036,N_13051);
or U18280 (N_18280,N_13141,N_10614);
or U18281 (N_18281,N_14343,N_11623);
or U18282 (N_18282,N_13252,N_10978);
or U18283 (N_18283,N_10497,N_11316);
nand U18284 (N_18284,N_13179,N_10409);
nor U18285 (N_18285,N_10314,N_13105);
or U18286 (N_18286,N_10103,N_11064);
nor U18287 (N_18287,N_11832,N_11304);
and U18288 (N_18288,N_14642,N_14975);
nor U18289 (N_18289,N_12305,N_12985);
or U18290 (N_18290,N_13908,N_11411);
and U18291 (N_18291,N_13200,N_12760);
and U18292 (N_18292,N_11826,N_14938);
xnor U18293 (N_18293,N_13534,N_10003);
nor U18294 (N_18294,N_12686,N_10745);
or U18295 (N_18295,N_12223,N_14976);
nand U18296 (N_18296,N_13373,N_10873);
or U18297 (N_18297,N_14961,N_10392);
xnor U18298 (N_18298,N_11712,N_12986);
nor U18299 (N_18299,N_13052,N_10735);
nor U18300 (N_18300,N_13649,N_11454);
nor U18301 (N_18301,N_12741,N_13974);
or U18302 (N_18302,N_14361,N_12706);
nand U18303 (N_18303,N_11492,N_10582);
and U18304 (N_18304,N_14857,N_12400);
xor U18305 (N_18305,N_10110,N_12875);
or U18306 (N_18306,N_11355,N_10821);
nor U18307 (N_18307,N_14216,N_13892);
or U18308 (N_18308,N_12138,N_11593);
and U18309 (N_18309,N_13742,N_11154);
or U18310 (N_18310,N_14712,N_12550);
and U18311 (N_18311,N_13212,N_11607);
nor U18312 (N_18312,N_14934,N_11481);
or U18313 (N_18313,N_14902,N_12087);
and U18314 (N_18314,N_10058,N_10638);
nor U18315 (N_18315,N_11196,N_14268);
or U18316 (N_18316,N_13102,N_11679);
nand U18317 (N_18317,N_10324,N_13070);
nand U18318 (N_18318,N_12447,N_14391);
nor U18319 (N_18319,N_10946,N_10959);
or U18320 (N_18320,N_10589,N_14223);
nand U18321 (N_18321,N_11198,N_10672);
xnor U18322 (N_18322,N_11553,N_12093);
nand U18323 (N_18323,N_10060,N_14780);
and U18324 (N_18324,N_14382,N_10427);
nor U18325 (N_18325,N_10141,N_14319);
or U18326 (N_18326,N_11813,N_14500);
xnor U18327 (N_18327,N_10157,N_12408);
nor U18328 (N_18328,N_10184,N_12419);
nor U18329 (N_18329,N_14510,N_12267);
nor U18330 (N_18330,N_12868,N_12809);
and U18331 (N_18331,N_13567,N_10685);
xnor U18332 (N_18332,N_12017,N_11141);
nand U18333 (N_18333,N_11345,N_11174);
and U18334 (N_18334,N_13501,N_13736);
or U18335 (N_18335,N_10357,N_12160);
and U18336 (N_18336,N_10581,N_13555);
and U18337 (N_18337,N_11952,N_12805);
or U18338 (N_18338,N_10847,N_10261);
nand U18339 (N_18339,N_14004,N_13074);
nand U18340 (N_18340,N_11983,N_11453);
or U18341 (N_18341,N_11397,N_14629);
nor U18342 (N_18342,N_14740,N_12620);
or U18343 (N_18343,N_11346,N_12895);
nand U18344 (N_18344,N_13197,N_14790);
nor U18345 (N_18345,N_12172,N_10848);
nand U18346 (N_18346,N_14287,N_12226);
nor U18347 (N_18347,N_12266,N_13643);
or U18348 (N_18348,N_11091,N_14190);
nand U18349 (N_18349,N_12962,N_13224);
nand U18350 (N_18350,N_13563,N_12915);
nor U18351 (N_18351,N_13673,N_12756);
or U18352 (N_18352,N_11248,N_12466);
and U18353 (N_18353,N_11915,N_10423);
or U18354 (N_18354,N_12935,N_13843);
nand U18355 (N_18355,N_12995,N_14417);
nor U18356 (N_18356,N_14755,N_13789);
or U18357 (N_18357,N_14122,N_10380);
or U18358 (N_18358,N_13123,N_14911);
or U18359 (N_18359,N_14837,N_10987);
nand U18360 (N_18360,N_10960,N_13050);
nand U18361 (N_18361,N_12169,N_11583);
nand U18362 (N_18362,N_11448,N_14423);
nor U18363 (N_18363,N_14667,N_13510);
nand U18364 (N_18364,N_11718,N_13020);
nand U18365 (N_18365,N_11684,N_10246);
nand U18366 (N_18366,N_12052,N_12773);
nor U18367 (N_18367,N_10175,N_13300);
nor U18368 (N_18368,N_13394,N_14852);
and U18369 (N_18369,N_14067,N_14104);
xnor U18370 (N_18370,N_10337,N_10393);
and U18371 (N_18371,N_12593,N_14880);
nand U18372 (N_18372,N_14184,N_10985);
or U18373 (N_18373,N_13684,N_11876);
nor U18374 (N_18374,N_14942,N_13536);
and U18375 (N_18375,N_11575,N_13252);
and U18376 (N_18376,N_12778,N_12467);
nor U18377 (N_18377,N_10517,N_14515);
nor U18378 (N_18378,N_12463,N_10202);
nor U18379 (N_18379,N_12690,N_11159);
and U18380 (N_18380,N_10428,N_11024);
nor U18381 (N_18381,N_14304,N_13023);
or U18382 (N_18382,N_13644,N_12916);
nor U18383 (N_18383,N_14196,N_14713);
or U18384 (N_18384,N_14946,N_11554);
nand U18385 (N_18385,N_13225,N_14898);
and U18386 (N_18386,N_12607,N_14018);
nand U18387 (N_18387,N_14431,N_11360);
xor U18388 (N_18388,N_14334,N_10882);
or U18389 (N_18389,N_12595,N_13954);
xor U18390 (N_18390,N_10845,N_10816);
and U18391 (N_18391,N_13302,N_14640);
xor U18392 (N_18392,N_10229,N_10917);
and U18393 (N_18393,N_14862,N_11439);
nand U18394 (N_18394,N_13365,N_12462);
nand U18395 (N_18395,N_13704,N_10764);
nand U18396 (N_18396,N_11628,N_12642);
and U18397 (N_18397,N_10748,N_12388);
nor U18398 (N_18398,N_10025,N_13540);
nor U18399 (N_18399,N_10375,N_13842);
nor U18400 (N_18400,N_11657,N_10999);
nor U18401 (N_18401,N_10249,N_11952);
and U18402 (N_18402,N_12795,N_14778);
nand U18403 (N_18403,N_12471,N_12973);
or U18404 (N_18404,N_12915,N_12989);
nand U18405 (N_18405,N_13407,N_13428);
and U18406 (N_18406,N_14607,N_11503);
nor U18407 (N_18407,N_14277,N_11740);
xnor U18408 (N_18408,N_12363,N_13019);
or U18409 (N_18409,N_13387,N_10536);
xor U18410 (N_18410,N_14141,N_11767);
and U18411 (N_18411,N_14574,N_10092);
nor U18412 (N_18412,N_13604,N_11156);
and U18413 (N_18413,N_12356,N_12152);
nand U18414 (N_18414,N_14054,N_11035);
nor U18415 (N_18415,N_14179,N_11352);
nor U18416 (N_18416,N_13634,N_13102);
nor U18417 (N_18417,N_14225,N_14207);
nor U18418 (N_18418,N_12424,N_13629);
xnor U18419 (N_18419,N_10327,N_12562);
xnor U18420 (N_18420,N_12082,N_13106);
nand U18421 (N_18421,N_10644,N_13733);
nand U18422 (N_18422,N_11269,N_10940);
and U18423 (N_18423,N_10069,N_10018);
nor U18424 (N_18424,N_11205,N_10666);
nor U18425 (N_18425,N_13093,N_13137);
nand U18426 (N_18426,N_13862,N_14544);
and U18427 (N_18427,N_11619,N_11518);
and U18428 (N_18428,N_12557,N_14330);
and U18429 (N_18429,N_13678,N_13407);
or U18430 (N_18430,N_11736,N_12448);
nor U18431 (N_18431,N_12364,N_13415);
nand U18432 (N_18432,N_10647,N_12730);
or U18433 (N_18433,N_13304,N_14496);
and U18434 (N_18434,N_12769,N_14851);
nor U18435 (N_18435,N_12254,N_13040);
or U18436 (N_18436,N_12746,N_10420);
nor U18437 (N_18437,N_14083,N_13757);
or U18438 (N_18438,N_10082,N_12710);
or U18439 (N_18439,N_10347,N_14191);
xor U18440 (N_18440,N_13908,N_10187);
nand U18441 (N_18441,N_12727,N_12411);
xor U18442 (N_18442,N_10737,N_10883);
and U18443 (N_18443,N_14957,N_10820);
nor U18444 (N_18444,N_10834,N_13145);
nand U18445 (N_18445,N_10779,N_14633);
and U18446 (N_18446,N_14620,N_12662);
and U18447 (N_18447,N_13074,N_10906);
nand U18448 (N_18448,N_10185,N_12130);
nor U18449 (N_18449,N_10444,N_10020);
nor U18450 (N_18450,N_11797,N_12084);
nand U18451 (N_18451,N_11175,N_10242);
and U18452 (N_18452,N_10186,N_13479);
or U18453 (N_18453,N_14601,N_14453);
nor U18454 (N_18454,N_14144,N_14862);
nand U18455 (N_18455,N_14844,N_10546);
xor U18456 (N_18456,N_11766,N_10761);
nor U18457 (N_18457,N_10079,N_13567);
nor U18458 (N_18458,N_13967,N_14935);
nand U18459 (N_18459,N_13352,N_14128);
and U18460 (N_18460,N_11339,N_12932);
nor U18461 (N_18461,N_10748,N_10480);
or U18462 (N_18462,N_13541,N_11058);
nand U18463 (N_18463,N_14460,N_10240);
or U18464 (N_18464,N_12000,N_13232);
nand U18465 (N_18465,N_13756,N_12580);
and U18466 (N_18466,N_14100,N_14329);
or U18467 (N_18467,N_10005,N_13477);
nor U18468 (N_18468,N_11729,N_12026);
xnor U18469 (N_18469,N_12335,N_13306);
xor U18470 (N_18470,N_14650,N_14425);
nor U18471 (N_18471,N_11010,N_10277);
nand U18472 (N_18472,N_10181,N_12139);
and U18473 (N_18473,N_14954,N_11813);
and U18474 (N_18474,N_10854,N_14777);
and U18475 (N_18475,N_13958,N_13768);
nor U18476 (N_18476,N_13113,N_12468);
nor U18477 (N_18477,N_14535,N_11122);
nor U18478 (N_18478,N_12330,N_13189);
and U18479 (N_18479,N_10883,N_13934);
or U18480 (N_18480,N_14834,N_10722);
or U18481 (N_18481,N_10674,N_14545);
or U18482 (N_18482,N_12734,N_12683);
and U18483 (N_18483,N_11818,N_11237);
or U18484 (N_18484,N_11865,N_14474);
or U18485 (N_18485,N_14910,N_13040);
nand U18486 (N_18486,N_11316,N_14487);
nor U18487 (N_18487,N_13189,N_12914);
or U18488 (N_18488,N_13224,N_12957);
nand U18489 (N_18489,N_11840,N_11942);
nor U18490 (N_18490,N_10923,N_10695);
nand U18491 (N_18491,N_12373,N_13402);
nor U18492 (N_18492,N_12486,N_11493);
and U18493 (N_18493,N_10311,N_13793);
and U18494 (N_18494,N_13972,N_12316);
and U18495 (N_18495,N_12079,N_12460);
and U18496 (N_18496,N_13940,N_11022);
nand U18497 (N_18497,N_12162,N_10468);
nand U18498 (N_18498,N_12253,N_13313);
nor U18499 (N_18499,N_13834,N_11584);
nand U18500 (N_18500,N_14414,N_12929);
or U18501 (N_18501,N_11268,N_11211);
nor U18502 (N_18502,N_11992,N_10608);
nor U18503 (N_18503,N_14222,N_14397);
or U18504 (N_18504,N_13243,N_13798);
and U18505 (N_18505,N_10970,N_14528);
nand U18506 (N_18506,N_10494,N_10828);
or U18507 (N_18507,N_11333,N_10840);
nand U18508 (N_18508,N_13944,N_11539);
nor U18509 (N_18509,N_11551,N_11732);
and U18510 (N_18510,N_14895,N_11879);
nor U18511 (N_18511,N_13874,N_13110);
or U18512 (N_18512,N_13951,N_12634);
nor U18513 (N_18513,N_14189,N_14715);
nor U18514 (N_18514,N_12380,N_14884);
nor U18515 (N_18515,N_13789,N_10403);
nor U18516 (N_18516,N_13023,N_14325);
nand U18517 (N_18517,N_11020,N_14880);
and U18518 (N_18518,N_14349,N_10379);
xnor U18519 (N_18519,N_10450,N_11802);
or U18520 (N_18520,N_14253,N_12758);
nand U18521 (N_18521,N_10548,N_13599);
or U18522 (N_18522,N_10254,N_13083);
and U18523 (N_18523,N_10312,N_14191);
or U18524 (N_18524,N_13087,N_10577);
nand U18525 (N_18525,N_13823,N_12184);
nand U18526 (N_18526,N_13349,N_13820);
nand U18527 (N_18527,N_14487,N_10894);
nor U18528 (N_18528,N_12635,N_11555);
nand U18529 (N_18529,N_13776,N_10787);
nand U18530 (N_18530,N_13582,N_13034);
and U18531 (N_18531,N_13328,N_13248);
or U18532 (N_18532,N_10705,N_14240);
and U18533 (N_18533,N_13592,N_10294);
xnor U18534 (N_18534,N_11907,N_12399);
nand U18535 (N_18535,N_14784,N_10893);
nand U18536 (N_18536,N_14797,N_12775);
nand U18537 (N_18537,N_10779,N_14230);
nand U18538 (N_18538,N_12243,N_13402);
and U18539 (N_18539,N_12475,N_11835);
nor U18540 (N_18540,N_10767,N_11768);
nand U18541 (N_18541,N_14110,N_12635);
nand U18542 (N_18542,N_12420,N_14966);
nand U18543 (N_18543,N_13955,N_14435);
and U18544 (N_18544,N_11377,N_11364);
and U18545 (N_18545,N_13558,N_14050);
nor U18546 (N_18546,N_12765,N_13153);
and U18547 (N_18547,N_14698,N_14333);
or U18548 (N_18548,N_10320,N_12194);
xor U18549 (N_18549,N_10131,N_12866);
nor U18550 (N_18550,N_11131,N_10198);
nor U18551 (N_18551,N_14857,N_10945);
and U18552 (N_18552,N_10249,N_14478);
nor U18553 (N_18553,N_11085,N_13265);
nor U18554 (N_18554,N_12649,N_14800);
nor U18555 (N_18555,N_11725,N_10641);
nor U18556 (N_18556,N_11521,N_13424);
or U18557 (N_18557,N_11886,N_14439);
xnor U18558 (N_18558,N_10774,N_13257);
nor U18559 (N_18559,N_12258,N_14470);
xnor U18560 (N_18560,N_14878,N_13344);
or U18561 (N_18561,N_10290,N_14068);
xnor U18562 (N_18562,N_12161,N_11474);
xnor U18563 (N_18563,N_10582,N_12699);
or U18564 (N_18564,N_13713,N_13633);
nor U18565 (N_18565,N_14215,N_14581);
and U18566 (N_18566,N_13773,N_10849);
and U18567 (N_18567,N_12057,N_14242);
xnor U18568 (N_18568,N_13665,N_12737);
nand U18569 (N_18569,N_12406,N_12564);
xnor U18570 (N_18570,N_12467,N_13595);
xor U18571 (N_18571,N_13174,N_13198);
and U18572 (N_18572,N_14639,N_14262);
nor U18573 (N_18573,N_14594,N_13456);
nand U18574 (N_18574,N_14293,N_12324);
or U18575 (N_18575,N_10432,N_14727);
or U18576 (N_18576,N_14013,N_14353);
xor U18577 (N_18577,N_12530,N_11996);
nor U18578 (N_18578,N_12613,N_13599);
and U18579 (N_18579,N_12848,N_13952);
or U18580 (N_18580,N_13743,N_13917);
and U18581 (N_18581,N_13542,N_13393);
nand U18582 (N_18582,N_12148,N_12809);
xor U18583 (N_18583,N_11597,N_10219);
nor U18584 (N_18584,N_13535,N_11542);
and U18585 (N_18585,N_14149,N_11948);
nand U18586 (N_18586,N_13913,N_13796);
or U18587 (N_18587,N_14237,N_11064);
nand U18588 (N_18588,N_12209,N_10897);
nor U18589 (N_18589,N_11740,N_13052);
nor U18590 (N_18590,N_14539,N_10916);
and U18591 (N_18591,N_13816,N_12962);
xor U18592 (N_18592,N_13197,N_12340);
nand U18593 (N_18593,N_14022,N_10485);
and U18594 (N_18594,N_11971,N_14764);
or U18595 (N_18595,N_13920,N_14076);
nor U18596 (N_18596,N_12028,N_10717);
and U18597 (N_18597,N_10355,N_10082);
or U18598 (N_18598,N_11458,N_12058);
xor U18599 (N_18599,N_13494,N_10933);
or U18600 (N_18600,N_14704,N_11676);
nor U18601 (N_18601,N_11346,N_14924);
nand U18602 (N_18602,N_11139,N_12223);
or U18603 (N_18603,N_12010,N_13933);
and U18604 (N_18604,N_10018,N_12470);
xor U18605 (N_18605,N_12530,N_13613);
xor U18606 (N_18606,N_14735,N_10961);
nor U18607 (N_18607,N_13189,N_12379);
nor U18608 (N_18608,N_11385,N_10567);
or U18609 (N_18609,N_11803,N_11615);
xnor U18610 (N_18610,N_13970,N_12140);
nand U18611 (N_18611,N_12571,N_14040);
nor U18612 (N_18612,N_10548,N_13330);
nor U18613 (N_18613,N_11247,N_11329);
nor U18614 (N_18614,N_10877,N_13869);
nand U18615 (N_18615,N_10854,N_10441);
nor U18616 (N_18616,N_13305,N_14230);
nand U18617 (N_18617,N_12140,N_11433);
or U18618 (N_18618,N_12007,N_11038);
or U18619 (N_18619,N_14718,N_12068);
or U18620 (N_18620,N_11514,N_11049);
or U18621 (N_18621,N_14212,N_10675);
and U18622 (N_18622,N_11667,N_10067);
or U18623 (N_18623,N_11611,N_10233);
or U18624 (N_18624,N_11155,N_10783);
or U18625 (N_18625,N_14294,N_12285);
nor U18626 (N_18626,N_10121,N_12709);
and U18627 (N_18627,N_13942,N_13951);
nor U18628 (N_18628,N_12268,N_10401);
and U18629 (N_18629,N_12956,N_10755);
or U18630 (N_18630,N_12562,N_14596);
xnor U18631 (N_18631,N_12386,N_12385);
nand U18632 (N_18632,N_13556,N_10981);
nor U18633 (N_18633,N_12608,N_14478);
and U18634 (N_18634,N_11741,N_11798);
or U18635 (N_18635,N_13414,N_11546);
nor U18636 (N_18636,N_11859,N_12529);
nor U18637 (N_18637,N_13604,N_13542);
nor U18638 (N_18638,N_13311,N_13105);
or U18639 (N_18639,N_10041,N_14225);
nor U18640 (N_18640,N_12413,N_10509);
nand U18641 (N_18641,N_12215,N_12893);
nand U18642 (N_18642,N_12993,N_10878);
xor U18643 (N_18643,N_11725,N_13706);
or U18644 (N_18644,N_12622,N_10280);
nand U18645 (N_18645,N_11951,N_10000);
nand U18646 (N_18646,N_10079,N_11289);
or U18647 (N_18647,N_10857,N_13686);
and U18648 (N_18648,N_13803,N_10447);
nor U18649 (N_18649,N_14422,N_13448);
or U18650 (N_18650,N_13137,N_12706);
nand U18651 (N_18651,N_12786,N_10019);
nand U18652 (N_18652,N_13828,N_11609);
or U18653 (N_18653,N_12131,N_11753);
or U18654 (N_18654,N_10990,N_13582);
or U18655 (N_18655,N_12166,N_11409);
nand U18656 (N_18656,N_10723,N_13836);
or U18657 (N_18657,N_13484,N_10248);
xor U18658 (N_18658,N_13713,N_13332);
nand U18659 (N_18659,N_13090,N_13360);
and U18660 (N_18660,N_10918,N_14628);
nor U18661 (N_18661,N_11512,N_13655);
xnor U18662 (N_18662,N_12921,N_10124);
or U18663 (N_18663,N_14255,N_11539);
and U18664 (N_18664,N_13666,N_12453);
and U18665 (N_18665,N_10865,N_11295);
nand U18666 (N_18666,N_13790,N_13850);
and U18667 (N_18667,N_13056,N_11693);
nand U18668 (N_18668,N_11183,N_13779);
nor U18669 (N_18669,N_10508,N_12410);
and U18670 (N_18670,N_14471,N_12496);
nor U18671 (N_18671,N_13372,N_12838);
xor U18672 (N_18672,N_13592,N_13417);
or U18673 (N_18673,N_11789,N_11916);
and U18674 (N_18674,N_12077,N_12155);
xnor U18675 (N_18675,N_13802,N_10915);
and U18676 (N_18676,N_14915,N_14544);
nor U18677 (N_18677,N_10599,N_13988);
nand U18678 (N_18678,N_12897,N_11283);
xnor U18679 (N_18679,N_14260,N_11773);
nand U18680 (N_18680,N_13692,N_12689);
and U18681 (N_18681,N_10398,N_14506);
nor U18682 (N_18682,N_12614,N_12612);
nand U18683 (N_18683,N_10014,N_10209);
nor U18684 (N_18684,N_13788,N_12870);
and U18685 (N_18685,N_11949,N_11946);
nand U18686 (N_18686,N_12658,N_12628);
nor U18687 (N_18687,N_11527,N_14740);
nor U18688 (N_18688,N_12490,N_13915);
nor U18689 (N_18689,N_11866,N_13086);
nand U18690 (N_18690,N_10537,N_10899);
xor U18691 (N_18691,N_11975,N_13529);
and U18692 (N_18692,N_13462,N_12723);
and U18693 (N_18693,N_14901,N_11670);
nor U18694 (N_18694,N_13626,N_13933);
or U18695 (N_18695,N_12233,N_11753);
nor U18696 (N_18696,N_10428,N_10453);
nand U18697 (N_18697,N_11055,N_10497);
nor U18698 (N_18698,N_10797,N_11945);
nor U18699 (N_18699,N_11068,N_14378);
nand U18700 (N_18700,N_14796,N_13752);
or U18701 (N_18701,N_11498,N_11719);
and U18702 (N_18702,N_13764,N_13236);
or U18703 (N_18703,N_10000,N_12061);
xor U18704 (N_18704,N_11341,N_11177);
and U18705 (N_18705,N_14239,N_14754);
nor U18706 (N_18706,N_14565,N_14132);
nor U18707 (N_18707,N_14709,N_11539);
or U18708 (N_18708,N_13122,N_14266);
nor U18709 (N_18709,N_12552,N_12137);
nand U18710 (N_18710,N_11620,N_12237);
nand U18711 (N_18711,N_14897,N_13375);
xor U18712 (N_18712,N_13360,N_12090);
or U18713 (N_18713,N_12748,N_13752);
nor U18714 (N_18714,N_13836,N_14870);
xnor U18715 (N_18715,N_10867,N_12038);
and U18716 (N_18716,N_10579,N_11636);
nand U18717 (N_18717,N_14606,N_12604);
nand U18718 (N_18718,N_12699,N_10359);
and U18719 (N_18719,N_10843,N_13477);
xor U18720 (N_18720,N_12344,N_12491);
or U18721 (N_18721,N_11869,N_11210);
nor U18722 (N_18722,N_10171,N_10138);
and U18723 (N_18723,N_12671,N_13607);
or U18724 (N_18724,N_14629,N_14610);
and U18725 (N_18725,N_14330,N_11814);
and U18726 (N_18726,N_11345,N_11868);
nand U18727 (N_18727,N_10405,N_13423);
and U18728 (N_18728,N_12254,N_11073);
nand U18729 (N_18729,N_10930,N_13133);
nand U18730 (N_18730,N_10982,N_10924);
nor U18731 (N_18731,N_10916,N_13478);
and U18732 (N_18732,N_13402,N_14763);
nand U18733 (N_18733,N_10265,N_11593);
and U18734 (N_18734,N_12841,N_10088);
nor U18735 (N_18735,N_10210,N_12635);
xor U18736 (N_18736,N_13358,N_11520);
and U18737 (N_18737,N_13718,N_11292);
nor U18738 (N_18738,N_12003,N_12740);
or U18739 (N_18739,N_11526,N_12896);
nor U18740 (N_18740,N_11781,N_11143);
nand U18741 (N_18741,N_12173,N_11077);
nand U18742 (N_18742,N_13283,N_10710);
and U18743 (N_18743,N_11463,N_11532);
and U18744 (N_18744,N_14603,N_11514);
nand U18745 (N_18745,N_12438,N_12471);
nand U18746 (N_18746,N_10918,N_14925);
or U18747 (N_18747,N_11746,N_10697);
and U18748 (N_18748,N_13597,N_10570);
or U18749 (N_18749,N_13554,N_13472);
nand U18750 (N_18750,N_13271,N_14865);
nand U18751 (N_18751,N_13167,N_13481);
or U18752 (N_18752,N_10863,N_11288);
and U18753 (N_18753,N_12589,N_13903);
and U18754 (N_18754,N_11629,N_10473);
nand U18755 (N_18755,N_11497,N_12685);
and U18756 (N_18756,N_10963,N_13771);
nor U18757 (N_18757,N_10374,N_13195);
nand U18758 (N_18758,N_14796,N_10233);
xor U18759 (N_18759,N_12784,N_13532);
xnor U18760 (N_18760,N_13110,N_13005);
or U18761 (N_18761,N_10984,N_14876);
nor U18762 (N_18762,N_11094,N_12034);
nand U18763 (N_18763,N_11128,N_12091);
and U18764 (N_18764,N_12400,N_13724);
nor U18765 (N_18765,N_13744,N_12477);
and U18766 (N_18766,N_12126,N_11406);
and U18767 (N_18767,N_11615,N_10357);
nor U18768 (N_18768,N_11704,N_12215);
nand U18769 (N_18769,N_12947,N_12032);
xor U18770 (N_18770,N_11131,N_12293);
or U18771 (N_18771,N_14555,N_11607);
nand U18772 (N_18772,N_14061,N_11280);
nand U18773 (N_18773,N_10763,N_10388);
nand U18774 (N_18774,N_10825,N_12960);
or U18775 (N_18775,N_11393,N_14628);
xnor U18776 (N_18776,N_11797,N_13230);
xnor U18777 (N_18777,N_10785,N_14153);
and U18778 (N_18778,N_12638,N_12487);
nand U18779 (N_18779,N_10034,N_10103);
and U18780 (N_18780,N_12170,N_13202);
or U18781 (N_18781,N_12657,N_14066);
nand U18782 (N_18782,N_12675,N_10371);
and U18783 (N_18783,N_14321,N_13647);
nor U18784 (N_18784,N_14506,N_10671);
xnor U18785 (N_18785,N_13752,N_12449);
nand U18786 (N_18786,N_11405,N_12109);
nand U18787 (N_18787,N_14339,N_12579);
nand U18788 (N_18788,N_13926,N_14797);
nor U18789 (N_18789,N_12029,N_10454);
nor U18790 (N_18790,N_11986,N_10743);
nand U18791 (N_18791,N_14962,N_11195);
and U18792 (N_18792,N_14994,N_14068);
nand U18793 (N_18793,N_12937,N_13798);
nand U18794 (N_18794,N_11704,N_10075);
and U18795 (N_18795,N_10782,N_11920);
nand U18796 (N_18796,N_11812,N_12787);
and U18797 (N_18797,N_10362,N_12863);
nand U18798 (N_18798,N_13502,N_13739);
nor U18799 (N_18799,N_10952,N_11966);
and U18800 (N_18800,N_10660,N_13479);
nand U18801 (N_18801,N_12751,N_12556);
nor U18802 (N_18802,N_11883,N_13078);
nand U18803 (N_18803,N_11725,N_11602);
nor U18804 (N_18804,N_11876,N_10457);
and U18805 (N_18805,N_13527,N_13520);
and U18806 (N_18806,N_11778,N_14009);
or U18807 (N_18807,N_14331,N_10403);
xnor U18808 (N_18808,N_11324,N_11311);
or U18809 (N_18809,N_13173,N_12926);
or U18810 (N_18810,N_12285,N_14123);
or U18811 (N_18811,N_13002,N_13182);
nand U18812 (N_18812,N_11786,N_11843);
or U18813 (N_18813,N_11555,N_14965);
nand U18814 (N_18814,N_12966,N_13409);
nand U18815 (N_18815,N_14178,N_10861);
nand U18816 (N_18816,N_12196,N_12245);
and U18817 (N_18817,N_11702,N_14041);
and U18818 (N_18818,N_13719,N_10582);
or U18819 (N_18819,N_11649,N_10404);
xnor U18820 (N_18820,N_12581,N_10190);
nand U18821 (N_18821,N_13509,N_13503);
nor U18822 (N_18822,N_11124,N_13283);
or U18823 (N_18823,N_12912,N_11150);
nand U18824 (N_18824,N_12864,N_11192);
nand U18825 (N_18825,N_12288,N_11639);
nor U18826 (N_18826,N_10312,N_13376);
or U18827 (N_18827,N_11509,N_13841);
or U18828 (N_18828,N_13956,N_11377);
nand U18829 (N_18829,N_11366,N_10987);
or U18830 (N_18830,N_12851,N_10122);
or U18831 (N_18831,N_13138,N_10701);
and U18832 (N_18832,N_10725,N_10506);
or U18833 (N_18833,N_11933,N_13715);
nand U18834 (N_18834,N_11833,N_13515);
and U18835 (N_18835,N_11346,N_12294);
nand U18836 (N_18836,N_14701,N_13282);
and U18837 (N_18837,N_13170,N_12138);
and U18838 (N_18838,N_11829,N_13035);
and U18839 (N_18839,N_12278,N_10035);
xor U18840 (N_18840,N_11502,N_11948);
xor U18841 (N_18841,N_11754,N_14061);
and U18842 (N_18842,N_11373,N_12863);
or U18843 (N_18843,N_12954,N_11525);
or U18844 (N_18844,N_13595,N_10391);
nor U18845 (N_18845,N_11949,N_12203);
or U18846 (N_18846,N_14447,N_10209);
nand U18847 (N_18847,N_13564,N_11409);
nand U18848 (N_18848,N_10873,N_13664);
xor U18849 (N_18849,N_11736,N_13037);
or U18850 (N_18850,N_12053,N_10437);
nor U18851 (N_18851,N_10971,N_12597);
nand U18852 (N_18852,N_10866,N_14661);
xnor U18853 (N_18853,N_11381,N_12800);
and U18854 (N_18854,N_11694,N_12260);
nand U18855 (N_18855,N_11961,N_14218);
nor U18856 (N_18856,N_12255,N_13715);
nand U18857 (N_18857,N_10810,N_12871);
or U18858 (N_18858,N_12567,N_14329);
and U18859 (N_18859,N_14935,N_12344);
xor U18860 (N_18860,N_12130,N_13797);
nand U18861 (N_18861,N_14174,N_13668);
or U18862 (N_18862,N_12575,N_14267);
nor U18863 (N_18863,N_12713,N_11156);
xor U18864 (N_18864,N_10914,N_14265);
xnor U18865 (N_18865,N_12434,N_12200);
nor U18866 (N_18866,N_12701,N_10857);
or U18867 (N_18867,N_11630,N_12288);
nor U18868 (N_18868,N_14305,N_14104);
nor U18869 (N_18869,N_14034,N_13971);
or U18870 (N_18870,N_10679,N_11652);
nand U18871 (N_18871,N_14424,N_14594);
nand U18872 (N_18872,N_13409,N_11209);
and U18873 (N_18873,N_12206,N_12027);
nand U18874 (N_18874,N_14786,N_14109);
nand U18875 (N_18875,N_12023,N_13245);
or U18876 (N_18876,N_11784,N_10658);
nand U18877 (N_18877,N_10518,N_10168);
nand U18878 (N_18878,N_13063,N_10468);
or U18879 (N_18879,N_11554,N_13703);
xnor U18880 (N_18880,N_12134,N_11602);
and U18881 (N_18881,N_11393,N_10913);
xnor U18882 (N_18882,N_14185,N_13215);
nor U18883 (N_18883,N_14942,N_13930);
nand U18884 (N_18884,N_13005,N_13809);
and U18885 (N_18885,N_14036,N_13997);
and U18886 (N_18886,N_12717,N_13371);
and U18887 (N_18887,N_14496,N_12965);
and U18888 (N_18888,N_14754,N_11164);
and U18889 (N_18889,N_10864,N_10882);
nor U18890 (N_18890,N_13509,N_14722);
nor U18891 (N_18891,N_11732,N_13889);
nor U18892 (N_18892,N_10593,N_10952);
nor U18893 (N_18893,N_12124,N_12341);
or U18894 (N_18894,N_12200,N_14057);
and U18895 (N_18895,N_12488,N_11070);
and U18896 (N_18896,N_13211,N_11978);
or U18897 (N_18897,N_10514,N_13308);
or U18898 (N_18898,N_13767,N_11024);
nand U18899 (N_18899,N_12145,N_10856);
nor U18900 (N_18900,N_11962,N_12875);
xnor U18901 (N_18901,N_10153,N_13526);
nand U18902 (N_18902,N_14772,N_14163);
or U18903 (N_18903,N_13833,N_12123);
nand U18904 (N_18904,N_10157,N_10226);
and U18905 (N_18905,N_14278,N_11221);
and U18906 (N_18906,N_13209,N_13707);
and U18907 (N_18907,N_11759,N_11091);
or U18908 (N_18908,N_10467,N_13089);
and U18909 (N_18909,N_11962,N_13068);
nand U18910 (N_18910,N_12378,N_13938);
and U18911 (N_18911,N_12440,N_12133);
or U18912 (N_18912,N_12477,N_13496);
xnor U18913 (N_18913,N_12421,N_10331);
or U18914 (N_18914,N_13452,N_12246);
and U18915 (N_18915,N_14484,N_13037);
or U18916 (N_18916,N_14579,N_12758);
and U18917 (N_18917,N_13907,N_10442);
and U18918 (N_18918,N_14568,N_10656);
and U18919 (N_18919,N_14122,N_12670);
or U18920 (N_18920,N_13316,N_12706);
or U18921 (N_18921,N_11665,N_11599);
nor U18922 (N_18922,N_10368,N_10431);
and U18923 (N_18923,N_14435,N_13724);
or U18924 (N_18924,N_13105,N_11364);
and U18925 (N_18925,N_12025,N_14903);
or U18926 (N_18926,N_11795,N_10708);
and U18927 (N_18927,N_13420,N_10026);
and U18928 (N_18928,N_11408,N_10840);
nor U18929 (N_18929,N_14698,N_10652);
and U18930 (N_18930,N_10349,N_12188);
nor U18931 (N_18931,N_11713,N_12862);
and U18932 (N_18932,N_12758,N_14590);
nor U18933 (N_18933,N_12482,N_14462);
or U18934 (N_18934,N_13924,N_14858);
xor U18935 (N_18935,N_12073,N_10118);
nor U18936 (N_18936,N_11406,N_12841);
and U18937 (N_18937,N_12857,N_14748);
nand U18938 (N_18938,N_13967,N_11596);
or U18939 (N_18939,N_10224,N_11676);
nor U18940 (N_18940,N_10364,N_13423);
xnor U18941 (N_18941,N_14423,N_10485);
nand U18942 (N_18942,N_13057,N_13646);
and U18943 (N_18943,N_10742,N_11090);
nor U18944 (N_18944,N_10538,N_10749);
and U18945 (N_18945,N_10904,N_14547);
or U18946 (N_18946,N_13097,N_12722);
nand U18947 (N_18947,N_13258,N_11386);
xor U18948 (N_18948,N_11781,N_10744);
or U18949 (N_18949,N_11747,N_11776);
nor U18950 (N_18950,N_10884,N_10136);
or U18951 (N_18951,N_14982,N_12784);
or U18952 (N_18952,N_14511,N_11059);
nand U18953 (N_18953,N_14182,N_13858);
nand U18954 (N_18954,N_10879,N_10691);
nor U18955 (N_18955,N_10724,N_14932);
nand U18956 (N_18956,N_12133,N_13189);
and U18957 (N_18957,N_12678,N_12600);
or U18958 (N_18958,N_10039,N_11502);
nor U18959 (N_18959,N_11904,N_13090);
nand U18960 (N_18960,N_14319,N_13928);
or U18961 (N_18961,N_10645,N_10736);
xnor U18962 (N_18962,N_13749,N_14498);
or U18963 (N_18963,N_13027,N_14081);
nand U18964 (N_18964,N_12876,N_12135);
nand U18965 (N_18965,N_11872,N_12085);
nand U18966 (N_18966,N_14724,N_10325);
or U18967 (N_18967,N_11374,N_10821);
nor U18968 (N_18968,N_14670,N_13359);
and U18969 (N_18969,N_10641,N_14092);
xor U18970 (N_18970,N_13439,N_11997);
and U18971 (N_18971,N_13947,N_12659);
nand U18972 (N_18972,N_12677,N_12629);
or U18973 (N_18973,N_11071,N_13336);
nand U18974 (N_18974,N_10524,N_12043);
or U18975 (N_18975,N_10527,N_11592);
nand U18976 (N_18976,N_12040,N_13855);
nor U18977 (N_18977,N_11936,N_13795);
xor U18978 (N_18978,N_13245,N_13132);
nor U18979 (N_18979,N_13048,N_12655);
or U18980 (N_18980,N_11556,N_10231);
nand U18981 (N_18981,N_10004,N_12516);
nand U18982 (N_18982,N_12816,N_10573);
or U18983 (N_18983,N_12431,N_12236);
or U18984 (N_18984,N_14921,N_14274);
xnor U18985 (N_18985,N_12436,N_10273);
and U18986 (N_18986,N_10895,N_11116);
nor U18987 (N_18987,N_11312,N_13867);
and U18988 (N_18988,N_10467,N_12951);
or U18989 (N_18989,N_10134,N_12392);
nand U18990 (N_18990,N_10112,N_10784);
and U18991 (N_18991,N_13871,N_10220);
and U18992 (N_18992,N_12983,N_12651);
nand U18993 (N_18993,N_12044,N_12181);
nor U18994 (N_18994,N_10108,N_14861);
or U18995 (N_18995,N_13946,N_13417);
nor U18996 (N_18996,N_12972,N_10251);
nand U18997 (N_18997,N_11893,N_14113);
nand U18998 (N_18998,N_13554,N_10589);
xor U18999 (N_18999,N_11280,N_13704);
or U19000 (N_19000,N_11920,N_10589);
nor U19001 (N_19001,N_11581,N_12880);
nor U19002 (N_19002,N_10466,N_13488);
xor U19003 (N_19003,N_11277,N_10501);
nor U19004 (N_19004,N_12809,N_14178);
and U19005 (N_19005,N_10533,N_12365);
and U19006 (N_19006,N_14575,N_14960);
nand U19007 (N_19007,N_12460,N_10283);
nand U19008 (N_19008,N_13117,N_11415);
nand U19009 (N_19009,N_10942,N_13512);
or U19010 (N_19010,N_12809,N_13962);
or U19011 (N_19011,N_14616,N_11512);
and U19012 (N_19012,N_13613,N_11828);
xnor U19013 (N_19013,N_10993,N_13761);
nand U19014 (N_19014,N_11340,N_12185);
nand U19015 (N_19015,N_10539,N_12694);
or U19016 (N_19016,N_13628,N_12660);
nand U19017 (N_19017,N_10244,N_10564);
nand U19018 (N_19018,N_11260,N_11199);
xnor U19019 (N_19019,N_10461,N_10966);
nor U19020 (N_19020,N_13797,N_12022);
or U19021 (N_19021,N_11011,N_12722);
xor U19022 (N_19022,N_14733,N_13409);
and U19023 (N_19023,N_13376,N_11011);
and U19024 (N_19024,N_14294,N_10674);
nor U19025 (N_19025,N_13340,N_13377);
nand U19026 (N_19026,N_13470,N_12254);
and U19027 (N_19027,N_14820,N_12681);
or U19028 (N_19028,N_12757,N_14891);
or U19029 (N_19029,N_12516,N_12179);
nor U19030 (N_19030,N_11348,N_11764);
and U19031 (N_19031,N_14228,N_12809);
and U19032 (N_19032,N_12533,N_10756);
and U19033 (N_19033,N_11269,N_12286);
and U19034 (N_19034,N_13905,N_11568);
nor U19035 (N_19035,N_12289,N_10320);
xnor U19036 (N_19036,N_14279,N_10208);
or U19037 (N_19037,N_13513,N_12354);
or U19038 (N_19038,N_13645,N_14614);
or U19039 (N_19039,N_10553,N_10049);
nand U19040 (N_19040,N_11364,N_11705);
or U19041 (N_19041,N_13053,N_13086);
or U19042 (N_19042,N_10218,N_11271);
nand U19043 (N_19043,N_11056,N_13621);
or U19044 (N_19044,N_12182,N_12147);
or U19045 (N_19045,N_10330,N_12379);
nor U19046 (N_19046,N_12764,N_13587);
nor U19047 (N_19047,N_11703,N_11545);
or U19048 (N_19048,N_13710,N_11355);
nand U19049 (N_19049,N_12304,N_12743);
nor U19050 (N_19050,N_13004,N_10509);
nand U19051 (N_19051,N_10206,N_11336);
nor U19052 (N_19052,N_14335,N_13235);
nand U19053 (N_19053,N_14117,N_12486);
or U19054 (N_19054,N_14252,N_12516);
and U19055 (N_19055,N_10590,N_11656);
nand U19056 (N_19056,N_13947,N_10046);
nand U19057 (N_19057,N_12748,N_14671);
xnor U19058 (N_19058,N_14061,N_12482);
nor U19059 (N_19059,N_11676,N_11811);
and U19060 (N_19060,N_11471,N_12782);
or U19061 (N_19061,N_12541,N_11793);
or U19062 (N_19062,N_14131,N_13502);
xor U19063 (N_19063,N_10003,N_11237);
or U19064 (N_19064,N_14595,N_11534);
nand U19065 (N_19065,N_12612,N_11612);
and U19066 (N_19066,N_14609,N_10672);
nor U19067 (N_19067,N_11555,N_11536);
xnor U19068 (N_19068,N_10078,N_13047);
xor U19069 (N_19069,N_12716,N_12343);
or U19070 (N_19070,N_11845,N_11352);
or U19071 (N_19071,N_10016,N_12532);
nand U19072 (N_19072,N_12120,N_11731);
or U19073 (N_19073,N_11214,N_10192);
nor U19074 (N_19074,N_14795,N_14539);
nand U19075 (N_19075,N_13858,N_10948);
or U19076 (N_19076,N_12321,N_13307);
and U19077 (N_19077,N_11823,N_11320);
nand U19078 (N_19078,N_11304,N_12884);
nor U19079 (N_19079,N_10334,N_10829);
xnor U19080 (N_19080,N_11337,N_14937);
nand U19081 (N_19081,N_14010,N_11195);
nor U19082 (N_19082,N_11908,N_10010);
nand U19083 (N_19083,N_11316,N_13460);
nor U19084 (N_19084,N_10858,N_14161);
or U19085 (N_19085,N_13906,N_10714);
or U19086 (N_19086,N_14952,N_12864);
nor U19087 (N_19087,N_14459,N_13231);
and U19088 (N_19088,N_13142,N_12962);
or U19089 (N_19089,N_11314,N_13881);
nand U19090 (N_19090,N_14110,N_13765);
or U19091 (N_19091,N_11030,N_12472);
nor U19092 (N_19092,N_14589,N_14243);
and U19093 (N_19093,N_10546,N_12017);
nand U19094 (N_19094,N_14277,N_11867);
or U19095 (N_19095,N_14674,N_14180);
xor U19096 (N_19096,N_14864,N_14059);
and U19097 (N_19097,N_10483,N_10285);
and U19098 (N_19098,N_13745,N_14297);
nor U19099 (N_19099,N_12219,N_14879);
or U19100 (N_19100,N_12169,N_14792);
nor U19101 (N_19101,N_11290,N_10250);
or U19102 (N_19102,N_13639,N_13481);
or U19103 (N_19103,N_10707,N_14165);
xnor U19104 (N_19104,N_12988,N_12400);
nand U19105 (N_19105,N_12369,N_13955);
or U19106 (N_19106,N_10987,N_11541);
or U19107 (N_19107,N_14424,N_12392);
nor U19108 (N_19108,N_12139,N_10040);
nand U19109 (N_19109,N_14453,N_12273);
xnor U19110 (N_19110,N_11231,N_13344);
xnor U19111 (N_19111,N_12530,N_13602);
nand U19112 (N_19112,N_11626,N_10038);
and U19113 (N_19113,N_10062,N_10544);
nand U19114 (N_19114,N_11734,N_12609);
and U19115 (N_19115,N_13618,N_13027);
nand U19116 (N_19116,N_12293,N_12151);
nor U19117 (N_19117,N_10850,N_13410);
nor U19118 (N_19118,N_11698,N_10802);
nor U19119 (N_19119,N_14946,N_13689);
nor U19120 (N_19120,N_13351,N_14233);
nor U19121 (N_19121,N_14448,N_10065);
nand U19122 (N_19122,N_10020,N_11309);
xor U19123 (N_19123,N_13750,N_14869);
or U19124 (N_19124,N_11475,N_10994);
nand U19125 (N_19125,N_12893,N_14190);
nor U19126 (N_19126,N_10446,N_14382);
nor U19127 (N_19127,N_13032,N_10608);
nand U19128 (N_19128,N_13214,N_10980);
nand U19129 (N_19129,N_13805,N_14209);
nor U19130 (N_19130,N_14015,N_10465);
and U19131 (N_19131,N_12936,N_12238);
nor U19132 (N_19132,N_14986,N_13292);
or U19133 (N_19133,N_13312,N_13648);
or U19134 (N_19134,N_13013,N_14302);
and U19135 (N_19135,N_14000,N_13028);
nand U19136 (N_19136,N_13105,N_14706);
xnor U19137 (N_19137,N_12772,N_14672);
and U19138 (N_19138,N_11962,N_14675);
nand U19139 (N_19139,N_11289,N_10781);
or U19140 (N_19140,N_11049,N_14620);
nand U19141 (N_19141,N_10942,N_13534);
nand U19142 (N_19142,N_14255,N_12253);
xnor U19143 (N_19143,N_11182,N_12866);
or U19144 (N_19144,N_14643,N_14528);
and U19145 (N_19145,N_11414,N_14878);
or U19146 (N_19146,N_11992,N_12306);
nor U19147 (N_19147,N_11619,N_11949);
nand U19148 (N_19148,N_11780,N_11329);
nand U19149 (N_19149,N_10571,N_10654);
nand U19150 (N_19150,N_13345,N_14844);
and U19151 (N_19151,N_12902,N_12730);
and U19152 (N_19152,N_12842,N_12811);
and U19153 (N_19153,N_13625,N_13667);
or U19154 (N_19154,N_11284,N_11937);
nand U19155 (N_19155,N_10198,N_11572);
and U19156 (N_19156,N_13199,N_10952);
xor U19157 (N_19157,N_14687,N_14536);
nand U19158 (N_19158,N_11281,N_13089);
and U19159 (N_19159,N_13959,N_14926);
and U19160 (N_19160,N_13016,N_13812);
nand U19161 (N_19161,N_10888,N_12164);
nand U19162 (N_19162,N_14497,N_10747);
or U19163 (N_19163,N_11600,N_10177);
nor U19164 (N_19164,N_13416,N_14897);
nand U19165 (N_19165,N_13524,N_11447);
nand U19166 (N_19166,N_14219,N_11281);
nand U19167 (N_19167,N_10804,N_13382);
or U19168 (N_19168,N_12704,N_14688);
xnor U19169 (N_19169,N_13620,N_12104);
nand U19170 (N_19170,N_13802,N_10014);
and U19171 (N_19171,N_13175,N_10754);
and U19172 (N_19172,N_10082,N_12081);
xor U19173 (N_19173,N_12445,N_10885);
nor U19174 (N_19174,N_14821,N_14744);
and U19175 (N_19175,N_13600,N_13934);
nand U19176 (N_19176,N_13594,N_14458);
nor U19177 (N_19177,N_10918,N_12819);
nand U19178 (N_19178,N_11351,N_11200);
nand U19179 (N_19179,N_14097,N_12193);
nand U19180 (N_19180,N_13255,N_13906);
xnor U19181 (N_19181,N_14216,N_12061);
and U19182 (N_19182,N_12099,N_13456);
xnor U19183 (N_19183,N_14153,N_12709);
and U19184 (N_19184,N_11635,N_11614);
nor U19185 (N_19185,N_10744,N_12105);
nand U19186 (N_19186,N_13426,N_10072);
and U19187 (N_19187,N_13294,N_11491);
xor U19188 (N_19188,N_10698,N_11525);
and U19189 (N_19189,N_14445,N_12229);
nor U19190 (N_19190,N_10388,N_11251);
nor U19191 (N_19191,N_13947,N_10886);
or U19192 (N_19192,N_11139,N_13650);
xnor U19193 (N_19193,N_11615,N_10944);
and U19194 (N_19194,N_11301,N_12306);
nor U19195 (N_19195,N_10218,N_14750);
nor U19196 (N_19196,N_12317,N_10241);
and U19197 (N_19197,N_10016,N_14485);
and U19198 (N_19198,N_12166,N_14923);
and U19199 (N_19199,N_12869,N_10716);
or U19200 (N_19200,N_13280,N_11413);
or U19201 (N_19201,N_10285,N_10813);
nand U19202 (N_19202,N_12359,N_12477);
nand U19203 (N_19203,N_13767,N_10001);
nor U19204 (N_19204,N_10801,N_12061);
or U19205 (N_19205,N_13808,N_13585);
or U19206 (N_19206,N_12837,N_13330);
or U19207 (N_19207,N_11107,N_12346);
nor U19208 (N_19208,N_12152,N_13031);
xnor U19209 (N_19209,N_11271,N_11516);
nor U19210 (N_19210,N_10947,N_10176);
and U19211 (N_19211,N_12304,N_11805);
or U19212 (N_19212,N_11524,N_14170);
nand U19213 (N_19213,N_11947,N_13153);
and U19214 (N_19214,N_10772,N_14269);
nand U19215 (N_19215,N_10941,N_13230);
or U19216 (N_19216,N_10639,N_12824);
and U19217 (N_19217,N_13504,N_11924);
or U19218 (N_19218,N_13092,N_14144);
nand U19219 (N_19219,N_12952,N_13724);
nand U19220 (N_19220,N_12775,N_14198);
and U19221 (N_19221,N_10236,N_12508);
nand U19222 (N_19222,N_12437,N_14779);
nand U19223 (N_19223,N_13964,N_11437);
nand U19224 (N_19224,N_12582,N_10784);
and U19225 (N_19225,N_12123,N_11504);
nand U19226 (N_19226,N_10587,N_14572);
nand U19227 (N_19227,N_12854,N_14836);
nor U19228 (N_19228,N_14728,N_13011);
nor U19229 (N_19229,N_14725,N_14301);
nor U19230 (N_19230,N_12518,N_12851);
nand U19231 (N_19231,N_13884,N_13691);
nor U19232 (N_19232,N_13625,N_14718);
and U19233 (N_19233,N_13733,N_14441);
and U19234 (N_19234,N_10058,N_11902);
nand U19235 (N_19235,N_13946,N_11110);
nand U19236 (N_19236,N_10187,N_14668);
and U19237 (N_19237,N_11463,N_10321);
xnor U19238 (N_19238,N_10324,N_12468);
nor U19239 (N_19239,N_12648,N_14329);
or U19240 (N_19240,N_14455,N_13862);
or U19241 (N_19241,N_13169,N_10391);
or U19242 (N_19242,N_11956,N_10434);
nor U19243 (N_19243,N_12248,N_11396);
nor U19244 (N_19244,N_10100,N_10499);
or U19245 (N_19245,N_12614,N_14698);
nor U19246 (N_19246,N_13851,N_13025);
nor U19247 (N_19247,N_10198,N_14348);
or U19248 (N_19248,N_11210,N_14804);
xnor U19249 (N_19249,N_11079,N_10547);
and U19250 (N_19250,N_14210,N_12581);
and U19251 (N_19251,N_10347,N_12754);
nor U19252 (N_19252,N_11323,N_10875);
or U19253 (N_19253,N_11893,N_12589);
and U19254 (N_19254,N_11076,N_13374);
or U19255 (N_19255,N_14323,N_12173);
or U19256 (N_19256,N_11093,N_12283);
and U19257 (N_19257,N_11839,N_10018);
xnor U19258 (N_19258,N_14201,N_13061);
xor U19259 (N_19259,N_12653,N_14483);
nor U19260 (N_19260,N_12923,N_11468);
and U19261 (N_19261,N_12467,N_13990);
and U19262 (N_19262,N_13543,N_10792);
and U19263 (N_19263,N_11556,N_14102);
and U19264 (N_19264,N_11082,N_12507);
nand U19265 (N_19265,N_11256,N_14804);
nand U19266 (N_19266,N_12163,N_14278);
and U19267 (N_19267,N_10706,N_10745);
nor U19268 (N_19268,N_11373,N_12218);
nand U19269 (N_19269,N_10491,N_11620);
or U19270 (N_19270,N_10444,N_11923);
or U19271 (N_19271,N_12272,N_12698);
nor U19272 (N_19272,N_11860,N_11500);
and U19273 (N_19273,N_12968,N_10034);
or U19274 (N_19274,N_10017,N_10123);
and U19275 (N_19275,N_12935,N_13226);
and U19276 (N_19276,N_13209,N_10245);
nor U19277 (N_19277,N_11753,N_14887);
nor U19278 (N_19278,N_11166,N_12929);
nor U19279 (N_19279,N_10077,N_11749);
xor U19280 (N_19280,N_11769,N_12561);
xor U19281 (N_19281,N_13806,N_12085);
nor U19282 (N_19282,N_12496,N_14072);
nand U19283 (N_19283,N_14810,N_14546);
nand U19284 (N_19284,N_13126,N_13927);
and U19285 (N_19285,N_10745,N_10569);
nand U19286 (N_19286,N_11653,N_14712);
or U19287 (N_19287,N_13055,N_14023);
or U19288 (N_19288,N_13223,N_10411);
xor U19289 (N_19289,N_14339,N_11810);
nand U19290 (N_19290,N_13074,N_10820);
nand U19291 (N_19291,N_10014,N_10714);
and U19292 (N_19292,N_14819,N_12763);
or U19293 (N_19293,N_11034,N_12660);
or U19294 (N_19294,N_11157,N_12082);
xnor U19295 (N_19295,N_11658,N_10732);
xnor U19296 (N_19296,N_11840,N_13344);
nand U19297 (N_19297,N_10735,N_14700);
or U19298 (N_19298,N_14513,N_10011);
and U19299 (N_19299,N_13393,N_11344);
nand U19300 (N_19300,N_12109,N_14210);
and U19301 (N_19301,N_13091,N_11738);
nand U19302 (N_19302,N_10224,N_14203);
and U19303 (N_19303,N_10013,N_11961);
nor U19304 (N_19304,N_10487,N_12058);
or U19305 (N_19305,N_12043,N_13028);
nor U19306 (N_19306,N_14059,N_13839);
xor U19307 (N_19307,N_12350,N_11788);
and U19308 (N_19308,N_10053,N_11996);
and U19309 (N_19309,N_12452,N_11553);
nor U19310 (N_19310,N_14736,N_14931);
and U19311 (N_19311,N_14782,N_12794);
nand U19312 (N_19312,N_13548,N_12843);
or U19313 (N_19313,N_12012,N_13748);
nand U19314 (N_19314,N_14699,N_13063);
nand U19315 (N_19315,N_10262,N_11645);
nand U19316 (N_19316,N_12874,N_14003);
and U19317 (N_19317,N_11281,N_11760);
and U19318 (N_19318,N_11081,N_11977);
nor U19319 (N_19319,N_10229,N_14552);
or U19320 (N_19320,N_11733,N_14472);
and U19321 (N_19321,N_12273,N_13950);
or U19322 (N_19322,N_14682,N_11089);
nand U19323 (N_19323,N_10744,N_12014);
and U19324 (N_19324,N_10986,N_13302);
nor U19325 (N_19325,N_12635,N_12857);
and U19326 (N_19326,N_10225,N_13854);
nand U19327 (N_19327,N_10793,N_14686);
nor U19328 (N_19328,N_14355,N_10382);
or U19329 (N_19329,N_14295,N_14575);
nor U19330 (N_19330,N_13026,N_12877);
or U19331 (N_19331,N_10045,N_14865);
and U19332 (N_19332,N_14522,N_12353);
nand U19333 (N_19333,N_14073,N_12309);
and U19334 (N_19334,N_10684,N_13237);
or U19335 (N_19335,N_12363,N_11780);
nor U19336 (N_19336,N_10494,N_10656);
nor U19337 (N_19337,N_11904,N_11779);
nor U19338 (N_19338,N_11556,N_12545);
and U19339 (N_19339,N_14091,N_13886);
nor U19340 (N_19340,N_13222,N_11280);
nor U19341 (N_19341,N_11761,N_14014);
and U19342 (N_19342,N_11306,N_10942);
nand U19343 (N_19343,N_10671,N_14803);
and U19344 (N_19344,N_12147,N_13819);
or U19345 (N_19345,N_13188,N_11699);
nand U19346 (N_19346,N_13127,N_12571);
nand U19347 (N_19347,N_10154,N_12168);
xnor U19348 (N_19348,N_11325,N_11264);
and U19349 (N_19349,N_10036,N_10069);
nor U19350 (N_19350,N_11705,N_12705);
nand U19351 (N_19351,N_12883,N_14826);
nand U19352 (N_19352,N_10660,N_12267);
and U19353 (N_19353,N_10537,N_11642);
xnor U19354 (N_19354,N_10481,N_10590);
or U19355 (N_19355,N_12482,N_12513);
and U19356 (N_19356,N_13523,N_10578);
nor U19357 (N_19357,N_12214,N_13332);
nor U19358 (N_19358,N_13435,N_12758);
or U19359 (N_19359,N_10099,N_12494);
or U19360 (N_19360,N_14626,N_14834);
and U19361 (N_19361,N_14533,N_14029);
nor U19362 (N_19362,N_13212,N_14520);
and U19363 (N_19363,N_10397,N_11977);
xor U19364 (N_19364,N_13701,N_12627);
nor U19365 (N_19365,N_10217,N_11716);
xor U19366 (N_19366,N_12516,N_12515);
nor U19367 (N_19367,N_13659,N_14570);
nand U19368 (N_19368,N_14808,N_10130);
nor U19369 (N_19369,N_11050,N_11915);
nand U19370 (N_19370,N_14683,N_11038);
nor U19371 (N_19371,N_12734,N_11687);
nor U19372 (N_19372,N_10029,N_13856);
and U19373 (N_19373,N_10740,N_13865);
nand U19374 (N_19374,N_14585,N_10856);
or U19375 (N_19375,N_13059,N_14147);
xor U19376 (N_19376,N_14008,N_12520);
or U19377 (N_19377,N_10600,N_10494);
nor U19378 (N_19378,N_14232,N_11710);
nand U19379 (N_19379,N_11516,N_10423);
nand U19380 (N_19380,N_13920,N_13501);
and U19381 (N_19381,N_10293,N_11811);
or U19382 (N_19382,N_14718,N_14171);
and U19383 (N_19383,N_13552,N_12543);
or U19384 (N_19384,N_14406,N_11781);
and U19385 (N_19385,N_14103,N_11621);
nand U19386 (N_19386,N_10315,N_10173);
nand U19387 (N_19387,N_13485,N_13896);
nor U19388 (N_19388,N_10664,N_10424);
nand U19389 (N_19389,N_13826,N_12159);
nand U19390 (N_19390,N_14710,N_13339);
nand U19391 (N_19391,N_10518,N_13581);
or U19392 (N_19392,N_10054,N_11504);
or U19393 (N_19393,N_10727,N_14201);
nand U19394 (N_19394,N_13133,N_14166);
xor U19395 (N_19395,N_12212,N_10016);
and U19396 (N_19396,N_12195,N_11208);
nand U19397 (N_19397,N_12017,N_12187);
and U19398 (N_19398,N_11875,N_12701);
and U19399 (N_19399,N_12435,N_13143);
or U19400 (N_19400,N_14889,N_11907);
nand U19401 (N_19401,N_12639,N_10088);
nor U19402 (N_19402,N_12333,N_12517);
or U19403 (N_19403,N_14334,N_13862);
nor U19404 (N_19404,N_11344,N_14026);
nor U19405 (N_19405,N_12169,N_11727);
or U19406 (N_19406,N_14514,N_12891);
nand U19407 (N_19407,N_11253,N_12539);
nor U19408 (N_19408,N_11878,N_13065);
and U19409 (N_19409,N_14543,N_10357);
and U19410 (N_19410,N_14698,N_12100);
nor U19411 (N_19411,N_13416,N_10224);
nor U19412 (N_19412,N_10549,N_14292);
and U19413 (N_19413,N_14528,N_14465);
or U19414 (N_19414,N_11255,N_12460);
xnor U19415 (N_19415,N_14764,N_14229);
nand U19416 (N_19416,N_11164,N_13308);
and U19417 (N_19417,N_10497,N_14280);
or U19418 (N_19418,N_10136,N_13456);
xor U19419 (N_19419,N_13974,N_13253);
and U19420 (N_19420,N_14765,N_14224);
and U19421 (N_19421,N_13108,N_12067);
or U19422 (N_19422,N_11582,N_11406);
and U19423 (N_19423,N_14916,N_11334);
or U19424 (N_19424,N_10280,N_12099);
nor U19425 (N_19425,N_10541,N_14390);
nor U19426 (N_19426,N_14626,N_13785);
nor U19427 (N_19427,N_11448,N_13400);
nor U19428 (N_19428,N_14939,N_12369);
nand U19429 (N_19429,N_13575,N_10938);
and U19430 (N_19430,N_10629,N_13533);
and U19431 (N_19431,N_11560,N_11576);
nor U19432 (N_19432,N_11252,N_12448);
nand U19433 (N_19433,N_12612,N_14604);
and U19434 (N_19434,N_11048,N_10184);
nor U19435 (N_19435,N_14469,N_14342);
xor U19436 (N_19436,N_10726,N_11341);
xor U19437 (N_19437,N_11134,N_14203);
and U19438 (N_19438,N_13587,N_13899);
and U19439 (N_19439,N_12895,N_10267);
nand U19440 (N_19440,N_13599,N_13016);
and U19441 (N_19441,N_13519,N_13254);
xnor U19442 (N_19442,N_11938,N_11156);
and U19443 (N_19443,N_14470,N_10827);
nand U19444 (N_19444,N_11025,N_12142);
nand U19445 (N_19445,N_14334,N_14570);
and U19446 (N_19446,N_12878,N_10378);
xor U19447 (N_19447,N_10762,N_11113);
nor U19448 (N_19448,N_13734,N_13736);
and U19449 (N_19449,N_11584,N_14915);
nor U19450 (N_19450,N_10631,N_11088);
or U19451 (N_19451,N_14903,N_14988);
nor U19452 (N_19452,N_13191,N_12539);
nor U19453 (N_19453,N_10370,N_10915);
or U19454 (N_19454,N_13510,N_14997);
or U19455 (N_19455,N_14772,N_13899);
nand U19456 (N_19456,N_12230,N_12451);
xnor U19457 (N_19457,N_12181,N_11278);
nand U19458 (N_19458,N_12867,N_11659);
and U19459 (N_19459,N_10604,N_10980);
nand U19460 (N_19460,N_14254,N_11823);
and U19461 (N_19461,N_11685,N_13779);
nand U19462 (N_19462,N_11820,N_11843);
and U19463 (N_19463,N_11625,N_11285);
xor U19464 (N_19464,N_11574,N_12300);
nor U19465 (N_19465,N_14049,N_14861);
nor U19466 (N_19466,N_14867,N_12306);
nor U19467 (N_19467,N_12259,N_11945);
nand U19468 (N_19468,N_12254,N_11021);
nand U19469 (N_19469,N_10757,N_11374);
or U19470 (N_19470,N_11857,N_10314);
nor U19471 (N_19471,N_12848,N_12509);
nand U19472 (N_19472,N_13098,N_12000);
nor U19473 (N_19473,N_13055,N_14449);
and U19474 (N_19474,N_14324,N_10396);
nand U19475 (N_19475,N_12934,N_11817);
nand U19476 (N_19476,N_13916,N_12401);
or U19477 (N_19477,N_11903,N_13091);
or U19478 (N_19478,N_11282,N_12768);
nor U19479 (N_19479,N_11593,N_11115);
or U19480 (N_19480,N_14899,N_13252);
nand U19481 (N_19481,N_12379,N_11640);
and U19482 (N_19482,N_13958,N_11664);
or U19483 (N_19483,N_10059,N_13945);
and U19484 (N_19484,N_12543,N_11538);
nand U19485 (N_19485,N_14905,N_13676);
nor U19486 (N_19486,N_12626,N_13222);
nand U19487 (N_19487,N_12076,N_14057);
and U19488 (N_19488,N_14160,N_12651);
nand U19489 (N_19489,N_11179,N_13349);
xor U19490 (N_19490,N_13101,N_14197);
nand U19491 (N_19491,N_10661,N_10941);
nor U19492 (N_19492,N_13654,N_14934);
nor U19493 (N_19493,N_13125,N_14982);
and U19494 (N_19494,N_10067,N_13396);
nor U19495 (N_19495,N_13994,N_13268);
xor U19496 (N_19496,N_10456,N_13208);
nor U19497 (N_19497,N_10972,N_10689);
and U19498 (N_19498,N_10873,N_14349);
or U19499 (N_19499,N_14780,N_14086);
nor U19500 (N_19500,N_10959,N_12701);
and U19501 (N_19501,N_13951,N_11677);
nor U19502 (N_19502,N_14573,N_11493);
nor U19503 (N_19503,N_11246,N_14608);
nand U19504 (N_19504,N_13646,N_14838);
and U19505 (N_19505,N_13996,N_11103);
nor U19506 (N_19506,N_14587,N_10166);
nor U19507 (N_19507,N_13447,N_11053);
or U19508 (N_19508,N_12398,N_10199);
and U19509 (N_19509,N_12726,N_11160);
or U19510 (N_19510,N_14814,N_12489);
nand U19511 (N_19511,N_11898,N_11121);
or U19512 (N_19512,N_11044,N_10439);
xor U19513 (N_19513,N_14390,N_14368);
and U19514 (N_19514,N_13573,N_10365);
nand U19515 (N_19515,N_14574,N_10664);
or U19516 (N_19516,N_13033,N_10163);
or U19517 (N_19517,N_11558,N_12031);
or U19518 (N_19518,N_13523,N_13197);
xor U19519 (N_19519,N_10862,N_14929);
nand U19520 (N_19520,N_14250,N_10721);
nor U19521 (N_19521,N_10279,N_13656);
or U19522 (N_19522,N_10473,N_14326);
xnor U19523 (N_19523,N_11733,N_11525);
nor U19524 (N_19524,N_13758,N_11926);
and U19525 (N_19525,N_12134,N_12001);
nand U19526 (N_19526,N_10448,N_12565);
nor U19527 (N_19527,N_14066,N_10423);
or U19528 (N_19528,N_13666,N_10949);
and U19529 (N_19529,N_10039,N_12480);
or U19530 (N_19530,N_13754,N_12159);
or U19531 (N_19531,N_12647,N_11094);
or U19532 (N_19532,N_10645,N_11495);
and U19533 (N_19533,N_14858,N_14662);
or U19534 (N_19534,N_13196,N_11210);
or U19535 (N_19535,N_12959,N_11022);
nand U19536 (N_19536,N_13678,N_12156);
and U19537 (N_19537,N_13422,N_12538);
and U19538 (N_19538,N_10709,N_13290);
and U19539 (N_19539,N_10281,N_10058);
xnor U19540 (N_19540,N_12001,N_11592);
nand U19541 (N_19541,N_11937,N_12946);
nor U19542 (N_19542,N_12033,N_13856);
nand U19543 (N_19543,N_12540,N_11016);
nand U19544 (N_19544,N_12385,N_12355);
xnor U19545 (N_19545,N_12486,N_11910);
and U19546 (N_19546,N_13517,N_10760);
nand U19547 (N_19547,N_11030,N_14388);
or U19548 (N_19548,N_10171,N_11681);
or U19549 (N_19549,N_11048,N_10891);
nor U19550 (N_19550,N_10132,N_11370);
and U19551 (N_19551,N_10813,N_13507);
nor U19552 (N_19552,N_12481,N_14588);
xnor U19553 (N_19553,N_11335,N_14733);
and U19554 (N_19554,N_10048,N_12510);
or U19555 (N_19555,N_11943,N_11695);
or U19556 (N_19556,N_10234,N_12842);
or U19557 (N_19557,N_10934,N_13752);
nand U19558 (N_19558,N_13802,N_12960);
and U19559 (N_19559,N_11663,N_12322);
nor U19560 (N_19560,N_11797,N_13247);
xnor U19561 (N_19561,N_12799,N_12024);
nor U19562 (N_19562,N_13454,N_12205);
or U19563 (N_19563,N_10560,N_13158);
xor U19564 (N_19564,N_11506,N_10007);
nand U19565 (N_19565,N_13430,N_12638);
nand U19566 (N_19566,N_13001,N_10671);
xnor U19567 (N_19567,N_10071,N_11493);
or U19568 (N_19568,N_10864,N_11925);
and U19569 (N_19569,N_13048,N_12827);
and U19570 (N_19570,N_14373,N_12471);
xnor U19571 (N_19571,N_10184,N_11421);
xnor U19572 (N_19572,N_12060,N_13159);
or U19573 (N_19573,N_12536,N_14898);
nor U19574 (N_19574,N_14597,N_12639);
xnor U19575 (N_19575,N_10291,N_12242);
or U19576 (N_19576,N_10471,N_10549);
nand U19577 (N_19577,N_10477,N_10652);
or U19578 (N_19578,N_14225,N_11206);
nor U19579 (N_19579,N_14872,N_12380);
or U19580 (N_19580,N_13208,N_14115);
and U19581 (N_19581,N_12421,N_12352);
nor U19582 (N_19582,N_14329,N_12435);
or U19583 (N_19583,N_11401,N_12743);
nand U19584 (N_19584,N_12921,N_11261);
or U19585 (N_19585,N_10515,N_12112);
nor U19586 (N_19586,N_10182,N_12655);
or U19587 (N_19587,N_10629,N_12878);
nand U19588 (N_19588,N_10727,N_13491);
nor U19589 (N_19589,N_14082,N_11153);
or U19590 (N_19590,N_13663,N_11128);
or U19591 (N_19591,N_13695,N_10757);
or U19592 (N_19592,N_13108,N_11286);
or U19593 (N_19593,N_12708,N_10412);
xnor U19594 (N_19594,N_14888,N_14592);
and U19595 (N_19595,N_13208,N_13493);
and U19596 (N_19596,N_10859,N_10850);
and U19597 (N_19597,N_14270,N_13308);
or U19598 (N_19598,N_11244,N_14002);
nand U19599 (N_19599,N_11344,N_13072);
and U19600 (N_19600,N_13955,N_13402);
nand U19601 (N_19601,N_14608,N_10353);
nand U19602 (N_19602,N_12330,N_14046);
nand U19603 (N_19603,N_12793,N_14550);
or U19604 (N_19604,N_10836,N_10033);
nor U19605 (N_19605,N_14151,N_10844);
nand U19606 (N_19606,N_11147,N_10152);
and U19607 (N_19607,N_14302,N_11962);
or U19608 (N_19608,N_14933,N_13957);
nand U19609 (N_19609,N_12963,N_12207);
and U19610 (N_19610,N_10669,N_11615);
and U19611 (N_19611,N_14830,N_10518);
or U19612 (N_19612,N_11960,N_12256);
or U19613 (N_19613,N_11254,N_13151);
nand U19614 (N_19614,N_10664,N_14111);
or U19615 (N_19615,N_11245,N_10830);
nor U19616 (N_19616,N_11281,N_11256);
nand U19617 (N_19617,N_13824,N_11878);
nand U19618 (N_19618,N_12749,N_11173);
nand U19619 (N_19619,N_12520,N_10745);
nor U19620 (N_19620,N_11955,N_12398);
nor U19621 (N_19621,N_13451,N_13320);
nor U19622 (N_19622,N_13849,N_14843);
and U19623 (N_19623,N_11004,N_14987);
and U19624 (N_19624,N_10967,N_13198);
or U19625 (N_19625,N_11115,N_13981);
or U19626 (N_19626,N_12494,N_12992);
or U19627 (N_19627,N_12791,N_13907);
or U19628 (N_19628,N_10964,N_14577);
or U19629 (N_19629,N_13632,N_12625);
and U19630 (N_19630,N_13801,N_10736);
and U19631 (N_19631,N_13558,N_10922);
or U19632 (N_19632,N_12369,N_13812);
or U19633 (N_19633,N_10140,N_14491);
or U19634 (N_19634,N_11422,N_13682);
xor U19635 (N_19635,N_14462,N_13861);
and U19636 (N_19636,N_10898,N_14394);
and U19637 (N_19637,N_14843,N_13151);
xnor U19638 (N_19638,N_13144,N_13902);
nand U19639 (N_19639,N_10088,N_10760);
nand U19640 (N_19640,N_13208,N_10753);
nor U19641 (N_19641,N_14542,N_10107);
or U19642 (N_19642,N_13101,N_13259);
nor U19643 (N_19643,N_13020,N_12055);
and U19644 (N_19644,N_11118,N_11396);
nor U19645 (N_19645,N_10638,N_10696);
or U19646 (N_19646,N_11217,N_10151);
and U19647 (N_19647,N_13922,N_10594);
or U19648 (N_19648,N_13486,N_14926);
or U19649 (N_19649,N_13249,N_14106);
and U19650 (N_19650,N_12679,N_13797);
nor U19651 (N_19651,N_14745,N_13229);
nand U19652 (N_19652,N_11512,N_11450);
and U19653 (N_19653,N_12846,N_11881);
and U19654 (N_19654,N_13785,N_14176);
nand U19655 (N_19655,N_14039,N_10072);
nor U19656 (N_19656,N_12506,N_10364);
nor U19657 (N_19657,N_11919,N_13999);
nand U19658 (N_19658,N_14126,N_11333);
and U19659 (N_19659,N_11632,N_10801);
and U19660 (N_19660,N_11473,N_10298);
and U19661 (N_19661,N_12922,N_14311);
and U19662 (N_19662,N_10396,N_10313);
and U19663 (N_19663,N_14293,N_13251);
nor U19664 (N_19664,N_12638,N_10574);
nor U19665 (N_19665,N_14316,N_13614);
nand U19666 (N_19666,N_10969,N_12634);
nand U19667 (N_19667,N_13318,N_14429);
nand U19668 (N_19668,N_13314,N_12845);
and U19669 (N_19669,N_11936,N_13126);
and U19670 (N_19670,N_14369,N_11608);
nor U19671 (N_19671,N_10845,N_10498);
nor U19672 (N_19672,N_11168,N_12228);
nor U19673 (N_19673,N_11197,N_14495);
nand U19674 (N_19674,N_10503,N_13658);
nand U19675 (N_19675,N_12299,N_13174);
nand U19676 (N_19676,N_11035,N_13037);
nand U19677 (N_19677,N_11029,N_14737);
nor U19678 (N_19678,N_13632,N_10979);
or U19679 (N_19679,N_10577,N_12487);
and U19680 (N_19680,N_10023,N_12511);
nor U19681 (N_19681,N_10404,N_13464);
nand U19682 (N_19682,N_12431,N_11779);
and U19683 (N_19683,N_10229,N_14846);
and U19684 (N_19684,N_10581,N_10424);
nand U19685 (N_19685,N_11943,N_13075);
nor U19686 (N_19686,N_11233,N_11271);
xor U19687 (N_19687,N_11303,N_14341);
or U19688 (N_19688,N_12999,N_12088);
and U19689 (N_19689,N_12338,N_14088);
or U19690 (N_19690,N_14737,N_13972);
nand U19691 (N_19691,N_11633,N_10738);
nand U19692 (N_19692,N_12162,N_12082);
nor U19693 (N_19693,N_10110,N_10583);
nand U19694 (N_19694,N_12439,N_11214);
or U19695 (N_19695,N_13292,N_13757);
xnor U19696 (N_19696,N_11851,N_10687);
nand U19697 (N_19697,N_14845,N_13246);
or U19698 (N_19698,N_12597,N_14362);
and U19699 (N_19699,N_10469,N_13217);
and U19700 (N_19700,N_10227,N_11536);
nor U19701 (N_19701,N_10489,N_12583);
or U19702 (N_19702,N_10901,N_13402);
nand U19703 (N_19703,N_10042,N_12800);
nor U19704 (N_19704,N_11126,N_12665);
nand U19705 (N_19705,N_11803,N_10134);
and U19706 (N_19706,N_11676,N_10166);
nand U19707 (N_19707,N_13246,N_12617);
and U19708 (N_19708,N_13737,N_12482);
nor U19709 (N_19709,N_13511,N_10747);
nor U19710 (N_19710,N_12267,N_11498);
xnor U19711 (N_19711,N_14761,N_14345);
xor U19712 (N_19712,N_12082,N_11723);
and U19713 (N_19713,N_13022,N_13179);
or U19714 (N_19714,N_11658,N_10066);
xor U19715 (N_19715,N_14336,N_11972);
nor U19716 (N_19716,N_10075,N_14554);
nand U19717 (N_19717,N_11909,N_14031);
nor U19718 (N_19718,N_13652,N_14074);
and U19719 (N_19719,N_13913,N_10215);
and U19720 (N_19720,N_14436,N_14727);
nor U19721 (N_19721,N_12058,N_11905);
nor U19722 (N_19722,N_13192,N_12860);
and U19723 (N_19723,N_11171,N_11298);
or U19724 (N_19724,N_11061,N_10488);
xor U19725 (N_19725,N_12721,N_13885);
or U19726 (N_19726,N_10771,N_11019);
and U19727 (N_19727,N_10329,N_14706);
and U19728 (N_19728,N_14757,N_12845);
nand U19729 (N_19729,N_10343,N_12105);
or U19730 (N_19730,N_12144,N_10281);
nand U19731 (N_19731,N_10318,N_14405);
or U19732 (N_19732,N_10251,N_10851);
and U19733 (N_19733,N_12223,N_10480);
and U19734 (N_19734,N_13165,N_12312);
or U19735 (N_19735,N_12000,N_11337);
xor U19736 (N_19736,N_13620,N_13741);
nor U19737 (N_19737,N_11741,N_11103);
nor U19738 (N_19738,N_10745,N_12290);
and U19739 (N_19739,N_12400,N_14784);
and U19740 (N_19740,N_10618,N_10679);
or U19741 (N_19741,N_12191,N_10795);
or U19742 (N_19742,N_11933,N_12353);
or U19743 (N_19743,N_13337,N_10666);
and U19744 (N_19744,N_11026,N_13749);
or U19745 (N_19745,N_12607,N_13093);
or U19746 (N_19746,N_13564,N_14540);
nor U19747 (N_19747,N_13037,N_11909);
or U19748 (N_19748,N_11908,N_11683);
nor U19749 (N_19749,N_13853,N_10173);
and U19750 (N_19750,N_10684,N_14624);
and U19751 (N_19751,N_11187,N_14917);
xor U19752 (N_19752,N_13414,N_13057);
or U19753 (N_19753,N_12911,N_12628);
nor U19754 (N_19754,N_10484,N_13525);
or U19755 (N_19755,N_12001,N_14845);
and U19756 (N_19756,N_10599,N_10461);
or U19757 (N_19757,N_10760,N_14875);
or U19758 (N_19758,N_13587,N_13008);
nand U19759 (N_19759,N_14409,N_10631);
nand U19760 (N_19760,N_13052,N_12248);
nand U19761 (N_19761,N_13672,N_11494);
or U19762 (N_19762,N_14344,N_12729);
and U19763 (N_19763,N_11789,N_13383);
nor U19764 (N_19764,N_12569,N_14120);
or U19765 (N_19765,N_10324,N_10953);
and U19766 (N_19766,N_11328,N_12560);
nand U19767 (N_19767,N_10933,N_11616);
nor U19768 (N_19768,N_12324,N_14799);
nand U19769 (N_19769,N_12530,N_12947);
or U19770 (N_19770,N_10170,N_12084);
and U19771 (N_19771,N_10418,N_10982);
or U19772 (N_19772,N_13620,N_11514);
nand U19773 (N_19773,N_12516,N_12699);
or U19774 (N_19774,N_14520,N_10097);
or U19775 (N_19775,N_14058,N_11795);
nand U19776 (N_19776,N_11718,N_14754);
nor U19777 (N_19777,N_12015,N_14820);
nor U19778 (N_19778,N_12477,N_14825);
nand U19779 (N_19779,N_12270,N_10246);
xor U19780 (N_19780,N_10531,N_13269);
nand U19781 (N_19781,N_10034,N_13078);
nor U19782 (N_19782,N_14939,N_11900);
or U19783 (N_19783,N_10111,N_11358);
nor U19784 (N_19784,N_12041,N_14265);
xnor U19785 (N_19785,N_11432,N_12990);
and U19786 (N_19786,N_13878,N_14228);
nor U19787 (N_19787,N_14235,N_13338);
or U19788 (N_19788,N_11996,N_10979);
and U19789 (N_19789,N_10865,N_13292);
nand U19790 (N_19790,N_13470,N_14396);
nand U19791 (N_19791,N_11678,N_14548);
xnor U19792 (N_19792,N_10975,N_12626);
or U19793 (N_19793,N_11535,N_14028);
xnor U19794 (N_19794,N_12595,N_12194);
or U19795 (N_19795,N_12597,N_13687);
nand U19796 (N_19796,N_13080,N_12230);
and U19797 (N_19797,N_10919,N_14689);
nand U19798 (N_19798,N_11152,N_11592);
nand U19799 (N_19799,N_12566,N_12919);
and U19800 (N_19800,N_11472,N_14335);
nor U19801 (N_19801,N_10664,N_12416);
nand U19802 (N_19802,N_11613,N_11709);
nand U19803 (N_19803,N_10327,N_12876);
nor U19804 (N_19804,N_13247,N_14701);
nor U19805 (N_19805,N_12189,N_13786);
and U19806 (N_19806,N_12786,N_12084);
or U19807 (N_19807,N_14628,N_12824);
and U19808 (N_19808,N_12775,N_11499);
nor U19809 (N_19809,N_10414,N_14393);
and U19810 (N_19810,N_13055,N_13911);
nand U19811 (N_19811,N_10392,N_10782);
nor U19812 (N_19812,N_11839,N_10410);
and U19813 (N_19813,N_11671,N_12556);
or U19814 (N_19814,N_14006,N_13780);
or U19815 (N_19815,N_12924,N_14404);
nand U19816 (N_19816,N_10826,N_10358);
nor U19817 (N_19817,N_10419,N_10152);
xor U19818 (N_19818,N_13615,N_14564);
nand U19819 (N_19819,N_11647,N_14372);
and U19820 (N_19820,N_14408,N_14466);
nand U19821 (N_19821,N_14887,N_12798);
nand U19822 (N_19822,N_12399,N_13808);
nor U19823 (N_19823,N_11310,N_11630);
nand U19824 (N_19824,N_10137,N_13812);
and U19825 (N_19825,N_14573,N_10256);
or U19826 (N_19826,N_14725,N_14468);
or U19827 (N_19827,N_11339,N_11018);
xor U19828 (N_19828,N_14522,N_13583);
or U19829 (N_19829,N_13459,N_13858);
and U19830 (N_19830,N_13785,N_13379);
nand U19831 (N_19831,N_14146,N_13254);
or U19832 (N_19832,N_13830,N_12568);
and U19833 (N_19833,N_14110,N_14140);
and U19834 (N_19834,N_13002,N_14145);
xnor U19835 (N_19835,N_11635,N_10370);
or U19836 (N_19836,N_11483,N_11393);
nor U19837 (N_19837,N_10220,N_13868);
nand U19838 (N_19838,N_11207,N_11938);
and U19839 (N_19839,N_10841,N_10950);
nand U19840 (N_19840,N_11787,N_14363);
nor U19841 (N_19841,N_11077,N_11409);
nor U19842 (N_19842,N_13671,N_11499);
and U19843 (N_19843,N_10129,N_10582);
and U19844 (N_19844,N_14588,N_11234);
or U19845 (N_19845,N_12703,N_12496);
nor U19846 (N_19846,N_10539,N_10574);
and U19847 (N_19847,N_12805,N_11303);
nand U19848 (N_19848,N_12669,N_14437);
nand U19849 (N_19849,N_13645,N_14735);
and U19850 (N_19850,N_12374,N_14009);
and U19851 (N_19851,N_10581,N_11501);
nand U19852 (N_19852,N_11777,N_10049);
xnor U19853 (N_19853,N_14564,N_14891);
or U19854 (N_19854,N_12204,N_10649);
nand U19855 (N_19855,N_12796,N_12188);
and U19856 (N_19856,N_12431,N_14164);
nand U19857 (N_19857,N_13406,N_14481);
or U19858 (N_19858,N_12253,N_11434);
and U19859 (N_19859,N_14388,N_12767);
or U19860 (N_19860,N_12823,N_12878);
and U19861 (N_19861,N_11566,N_13670);
or U19862 (N_19862,N_12980,N_12309);
nor U19863 (N_19863,N_10755,N_12891);
nand U19864 (N_19864,N_12850,N_11141);
or U19865 (N_19865,N_11447,N_12997);
and U19866 (N_19866,N_14878,N_12924);
nor U19867 (N_19867,N_14222,N_14699);
nor U19868 (N_19868,N_10545,N_10300);
nor U19869 (N_19869,N_11291,N_10611);
nand U19870 (N_19870,N_12380,N_10954);
nand U19871 (N_19871,N_13208,N_11023);
nor U19872 (N_19872,N_11038,N_11599);
and U19873 (N_19873,N_12629,N_12067);
nor U19874 (N_19874,N_14924,N_12449);
and U19875 (N_19875,N_12869,N_13757);
xor U19876 (N_19876,N_14786,N_14955);
or U19877 (N_19877,N_14680,N_10336);
or U19878 (N_19878,N_13804,N_11237);
nor U19879 (N_19879,N_10441,N_10028);
nor U19880 (N_19880,N_12660,N_13694);
and U19881 (N_19881,N_11971,N_12980);
xor U19882 (N_19882,N_12069,N_13153);
and U19883 (N_19883,N_13641,N_10030);
nand U19884 (N_19884,N_11908,N_13966);
nand U19885 (N_19885,N_12948,N_14113);
or U19886 (N_19886,N_13509,N_11111);
xnor U19887 (N_19887,N_14818,N_10321);
and U19888 (N_19888,N_12476,N_13205);
xnor U19889 (N_19889,N_11992,N_13699);
and U19890 (N_19890,N_13212,N_11992);
and U19891 (N_19891,N_13879,N_11066);
and U19892 (N_19892,N_10486,N_13152);
or U19893 (N_19893,N_13166,N_14981);
nor U19894 (N_19894,N_14156,N_10420);
nand U19895 (N_19895,N_14380,N_12497);
xor U19896 (N_19896,N_13972,N_14355);
or U19897 (N_19897,N_12378,N_12720);
or U19898 (N_19898,N_12442,N_13241);
and U19899 (N_19899,N_10190,N_14712);
nand U19900 (N_19900,N_10627,N_14228);
nand U19901 (N_19901,N_12198,N_13818);
and U19902 (N_19902,N_12745,N_12415);
and U19903 (N_19903,N_13682,N_12958);
or U19904 (N_19904,N_14212,N_11078);
and U19905 (N_19905,N_13995,N_13264);
nor U19906 (N_19906,N_10347,N_12147);
and U19907 (N_19907,N_10888,N_13373);
nor U19908 (N_19908,N_13399,N_10703);
or U19909 (N_19909,N_12393,N_11841);
nor U19910 (N_19910,N_12972,N_12893);
and U19911 (N_19911,N_14157,N_13507);
or U19912 (N_19912,N_10959,N_12380);
nor U19913 (N_19913,N_13885,N_12566);
nand U19914 (N_19914,N_11427,N_11259);
nor U19915 (N_19915,N_11676,N_12649);
nor U19916 (N_19916,N_12234,N_14746);
or U19917 (N_19917,N_11850,N_12299);
nand U19918 (N_19918,N_10397,N_10968);
and U19919 (N_19919,N_11445,N_10698);
or U19920 (N_19920,N_14625,N_13429);
or U19921 (N_19921,N_14367,N_10202);
and U19922 (N_19922,N_10560,N_13930);
nand U19923 (N_19923,N_10671,N_11184);
nor U19924 (N_19924,N_11618,N_13446);
and U19925 (N_19925,N_12247,N_11206);
nor U19926 (N_19926,N_11140,N_10795);
and U19927 (N_19927,N_10006,N_14728);
nor U19928 (N_19928,N_13811,N_14241);
or U19929 (N_19929,N_12240,N_12872);
or U19930 (N_19930,N_10032,N_14526);
nor U19931 (N_19931,N_11387,N_12759);
nor U19932 (N_19932,N_13494,N_12227);
nand U19933 (N_19933,N_11930,N_10889);
xor U19934 (N_19934,N_10090,N_11413);
or U19935 (N_19935,N_13679,N_13129);
or U19936 (N_19936,N_13567,N_14855);
and U19937 (N_19937,N_13089,N_11054);
and U19938 (N_19938,N_10913,N_11686);
and U19939 (N_19939,N_11019,N_13317);
and U19940 (N_19940,N_14483,N_11505);
nor U19941 (N_19941,N_11570,N_13930);
nor U19942 (N_19942,N_10554,N_10547);
and U19943 (N_19943,N_10626,N_14505);
and U19944 (N_19944,N_11256,N_10241);
or U19945 (N_19945,N_12809,N_14388);
and U19946 (N_19946,N_10961,N_14465);
nor U19947 (N_19947,N_13344,N_10205);
or U19948 (N_19948,N_13327,N_11358);
and U19949 (N_19949,N_12696,N_14770);
and U19950 (N_19950,N_14651,N_12144);
and U19951 (N_19951,N_12106,N_11818);
or U19952 (N_19952,N_10763,N_13769);
and U19953 (N_19953,N_14402,N_14651);
nor U19954 (N_19954,N_10137,N_13277);
nor U19955 (N_19955,N_12524,N_13069);
xnor U19956 (N_19956,N_12353,N_12080);
and U19957 (N_19957,N_11556,N_12706);
nor U19958 (N_19958,N_12908,N_13170);
nand U19959 (N_19959,N_14350,N_13053);
nand U19960 (N_19960,N_10199,N_14475);
or U19961 (N_19961,N_14170,N_10688);
nor U19962 (N_19962,N_10113,N_14630);
or U19963 (N_19963,N_10984,N_11435);
nor U19964 (N_19964,N_14089,N_12653);
xnor U19965 (N_19965,N_14131,N_14852);
nor U19966 (N_19966,N_12123,N_13536);
xnor U19967 (N_19967,N_12226,N_13791);
nand U19968 (N_19968,N_10221,N_13753);
nand U19969 (N_19969,N_13837,N_11265);
and U19970 (N_19970,N_13933,N_10921);
nor U19971 (N_19971,N_13111,N_11719);
or U19972 (N_19972,N_11569,N_13908);
and U19973 (N_19973,N_13894,N_12804);
or U19974 (N_19974,N_12369,N_10079);
or U19975 (N_19975,N_11207,N_10844);
xor U19976 (N_19976,N_14974,N_12263);
and U19977 (N_19977,N_10706,N_10111);
nor U19978 (N_19978,N_13728,N_14715);
and U19979 (N_19979,N_11708,N_12681);
nand U19980 (N_19980,N_11406,N_14915);
and U19981 (N_19981,N_12432,N_12316);
nand U19982 (N_19982,N_11345,N_13441);
and U19983 (N_19983,N_13280,N_13380);
and U19984 (N_19984,N_13762,N_12485);
nor U19985 (N_19985,N_13481,N_10405);
and U19986 (N_19986,N_10708,N_12814);
nor U19987 (N_19987,N_12986,N_13547);
and U19988 (N_19988,N_14186,N_12589);
nor U19989 (N_19989,N_13606,N_14845);
nor U19990 (N_19990,N_14680,N_11567);
nor U19991 (N_19991,N_11652,N_14412);
nor U19992 (N_19992,N_13250,N_14326);
xnor U19993 (N_19993,N_13174,N_12277);
nand U19994 (N_19994,N_14597,N_13577);
nand U19995 (N_19995,N_14704,N_14303);
or U19996 (N_19996,N_12738,N_12511);
xor U19997 (N_19997,N_11881,N_14138);
xnor U19998 (N_19998,N_12040,N_11584);
and U19999 (N_19999,N_12513,N_14255);
and UO_0 (O_0,N_19328,N_15841);
nor UO_1 (O_1,N_17033,N_18188);
and UO_2 (O_2,N_19107,N_19555);
and UO_3 (O_3,N_18170,N_16933);
and UO_4 (O_4,N_16039,N_19904);
or UO_5 (O_5,N_15246,N_16961);
or UO_6 (O_6,N_19611,N_15745);
or UO_7 (O_7,N_17347,N_15895);
and UO_8 (O_8,N_16443,N_16553);
nor UO_9 (O_9,N_16572,N_19286);
nand UO_10 (O_10,N_19819,N_16848);
xor UO_11 (O_11,N_15078,N_16918);
or UO_12 (O_12,N_15660,N_19241);
xnor UO_13 (O_13,N_16878,N_17631);
or UO_14 (O_14,N_18720,N_15969);
or UO_15 (O_15,N_17513,N_17079);
nand UO_16 (O_16,N_18364,N_15467);
and UO_17 (O_17,N_18892,N_18930);
and UO_18 (O_18,N_16737,N_15164);
and UO_19 (O_19,N_15489,N_19367);
and UO_20 (O_20,N_15705,N_16482);
or UO_21 (O_21,N_17633,N_16461);
and UO_22 (O_22,N_16895,N_19894);
nand UO_23 (O_23,N_15444,N_18347);
nor UO_24 (O_24,N_19086,N_19934);
nor UO_25 (O_25,N_15712,N_17086);
and UO_26 (O_26,N_19280,N_15798);
nor UO_27 (O_27,N_19251,N_18527);
nand UO_28 (O_28,N_18161,N_19988);
and UO_29 (O_29,N_18145,N_19604);
xnor UO_30 (O_30,N_15183,N_15018);
or UO_31 (O_31,N_16199,N_19689);
nand UO_32 (O_32,N_19545,N_15089);
nor UO_33 (O_33,N_15657,N_15172);
and UO_34 (O_34,N_15837,N_18244);
nor UO_35 (O_35,N_17746,N_19309);
or UO_36 (O_36,N_17630,N_15939);
nand UO_37 (O_37,N_19794,N_17139);
nand UO_38 (O_38,N_15200,N_19900);
nor UO_39 (O_39,N_19989,N_17761);
and UO_40 (O_40,N_15612,N_18653);
xnor UO_41 (O_41,N_16323,N_16021);
or UO_42 (O_42,N_16987,N_18210);
and UO_43 (O_43,N_15131,N_18383);
and UO_44 (O_44,N_17243,N_18701);
xnor UO_45 (O_45,N_18471,N_19351);
nand UO_46 (O_46,N_18135,N_15373);
nand UO_47 (O_47,N_16359,N_19722);
and UO_48 (O_48,N_18676,N_15214);
nor UO_49 (O_49,N_18013,N_17219);
and UO_50 (O_50,N_16787,N_16285);
or UO_51 (O_51,N_17453,N_18940);
nor UO_52 (O_52,N_17135,N_19256);
nand UO_53 (O_53,N_17790,N_15258);
xor UO_54 (O_54,N_19986,N_16023);
nand UO_55 (O_55,N_15976,N_17388);
and UO_56 (O_56,N_15479,N_19291);
nor UO_57 (O_57,N_17977,N_17458);
and UO_58 (O_58,N_16405,N_16994);
nand UO_59 (O_59,N_19433,N_15898);
or UO_60 (O_60,N_18158,N_18057);
and UO_61 (O_61,N_17339,N_18163);
or UO_62 (O_62,N_17938,N_19198);
or UO_63 (O_63,N_16432,N_19752);
nand UO_64 (O_64,N_19508,N_19719);
and UO_65 (O_65,N_19737,N_17333);
or UO_66 (O_66,N_19909,N_16583);
or UO_67 (O_67,N_18618,N_17559);
or UO_68 (O_68,N_18632,N_17989);
nand UO_69 (O_69,N_15516,N_17676);
or UO_70 (O_70,N_15577,N_16701);
and UO_71 (O_71,N_16828,N_19827);
and UO_72 (O_72,N_18900,N_18438);
nand UO_73 (O_73,N_19124,N_19503);
nor UO_74 (O_74,N_15344,N_19780);
or UO_75 (O_75,N_15377,N_18523);
nor UO_76 (O_76,N_17907,N_16166);
nand UO_77 (O_77,N_19427,N_18081);
and UO_78 (O_78,N_19963,N_18556);
or UO_79 (O_79,N_19961,N_17999);
or UO_80 (O_80,N_18528,N_18571);
and UO_81 (O_81,N_16379,N_15253);
or UO_82 (O_82,N_18704,N_17853);
nor UO_83 (O_83,N_18146,N_17164);
nand UO_84 (O_84,N_18069,N_19535);
and UO_85 (O_85,N_18726,N_18659);
nand UO_86 (O_86,N_15825,N_17315);
nor UO_87 (O_87,N_18834,N_19643);
xnor UO_88 (O_88,N_18058,N_19495);
or UO_89 (O_89,N_19873,N_18519);
or UO_90 (O_90,N_15958,N_18059);
xor UO_91 (O_91,N_17457,N_18633);
or UO_92 (O_92,N_18225,N_15379);
or UO_93 (O_93,N_17175,N_19959);
nor UO_94 (O_94,N_19239,N_17272);
xor UO_95 (O_95,N_17779,N_18533);
xnor UO_96 (O_96,N_19553,N_16508);
or UO_97 (O_97,N_16065,N_15213);
nand UO_98 (O_98,N_19790,N_19217);
nor UO_99 (O_99,N_18048,N_19592);
xor UO_100 (O_100,N_19522,N_17495);
nor UO_101 (O_101,N_16084,N_18344);
nand UO_102 (O_102,N_16634,N_16739);
and UO_103 (O_103,N_15486,N_18989);
nand UO_104 (O_104,N_15238,N_19352);
and UO_105 (O_105,N_19143,N_18508);
nand UO_106 (O_106,N_16451,N_16160);
nor UO_107 (O_107,N_15284,N_17529);
nor UO_108 (O_108,N_18346,N_18790);
nor UO_109 (O_109,N_16085,N_16757);
and UO_110 (O_110,N_15404,N_17193);
nor UO_111 (O_111,N_15628,N_16389);
nor UO_112 (O_112,N_15362,N_18299);
nand UO_113 (O_113,N_16398,N_17072);
and UO_114 (O_114,N_17891,N_17874);
nand UO_115 (O_115,N_19785,N_19945);
xnor UO_116 (O_116,N_16712,N_15747);
and UO_117 (O_117,N_16666,N_19318);
and UO_118 (O_118,N_16804,N_17307);
or UO_119 (O_119,N_18159,N_15891);
and UO_120 (O_120,N_17183,N_15600);
nand UO_121 (O_121,N_18501,N_17961);
nand UO_122 (O_122,N_15524,N_15610);
xor UO_123 (O_123,N_17334,N_17739);
and UO_124 (O_124,N_18491,N_15512);
and UO_125 (O_125,N_19551,N_15527);
nand UO_126 (O_126,N_16346,N_19577);
nand UO_127 (O_127,N_17492,N_16514);
and UO_128 (O_128,N_16022,N_15729);
nor UO_129 (O_129,N_17295,N_18055);
xor UO_130 (O_130,N_19225,N_18702);
nor UO_131 (O_131,N_16148,N_16274);
and UO_132 (O_132,N_16251,N_16955);
nor UO_133 (O_133,N_15796,N_16853);
nor UO_134 (O_134,N_19080,N_15926);
or UO_135 (O_135,N_18875,N_17800);
or UO_136 (O_136,N_18411,N_16225);
and UO_137 (O_137,N_15053,N_18607);
nand UO_138 (O_138,N_18601,N_15268);
or UO_139 (O_139,N_18967,N_15643);
nand UO_140 (O_140,N_15445,N_18973);
nand UO_141 (O_141,N_15616,N_17301);
and UO_142 (O_142,N_19154,N_17053);
nor UO_143 (O_143,N_16256,N_17312);
or UO_144 (O_144,N_15782,N_17268);
or UO_145 (O_145,N_17979,N_19046);
and UO_146 (O_146,N_17925,N_15582);
nand UO_147 (O_147,N_18128,N_18304);
nor UO_148 (O_148,N_17768,N_17230);
and UO_149 (O_149,N_15573,N_15222);
and UO_150 (O_150,N_17256,N_19303);
nor UO_151 (O_151,N_18788,N_18157);
nor UO_152 (O_152,N_15431,N_17075);
nor UO_153 (O_153,N_18578,N_15276);
nand UO_154 (O_154,N_16880,N_19890);
and UO_155 (O_155,N_15642,N_17255);
and UO_156 (O_156,N_15171,N_16009);
nand UO_157 (O_157,N_19725,N_19081);
nand UO_158 (O_158,N_15567,N_15843);
and UO_159 (O_159,N_17832,N_15069);
nand UO_160 (O_160,N_19616,N_16462);
nand UO_161 (O_161,N_18511,N_19159);
or UO_162 (O_162,N_15039,N_18339);
and UO_163 (O_163,N_16178,N_16203);
nand UO_164 (O_164,N_18742,N_15314);
nand UO_165 (O_165,N_17618,N_17187);
or UO_166 (O_166,N_17305,N_18166);
and UO_167 (O_167,N_19369,N_18851);
nor UO_168 (O_168,N_17246,N_19492);
and UO_169 (O_169,N_17881,N_18454);
or UO_170 (O_170,N_16117,N_18390);
or UO_171 (O_171,N_17944,N_18382);
nand UO_172 (O_172,N_16344,N_17261);
nor UO_173 (O_173,N_16399,N_19777);
and UO_174 (O_174,N_18015,N_15033);
nand UO_175 (O_175,N_19110,N_19304);
nand UO_176 (O_176,N_18806,N_16381);
nand UO_177 (O_177,N_19717,N_18588);
or UO_178 (O_178,N_17990,N_17705);
nor UO_179 (O_179,N_18760,N_15149);
and UO_180 (O_180,N_15371,N_15700);
or UO_181 (O_181,N_18557,N_17461);
nand UO_182 (O_182,N_17600,N_16920);
or UO_183 (O_183,N_16352,N_18494);
nor UO_184 (O_184,N_19911,N_17915);
nor UO_185 (O_185,N_18634,N_15988);
nor UO_186 (O_186,N_19798,N_16005);
nand UO_187 (O_187,N_15147,N_18253);
or UO_188 (O_188,N_16836,N_15071);
or UO_189 (O_189,N_17273,N_19603);
nor UO_190 (O_190,N_17992,N_15230);
nor UO_191 (O_191,N_15332,N_19035);
or UO_192 (O_192,N_15739,N_15795);
nor UO_193 (O_193,N_15182,N_15554);
nand UO_194 (O_194,N_18456,N_17632);
or UO_195 (O_195,N_18071,N_16056);
and UO_196 (O_196,N_16128,N_18190);
nand UO_197 (O_197,N_19467,N_16142);
or UO_198 (O_198,N_18833,N_15493);
and UO_199 (O_199,N_18045,N_16149);
and UO_200 (O_200,N_15336,N_18223);
or UO_201 (O_201,N_18226,N_18078);
xor UO_202 (O_202,N_15542,N_15596);
nor UO_203 (O_203,N_19997,N_17393);
and UO_204 (O_204,N_19138,N_15828);
xor UO_205 (O_205,N_19131,N_16717);
and UO_206 (O_206,N_15394,N_15264);
nand UO_207 (O_207,N_17982,N_16331);
nand UO_208 (O_208,N_17427,N_19388);
and UO_209 (O_209,N_19916,N_17332);
and UO_210 (O_210,N_19812,N_17593);
xor UO_211 (O_211,N_19016,N_15223);
nor UO_212 (O_212,N_19339,N_19899);
and UO_213 (O_213,N_16301,N_19970);
or UO_214 (O_214,N_19552,N_19126);
and UO_215 (O_215,N_16893,N_16146);
nand UO_216 (O_216,N_18999,N_18970);
and UO_217 (O_217,N_17698,N_19956);
nor UO_218 (O_218,N_17184,N_19041);
or UO_219 (O_219,N_19704,N_18737);
xor UO_220 (O_220,N_16721,N_15821);
and UO_221 (O_221,N_18112,N_19820);
nor UO_222 (O_222,N_17935,N_19562);
nand UO_223 (O_223,N_18904,N_15154);
nor UO_224 (O_224,N_16358,N_15101);
or UO_225 (O_225,N_19636,N_17744);
nor UO_226 (O_226,N_15429,N_15911);
nand UO_227 (O_227,N_19377,N_16280);
or UO_228 (O_228,N_17387,N_18040);
xnor UO_229 (O_229,N_18958,N_15991);
xor UO_230 (O_230,N_19343,N_17176);
or UO_231 (O_231,N_17238,N_19773);
and UO_232 (O_232,N_15529,N_15664);
nor UO_233 (O_233,N_19907,N_18336);
nor UO_234 (O_234,N_18895,N_19795);
or UO_235 (O_235,N_17823,N_17249);
nand UO_236 (O_236,N_18481,N_16778);
and UO_237 (O_237,N_15631,N_15060);
xor UO_238 (O_238,N_18110,N_15714);
nand UO_239 (O_239,N_15094,N_18550);
xor UO_240 (O_240,N_19826,N_18888);
xnor UO_241 (O_241,N_18100,N_17995);
xnor UO_242 (O_242,N_17488,N_16179);
nand UO_243 (O_243,N_17740,N_15755);
nand UO_244 (O_244,N_18591,N_16490);
nand UO_245 (O_245,N_16977,N_17251);
nor UO_246 (O_246,N_16281,N_19664);
and UO_247 (O_247,N_15923,N_15565);
nor UO_248 (O_248,N_15966,N_17479);
and UO_249 (O_249,N_15557,N_18484);
xnor UO_250 (O_250,N_17099,N_17627);
nor UO_251 (O_251,N_17793,N_17693);
or UO_252 (O_252,N_18093,N_19836);
nor UO_253 (O_253,N_15945,N_18010);
xnor UO_254 (O_254,N_19585,N_19044);
and UO_255 (O_255,N_16581,N_18130);
and UO_256 (O_256,N_18692,N_16187);
or UO_257 (O_257,N_15023,N_19075);
nand UO_258 (O_258,N_16485,N_15068);
nand UO_259 (O_259,N_17808,N_19702);
and UO_260 (O_260,N_17549,N_17406);
nor UO_261 (O_261,N_15417,N_19236);
xor UO_262 (O_262,N_18937,N_15629);
and UO_263 (O_263,N_18766,N_18265);
nand UO_264 (O_264,N_15648,N_18290);
nor UO_265 (O_265,N_15772,N_18561);
and UO_266 (O_266,N_15749,N_17362);
or UO_267 (O_267,N_18509,N_17769);
nor UO_268 (O_268,N_18477,N_19036);
and UO_269 (O_269,N_17550,N_17004);
nor UO_270 (O_270,N_15405,N_18635);
xor UO_271 (O_271,N_15269,N_18736);
nor UO_272 (O_272,N_19308,N_16913);
and UO_273 (O_273,N_18427,N_15151);
nor UO_274 (O_274,N_18639,N_16667);
nor UO_275 (O_275,N_19457,N_15451);
and UO_276 (O_276,N_18710,N_15408);
and UO_277 (O_277,N_19314,N_15982);
nand UO_278 (O_278,N_16713,N_18312);
nor UO_279 (O_279,N_15838,N_16515);
or UO_280 (O_280,N_18001,N_15402);
or UO_281 (O_281,N_18345,N_15862);
nor UO_282 (O_282,N_19385,N_17998);
and UO_283 (O_283,N_19077,N_17847);
and UO_284 (O_284,N_18132,N_16525);
nand UO_285 (O_285,N_19647,N_16540);
nor UO_286 (O_286,N_18552,N_19902);
xnor UO_287 (O_287,N_16560,N_19432);
nor UO_288 (O_288,N_17002,N_16590);
and UO_289 (O_289,N_18577,N_16397);
xor UO_290 (O_290,N_18952,N_18106);
xnor UO_291 (O_291,N_18263,N_15196);
xor UO_292 (O_292,N_19881,N_16248);
and UO_293 (O_293,N_15770,N_16837);
or UO_294 (O_294,N_18986,N_16332);
nor UO_295 (O_295,N_18053,N_17781);
nand UO_296 (O_296,N_18361,N_19865);
nand UO_297 (O_297,N_16830,N_15502);
nand UO_298 (O_298,N_19823,N_15879);
nor UO_299 (O_299,N_16219,N_19923);
or UO_300 (O_300,N_19207,N_16827);
nand UO_301 (O_301,N_17599,N_17217);
nor UO_302 (O_302,N_16580,N_17590);
nor UO_303 (O_303,N_19735,N_16137);
nand UO_304 (O_304,N_18211,N_19515);
nand UO_305 (O_305,N_18934,N_18960);
or UO_306 (O_306,N_18352,N_17519);
and UO_307 (O_307,N_19056,N_19258);
nand UO_308 (O_308,N_18379,N_18741);
or UO_309 (O_309,N_15312,N_19676);
nand UO_310 (O_310,N_16992,N_15024);
nor UO_311 (O_311,N_18683,N_17097);
nor UO_312 (O_312,N_17379,N_19335);
and UO_313 (O_313,N_17207,N_16158);
nand UO_314 (O_314,N_18184,N_16528);
nand UO_315 (O_315,N_19268,N_19279);
xnor UO_316 (O_316,N_19320,N_19638);
or UO_317 (O_317,N_15615,N_19569);
or UO_318 (O_318,N_15849,N_17205);
nand UO_319 (O_319,N_16211,N_17724);
xnor UO_320 (O_320,N_17893,N_18232);
xor UO_321 (O_321,N_17530,N_17515);
nor UO_322 (O_322,N_17786,N_19749);
xnor UO_323 (O_323,N_17770,N_15418);
or UO_324 (O_324,N_17497,N_16760);
or UO_325 (O_325,N_19912,N_17959);
and UO_326 (O_326,N_17442,N_18972);
and UO_327 (O_327,N_16619,N_15986);
or UO_328 (O_328,N_17277,N_17372);
and UO_329 (O_329,N_15128,N_18275);
xnor UO_330 (O_330,N_19982,N_17452);
nor UO_331 (O_331,N_19891,N_15971);
and UO_332 (O_332,N_19629,N_19858);
nand UO_333 (O_333,N_18175,N_19549);
or UO_334 (O_334,N_15801,N_19195);
nand UO_335 (O_335,N_17023,N_18668);
or UO_336 (O_336,N_18418,N_16147);
and UO_337 (O_337,N_19696,N_19511);
and UO_338 (O_338,N_17532,N_19175);
nor UO_339 (O_339,N_18472,N_17250);
nand UO_340 (O_340,N_17548,N_18302);
nand UO_341 (O_341,N_16218,N_16202);
or UO_342 (O_342,N_18763,N_16373);
and UO_343 (O_343,N_19659,N_16393);
nand UO_344 (O_344,N_18532,N_16569);
nor UO_345 (O_345,N_15446,N_16229);
or UO_346 (O_346,N_19142,N_17358);
or UO_347 (O_347,N_19979,N_17008);
or UO_348 (O_348,N_17446,N_15623);
xnor UO_349 (O_349,N_17066,N_15523);
nand UO_350 (O_350,N_18306,N_15834);
and UO_351 (O_351,N_15165,N_17748);
and UO_352 (O_352,N_16134,N_17665);
or UO_353 (O_353,N_18560,N_15924);
nand UO_354 (O_354,N_16777,N_16557);
nand UO_355 (O_355,N_16078,N_17049);
nand UO_356 (O_356,N_16050,N_16896);
or UO_357 (O_357,N_16849,N_17120);
and UO_358 (O_358,N_16466,N_17303);
xnor UO_359 (O_359,N_17240,N_17540);
nand UO_360 (O_360,N_17395,N_15630);
and UO_361 (O_361,N_18991,N_16240);
or UO_362 (O_362,N_19300,N_19797);
nor UO_363 (O_363,N_16457,N_18630);
xnor UO_364 (O_364,N_15427,N_16965);
or UO_365 (O_365,N_19205,N_16136);
or UO_366 (O_366,N_15166,N_17192);
nand UO_367 (O_367,N_17487,N_17162);
xnor UO_368 (O_368,N_19751,N_18419);
nand UO_369 (O_369,N_18370,N_18152);
nand UO_370 (O_370,N_17241,N_18753);
nor UO_371 (O_371,N_19344,N_16618);
nand UO_372 (O_372,N_17719,N_15586);
nor UO_373 (O_373,N_19017,N_15548);
or UO_374 (O_374,N_19188,N_16150);
and UO_375 (O_375,N_15706,N_17143);
nand UO_376 (O_376,N_19333,N_16861);
or UO_377 (O_377,N_16646,N_19209);
xnor UO_378 (O_378,N_18899,N_17258);
nor UO_379 (O_379,N_15666,N_19048);
nand UO_380 (O_380,N_16803,N_15295);
and UO_381 (O_381,N_17582,N_18220);
or UO_382 (O_382,N_17280,N_15977);
or UO_383 (O_383,N_18317,N_18745);
nor UO_384 (O_384,N_18880,N_19257);
nand UO_385 (O_385,N_15607,N_16247);
and UO_386 (O_386,N_17010,N_15127);
nor UO_387 (O_387,N_15979,N_18727);
xor UO_388 (O_388,N_19224,N_19399);
and UO_389 (O_389,N_15719,N_16386);
nand UO_390 (O_390,N_17991,N_16745);
xor UO_391 (O_391,N_17366,N_19960);
xor UO_392 (O_392,N_15448,N_15870);
nor UO_393 (O_393,N_19509,N_16885);
and UO_394 (O_394,N_15475,N_18890);
xor UO_395 (O_395,N_18927,N_17730);
or UO_396 (O_396,N_15647,N_15217);
nand UO_397 (O_397,N_16636,N_15231);
nor UO_398 (O_398,N_15494,N_15140);
nor UO_399 (O_399,N_17024,N_15964);
and UO_400 (O_400,N_16173,N_17231);
nand UO_401 (O_401,N_18043,N_19254);
nor UO_402 (O_402,N_17782,N_18358);
and UO_403 (O_403,N_18311,N_17602);
and UO_404 (O_404,N_15161,N_18708);
or UO_405 (O_405,N_17741,N_16756);
nand UO_406 (O_406,N_16840,N_15360);
and UO_407 (O_407,N_16270,N_17063);
xnor UO_408 (O_408,N_15084,N_17531);
nand UO_409 (O_409,N_18155,N_15370);
or UO_410 (O_410,N_17073,N_19134);
nor UO_411 (O_411,N_19578,N_19738);
nor UO_412 (O_412,N_17061,N_16626);
or UO_413 (O_413,N_19615,N_19029);
and UO_414 (O_414,N_19178,N_16384);
or UO_415 (O_415,N_16582,N_18993);
nor UO_416 (O_416,N_15345,N_18307);
or UO_417 (O_417,N_18950,N_17096);
and UO_418 (O_418,N_19071,N_15918);
and UO_419 (O_419,N_15818,N_19831);
nor UO_420 (O_420,N_19893,N_19830);
and UO_421 (O_421,N_18463,N_17279);
xor UO_422 (O_422,N_18629,N_17996);
and UO_423 (O_423,N_16174,N_15163);
and UO_424 (O_424,N_18261,N_17521);
xnor UO_425 (O_425,N_15454,N_18474);
or UO_426 (O_426,N_16703,N_17860);
nor UO_427 (O_427,N_17344,N_18848);
nand UO_428 (O_428,N_16228,N_18118);
or UO_429 (O_429,N_16993,N_19272);
nand UO_430 (O_430,N_16551,N_15595);
nor UO_431 (O_431,N_15889,N_18189);
nor UO_432 (O_432,N_16894,N_17975);
nor UO_433 (O_433,N_19665,N_15553);
or UO_434 (O_434,N_19033,N_16753);
and UO_435 (O_435,N_18531,N_16113);
nand UO_436 (O_436,N_15287,N_17262);
or UO_437 (O_437,N_18156,N_18667);
or UO_438 (O_438,N_16099,N_16017);
nand UO_439 (O_439,N_17364,N_17114);
and UO_440 (O_440,N_16130,N_15177);
or UO_441 (O_441,N_19929,N_19116);
and UO_442 (O_442,N_19828,N_15014);
or UO_443 (O_443,N_18054,N_17651);
nand UO_444 (O_444,N_17952,N_18380);
and UO_445 (O_445,N_15376,N_15936);
xor UO_446 (O_446,N_15420,N_15040);
nand UO_447 (O_447,N_16206,N_19480);
nand UO_448 (O_448,N_16092,N_19087);
or UO_449 (O_449,N_16531,N_18609);
or UO_450 (O_450,N_18038,N_18917);
or UO_451 (O_451,N_15593,N_17351);
or UO_452 (O_452,N_15083,N_17950);
or UO_453 (O_453,N_18205,N_17572);
and UO_454 (O_454,N_17357,N_18612);
and UO_455 (O_455,N_16823,N_17677);
nor UO_456 (O_456,N_17286,N_19531);
nor UO_457 (O_457,N_17958,N_17363);
or UO_458 (O_458,N_15187,N_15132);
xor UO_459 (O_459,N_18896,N_18032);
and UO_460 (O_460,N_15407,N_18871);
and UO_461 (O_461,N_19267,N_15572);
or UO_462 (O_462,N_19245,N_17359);
xor UO_463 (O_463,N_19684,N_16963);
nor UO_464 (O_464,N_16656,N_16048);
nor UO_465 (O_465,N_18003,N_17186);
nor UO_466 (O_466,N_19864,N_15469);
or UO_467 (O_467,N_16338,N_15724);
or UO_468 (O_468,N_15564,N_18009);
and UO_469 (O_469,N_17983,N_16730);
nand UO_470 (O_470,N_17133,N_17340);
xor UO_471 (O_471,N_15682,N_18689);
or UO_472 (O_472,N_19583,N_15728);
or UO_473 (O_473,N_19059,N_16500);
nand UO_474 (O_474,N_16817,N_19897);
and UO_475 (O_475,N_16923,N_15233);
and UO_476 (O_476,N_16503,N_17624);
nand UO_477 (O_477,N_18926,N_15297);
and UO_478 (O_478,N_15681,N_16024);
nor UO_479 (O_479,N_15704,N_15257);
and UO_480 (O_480,N_19949,N_19550);
and UO_481 (O_481,N_19011,N_16732);
nand UO_482 (O_482,N_17887,N_16436);
and UO_483 (O_483,N_19203,N_17003);
nand UO_484 (O_484,N_15216,N_15435);
and UO_485 (O_485,N_19430,N_19591);
and UO_486 (O_486,N_18310,N_18626);
or UO_487 (O_487,N_16808,N_17325);
xor UO_488 (O_488,N_16652,N_16741);
nor UO_489 (O_489,N_19253,N_15288);
nand UO_490 (O_490,N_15474,N_18031);
nor UO_491 (O_491,N_17976,N_15589);
nand UO_492 (O_492,N_19112,N_15423);
nand UO_493 (O_493,N_19487,N_16435);
or UO_494 (O_494,N_18237,N_18587);
xnor UO_495 (O_495,N_15234,N_16625);
nor UO_496 (O_496,N_17502,N_15515);
nand UO_497 (O_497,N_17311,N_16608);
or UO_498 (O_498,N_15031,N_17182);
nand UO_499 (O_499,N_18091,N_19484);
or UO_500 (O_500,N_15218,N_16140);
nand UO_501 (O_501,N_15789,N_15960);
or UO_502 (O_502,N_15640,N_15260);
nand UO_503 (O_503,N_16013,N_17160);
and UO_504 (O_504,N_18497,N_16843);
nand UO_505 (O_505,N_18264,N_17439);
xnor UO_506 (O_506,N_17145,N_18060);
nor UO_507 (O_507,N_15561,N_17791);
nor UO_508 (O_508,N_15272,N_19255);
xor UO_509 (O_509,N_18242,N_19396);
and UO_510 (O_510,N_18912,N_18298);
nor UO_511 (O_511,N_15366,N_16882);
nor UO_512 (O_512,N_16366,N_17799);
nor UO_513 (O_513,N_18536,N_16273);
xor UO_514 (O_514,N_15141,N_15698);
or UO_515 (O_515,N_15780,N_16139);
nor UO_516 (O_516,N_18330,N_16644);
and UO_517 (O_517,N_19976,N_18898);
or UO_518 (O_518,N_19715,N_19564);
nand UO_519 (O_519,N_15036,N_18897);
and UO_520 (O_520,N_17391,N_19772);
nand UO_521 (O_521,N_19944,N_15856);
nand UO_522 (O_522,N_15546,N_19227);
nor UO_523 (O_523,N_18136,N_18328);
nand UO_524 (O_524,N_15436,N_18584);
or UO_525 (O_525,N_16989,N_18075);
nand UO_526 (O_526,N_19324,N_17663);
and UO_527 (O_527,N_19774,N_19867);
or UO_528 (O_528,N_17478,N_19221);
nor UO_529 (O_529,N_19387,N_16034);
and UO_530 (O_530,N_15584,N_15532);
xnor UO_531 (O_531,N_19456,N_16996);
nand UO_532 (O_532,N_19803,N_17123);
nor UO_533 (O_533,N_17342,N_17200);
nand UO_534 (O_534,N_15395,N_18843);
nor UO_535 (O_535,N_19718,N_17011);
or UO_536 (O_536,N_19401,N_18705);
nand UO_537 (O_537,N_17963,N_19910);
and UO_538 (O_538,N_15815,N_19152);
nand UO_539 (O_539,N_19202,N_17244);
or UO_540 (O_540,N_17681,N_15481);
xor UO_541 (O_541,N_15020,N_16220);
and UO_542 (O_542,N_16241,N_15937);
and UO_543 (O_543,N_15226,N_15846);
or UO_544 (O_544,N_16854,N_16949);
and UO_545 (O_545,N_16479,N_19452);
nand UO_546 (O_546,N_17022,N_17702);
or UO_547 (O_547,N_19400,N_17957);
or UO_548 (O_548,N_15134,N_18281);
nand UO_549 (O_549,N_18809,N_15348);
nand UO_550 (O_550,N_18460,N_16495);
nand UO_551 (O_551,N_18061,N_18012);
and UO_552 (O_552,N_18289,N_17758);
or UO_553 (O_553,N_16546,N_17190);
or UO_554 (O_554,N_18096,N_16093);
nand UO_555 (O_555,N_16105,N_15508);
xnor UO_556 (O_556,N_19164,N_15890);
and UO_557 (O_557,N_15178,N_17728);
and UO_558 (O_558,N_18810,N_17071);
or UO_559 (O_559,N_16086,N_18749);
and UO_560 (O_560,N_15679,N_19058);
nor UO_561 (O_561,N_16798,N_16064);
nor UO_562 (O_562,N_16232,N_18805);
nor UO_563 (O_563,N_19957,N_17416);
and UO_564 (O_564,N_19482,N_19406);
nor UO_565 (O_565,N_16914,N_16586);
and UO_566 (O_566,N_18105,N_19398);
or UO_567 (O_567,N_18824,N_19952);
or UO_568 (O_568,N_19171,N_19346);
xor UO_569 (O_569,N_16018,N_19447);
and UO_570 (O_570,N_16079,N_17517);
or UO_571 (O_571,N_17282,N_16988);
nor UO_572 (O_572,N_18641,N_16375);
nor UO_573 (O_573,N_15041,N_17619);
nand UO_574 (O_574,N_19453,N_17668);
or UO_575 (O_575,N_16956,N_18688);
nor UO_576 (O_576,N_15763,N_19372);
nor UO_577 (O_577,N_15293,N_16330);
nor UO_578 (O_578,N_19848,N_15511);
and UO_579 (O_579,N_18617,N_19630);
nor UO_580 (O_580,N_16061,N_16189);
and UO_581 (O_581,N_15346,N_17937);
nor UO_582 (O_582,N_17660,N_18545);
or UO_583 (O_583,N_18876,N_17689);
or UO_584 (O_584,N_19434,N_17577);
nor UO_585 (O_585,N_16051,N_17954);
and UO_586 (O_586,N_19727,N_17628);
and UO_587 (O_587,N_19670,N_16289);
and UO_588 (O_588,N_19246,N_19039);
nor UO_589 (O_589,N_18309,N_16188);
nand UO_590 (O_590,N_17655,N_19594);
and UO_591 (O_591,N_18814,N_15916);
nor UO_592 (O_592,N_19182,N_17222);
nand UO_593 (O_593,N_15055,N_17554);
nand UO_594 (O_594,N_18359,N_16244);
xor UO_595 (O_595,N_15343,N_19658);
or UO_596 (O_596,N_18036,N_19414);
nand UO_597 (O_597,N_19927,N_17245);
nand UO_598 (O_598,N_15784,N_18221);
nor UO_599 (O_599,N_17105,N_18686);
and UO_600 (O_600,N_16311,N_16665);
nand UO_601 (O_601,N_19391,N_18698);
nand UO_602 (O_602,N_16176,N_17713);
nand UO_603 (O_603,N_15175,N_15606);
or UO_604 (O_604,N_15742,N_16810);
xnor UO_605 (O_605,N_18624,N_15307);
nand UO_606 (O_606,N_16083,N_17021);
nor UO_607 (O_607,N_15569,N_19468);
nand UO_608 (O_608,N_19502,N_18526);
or UO_609 (O_609,N_15574,N_15570);
nand UO_610 (O_610,N_19614,N_16671);
xor UO_611 (O_611,N_15622,N_16308);
nor UO_612 (O_612,N_15954,N_17005);
nor UO_613 (O_613,N_17012,N_16478);
nand UO_614 (O_614,N_18729,N_17514);
nor UO_615 (O_615,N_16058,N_18355);
or UO_616 (O_616,N_19706,N_16681);
or UO_617 (O_617,N_16772,N_15438);
xor UO_618 (O_618,N_17759,N_18719);
nor UO_619 (O_619,N_19524,N_19632);
xor UO_620 (O_620,N_17153,N_17078);
xnor UO_621 (O_621,N_19975,N_15152);
nand UO_622 (O_622,N_16770,N_19847);
nor UO_623 (O_623,N_16257,N_17725);
xnor UO_624 (O_624,N_19703,N_16440);
nor UO_625 (O_625,N_19102,N_15201);
xor UO_626 (O_626,N_19623,N_15008);
nand UO_627 (O_627,N_17674,N_17922);
xor UO_628 (O_628,N_15951,N_17468);
nand UO_629 (O_629,N_16427,N_19600);
or UO_630 (O_630,N_18740,N_16859);
or UO_631 (O_631,N_17009,N_17829);
or UO_632 (O_632,N_17967,N_18277);
nor UO_633 (O_633,N_18794,N_19330);
and UO_634 (O_634,N_19498,N_17386);
or UO_635 (O_635,N_19789,N_19065);
nand UO_636 (O_636,N_15806,N_15588);
nor UO_637 (O_637,N_17371,N_15820);
nand UO_638 (O_638,N_15316,N_19162);
nor UO_639 (O_639,N_16562,N_19536);
and UO_640 (O_640,N_19288,N_18301);
xor UO_641 (O_641,N_17551,N_18476);
nand UO_642 (O_642,N_19311,N_18176);
nor UO_643 (O_643,N_15167,N_17897);
xor UO_644 (O_644,N_19728,N_19359);
and UO_645 (O_645,N_18971,N_18723);
or UO_646 (O_646,N_17352,N_18797);
or UO_647 (O_647,N_19034,N_16182);
xor UO_648 (O_648,N_17103,N_15380);
nand UO_649 (O_649,N_19050,N_18206);
or UO_650 (O_650,N_18260,N_16489);
xnor UO_651 (O_651,N_18337,N_19682);
and UO_652 (O_652,N_17435,N_16294);
xnor UO_653 (O_653,N_15519,N_17840);
nand UO_654 (O_654,N_17984,N_16276);
or UO_655 (O_655,N_15453,N_18392);
or UO_656 (O_656,N_18944,N_19094);
nor UO_657 (O_657,N_17943,N_17199);
xor UO_658 (O_658,N_16628,N_16438);
nand UO_659 (O_659,N_18540,N_16929);
xnor UO_660 (O_660,N_19587,N_19074);
nand UO_661 (O_661,N_17014,N_17173);
nand UO_662 (O_662,N_16534,N_19791);
nand UO_663 (O_663,N_16237,N_17252);
and UO_664 (O_664,N_17144,N_19109);
or UO_665 (O_665,N_17221,N_17535);
or UO_666 (O_666,N_16098,N_18516);
nand UO_667 (O_667,N_15021,N_17867);
nor UO_668 (O_668,N_19417,N_16765);
or UO_669 (O_669,N_17378,N_19394);
or UO_670 (O_670,N_18180,N_18269);
nor UO_671 (O_671,N_15363,N_18147);
or UO_672 (O_672,N_17803,N_19357);
or UO_673 (O_673,N_17703,N_18590);
xnor UO_674 (O_674,N_16694,N_15670);
nand UO_675 (O_675,N_19390,N_16735);
xnor UO_676 (O_676,N_16922,N_16615);
nand UO_677 (O_677,N_19052,N_18125);
and UO_678 (O_678,N_19538,N_15080);
xor UO_679 (O_679,N_16607,N_15756);
and UO_680 (O_680,N_16459,N_18083);
nor UO_681 (O_681,N_19935,N_18340);
and UO_682 (O_682,N_15871,N_16786);
and UO_683 (O_683,N_18551,N_19123);
and UO_684 (O_684,N_18558,N_18487);
and UO_685 (O_685,N_15224,N_16167);
nor UO_686 (O_686,N_18724,N_17436);
nor UO_687 (O_687,N_16567,N_16851);
or UO_688 (O_688,N_18746,N_17511);
nand UO_689 (O_689,N_16932,N_17885);
xor UO_690 (O_690,N_16637,N_15211);
nand UO_691 (O_691,N_16448,N_17141);
xnor UO_692 (O_692,N_17045,N_15944);
or UO_693 (O_693,N_16497,N_15555);
nor UO_694 (O_694,N_17294,N_18808);
nand UO_695 (O_695,N_15685,N_16950);
xor UO_696 (O_696,N_15123,N_16679);
nand UO_697 (O_697,N_17289,N_16222);
nand UO_698 (O_698,N_17764,N_17422);
nor UO_699 (O_699,N_19069,N_17101);
or UO_700 (O_700,N_18524,N_17929);
nor UO_701 (O_701,N_17694,N_17671);
nand UO_702 (O_702,N_18020,N_16788);
nand UO_703 (O_703,N_16074,N_17034);
nor UO_704 (O_704,N_18412,N_18039);
and UO_705 (O_705,N_18666,N_18847);
or UO_706 (O_706,N_18610,N_16277);
nor UO_707 (O_707,N_19249,N_15671);
and UO_708 (O_708,N_15074,N_18499);
and UO_709 (O_709,N_16133,N_19666);
or UO_710 (O_710,N_15419,N_16286);
nand UO_711 (O_711,N_15057,N_17215);
nand UO_712 (O_712,N_19686,N_15752);
nor UO_713 (O_713,N_16708,N_15690);
xnor UO_714 (O_714,N_16347,N_17927);
nand UO_715 (O_715,N_15480,N_16343);
nand UO_716 (O_716,N_19007,N_18341);
or UO_717 (O_717,N_17766,N_19788);
nor UO_718 (O_718,N_18541,N_17288);
nor UO_719 (O_719,N_17147,N_15186);
nand UO_720 (O_720,N_17318,N_17356);
nand UO_721 (O_721,N_18002,N_16782);
nand UO_722 (O_722,N_18915,N_16210);
and UO_723 (O_723,N_16376,N_19281);
nand UO_724 (O_724,N_16548,N_15245);
nand UO_725 (O_725,N_19903,N_19090);
nor UO_726 (O_726,N_19479,N_16887);
and UO_727 (O_727,N_15783,N_15305);
nor UO_728 (O_728,N_15052,N_16597);
nor UO_729 (O_729,N_16409,N_18461);
nor UO_730 (O_730,N_16114,N_17484);
nor UO_731 (O_731,N_19883,N_17130);
nor UO_732 (O_732,N_17365,N_17195);
and UO_733 (O_733,N_18444,N_18595);
xor UO_734 (O_734,N_15592,N_15853);
nand UO_735 (O_735,N_18168,N_17879);
or UO_736 (O_736,N_17753,N_19769);
or UO_737 (O_737,N_17603,N_16519);
xor UO_738 (O_738,N_19607,N_19921);
nor UO_739 (O_739,N_17269,N_19402);
and UO_740 (O_740,N_19544,N_17156);
nor UO_741 (O_741,N_16506,N_16639);
or UO_742 (O_742,N_18955,N_19442);
and UO_743 (O_743,N_15247,N_16090);
or UO_744 (O_744,N_19854,N_15354);
and UO_745 (O_745,N_17675,N_15892);
and UO_746 (O_746,N_18959,N_16411);
nand UO_747 (O_747,N_18181,N_19525);
xnor UO_748 (O_748,N_19460,N_16439);
and UO_749 (O_749,N_15235,N_16036);
nand UO_750 (O_750,N_16380,N_17933);
and UO_751 (O_751,N_16318,N_15914);
or UO_752 (O_752,N_19884,N_16831);
nand UO_753 (O_753,N_17110,N_17914);
nand UO_754 (O_754,N_18730,N_17025);
nor UO_755 (O_755,N_19445,N_15978);
nand UO_756 (O_756,N_19356,N_17275);
nand UO_757 (O_757,N_18530,N_19882);
nor UO_758 (O_758,N_17634,N_17733);
and UO_759 (O_759,N_16412,N_15328);
and UO_760 (O_760,N_15100,N_19701);
nand UO_761 (O_761,N_17212,N_15568);
nor UO_762 (O_762,N_18818,N_15303);
xnor UO_763 (O_763,N_19266,N_16445);
nor UO_764 (O_764,N_19537,N_19855);
nor UO_765 (O_765,N_18120,N_16846);
nor UO_766 (O_766,N_17509,N_16307);
and UO_767 (O_767,N_16883,N_19470);
and UO_768 (O_768,N_18224,N_16334);
nor UO_769 (O_769,N_15478,N_19341);
nor UO_770 (O_770,N_16604,N_17526);
or UO_771 (O_771,N_17811,N_15198);
and UO_772 (O_772,N_18565,N_15678);
nand UO_773 (O_773,N_19380,N_16952);
xor UO_774 (O_774,N_19003,N_19350);
nand UO_775 (O_775,N_16650,N_16606);
xnor UO_776 (O_776,N_19098,N_18142);
or UO_777 (O_777,N_17508,N_19995);
or UO_778 (O_778,N_15536,N_15387);
or UO_779 (O_779,N_17421,N_16156);
and UO_780 (O_780,N_17006,N_17444);
or UO_781 (O_781,N_19842,N_17964);
nand UO_782 (O_782,N_16110,N_19817);
nor UO_783 (O_783,N_17726,N_19519);
nand UO_784 (O_784,N_17538,N_17507);
xnor UO_785 (O_785,N_18660,N_18870);
or UO_786 (O_786,N_17191,N_17831);
nor UO_787 (O_787,N_17656,N_18367);
nor UO_788 (O_788,N_16377,N_17410);
nand UO_789 (O_789,N_19443,N_19532);
or UO_790 (O_790,N_16456,N_16800);
nand UO_791 (O_791,N_19261,N_16419);
and UO_792 (O_792,N_18542,N_15081);
or UO_793 (O_793,N_15280,N_18980);
nor UO_794 (O_794,N_18452,N_17224);
or UO_795 (O_795,N_16315,N_16928);
nand UO_796 (O_796,N_17661,N_19688);
and UO_797 (O_797,N_17345,N_17106);
nand UO_798 (O_798,N_19527,N_18762);
or UO_799 (O_799,N_19764,N_15759);
or UO_800 (O_800,N_19877,N_17523);
nor UO_801 (O_801,N_16387,N_15802);
and UO_802 (O_802,N_18250,N_19213);
and UO_803 (O_803,N_17402,N_16621);
nand UO_804 (O_804,N_15414,N_17131);
and UO_805 (O_805,N_18665,N_19194);
xor UO_806 (O_806,N_17274,N_19793);
and UO_807 (O_807,N_18011,N_16350);
and UO_808 (O_808,N_16940,N_19889);
and UO_809 (O_809,N_18906,N_19214);
nor UO_810 (O_810,N_18202,N_16775);
nand UO_811 (O_811,N_17134,N_15065);
nor UO_812 (O_812,N_19599,N_17233);
nand UO_813 (O_813,N_15315,N_18504);
nand UO_814 (O_814,N_15733,N_15338);
nor UO_815 (O_815,N_19156,N_17787);
xor UO_816 (O_816,N_15425,N_15762);
nand UO_817 (O_817,N_15882,N_17413);
xor UO_818 (O_818,N_19187,N_18658);
nor UO_819 (O_819,N_15397,N_19763);
nor UO_820 (O_820,N_19180,N_17716);
or UO_821 (O_821,N_19815,N_16547);
and UO_822 (O_822,N_19108,N_17126);
xor UO_823 (O_823,N_18743,N_16924);
or UO_824 (O_824,N_17841,N_16325);
nand UO_825 (O_825,N_19940,N_17171);
and UO_826 (O_826,N_17919,N_17516);
or UO_827 (O_827,N_16159,N_16881);
and UO_828 (O_828,N_15252,N_17210);
or UO_829 (O_829,N_15768,N_19166);
nor UO_830 (O_830,N_18033,N_18097);
nor UO_831 (O_831,N_15618,N_19062);
and UO_832 (O_832,N_16321,N_17835);
nand UO_833 (O_833,N_19045,N_15952);
nor UO_834 (O_834,N_19620,N_18750);
xor UO_835 (O_835,N_17854,N_16364);
or UO_836 (O_836,N_17953,N_17293);
or UO_837 (O_837,N_16095,N_17652);
nand UO_838 (O_838,N_17560,N_16480);
nand UO_839 (O_839,N_17058,N_16069);
nor UO_840 (O_840,N_19709,N_17247);
xnor UO_841 (O_841,N_17745,N_16871);
nor UO_842 (O_842,N_18977,N_18443);
nor UO_843 (O_843,N_17833,N_16475);
and UO_844 (O_844,N_17972,N_16309);
nor UO_845 (O_845,N_16793,N_16368);
or UO_846 (O_846,N_16631,N_19337);
and UO_847 (O_847,N_19243,N_16879);
nand UO_848 (O_848,N_16747,N_19464);
nor UO_849 (O_849,N_17463,N_18368);
nand UO_850 (O_850,N_19810,N_16696);
or UO_851 (O_851,N_15726,N_16312);
nor UO_852 (O_852,N_16638,N_19084);
nand UO_853 (O_853,N_16360,N_19622);
nand UO_854 (O_854,N_17743,N_17747);
or UO_855 (O_855,N_17329,N_19136);
and UO_856 (O_856,N_18566,N_15079);
nor UO_857 (O_857,N_17265,N_16410);
nor UO_858 (O_858,N_18943,N_19560);
nand UO_859 (O_859,N_18781,N_16890);
or UO_860 (O_860,N_17910,N_18303);
nand UO_861 (O_861,N_18270,N_19833);
and UO_862 (O_862,N_15403,N_19660);
or UO_863 (O_863,N_16792,N_19993);
nand UO_864 (O_864,N_16385,N_15959);
and UO_865 (O_865,N_19005,N_15848);
nand UO_866 (O_866,N_15910,N_15694);
xor UO_867 (O_867,N_18715,N_16236);
or UO_868 (O_868,N_16751,N_19723);
and UO_869 (O_869,N_19193,N_18802);
or UO_870 (O_870,N_18139,N_19695);
nor UO_871 (O_871,N_17360,N_15654);
xor UO_872 (O_872,N_18445,N_19189);
nor UO_873 (O_873,N_16524,N_16729);
nand UO_874 (O_874,N_17888,N_19754);
nand UO_875 (O_875,N_17622,N_19145);
xnor UO_876 (O_876,N_18286,N_18044);
nand UO_877 (O_877,N_18021,N_18925);
or UO_878 (O_878,N_16392,N_19200);
nor UO_879 (O_879,N_17960,N_15388);
nand UO_880 (O_880,N_19197,N_17870);
or UO_881 (O_881,N_17292,N_15697);
nor UO_882 (O_882,N_17037,N_17645);
nor UO_883 (O_883,N_16129,N_17163);
and UO_884 (O_884,N_15541,N_19450);
nand UO_885 (O_885,N_17015,N_16509);
and UO_886 (O_886,N_16291,N_18230);
nand UO_887 (O_887,N_16383,N_16875);
nand UO_888 (O_888,N_17172,N_16304);
and UO_889 (O_889,N_18649,N_17380);
or UO_890 (O_890,N_16692,N_16181);
and UO_891 (O_891,N_18027,N_18143);
and UO_892 (O_892,N_18800,N_19458);
or UO_893 (O_893,N_18219,N_18282);
nor UO_894 (O_894,N_16238,N_17248);
and UO_895 (O_895,N_15816,N_15306);
or UO_896 (O_896,N_17541,N_16265);
or UO_897 (O_897,N_19783,N_19984);
or UO_898 (O_898,N_17412,N_19516);
and UO_899 (O_899,N_18485,N_16738);
nor UO_900 (O_900,N_17044,N_18196);
nand UO_901 (O_901,N_17338,N_17842);
nor UO_902 (O_902,N_17081,N_16706);
and UO_903 (O_903,N_17119,N_19641);
or UO_904 (O_904,N_19477,N_19358);
xnor UO_905 (O_905,N_18308,N_16391);
nand UO_906 (O_906,N_15352,N_19128);
nand UO_907 (O_907,N_16687,N_19748);
or UO_908 (O_908,N_18357,N_16168);
nor UO_909 (O_909,N_18911,N_15624);
and UO_910 (O_910,N_15457,N_18582);
or UO_911 (O_911,N_18424,N_15566);
nand UO_912 (O_912,N_16773,N_17223);
xnor UO_913 (O_913,N_16599,N_18267);
xnor UO_914 (O_914,N_19530,N_15289);
or UO_915 (O_915,N_18320,N_16075);
or UO_916 (O_916,N_17179,N_19650);
nand UO_917 (O_917,N_18258,N_18077);
and UO_918 (O_918,N_15492,N_19861);
and UO_919 (O_919,N_19707,N_16790);
or UO_920 (O_920,N_18182,N_18462);
or UO_921 (O_921,N_15007,N_17100);
nor UO_922 (O_922,N_15072,N_17900);
nand UO_923 (O_923,N_15433,N_16869);
xor UO_924 (O_924,N_18791,N_19724);
or UO_925 (O_925,N_19656,N_18722);
or UO_926 (O_926,N_18385,N_16816);
nand UO_927 (O_927,N_18864,N_17613);
or UO_928 (O_928,N_15090,N_19946);
nor UO_929 (O_929,N_18086,N_17988);
or UO_930 (O_930,N_19362,N_16683);
and UO_931 (O_931,N_17684,N_17122);
nor UO_932 (O_932,N_16345,N_19759);
xnor UO_933 (O_933,N_19349,N_17917);
or UO_934 (O_934,N_19765,N_15731);
nor UO_935 (O_935,N_19771,N_19863);
nor UO_936 (O_936,N_17575,N_15999);
nor UO_937 (O_937,N_16655,N_19411);
or UO_938 (O_938,N_18924,N_15653);
and UO_939 (O_939,N_18349,N_19733);
nand UO_940 (O_940,N_16552,N_19153);
or UO_941 (O_941,N_19621,N_18716);
nand UO_942 (O_942,N_18751,N_17734);
nand UO_943 (O_943,N_18447,N_16266);
and UO_944 (O_944,N_16041,N_17491);
xor UO_945 (O_945,N_17367,N_18812);
or UO_946 (O_946,N_16258,N_15751);
nand UO_947 (O_947,N_15985,N_17257);
nand UO_948 (O_948,N_18908,N_17948);
and UO_949 (O_949,N_19612,N_19917);
or UO_950 (O_950,N_16910,N_17041);
or UO_951 (O_951,N_16424,N_17806);
nand UO_952 (O_952,N_18007,N_16322);
nand UO_953 (O_953,N_19644,N_17201);
nand UO_954 (O_954,N_19317,N_19805);
or UO_955 (O_955,N_16272,N_19990);
or UO_956 (O_956,N_19747,N_15077);
or UO_957 (O_957,N_17260,N_17149);
or UO_958 (O_958,N_17404,N_15013);
or UO_959 (O_959,N_17203,N_19685);
or UO_960 (O_960,N_15517,N_16372);
nor UO_961 (O_961,N_15636,N_17534);
and UO_962 (O_962,N_15384,N_16673);
nand UO_963 (O_963,N_19466,N_15980);
nand UO_964 (O_964,N_17774,N_17928);
and UO_965 (O_965,N_18569,N_16152);
or UO_966 (O_966,N_19489,N_19260);
and UO_967 (O_967,N_17168,N_16591);
and UO_968 (O_968,N_16026,N_19132);
nand UO_969 (O_969,N_19675,N_18598);
and UO_970 (O_970,N_18342,N_19091);
or UO_971 (O_971,N_15426,N_17899);
and UO_972 (O_972,N_16042,N_18343);
nand UO_973 (O_973,N_17481,N_17471);
and UO_974 (O_974,N_18235,N_15735);
nand UO_975 (O_975,N_16601,N_15956);
nor UO_976 (O_976,N_18148,N_15585);
nand UO_977 (O_977,N_19160,N_16483);
nor UO_978 (O_978,N_16324,N_18643);
xnor UO_979 (O_979,N_19032,N_17667);
nor UO_980 (O_980,N_17181,N_19139);
nor UO_981 (O_981,N_16259,N_15649);
nor UO_982 (O_982,N_16204,N_16693);
nor UO_983 (O_983,N_18885,N_18493);
nor UO_984 (O_984,N_18605,N_16231);
and UO_985 (O_985,N_18514,N_18535);
nor UO_986 (O_986,N_15617,N_19174);
nor UO_987 (O_987,N_18423,N_18775);
or UO_988 (O_988,N_15109,N_15830);
or UO_989 (O_989,N_16401,N_16402);
or UO_990 (O_990,N_17949,N_19657);
and UO_991 (O_991,N_17707,N_15840);
nand UO_992 (O_992,N_18661,N_16543);
xor UO_993 (O_993,N_19857,N_19021);
and UO_994 (O_994,N_16153,N_15458);
and UO_995 (O_995,N_19782,N_18798);
nor UO_996 (O_996,N_18863,N_15473);
and UO_997 (O_997,N_19843,N_18622);
nor UO_998 (O_998,N_15718,N_16233);
nor UO_999 (O_999,N_16555,N_18842);
and UO_1000 (O_1000,N_18114,N_18599);
nand UO_1001 (O_1001,N_15787,N_16512);
nand UO_1002 (O_1002,N_19635,N_16662);
and UO_1003 (O_1003,N_17569,N_17430);
nand UO_1004 (O_1004,N_18520,N_15965);
or UO_1005 (O_1005,N_17920,N_16718);
nand UO_1006 (O_1006,N_15766,N_19667);
and UO_1007 (O_1007,N_15374,N_15406);
nand UO_1008 (O_1008,N_18271,N_17428);
or UO_1009 (O_1009,N_19597,N_17796);
or UO_1010 (O_1010,N_18987,N_17493);
xor UO_1011 (O_1011,N_15562,N_17872);
nor UO_1012 (O_1012,N_18920,N_19654);
nor UO_1013 (O_1013,N_19588,N_17306);
and UO_1014 (O_1014,N_15842,N_18386);
nand UO_1015 (O_1015,N_19177,N_18874);
nor UO_1016 (O_1016,N_17649,N_17650);
and UO_1017 (O_1017,N_18376,N_18821);
or UO_1018 (O_1018,N_17851,N_17807);
and UO_1019 (O_1019,N_15076,N_16657);
and UO_1020 (O_1020,N_16043,N_18593);
and UO_1021 (O_1021,N_18836,N_16037);
and UO_1022 (O_1022,N_16613,N_18273);
nand UO_1023 (O_1023,N_19473,N_15490);
xor UO_1024 (O_1024,N_17527,N_15669);
xnor UO_1025 (O_1025,N_18496,N_18014);
nor UO_1026 (O_1026,N_18795,N_16820);
nor UO_1027 (O_1027,N_15507,N_16487);
nor UO_1028 (O_1028,N_16261,N_17368);
nand UO_1029 (O_1029,N_17968,N_17059);
and UO_1030 (O_1030,N_15975,N_18792);
nand UO_1031 (O_1031,N_19111,N_16872);
xnor UO_1032 (O_1032,N_19928,N_15440);
nor UO_1033 (O_1033,N_16477,N_17409);
and UO_1034 (O_1034,N_15091,N_17062);
nor UO_1035 (O_1035,N_17065,N_18314);
nor UO_1036 (O_1036,N_17042,N_17616);
nand UO_1037 (O_1037,N_16423,N_19023);
nor UO_1038 (O_1038,N_19931,N_18939);
nor UO_1039 (O_1039,N_15281,N_16096);
and UO_1040 (O_1040,N_15487,N_17095);
and UO_1041 (O_1041,N_15017,N_16327);
nand UO_1042 (O_1042,N_17697,N_17384);
and UO_1043 (O_1043,N_17324,N_18517);
and UO_1044 (O_1044,N_18111,N_19554);
nand UO_1045 (O_1045,N_16942,N_16684);
and UO_1046 (O_1046,N_17985,N_17912);
xnor UO_1047 (O_1047,N_17226,N_19294);
nand UO_1048 (O_1048,N_16060,N_15900);
nand UO_1049 (O_1049,N_19850,N_18546);
and UO_1050 (O_1050,N_19958,N_19602);
and UO_1051 (O_1051,N_17196,N_19566);
or UO_1052 (O_1052,N_17612,N_19201);
nand UO_1053 (O_1053,N_17235,N_18420);
nor UO_1054 (O_1054,N_15184,N_18868);
and UO_1055 (O_1055,N_17556,N_16494);
nand UO_1056 (O_1056,N_17498,N_15822);
nor UO_1057 (O_1057,N_18217,N_18300);
nand UO_1058 (O_1058,N_19490,N_17890);
or UO_1059 (O_1059,N_17328,N_16348);
and UO_1060 (O_1060,N_18910,N_17868);
and UO_1061 (O_1061,N_18439,N_18799);
nand UO_1062 (O_1062,N_18909,N_17091);
and UO_1063 (O_1063,N_18650,N_19953);
nor UO_1064 (O_1064,N_15411,N_18579);
nor UO_1065 (O_1065,N_15935,N_15422);
nor UO_1066 (O_1066,N_17838,N_15194);
nor UO_1067 (O_1067,N_16510,N_15028);
and UO_1068 (O_1068,N_15725,N_16175);
or UO_1069 (O_1069,N_17486,N_17115);
and UO_1070 (O_1070,N_15893,N_17094);
and UO_1071 (O_1071,N_19043,N_17776);
and UO_1072 (O_1072,N_16460,N_18201);
nand UO_1073 (O_1073,N_19325,N_18711);
and UO_1074 (O_1074,N_17376,N_17052);
nand UO_1075 (O_1075,N_16028,N_15987);
or UO_1076 (O_1076,N_19395,N_17361);
or UO_1077 (O_1077,N_19478,N_17170);
or UO_1078 (O_1078,N_16416,N_15042);
and UO_1079 (O_1079,N_16974,N_16118);
and UO_1080 (O_1080,N_18480,N_17849);
or UO_1081 (O_1081,N_15506,N_16455);
or UO_1082 (O_1082,N_16407,N_18316);
and UO_1083 (O_1083,N_17525,N_19129);
nand UO_1084 (O_1084,N_19822,N_19155);
nand UO_1085 (O_1085,N_18458,N_16484);
or UO_1086 (O_1086,N_19720,N_17494);
xor UO_1087 (O_1087,N_17798,N_18056);
nor UO_1088 (O_1088,N_15353,N_15461);
nor UO_1089 (O_1089,N_19936,N_16814);
nor UO_1090 (O_1090,N_16761,N_19408);
or UO_1091 (O_1091,N_16698,N_17771);
nor UO_1092 (O_1092,N_15957,N_19521);
xnor UO_1093 (O_1093,N_17884,N_18327);
nand UO_1094 (O_1094,N_15962,N_17852);
or UO_1095 (O_1095,N_15941,N_19781);
nor UO_1096 (O_1096,N_17971,N_17686);
and UO_1097 (O_1097,N_16071,N_18570);
and UO_1098 (O_1098,N_17466,N_15189);
and UO_1099 (O_1099,N_16857,N_19118);
and UO_1100 (O_1100,N_15120,N_16335);
nor UO_1101 (O_1101,N_18544,N_19712);
xor UO_1102 (O_1102,N_18154,N_15340);
and UO_1103 (O_1103,N_16101,N_15667);
and UO_1104 (O_1104,N_15791,N_17029);
nor UO_1105 (O_1105,N_16504,N_15110);
nor UO_1106 (O_1106,N_17330,N_17157);
and UO_1107 (O_1107,N_15319,N_17858);
and UO_1108 (O_1108,N_16978,N_18663);
or UO_1109 (O_1109,N_17839,N_18062);
xnor UO_1110 (O_1110,N_16825,N_16663);
nor UO_1111 (O_1111,N_17225,N_19355);
or UO_1112 (O_1112,N_18923,N_18465);
or UO_1113 (O_1113,N_15499,N_16473);
nand UO_1114 (O_1114,N_16578,N_17715);
or UO_1115 (O_1115,N_18080,N_17825);
nor UO_1116 (O_1116,N_19653,N_18388);
and UO_1117 (O_1117,N_18004,N_17159);
or UO_1118 (O_1118,N_17621,N_18198);
and UO_1119 (O_1119,N_15415,N_19024);
xor UO_1120 (O_1120,N_15356,N_18589);
and UO_1121 (O_1121,N_15847,N_18268);
nand UO_1122 (O_1122,N_17729,N_17876);
and UO_1123 (O_1123,N_16035,N_15321);
xor UO_1124 (O_1124,N_18262,N_17370);
nand UO_1125 (O_1125,N_19998,N_15510);
nor UO_1126 (O_1126,N_16796,N_18008);
nor UO_1127 (O_1127,N_15580,N_19299);
nand UO_1128 (O_1128,N_16622,N_17820);
or UO_1129 (O_1129,N_16496,N_17940);
nand UO_1130 (O_1130,N_15112,N_18052);
nand UO_1131 (O_1131,N_19811,N_18903);
and UO_1132 (O_1132,N_16838,N_18538);
xnor UO_1133 (O_1133,N_19491,N_18284);
nor UO_1134 (O_1134,N_17889,N_15571);
and UO_1135 (O_1135,N_16297,N_18953);
nand UO_1136 (O_1136,N_17239,N_18266);
nand UO_1137 (O_1137,N_17189,N_18127);
nor UO_1138 (O_1138,N_16063,N_19840);
and UO_1139 (O_1139,N_19121,N_18703);
nor UO_1140 (O_1140,N_17731,N_16771);
nand UO_1141 (O_1141,N_16371,N_17545);
nand UO_1142 (O_1142,N_17180,N_15114);
nor UO_1143 (O_1143,N_17394,N_19731);
nand UO_1144 (O_1144,N_19807,N_18657);
nor UO_1145 (O_1145,N_19878,N_18490);
and UO_1146 (O_1146,N_17565,N_15604);
or UO_1147 (O_1147,N_19496,N_19559);
and UO_1148 (O_1148,N_16934,N_15160);
and UO_1149 (O_1149,N_19006,N_17896);
nand UO_1150 (O_1150,N_16649,N_19514);
and UO_1151 (O_1151,N_15243,N_17877);
xor UO_1152 (O_1152,N_15019,N_19407);
xor UO_1153 (O_1153,N_16102,N_15302);
and UO_1154 (O_1154,N_18905,N_17161);
xnor UO_1155 (O_1155,N_15488,N_15687);
xnor UO_1156 (O_1156,N_17903,N_15455);
nor UO_1157 (O_1157,N_19839,N_16103);
or UO_1158 (O_1158,N_16400,N_19412);
nand UO_1159 (O_1159,N_16527,N_16844);
and UO_1160 (O_1160,N_19019,N_16664);
xnor UO_1161 (O_1161,N_17755,N_17544);
or UO_1162 (O_1162,N_17735,N_15116);
nor UO_1163 (O_1163,N_16623,N_17117);
nor UO_1164 (O_1164,N_19378,N_17802);
and UO_1165 (O_1165,N_19639,N_17198);
and UO_1166 (O_1166,N_16629,N_17185);
nor UO_1167 (O_1167,N_15324,N_17558);
and UO_1168 (O_1168,N_19590,N_18140);
and UO_1169 (O_1169,N_18922,N_18642);
or UO_1170 (O_1170,N_17407,N_19105);
xor UO_1171 (O_1171,N_19106,N_15044);
xor UO_1172 (O_1172,N_15093,N_17947);
and UO_1173 (O_1173,N_15327,N_19974);
xnor UO_1174 (O_1174,N_17267,N_16250);
or UO_1175 (O_1175,N_18759,N_17477);
or UO_1176 (O_1176,N_18913,N_17089);
xnor UO_1177 (O_1177,N_17869,N_16542);
and UO_1178 (O_1178,N_16164,N_16653);
or UO_1179 (O_1179,N_19925,N_18213);
nand UO_1180 (O_1180,N_15730,N_16365);
and UO_1181 (O_1181,N_16902,N_17087);
nand UO_1182 (O_1182,N_18849,N_16697);
nand UO_1183 (O_1183,N_16328,N_16986);
nand UO_1184 (O_1184,N_18350,N_19354);
nor UO_1185 (O_1185,N_15646,N_15067);
nor UO_1186 (O_1186,N_18025,N_18410);
xor UO_1187 (O_1187,N_19493,N_15919);
and UO_1188 (O_1188,N_15734,N_16239);
nand UO_1189 (O_1189,N_19880,N_18534);
xor UO_1190 (O_1190,N_19673,N_18754);
or UO_1191 (O_1191,N_19083,N_18928);
nand UO_1192 (O_1192,N_19418,N_17232);
nor UO_1193 (O_1193,N_16767,N_16403);
or UO_1194 (O_1194,N_16271,N_16997);
xnor UO_1195 (O_1195,N_15259,N_16818);
nor UO_1196 (O_1196,N_15220,N_19608);
or UO_1197 (O_1197,N_18638,N_19541);
and UO_1198 (O_1198,N_17373,N_16044);
and UO_1199 (O_1199,N_18518,N_16784);
nand UO_1200 (O_1200,N_15695,N_16170);
and UO_1201 (O_1201,N_18628,N_15249);
nor UO_1202 (O_1202,N_16841,N_17271);
or UO_1203 (O_1203,N_18228,N_18398);
and UO_1204 (O_1204,N_18047,N_18664);
xor UO_1205 (O_1205,N_18107,N_18291);
xnor UO_1206 (O_1206,N_15819,N_19892);
and UO_1207 (O_1207,N_15049,N_16449);
or UO_1208 (O_1208,N_16794,N_18539);
nor UO_1209 (O_1209,N_15450,N_18064);
nand UO_1210 (O_1210,N_18331,N_18203);
and UO_1211 (O_1211,N_18429,N_16865);
nor UO_1212 (O_1212,N_15291,N_16299);
nor UO_1213 (O_1213,N_19528,N_18513);
and UO_1214 (O_1214,N_16201,N_16845);
and UO_1215 (O_1215,N_18756,N_19263);
nor UO_1216 (O_1216,N_15210,N_18616);
or UO_1217 (O_1217,N_17871,N_16743);
nor UO_1218 (O_1218,N_17426,N_18005);
and UO_1219 (O_1219,N_16594,N_15899);
nand UO_1220 (O_1220,N_18725,N_17601);
nor UO_1221 (O_1221,N_15800,N_16565);
nor UO_1222 (O_1222,N_18194,N_15709);
xor UO_1223 (O_1223,N_19381,N_17326);
or UO_1224 (O_1224,N_18969,N_18537);
xor UO_1225 (O_1225,N_17701,N_18467);
nor UO_1226 (O_1226,N_15927,N_15788);
nand UO_1227 (O_1227,N_15005,N_16884);
and UO_1228 (O_1228,N_15792,N_15313);
nand UO_1229 (O_1229,N_19455,N_19584);
and UO_1230 (O_1230,N_18783,N_19292);
or UO_1231 (O_1231,N_18257,N_18853);
nand UO_1232 (O_1232,N_19837,N_18115);
and UO_1233 (O_1233,N_17447,N_15113);
nor UO_1234 (O_1234,N_19799,N_16355);
nor UO_1235 (O_1235,N_15368,N_15683);
nand UO_1236 (O_1236,N_19708,N_15696);
and UO_1237 (O_1237,N_18124,N_18778);
and UO_1238 (O_1238,N_19421,N_19095);
or UO_1239 (O_1239,N_19939,N_18141);
nand UO_1240 (O_1240,N_18581,N_16161);
or UO_1241 (O_1241,N_15576,N_19425);
or UO_1242 (O_1242,N_17510,N_19282);
nand UO_1243 (O_1243,N_18656,N_16876);
and UO_1244 (O_1244,N_19101,N_18436);
nor UO_1245 (O_1245,N_18942,N_15777);
and UO_1246 (O_1246,N_15638,N_16661);
nand UO_1247 (O_1247,N_17615,N_19092);
or UO_1248 (O_1248,N_18933,N_15317);
or UO_1249 (O_1249,N_19693,N_19919);
nand UO_1250 (O_1250,N_18878,N_17213);
nand UO_1251 (O_1251,N_15867,N_16791);
xor UO_1252 (O_1252,N_15375,N_17040);
or UO_1253 (O_1253,N_18360,N_16959);
and UO_1254 (O_1254,N_17125,N_18498);
xnor UO_1255 (O_1255,N_18448,N_15809);
nand UO_1256 (O_1256,N_16651,N_15326);
nor UO_1257 (O_1257,N_18623,N_16326);
or UO_1258 (O_1258,N_16186,N_16354);
and UO_1259 (O_1259,N_16758,N_18620);
and UO_1260 (O_1260,N_19028,N_16163);
nor UO_1261 (O_1261,N_16764,N_16388);
nor UO_1262 (O_1262,N_15970,N_18351);
nand UO_1263 (O_1263,N_19700,N_18197);
nand UO_1264 (O_1264,N_15673,N_19321);
and UO_1265 (O_1265,N_16180,N_19996);
xor UO_1266 (O_1266,N_18956,N_15885);
and UO_1267 (O_1267,N_18373,N_19298);
nor UO_1268 (O_1268,N_17859,N_18104);
or UO_1269 (O_1269,N_17591,N_15117);
nand UO_1270 (O_1270,N_17148,N_15535);
and UO_1271 (O_1271,N_17658,N_15563);
and UO_1272 (O_1272,N_16829,N_16172);
xnor UO_1273 (O_1273,N_17643,N_18681);
and UO_1274 (O_1274,N_17862,N_19951);
nor UO_1275 (O_1275,N_15012,N_15159);
xnor UO_1276 (O_1276,N_18117,N_17129);
or UO_1277 (O_1277,N_19859,N_18881);
and UO_1278 (O_1278,N_16873,N_17638);
and UO_1279 (O_1279,N_15102,N_18067);
nor UO_1280 (O_1280,N_19247,N_18153);
and UO_1281 (O_1281,N_16561,N_16850);
or UO_1282 (O_1282,N_17738,N_16040);
and UO_1283 (O_1283,N_17706,N_19376);
and UO_1284 (O_1284,N_17067,N_17227);
or UO_1285 (O_1285,N_18240,N_19097);
and UO_1286 (O_1286,N_18929,N_18640);
nor UO_1287 (O_1287,N_15292,N_16121);
nor UO_1288 (O_1288,N_15274,N_19888);
or UO_1289 (O_1289,N_18998,N_17298);
or UO_1290 (O_1290,N_18755,N_16536);
xor UO_1291 (O_1291,N_16905,N_17349);
xor UO_1292 (O_1292,N_17035,N_18564);
or UO_1293 (O_1293,N_18830,N_18945);
nand UO_1294 (O_1294,N_19481,N_16080);
nand UO_1295 (O_1295,N_18886,N_15608);
and UO_1296 (O_1296,N_16867,N_19971);
and UO_1297 (O_1297,N_18050,N_15794);
nand UO_1298 (O_1298,N_16088,N_16915);
xnor UO_1299 (O_1299,N_15412,N_19262);
xnor UO_1300 (O_1300,N_18455,N_16891);
and UO_1301 (O_1301,N_15886,N_18431);
nand UO_1302 (O_1302,N_15413,N_19978);
nand UO_1303 (O_1303,N_15736,N_18844);
or UO_1304 (O_1304,N_19896,N_18022);
nand UO_1305 (O_1305,N_15335,N_19662);
nor UO_1306 (O_1306,N_15129,N_15711);
nor UO_1307 (O_1307,N_16744,N_18079);
nand UO_1308 (O_1308,N_15334,N_19633);
nand UO_1309 (O_1309,N_17557,N_18784);
and UO_1310 (O_1310,N_17936,N_19619);
and UO_1311 (O_1311,N_18771,N_18651);
nor UO_1312 (O_1312,N_15865,N_19148);
nor UO_1313 (O_1313,N_15656,N_16980);
nand UO_1314 (O_1314,N_16550,N_17169);
and UO_1315 (O_1315,N_16055,N_18613);
nor UO_1316 (O_1316,N_18529,N_18984);
or UO_1317 (O_1317,N_19740,N_16196);
nand UO_1318 (O_1318,N_18687,N_15330);
nor UO_1319 (O_1319,N_19821,N_18608);
or UO_1320 (O_1320,N_15075,N_19841);
nand UO_1321 (O_1321,N_18507,N_15158);
nand UO_1322 (O_1322,N_18294,N_17696);
and UO_1323 (O_1323,N_15632,N_17127);
nor UO_1324 (O_1324,N_15208,N_17390);
and UO_1325 (O_1325,N_18803,N_16749);
and UO_1326 (O_1326,N_16654,N_18968);
xor UO_1327 (O_1327,N_18365,N_17299);
nand UO_1328 (O_1328,N_15174,N_17909);
and UO_1329 (O_1329,N_19440,N_16493);
or UO_1330 (O_1330,N_15027,N_18521);
or UO_1331 (O_1331,N_19038,N_17873);
or UO_1332 (O_1332,N_17784,N_17283);
nor UO_1333 (O_1333,N_16957,N_15738);
nand UO_1334 (O_1334,N_16563,N_19968);
nand UO_1335 (O_1335,N_17374,N_15655);
nor UO_1336 (O_1336,N_17679,N_15998);
and UO_1337 (O_1337,N_18274,N_19750);
nor UO_1338 (O_1338,N_18963,N_19862);
or UO_1339 (O_1339,N_17767,N_19191);
nor UO_1340 (O_1340,N_15205,N_15786);
nand UO_1341 (O_1341,N_19269,N_16700);
xor UO_1342 (O_1342,N_15255,N_17464);
and UO_1343 (O_1343,N_17866,N_18748);
nand UO_1344 (O_1344,N_18840,N_15046);
or UO_1345 (O_1345,N_15396,N_15909);
nand UO_1346 (O_1346,N_16027,N_15432);
or UO_1347 (O_1347,N_18949,N_19879);
or UO_1348 (O_1348,N_18072,N_16421);
and UO_1349 (O_1349,N_16263,N_15881);
xor UO_1350 (O_1350,N_16645,N_15092);
or UO_1351 (O_1351,N_17111,N_19824);
nor UO_1352 (O_1352,N_18832,N_15598);
nor UO_1353 (O_1353,N_17780,N_15858);
and UO_1354 (O_1354,N_15992,N_16962);
or UO_1355 (O_1355,N_19051,N_15776);
or UO_1356 (O_1356,N_18193,N_19924);
nor UO_1357 (O_1357,N_16282,N_17680);
nor UO_1358 (O_1358,N_16278,N_18647);
and UO_1359 (O_1359,N_17857,N_17902);
nor UO_1360 (O_1360,N_16057,N_19190);
xnor UO_1361 (O_1361,N_15855,N_19424);
or UO_1362 (O_1362,N_17678,N_17809);
xor UO_1363 (O_1363,N_17445,N_17382);
or UO_1364 (O_1364,N_18470,N_16685);
or UO_1365 (O_1365,N_17433,N_16822);
or UO_1366 (O_1366,N_18409,N_15526);
and UO_1367 (O_1367,N_19500,N_15190);
nor UO_1368 (O_1368,N_18231,N_15261);
and UO_1369 (O_1369,N_16109,N_16642);
and UO_1370 (O_1370,N_18673,N_16429);
nor UO_1371 (O_1371,N_17385,N_17055);
nor UO_1372 (O_1372,N_16672,N_18850);
or UO_1373 (O_1373,N_16931,N_19437);
or UO_1374 (O_1374,N_15880,N_19595);
nor UO_1375 (O_1375,N_16954,N_15953);
and UO_1376 (O_1376,N_15525,N_16995);
xor UO_1377 (O_1377,N_16019,N_18378);
or UO_1378 (O_1378,N_19800,N_16624);
nor UO_1379 (O_1379,N_17580,N_19042);
or UO_1380 (O_1380,N_16864,N_19252);
nor UO_1381 (O_1381,N_17797,N_16926);
or UO_1382 (O_1382,N_19250,N_18994);
nor UO_1383 (O_1383,N_19025,N_15308);
or UO_1384 (O_1384,N_17327,N_19582);
nand UO_1385 (O_1385,N_16230,N_16418);
and UO_1386 (O_1386,N_19120,N_17605);
and UO_1387 (O_1387,N_16856,N_19219);
and UO_1388 (O_1388,N_15135,N_18889);
or UO_1389 (O_1389,N_19784,N_16246);
and UO_1390 (O_1390,N_16886,N_18028);
nor UO_1391 (O_1391,N_16596,N_19336);
nor UO_1392 (O_1392,N_19994,N_16558);
nand UO_1393 (O_1393,N_18272,N_15239);
nand UO_1394 (O_1394,N_18951,N_17403);
or UO_1395 (O_1395,N_16339,N_15472);
or UO_1396 (O_1396,N_15339,N_18854);
and UO_1397 (O_1397,N_17709,N_19439);
nand UO_1398 (O_1398,N_19808,N_15225);
nor UO_1399 (O_1399,N_18879,N_17895);
or UO_1400 (O_1400,N_15361,N_18451);
nor UO_1401 (O_1401,N_18207,N_19548);
or UO_1402 (O_1402,N_17585,N_18276);
or UO_1403 (O_1403,N_19699,N_17682);
and UO_1404 (O_1404,N_16249,N_19648);
or UO_1405 (O_1405,N_19117,N_19022);
xor UO_1406 (O_1406,N_18051,N_16824);
nand UO_1407 (O_1407,N_18654,N_16126);
nor UO_1408 (O_1408,N_18259,N_15605);
nor UO_1409 (O_1409,N_17856,N_15251);
xnor UO_1410 (O_1410,N_19901,N_17450);
nor UO_1411 (O_1411,N_15868,N_15398);
and UO_1412 (O_1412,N_16763,N_15500);
nor UO_1413 (O_1413,N_15753,N_18063);
and UO_1414 (O_1414,N_18466,N_17827);
and UO_1415 (O_1415,N_18573,N_19852);
nand UO_1416 (O_1416,N_15130,N_19529);
nand UO_1417 (O_1417,N_18975,N_19567);
nor UO_1418 (O_1418,N_16006,N_19419);
nor UO_1419 (O_1419,N_16635,N_15263);
and UO_1420 (O_1420,N_19651,N_18636);
nor UO_1421 (O_1421,N_15619,N_16077);
nor UO_1422 (O_1422,N_18576,N_15599);
nor UO_1423 (O_1423,N_15513,N_15048);
xnor UO_1424 (O_1424,N_19829,N_18921);
nor UO_1425 (O_1425,N_16144,N_18399);
xor UO_1426 (O_1426,N_17092,N_17837);
nand UO_1427 (O_1427,N_19141,N_16975);
nand UO_1428 (O_1428,N_16589,N_15680);
nor UO_1429 (O_1429,N_19389,N_15591);
nand UO_1430 (O_1430,N_18757,N_18046);
nand UO_1431 (O_1431,N_15342,N_19423);
nand UO_1432 (O_1432,N_15275,N_17875);
and UO_1433 (O_1433,N_18988,N_17752);
nand UO_1434 (O_1434,N_17568,N_19849);
xnor UO_1435 (O_1435,N_16731,N_15294);
xor UO_1436 (O_1436,N_15086,N_15273);
or UO_1437 (O_1437,N_19149,N_15930);
and UO_1438 (O_1438,N_18631,N_17962);
and UO_1439 (O_1439,N_19905,N_16003);
nand UO_1440 (O_1440,N_18209,N_19825);
nor UO_1441 (O_1441,N_15637,N_16157);
or UO_1442 (O_1442,N_17068,N_18835);
xnor UO_1443 (O_1443,N_19671,N_17425);
or UO_1444 (O_1444,N_16960,N_16953);
and UO_1445 (O_1445,N_19716,N_17060);
nor UO_1446 (O_1446,N_18468,N_17432);
or UO_1447 (O_1447,N_17443,N_18891);
xor UO_1448 (O_1448,N_17174,N_17398);
and UO_1449 (O_1449,N_18965,N_19004);
nand UO_1450 (O_1450,N_18362,N_16200);
xor UO_1451 (O_1451,N_19374,N_15859);
nand UO_1452 (O_1452,N_15401,N_18600);
nor UO_1453 (O_1453,N_15202,N_17155);
nor UO_1454 (O_1454,N_15296,N_18873);
and UO_1455 (O_1455,N_19366,N_18162);
nand UO_1456 (O_1456,N_19284,N_16283);
nand UO_1457 (O_1457,N_18954,N_16351);
and UO_1458 (O_1458,N_16690,N_16603);
nand UO_1459 (O_1459,N_19534,N_16617);
and UO_1460 (O_1460,N_16267,N_18717);
or UO_1461 (O_1461,N_17165,N_15601);
or UO_1462 (O_1462,N_16212,N_18381);
nand UO_1463 (O_1463,N_15538,N_17462);
nor UO_1464 (O_1464,N_16847,N_17030);
nor UO_1465 (O_1465,N_17090,N_16930);
nor UO_1466 (O_1466,N_19475,N_19242);
nor UO_1467 (O_1467,N_17177,N_15955);
nor UO_1468 (O_1468,N_16911,N_16526);
nor UO_1469 (O_1469,N_15381,N_16162);
xor UO_1470 (O_1470,N_16073,N_16537);
and UO_1471 (O_1471,N_17383,N_17801);
nor UO_1472 (O_1472,N_17242,N_17151);
and UO_1473 (O_1473,N_16135,N_18137);
nand UO_1474 (O_1474,N_16049,N_19057);
or UO_1475 (O_1475,N_19730,N_15720);
or UO_1476 (O_1476,N_19089,N_17080);
nand UO_1477 (O_1477,N_16205,N_19199);
and UO_1478 (O_1478,N_17547,N_15331);
or UO_1479 (O_1479,N_19040,N_16059);
xnor UO_1480 (O_1480,N_19645,N_18204);
and UO_1481 (O_1481,N_18408,N_17038);
and UO_1482 (O_1482,N_17880,N_15447);
nand UO_1483 (O_1483,N_17941,N_16585);
or UO_1484 (O_1484,N_18761,N_17673);
and UO_1485 (O_1485,N_19937,N_17710);
or UO_1486 (O_1486,N_18680,N_18229);
nor UO_1487 (O_1487,N_18108,N_18183);
nor UO_1488 (O_1488,N_16813,N_19866);
nand UO_1489 (O_1489,N_15144,N_16032);
nand UO_1490 (O_1490,N_16752,N_16115);
or UO_1491 (O_1491,N_19273,N_16217);
and UO_1492 (O_1492,N_18432,N_16406);
or UO_1493 (O_1493,N_15540,N_19158);
or UO_1494 (O_1494,N_15520,N_16305);
or UO_1495 (O_1495,N_15760,N_15121);
or UO_1496 (O_1496,N_18348,N_17828);
nor UO_1497 (O_1497,N_15025,N_15727);
and UO_1498 (O_1498,N_16785,N_16670);
or UO_1499 (O_1499,N_17956,N_16579);
nand UO_1500 (O_1500,N_15105,N_17901);
or UO_1501 (O_1501,N_17736,N_15085);
or UO_1502 (O_1502,N_17723,N_17886);
nor UO_1503 (O_1503,N_16474,N_17489);
nor UO_1504 (O_1504,N_19543,N_17137);
and UO_1505 (O_1505,N_19786,N_16016);
and UO_1506 (O_1506,N_19661,N_19015);
nand UO_1507 (O_1507,N_17978,N_17980);
or UO_1508 (O_1508,N_15051,N_18442);
and UO_1509 (O_1509,N_16505,N_15807);
nor UO_1510 (O_1510,N_19167,N_16577);
or UO_1511 (O_1511,N_16498,N_18978);
nor UO_1512 (O_1512,N_17594,N_16463);
nand UO_1513 (O_1513,N_18774,N_15232);
or UO_1514 (O_1514,N_16268,N_19382);
nand UO_1515 (O_1515,N_17911,N_17050);
and UO_1516 (O_1516,N_17302,N_15262);
or UO_1517 (O_1517,N_15495,N_19306);
or UO_1518 (O_1518,N_16112,N_15824);
or UO_1519 (O_1519,N_15188,N_16695);
nor UO_1520 (O_1520,N_18172,N_19649);
and UO_1521 (O_1521,N_15767,N_16287);
nor UO_1522 (O_1522,N_17749,N_17646);
nand UO_1523 (O_1523,N_16889,N_15552);
or UO_1524 (O_1524,N_16207,N_18065);
or UO_1525 (O_1525,N_15082,N_16104);
nor UO_1526 (O_1526,N_16588,N_18389);
nor UO_1527 (O_1527,N_19792,N_17865);
nor UO_1528 (O_1528,N_17317,N_18819);
xor UO_1529 (O_1529,N_18869,N_15668);
nor UO_1530 (O_1530,N_19302,N_19485);
xor UO_1531 (O_1531,N_18248,N_18094);
or UO_1532 (O_1532,N_16826,N_19031);
or UO_1533 (O_1533,N_18706,N_15118);
xor UO_1534 (O_1534,N_18553,N_18662);
and UO_1535 (O_1535,N_19206,N_19679);
nor UO_1536 (O_1536,N_18862,N_19037);
or UO_1537 (O_1537,N_16755,N_15534);
and UO_1538 (O_1538,N_15922,N_15180);
xor UO_1539 (O_1539,N_19360,N_17763);
nand UO_1540 (O_1540,N_19297,N_15740);
nor UO_1541 (O_1541,N_15195,N_19122);
nor UO_1542 (O_1542,N_17691,N_16762);
nor UO_1543 (O_1543,N_18747,N_15950);
nor UO_1544 (O_1544,N_17064,N_16866);
xor UO_1545 (O_1545,N_17586,N_19345);
nor UO_1546 (O_1546,N_15839,N_19871);
xnor UO_1547 (O_1547,N_19601,N_16107);
nor UO_1548 (O_1548,N_16120,N_15917);
xnor UO_1549 (O_1549,N_16227,N_18179);
or UO_1550 (O_1550,N_16707,N_18116);
nor UO_1551 (O_1551,N_15906,N_17132);
and UO_1552 (O_1552,N_18160,N_18322);
and UO_1553 (O_1553,N_15096,N_17399);
or UO_1554 (O_1554,N_17276,N_15901);
nor UO_1555 (O_1555,N_17354,N_17934);
and UO_1556 (O_1556,N_15778,N_18793);
and UO_1557 (O_1557,N_19721,N_16680);
nand UO_1558 (O_1558,N_15437,N_19875);
or UO_1559 (O_1559,N_17812,N_17188);
nand UO_1560 (O_1560,N_17441,N_19908);
nor UO_1561 (O_1561,N_16193,N_15227);
nand UO_1562 (O_1562,N_18174,N_15634);
nand UO_1563 (O_1563,N_16802,N_17253);
or UO_1564 (O_1564,N_18101,N_19326);
nor UO_1565 (O_1565,N_16750,N_17501);
nand UO_1566 (O_1566,N_17695,N_17031);
nand UO_1567 (O_1567,N_18627,N_18684);
and UO_1568 (O_1568,N_18735,N_15170);
nand UO_1569 (O_1569,N_18138,N_16446);
and UO_1570 (O_1570,N_17264,N_16317);
or UO_1571 (O_1571,N_18280,N_15545);
or UO_1572 (O_1572,N_18133,N_15716);
or UO_1573 (O_1573,N_18682,N_19540);
nand UO_1574 (O_1574,N_17623,N_16630);
nor UO_1575 (O_1575,N_17537,N_16852);
nand UO_1576 (O_1576,N_17026,N_19397);
and UO_1577 (O_1577,N_19895,N_19150);
nand UO_1578 (O_1578,N_18948,N_18811);
nor UO_1579 (O_1579,N_16426,N_15651);
or UO_1580 (O_1580,N_15237,N_15477);
or UO_1581 (O_1581,N_16316,N_16781);
and UO_1582 (O_1582,N_18728,N_15241);
xor UO_1583 (O_1583,N_16465,N_17355);
nor UO_1584 (O_1584,N_15400,N_15248);
or UO_1585 (O_1585,N_15717,N_19234);
nor UO_1586 (O_1586,N_16468,N_18024);
nor UO_1587 (O_1587,N_16699,N_19868);
nand UO_1588 (O_1588,N_16564,N_19874);
and UO_1589 (O_1589,N_15026,N_19449);
or UO_1590 (O_1590,N_18549,N_16290);
or UO_1591 (O_1591,N_15587,N_17108);
and UO_1592 (O_1592,N_18249,N_16434);
and UO_1593 (O_1593,N_18936,N_17821);
nand UO_1594 (O_1594,N_16554,N_15267);
and UO_1595 (O_1595,N_16264,N_16123);
nand UO_1596 (O_1596,N_17659,N_18254);
nor UO_1597 (O_1597,N_18712,N_18678);
or UO_1598 (O_1598,N_15544,N_19176);
or UO_1599 (O_1599,N_16361,N_18126);
nor UO_1600 (O_1600,N_15242,N_19295);
xor UO_1601 (O_1601,N_15009,N_15877);
nor UO_1602 (O_1602,N_16357,N_18406);
xor UO_1603 (O_1603,N_19969,N_19002);
nor UO_1604 (O_1604,N_17732,N_15661);
and UO_1605 (O_1605,N_15537,N_16444);
nand UO_1606 (O_1606,N_16066,N_17046);
or UO_1607 (O_1607,N_17939,N_16119);
or UO_1608 (O_1608,N_19691,N_17506);
xor UO_1609 (O_1609,N_19499,N_16855);
nand UO_1610 (O_1610,N_18326,N_18256);
nor UO_1611 (O_1611,N_17855,N_16242);
nor UO_1612 (O_1612,N_17314,N_18974);
and UO_1613 (O_1613,N_15456,N_19476);
and UO_1614 (O_1614,N_15391,N_17013);
and UO_1615 (O_1615,N_19444,N_19640);
or UO_1616 (O_1616,N_19240,N_19845);
or UO_1617 (O_1617,N_16669,N_16374);
xnor UO_1618 (O_1618,N_17614,N_19441);
and UO_1619 (O_1619,N_15692,N_17805);
or UO_1620 (O_1620,N_17818,N_17595);
nor UO_1621 (O_1621,N_18416,N_19742);
and UO_1622 (O_1622,N_16904,N_19054);
or UO_1623 (O_1623,N_15464,N_19853);
nand UO_1624 (O_1624,N_16522,N_17353);
or UO_1625 (O_1625,N_15265,N_18675);
and UO_1626 (O_1626,N_16284,N_18713);
nand UO_1627 (O_1627,N_16116,N_15016);
nand UO_1628 (O_1628,N_19472,N_17966);
and UO_1629 (O_1629,N_15866,N_16378);
nor UO_1630 (O_1630,N_16877,N_15850);
nand UO_1631 (O_1631,N_17576,N_19231);
or UO_1632 (O_1632,N_16938,N_16215);
and UO_1633 (O_1633,N_19347,N_19233);
and UO_1634 (O_1634,N_16275,N_15104);
or UO_1635 (O_1635,N_16610,N_18095);
nor UO_1636 (O_1636,N_16031,N_19987);
or UO_1637 (O_1637,N_19628,N_15551);
nand UO_1638 (O_1638,N_19547,N_18677);
and UO_1639 (O_1639,N_15761,N_15460);
and UO_1640 (O_1640,N_18404,N_15115);
and UO_1641 (O_1641,N_19436,N_16087);
or UO_1642 (O_1642,N_15614,N_15558);
xor UO_1643 (O_1643,N_15578,N_18395);
nor UO_1644 (O_1644,N_18916,N_18946);
or UO_1645 (O_1645,N_16052,N_15547);
nand UO_1646 (O_1646,N_19506,N_15672);
nor UO_1647 (O_1647,N_15192,N_18296);
and UO_1648 (O_1648,N_16806,N_18092);
and UO_1649 (O_1649,N_16916,N_16417);
or UO_1650 (O_1650,N_17848,N_18192);
xor UO_1651 (O_1651,N_17892,N_17070);
or UO_1652 (O_1652,N_15030,N_18721);
or UO_1653 (O_1653,N_15860,N_19290);
and UO_1654 (O_1654,N_19624,N_16507);
and UO_1655 (O_1655,N_16668,N_17414);
xor UO_1656 (O_1656,N_19539,N_19008);
or UO_1657 (O_1657,N_18492,N_16010);
and UO_1658 (O_1658,N_19030,N_19942);
or UO_1659 (O_1659,N_15639,N_18070);
nor UO_1660 (O_1660,N_16769,N_17424);
nand UO_1661 (O_1661,N_18621,N_18575);
or UO_1662 (O_1662,N_19744,N_19409);
nand UO_1663 (O_1663,N_16279,N_17287);
xnor UO_1664 (O_1664,N_17861,N_17142);
nor UO_1665 (O_1665,N_17297,N_17926);
nor UO_1666 (O_1666,N_16314,N_19488);
and UO_1667 (O_1667,N_16863,N_16783);
nor UO_1668 (O_1668,N_17474,N_17211);
xor UO_1669 (O_1669,N_19448,N_18430);
xor UO_1670 (O_1670,N_19991,N_16815);
and UO_1671 (O_1671,N_18134,N_19669);
nand UO_1672 (O_1672,N_19618,N_18674);
nand UO_1673 (O_1673,N_16616,N_17597);
nand UO_1674 (O_1674,N_18901,N_18446);
nor UO_1675 (O_1675,N_19161,N_19711);
and UO_1676 (O_1676,N_17496,N_18966);
and UO_1677 (O_1677,N_16209,N_18941);
nand UO_1678 (O_1678,N_17308,N_19373);
nor UO_1679 (O_1679,N_16053,N_16643);
and UO_1680 (O_1680,N_15199,N_15684);
and UO_1681 (O_1681,N_17152,N_16686);
nor UO_1682 (O_1682,N_16832,N_18123);
and UO_1683 (O_1683,N_19698,N_17146);
and UO_1684 (O_1684,N_19375,N_18855);
and UO_1685 (O_1685,N_17815,N_19416);
xor UO_1686 (O_1686,N_17418,N_15139);
or UO_1687 (O_1687,N_15050,N_19053);
nor UO_1688 (O_1688,N_19710,N_16070);
nand UO_1689 (O_1689,N_18315,N_16789);
and UO_1690 (O_1690,N_17574,N_18150);
or UO_1691 (O_1691,N_16390,N_18278);
xnor UO_1692 (O_1692,N_17777,N_18779);
nand UO_1693 (O_1693,N_19329,N_19338);
nor UO_1694 (O_1694,N_15064,N_15409);
or UO_1695 (O_1695,N_19127,N_15878);
nand UO_1696 (O_1696,N_17754,N_15207);
xnor UO_1697 (O_1697,N_15677,N_17606);
nor UO_1698 (O_1698,N_18592,N_17760);
nor UO_1699 (O_1699,N_15702,N_19264);
or UO_1700 (O_1700,N_19736,N_16571);
nor UO_1701 (O_1701,N_15814,N_15058);
and UO_1702 (O_1702,N_18606,N_19713);
nor UO_1703 (O_1703,N_15905,N_15688);
and UO_1704 (O_1704,N_17563,N_18428);
nand UO_1705 (O_1705,N_15185,N_15310);
nor UO_1706 (O_1706,N_15896,N_17124);
or UO_1707 (O_1707,N_15056,N_15902);
nor UO_1708 (O_1708,N_18964,N_17688);
nor UO_1709 (O_1709,N_15994,N_15773);
nor UO_1710 (O_1710,N_19368,N_15947);
nor UO_1711 (O_1711,N_15125,N_18034);
nand UO_1712 (O_1712,N_15466,N_18615);
xnor UO_1713 (O_1713,N_19220,N_19766);
or UO_1714 (O_1714,N_15355,N_18102);
or UO_1715 (O_1715,N_19319,N_18469);
nand UO_1716 (O_1716,N_18457,N_16719);
nor UO_1717 (O_1717,N_15037,N_18877);
and UO_1718 (O_1718,N_16082,N_16981);
and UO_1719 (O_1719,N_17448,N_17863);
and UO_1720 (O_1720,N_17878,N_19846);
nand UO_1721 (O_1721,N_16944,N_19851);
nor UO_1722 (O_1722,N_16677,N_18691);
nand UO_1723 (O_1723,N_18285,N_18990);
nor UO_1724 (O_1724,N_16939,N_16089);
nor UO_1725 (O_1725,N_15808,N_19461);
nor UO_1726 (O_1726,N_15449,N_19497);
or UO_1727 (O_1727,N_19204,N_15940);
and UO_1728 (O_1728,N_15279,N_17589);
nand UO_1729 (O_1729,N_19088,N_15663);
xor UO_1730 (O_1730,N_19218,N_19732);
xnor UO_1731 (O_1731,N_16269,N_15579);
xor UO_1732 (O_1732,N_15938,N_17381);
and UO_1733 (O_1733,N_17581,N_17331);
nor UO_1734 (O_1734,N_17440,N_17555);
or UO_1735 (O_1735,N_16544,N_18109);
and UO_1736 (O_1736,N_19055,N_17396);
nor UO_1737 (O_1737,N_18554,N_16958);
xor UO_1738 (O_1738,N_16197,N_15963);
nor UO_1739 (O_1739,N_15108,N_16874);
nand UO_1740 (O_1740,N_15318,N_19212);
nand UO_1741 (O_1741,N_18313,N_16746);
nor UO_1742 (O_1742,N_15323,N_17512);
nand UO_1743 (O_1743,N_19796,N_18222);
or UO_1744 (O_1744,N_16111,N_18804);
nor UO_1745 (O_1745,N_19216,N_15854);
nor UO_1746 (O_1746,N_19361,N_17423);
and UO_1747 (O_1747,N_15244,N_16452);
and UO_1748 (O_1748,N_15389,N_19275);
or UO_1749 (O_1749,N_19293,N_15382);
nand UO_1750 (O_1750,N_18255,N_19010);
xor UO_1751 (O_1751,N_19605,N_19185);
or UO_1752 (O_1752,N_19999,N_15256);
or UO_1753 (O_1753,N_18866,N_18356);
or UO_1754 (O_1754,N_15365,N_18860);
nand UO_1755 (O_1755,N_19315,N_18017);
nor UO_1756 (O_1756,N_19384,N_17320);
or UO_1757 (O_1757,N_15032,N_17567);
and UO_1758 (O_1758,N_18371,N_19572);
or UO_1759 (O_1759,N_17533,N_17819);
nand UO_1760 (O_1760,N_15385,N_17714);
xor UO_1761 (O_1761,N_15946,N_18856);
nor UO_1762 (O_1762,N_19571,N_19985);
xnor UO_1763 (O_1763,N_18321,N_16422);
and UO_1764 (O_1764,N_18772,N_19137);
and UO_1765 (O_1765,N_17107,N_15715);
nand UO_1766 (O_1766,N_17951,N_15943);
nor UO_1767 (O_1767,N_15915,N_15173);
nor UO_1768 (O_1768,N_15662,N_15501);
nand UO_1769 (O_1769,N_18914,N_18679);
nor UO_1770 (O_1770,N_17369,N_19422);
nor UO_1771 (O_1771,N_18611,N_18283);
or UO_1772 (O_1772,N_15484,N_18707);
and UO_1773 (O_1773,N_16575,N_15228);
or UO_1774 (O_1774,N_16340,N_17843);
nor UO_1775 (O_1775,N_19746,N_15693);
nor UO_1776 (O_1776,N_16903,N_18645);
or UO_1777 (O_1777,N_18486,N_19146);
nand UO_1778 (O_1778,N_19627,N_19558);
xnor UO_1779 (O_1779,N_15000,N_16306);
or UO_1780 (O_1780,N_17664,N_19806);
or UO_1781 (O_1781,N_15011,N_17480);
nand UO_1782 (O_1782,N_18838,N_18218);
or UO_1783 (O_1783,N_15421,N_17762);
xor UO_1784 (O_1784,N_19775,N_15462);
xnor UO_1785 (O_1785,N_17459,N_19305);
nor UO_1786 (O_1786,N_15476,N_19586);
nor UO_1787 (O_1787,N_19278,N_19494);
nand UO_1788 (O_1788,N_16612,N_15010);
and UO_1789 (O_1789,N_18252,N_15689);
nand UO_1790 (O_1790,N_19223,N_19342);
or UO_1791 (O_1791,N_16516,N_16641);
nand UO_1792 (O_1792,N_15827,N_19463);
nand UO_1793 (O_1793,N_18935,N_19761);
nor UO_1794 (O_1794,N_19163,N_18246);
nand UO_1795 (O_1795,N_18103,N_15470);
or UO_1796 (O_1796,N_17608,N_17483);
or UO_1797 (O_1797,N_15497,N_16454);
and UO_1798 (O_1798,N_15645,N_17051);
nor UO_1799 (O_1799,N_15179,N_15145);
or UO_1800 (O_1800,N_15212,N_15804);
nor UO_1801 (O_1801,N_16927,N_19323);
nor UO_1802 (O_1802,N_15857,N_16363);
or UO_1803 (O_1803,N_19192,N_19353);
nor UO_1804 (O_1804,N_15633,N_19060);
or UO_1805 (O_1805,N_17460,N_17718);
and UO_1806 (O_1806,N_18164,N_18018);
nor UO_1807 (O_1807,N_18652,N_16521);
or UO_1808 (O_1808,N_17202,N_16658);
nand UO_1809 (O_1809,N_16015,N_19626);
and UO_1810 (O_1810,N_18026,N_19068);
and UO_1811 (O_1811,N_16008,N_16303);
nor UO_1812 (O_1812,N_15635,N_18574);
and UO_1813 (O_1813,N_17636,N_17969);
and UO_1814 (O_1814,N_18495,N_17587);
xor UO_1815 (O_1815,N_16467,N_18586);
nor UO_1816 (O_1816,N_18997,N_19832);
xnor UO_1817 (O_1817,N_17836,N_16145);
nand UO_1818 (O_1818,N_15337,N_15549);
or UO_1819 (O_1819,N_16964,N_16766);
and UO_1820 (O_1820,N_18173,N_19125);
or UO_1821 (O_1821,N_16935,N_18503);
xor UO_1822 (O_1822,N_16710,N_19950);
nand UO_1823 (O_1823,N_17336,N_16288);
nand UO_1824 (O_1824,N_17641,N_18709);
or UO_1825 (O_1825,N_16907,N_16486);
and UO_1826 (O_1826,N_16921,N_16776);
or UO_1827 (O_1827,N_15897,N_15299);
or UO_1828 (O_1828,N_17438,N_15073);
or UO_1829 (O_1829,N_18597,N_18996);
nand UO_1830 (O_1830,N_18505,N_15416);
or UO_1831 (O_1831,N_16556,N_18482);
nor UO_1832 (O_1832,N_18400,N_15625);
and UO_1833 (O_1833,N_15509,N_15122);
nor UO_1834 (O_1834,N_16570,N_18522);
nor UO_1835 (O_1835,N_15888,N_16224);
and UO_1836 (O_1836,N_19413,N_15181);
and UO_1837 (O_1837,N_16532,N_16632);
or UO_1838 (O_1838,N_18090,N_19363);
and UO_1839 (O_1839,N_19778,N_17467);
and UO_1840 (O_1840,N_19133,N_19312);
nand UO_1841 (O_1841,N_19340,N_17138);
nand UO_1842 (O_1842,N_18074,N_18637);
nor UO_1843 (O_1843,N_18214,N_15111);
xor UO_1844 (O_1844,N_17451,N_18846);
and UO_1845 (O_1845,N_16559,N_15997);
nand UO_1846 (O_1846,N_18437,N_15757);
nor UO_1847 (O_1847,N_18297,N_17598);
nand UO_1848 (O_1848,N_18338,N_16499);
or UO_1849 (O_1849,N_18167,N_18119);
nor UO_1850 (O_1850,N_18697,N_15852);
and UO_1851 (O_1851,N_19170,N_16513);
xor UO_1852 (O_1852,N_19755,N_15176);
nor UO_1853 (O_1853,N_15367,N_19510);
and UO_1854 (O_1854,N_19692,N_18902);
nor UO_1855 (O_1855,N_15942,N_15045);
or UO_1856 (O_1856,N_17337,N_16253);
or UO_1857 (O_1857,N_17316,N_17321);
or UO_1858 (O_1858,N_15364,N_19575);
nand UO_1859 (O_1859,N_15699,N_17542);
nor UO_1860 (O_1860,N_18084,N_15833);
nor UO_1861 (O_1861,N_15823,N_18324);
and UO_1862 (O_1862,N_15498,N_16704);
nor UO_1863 (O_1863,N_15119,N_16518);
nor UO_1864 (O_1864,N_19383,N_18547);
nor UO_1865 (O_1865,N_19454,N_17579);
xnor UO_1866 (O_1866,N_19714,N_19000);
nand UO_1867 (O_1867,N_18402,N_19581);
or UO_1868 (O_1868,N_16807,N_17490);
or UO_1869 (O_1869,N_16020,N_16811);
and UO_1870 (O_1870,N_17584,N_16502);
and UO_1871 (O_1871,N_17845,N_19504);
and UO_1872 (O_1872,N_19287,N_16541);
and UO_1873 (O_1873,N_18247,N_17546);
nand UO_1874 (O_1874,N_18502,N_16736);
or UO_1875 (O_1875,N_15949,N_18066);
nor UO_1876 (O_1876,N_17465,N_17850);
nand UO_1877 (O_1877,N_17596,N_18604);
and UO_1878 (O_1878,N_16805,N_16216);
nand UO_1879 (O_1879,N_17685,N_16972);
and UO_1880 (O_1880,N_15813,N_18823);
and UO_1881 (O_1881,N_19915,N_17167);
and UO_1882 (O_1882,N_17639,N_18585);
nor UO_1883 (O_1883,N_18372,N_15459);
nor UO_1884 (O_1884,N_19668,N_17056);
nand UO_1885 (O_1885,N_18000,N_15785);
nand UO_1886 (O_1886,N_15359,N_16367);
nand UO_1887 (O_1887,N_16517,N_18884);
or UO_1888 (O_1888,N_16676,N_17712);
nand UO_1889 (O_1889,N_19334,N_16341);
and UO_1890 (O_1890,N_18932,N_16141);
and UO_1891 (O_1891,N_15468,N_18335);
and UO_1892 (O_1892,N_18603,N_16469);
and UO_1893 (O_1893,N_16535,N_19814);
xnor UO_1894 (O_1894,N_19642,N_18816);
nand UO_1895 (O_1895,N_16450,N_17377);
nand UO_1896 (O_1896,N_18369,N_18425);
or UO_1897 (O_1897,N_17310,N_18169);
xor UO_1898 (O_1898,N_15797,N_16437);
and UO_1899 (O_1899,N_19316,N_15972);
or UO_1900 (O_1900,N_19064,N_17278);
nand UO_1901 (O_1901,N_19523,N_16835);
and UO_1902 (O_1902,N_15349,N_17775);
nand UO_1903 (O_1903,N_16298,N_19076);
and UO_1904 (O_1904,N_18773,N_19001);
and UO_1905 (O_1905,N_16045,N_19151);
nor UO_1906 (O_1906,N_16097,N_15424);
and UO_1907 (O_1907,N_15650,N_18957);
nor UO_1908 (O_1908,N_16539,N_17625);
nand UO_1909 (O_1909,N_15528,N_19920);
and UO_1910 (O_1910,N_19705,N_17721);
xnor UO_1911 (O_1911,N_15781,N_15485);
xnor UO_1912 (O_1912,N_19393,N_16221);
nor UO_1913 (O_1913,N_16420,N_19070);
nand UO_1914 (O_1914,N_17789,N_19576);
or UO_1915 (O_1915,N_18478,N_15070);
xnor UO_1916 (O_1916,N_18187,N_16748);
and UO_1917 (O_1917,N_15463,N_16917);
nand UO_1918 (O_1918,N_17970,N_15156);
or UO_1919 (O_1919,N_15626,N_19420);
or UO_1920 (O_1920,N_19757,N_16171);
xnor UO_1921 (O_1921,N_19066,N_19526);
xor UO_1922 (O_1922,N_17083,N_15386);
nand UO_1923 (O_1923,N_18815,N_17571);
nand UO_1924 (O_1924,N_17742,N_17543);
nand UO_1925 (O_1925,N_17216,N_15993);
and UO_1926 (O_1926,N_17830,N_15981);
and UO_1927 (O_1927,N_16595,N_18236);
or UO_1928 (O_1928,N_17834,N_17923);
or UO_1929 (O_1929,N_19119,N_18887);
or UO_1930 (O_1930,N_17604,N_17640);
nor UO_1931 (O_1931,N_15627,N_16151);
xor UO_1932 (O_1932,N_15465,N_17908);
and UO_1933 (O_1933,N_16046,N_19922);
nor UO_1934 (O_1934,N_17924,N_15732);
or UO_1935 (O_1935,N_19196,N_16415);
nand UO_1936 (O_1936,N_18852,N_15531);
nor UO_1937 (O_1937,N_16976,N_16809);
xor UO_1938 (O_1938,N_18786,N_17218);
nor UO_1939 (O_1939,N_19966,N_18251);
and UO_1940 (O_1940,N_15378,N_19981);
and UO_1941 (O_1941,N_16970,N_15713);
nor UO_1942 (O_1942,N_17350,N_18644);
and UO_1943 (O_1943,N_17082,N_15887);
or UO_1944 (O_1944,N_18403,N_19168);
or UO_1945 (O_1945,N_18510,N_16682);
nor UO_1946 (O_1946,N_19512,N_16593);
or UO_1947 (O_1947,N_17648,N_19244);
or UO_1948 (O_1948,N_16858,N_17220);
and UO_1949 (O_1949,N_17644,N_16660);
and UO_1950 (O_1950,N_19955,N_18421);
or UO_1951 (O_1951,N_19501,N_16991);
xnor UO_1952 (O_1952,N_19964,N_18113);
or UO_1953 (O_1953,N_19265,N_19779);
nor UO_1954 (O_1954,N_15215,N_16726);
nand UO_1955 (O_1955,N_16714,N_16481);
nor UO_1956 (O_1956,N_15138,N_16492);
nor UO_1957 (O_1957,N_18422,N_19259);
nor UO_1958 (O_1958,N_16208,N_19926);
and UO_1959 (O_1959,N_19517,N_19743);
nand UO_1960 (O_1960,N_17566,N_15043);
xnor UO_1961 (O_1961,N_19228,N_17894);
or UO_1962 (O_1962,N_15061,N_15022);
nand UO_1963 (O_1963,N_19067,N_18872);
and UO_1964 (O_1964,N_17662,N_16054);
nor UO_1965 (O_1965,N_17434,N_16900);
or UO_1966 (O_1966,N_19672,N_16124);
nand UO_1967 (O_1967,N_16441,N_19565);
or UO_1968 (O_1968,N_17470,N_16245);
or UO_1969 (O_1969,N_17228,N_15002);
and UO_1970 (O_1970,N_18813,N_18049);
and UO_1971 (O_1971,N_19767,N_15710);
nor UO_1972 (O_1972,N_18596,N_15357);
and UO_1973 (O_1973,N_15285,N_18580);
and UO_1974 (O_1974,N_16296,N_18035);
or UO_1975 (O_1975,N_16030,N_16214);
nor UO_1976 (O_1976,N_17285,N_15550);
nor UO_1977 (O_1977,N_19898,N_17214);
nor UO_1978 (O_1978,N_18401,N_17687);
or UO_1979 (O_1979,N_19533,N_15390);
nand UO_1980 (O_1980,N_15581,N_18413);
or UO_1981 (O_1981,N_16169,N_19914);
nand UO_1982 (O_1982,N_15358,N_18318);
and UO_1983 (O_1983,N_16370,N_17178);
and UO_1984 (O_1984,N_17469,N_16262);
or UO_1985 (O_1985,N_15817,N_17757);
or UO_1986 (O_1986,N_16627,N_16689);
nor UO_1987 (O_1987,N_19410,N_18089);
and UO_1988 (O_1988,N_18353,N_17737);
nand UO_1989 (O_1989,N_15107,N_18672);
or UO_1990 (O_1990,N_18828,N_18861);
nor UO_1991 (O_1991,N_19887,N_17389);
and UO_1992 (O_1992,N_17208,N_19918);
or UO_1993 (O_1993,N_18961,N_17309);
and UO_1994 (O_1994,N_16566,N_18295);
nor UO_1995 (O_1995,N_15283,N_18433);
and UO_1996 (O_1996,N_17118,N_17346);
nand UO_1997 (O_1997,N_18733,N_15392);
xnor UO_1998 (O_1998,N_17503,N_19049);
nor UO_1999 (O_1999,N_18831,N_17794);
and UO_2000 (O_2000,N_18397,N_16001);
nand UO_2001 (O_2001,N_19428,N_19237);
or UO_2002 (O_2002,N_19546,N_16797);
nand UO_2003 (O_2003,N_16870,N_15931);
nand UO_2004 (O_2004,N_17411,N_17098);
or UO_2005 (O_2005,N_19680,N_15845);
nor UO_2006 (O_2006,N_15750,N_16716);
nor UO_2007 (O_2007,N_15912,N_17121);
or UO_2008 (O_2008,N_15948,N_18199);
and UO_2009 (O_2009,N_15771,N_16319);
nand UO_2010 (O_2010,N_15533,N_19438);
nor UO_2011 (O_2011,N_16395,N_19248);
or UO_2012 (O_2012,N_18475,N_18825);
nor UO_2013 (O_2013,N_19809,N_15884);
nor UO_2014 (O_2014,N_19838,N_18464);
nand UO_2015 (O_2015,N_17158,N_19610);
nand UO_2016 (O_2016,N_18568,N_16029);
nand UO_2017 (O_2017,N_16529,N_19933);
nand UO_2018 (O_2018,N_19818,N_17955);
nand UO_2019 (O_2019,N_15266,N_16600);
nor UO_2020 (O_2020,N_18030,N_19486);
and UO_2021 (O_2021,N_16538,N_18646);
and UO_2022 (O_2022,N_15143,N_17128);
nor UO_2023 (O_2023,N_17524,N_17965);
and UO_2024 (O_2024,N_18744,N_17500);
nand UO_2025 (O_2025,N_15029,N_18865);
nor UO_2026 (O_2026,N_17518,N_18883);
or UO_2027 (O_2027,N_16740,N_18826);
nand UO_2028 (O_2028,N_18122,N_15775);
and UO_2029 (O_2029,N_17291,N_19802);
nor UO_2030 (O_2030,N_19415,N_17505);
or UO_2031 (O_2031,N_15883,N_19518);
nor UO_2032 (O_2032,N_16125,N_15765);
and UO_2033 (O_2033,N_17000,N_17116);
or UO_2034 (O_2034,N_17942,N_17987);
and UO_2035 (O_2035,N_19392,N_19941);
and UO_2036 (O_2036,N_19348,N_17236);
xor UO_2037 (O_2037,N_19542,N_15350);
nor UO_2038 (O_2038,N_15741,N_16774);
xor UO_2039 (O_2039,N_19289,N_19631);
nand UO_2040 (O_2040,N_17717,N_15098);
xor UO_2041 (O_2041,N_17788,N_18506);
or UO_2042 (O_2042,N_16431,N_16428);
xor UO_2043 (O_2043,N_17020,N_15559);
nand UO_2044 (O_2044,N_19593,N_17609);
xor UO_2045 (O_2045,N_18426,N_19215);
nand UO_2046 (O_2046,N_17323,N_17905);
nand UO_2047 (O_2047,N_17048,N_15920);
nor UO_2048 (O_2048,N_16674,N_15347);
nor UO_2049 (O_2049,N_17263,N_16842);
nand UO_2050 (O_2050,N_15835,N_19365);
or UO_2051 (O_2051,N_18500,N_17415);
nor UO_2052 (O_2052,N_15087,N_17043);
nor UO_2053 (O_2053,N_15779,N_15701);
and UO_2054 (O_2054,N_16754,N_18029);
or UO_2055 (O_2055,N_17194,N_16226);
nand UO_2056 (O_2056,N_17637,N_17007);
and UO_2057 (O_2057,N_19573,N_17019);
nand UO_2058 (O_2058,N_18782,N_17997);
nor UO_2059 (O_2059,N_17069,N_17846);
nand UO_2060 (O_2060,N_16177,N_19313);
nand UO_2061 (O_2061,N_17824,N_17209);
nor UO_2062 (O_2062,N_17528,N_15155);
nand UO_2063 (O_2063,N_15038,N_19760);
nor UO_2064 (O_2064,N_17296,N_18625);
nor UO_2065 (O_2065,N_18817,N_19580);
nand UO_2066 (O_2066,N_19222,N_15278);
or UO_2067 (O_2067,N_17290,N_16235);
and UO_2068 (O_2068,N_16068,N_17204);
nor UO_2069 (O_2069,N_15300,N_18907);
xnor UO_2070 (O_2070,N_16408,N_17027);
nand UO_2071 (O_2071,N_17028,N_17826);
xor UO_2072 (O_2072,N_16333,N_19596);
nor UO_2073 (O_2073,N_15594,N_17626);
nand UO_2074 (O_2074,N_18099,N_16734);
xnor UO_2075 (O_2075,N_18151,N_19082);
nand UO_2076 (O_2076,N_15206,N_19104);
and UO_2077 (O_2077,N_18434,N_18548);
nor UO_2078 (O_2078,N_16047,N_16947);
and UO_2079 (O_2079,N_19739,N_15758);
and UO_2080 (O_2080,N_15137,N_19568);
and UO_2081 (O_2081,N_15505,N_16724);
and UO_2082 (O_2082,N_19079,N_17539);
nor UO_2083 (O_2083,N_18789,N_17931);
and UO_2084 (O_2084,N_15062,N_19886);
nor UO_2085 (O_2085,N_16453,N_17420);
or UO_2086 (O_2086,N_19745,N_18333);
nor UO_2087 (O_2087,N_16574,N_15929);
xnor UO_2088 (O_2088,N_15873,N_15990);
or UO_2089 (O_2089,N_17437,N_18563);
nand UO_2090 (O_2090,N_16007,N_18149);
xnor UO_2091 (O_2091,N_17751,N_18417);
nor UO_2092 (O_2092,N_18976,N_18391);
and UO_2093 (O_2093,N_15925,N_19563);
nand UO_2094 (O_2094,N_19876,N_16862);
and UO_2095 (O_2095,N_16705,N_19557);
nor UO_2096 (O_2096,N_17113,N_17883);
and UO_2097 (O_2097,N_15209,N_16983);
nor UO_2098 (O_2098,N_19147,N_15298);
or UO_2099 (O_2099,N_19943,N_15399);
or UO_2100 (O_2100,N_16573,N_16414);
nor UO_2101 (O_2101,N_15004,N_18396);
or UO_2102 (O_2102,N_19379,N_17792);
and UO_2103 (O_2103,N_18583,N_17804);
xor UO_2104 (O_2104,N_16369,N_15863);
and UO_2105 (O_2105,N_15812,N_16720);
and UO_2106 (O_2106,N_15836,N_19026);
or UO_2107 (O_2107,N_16946,N_17921);
nand UO_2108 (O_2108,N_16106,N_16611);
nand UO_2109 (O_2109,N_19370,N_17032);
nand UO_2110 (O_2110,N_18690,N_15603);
or UO_2111 (O_2111,N_16002,N_18453);
nand UO_2112 (O_2112,N_15968,N_19429);
or UO_2113 (O_2113,N_17400,N_15236);
and UO_2114 (O_2114,N_18614,N_15066);
xor UO_2115 (O_2115,N_18525,N_17882);
nor UO_2116 (O_2116,N_18375,N_15620);
and UO_2117 (O_2117,N_19579,N_17553);
nand UO_2118 (O_2118,N_18699,N_19965);
xor UO_2119 (O_2119,N_18414,N_18191);
nand UO_2120 (O_2120,N_16195,N_17647);
nand UO_2121 (O_2121,N_17017,N_18655);
or UO_2122 (O_2122,N_18293,N_16780);
and UO_2123 (O_2123,N_16909,N_18670);
and UO_2124 (O_2124,N_17720,N_16759);
nor UO_2125 (O_2125,N_17281,N_15613);
nand UO_2126 (O_2126,N_16183,N_16198);
or UO_2127 (O_2127,N_17708,N_15560);
or UO_2128 (O_2128,N_19598,N_17455);
nor UO_2129 (O_2129,N_19770,N_15329);
xnor UO_2130 (O_2130,N_18979,N_15995);
nor UO_2131 (O_2131,N_18212,N_16990);
and UO_2132 (O_2132,N_17270,N_15003);
nand UO_2133 (O_2133,N_17520,N_16491);
nand UO_2134 (O_2134,N_16108,N_15674);
and UO_2135 (O_2135,N_16062,N_19690);
nor UO_2136 (O_2136,N_19471,N_19787);
and UO_2137 (O_2137,N_19469,N_17419);
nand UO_2138 (O_2138,N_17607,N_16779);
and UO_2139 (O_2139,N_16966,N_17088);
or UO_2140 (O_2140,N_19063,N_16255);
and UO_2141 (O_2141,N_16609,N_17822);
nand UO_2142 (O_2142,N_18841,N_19274);
nor UO_2143 (O_2143,N_15908,N_18962);
xnor UO_2144 (O_2144,N_19386,N_17700);
nor UO_2145 (O_2145,N_18085,N_16185);
nor UO_2146 (O_2146,N_18076,N_16523);
nor UO_2147 (O_2147,N_16568,N_18515);
or UO_2148 (O_2148,N_18016,N_17916);
nor UO_2149 (O_2149,N_15372,N_17259);
nand UO_2150 (O_2150,N_15658,N_16812);
or UO_2151 (O_2151,N_18770,N_17077);
nand UO_2152 (O_2152,N_19932,N_15832);
and UO_2153 (O_2153,N_18732,N_18867);
or UO_2154 (O_2154,N_18489,N_19210);
nand UO_2155 (O_2155,N_16511,N_19173);
or UO_2156 (O_2156,N_19678,N_15504);
or UO_2157 (O_2157,N_17666,N_19100);
nor UO_2158 (O_2158,N_17016,N_19322);
nand UO_2159 (O_2159,N_15793,N_16768);
and UO_2160 (O_2160,N_16122,N_19637);
and UO_2161 (O_2161,N_16998,N_16292);
or UO_2162 (O_2162,N_15708,N_15491);
nand UO_2163 (O_2163,N_16795,N_15602);
nand UO_2164 (O_2164,N_18131,N_19405);
nand UO_2165 (O_2165,N_16471,N_15351);
or UO_2166 (O_2166,N_16025,N_17561);
or UO_2167 (O_2167,N_18384,N_17341);
nand UO_2168 (O_2168,N_19235,N_18919);
or UO_2169 (O_2169,N_16154,N_18042);
nand UO_2170 (O_2170,N_16464,N_19947);
xnor UO_2171 (O_2171,N_19860,N_17054);
nand UO_2172 (O_2172,N_16801,N_18694);
xor UO_2173 (O_2173,N_18619,N_19130);
nand UO_2174 (O_2174,N_16260,N_17392);
nand UO_2175 (O_2175,N_16868,N_16985);
xor UO_2176 (O_2176,N_16648,N_18366);
and UO_2177 (O_2177,N_15799,N_19609);
nand UO_2178 (O_2178,N_17692,N_15831);
nor UO_2179 (O_2179,N_18731,N_16100);
nand UO_2180 (O_2180,N_19663,N_17140);
nand UO_2181 (O_2181,N_17783,N_17670);
xor UO_2182 (O_2182,N_19061,N_19967);
or UO_2183 (O_2183,N_17039,N_15047);
or UO_2184 (O_2184,N_16941,N_19172);
or UO_2185 (O_2185,N_19753,N_19813);
and UO_2186 (O_2186,N_17592,N_15803);
and UO_2187 (O_2187,N_18177,N_17047);
nand UO_2188 (O_2188,N_15984,N_15764);
nor UO_2189 (O_2189,N_19980,N_15928);
and UO_2190 (O_2190,N_15875,N_17136);
nor UO_2191 (O_2191,N_19513,N_19027);
or UO_2192 (O_2192,N_17993,N_17036);
nor UO_2193 (O_2193,N_19834,N_18767);
xor UO_2194 (O_2194,N_15722,N_19230);
and UO_2195 (O_2195,N_16919,N_18245);
xnor UO_2196 (O_2196,N_15876,N_15270);
nand UO_2197 (O_2197,N_17816,N_16892);
nand UO_2198 (O_2198,N_17810,N_19655);
nand UO_2199 (O_2199,N_17657,N_18088);
nand UO_2200 (O_2200,N_16936,N_16223);
xnor UO_2201 (O_2201,N_16973,N_15430);
or UO_2202 (O_2202,N_16252,N_16382);
and UO_2203 (O_2203,N_17669,N_19211);
and UO_2204 (O_2204,N_16349,N_15240);
or UO_2205 (O_2205,N_15369,N_16353);
and UO_2206 (O_2206,N_15790,N_17930);
nand UO_2207 (O_2207,N_19613,N_17322);
xnor UO_2208 (O_2208,N_18178,N_17472);
nand UO_2209 (O_2209,N_17620,N_15203);
or UO_2210 (O_2210,N_19135,N_17504);
and UO_2211 (O_2211,N_19758,N_18121);
or UO_2212 (O_2212,N_17690,N_17150);
nor UO_2213 (O_2213,N_18473,N_18764);
and UO_2214 (O_2214,N_17266,N_19483);
xnor UO_2215 (O_2215,N_17057,N_19729);
nand UO_2216 (O_2216,N_17085,N_17946);
xor UO_2217 (O_2217,N_15106,N_17401);
and UO_2218 (O_2218,N_15974,N_18171);
nand UO_2219 (O_2219,N_19332,N_18594);
and UO_2220 (O_2220,N_18718,N_18234);
or UO_2221 (O_2221,N_16313,N_15063);
and UO_2222 (O_2222,N_15428,N_17552);
nor UO_2223 (O_2223,N_15271,N_17429);
and UO_2224 (O_2224,N_19078,N_17765);
xnor UO_2225 (O_2225,N_18780,N_15169);
and UO_2226 (O_2226,N_17635,N_15933);
nand UO_2227 (O_2227,N_16951,N_16243);
nor UO_2228 (O_2228,N_15913,N_16442);
nand UO_2229 (O_2229,N_19762,N_18087);
nor UO_2230 (O_2230,N_18985,N_15124);
or UO_2231 (O_2231,N_19208,N_17348);
xnor UO_2232 (O_2232,N_15723,N_19556);
or UO_2233 (O_2233,N_16587,N_16968);
nand UO_2234 (O_2234,N_16394,N_15204);
nand UO_2235 (O_2235,N_16971,N_17076);
xor UO_2236 (O_2236,N_15805,N_18734);
nor UO_2237 (O_2237,N_16691,N_17093);
or UO_2238 (O_2238,N_17109,N_19404);
and UO_2239 (O_2239,N_19277,N_18685);
nand UO_2240 (O_2240,N_19776,N_18387);
or UO_2241 (O_2241,N_16501,N_18752);
or UO_2242 (O_2242,N_17104,N_18714);
and UO_2243 (O_2243,N_17727,N_18555);
nor UO_2244 (O_2244,N_17756,N_19816);
nand UO_2245 (O_2245,N_19331,N_16727);
nor UO_2246 (O_2246,N_19869,N_17785);
or UO_2247 (O_2247,N_19948,N_16839);
nand UO_2248 (O_2248,N_15864,N_16430);
nand UO_2249 (O_2249,N_15707,N_15254);
nor UO_2250 (O_2250,N_18559,N_17722);
or UO_2251 (O_2251,N_17588,N_17001);
and UO_2252 (O_2252,N_16213,N_16138);
or UO_2253 (O_2253,N_19835,N_15644);
or UO_2254 (O_2254,N_19726,N_19505);
or UO_2255 (O_2255,N_17564,N_18983);
nor UO_2256 (O_2256,N_15659,N_19229);
nor UO_2257 (O_2257,N_16999,N_16688);
and UO_2258 (O_2258,N_16984,N_16413);
nand UO_2259 (O_2259,N_18233,N_15193);
nor UO_2260 (O_2260,N_16520,N_15503);
nor UO_2261 (O_2261,N_15443,N_15282);
xor UO_2262 (O_2262,N_18938,N_15341);
nand UO_2263 (O_2263,N_18693,N_18449);
or UO_2264 (O_2264,N_15989,N_16155);
and UO_2265 (O_2265,N_15826,N_16458);
nand UO_2266 (O_2266,N_15333,N_15748);
or UO_2267 (O_2267,N_19114,N_18785);
nor UO_2268 (O_2268,N_16295,N_16834);
and UO_2269 (O_2269,N_18981,N_17583);
or UO_2270 (O_2270,N_16647,N_15810);
or UO_2271 (O_2271,N_17237,N_17405);
nor UO_2272 (O_2272,N_16833,N_15434);
or UO_2273 (O_2273,N_15383,N_15543);
or UO_2274 (O_2274,N_17074,N_16821);
and UO_2275 (O_2275,N_17610,N_19013);
nand UO_2276 (O_2276,N_19844,N_18073);
nor UO_2277 (O_2277,N_18829,N_15518);
and UO_2278 (O_2278,N_16184,N_17906);
and UO_2279 (O_2279,N_15441,N_15743);
xor UO_2280 (O_2280,N_18144,N_19801);
or UO_2281 (O_2281,N_17417,N_15162);
nor UO_2282 (O_2282,N_16898,N_17431);
and UO_2283 (O_2283,N_17343,N_18807);
or UO_2284 (O_2284,N_19283,N_15034);
nor UO_2285 (O_2285,N_16011,N_15609);
or UO_2286 (O_2286,N_15869,N_16675);
or UO_2287 (O_2287,N_15829,N_16132);
or UO_2288 (O_2288,N_15675,N_19009);
or UO_2289 (O_2289,N_19474,N_18334);
nand UO_2290 (O_2290,N_17375,N_19617);
nor UO_2291 (O_2291,N_18567,N_16356);
or UO_2292 (O_2292,N_18165,N_16602);
or UO_2293 (O_2293,N_18696,N_15322);
xor UO_2294 (O_2294,N_16194,N_16472);
nor UO_2295 (O_2295,N_19103,N_18216);
or UO_2296 (O_2296,N_16967,N_18992);
or UO_2297 (O_2297,N_18857,N_15539);
nand UO_2298 (O_2298,N_19140,N_19589);
or UO_2299 (O_2299,N_18239,N_15452);
nor UO_2300 (O_2300,N_17482,N_16072);
and UO_2301 (O_2301,N_15861,N_16191);
nor UO_2302 (O_2302,N_18882,N_18405);
nand UO_2303 (O_2303,N_16000,N_18602);
nor UO_2304 (O_2304,N_18374,N_18858);
and UO_2305 (O_2305,N_19992,N_19913);
or UO_2306 (O_2306,N_19872,N_17814);
or UO_2307 (O_2307,N_19186,N_15754);
or UO_2308 (O_2308,N_16033,N_15309);
xnor UO_2309 (O_2309,N_17629,N_19646);
or UO_2310 (O_2310,N_19465,N_16300);
nand UO_2311 (O_2311,N_17672,N_19364);
or UO_2312 (O_2312,N_19226,N_18200);
and UO_2313 (O_2313,N_18393,N_19930);
nor UO_2314 (O_2314,N_16711,N_17454);
nand UO_2315 (O_2315,N_16396,N_17844);
or UO_2316 (O_2316,N_17499,N_17166);
nor UO_2317 (O_2317,N_16254,N_17229);
nand UO_2318 (O_2318,N_15961,N_16897);
nor UO_2319 (O_2319,N_19181,N_15996);
xor UO_2320 (O_2320,N_19276,N_18765);
nand UO_2321 (O_2321,N_15746,N_18787);
and UO_2322 (O_2322,N_19371,N_16620);
xor UO_2323 (O_2323,N_15103,N_16969);
xor UO_2324 (O_2324,N_18305,N_16888);
and UO_2325 (O_2325,N_15496,N_15099);
nand UO_2326 (O_2326,N_17617,N_15482);
nor UO_2327 (O_2327,N_18279,N_15059);
or UO_2328 (O_2328,N_16076,N_18325);
nand UO_2329 (O_2329,N_16819,N_16530);
or UO_2330 (O_2330,N_18777,N_19677);
and UO_2331 (O_2331,N_17154,N_15320);
nand UO_2332 (O_2332,N_16979,N_17711);
xor UO_2333 (O_2333,N_18068,N_18796);
and UO_2334 (O_2334,N_17254,N_18215);
nor UO_2335 (O_2335,N_15229,N_18845);
and UO_2336 (O_2336,N_15410,N_19157);
nand UO_2337 (O_2337,N_17570,N_15191);
nand UO_2338 (O_2338,N_16723,N_16404);
xnor UO_2339 (O_2339,N_15521,N_19014);
nor UO_2340 (O_2340,N_15872,N_16293);
and UO_2341 (O_2341,N_17932,N_19270);
nand UO_2342 (O_2342,N_17642,N_18082);
nor UO_2343 (O_2343,N_16614,N_19977);
or UO_2344 (O_2344,N_15691,N_19462);
nor UO_2345 (O_2345,N_19301,N_16709);
nand UO_2346 (O_2346,N_15874,N_15168);
nand UO_2347 (O_2347,N_16192,N_17981);
nand UO_2348 (O_2348,N_19962,N_19085);
nand UO_2349 (O_2349,N_16337,N_19115);
nand UO_2350 (O_2350,N_18669,N_17778);
nand UO_2351 (O_2351,N_18768,N_16722);
nand UO_2352 (O_2352,N_17945,N_18931);
nand UO_2353 (O_2353,N_15904,N_16576);
nor UO_2354 (O_2354,N_18415,N_16094);
nor UO_2355 (O_2355,N_18947,N_19296);
or UO_2356 (O_2356,N_18227,N_17456);
or UO_2357 (O_2357,N_18019,N_19459);
xnor UO_2358 (O_2358,N_18363,N_18129);
nand UO_2359 (O_2359,N_18329,N_19327);
xor UO_2360 (O_2360,N_16081,N_18023);
and UO_2361 (O_2361,N_15146,N_17449);
or UO_2362 (O_2362,N_18459,N_19681);
and UO_2363 (O_2363,N_16336,N_17313);
and UO_2364 (O_2364,N_17654,N_15556);
xor UO_2365 (O_2365,N_18695,N_19096);
nand UO_2366 (O_2366,N_17475,N_15665);
nand UO_2367 (O_2367,N_18435,N_19683);
nor UO_2368 (O_2368,N_16659,N_18186);
and UO_2369 (O_2369,N_18377,N_19169);
and UO_2370 (O_2370,N_19403,N_15301);
or UO_2371 (O_2371,N_19271,N_18332);
nand UO_2372 (O_2372,N_19431,N_17772);
nand UO_2373 (O_2373,N_15197,N_16067);
xor UO_2374 (O_2374,N_16733,N_15006);
nand UO_2375 (O_2375,N_16470,N_18041);
nand UO_2376 (O_2376,N_19507,N_18995);
and UO_2377 (O_2377,N_17750,N_19983);
nand UO_2378 (O_2378,N_16012,N_15621);
or UO_2379 (O_2379,N_18208,N_16320);
or UO_2380 (O_2380,N_18479,N_19972);
or UO_2381 (O_2381,N_18323,N_18319);
xnor UO_2382 (O_2382,N_16945,N_17573);
or UO_2383 (O_2383,N_17206,N_19885);
or UO_2384 (O_2384,N_17319,N_15148);
nor UO_2385 (O_2385,N_17704,N_17284);
nor UO_2386 (O_2386,N_18238,N_17112);
and UO_2387 (O_2387,N_15590,N_16605);
nor UO_2388 (O_2388,N_18037,N_15934);
and UO_2389 (O_2389,N_19741,N_19870);
xnor UO_2390 (O_2390,N_15894,N_18407);
or UO_2391 (O_2391,N_15136,N_15597);
nor UO_2392 (O_2392,N_18837,N_15932);
nand UO_2393 (O_2393,N_19099,N_16899);
nand UO_2394 (O_2394,N_16433,N_15304);
xnor UO_2395 (O_2395,N_16234,N_15522);
nand UO_2396 (O_2396,N_15844,N_19232);
nor UO_2397 (O_2397,N_15983,N_17476);
nand UO_2398 (O_2398,N_16533,N_19768);
and UO_2399 (O_2399,N_18185,N_19652);
or UO_2400 (O_2400,N_19574,N_19674);
and UO_2401 (O_2401,N_19307,N_17913);
or UO_2402 (O_2402,N_19179,N_16592);
or UO_2403 (O_2403,N_18288,N_19734);
xor UO_2404 (O_2404,N_19804,N_18820);
and UO_2405 (O_2405,N_17234,N_18098);
nand UO_2406 (O_2406,N_16038,N_15157);
xnor UO_2407 (O_2407,N_18700,N_16906);
or UO_2408 (O_2408,N_15035,N_15095);
nor UO_2409 (O_2409,N_17773,N_15744);
xnor UO_2410 (O_2410,N_18562,N_18006);
and UO_2411 (O_2411,N_17102,N_17986);
xnor UO_2412 (O_2412,N_17562,N_19238);
or UO_2413 (O_2413,N_16425,N_17813);
nand UO_2414 (O_2414,N_16549,N_15439);
nor UO_2415 (O_2415,N_16633,N_15088);
and UO_2416 (O_2416,N_19561,N_18769);
nor UO_2417 (O_2417,N_16143,N_15907);
and UO_2418 (O_2418,N_19906,N_19165);
nand UO_2419 (O_2419,N_15921,N_18671);
nand UO_2420 (O_2420,N_16342,N_17197);
or UO_2421 (O_2421,N_18483,N_19451);
nor UO_2422 (O_2422,N_17578,N_19756);
nor UO_2423 (O_2423,N_18827,N_17335);
and UO_2424 (O_2424,N_16476,N_19144);
nor UO_2425 (O_2425,N_15514,N_15471);
and UO_2426 (O_2426,N_16014,N_16190);
and UO_2427 (O_2427,N_15001,N_18918);
and UO_2428 (O_2428,N_15142,N_15015);
or UO_2429 (O_2429,N_15442,N_17918);
or UO_2430 (O_2430,N_16584,N_16131);
xor UO_2431 (O_2431,N_18195,N_19018);
or UO_2432 (O_2432,N_16488,N_17611);
nor UO_2433 (O_2433,N_15277,N_18450);
nand UO_2434 (O_2434,N_18440,N_17898);
nand UO_2435 (O_2435,N_16310,N_17522);
nand UO_2436 (O_2436,N_18292,N_18241);
or UO_2437 (O_2437,N_18543,N_15286);
or UO_2438 (O_2438,N_19634,N_19285);
nor UO_2439 (O_2439,N_15483,N_17397);
nand UO_2440 (O_2440,N_15126,N_16799);
and UO_2441 (O_2441,N_17795,N_16948);
xnor UO_2442 (O_2442,N_18648,N_18894);
and UO_2443 (O_2443,N_15221,N_17817);
nand UO_2444 (O_2444,N_15769,N_16127);
and UO_2445 (O_2445,N_15737,N_15575);
and UO_2446 (O_2446,N_18354,N_17536);
nand UO_2447 (O_2447,N_16912,N_15219);
nor UO_2448 (O_2448,N_15153,N_18572);
or UO_2449 (O_2449,N_19113,N_18739);
xor UO_2450 (O_2450,N_16598,N_19093);
nor UO_2451 (O_2451,N_17994,N_15721);
and UO_2452 (O_2452,N_16447,N_16545);
nor UO_2453 (O_2453,N_15097,N_19687);
and UO_2454 (O_2454,N_16925,N_17699);
or UO_2455 (O_2455,N_17864,N_16943);
and UO_2456 (O_2456,N_15703,N_16982);
nand UO_2457 (O_2457,N_17653,N_15903);
or UO_2458 (O_2458,N_16742,N_19954);
or UO_2459 (O_2459,N_15641,N_18243);
or UO_2460 (O_2460,N_15652,N_18441);
or UO_2461 (O_2461,N_19310,N_18982);
and UO_2462 (O_2462,N_15851,N_17973);
and UO_2463 (O_2463,N_19570,N_15133);
and UO_2464 (O_2464,N_17473,N_18893);
nand UO_2465 (O_2465,N_16091,N_17084);
nand UO_2466 (O_2466,N_16678,N_19446);
nor UO_2467 (O_2467,N_16937,N_19938);
nor UO_2468 (O_2468,N_18839,N_19697);
or UO_2469 (O_2469,N_16329,N_15774);
and UO_2470 (O_2470,N_19625,N_15530);
or UO_2471 (O_2471,N_15973,N_15967);
nand UO_2472 (O_2472,N_16860,N_16908);
or UO_2473 (O_2473,N_18758,N_18488);
or UO_2474 (O_2474,N_17683,N_15676);
or UO_2475 (O_2475,N_16004,N_15150);
nor UO_2476 (O_2476,N_18801,N_19184);
and UO_2477 (O_2477,N_15290,N_19856);
nor UO_2478 (O_2478,N_18859,N_19020);
and UO_2479 (O_2479,N_19183,N_15611);
and UO_2480 (O_2480,N_19973,N_17485);
nand UO_2481 (O_2481,N_17304,N_18394);
xnor UO_2482 (O_2482,N_19435,N_16302);
nand UO_2483 (O_2483,N_15393,N_19072);
or UO_2484 (O_2484,N_19606,N_15686);
nor UO_2485 (O_2485,N_17974,N_19520);
and UO_2486 (O_2486,N_17300,N_16362);
or UO_2487 (O_2487,N_16165,N_16728);
nand UO_2488 (O_2488,N_15250,N_15054);
nand UO_2489 (O_2489,N_17408,N_19012);
nand UO_2490 (O_2490,N_16702,N_19694);
nand UO_2491 (O_2491,N_16715,N_18287);
or UO_2492 (O_2492,N_16725,N_19073);
and UO_2493 (O_2493,N_18512,N_15811);
and UO_2494 (O_2494,N_19426,N_17018);
and UO_2495 (O_2495,N_15325,N_17904);
and UO_2496 (O_2496,N_18738,N_18776);
nand UO_2497 (O_2497,N_16640,N_15311);
nor UO_2498 (O_2498,N_15583,N_16901);
and UO_2499 (O_2499,N_18822,N_19047);
endmodule